

module top
(
  data_i,
  sel_i,
  data_o
);

  input [8191:0] data_i;
  input [5:0] sel_i;
  output [8191:0] data_o;

  bsg_mux_butterfly
  wrapper
  (
    .data_i(data_i),
    .sel_i(sel_i),
    .data_o(data_o)
  );


endmodule



module bsg_swap_width_p128
(
  data_i,
  swap_i,
  data_o
);

  input [255:0] data_i;
  output [255:0] data_o;
  input swap_i;
  wire [255:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[127:0], data_i[255:128] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p256
(
  data_i,
  swap_i,
  data_o
);

  input [511:0] data_i;
  output [511:0] data_o;
  input swap_i;
  wire [511:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[255:0], data_i[511:256] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p512
(
  data_i,
  swap_i,
  data_o
);

  input [1023:0] data_i;
  output [1023:0] data_o;
  input swap_i;
  wire [1023:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[511:0], data_i[1023:512] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p1024
(
  data_i,
  swap_i,
  data_o
);

  input [2047:0] data_i;
  output [2047:0] data_o;
  input swap_i;
  wire [2047:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[1023:0], data_i[2047:1024] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p2048
(
  data_i,
  swap_i,
  data_o
);

  input [4095:0] data_i;
  output [4095:0] data_o;
  input swap_i;
  wire [4095:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[2047:0], data_i[4095:2048] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p4096
(
  data_i,
  swap_i,
  data_o
);

  input [8191:0] data_i;
  output [8191:0] data_o;
  input swap_i;
  wire [8191:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[4095:0], data_i[8191:4096] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_mux_butterfly
(
  data_i,
  sel_i,
  data_o
);

  input [8191:0] data_i;
  input [5:0] sel_i;
  output [8191:0] data_o;
  wire [8191:0] data_o;
  wire data_stage_1__8191_,data_stage_1__8190_,data_stage_1__8189_,data_stage_1__8188_,
  data_stage_1__8187_,data_stage_1__8186_,data_stage_1__8185_,data_stage_1__8184_,
  data_stage_1__8183_,data_stage_1__8182_,data_stage_1__8181_,data_stage_1__8180_,
  data_stage_1__8179_,data_stage_1__8178_,data_stage_1__8177_,data_stage_1__8176_,
  data_stage_1__8175_,data_stage_1__8174_,data_stage_1__8173_,data_stage_1__8172_,
  data_stage_1__8171_,data_stage_1__8170_,data_stage_1__8169_,data_stage_1__8168_,
  data_stage_1__8167_,data_stage_1__8166_,data_stage_1__8165_,data_stage_1__8164_,
  data_stage_1__8163_,data_stage_1__8162_,data_stage_1__8161_,data_stage_1__8160_,
  data_stage_1__8159_,data_stage_1__8158_,data_stage_1__8157_,data_stage_1__8156_,
  data_stage_1__8155_,data_stage_1__8154_,data_stage_1__8153_,data_stage_1__8152_,
  data_stage_1__8151_,data_stage_1__8150_,data_stage_1__8149_,data_stage_1__8148_,
  data_stage_1__8147_,data_stage_1__8146_,data_stage_1__8145_,data_stage_1__8144_,
  data_stage_1__8143_,data_stage_1__8142_,data_stage_1__8141_,data_stage_1__8140_,
  data_stage_1__8139_,data_stage_1__8138_,data_stage_1__8137_,data_stage_1__8136_,
  data_stage_1__8135_,data_stage_1__8134_,data_stage_1__8133_,data_stage_1__8132_,
  data_stage_1__8131_,data_stage_1__8130_,data_stage_1__8129_,data_stage_1__8128_,
  data_stage_1__8127_,data_stage_1__8126_,data_stage_1__8125_,data_stage_1__8124_,
  data_stage_1__8123_,data_stage_1__8122_,data_stage_1__8121_,data_stage_1__8120_,
  data_stage_1__8119_,data_stage_1__8118_,data_stage_1__8117_,data_stage_1__8116_,
  data_stage_1__8115_,data_stage_1__8114_,data_stage_1__8113_,data_stage_1__8112_,
  data_stage_1__8111_,data_stage_1__8110_,data_stage_1__8109_,data_stage_1__8108_,
  data_stage_1__8107_,data_stage_1__8106_,data_stage_1__8105_,data_stage_1__8104_,
  data_stage_1__8103_,data_stage_1__8102_,data_stage_1__8101_,data_stage_1__8100_,
  data_stage_1__8099_,data_stage_1__8098_,data_stage_1__8097_,data_stage_1__8096_,
  data_stage_1__8095_,data_stage_1__8094_,data_stage_1__8093_,data_stage_1__8092_,
  data_stage_1__8091_,data_stage_1__8090_,data_stage_1__8089_,data_stage_1__8088_,
  data_stage_1__8087_,data_stage_1__8086_,data_stage_1__8085_,data_stage_1__8084_,
  data_stage_1__8083_,data_stage_1__8082_,data_stage_1__8081_,data_stage_1__8080_,
  data_stage_1__8079_,data_stage_1__8078_,data_stage_1__8077_,data_stage_1__8076_,
  data_stage_1__8075_,data_stage_1__8074_,data_stage_1__8073_,data_stage_1__8072_,
  data_stage_1__8071_,data_stage_1__8070_,data_stage_1__8069_,data_stage_1__8068_,
  data_stage_1__8067_,data_stage_1__8066_,data_stage_1__8065_,data_stage_1__8064_,
  data_stage_1__8063_,data_stage_1__8062_,data_stage_1__8061_,data_stage_1__8060_,
  data_stage_1__8059_,data_stage_1__8058_,data_stage_1__8057_,data_stage_1__8056_,
  data_stage_1__8055_,data_stage_1__8054_,data_stage_1__8053_,data_stage_1__8052_,
  data_stage_1__8051_,data_stage_1__8050_,data_stage_1__8049_,data_stage_1__8048_,
  data_stage_1__8047_,data_stage_1__8046_,data_stage_1__8045_,data_stage_1__8044_,
  data_stage_1__8043_,data_stage_1__8042_,data_stage_1__8041_,data_stage_1__8040_,
  data_stage_1__8039_,data_stage_1__8038_,data_stage_1__8037_,data_stage_1__8036_,
  data_stage_1__8035_,data_stage_1__8034_,data_stage_1__8033_,data_stage_1__8032_,
  data_stage_1__8031_,data_stage_1__8030_,data_stage_1__8029_,data_stage_1__8028_,
  data_stage_1__8027_,data_stage_1__8026_,data_stage_1__8025_,data_stage_1__8024_,
  data_stage_1__8023_,data_stage_1__8022_,data_stage_1__8021_,data_stage_1__8020_,
  data_stage_1__8019_,data_stage_1__8018_,data_stage_1__8017_,data_stage_1__8016_,
  data_stage_1__8015_,data_stage_1__8014_,data_stage_1__8013_,data_stage_1__8012_,
  data_stage_1__8011_,data_stage_1__8010_,data_stage_1__8009_,data_stage_1__8008_,
  data_stage_1__8007_,data_stage_1__8006_,data_stage_1__8005_,data_stage_1__8004_,
  data_stage_1__8003_,data_stage_1__8002_,data_stage_1__8001_,data_stage_1__8000_,
  data_stage_1__7999_,data_stage_1__7998_,data_stage_1__7997_,data_stage_1__7996_,
  data_stage_1__7995_,data_stage_1__7994_,data_stage_1__7993_,data_stage_1__7992_,
  data_stage_1__7991_,data_stage_1__7990_,data_stage_1__7989_,data_stage_1__7988_,
  data_stage_1__7987_,data_stage_1__7986_,data_stage_1__7985_,data_stage_1__7984_,
  data_stage_1__7983_,data_stage_1__7982_,data_stage_1__7981_,data_stage_1__7980_,
  data_stage_1__7979_,data_stage_1__7978_,data_stage_1__7977_,data_stage_1__7976_,
  data_stage_1__7975_,data_stage_1__7974_,data_stage_1__7973_,data_stage_1__7972_,
  data_stage_1__7971_,data_stage_1__7970_,data_stage_1__7969_,data_stage_1__7968_,
  data_stage_1__7967_,data_stage_1__7966_,data_stage_1__7965_,data_stage_1__7964_,
  data_stage_1__7963_,data_stage_1__7962_,data_stage_1__7961_,data_stage_1__7960_,
  data_stage_1__7959_,data_stage_1__7958_,data_stage_1__7957_,data_stage_1__7956_,
  data_stage_1__7955_,data_stage_1__7954_,data_stage_1__7953_,data_stage_1__7952_,
  data_stage_1__7951_,data_stage_1__7950_,data_stage_1__7949_,data_stage_1__7948_,
  data_stage_1__7947_,data_stage_1__7946_,data_stage_1__7945_,data_stage_1__7944_,
  data_stage_1__7943_,data_stage_1__7942_,data_stage_1__7941_,data_stage_1__7940_,
  data_stage_1__7939_,data_stage_1__7938_,data_stage_1__7937_,data_stage_1__7936_,
  data_stage_1__7935_,data_stage_1__7934_,data_stage_1__7933_,data_stage_1__7932_,
  data_stage_1__7931_,data_stage_1__7930_,data_stage_1__7929_,data_stage_1__7928_,
  data_stage_1__7927_,data_stage_1__7926_,data_stage_1__7925_,data_stage_1__7924_,
  data_stage_1__7923_,data_stage_1__7922_,data_stage_1__7921_,data_stage_1__7920_,
  data_stage_1__7919_,data_stage_1__7918_,data_stage_1__7917_,data_stage_1__7916_,
  data_stage_1__7915_,data_stage_1__7914_,data_stage_1__7913_,data_stage_1__7912_,
  data_stage_1__7911_,data_stage_1__7910_,data_stage_1__7909_,data_stage_1__7908_,
  data_stage_1__7907_,data_stage_1__7906_,data_stage_1__7905_,data_stage_1__7904_,
  data_stage_1__7903_,data_stage_1__7902_,data_stage_1__7901_,data_stage_1__7900_,
  data_stage_1__7899_,data_stage_1__7898_,data_stage_1__7897_,data_stage_1__7896_,
  data_stage_1__7895_,data_stage_1__7894_,data_stage_1__7893_,data_stage_1__7892_,
  data_stage_1__7891_,data_stage_1__7890_,data_stage_1__7889_,data_stage_1__7888_,
  data_stage_1__7887_,data_stage_1__7886_,data_stage_1__7885_,data_stage_1__7884_,
  data_stage_1__7883_,data_stage_1__7882_,data_stage_1__7881_,data_stage_1__7880_,
  data_stage_1__7879_,data_stage_1__7878_,data_stage_1__7877_,data_stage_1__7876_,
  data_stage_1__7875_,data_stage_1__7874_,data_stage_1__7873_,data_stage_1__7872_,
  data_stage_1__7871_,data_stage_1__7870_,data_stage_1__7869_,data_stage_1__7868_,
  data_stage_1__7867_,data_stage_1__7866_,data_stage_1__7865_,data_stage_1__7864_,
  data_stage_1__7863_,data_stage_1__7862_,data_stage_1__7861_,data_stage_1__7860_,
  data_stage_1__7859_,data_stage_1__7858_,data_stage_1__7857_,data_stage_1__7856_,
  data_stage_1__7855_,data_stage_1__7854_,data_stage_1__7853_,data_stage_1__7852_,
  data_stage_1__7851_,data_stage_1__7850_,data_stage_1__7849_,data_stage_1__7848_,
  data_stage_1__7847_,data_stage_1__7846_,data_stage_1__7845_,data_stage_1__7844_,
  data_stage_1__7843_,data_stage_1__7842_,data_stage_1__7841_,data_stage_1__7840_,
  data_stage_1__7839_,data_stage_1__7838_,data_stage_1__7837_,data_stage_1__7836_,
  data_stage_1__7835_,data_stage_1__7834_,data_stage_1__7833_,data_stage_1__7832_,
  data_stage_1__7831_,data_stage_1__7830_,data_stage_1__7829_,data_stage_1__7828_,
  data_stage_1__7827_,data_stage_1__7826_,data_stage_1__7825_,data_stage_1__7824_,
  data_stage_1__7823_,data_stage_1__7822_,data_stage_1__7821_,data_stage_1__7820_,
  data_stage_1__7819_,data_stage_1__7818_,data_stage_1__7817_,data_stage_1__7816_,
  data_stage_1__7815_,data_stage_1__7814_,data_stage_1__7813_,data_stage_1__7812_,
  data_stage_1__7811_,data_stage_1__7810_,data_stage_1__7809_,data_stage_1__7808_,
  data_stage_1__7807_,data_stage_1__7806_,data_stage_1__7805_,data_stage_1__7804_,
  data_stage_1__7803_,data_stage_1__7802_,data_stage_1__7801_,data_stage_1__7800_,
  data_stage_1__7799_,data_stage_1__7798_,data_stage_1__7797_,data_stage_1__7796_,
  data_stage_1__7795_,data_stage_1__7794_,data_stage_1__7793_,data_stage_1__7792_,
  data_stage_1__7791_,data_stage_1__7790_,data_stage_1__7789_,data_stage_1__7788_,
  data_stage_1__7787_,data_stage_1__7786_,data_stage_1__7785_,data_stage_1__7784_,
  data_stage_1__7783_,data_stage_1__7782_,data_stage_1__7781_,data_stage_1__7780_,
  data_stage_1__7779_,data_stage_1__7778_,data_stage_1__7777_,data_stage_1__7776_,
  data_stage_1__7775_,data_stage_1__7774_,data_stage_1__7773_,data_stage_1__7772_,
  data_stage_1__7771_,data_stage_1__7770_,data_stage_1__7769_,data_stage_1__7768_,
  data_stage_1__7767_,data_stage_1__7766_,data_stage_1__7765_,data_stage_1__7764_,
  data_stage_1__7763_,data_stage_1__7762_,data_stage_1__7761_,data_stage_1__7760_,
  data_stage_1__7759_,data_stage_1__7758_,data_stage_1__7757_,data_stage_1__7756_,
  data_stage_1__7755_,data_stage_1__7754_,data_stage_1__7753_,data_stage_1__7752_,
  data_stage_1__7751_,data_stage_1__7750_,data_stage_1__7749_,data_stage_1__7748_,
  data_stage_1__7747_,data_stage_1__7746_,data_stage_1__7745_,data_stage_1__7744_,
  data_stage_1__7743_,data_stage_1__7742_,data_stage_1__7741_,data_stage_1__7740_,
  data_stage_1__7739_,data_stage_1__7738_,data_stage_1__7737_,data_stage_1__7736_,
  data_stage_1__7735_,data_stage_1__7734_,data_stage_1__7733_,data_stage_1__7732_,
  data_stage_1__7731_,data_stage_1__7730_,data_stage_1__7729_,data_stage_1__7728_,
  data_stage_1__7727_,data_stage_1__7726_,data_stage_1__7725_,data_stage_1__7724_,
  data_stage_1__7723_,data_stage_1__7722_,data_stage_1__7721_,data_stage_1__7720_,
  data_stage_1__7719_,data_stage_1__7718_,data_stage_1__7717_,data_stage_1__7716_,
  data_stage_1__7715_,data_stage_1__7714_,data_stage_1__7713_,data_stage_1__7712_,
  data_stage_1__7711_,data_stage_1__7710_,data_stage_1__7709_,data_stage_1__7708_,
  data_stage_1__7707_,data_stage_1__7706_,data_stage_1__7705_,data_stage_1__7704_,
  data_stage_1__7703_,data_stage_1__7702_,data_stage_1__7701_,data_stage_1__7700_,
  data_stage_1__7699_,data_stage_1__7698_,data_stage_1__7697_,data_stage_1__7696_,
  data_stage_1__7695_,data_stage_1__7694_,data_stage_1__7693_,data_stage_1__7692_,
  data_stage_1__7691_,data_stage_1__7690_,data_stage_1__7689_,data_stage_1__7688_,
  data_stage_1__7687_,data_stage_1__7686_,data_stage_1__7685_,data_stage_1__7684_,
  data_stage_1__7683_,data_stage_1__7682_,data_stage_1__7681_,data_stage_1__7680_,
  data_stage_1__7679_,data_stage_1__7678_,data_stage_1__7677_,data_stage_1__7676_,
  data_stage_1__7675_,data_stage_1__7674_,data_stage_1__7673_,data_stage_1__7672_,
  data_stage_1__7671_,data_stage_1__7670_,data_stage_1__7669_,data_stage_1__7668_,
  data_stage_1__7667_,data_stage_1__7666_,data_stage_1__7665_,data_stage_1__7664_,
  data_stage_1__7663_,data_stage_1__7662_,data_stage_1__7661_,data_stage_1__7660_,
  data_stage_1__7659_,data_stage_1__7658_,data_stage_1__7657_,data_stage_1__7656_,
  data_stage_1__7655_,data_stage_1__7654_,data_stage_1__7653_,data_stage_1__7652_,
  data_stage_1__7651_,data_stage_1__7650_,data_stage_1__7649_,data_stage_1__7648_,
  data_stage_1__7647_,data_stage_1__7646_,data_stage_1__7645_,data_stage_1__7644_,
  data_stage_1__7643_,data_stage_1__7642_,data_stage_1__7641_,data_stage_1__7640_,
  data_stage_1__7639_,data_stage_1__7638_,data_stage_1__7637_,data_stage_1__7636_,
  data_stage_1__7635_,data_stage_1__7634_,data_stage_1__7633_,data_stage_1__7632_,
  data_stage_1__7631_,data_stage_1__7630_,data_stage_1__7629_,data_stage_1__7628_,
  data_stage_1__7627_,data_stage_1__7626_,data_stage_1__7625_,data_stage_1__7624_,
  data_stage_1__7623_,data_stage_1__7622_,data_stage_1__7621_,data_stage_1__7620_,
  data_stage_1__7619_,data_stage_1__7618_,data_stage_1__7617_,data_stage_1__7616_,
  data_stage_1__7615_,data_stage_1__7614_,data_stage_1__7613_,data_stage_1__7612_,
  data_stage_1__7611_,data_stage_1__7610_,data_stage_1__7609_,data_stage_1__7608_,
  data_stage_1__7607_,data_stage_1__7606_,data_stage_1__7605_,data_stage_1__7604_,
  data_stage_1__7603_,data_stage_1__7602_,data_stage_1__7601_,data_stage_1__7600_,
  data_stage_1__7599_,data_stage_1__7598_,data_stage_1__7597_,data_stage_1__7596_,
  data_stage_1__7595_,data_stage_1__7594_,data_stage_1__7593_,data_stage_1__7592_,
  data_stage_1__7591_,data_stage_1__7590_,data_stage_1__7589_,data_stage_1__7588_,
  data_stage_1__7587_,data_stage_1__7586_,data_stage_1__7585_,data_stage_1__7584_,
  data_stage_1__7583_,data_stage_1__7582_,data_stage_1__7581_,data_stage_1__7580_,
  data_stage_1__7579_,data_stage_1__7578_,data_stage_1__7577_,data_stage_1__7576_,
  data_stage_1__7575_,data_stage_1__7574_,data_stage_1__7573_,data_stage_1__7572_,
  data_stage_1__7571_,data_stage_1__7570_,data_stage_1__7569_,data_stage_1__7568_,
  data_stage_1__7567_,data_stage_1__7566_,data_stage_1__7565_,data_stage_1__7564_,
  data_stage_1__7563_,data_stage_1__7562_,data_stage_1__7561_,data_stage_1__7560_,
  data_stage_1__7559_,data_stage_1__7558_,data_stage_1__7557_,data_stage_1__7556_,
  data_stage_1__7555_,data_stage_1__7554_,data_stage_1__7553_,data_stage_1__7552_,
  data_stage_1__7551_,data_stage_1__7550_,data_stage_1__7549_,data_stage_1__7548_,
  data_stage_1__7547_,data_stage_1__7546_,data_stage_1__7545_,data_stage_1__7544_,
  data_stage_1__7543_,data_stage_1__7542_,data_stage_1__7541_,data_stage_1__7540_,
  data_stage_1__7539_,data_stage_1__7538_,data_stage_1__7537_,data_stage_1__7536_,
  data_stage_1__7535_,data_stage_1__7534_,data_stage_1__7533_,data_stage_1__7532_,
  data_stage_1__7531_,data_stage_1__7530_,data_stage_1__7529_,data_stage_1__7528_,
  data_stage_1__7527_,data_stage_1__7526_,data_stage_1__7525_,data_stage_1__7524_,
  data_stage_1__7523_,data_stage_1__7522_,data_stage_1__7521_,data_stage_1__7520_,
  data_stage_1__7519_,data_stage_1__7518_,data_stage_1__7517_,data_stage_1__7516_,
  data_stage_1__7515_,data_stage_1__7514_,data_stage_1__7513_,data_stage_1__7512_,
  data_stage_1__7511_,data_stage_1__7510_,data_stage_1__7509_,data_stage_1__7508_,
  data_stage_1__7507_,data_stage_1__7506_,data_stage_1__7505_,data_stage_1__7504_,
  data_stage_1__7503_,data_stage_1__7502_,data_stage_1__7501_,data_stage_1__7500_,
  data_stage_1__7499_,data_stage_1__7498_,data_stage_1__7497_,data_stage_1__7496_,
  data_stage_1__7495_,data_stage_1__7494_,data_stage_1__7493_,data_stage_1__7492_,
  data_stage_1__7491_,data_stage_1__7490_,data_stage_1__7489_,data_stage_1__7488_,
  data_stage_1__7487_,data_stage_1__7486_,data_stage_1__7485_,data_stage_1__7484_,
  data_stage_1__7483_,data_stage_1__7482_,data_stage_1__7481_,data_stage_1__7480_,
  data_stage_1__7479_,data_stage_1__7478_,data_stage_1__7477_,data_stage_1__7476_,
  data_stage_1__7475_,data_stage_1__7474_,data_stage_1__7473_,data_stage_1__7472_,
  data_stage_1__7471_,data_stage_1__7470_,data_stage_1__7469_,data_stage_1__7468_,
  data_stage_1__7467_,data_stage_1__7466_,data_stage_1__7465_,data_stage_1__7464_,
  data_stage_1__7463_,data_stage_1__7462_,data_stage_1__7461_,data_stage_1__7460_,
  data_stage_1__7459_,data_stage_1__7458_,data_stage_1__7457_,data_stage_1__7456_,
  data_stage_1__7455_,data_stage_1__7454_,data_stage_1__7453_,data_stage_1__7452_,
  data_stage_1__7451_,data_stage_1__7450_,data_stage_1__7449_,data_stage_1__7448_,
  data_stage_1__7447_,data_stage_1__7446_,data_stage_1__7445_,data_stage_1__7444_,
  data_stage_1__7443_,data_stage_1__7442_,data_stage_1__7441_,data_stage_1__7440_,
  data_stage_1__7439_,data_stage_1__7438_,data_stage_1__7437_,data_stage_1__7436_,
  data_stage_1__7435_,data_stage_1__7434_,data_stage_1__7433_,data_stage_1__7432_,
  data_stage_1__7431_,data_stage_1__7430_,data_stage_1__7429_,data_stage_1__7428_,
  data_stage_1__7427_,data_stage_1__7426_,data_stage_1__7425_,data_stage_1__7424_,
  data_stage_1__7423_,data_stage_1__7422_,data_stage_1__7421_,data_stage_1__7420_,
  data_stage_1__7419_,data_stage_1__7418_,data_stage_1__7417_,data_stage_1__7416_,
  data_stage_1__7415_,data_stage_1__7414_,data_stage_1__7413_,data_stage_1__7412_,
  data_stage_1__7411_,data_stage_1__7410_,data_stage_1__7409_,data_stage_1__7408_,
  data_stage_1__7407_,data_stage_1__7406_,data_stage_1__7405_,data_stage_1__7404_,
  data_stage_1__7403_,data_stage_1__7402_,data_stage_1__7401_,data_stage_1__7400_,
  data_stage_1__7399_,data_stage_1__7398_,data_stage_1__7397_,data_stage_1__7396_,
  data_stage_1__7395_,data_stage_1__7394_,data_stage_1__7393_,data_stage_1__7392_,
  data_stage_1__7391_,data_stage_1__7390_,data_stage_1__7389_,data_stage_1__7388_,
  data_stage_1__7387_,data_stage_1__7386_,data_stage_1__7385_,data_stage_1__7384_,
  data_stage_1__7383_,data_stage_1__7382_,data_stage_1__7381_,data_stage_1__7380_,
  data_stage_1__7379_,data_stage_1__7378_,data_stage_1__7377_,data_stage_1__7376_,
  data_stage_1__7375_,data_stage_1__7374_,data_stage_1__7373_,data_stage_1__7372_,
  data_stage_1__7371_,data_stage_1__7370_,data_stage_1__7369_,data_stage_1__7368_,
  data_stage_1__7367_,data_stage_1__7366_,data_stage_1__7365_,data_stage_1__7364_,
  data_stage_1__7363_,data_stage_1__7362_,data_stage_1__7361_,data_stage_1__7360_,
  data_stage_1__7359_,data_stage_1__7358_,data_stage_1__7357_,data_stage_1__7356_,
  data_stage_1__7355_,data_stage_1__7354_,data_stage_1__7353_,data_stage_1__7352_,
  data_stage_1__7351_,data_stage_1__7350_,data_stage_1__7349_,data_stage_1__7348_,
  data_stage_1__7347_,data_stage_1__7346_,data_stage_1__7345_,data_stage_1__7344_,
  data_stage_1__7343_,data_stage_1__7342_,data_stage_1__7341_,data_stage_1__7340_,
  data_stage_1__7339_,data_stage_1__7338_,data_stage_1__7337_,data_stage_1__7336_,
  data_stage_1__7335_,data_stage_1__7334_,data_stage_1__7333_,data_stage_1__7332_,
  data_stage_1__7331_,data_stage_1__7330_,data_stage_1__7329_,data_stage_1__7328_,
  data_stage_1__7327_,data_stage_1__7326_,data_stage_1__7325_,data_stage_1__7324_,
  data_stage_1__7323_,data_stage_1__7322_,data_stage_1__7321_,data_stage_1__7320_,
  data_stage_1__7319_,data_stage_1__7318_,data_stage_1__7317_,data_stage_1__7316_,
  data_stage_1__7315_,data_stage_1__7314_,data_stage_1__7313_,data_stage_1__7312_,
  data_stage_1__7311_,data_stage_1__7310_,data_stage_1__7309_,data_stage_1__7308_,
  data_stage_1__7307_,data_stage_1__7306_,data_stage_1__7305_,data_stage_1__7304_,
  data_stage_1__7303_,data_stage_1__7302_,data_stage_1__7301_,data_stage_1__7300_,
  data_stage_1__7299_,data_stage_1__7298_,data_stage_1__7297_,data_stage_1__7296_,
  data_stage_1__7295_,data_stage_1__7294_,data_stage_1__7293_,data_stage_1__7292_,
  data_stage_1__7291_,data_stage_1__7290_,data_stage_1__7289_,data_stage_1__7288_,
  data_stage_1__7287_,data_stage_1__7286_,data_stage_1__7285_,data_stage_1__7284_,
  data_stage_1__7283_,data_stage_1__7282_,data_stage_1__7281_,data_stage_1__7280_,
  data_stage_1__7279_,data_stage_1__7278_,data_stage_1__7277_,data_stage_1__7276_,
  data_stage_1__7275_,data_stage_1__7274_,data_stage_1__7273_,data_stage_1__7272_,
  data_stage_1__7271_,data_stage_1__7270_,data_stage_1__7269_,data_stage_1__7268_,
  data_stage_1__7267_,data_stage_1__7266_,data_stage_1__7265_,data_stage_1__7264_,
  data_stage_1__7263_,data_stage_1__7262_,data_stage_1__7261_,data_stage_1__7260_,
  data_stage_1__7259_,data_stage_1__7258_,data_stage_1__7257_,data_stage_1__7256_,
  data_stage_1__7255_,data_stage_1__7254_,data_stage_1__7253_,data_stage_1__7252_,
  data_stage_1__7251_,data_stage_1__7250_,data_stage_1__7249_,data_stage_1__7248_,
  data_stage_1__7247_,data_stage_1__7246_,data_stage_1__7245_,data_stage_1__7244_,
  data_stage_1__7243_,data_stage_1__7242_,data_stage_1__7241_,data_stage_1__7240_,
  data_stage_1__7239_,data_stage_1__7238_,data_stage_1__7237_,data_stage_1__7236_,
  data_stage_1__7235_,data_stage_1__7234_,data_stage_1__7233_,data_stage_1__7232_,
  data_stage_1__7231_,data_stage_1__7230_,data_stage_1__7229_,data_stage_1__7228_,
  data_stage_1__7227_,data_stage_1__7226_,data_stage_1__7225_,data_stage_1__7224_,
  data_stage_1__7223_,data_stage_1__7222_,data_stage_1__7221_,data_stage_1__7220_,
  data_stage_1__7219_,data_stage_1__7218_,data_stage_1__7217_,data_stage_1__7216_,
  data_stage_1__7215_,data_stage_1__7214_,data_stage_1__7213_,data_stage_1__7212_,
  data_stage_1__7211_,data_stage_1__7210_,data_stage_1__7209_,data_stage_1__7208_,
  data_stage_1__7207_,data_stage_1__7206_,data_stage_1__7205_,data_stage_1__7204_,
  data_stage_1__7203_,data_stage_1__7202_,data_stage_1__7201_,data_stage_1__7200_,
  data_stage_1__7199_,data_stage_1__7198_,data_stage_1__7197_,data_stage_1__7196_,
  data_stage_1__7195_,data_stage_1__7194_,data_stage_1__7193_,data_stage_1__7192_,
  data_stage_1__7191_,data_stage_1__7190_,data_stage_1__7189_,data_stage_1__7188_,
  data_stage_1__7187_,data_stage_1__7186_,data_stage_1__7185_,data_stage_1__7184_,
  data_stage_1__7183_,data_stage_1__7182_,data_stage_1__7181_,data_stage_1__7180_,
  data_stage_1__7179_,data_stage_1__7178_,data_stage_1__7177_,data_stage_1__7176_,
  data_stage_1__7175_,data_stage_1__7174_,data_stage_1__7173_,data_stage_1__7172_,
  data_stage_1__7171_,data_stage_1__7170_,data_stage_1__7169_,data_stage_1__7168_,
  data_stage_1__7167_,data_stage_1__7166_,data_stage_1__7165_,data_stage_1__7164_,
  data_stage_1__7163_,data_stage_1__7162_,data_stage_1__7161_,data_stage_1__7160_,
  data_stage_1__7159_,data_stage_1__7158_,data_stage_1__7157_,data_stage_1__7156_,
  data_stage_1__7155_,data_stage_1__7154_,data_stage_1__7153_,data_stage_1__7152_,
  data_stage_1__7151_,data_stage_1__7150_,data_stage_1__7149_,data_stage_1__7148_,
  data_stage_1__7147_,data_stage_1__7146_,data_stage_1__7145_,data_stage_1__7144_,
  data_stage_1__7143_,data_stage_1__7142_,data_stage_1__7141_,data_stage_1__7140_,
  data_stage_1__7139_,data_stage_1__7138_,data_stage_1__7137_,data_stage_1__7136_,
  data_stage_1__7135_,data_stage_1__7134_,data_stage_1__7133_,data_stage_1__7132_,
  data_stage_1__7131_,data_stage_1__7130_,data_stage_1__7129_,data_stage_1__7128_,
  data_stage_1__7127_,data_stage_1__7126_,data_stage_1__7125_,data_stage_1__7124_,
  data_stage_1__7123_,data_stage_1__7122_,data_stage_1__7121_,data_stage_1__7120_,
  data_stage_1__7119_,data_stage_1__7118_,data_stage_1__7117_,data_stage_1__7116_,
  data_stage_1__7115_,data_stage_1__7114_,data_stage_1__7113_,data_stage_1__7112_,
  data_stage_1__7111_,data_stage_1__7110_,data_stage_1__7109_,data_stage_1__7108_,
  data_stage_1__7107_,data_stage_1__7106_,data_stage_1__7105_,data_stage_1__7104_,
  data_stage_1__7103_,data_stage_1__7102_,data_stage_1__7101_,data_stage_1__7100_,
  data_stage_1__7099_,data_stage_1__7098_,data_stage_1__7097_,data_stage_1__7096_,
  data_stage_1__7095_,data_stage_1__7094_,data_stage_1__7093_,data_stage_1__7092_,
  data_stage_1__7091_,data_stage_1__7090_,data_stage_1__7089_,data_stage_1__7088_,
  data_stage_1__7087_,data_stage_1__7086_,data_stage_1__7085_,data_stage_1__7084_,
  data_stage_1__7083_,data_stage_1__7082_,data_stage_1__7081_,data_stage_1__7080_,
  data_stage_1__7079_,data_stage_1__7078_,data_stage_1__7077_,data_stage_1__7076_,
  data_stage_1__7075_,data_stage_1__7074_,data_stage_1__7073_,data_stage_1__7072_,
  data_stage_1__7071_,data_stage_1__7070_,data_stage_1__7069_,data_stage_1__7068_,
  data_stage_1__7067_,data_stage_1__7066_,data_stage_1__7065_,data_stage_1__7064_,
  data_stage_1__7063_,data_stage_1__7062_,data_stage_1__7061_,data_stage_1__7060_,
  data_stage_1__7059_,data_stage_1__7058_,data_stage_1__7057_,data_stage_1__7056_,
  data_stage_1__7055_,data_stage_1__7054_,data_stage_1__7053_,data_stage_1__7052_,
  data_stage_1__7051_,data_stage_1__7050_,data_stage_1__7049_,data_stage_1__7048_,
  data_stage_1__7047_,data_stage_1__7046_,data_stage_1__7045_,data_stage_1__7044_,
  data_stage_1__7043_,data_stage_1__7042_,data_stage_1__7041_,data_stage_1__7040_,
  data_stage_1__7039_,data_stage_1__7038_,data_stage_1__7037_,data_stage_1__7036_,
  data_stage_1__7035_,data_stage_1__7034_,data_stage_1__7033_,data_stage_1__7032_,
  data_stage_1__7031_,data_stage_1__7030_,data_stage_1__7029_,data_stage_1__7028_,
  data_stage_1__7027_,data_stage_1__7026_,data_stage_1__7025_,data_stage_1__7024_,
  data_stage_1__7023_,data_stage_1__7022_,data_stage_1__7021_,data_stage_1__7020_,
  data_stage_1__7019_,data_stage_1__7018_,data_stage_1__7017_,data_stage_1__7016_,
  data_stage_1__7015_,data_stage_1__7014_,data_stage_1__7013_,data_stage_1__7012_,
  data_stage_1__7011_,data_stage_1__7010_,data_stage_1__7009_,data_stage_1__7008_,
  data_stage_1__7007_,data_stage_1__7006_,data_stage_1__7005_,data_stage_1__7004_,
  data_stage_1__7003_,data_stage_1__7002_,data_stage_1__7001_,data_stage_1__7000_,
  data_stage_1__6999_,data_stage_1__6998_,data_stage_1__6997_,data_stage_1__6996_,
  data_stage_1__6995_,data_stage_1__6994_,data_stage_1__6993_,data_stage_1__6992_,
  data_stage_1__6991_,data_stage_1__6990_,data_stage_1__6989_,data_stage_1__6988_,
  data_stage_1__6987_,data_stage_1__6986_,data_stage_1__6985_,data_stage_1__6984_,
  data_stage_1__6983_,data_stage_1__6982_,data_stage_1__6981_,data_stage_1__6980_,
  data_stage_1__6979_,data_stage_1__6978_,data_stage_1__6977_,data_stage_1__6976_,
  data_stage_1__6975_,data_stage_1__6974_,data_stage_1__6973_,data_stage_1__6972_,
  data_stage_1__6971_,data_stage_1__6970_,data_stage_1__6969_,data_stage_1__6968_,
  data_stage_1__6967_,data_stage_1__6966_,data_stage_1__6965_,data_stage_1__6964_,
  data_stage_1__6963_,data_stage_1__6962_,data_stage_1__6961_,data_stage_1__6960_,
  data_stage_1__6959_,data_stage_1__6958_,data_stage_1__6957_,data_stage_1__6956_,
  data_stage_1__6955_,data_stage_1__6954_,data_stage_1__6953_,data_stage_1__6952_,
  data_stage_1__6951_,data_stage_1__6950_,data_stage_1__6949_,data_stage_1__6948_,
  data_stage_1__6947_,data_stage_1__6946_,data_stage_1__6945_,data_stage_1__6944_,
  data_stage_1__6943_,data_stage_1__6942_,data_stage_1__6941_,data_stage_1__6940_,
  data_stage_1__6939_,data_stage_1__6938_,data_stage_1__6937_,data_stage_1__6936_,
  data_stage_1__6935_,data_stage_1__6934_,data_stage_1__6933_,data_stage_1__6932_,
  data_stage_1__6931_,data_stage_1__6930_,data_stage_1__6929_,data_stage_1__6928_,
  data_stage_1__6927_,data_stage_1__6926_,data_stage_1__6925_,data_stage_1__6924_,
  data_stage_1__6923_,data_stage_1__6922_,data_stage_1__6921_,data_stage_1__6920_,
  data_stage_1__6919_,data_stage_1__6918_,data_stage_1__6917_,data_stage_1__6916_,
  data_stage_1__6915_,data_stage_1__6914_,data_stage_1__6913_,data_stage_1__6912_,
  data_stage_1__6911_,data_stage_1__6910_,data_stage_1__6909_,data_stage_1__6908_,
  data_stage_1__6907_,data_stage_1__6906_,data_stage_1__6905_,data_stage_1__6904_,
  data_stage_1__6903_,data_stage_1__6902_,data_stage_1__6901_,data_stage_1__6900_,
  data_stage_1__6899_,data_stage_1__6898_,data_stage_1__6897_,data_stage_1__6896_,
  data_stage_1__6895_,data_stage_1__6894_,data_stage_1__6893_,data_stage_1__6892_,
  data_stage_1__6891_,data_stage_1__6890_,data_stage_1__6889_,data_stage_1__6888_,
  data_stage_1__6887_,data_stage_1__6886_,data_stage_1__6885_,data_stage_1__6884_,
  data_stage_1__6883_,data_stage_1__6882_,data_stage_1__6881_,data_stage_1__6880_,
  data_stage_1__6879_,data_stage_1__6878_,data_stage_1__6877_,data_stage_1__6876_,
  data_stage_1__6875_,data_stage_1__6874_,data_stage_1__6873_,data_stage_1__6872_,
  data_stage_1__6871_,data_stage_1__6870_,data_stage_1__6869_,data_stage_1__6868_,
  data_stage_1__6867_,data_stage_1__6866_,data_stage_1__6865_,data_stage_1__6864_,
  data_stage_1__6863_,data_stage_1__6862_,data_stage_1__6861_,data_stage_1__6860_,
  data_stage_1__6859_,data_stage_1__6858_,data_stage_1__6857_,data_stage_1__6856_,
  data_stage_1__6855_,data_stage_1__6854_,data_stage_1__6853_,data_stage_1__6852_,
  data_stage_1__6851_,data_stage_1__6850_,data_stage_1__6849_,data_stage_1__6848_,
  data_stage_1__6847_,data_stage_1__6846_,data_stage_1__6845_,data_stage_1__6844_,
  data_stage_1__6843_,data_stage_1__6842_,data_stage_1__6841_,data_stage_1__6840_,
  data_stage_1__6839_,data_stage_1__6838_,data_stage_1__6837_,data_stage_1__6836_,
  data_stage_1__6835_,data_stage_1__6834_,data_stage_1__6833_,data_stage_1__6832_,
  data_stage_1__6831_,data_stage_1__6830_,data_stage_1__6829_,data_stage_1__6828_,
  data_stage_1__6827_,data_stage_1__6826_,data_stage_1__6825_,data_stage_1__6824_,
  data_stage_1__6823_,data_stage_1__6822_,data_stage_1__6821_,data_stage_1__6820_,
  data_stage_1__6819_,data_stage_1__6818_,data_stage_1__6817_,data_stage_1__6816_,
  data_stage_1__6815_,data_stage_1__6814_,data_stage_1__6813_,data_stage_1__6812_,
  data_stage_1__6811_,data_stage_1__6810_,data_stage_1__6809_,data_stage_1__6808_,
  data_stage_1__6807_,data_stage_1__6806_,data_stage_1__6805_,data_stage_1__6804_,
  data_stage_1__6803_,data_stage_1__6802_,data_stage_1__6801_,data_stage_1__6800_,
  data_stage_1__6799_,data_stage_1__6798_,data_stage_1__6797_,data_stage_1__6796_,
  data_stage_1__6795_,data_stage_1__6794_,data_stage_1__6793_,data_stage_1__6792_,
  data_stage_1__6791_,data_stage_1__6790_,data_stage_1__6789_,data_stage_1__6788_,
  data_stage_1__6787_,data_stage_1__6786_,data_stage_1__6785_,data_stage_1__6784_,
  data_stage_1__6783_,data_stage_1__6782_,data_stage_1__6781_,data_stage_1__6780_,
  data_stage_1__6779_,data_stage_1__6778_,data_stage_1__6777_,data_stage_1__6776_,
  data_stage_1__6775_,data_stage_1__6774_,data_stage_1__6773_,data_stage_1__6772_,
  data_stage_1__6771_,data_stage_1__6770_,data_stage_1__6769_,data_stage_1__6768_,
  data_stage_1__6767_,data_stage_1__6766_,data_stage_1__6765_,data_stage_1__6764_,
  data_stage_1__6763_,data_stage_1__6762_,data_stage_1__6761_,data_stage_1__6760_,
  data_stage_1__6759_,data_stage_1__6758_,data_stage_1__6757_,data_stage_1__6756_,
  data_stage_1__6755_,data_stage_1__6754_,data_stage_1__6753_,data_stage_1__6752_,
  data_stage_1__6751_,data_stage_1__6750_,data_stage_1__6749_,data_stage_1__6748_,
  data_stage_1__6747_,data_stage_1__6746_,data_stage_1__6745_,data_stage_1__6744_,
  data_stage_1__6743_,data_stage_1__6742_,data_stage_1__6741_,data_stage_1__6740_,
  data_stage_1__6739_,data_stage_1__6738_,data_stage_1__6737_,data_stage_1__6736_,
  data_stage_1__6735_,data_stage_1__6734_,data_stage_1__6733_,data_stage_1__6732_,
  data_stage_1__6731_,data_stage_1__6730_,data_stage_1__6729_,data_stage_1__6728_,
  data_stage_1__6727_,data_stage_1__6726_,data_stage_1__6725_,data_stage_1__6724_,
  data_stage_1__6723_,data_stage_1__6722_,data_stage_1__6721_,data_stage_1__6720_,
  data_stage_1__6719_,data_stage_1__6718_,data_stage_1__6717_,data_stage_1__6716_,
  data_stage_1__6715_,data_stage_1__6714_,data_stage_1__6713_,data_stage_1__6712_,
  data_stage_1__6711_,data_stage_1__6710_,data_stage_1__6709_,data_stage_1__6708_,
  data_stage_1__6707_,data_stage_1__6706_,data_stage_1__6705_,data_stage_1__6704_,
  data_stage_1__6703_,data_stage_1__6702_,data_stage_1__6701_,data_stage_1__6700_,
  data_stage_1__6699_,data_stage_1__6698_,data_stage_1__6697_,data_stage_1__6696_,
  data_stage_1__6695_,data_stage_1__6694_,data_stage_1__6693_,data_stage_1__6692_,
  data_stage_1__6691_,data_stage_1__6690_,data_stage_1__6689_,data_stage_1__6688_,
  data_stage_1__6687_,data_stage_1__6686_,data_stage_1__6685_,data_stage_1__6684_,
  data_stage_1__6683_,data_stage_1__6682_,data_stage_1__6681_,data_stage_1__6680_,
  data_stage_1__6679_,data_stage_1__6678_,data_stage_1__6677_,data_stage_1__6676_,
  data_stage_1__6675_,data_stage_1__6674_,data_stage_1__6673_,data_stage_1__6672_,
  data_stage_1__6671_,data_stage_1__6670_,data_stage_1__6669_,data_stage_1__6668_,
  data_stage_1__6667_,data_stage_1__6666_,data_stage_1__6665_,data_stage_1__6664_,
  data_stage_1__6663_,data_stage_1__6662_,data_stage_1__6661_,data_stage_1__6660_,
  data_stage_1__6659_,data_stage_1__6658_,data_stage_1__6657_,data_stage_1__6656_,
  data_stage_1__6655_,data_stage_1__6654_,data_stage_1__6653_,data_stage_1__6652_,
  data_stage_1__6651_,data_stage_1__6650_,data_stage_1__6649_,data_stage_1__6648_,
  data_stage_1__6647_,data_stage_1__6646_,data_stage_1__6645_,data_stage_1__6644_,
  data_stage_1__6643_,data_stage_1__6642_,data_stage_1__6641_,data_stage_1__6640_,
  data_stage_1__6639_,data_stage_1__6638_,data_stage_1__6637_,data_stage_1__6636_,
  data_stage_1__6635_,data_stage_1__6634_,data_stage_1__6633_,data_stage_1__6632_,
  data_stage_1__6631_,data_stage_1__6630_,data_stage_1__6629_,data_stage_1__6628_,
  data_stage_1__6627_,data_stage_1__6626_,data_stage_1__6625_,data_stage_1__6624_,
  data_stage_1__6623_,data_stage_1__6622_,data_stage_1__6621_,data_stage_1__6620_,
  data_stage_1__6619_,data_stage_1__6618_,data_stage_1__6617_,data_stage_1__6616_,
  data_stage_1__6615_,data_stage_1__6614_,data_stage_1__6613_,data_stage_1__6612_,
  data_stage_1__6611_,data_stage_1__6610_,data_stage_1__6609_,data_stage_1__6608_,
  data_stage_1__6607_,data_stage_1__6606_,data_stage_1__6605_,data_stage_1__6604_,
  data_stage_1__6603_,data_stage_1__6602_,data_stage_1__6601_,data_stage_1__6600_,
  data_stage_1__6599_,data_stage_1__6598_,data_stage_1__6597_,data_stage_1__6596_,
  data_stage_1__6595_,data_stage_1__6594_,data_stage_1__6593_,data_stage_1__6592_,
  data_stage_1__6591_,data_stage_1__6590_,data_stage_1__6589_,data_stage_1__6588_,
  data_stage_1__6587_,data_stage_1__6586_,data_stage_1__6585_,data_stage_1__6584_,
  data_stage_1__6583_,data_stage_1__6582_,data_stage_1__6581_,data_stage_1__6580_,
  data_stage_1__6579_,data_stage_1__6578_,data_stage_1__6577_,data_stage_1__6576_,
  data_stage_1__6575_,data_stage_1__6574_,data_stage_1__6573_,data_stage_1__6572_,
  data_stage_1__6571_,data_stage_1__6570_,data_stage_1__6569_,data_stage_1__6568_,
  data_stage_1__6567_,data_stage_1__6566_,data_stage_1__6565_,data_stage_1__6564_,
  data_stage_1__6563_,data_stage_1__6562_,data_stage_1__6561_,data_stage_1__6560_,
  data_stage_1__6559_,data_stage_1__6558_,data_stage_1__6557_,data_stage_1__6556_,
  data_stage_1__6555_,data_stage_1__6554_,data_stage_1__6553_,data_stage_1__6552_,
  data_stage_1__6551_,data_stage_1__6550_,data_stage_1__6549_,data_stage_1__6548_,
  data_stage_1__6547_,data_stage_1__6546_,data_stage_1__6545_,data_stage_1__6544_,
  data_stage_1__6543_,data_stage_1__6542_,data_stage_1__6541_,data_stage_1__6540_,
  data_stage_1__6539_,data_stage_1__6538_,data_stage_1__6537_,data_stage_1__6536_,
  data_stage_1__6535_,data_stage_1__6534_,data_stage_1__6533_,data_stage_1__6532_,
  data_stage_1__6531_,data_stage_1__6530_,data_stage_1__6529_,data_stage_1__6528_,
  data_stage_1__6527_,data_stage_1__6526_,data_stage_1__6525_,data_stage_1__6524_,
  data_stage_1__6523_,data_stage_1__6522_,data_stage_1__6521_,data_stage_1__6520_,
  data_stage_1__6519_,data_stage_1__6518_,data_stage_1__6517_,data_stage_1__6516_,
  data_stage_1__6515_,data_stage_1__6514_,data_stage_1__6513_,data_stage_1__6512_,
  data_stage_1__6511_,data_stage_1__6510_,data_stage_1__6509_,data_stage_1__6508_,
  data_stage_1__6507_,data_stage_1__6506_,data_stage_1__6505_,data_stage_1__6504_,
  data_stage_1__6503_,data_stage_1__6502_,data_stage_1__6501_,data_stage_1__6500_,
  data_stage_1__6499_,data_stage_1__6498_,data_stage_1__6497_,data_stage_1__6496_,
  data_stage_1__6495_,data_stage_1__6494_,data_stage_1__6493_,data_stage_1__6492_,
  data_stage_1__6491_,data_stage_1__6490_,data_stage_1__6489_,data_stage_1__6488_,
  data_stage_1__6487_,data_stage_1__6486_,data_stage_1__6485_,data_stage_1__6484_,
  data_stage_1__6483_,data_stage_1__6482_,data_stage_1__6481_,data_stage_1__6480_,
  data_stage_1__6479_,data_stage_1__6478_,data_stage_1__6477_,data_stage_1__6476_,
  data_stage_1__6475_,data_stage_1__6474_,data_stage_1__6473_,data_stage_1__6472_,
  data_stage_1__6471_,data_stage_1__6470_,data_stage_1__6469_,data_stage_1__6468_,
  data_stage_1__6467_,data_stage_1__6466_,data_stage_1__6465_,data_stage_1__6464_,
  data_stage_1__6463_,data_stage_1__6462_,data_stage_1__6461_,data_stage_1__6460_,
  data_stage_1__6459_,data_stage_1__6458_,data_stage_1__6457_,data_stage_1__6456_,
  data_stage_1__6455_,data_stage_1__6454_,data_stage_1__6453_,data_stage_1__6452_,
  data_stage_1__6451_,data_stage_1__6450_,data_stage_1__6449_,data_stage_1__6448_,
  data_stage_1__6447_,data_stage_1__6446_,data_stage_1__6445_,data_stage_1__6444_,
  data_stage_1__6443_,data_stage_1__6442_,data_stage_1__6441_,data_stage_1__6440_,
  data_stage_1__6439_,data_stage_1__6438_,data_stage_1__6437_,data_stage_1__6436_,
  data_stage_1__6435_,data_stage_1__6434_,data_stage_1__6433_,data_stage_1__6432_,
  data_stage_1__6431_,data_stage_1__6430_,data_stage_1__6429_,data_stage_1__6428_,
  data_stage_1__6427_,data_stage_1__6426_,data_stage_1__6425_,data_stage_1__6424_,
  data_stage_1__6423_,data_stage_1__6422_,data_stage_1__6421_,data_stage_1__6420_,
  data_stage_1__6419_,data_stage_1__6418_,data_stage_1__6417_,data_stage_1__6416_,
  data_stage_1__6415_,data_stage_1__6414_,data_stage_1__6413_,data_stage_1__6412_,
  data_stage_1__6411_,data_stage_1__6410_,data_stage_1__6409_,data_stage_1__6408_,
  data_stage_1__6407_,data_stage_1__6406_,data_stage_1__6405_,data_stage_1__6404_,
  data_stage_1__6403_,data_stage_1__6402_,data_stage_1__6401_,data_stage_1__6400_,
  data_stage_1__6399_,data_stage_1__6398_,data_stage_1__6397_,data_stage_1__6396_,
  data_stage_1__6395_,data_stage_1__6394_,data_stage_1__6393_,data_stage_1__6392_,
  data_stage_1__6391_,data_stage_1__6390_,data_stage_1__6389_,data_stage_1__6388_,
  data_stage_1__6387_,data_stage_1__6386_,data_stage_1__6385_,data_stage_1__6384_,
  data_stage_1__6383_,data_stage_1__6382_,data_stage_1__6381_,data_stage_1__6380_,
  data_stage_1__6379_,data_stage_1__6378_,data_stage_1__6377_,data_stage_1__6376_,
  data_stage_1__6375_,data_stage_1__6374_,data_stage_1__6373_,data_stage_1__6372_,
  data_stage_1__6371_,data_stage_1__6370_,data_stage_1__6369_,data_stage_1__6368_,
  data_stage_1__6367_,data_stage_1__6366_,data_stage_1__6365_,data_stage_1__6364_,
  data_stage_1__6363_,data_stage_1__6362_,data_stage_1__6361_,data_stage_1__6360_,
  data_stage_1__6359_,data_stage_1__6358_,data_stage_1__6357_,data_stage_1__6356_,
  data_stage_1__6355_,data_stage_1__6354_,data_stage_1__6353_,data_stage_1__6352_,
  data_stage_1__6351_,data_stage_1__6350_,data_stage_1__6349_,data_stage_1__6348_,
  data_stage_1__6347_,data_stage_1__6346_,data_stage_1__6345_,data_stage_1__6344_,
  data_stage_1__6343_,data_stage_1__6342_,data_stage_1__6341_,data_stage_1__6340_,
  data_stage_1__6339_,data_stage_1__6338_,data_stage_1__6337_,data_stage_1__6336_,
  data_stage_1__6335_,data_stage_1__6334_,data_stage_1__6333_,data_stage_1__6332_,
  data_stage_1__6331_,data_stage_1__6330_,data_stage_1__6329_,data_stage_1__6328_,
  data_stage_1__6327_,data_stage_1__6326_,data_stage_1__6325_,data_stage_1__6324_,
  data_stage_1__6323_,data_stage_1__6322_,data_stage_1__6321_,data_stage_1__6320_,
  data_stage_1__6319_,data_stage_1__6318_,data_stage_1__6317_,data_stage_1__6316_,
  data_stage_1__6315_,data_stage_1__6314_,data_stage_1__6313_,data_stage_1__6312_,
  data_stage_1__6311_,data_stage_1__6310_,data_stage_1__6309_,data_stage_1__6308_,
  data_stage_1__6307_,data_stage_1__6306_,data_stage_1__6305_,data_stage_1__6304_,
  data_stage_1__6303_,data_stage_1__6302_,data_stage_1__6301_,data_stage_1__6300_,
  data_stage_1__6299_,data_stage_1__6298_,data_stage_1__6297_,data_stage_1__6296_,
  data_stage_1__6295_,data_stage_1__6294_,data_stage_1__6293_,data_stage_1__6292_,
  data_stage_1__6291_,data_stage_1__6290_,data_stage_1__6289_,data_stage_1__6288_,
  data_stage_1__6287_,data_stage_1__6286_,data_stage_1__6285_,data_stage_1__6284_,
  data_stage_1__6283_,data_stage_1__6282_,data_stage_1__6281_,data_stage_1__6280_,
  data_stage_1__6279_,data_stage_1__6278_,data_stage_1__6277_,data_stage_1__6276_,
  data_stage_1__6275_,data_stage_1__6274_,data_stage_1__6273_,data_stage_1__6272_,
  data_stage_1__6271_,data_stage_1__6270_,data_stage_1__6269_,data_stage_1__6268_,
  data_stage_1__6267_,data_stage_1__6266_,data_stage_1__6265_,data_stage_1__6264_,
  data_stage_1__6263_,data_stage_1__6262_,data_stage_1__6261_,data_stage_1__6260_,
  data_stage_1__6259_,data_stage_1__6258_,data_stage_1__6257_,data_stage_1__6256_,
  data_stage_1__6255_,data_stage_1__6254_,data_stage_1__6253_,data_stage_1__6252_,
  data_stage_1__6251_,data_stage_1__6250_,data_stage_1__6249_,data_stage_1__6248_,
  data_stage_1__6247_,data_stage_1__6246_,data_stage_1__6245_,data_stage_1__6244_,
  data_stage_1__6243_,data_stage_1__6242_,data_stage_1__6241_,data_stage_1__6240_,
  data_stage_1__6239_,data_stage_1__6238_,data_stage_1__6237_,data_stage_1__6236_,
  data_stage_1__6235_,data_stage_1__6234_,data_stage_1__6233_,data_stage_1__6232_,
  data_stage_1__6231_,data_stage_1__6230_,data_stage_1__6229_,data_stage_1__6228_,
  data_stage_1__6227_,data_stage_1__6226_,data_stage_1__6225_,data_stage_1__6224_,
  data_stage_1__6223_,data_stage_1__6222_,data_stage_1__6221_,data_stage_1__6220_,
  data_stage_1__6219_,data_stage_1__6218_,data_stage_1__6217_,data_stage_1__6216_,
  data_stage_1__6215_,data_stage_1__6214_,data_stage_1__6213_,data_stage_1__6212_,
  data_stage_1__6211_,data_stage_1__6210_,data_stage_1__6209_,data_stage_1__6208_,
  data_stage_1__6207_,data_stage_1__6206_,data_stage_1__6205_,data_stage_1__6204_,
  data_stage_1__6203_,data_stage_1__6202_,data_stage_1__6201_,data_stage_1__6200_,
  data_stage_1__6199_,data_stage_1__6198_,data_stage_1__6197_,data_stage_1__6196_,
  data_stage_1__6195_,data_stage_1__6194_,data_stage_1__6193_,data_stage_1__6192_,
  data_stage_1__6191_,data_stage_1__6190_,data_stage_1__6189_,data_stage_1__6188_,
  data_stage_1__6187_,data_stage_1__6186_,data_stage_1__6185_,data_stage_1__6184_,
  data_stage_1__6183_,data_stage_1__6182_,data_stage_1__6181_,data_stage_1__6180_,
  data_stage_1__6179_,data_stage_1__6178_,data_stage_1__6177_,data_stage_1__6176_,
  data_stage_1__6175_,data_stage_1__6174_,data_stage_1__6173_,data_stage_1__6172_,
  data_stage_1__6171_,data_stage_1__6170_,data_stage_1__6169_,data_stage_1__6168_,
  data_stage_1__6167_,data_stage_1__6166_,data_stage_1__6165_,data_stage_1__6164_,
  data_stage_1__6163_,data_stage_1__6162_,data_stage_1__6161_,data_stage_1__6160_,
  data_stage_1__6159_,data_stage_1__6158_,data_stage_1__6157_,data_stage_1__6156_,
  data_stage_1__6155_,data_stage_1__6154_,data_stage_1__6153_,data_stage_1__6152_,
  data_stage_1__6151_,data_stage_1__6150_,data_stage_1__6149_,data_stage_1__6148_,
  data_stage_1__6147_,data_stage_1__6146_,data_stage_1__6145_,data_stage_1__6144_,
  data_stage_1__6143_,data_stage_1__6142_,data_stage_1__6141_,data_stage_1__6140_,
  data_stage_1__6139_,data_stage_1__6138_,data_stage_1__6137_,data_stage_1__6136_,
  data_stage_1__6135_,data_stage_1__6134_,data_stage_1__6133_,data_stage_1__6132_,
  data_stage_1__6131_,data_stage_1__6130_,data_stage_1__6129_,data_stage_1__6128_,
  data_stage_1__6127_,data_stage_1__6126_,data_stage_1__6125_,data_stage_1__6124_,
  data_stage_1__6123_,data_stage_1__6122_,data_stage_1__6121_,data_stage_1__6120_,
  data_stage_1__6119_,data_stage_1__6118_,data_stage_1__6117_,data_stage_1__6116_,
  data_stage_1__6115_,data_stage_1__6114_,data_stage_1__6113_,data_stage_1__6112_,
  data_stage_1__6111_,data_stage_1__6110_,data_stage_1__6109_,data_stage_1__6108_,
  data_stage_1__6107_,data_stage_1__6106_,data_stage_1__6105_,data_stage_1__6104_,
  data_stage_1__6103_,data_stage_1__6102_,data_stage_1__6101_,data_stage_1__6100_,
  data_stage_1__6099_,data_stage_1__6098_,data_stage_1__6097_,data_stage_1__6096_,
  data_stage_1__6095_,data_stage_1__6094_,data_stage_1__6093_,data_stage_1__6092_,
  data_stage_1__6091_,data_stage_1__6090_,data_stage_1__6089_,data_stage_1__6088_,
  data_stage_1__6087_,data_stage_1__6086_,data_stage_1__6085_,data_stage_1__6084_,
  data_stage_1__6083_,data_stage_1__6082_,data_stage_1__6081_,data_stage_1__6080_,
  data_stage_1__6079_,data_stage_1__6078_,data_stage_1__6077_,data_stage_1__6076_,
  data_stage_1__6075_,data_stage_1__6074_,data_stage_1__6073_,data_stage_1__6072_,
  data_stage_1__6071_,data_stage_1__6070_,data_stage_1__6069_,data_stage_1__6068_,
  data_stage_1__6067_,data_stage_1__6066_,data_stage_1__6065_,data_stage_1__6064_,
  data_stage_1__6063_,data_stage_1__6062_,data_stage_1__6061_,data_stage_1__6060_,
  data_stage_1__6059_,data_stage_1__6058_,data_stage_1__6057_,data_stage_1__6056_,
  data_stage_1__6055_,data_stage_1__6054_,data_stage_1__6053_,data_stage_1__6052_,
  data_stage_1__6051_,data_stage_1__6050_,data_stage_1__6049_,data_stage_1__6048_,
  data_stage_1__6047_,data_stage_1__6046_,data_stage_1__6045_,data_stage_1__6044_,
  data_stage_1__6043_,data_stage_1__6042_,data_stage_1__6041_,data_stage_1__6040_,
  data_stage_1__6039_,data_stage_1__6038_,data_stage_1__6037_,data_stage_1__6036_,
  data_stage_1__6035_,data_stage_1__6034_,data_stage_1__6033_,data_stage_1__6032_,
  data_stage_1__6031_,data_stage_1__6030_,data_stage_1__6029_,data_stage_1__6028_,
  data_stage_1__6027_,data_stage_1__6026_,data_stage_1__6025_,data_stage_1__6024_,
  data_stage_1__6023_,data_stage_1__6022_,data_stage_1__6021_,data_stage_1__6020_,
  data_stage_1__6019_,data_stage_1__6018_,data_stage_1__6017_,data_stage_1__6016_,
  data_stage_1__6015_,data_stage_1__6014_,data_stage_1__6013_,data_stage_1__6012_,
  data_stage_1__6011_,data_stage_1__6010_,data_stage_1__6009_,data_stage_1__6008_,
  data_stage_1__6007_,data_stage_1__6006_,data_stage_1__6005_,data_stage_1__6004_,
  data_stage_1__6003_,data_stage_1__6002_,data_stage_1__6001_,data_stage_1__6000_,
  data_stage_1__5999_,data_stage_1__5998_,data_stage_1__5997_,data_stage_1__5996_,
  data_stage_1__5995_,data_stage_1__5994_,data_stage_1__5993_,data_stage_1__5992_,
  data_stage_1__5991_,data_stage_1__5990_,data_stage_1__5989_,data_stage_1__5988_,
  data_stage_1__5987_,data_stage_1__5986_,data_stage_1__5985_,data_stage_1__5984_,
  data_stage_1__5983_,data_stage_1__5982_,data_stage_1__5981_,data_stage_1__5980_,
  data_stage_1__5979_,data_stage_1__5978_,data_stage_1__5977_,data_stage_1__5976_,
  data_stage_1__5975_,data_stage_1__5974_,data_stage_1__5973_,data_stage_1__5972_,
  data_stage_1__5971_,data_stage_1__5970_,data_stage_1__5969_,data_stage_1__5968_,
  data_stage_1__5967_,data_stage_1__5966_,data_stage_1__5965_,data_stage_1__5964_,
  data_stage_1__5963_,data_stage_1__5962_,data_stage_1__5961_,data_stage_1__5960_,
  data_stage_1__5959_,data_stage_1__5958_,data_stage_1__5957_,data_stage_1__5956_,
  data_stage_1__5955_,data_stage_1__5954_,data_stage_1__5953_,data_stage_1__5952_,
  data_stage_1__5951_,data_stage_1__5950_,data_stage_1__5949_,data_stage_1__5948_,
  data_stage_1__5947_,data_stage_1__5946_,data_stage_1__5945_,data_stage_1__5944_,
  data_stage_1__5943_,data_stage_1__5942_,data_stage_1__5941_,data_stage_1__5940_,
  data_stage_1__5939_,data_stage_1__5938_,data_stage_1__5937_,data_stage_1__5936_,
  data_stage_1__5935_,data_stage_1__5934_,data_stage_1__5933_,data_stage_1__5932_,
  data_stage_1__5931_,data_stage_1__5930_,data_stage_1__5929_,data_stage_1__5928_,
  data_stage_1__5927_,data_stage_1__5926_,data_stage_1__5925_,data_stage_1__5924_,
  data_stage_1__5923_,data_stage_1__5922_,data_stage_1__5921_,data_stage_1__5920_,
  data_stage_1__5919_,data_stage_1__5918_,data_stage_1__5917_,data_stage_1__5916_,
  data_stage_1__5915_,data_stage_1__5914_,data_stage_1__5913_,data_stage_1__5912_,
  data_stage_1__5911_,data_stage_1__5910_,data_stage_1__5909_,data_stage_1__5908_,
  data_stage_1__5907_,data_stage_1__5906_,data_stage_1__5905_,data_stage_1__5904_,
  data_stage_1__5903_,data_stage_1__5902_,data_stage_1__5901_,data_stage_1__5900_,
  data_stage_1__5899_,data_stage_1__5898_,data_stage_1__5897_,data_stage_1__5896_,
  data_stage_1__5895_,data_stage_1__5894_,data_stage_1__5893_,data_stage_1__5892_,
  data_stage_1__5891_,data_stage_1__5890_,data_stage_1__5889_,data_stage_1__5888_,
  data_stage_1__5887_,data_stage_1__5886_,data_stage_1__5885_,data_stage_1__5884_,
  data_stage_1__5883_,data_stage_1__5882_,data_stage_1__5881_,data_stage_1__5880_,
  data_stage_1__5879_,data_stage_1__5878_,data_stage_1__5877_,data_stage_1__5876_,
  data_stage_1__5875_,data_stage_1__5874_,data_stage_1__5873_,data_stage_1__5872_,
  data_stage_1__5871_,data_stage_1__5870_,data_stage_1__5869_,data_stage_1__5868_,
  data_stage_1__5867_,data_stage_1__5866_,data_stage_1__5865_,data_stage_1__5864_,
  data_stage_1__5863_,data_stage_1__5862_,data_stage_1__5861_,data_stage_1__5860_,
  data_stage_1__5859_,data_stage_1__5858_,data_stage_1__5857_,data_stage_1__5856_,
  data_stage_1__5855_,data_stage_1__5854_,data_stage_1__5853_,data_stage_1__5852_,
  data_stage_1__5851_,data_stage_1__5850_,data_stage_1__5849_,data_stage_1__5848_,
  data_stage_1__5847_,data_stage_1__5846_,data_stage_1__5845_,data_stage_1__5844_,
  data_stage_1__5843_,data_stage_1__5842_,data_stage_1__5841_,data_stage_1__5840_,
  data_stage_1__5839_,data_stage_1__5838_,data_stage_1__5837_,data_stage_1__5836_,
  data_stage_1__5835_,data_stage_1__5834_,data_stage_1__5833_,data_stage_1__5832_,
  data_stage_1__5831_,data_stage_1__5830_,data_stage_1__5829_,data_stage_1__5828_,
  data_stage_1__5827_,data_stage_1__5826_,data_stage_1__5825_,data_stage_1__5824_,
  data_stage_1__5823_,data_stage_1__5822_,data_stage_1__5821_,data_stage_1__5820_,
  data_stage_1__5819_,data_stage_1__5818_,data_stage_1__5817_,data_stage_1__5816_,
  data_stage_1__5815_,data_stage_1__5814_,data_stage_1__5813_,data_stage_1__5812_,
  data_stage_1__5811_,data_stage_1__5810_,data_stage_1__5809_,data_stage_1__5808_,
  data_stage_1__5807_,data_stage_1__5806_,data_stage_1__5805_,data_stage_1__5804_,
  data_stage_1__5803_,data_stage_1__5802_,data_stage_1__5801_,data_stage_1__5800_,
  data_stage_1__5799_,data_stage_1__5798_,data_stage_1__5797_,data_stage_1__5796_,
  data_stage_1__5795_,data_stage_1__5794_,data_stage_1__5793_,data_stage_1__5792_,
  data_stage_1__5791_,data_stage_1__5790_,data_stage_1__5789_,data_stage_1__5788_,
  data_stage_1__5787_,data_stage_1__5786_,data_stage_1__5785_,data_stage_1__5784_,
  data_stage_1__5783_,data_stage_1__5782_,data_stage_1__5781_,data_stage_1__5780_,
  data_stage_1__5779_,data_stage_1__5778_,data_stage_1__5777_,data_stage_1__5776_,
  data_stage_1__5775_,data_stage_1__5774_,data_stage_1__5773_,data_stage_1__5772_,
  data_stage_1__5771_,data_stage_1__5770_,data_stage_1__5769_,data_stage_1__5768_,
  data_stage_1__5767_,data_stage_1__5766_,data_stage_1__5765_,data_stage_1__5764_,
  data_stage_1__5763_,data_stage_1__5762_,data_stage_1__5761_,data_stage_1__5760_,
  data_stage_1__5759_,data_stage_1__5758_,data_stage_1__5757_,data_stage_1__5756_,
  data_stage_1__5755_,data_stage_1__5754_,data_stage_1__5753_,data_stage_1__5752_,
  data_stage_1__5751_,data_stage_1__5750_,data_stage_1__5749_,data_stage_1__5748_,
  data_stage_1__5747_,data_stage_1__5746_,data_stage_1__5745_,data_stage_1__5744_,
  data_stage_1__5743_,data_stage_1__5742_,data_stage_1__5741_,data_stage_1__5740_,
  data_stage_1__5739_,data_stage_1__5738_,data_stage_1__5737_,data_stage_1__5736_,
  data_stage_1__5735_,data_stage_1__5734_,data_stage_1__5733_,data_stage_1__5732_,
  data_stage_1__5731_,data_stage_1__5730_,data_stage_1__5729_,data_stage_1__5728_,
  data_stage_1__5727_,data_stage_1__5726_,data_stage_1__5725_,data_stage_1__5724_,
  data_stage_1__5723_,data_stage_1__5722_,data_stage_1__5721_,data_stage_1__5720_,
  data_stage_1__5719_,data_stage_1__5718_,data_stage_1__5717_,data_stage_1__5716_,
  data_stage_1__5715_,data_stage_1__5714_,data_stage_1__5713_,data_stage_1__5712_,
  data_stage_1__5711_,data_stage_1__5710_,data_stage_1__5709_,data_stage_1__5708_,
  data_stage_1__5707_,data_stage_1__5706_,data_stage_1__5705_,data_stage_1__5704_,
  data_stage_1__5703_,data_stage_1__5702_,data_stage_1__5701_,data_stage_1__5700_,
  data_stage_1__5699_,data_stage_1__5698_,data_stage_1__5697_,data_stage_1__5696_,
  data_stage_1__5695_,data_stage_1__5694_,data_stage_1__5693_,data_stage_1__5692_,
  data_stage_1__5691_,data_stage_1__5690_,data_stage_1__5689_,data_stage_1__5688_,
  data_stage_1__5687_,data_stage_1__5686_,data_stage_1__5685_,data_stage_1__5684_,
  data_stage_1__5683_,data_stage_1__5682_,data_stage_1__5681_,data_stage_1__5680_,
  data_stage_1__5679_,data_stage_1__5678_,data_stage_1__5677_,data_stage_1__5676_,
  data_stage_1__5675_,data_stage_1__5674_,data_stage_1__5673_,data_stage_1__5672_,
  data_stage_1__5671_,data_stage_1__5670_,data_stage_1__5669_,data_stage_1__5668_,
  data_stage_1__5667_,data_stage_1__5666_,data_stage_1__5665_,data_stage_1__5664_,
  data_stage_1__5663_,data_stage_1__5662_,data_stage_1__5661_,data_stage_1__5660_,
  data_stage_1__5659_,data_stage_1__5658_,data_stage_1__5657_,data_stage_1__5656_,
  data_stage_1__5655_,data_stage_1__5654_,data_stage_1__5653_,data_stage_1__5652_,
  data_stage_1__5651_,data_stage_1__5650_,data_stage_1__5649_,data_stage_1__5648_,
  data_stage_1__5647_,data_stage_1__5646_,data_stage_1__5645_,data_stage_1__5644_,
  data_stage_1__5643_,data_stage_1__5642_,data_stage_1__5641_,data_stage_1__5640_,
  data_stage_1__5639_,data_stage_1__5638_,data_stage_1__5637_,data_stage_1__5636_,
  data_stage_1__5635_,data_stage_1__5634_,data_stage_1__5633_,data_stage_1__5632_,
  data_stage_1__5631_,data_stage_1__5630_,data_stage_1__5629_,data_stage_1__5628_,
  data_stage_1__5627_,data_stage_1__5626_,data_stage_1__5625_,data_stage_1__5624_,
  data_stage_1__5623_,data_stage_1__5622_,data_stage_1__5621_,data_stage_1__5620_,
  data_stage_1__5619_,data_stage_1__5618_,data_stage_1__5617_,data_stage_1__5616_,
  data_stage_1__5615_,data_stage_1__5614_,data_stage_1__5613_,data_stage_1__5612_,
  data_stage_1__5611_,data_stage_1__5610_,data_stage_1__5609_,data_stage_1__5608_,
  data_stage_1__5607_,data_stage_1__5606_,data_stage_1__5605_,data_stage_1__5604_,
  data_stage_1__5603_,data_stage_1__5602_,data_stage_1__5601_,data_stage_1__5600_,
  data_stage_1__5599_,data_stage_1__5598_,data_stage_1__5597_,data_stage_1__5596_,
  data_stage_1__5595_,data_stage_1__5594_,data_stage_1__5593_,data_stage_1__5592_,
  data_stage_1__5591_,data_stage_1__5590_,data_stage_1__5589_,data_stage_1__5588_,
  data_stage_1__5587_,data_stage_1__5586_,data_stage_1__5585_,data_stage_1__5584_,
  data_stage_1__5583_,data_stage_1__5582_,data_stage_1__5581_,data_stage_1__5580_,
  data_stage_1__5579_,data_stage_1__5578_,data_stage_1__5577_,data_stage_1__5576_,
  data_stage_1__5575_,data_stage_1__5574_,data_stage_1__5573_,data_stage_1__5572_,
  data_stage_1__5571_,data_stage_1__5570_,data_stage_1__5569_,data_stage_1__5568_,
  data_stage_1__5567_,data_stage_1__5566_,data_stage_1__5565_,data_stage_1__5564_,
  data_stage_1__5563_,data_stage_1__5562_,data_stage_1__5561_,data_stage_1__5560_,
  data_stage_1__5559_,data_stage_1__5558_,data_stage_1__5557_,data_stage_1__5556_,
  data_stage_1__5555_,data_stage_1__5554_,data_stage_1__5553_,data_stage_1__5552_,
  data_stage_1__5551_,data_stage_1__5550_,data_stage_1__5549_,data_stage_1__5548_,
  data_stage_1__5547_,data_stage_1__5546_,data_stage_1__5545_,data_stage_1__5544_,
  data_stage_1__5543_,data_stage_1__5542_,data_stage_1__5541_,data_stage_1__5540_,
  data_stage_1__5539_,data_stage_1__5538_,data_stage_1__5537_,data_stage_1__5536_,
  data_stage_1__5535_,data_stage_1__5534_,data_stage_1__5533_,data_stage_1__5532_,
  data_stage_1__5531_,data_stage_1__5530_,data_stage_1__5529_,data_stage_1__5528_,
  data_stage_1__5527_,data_stage_1__5526_,data_stage_1__5525_,data_stage_1__5524_,
  data_stage_1__5523_,data_stage_1__5522_,data_stage_1__5521_,data_stage_1__5520_,
  data_stage_1__5519_,data_stage_1__5518_,data_stage_1__5517_,data_stage_1__5516_,
  data_stage_1__5515_,data_stage_1__5514_,data_stage_1__5513_,data_stage_1__5512_,
  data_stage_1__5511_,data_stage_1__5510_,data_stage_1__5509_,data_stage_1__5508_,
  data_stage_1__5507_,data_stage_1__5506_,data_stage_1__5505_,data_stage_1__5504_,
  data_stage_1__5503_,data_stage_1__5502_,data_stage_1__5501_,data_stage_1__5500_,
  data_stage_1__5499_,data_stage_1__5498_,data_stage_1__5497_,data_stage_1__5496_,
  data_stage_1__5495_,data_stage_1__5494_,data_stage_1__5493_,data_stage_1__5492_,
  data_stage_1__5491_,data_stage_1__5490_,data_stage_1__5489_,data_stage_1__5488_,
  data_stage_1__5487_,data_stage_1__5486_,data_stage_1__5485_,data_stage_1__5484_,
  data_stage_1__5483_,data_stage_1__5482_,data_stage_1__5481_,data_stage_1__5480_,
  data_stage_1__5479_,data_stage_1__5478_,data_stage_1__5477_,data_stage_1__5476_,
  data_stage_1__5475_,data_stage_1__5474_,data_stage_1__5473_,data_stage_1__5472_,
  data_stage_1__5471_,data_stage_1__5470_,data_stage_1__5469_,data_stage_1__5468_,
  data_stage_1__5467_,data_stage_1__5466_,data_stage_1__5465_,data_stage_1__5464_,
  data_stage_1__5463_,data_stage_1__5462_,data_stage_1__5461_,data_stage_1__5460_,
  data_stage_1__5459_,data_stage_1__5458_,data_stage_1__5457_,data_stage_1__5456_,
  data_stage_1__5455_,data_stage_1__5454_,data_stage_1__5453_,data_stage_1__5452_,
  data_stage_1__5451_,data_stage_1__5450_,data_stage_1__5449_,data_stage_1__5448_,
  data_stage_1__5447_,data_stage_1__5446_,data_stage_1__5445_,data_stage_1__5444_,
  data_stage_1__5443_,data_stage_1__5442_,data_stage_1__5441_,data_stage_1__5440_,
  data_stage_1__5439_,data_stage_1__5438_,data_stage_1__5437_,data_stage_1__5436_,
  data_stage_1__5435_,data_stage_1__5434_,data_stage_1__5433_,data_stage_1__5432_,
  data_stage_1__5431_,data_stage_1__5430_,data_stage_1__5429_,data_stage_1__5428_,
  data_stage_1__5427_,data_stage_1__5426_,data_stage_1__5425_,data_stage_1__5424_,
  data_stage_1__5423_,data_stage_1__5422_,data_stage_1__5421_,data_stage_1__5420_,
  data_stage_1__5419_,data_stage_1__5418_,data_stage_1__5417_,data_stage_1__5416_,
  data_stage_1__5415_,data_stage_1__5414_,data_stage_1__5413_,data_stage_1__5412_,
  data_stage_1__5411_,data_stage_1__5410_,data_stage_1__5409_,data_stage_1__5408_,
  data_stage_1__5407_,data_stage_1__5406_,data_stage_1__5405_,data_stage_1__5404_,
  data_stage_1__5403_,data_stage_1__5402_,data_stage_1__5401_,data_stage_1__5400_,
  data_stage_1__5399_,data_stage_1__5398_,data_stage_1__5397_,data_stage_1__5396_,
  data_stage_1__5395_,data_stage_1__5394_,data_stage_1__5393_,data_stage_1__5392_,
  data_stage_1__5391_,data_stage_1__5390_,data_stage_1__5389_,data_stage_1__5388_,
  data_stage_1__5387_,data_stage_1__5386_,data_stage_1__5385_,data_stage_1__5384_,
  data_stage_1__5383_,data_stage_1__5382_,data_stage_1__5381_,data_stage_1__5380_,
  data_stage_1__5379_,data_stage_1__5378_,data_stage_1__5377_,data_stage_1__5376_,
  data_stage_1__5375_,data_stage_1__5374_,data_stage_1__5373_,data_stage_1__5372_,
  data_stage_1__5371_,data_stage_1__5370_,data_stage_1__5369_,data_stage_1__5368_,
  data_stage_1__5367_,data_stage_1__5366_,data_stage_1__5365_,data_stage_1__5364_,
  data_stage_1__5363_,data_stage_1__5362_,data_stage_1__5361_,data_stage_1__5360_,
  data_stage_1__5359_,data_stage_1__5358_,data_stage_1__5357_,data_stage_1__5356_,
  data_stage_1__5355_,data_stage_1__5354_,data_stage_1__5353_,data_stage_1__5352_,
  data_stage_1__5351_,data_stage_1__5350_,data_stage_1__5349_,data_stage_1__5348_,
  data_stage_1__5347_,data_stage_1__5346_,data_stage_1__5345_,data_stage_1__5344_,
  data_stage_1__5343_,data_stage_1__5342_,data_stage_1__5341_,data_stage_1__5340_,
  data_stage_1__5339_,data_stage_1__5338_,data_stage_1__5337_,data_stage_1__5336_,
  data_stage_1__5335_,data_stage_1__5334_,data_stage_1__5333_,data_stage_1__5332_,
  data_stage_1__5331_,data_stage_1__5330_,data_stage_1__5329_,data_stage_1__5328_,
  data_stage_1__5327_,data_stage_1__5326_,data_stage_1__5325_,data_stage_1__5324_,
  data_stage_1__5323_,data_stage_1__5322_,data_stage_1__5321_,data_stage_1__5320_,
  data_stage_1__5319_,data_stage_1__5318_,data_stage_1__5317_,data_stage_1__5316_,
  data_stage_1__5315_,data_stage_1__5314_,data_stage_1__5313_,data_stage_1__5312_,
  data_stage_1__5311_,data_stage_1__5310_,data_stage_1__5309_,data_stage_1__5308_,
  data_stage_1__5307_,data_stage_1__5306_,data_stage_1__5305_,data_stage_1__5304_,
  data_stage_1__5303_,data_stage_1__5302_,data_stage_1__5301_,data_stage_1__5300_,
  data_stage_1__5299_,data_stage_1__5298_,data_stage_1__5297_,data_stage_1__5296_,
  data_stage_1__5295_,data_stage_1__5294_,data_stage_1__5293_,data_stage_1__5292_,
  data_stage_1__5291_,data_stage_1__5290_,data_stage_1__5289_,data_stage_1__5288_,
  data_stage_1__5287_,data_stage_1__5286_,data_stage_1__5285_,data_stage_1__5284_,
  data_stage_1__5283_,data_stage_1__5282_,data_stage_1__5281_,data_stage_1__5280_,
  data_stage_1__5279_,data_stage_1__5278_,data_stage_1__5277_,data_stage_1__5276_,
  data_stage_1__5275_,data_stage_1__5274_,data_stage_1__5273_,data_stage_1__5272_,
  data_stage_1__5271_,data_stage_1__5270_,data_stage_1__5269_,data_stage_1__5268_,
  data_stage_1__5267_,data_stage_1__5266_,data_stage_1__5265_,data_stage_1__5264_,
  data_stage_1__5263_,data_stage_1__5262_,data_stage_1__5261_,data_stage_1__5260_,
  data_stage_1__5259_,data_stage_1__5258_,data_stage_1__5257_,data_stage_1__5256_,
  data_stage_1__5255_,data_stage_1__5254_,data_stage_1__5253_,data_stage_1__5252_,
  data_stage_1__5251_,data_stage_1__5250_,data_stage_1__5249_,data_stage_1__5248_,
  data_stage_1__5247_,data_stage_1__5246_,data_stage_1__5245_,data_stage_1__5244_,
  data_stage_1__5243_,data_stage_1__5242_,data_stage_1__5241_,data_stage_1__5240_,
  data_stage_1__5239_,data_stage_1__5238_,data_stage_1__5237_,data_stage_1__5236_,
  data_stage_1__5235_,data_stage_1__5234_,data_stage_1__5233_,data_stage_1__5232_,
  data_stage_1__5231_,data_stage_1__5230_,data_stage_1__5229_,data_stage_1__5228_,
  data_stage_1__5227_,data_stage_1__5226_,data_stage_1__5225_,data_stage_1__5224_,
  data_stage_1__5223_,data_stage_1__5222_,data_stage_1__5221_,data_stage_1__5220_,
  data_stage_1__5219_,data_stage_1__5218_,data_stage_1__5217_,data_stage_1__5216_,
  data_stage_1__5215_,data_stage_1__5214_,data_stage_1__5213_,data_stage_1__5212_,
  data_stage_1__5211_,data_stage_1__5210_,data_stage_1__5209_,data_stage_1__5208_,
  data_stage_1__5207_,data_stage_1__5206_,data_stage_1__5205_,data_stage_1__5204_,
  data_stage_1__5203_,data_stage_1__5202_,data_stage_1__5201_,data_stage_1__5200_,
  data_stage_1__5199_,data_stage_1__5198_,data_stage_1__5197_,data_stage_1__5196_,
  data_stage_1__5195_,data_stage_1__5194_,data_stage_1__5193_,data_stage_1__5192_,
  data_stage_1__5191_,data_stage_1__5190_,data_stage_1__5189_,data_stage_1__5188_,
  data_stage_1__5187_,data_stage_1__5186_,data_stage_1__5185_,data_stage_1__5184_,
  data_stage_1__5183_,data_stage_1__5182_,data_stage_1__5181_,data_stage_1__5180_,
  data_stage_1__5179_,data_stage_1__5178_,data_stage_1__5177_,data_stage_1__5176_,
  data_stage_1__5175_,data_stage_1__5174_,data_stage_1__5173_,data_stage_1__5172_,
  data_stage_1__5171_,data_stage_1__5170_,data_stage_1__5169_,data_stage_1__5168_,
  data_stage_1__5167_,data_stage_1__5166_,data_stage_1__5165_,data_stage_1__5164_,
  data_stage_1__5163_,data_stage_1__5162_,data_stage_1__5161_,data_stage_1__5160_,
  data_stage_1__5159_,data_stage_1__5158_,data_stage_1__5157_,data_stage_1__5156_,
  data_stage_1__5155_,data_stage_1__5154_,data_stage_1__5153_,data_stage_1__5152_,
  data_stage_1__5151_,data_stage_1__5150_,data_stage_1__5149_,data_stage_1__5148_,
  data_stage_1__5147_,data_stage_1__5146_,data_stage_1__5145_,data_stage_1__5144_,
  data_stage_1__5143_,data_stage_1__5142_,data_stage_1__5141_,data_stage_1__5140_,
  data_stage_1__5139_,data_stage_1__5138_,data_stage_1__5137_,data_stage_1__5136_,
  data_stage_1__5135_,data_stage_1__5134_,data_stage_1__5133_,data_stage_1__5132_,
  data_stage_1__5131_,data_stage_1__5130_,data_stage_1__5129_,data_stage_1__5128_,
  data_stage_1__5127_,data_stage_1__5126_,data_stage_1__5125_,data_stage_1__5124_,
  data_stage_1__5123_,data_stage_1__5122_,data_stage_1__5121_,data_stage_1__5120_,
  data_stage_1__5119_,data_stage_1__5118_,data_stage_1__5117_,data_stage_1__5116_,
  data_stage_1__5115_,data_stage_1__5114_,data_stage_1__5113_,data_stage_1__5112_,
  data_stage_1__5111_,data_stage_1__5110_,data_stage_1__5109_,data_stage_1__5108_,
  data_stage_1__5107_,data_stage_1__5106_,data_stage_1__5105_,data_stage_1__5104_,
  data_stage_1__5103_,data_stage_1__5102_,data_stage_1__5101_,data_stage_1__5100_,
  data_stage_1__5099_,data_stage_1__5098_,data_stage_1__5097_,data_stage_1__5096_,
  data_stage_1__5095_,data_stage_1__5094_,data_stage_1__5093_,data_stage_1__5092_,
  data_stage_1__5091_,data_stage_1__5090_,data_stage_1__5089_,data_stage_1__5088_,
  data_stage_1__5087_,data_stage_1__5086_,data_stage_1__5085_,data_stage_1__5084_,
  data_stage_1__5083_,data_stage_1__5082_,data_stage_1__5081_,data_stage_1__5080_,
  data_stage_1__5079_,data_stage_1__5078_,data_stage_1__5077_,data_stage_1__5076_,
  data_stage_1__5075_,data_stage_1__5074_,data_stage_1__5073_,data_stage_1__5072_,
  data_stage_1__5071_,data_stage_1__5070_,data_stage_1__5069_,data_stage_1__5068_,
  data_stage_1__5067_,data_stage_1__5066_,data_stage_1__5065_,data_stage_1__5064_,
  data_stage_1__5063_,data_stage_1__5062_,data_stage_1__5061_,data_stage_1__5060_,
  data_stage_1__5059_,data_stage_1__5058_,data_stage_1__5057_,data_stage_1__5056_,
  data_stage_1__5055_,data_stage_1__5054_,data_stage_1__5053_,data_stage_1__5052_,
  data_stage_1__5051_,data_stage_1__5050_,data_stage_1__5049_,data_stage_1__5048_,
  data_stage_1__5047_,data_stage_1__5046_,data_stage_1__5045_,data_stage_1__5044_,
  data_stage_1__5043_,data_stage_1__5042_,data_stage_1__5041_,data_stage_1__5040_,
  data_stage_1__5039_,data_stage_1__5038_,data_stage_1__5037_,data_stage_1__5036_,
  data_stage_1__5035_,data_stage_1__5034_,data_stage_1__5033_,data_stage_1__5032_,
  data_stage_1__5031_,data_stage_1__5030_,data_stage_1__5029_,data_stage_1__5028_,
  data_stage_1__5027_,data_stage_1__5026_,data_stage_1__5025_,data_stage_1__5024_,
  data_stage_1__5023_,data_stage_1__5022_,data_stage_1__5021_,data_stage_1__5020_,
  data_stage_1__5019_,data_stage_1__5018_,data_stage_1__5017_,data_stage_1__5016_,
  data_stage_1__5015_,data_stage_1__5014_,data_stage_1__5013_,data_stage_1__5012_,
  data_stage_1__5011_,data_stage_1__5010_,data_stage_1__5009_,data_stage_1__5008_,
  data_stage_1__5007_,data_stage_1__5006_,data_stage_1__5005_,data_stage_1__5004_,
  data_stage_1__5003_,data_stage_1__5002_,data_stage_1__5001_,data_stage_1__5000_,
  data_stage_1__4999_,data_stage_1__4998_,data_stage_1__4997_,data_stage_1__4996_,
  data_stage_1__4995_,data_stage_1__4994_,data_stage_1__4993_,data_stage_1__4992_,
  data_stage_1__4991_,data_stage_1__4990_,data_stage_1__4989_,data_stage_1__4988_,
  data_stage_1__4987_,data_stage_1__4986_,data_stage_1__4985_,data_stage_1__4984_,
  data_stage_1__4983_,data_stage_1__4982_,data_stage_1__4981_,data_stage_1__4980_,
  data_stage_1__4979_,data_stage_1__4978_,data_stage_1__4977_,data_stage_1__4976_,
  data_stage_1__4975_,data_stage_1__4974_,data_stage_1__4973_,data_stage_1__4972_,
  data_stage_1__4971_,data_stage_1__4970_,data_stage_1__4969_,data_stage_1__4968_,
  data_stage_1__4967_,data_stage_1__4966_,data_stage_1__4965_,data_stage_1__4964_,
  data_stage_1__4963_,data_stage_1__4962_,data_stage_1__4961_,data_stage_1__4960_,
  data_stage_1__4959_,data_stage_1__4958_,data_stage_1__4957_,data_stage_1__4956_,
  data_stage_1__4955_,data_stage_1__4954_,data_stage_1__4953_,data_stage_1__4952_,
  data_stage_1__4951_,data_stage_1__4950_,data_stage_1__4949_,data_stage_1__4948_,
  data_stage_1__4947_,data_stage_1__4946_,data_stage_1__4945_,data_stage_1__4944_,
  data_stage_1__4943_,data_stage_1__4942_,data_stage_1__4941_,data_stage_1__4940_,
  data_stage_1__4939_,data_stage_1__4938_,data_stage_1__4937_,data_stage_1__4936_,
  data_stage_1__4935_,data_stage_1__4934_,data_stage_1__4933_,data_stage_1__4932_,
  data_stage_1__4931_,data_stage_1__4930_,data_stage_1__4929_,data_stage_1__4928_,
  data_stage_1__4927_,data_stage_1__4926_,data_stage_1__4925_,data_stage_1__4924_,
  data_stage_1__4923_,data_stage_1__4922_,data_stage_1__4921_,data_stage_1__4920_,
  data_stage_1__4919_,data_stage_1__4918_,data_stage_1__4917_,data_stage_1__4916_,
  data_stage_1__4915_,data_stage_1__4914_,data_stage_1__4913_,data_stage_1__4912_,
  data_stage_1__4911_,data_stage_1__4910_,data_stage_1__4909_,data_stage_1__4908_,
  data_stage_1__4907_,data_stage_1__4906_,data_stage_1__4905_,data_stage_1__4904_,
  data_stage_1__4903_,data_stage_1__4902_,data_stage_1__4901_,data_stage_1__4900_,
  data_stage_1__4899_,data_stage_1__4898_,data_stage_1__4897_,data_stage_1__4896_,
  data_stage_1__4895_,data_stage_1__4894_,data_stage_1__4893_,data_stage_1__4892_,
  data_stage_1__4891_,data_stage_1__4890_,data_stage_1__4889_,data_stage_1__4888_,
  data_stage_1__4887_,data_stage_1__4886_,data_stage_1__4885_,data_stage_1__4884_,
  data_stage_1__4883_,data_stage_1__4882_,data_stage_1__4881_,data_stage_1__4880_,
  data_stage_1__4879_,data_stage_1__4878_,data_stage_1__4877_,data_stage_1__4876_,
  data_stage_1__4875_,data_stage_1__4874_,data_stage_1__4873_,data_stage_1__4872_,
  data_stage_1__4871_,data_stage_1__4870_,data_stage_1__4869_,data_stage_1__4868_,
  data_stage_1__4867_,data_stage_1__4866_,data_stage_1__4865_,data_stage_1__4864_,
  data_stage_1__4863_,data_stage_1__4862_,data_stage_1__4861_,data_stage_1__4860_,
  data_stage_1__4859_,data_stage_1__4858_,data_stage_1__4857_,data_stage_1__4856_,
  data_stage_1__4855_,data_stage_1__4854_,data_stage_1__4853_,data_stage_1__4852_,
  data_stage_1__4851_,data_stage_1__4850_,data_stage_1__4849_,data_stage_1__4848_,
  data_stage_1__4847_,data_stage_1__4846_,data_stage_1__4845_,data_stage_1__4844_,
  data_stage_1__4843_,data_stage_1__4842_,data_stage_1__4841_,data_stage_1__4840_,
  data_stage_1__4839_,data_stage_1__4838_,data_stage_1__4837_,data_stage_1__4836_,
  data_stage_1__4835_,data_stage_1__4834_,data_stage_1__4833_,data_stage_1__4832_,
  data_stage_1__4831_,data_stage_1__4830_,data_stage_1__4829_,data_stage_1__4828_,
  data_stage_1__4827_,data_stage_1__4826_,data_stage_1__4825_,data_stage_1__4824_,
  data_stage_1__4823_,data_stage_1__4822_,data_stage_1__4821_,data_stage_1__4820_,
  data_stage_1__4819_,data_stage_1__4818_,data_stage_1__4817_,data_stage_1__4816_,
  data_stage_1__4815_,data_stage_1__4814_,data_stage_1__4813_,data_stage_1__4812_,
  data_stage_1__4811_,data_stage_1__4810_,data_stage_1__4809_,data_stage_1__4808_,
  data_stage_1__4807_,data_stage_1__4806_,data_stage_1__4805_,data_stage_1__4804_,
  data_stage_1__4803_,data_stage_1__4802_,data_stage_1__4801_,data_stage_1__4800_,
  data_stage_1__4799_,data_stage_1__4798_,data_stage_1__4797_,data_stage_1__4796_,
  data_stage_1__4795_,data_stage_1__4794_,data_stage_1__4793_,data_stage_1__4792_,
  data_stage_1__4791_,data_stage_1__4790_,data_stage_1__4789_,data_stage_1__4788_,
  data_stage_1__4787_,data_stage_1__4786_,data_stage_1__4785_,data_stage_1__4784_,
  data_stage_1__4783_,data_stage_1__4782_,data_stage_1__4781_,data_stage_1__4780_,
  data_stage_1__4779_,data_stage_1__4778_,data_stage_1__4777_,data_stage_1__4776_,
  data_stage_1__4775_,data_stage_1__4774_,data_stage_1__4773_,data_stage_1__4772_,
  data_stage_1__4771_,data_stage_1__4770_,data_stage_1__4769_,data_stage_1__4768_,
  data_stage_1__4767_,data_stage_1__4766_,data_stage_1__4765_,data_stage_1__4764_,
  data_stage_1__4763_,data_stage_1__4762_,data_stage_1__4761_,data_stage_1__4760_,
  data_stage_1__4759_,data_stage_1__4758_,data_stage_1__4757_,data_stage_1__4756_,
  data_stage_1__4755_,data_stage_1__4754_,data_stage_1__4753_,data_stage_1__4752_,
  data_stage_1__4751_,data_stage_1__4750_,data_stage_1__4749_,data_stage_1__4748_,
  data_stage_1__4747_,data_stage_1__4746_,data_stage_1__4745_,data_stage_1__4744_,
  data_stage_1__4743_,data_stage_1__4742_,data_stage_1__4741_,data_stage_1__4740_,
  data_stage_1__4739_,data_stage_1__4738_,data_stage_1__4737_,data_stage_1__4736_,
  data_stage_1__4735_,data_stage_1__4734_,data_stage_1__4733_,data_stage_1__4732_,
  data_stage_1__4731_,data_stage_1__4730_,data_stage_1__4729_,data_stage_1__4728_,
  data_stage_1__4727_,data_stage_1__4726_,data_stage_1__4725_,data_stage_1__4724_,
  data_stage_1__4723_,data_stage_1__4722_,data_stage_1__4721_,data_stage_1__4720_,
  data_stage_1__4719_,data_stage_1__4718_,data_stage_1__4717_,data_stage_1__4716_,
  data_stage_1__4715_,data_stage_1__4714_,data_stage_1__4713_,data_stage_1__4712_,
  data_stage_1__4711_,data_stage_1__4710_,data_stage_1__4709_,data_stage_1__4708_,
  data_stage_1__4707_,data_stage_1__4706_,data_stage_1__4705_,data_stage_1__4704_,
  data_stage_1__4703_,data_stage_1__4702_,data_stage_1__4701_,data_stage_1__4700_,
  data_stage_1__4699_,data_stage_1__4698_,data_stage_1__4697_,data_stage_1__4696_,
  data_stage_1__4695_,data_stage_1__4694_,data_stage_1__4693_,data_stage_1__4692_,
  data_stage_1__4691_,data_stage_1__4690_,data_stage_1__4689_,data_stage_1__4688_,
  data_stage_1__4687_,data_stage_1__4686_,data_stage_1__4685_,data_stage_1__4684_,
  data_stage_1__4683_,data_stage_1__4682_,data_stage_1__4681_,data_stage_1__4680_,
  data_stage_1__4679_,data_stage_1__4678_,data_stage_1__4677_,data_stage_1__4676_,
  data_stage_1__4675_,data_stage_1__4674_,data_stage_1__4673_,data_stage_1__4672_,
  data_stage_1__4671_,data_stage_1__4670_,data_stage_1__4669_,data_stage_1__4668_,
  data_stage_1__4667_,data_stage_1__4666_,data_stage_1__4665_,data_stage_1__4664_,
  data_stage_1__4663_,data_stage_1__4662_,data_stage_1__4661_,data_stage_1__4660_,
  data_stage_1__4659_,data_stage_1__4658_,data_stage_1__4657_,data_stage_1__4656_,
  data_stage_1__4655_,data_stage_1__4654_,data_stage_1__4653_,data_stage_1__4652_,
  data_stage_1__4651_,data_stage_1__4650_,data_stage_1__4649_,data_stage_1__4648_,
  data_stage_1__4647_,data_stage_1__4646_,data_stage_1__4645_,data_stage_1__4644_,
  data_stage_1__4643_,data_stage_1__4642_,data_stage_1__4641_,data_stage_1__4640_,
  data_stage_1__4639_,data_stage_1__4638_,data_stage_1__4637_,data_stage_1__4636_,
  data_stage_1__4635_,data_stage_1__4634_,data_stage_1__4633_,data_stage_1__4632_,
  data_stage_1__4631_,data_stage_1__4630_,data_stage_1__4629_,data_stage_1__4628_,
  data_stage_1__4627_,data_stage_1__4626_,data_stage_1__4625_,data_stage_1__4624_,
  data_stage_1__4623_,data_stage_1__4622_,data_stage_1__4621_,data_stage_1__4620_,
  data_stage_1__4619_,data_stage_1__4618_,data_stage_1__4617_,data_stage_1__4616_,
  data_stage_1__4615_,data_stage_1__4614_,data_stage_1__4613_,data_stage_1__4612_,
  data_stage_1__4611_,data_stage_1__4610_,data_stage_1__4609_,data_stage_1__4608_,
  data_stage_1__4607_,data_stage_1__4606_,data_stage_1__4605_,data_stage_1__4604_,
  data_stage_1__4603_,data_stage_1__4602_,data_stage_1__4601_,data_stage_1__4600_,
  data_stage_1__4599_,data_stage_1__4598_,data_stage_1__4597_,data_stage_1__4596_,
  data_stage_1__4595_,data_stage_1__4594_,data_stage_1__4593_,data_stage_1__4592_,
  data_stage_1__4591_,data_stage_1__4590_,data_stage_1__4589_,data_stage_1__4588_,
  data_stage_1__4587_,data_stage_1__4586_,data_stage_1__4585_,data_stage_1__4584_,
  data_stage_1__4583_,data_stage_1__4582_,data_stage_1__4581_,data_stage_1__4580_,
  data_stage_1__4579_,data_stage_1__4578_,data_stage_1__4577_,data_stage_1__4576_,
  data_stage_1__4575_,data_stage_1__4574_,data_stage_1__4573_,data_stage_1__4572_,
  data_stage_1__4571_,data_stage_1__4570_,data_stage_1__4569_,data_stage_1__4568_,
  data_stage_1__4567_,data_stage_1__4566_,data_stage_1__4565_,data_stage_1__4564_,
  data_stage_1__4563_,data_stage_1__4562_,data_stage_1__4561_,data_stage_1__4560_,
  data_stage_1__4559_,data_stage_1__4558_,data_stage_1__4557_,data_stage_1__4556_,
  data_stage_1__4555_,data_stage_1__4554_,data_stage_1__4553_,data_stage_1__4552_,
  data_stage_1__4551_,data_stage_1__4550_,data_stage_1__4549_,data_stage_1__4548_,
  data_stage_1__4547_,data_stage_1__4546_,data_stage_1__4545_,data_stage_1__4544_,
  data_stage_1__4543_,data_stage_1__4542_,data_stage_1__4541_,data_stage_1__4540_,
  data_stage_1__4539_,data_stage_1__4538_,data_stage_1__4537_,data_stage_1__4536_,
  data_stage_1__4535_,data_stage_1__4534_,data_stage_1__4533_,data_stage_1__4532_,
  data_stage_1__4531_,data_stage_1__4530_,data_stage_1__4529_,data_stage_1__4528_,
  data_stage_1__4527_,data_stage_1__4526_,data_stage_1__4525_,data_stage_1__4524_,
  data_stage_1__4523_,data_stage_1__4522_,data_stage_1__4521_,data_stage_1__4520_,
  data_stage_1__4519_,data_stage_1__4518_,data_stage_1__4517_,data_stage_1__4516_,
  data_stage_1__4515_,data_stage_1__4514_,data_stage_1__4513_,data_stage_1__4512_,
  data_stage_1__4511_,data_stage_1__4510_,data_stage_1__4509_,data_stage_1__4508_,
  data_stage_1__4507_,data_stage_1__4506_,data_stage_1__4505_,data_stage_1__4504_,
  data_stage_1__4503_,data_stage_1__4502_,data_stage_1__4501_,data_stage_1__4500_,
  data_stage_1__4499_,data_stage_1__4498_,data_stage_1__4497_,data_stage_1__4496_,
  data_stage_1__4495_,data_stage_1__4494_,data_stage_1__4493_,data_stage_1__4492_,
  data_stage_1__4491_,data_stage_1__4490_,data_stage_1__4489_,data_stage_1__4488_,
  data_stage_1__4487_,data_stage_1__4486_,data_stage_1__4485_,data_stage_1__4484_,
  data_stage_1__4483_,data_stage_1__4482_,data_stage_1__4481_,data_stage_1__4480_,
  data_stage_1__4479_,data_stage_1__4478_,data_stage_1__4477_,data_stage_1__4476_,
  data_stage_1__4475_,data_stage_1__4474_,data_stage_1__4473_,data_stage_1__4472_,
  data_stage_1__4471_,data_stage_1__4470_,data_stage_1__4469_,data_stage_1__4468_,
  data_stage_1__4467_,data_stage_1__4466_,data_stage_1__4465_,data_stage_1__4464_,
  data_stage_1__4463_,data_stage_1__4462_,data_stage_1__4461_,data_stage_1__4460_,
  data_stage_1__4459_,data_stage_1__4458_,data_stage_1__4457_,data_stage_1__4456_,
  data_stage_1__4455_,data_stage_1__4454_,data_stage_1__4453_,data_stage_1__4452_,
  data_stage_1__4451_,data_stage_1__4450_,data_stage_1__4449_,data_stage_1__4448_,
  data_stage_1__4447_,data_stage_1__4446_,data_stage_1__4445_,data_stage_1__4444_,
  data_stage_1__4443_,data_stage_1__4442_,data_stage_1__4441_,data_stage_1__4440_,
  data_stage_1__4439_,data_stage_1__4438_,data_stage_1__4437_,data_stage_1__4436_,
  data_stage_1__4435_,data_stage_1__4434_,data_stage_1__4433_,data_stage_1__4432_,
  data_stage_1__4431_,data_stage_1__4430_,data_stage_1__4429_,data_stage_1__4428_,
  data_stage_1__4427_,data_stage_1__4426_,data_stage_1__4425_,data_stage_1__4424_,
  data_stage_1__4423_,data_stage_1__4422_,data_stage_1__4421_,data_stage_1__4420_,
  data_stage_1__4419_,data_stage_1__4418_,data_stage_1__4417_,data_stage_1__4416_,
  data_stage_1__4415_,data_stage_1__4414_,data_stage_1__4413_,data_stage_1__4412_,
  data_stage_1__4411_,data_stage_1__4410_,data_stage_1__4409_,data_stage_1__4408_,
  data_stage_1__4407_,data_stage_1__4406_,data_stage_1__4405_,data_stage_1__4404_,
  data_stage_1__4403_,data_stage_1__4402_,data_stage_1__4401_,data_stage_1__4400_,
  data_stage_1__4399_,data_stage_1__4398_,data_stage_1__4397_,data_stage_1__4396_,
  data_stage_1__4395_,data_stage_1__4394_,data_stage_1__4393_,data_stage_1__4392_,
  data_stage_1__4391_,data_stage_1__4390_,data_stage_1__4389_,data_stage_1__4388_,
  data_stage_1__4387_,data_stage_1__4386_,data_stage_1__4385_,data_stage_1__4384_,
  data_stage_1__4383_,data_stage_1__4382_,data_stage_1__4381_,data_stage_1__4380_,
  data_stage_1__4379_,data_stage_1__4378_,data_stage_1__4377_,data_stage_1__4376_,
  data_stage_1__4375_,data_stage_1__4374_,data_stage_1__4373_,data_stage_1__4372_,
  data_stage_1__4371_,data_stage_1__4370_,data_stage_1__4369_,data_stage_1__4368_,
  data_stage_1__4367_,data_stage_1__4366_,data_stage_1__4365_,data_stage_1__4364_,
  data_stage_1__4363_,data_stage_1__4362_,data_stage_1__4361_,data_stage_1__4360_,
  data_stage_1__4359_,data_stage_1__4358_,data_stage_1__4357_,data_stage_1__4356_,
  data_stage_1__4355_,data_stage_1__4354_,data_stage_1__4353_,data_stage_1__4352_,
  data_stage_1__4351_,data_stage_1__4350_,data_stage_1__4349_,data_stage_1__4348_,
  data_stage_1__4347_,data_stage_1__4346_,data_stage_1__4345_,data_stage_1__4344_,
  data_stage_1__4343_,data_stage_1__4342_,data_stage_1__4341_,data_stage_1__4340_,
  data_stage_1__4339_,data_stage_1__4338_,data_stage_1__4337_,data_stage_1__4336_,
  data_stage_1__4335_,data_stage_1__4334_,data_stage_1__4333_,data_stage_1__4332_,
  data_stage_1__4331_,data_stage_1__4330_,data_stage_1__4329_,data_stage_1__4328_,
  data_stage_1__4327_,data_stage_1__4326_,data_stage_1__4325_,data_stage_1__4324_,
  data_stage_1__4323_,data_stage_1__4322_,data_stage_1__4321_,data_stage_1__4320_,
  data_stage_1__4319_,data_stage_1__4318_,data_stage_1__4317_,data_stage_1__4316_,
  data_stage_1__4315_,data_stage_1__4314_,data_stage_1__4313_,data_stage_1__4312_,
  data_stage_1__4311_,data_stage_1__4310_,data_stage_1__4309_,data_stage_1__4308_,
  data_stage_1__4307_,data_stage_1__4306_,data_stage_1__4305_,data_stage_1__4304_,
  data_stage_1__4303_,data_stage_1__4302_,data_stage_1__4301_,data_stage_1__4300_,
  data_stage_1__4299_,data_stage_1__4298_,data_stage_1__4297_,data_stage_1__4296_,
  data_stage_1__4295_,data_stage_1__4294_,data_stage_1__4293_,data_stage_1__4292_,
  data_stage_1__4291_,data_stage_1__4290_,data_stage_1__4289_,data_stage_1__4288_,
  data_stage_1__4287_,data_stage_1__4286_,data_stage_1__4285_,data_stage_1__4284_,
  data_stage_1__4283_,data_stage_1__4282_,data_stage_1__4281_,data_stage_1__4280_,
  data_stage_1__4279_,data_stage_1__4278_,data_stage_1__4277_,data_stage_1__4276_,
  data_stage_1__4275_,data_stage_1__4274_,data_stage_1__4273_,data_stage_1__4272_,
  data_stage_1__4271_,data_stage_1__4270_,data_stage_1__4269_,data_stage_1__4268_,
  data_stage_1__4267_,data_stage_1__4266_,data_stage_1__4265_,data_stage_1__4264_,
  data_stage_1__4263_,data_stage_1__4262_,data_stage_1__4261_,data_stage_1__4260_,
  data_stage_1__4259_,data_stage_1__4258_,data_stage_1__4257_,data_stage_1__4256_,
  data_stage_1__4255_,data_stage_1__4254_,data_stage_1__4253_,data_stage_1__4252_,
  data_stage_1__4251_,data_stage_1__4250_,data_stage_1__4249_,data_stage_1__4248_,
  data_stage_1__4247_,data_stage_1__4246_,data_stage_1__4245_,data_stage_1__4244_,
  data_stage_1__4243_,data_stage_1__4242_,data_stage_1__4241_,data_stage_1__4240_,
  data_stage_1__4239_,data_stage_1__4238_,data_stage_1__4237_,data_stage_1__4236_,
  data_stage_1__4235_,data_stage_1__4234_,data_stage_1__4233_,data_stage_1__4232_,
  data_stage_1__4231_,data_stage_1__4230_,data_stage_1__4229_,data_stage_1__4228_,
  data_stage_1__4227_,data_stage_1__4226_,data_stage_1__4225_,data_stage_1__4224_,
  data_stage_1__4223_,data_stage_1__4222_,data_stage_1__4221_,data_stage_1__4220_,
  data_stage_1__4219_,data_stage_1__4218_,data_stage_1__4217_,data_stage_1__4216_,
  data_stage_1__4215_,data_stage_1__4214_,data_stage_1__4213_,data_stage_1__4212_,
  data_stage_1__4211_,data_stage_1__4210_,data_stage_1__4209_,data_stage_1__4208_,
  data_stage_1__4207_,data_stage_1__4206_,data_stage_1__4205_,data_stage_1__4204_,
  data_stage_1__4203_,data_stage_1__4202_,data_stage_1__4201_,data_stage_1__4200_,
  data_stage_1__4199_,data_stage_1__4198_,data_stage_1__4197_,data_stage_1__4196_,
  data_stage_1__4195_,data_stage_1__4194_,data_stage_1__4193_,data_stage_1__4192_,
  data_stage_1__4191_,data_stage_1__4190_,data_stage_1__4189_,data_stage_1__4188_,
  data_stage_1__4187_,data_stage_1__4186_,data_stage_1__4185_,data_stage_1__4184_,
  data_stage_1__4183_,data_stage_1__4182_,data_stage_1__4181_,data_stage_1__4180_,
  data_stage_1__4179_,data_stage_1__4178_,data_stage_1__4177_,data_stage_1__4176_,
  data_stage_1__4175_,data_stage_1__4174_,data_stage_1__4173_,data_stage_1__4172_,
  data_stage_1__4171_,data_stage_1__4170_,data_stage_1__4169_,data_stage_1__4168_,
  data_stage_1__4167_,data_stage_1__4166_,data_stage_1__4165_,data_stage_1__4164_,
  data_stage_1__4163_,data_stage_1__4162_,data_stage_1__4161_,data_stage_1__4160_,
  data_stage_1__4159_,data_stage_1__4158_,data_stage_1__4157_,data_stage_1__4156_,
  data_stage_1__4155_,data_stage_1__4154_,data_stage_1__4153_,data_stage_1__4152_,
  data_stage_1__4151_,data_stage_1__4150_,data_stage_1__4149_,data_stage_1__4148_,
  data_stage_1__4147_,data_stage_1__4146_,data_stage_1__4145_,data_stage_1__4144_,
  data_stage_1__4143_,data_stage_1__4142_,data_stage_1__4141_,data_stage_1__4140_,
  data_stage_1__4139_,data_stage_1__4138_,data_stage_1__4137_,data_stage_1__4136_,
  data_stage_1__4135_,data_stage_1__4134_,data_stage_1__4133_,data_stage_1__4132_,
  data_stage_1__4131_,data_stage_1__4130_,data_stage_1__4129_,data_stage_1__4128_,
  data_stage_1__4127_,data_stage_1__4126_,data_stage_1__4125_,data_stage_1__4124_,
  data_stage_1__4123_,data_stage_1__4122_,data_stage_1__4121_,data_stage_1__4120_,
  data_stage_1__4119_,data_stage_1__4118_,data_stage_1__4117_,data_stage_1__4116_,
  data_stage_1__4115_,data_stage_1__4114_,data_stage_1__4113_,data_stage_1__4112_,
  data_stage_1__4111_,data_stage_1__4110_,data_stage_1__4109_,data_stage_1__4108_,
  data_stage_1__4107_,data_stage_1__4106_,data_stage_1__4105_,data_stage_1__4104_,
  data_stage_1__4103_,data_stage_1__4102_,data_stage_1__4101_,data_stage_1__4100_,
  data_stage_1__4099_,data_stage_1__4098_,data_stage_1__4097_,data_stage_1__4096_,
  data_stage_1__4095_,data_stage_1__4094_,data_stage_1__4093_,data_stage_1__4092_,
  data_stage_1__4091_,data_stage_1__4090_,data_stage_1__4089_,data_stage_1__4088_,
  data_stage_1__4087_,data_stage_1__4086_,data_stage_1__4085_,data_stage_1__4084_,
  data_stage_1__4083_,data_stage_1__4082_,data_stage_1__4081_,data_stage_1__4080_,
  data_stage_1__4079_,data_stage_1__4078_,data_stage_1__4077_,data_stage_1__4076_,
  data_stage_1__4075_,data_stage_1__4074_,data_stage_1__4073_,data_stage_1__4072_,
  data_stage_1__4071_,data_stage_1__4070_,data_stage_1__4069_,data_stage_1__4068_,
  data_stage_1__4067_,data_stage_1__4066_,data_stage_1__4065_,data_stage_1__4064_,
  data_stage_1__4063_,data_stage_1__4062_,data_stage_1__4061_,data_stage_1__4060_,
  data_stage_1__4059_,data_stage_1__4058_,data_stage_1__4057_,data_stage_1__4056_,
  data_stage_1__4055_,data_stage_1__4054_,data_stage_1__4053_,data_stage_1__4052_,
  data_stage_1__4051_,data_stage_1__4050_,data_stage_1__4049_,data_stage_1__4048_,
  data_stage_1__4047_,data_stage_1__4046_,data_stage_1__4045_,data_stage_1__4044_,
  data_stage_1__4043_,data_stage_1__4042_,data_stage_1__4041_,data_stage_1__4040_,
  data_stage_1__4039_,data_stage_1__4038_,data_stage_1__4037_,data_stage_1__4036_,
  data_stage_1__4035_,data_stage_1__4034_,data_stage_1__4033_,data_stage_1__4032_,
  data_stage_1__4031_,data_stage_1__4030_,data_stage_1__4029_,data_stage_1__4028_,
  data_stage_1__4027_,data_stage_1__4026_,data_stage_1__4025_,data_stage_1__4024_,
  data_stage_1__4023_,data_stage_1__4022_,data_stage_1__4021_,data_stage_1__4020_,
  data_stage_1__4019_,data_stage_1__4018_,data_stage_1__4017_,data_stage_1__4016_,
  data_stage_1__4015_,data_stage_1__4014_,data_stage_1__4013_,data_stage_1__4012_,
  data_stage_1__4011_,data_stage_1__4010_,data_stage_1__4009_,data_stage_1__4008_,
  data_stage_1__4007_,data_stage_1__4006_,data_stage_1__4005_,data_stage_1__4004_,
  data_stage_1__4003_,data_stage_1__4002_,data_stage_1__4001_,data_stage_1__4000_,
  data_stage_1__3999_,data_stage_1__3998_,data_stage_1__3997_,data_stage_1__3996_,
  data_stage_1__3995_,data_stage_1__3994_,data_stage_1__3993_,data_stage_1__3992_,
  data_stage_1__3991_,data_stage_1__3990_,data_stage_1__3989_,data_stage_1__3988_,
  data_stage_1__3987_,data_stage_1__3986_,data_stage_1__3985_,data_stage_1__3984_,
  data_stage_1__3983_,data_stage_1__3982_,data_stage_1__3981_,data_stage_1__3980_,
  data_stage_1__3979_,data_stage_1__3978_,data_stage_1__3977_,data_stage_1__3976_,
  data_stage_1__3975_,data_stage_1__3974_,data_stage_1__3973_,data_stage_1__3972_,
  data_stage_1__3971_,data_stage_1__3970_,data_stage_1__3969_,data_stage_1__3968_,
  data_stage_1__3967_,data_stage_1__3966_,data_stage_1__3965_,data_stage_1__3964_,
  data_stage_1__3963_,data_stage_1__3962_,data_stage_1__3961_,data_stage_1__3960_,
  data_stage_1__3959_,data_stage_1__3958_,data_stage_1__3957_,data_stage_1__3956_,
  data_stage_1__3955_,data_stage_1__3954_,data_stage_1__3953_,data_stage_1__3952_,
  data_stage_1__3951_,data_stage_1__3950_,data_stage_1__3949_,data_stage_1__3948_,
  data_stage_1__3947_,data_stage_1__3946_,data_stage_1__3945_,data_stage_1__3944_,
  data_stage_1__3943_,data_stage_1__3942_,data_stage_1__3941_,data_stage_1__3940_,
  data_stage_1__3939_,data_stage_1__3938_,data_stage_1__3937_,data_stage_1__3936_,
  data_stage_1__3935_,data_stage_1__3934_,data_stage_1__3933_,data_stage_1__3932_,
  data_stage_1__3931_,data_stage_1__3930_,data_stage_1__3929_,data_stage_1__3928_,
  data_stage_1__3927_,data_stage_1__3926_,data_stage_1__3925_,data_stage_1__3924_,
  data_stage_1__3923_,data_stage_1__3922_,data_stage_1__3921_,data_stage_1__3920_,
  data_stage_1__3919_,data_stage_1__3918_,data_stage_1__3917_,data_stage_1__3916_,
  data_stage_1__3915_,data_stage_1__3914_,data_stage_1__3913_,data_stage_1__3912_,
  data_stage_1__3911_,data_stage_1__3910_,data_stage_1__3909_,data_stage_1__3908_,
  data_stage_1__3907_,data_stage_1__3906_,data_stage_1__3905_,data_stage_1__3904_,
  data_stage_1__3903_,data_stage_1__3902_,data_stage_1__3901_,data_stage_1__3900_,
  data_stage_1__3899_,data_stage_1__3898_,data_stage_1__3897_,data_stage_1__3896_,
  data_stage_1__3895_,data_stage_1__3894_,data_stage_1__3893_,data_stage_1__3892_,
  data_stage_1__3891_,data_stage_1__3890_,data_stage_1__3889_,data_stage_1__3888_,
  data_stage_1__3887_,data_stage_1__3886_,data_stage_1__3885_,data_stage_1__3884_,
  data_stage_1__3883_,data_stage_1__3882_,data_stage_1__3881_,data_stage_1__3880_,
  data_stage_1__3879_,data_stage_1__3878_,data_stage_1__3877_,data_stage_1__3876_,
  data_stage_1__3875_,data_stage_1__3874_,data_stage_1__3873_,data_stage_1__3872_,
  data_stage_1__3871_,data_stage_1__3870_,data_stage_1__3869_,data_stage_1__3868_,
  data_stage_1__3867_,data_stage_1__3866_,data_stage_1__3865_,data_stage_1__3864_,
  data_stage_1__3863_,data_stage_1__3862_,data_stage_1__3861_,data_stage_1__3860_,
  data_stage_1__3859_,data_stage_1__3858_,data_stage_1__3857_,data_stage_1__3856_,
  data_stage_1__3855_,data_stage_1__3854_,data_stage_1__3853_,data_stage_1__3852_,
  data_stage_1__3851_,data_stage_1__3850_,data_stage_1__3849_,data_stage_1__3848_,
  data_stage_1__3847_,data_stage_1__3846_,data_stage_1__3845_,data_stage_1__3844_,
  data_stage_1__3843_,data_stage_1__3842_,data_stage_1__3841_,data_stage_1__3840_,
  data_stage_1__3839_,data_stage_1__3838_,data_stage_1__3837_,data_stage_1__3836_,
  data_stage_1__3835_,data_stage_1__3834_,data_stage_1__3833_,data_stage_1__3832_,
  data_stage_1__3831_,data_stage_1__3830_,data_stage_1__3829_,data_stage_1__3828_,
  data_stage_1__3827_,data_stage_1__3826_,data_stage_1__3825_,data_stage_1__3824_,
  data_stage_1__3823_,data_stage_1__3822_,data_stage_1__3821_,data_stage_1__3820_,
  data_stage_1__3819_,data_stage_1__3818_,data_stage_1__3817_,data_stage_1__3816_,
  data_stage_1__3815_,data_stage_1__3814_,data_stage_1__3813_,data_stage_1__3812_,
  data_stage_1__3811_,data_stage_1__3810_,data_stage_1__3809_,data_stage_1__3808_,
  data_stage_1__3807_,data_stage_1__3806_,data_stage_1__3805_,data_stage_1__3804_,
  data_stage_1__3803_,data_stage_1__3802_,data_stage_1__3801_,data_stage_1__3800_,
  data_stage_1__3799_,data_stage_1__3798_,data_stage_1__3797_,data_stage_1__3796_,
  data_stage_1__3795_,data_stage_1__3794_,data_stage_1__3793_,data_stage_1__3792_,
  data_stage_1__3791_,data_stage_1__3790_,data_stage_1__3789_,data_stage_1__3788_,
  data_stage_1__3787_,data_stage_1__3786_,data_stage_1__3785_,data_stage_1__3784_,
  data_stage_1__3783_,data_stage_1__3782_,data_stage_1__3781_,data_stage_1__3780_,
  data_stage_1__3779_,data_stage_1__3778_,data_stage_1__3777_,data_stage_1__3776_,
  data_stage_1__3775_,data_stage_1__3774_,data_stage_1__3773_,data_stage_1__3772_,
  data_stage_1__3771_,data_stage_1__3770_,data_stage_1__3769_,data_stage_1__3768_,
  data_stage_1__3767_,data_stage_1__3766_,data_stage_1__3765_,data_stage_1__3764_,
  data_stage_1__3763_,data_stage_1__3762_,data_stage_1__3761_,data_stage_1__3760_,
  data_stage_1__3759_,data_stage_1__3758_,data_stage_1__3757_,data_stage_1__3756_,
  data_stage_1__3755_,data_stage_1__3754_,data_stage_1__3753_,data_stage_1__3752_,
  data_stage_1__3751_,data_stage_1__3750_,data_stage_1__3749_,data_stage_1__3748_,
  data_stage_1__3747_,data_stage_1__3746_,data_stage_1__3745_,data_stage_1__3744_,
  data_stage_1__3743_,data_stage_1__3742_,data_stage_1__3741_,data_stage_1__3740_,
  data_stage_1__3739_,data_stage_1__3738_,data_stage_1__3737_,data_stage_1__3736_,
  data_stage_1__3735_,data_stage_1__3734_,data_stage_1__3733_,data_stage_1__3732_,
  data_stage_1__3731_,data_stage_1__3730_,data_stage_1__3729_,data_stage_1__3728_,
  data_stage_1__3727_,data_stage_1__3726_,data_stage_1__3725_,data_stage_1__3724_,
  data_stage_1__3723_,data_stage_1__3722_,data_stage_1__3721_,data_stage_1__3720_,
  data_stage_1__3719_,data_stage_1__3718_,data_stage_1__3717_,data_stage_1__3716_,
  data_stage_1__3715_,data_stage_1__3714_,data_stage_1__3713_,data_stage_1__3712_,
  data_stage_1__3711_,data_stage_1__3710_,data_stage_1__3709_,data_stage_1__3708_,
  data_stage_1__3707_,data_stage_1__3706_,data_stage_1__3705_,data_stage_1__3704_,
  data_stage_1__3703_,data_stage_1__3702_,data_stage_1__3701_,data_stage_1__3700_,
  data_stage_1__3699_,data_stage_1__3698_,data_stage_1__3697_,data_stage_1__3696_,
  data_stage_1__3695_,data_stage_1__3694_,data_stage_1__3693_,data_stage_1__3692_,
  data_stage_1__3691_,data_stage_1__3690_,data_stage_1__3689_,data_stage_1__3688_,
  data_stage_1__3687_,data_stage_1__3686_,data_stage_1__3685_,data_stage_1__3684_,
  data_stage_1__3683_,data_stage_1__3682_,data_stage_1__3681_,data_stage_1__3680_,
  data_stage_1__3679_,data_stage_1__3678_,data_stage_1__3677_,data_stage_1__3676_,
  data_stage_1__3675_,data_stage_1__3674_,data_stage_1__3673_,data_stage_1__3672_,
  data_stage_1__3671_,data_stage_1__3670_,data_stage_1__3669_,data_stage_1__3668_,
  data_stage_1__3667_,data_stage_1__3666_,data_stage_1__3665_,data_stage_1__3664_,
  data_stage_1__3663_,data_stage_1__3662_,data_stage_1__3661_,data_stage_1__3660_,
  data_stage_1__3659_,data_stage_1__3658_,data_stage_1__3657_,data_stage_1__3656_,
  data_stage_1__3655_,data_stage_1__3654_,data_stage_1__3653_,data_stage_1__3652_,
  data_stage_1__3651_,data_stage_1__3650_,data_stage_1__3649_,data_stage_1__3648_,
  data_stage_1__3647_,data_stage_1__3646_,data_stage_1__3645_,data_stage_1__3644_,
  data_stage_1__3643_,data_stage_1__3642_,data_stage_1__3641_,data_stage_1__3640_,
  data_stage_1__3639_,data_stage_1__3638_,data_stage_1__3637_,data_stage_1__3636_,
  data_stage_1__3635_,data_stage_1__3634_,data_stage_1__3633_,data_stage_1__3632_,
  data_stage_1__3631_,data_stage_1__3630_,data_stage_1__3629_,data_stage_1__3628_,
  data_stage_1__3627_,data_stage_1__3626_,data_stage_1__3625_,data_stage_1__3624_,
  data_stage_1__3623_,data_stage_1__3622_,data_stage_1__3621_,data_stage_1__3620_,
  data_stage_1__3619_,data_stage_1__3618_,data_stage_1__3617_,data_stage_1__3616_,
  data_stage_1__3615_,data_stage_1__3614_,data_stage_1__3613_,data_stage_1__3612_,
  data_stage_1__3611_,data_stage_1__3610_,data_stage_1__3609_,data_stage_1__3608_,
  data_stage_1__3607_,data_stage_1__3606_,data_stage_1__3605_,data_stage_1__3604_,
  data_stage_1__3603_,data_stage_1__3602_,data_stage_1__3601_,data_stage_1__3600_,
  data_stage_1__3599_,data_stage_1__3598_,data_stage_1__3597_,data_stage_1__3596_,
  data_stage_1__3595_,data_stage_1__3594_,data_stage_1__3593_,data_stage_1__3592_,
  data_stage_1__3591_,data_stage_1__3590_,data_stage_1__3589_,data_stage_1__3588_,
  data_stage_1__3587_,data_stage_1__3586_,data_stage_1__3585_,data_stage_1__3584_,
  data_stage_1__3583_,data_stage_1__3582_,data_stage_1__3581_,data_stage_1__3580_,
  data_stage_1__3579_,data_stage_1__3578_,data_stage_1__3577_,data_stage_1__3576_,
  data_stage_1__3575_,data_stage_1__3574_,data_stage_1__3573_,data_stage_1__3572_,
  data_stage_1__3571_,data_stage_1__3570_,data_stage_1__3569_,data_stage_1__3568_,
  data_stage_1__3567_,data_stage_1__3566_,data_stage_1__3565_,data_stage_1__3564_,
  data_stage_1__3563_,data_stage_1__3562_,data_stage_1__3561_,data_stage_1__3560_,
  data_stage_1__3559_,data_stage_1__3558_,data_stage_1__3557_,data_stage_1__3556_,
  data_stage_1__3555_,data_stage_1__3554_,data_stage_1__3553_,data_stage_1__3552_,
  data_stage_1__3551_,data_stage_1__3550_,data_stage_1__3549_,data_stage_1__3548_,
  data_stage_1__3547_,data_stage_1__3546_,data_stage_1__3545_,data_stage_1__3544_,
  data_stage_1__3543_,data_stage_1__3542_,data_stage_1__3541_,data_stage_1__3540_,
  data_stage_1__3539_,data_stage_1__3538_,data_stage_1__3537_,data_stage_1__3536_,
  data_stage_1__3535_,data_stage_1__3534_,data_stage_1__3533_,data_stage_1__3532_,
  data_stage_1__3531_,data_stage_1__3530_,data_stage_1__3529_,data_stage_1__3528_,
  data_stage_1__3527_,data_stage_1__3526_,data_stage_1__3525_,data_stage_1__3524_,
  data_stage_1__3523_,data_stage_1__3522_,data_stage_1__3521_,data_stage_1__3520_,
  data_stage_1__3519_,data_stage_1__3518_,data_stage_1__3517_,data_stage_1__3516_,
  data_stage_1__3515_,data_stage_1__3514_,data_stage_1__3513_,data_stage_1__3512_,
  data_stage_1__3511_,data_stage_1__3510_,data_stage_1__3509_,data_stage_1__3508_,
  data_stage_1__3507_,data_stage_1__3506_,data_stage_1__3505_,data_stage_1__3504_,
  data_stage_1__3503_,data_stage_1__3502_,data_stage_1__3501_,data_stage_1__3500_,
  data_stage_1__3499_,data_stage_1__3498_,data_stage_1__3497_,data_stage_1__3496_,
  data_stage_1__3495_,data_stage_1__3494_,data_stage_1__3493_,data_stage_1__3492_,
  data_stage_1__3491_,data_stage_1__3490_,data_stage_1__3489_,data_stage_1__3488_,
  data_stage_1__3487_,data_stage_1__3486_,data_stage_1__3485_,data_stage_1__3484_,
  data_stage_1__3483_,data_stage_1__3482_,data_stage_1__3481_,data_stage_1__3480_,
  data_stage_1__3479_,data_stage_1__3478_,data_stage_1__3477_,data_stage_1__3476_,
  data_stage_1__3475_,data_stage_1__3474_,data_stage_1__3473_,data_stage_1__3472_,
  data_stage_1__3471_,data_stage_1__3470_,data_stage_1__3469_,data_stage_1__3468_,
  data_stage_1__3467_,data_stage_1__3466_,data_stage_1__3465_,data_stage_1__3464_,
  data_stage_1__3463_,data_stage_1__3462_,data_stage_1__3461_,data_stage_1__3460_,
  data_stage_1__3459_,data_stage_1__3458_,data_stage_1__3457_,data_stage_1__3456_,
  data_stage_1__3455_,data_stage_1__3454_,data_stage_1__3453_,data_stage_1__3452_,
  data_stage_1__3451_,data_stage_1__3450_,data_stage_1__3449_,data_stage_1__3448_,
  data_stage_1__3447_,data_stage_1__3446_,data_stage_1__3445_,data_stage_1__3444_,
  data_stage_1__3443_,data_stage_1__3442_,data_stage_1__3441_,data_stage_1__3440_,
  data_stage_1__3439_,data_stage_1__3438_,data_stage_1__3437_,data_stage_1__3436_,
  data_stage_1__3435_,data_stage_1__3434_,data_stage_1__3433_,data_stage_1__3432_,
  data_stage_1__3431_,data_stage_1__3430_,data_stage_1__3429_,data_stage_1__3428_,
  data_stage_1__3427_,data_stage_1__3426_,data_stage_1__3425_,data_stage_1__3424_,
  data_stage_1__3423_,data_stage_1__3422_,data_stage_1__3421_,data_stage_1__3420_,
  data_stage_1__3419_,data_stage_1__3418_,data_stage_1__3417_,data_stage_1__3416_,
  data_stage_1__3415_,data_stage_1__3414_,data_stage_1__3413_,data_stage_1__3412_,
  data_stage_1__3411_,data_stage_1__3410_,data_stage_1__3409_,data_stage_1__3408_,
  data_stage_1__3407_,data_stage_1__3406_,data_stage_1__3405_,data_stage_1__3404_,
  data_stage_1__3403_,data_stage_1__3402_,data_stage_1__3401_,data_stage_1__3400_,
  data_stage_1__3399_,data_stage_1__3398_,data_stage_1__3397_,data_stage_1__3396_,
  data_stage_1__3395_,data_stage_1__3394_,data_stage_1__3393_,data_stage_1__3392_,
  data_stage_1__3391_,data_stage_1__3390_,data_stage_1__3389_,data_stage_1__3388_,
  data_stage_1__3387_,data_stage_1__3386_,data_stage_1__3385_,data_stage_1__3384_,
  data_stage_1__3383_,data_stage_1__3382_,data_stage_1__3381_,data_stage_1__3380_,
  data_stage_1__3379_,data_stage_1__3378_,data_stage_1__3377_,data_stage_1__3376_,
  data_stage_1__3375_,data_stage_1__3374_,data_stage_1__3373_,data_stage_1__3372_,
  data_stage_1__3371_,data_stage_1__3370_,data_stage_1__3369_,data_stage_1__3368_,
  data_stage_1__3367_,data_stage_1__3366_,data_stage_1__3365_,data_stage_1__3364_,
  data_stage_1__3363_,data_stage_1__3362_,data_stage_1__3361_,data_stage_1__3360_,
  data_stage_1__3359_,data_stage_1__3358_,data_stage_1__3357_,data_stage_1__3356_,
  data_stage_1__3355_,data_stage_1__3354_,data_stage_1__3353_,data_stage_1__3352_,
  data_stage_1__3351_,data_stage_1__3350_,data_stage_1__3349_,data_stage_1__3348_,
  data_stage_1__3347_,data_stage_1__3346_,data_stage_1__3345_,data_stage_1__3344_,
  data_stage_1__3343_,data_stage_1__3342_,data_stage_1__3341_,data_stage_1__3340_,
  data_stage_1__3339_,data_stage_1__3338_,data_stage_1__3337_,data_stage_1__3336_,
  data_stage_1__3335_,data_stage_1__3334_,data_stage_1__3333_,data_stage_1__3332_,
  data_stage_1__3331_,data_stage_1__3330_,data_stage_1__3329_,data_stage_1__3328_,
  data_stage_1__3327_,data_stage_1__3326_,data_stage_1__3325_,data_stage_1__3324_,
  data_stage_1__3323_,data_stage_1__3322_,data_stage_1__3321_,data_stage_1__3320_,
  data_stage_1__3319_,data_stage_1__3318_,data_stage_1__3317_,data_stage_1__3316_,
  data_stage_1__3315_,data_stage_1__3314_,data_stage_1__3313_,data_stage_1__3312_,
  data_stage_1__3311_,data_stage_1__3310_,data_stage_1__3309_,data_stage_1__3308_,
  data_stage_1__3307_,data_stage_1__3306_,data_stage_1__3305_,data_stage_1__3304_,
  data_stage_1__3303_,data_stage_1__3302_,data_stage_1__3301_,data_stage_1__3300_,
  data_stage_1__3299_,data_stage_1__3298_,data_stage_1__3297_,data_stage_1__3296_,
  data_stage_1__3295_,data_stage_1__3294_,data_stage_1__3293_,data_stage_1__3292_,
  data_stage_1__3291_,data_stage_1__3290_,data_stage_1__3289_,data_stage_1__3288_,
  data_stage_1__3287_,data_stage_1__3286_,data_stage_1__3285_,data_stage_1__3284_,
  data_stage_1__3283_,data_stage_1__3282_,data_stage_1__3281_,data_stage_1__3280_,
  data_stage_1__3279_,data_stage_1__3278_,data_stage_1__3277_,data_stage_1__3276_,
  data_stage_1__3275_,data_stage_1__3274_,data_stage_1__3273_,data_stage_1__3272_,
  data_stage_1__3271_,data_stage_1__3270_,data_stage_1__3269_,data_stage_1__3268_,
  data_stage_1__3267_,data_stage_1__3266_,data_stage_1__3265_,data_stage_1__3264_,
  data_stage_1__3263_,data_stage_1__3262_,data_stage_1__3261_,data_stage_1__3260_,
  data_stage_1__3259_,data_stage_1__3258_,data_stage_1__3257_,data_stage_1__3256_,
  data_stage_1__3255_,data_stage_1__3254_,data_stage_1__3253_,data_stage_1__3252_,
  data_stage_1__3251_,data_stage_1__3250_,data_stage_1__3249_,data_stage_1__3248_,
  data_stage_1__3247_,data_stage_1__3246_,data_stage_1__3245_,data_stage_1__3244_,
  data_stage_1__3243_,data_stage_1__3242_,data_stage_1__3241_,data_stage_1__3240_,
  data_stage_1__3239_,data_stage_1__3238_,data_stage_1__3237_,data_stage_1__3236_,
  data_stage_1__3235_,data_stage_1__3234_,data_stage_1__3233_,data_stage_1__3232_,
  data_stage_1__3231_,data_stage_1__3230_,data_stage_1__3229_,data_stage_1__3228_,
  data_stage_1__3227_,data_stage_1__3226_,data_stage_1__3225_,data_stage_1__3224_,
  data_stage_1__3223_,data_stage_1__3222_,data_stage_1__3221_,data_stage_1__3220_,
  data_stage_1__3219_,data_stage_1__3218_,data_stage_1__3217_,data_stage_1__3216_,
  data_stage_1__3215_,data_stage_1__3214_,data_stage_1__3213_,data_stage_1__3212_,
  data_stage_1__3211_,data_stage_1__3210_,data_stage_1__3209_,data_stage_1__3208_,
  data_stage_1__3207_,data_stage_1__3206_,data_stage_1__3205_,data_stage_1__3204_,
  data_stage_1__3203_,data_stage_1__3202_,data_stage_1__3201_,data_stage_1__3200_,
  data_stage_1__3199_,data_stage_1__3198_,data_stage_1__3197_,data_stage_1__3196_,
  data_stage_1__3195_,data_stage_1__3194_,data_stage_1__3193_,data_stage_1__3192_,
  data_stage_1__3191_,data_stage_1__3190_,data_stage_1__3189_,data_stage_1__3188_,
  data_stage_1__3187_,data_stage_1__3186_,data_stage_1__3185_,data_stage_1__3184_,
  data_stage_1__3183_,data_stage_1__3182_,data_stage_1__3181_,data_stage_1__3180_,
  data_stage_1__3179_,data_stage_1__3178_,data_stage_1__3177_,data_stage_1__3176_,
  data_stage_1__3175_,data_stage_1__3174_,data_stage_1__3173_,data_stage_1__3172_,
  data_stage_1__3171_,data_stage_1__3170_,data_stage_1__3169_,data_stage_1__3168_,
  data_stage_1__3167_,data_stage_1__3166_,data_stage_1__3165_,data_stage_1__3164_,
  data_stage_1__3163_,data_stage_1__3162_,data_stage_1__3161_,data_stage_1__3160_,
  data_stage_1__3159_,data_stage_1__3158_,data_stage_1__3157_,data_stage_1__3156_,
  data_stage_1__3155_,data_stage_1__3154_,data_stage_1__3153_,data_stage_1__3152_,
  data_stage_1__3151_,data_stage_1__3150_,data_stage_1__3149_,data_stage_1__3148_,
  data_stage_1__3147_,data_stage_1__3146_,data_stage_1__3145_,data_stage_1__3144_,
  data_stage_1__3143_,data_stage_1__3142_,data_stage_1__3141_,data_stage_1__3140_,
  data_stage_1__3139_,data_stage_1__3138_,data_stage_1__3137_,data_stage_1__3136_,
  data_stage_1__3135_,data_stage_1__3134_,data_stage_1__3133_,data_stage_1__3132_,
  data_stage_1__3131_,data_stage_1__3130_,data_stage_1__3129_,data_stage_1__3128_,
  data_stage_1__3127_,data_stage_1__3126_,data_stage_1__3125_,data_stage_1__3124_,
  data_stage_1__3123_,data_stage_1__3122_,data_stage_1__3121_,data_stage_1__3120_,
  data_stage_1__3119_,data_stage_1__3118_,data_stage_1__3117_,data_stage_1__3116_,
  data_stage_1__3115_,data_stage_1__3114_,data_stage_1__3113_,data_stage_1__3112_,
  data_stage_1__3111_,data_stage_1__3110_,data_stage_1__3109_,data_stage_1__3108_,
  data_stage_1__3107_,data_stage_1__3106_,data_stage_1__3105_,data_stage_1__3104_,
  data_stage_1__3103_,data_stage_1__3102_,data_stage_1__3101_,data_stage_1__3100_,
  data_stage_1__3099_,data_stage_1__3098_,data_stage_1__3097_,data_stage_1__3096_,
  data_stage_1__3095_,data_stage_1__3094_,data_stage_1__3093_,data_stage_1__3092_,
  data_stage_1__3091_,data_stage_1__3090_,data_stage_1__3089_,data_stage_1__3088_,
  data_stage_1__3087_,data_stage_1__3086_,data_stage_1__3085_,data_stage_1__3084_,
  data_stage_1__3083_,data_stage_1__3082_,data_stage_1__3081_,data_stage_1__3080_,
  data_stage_1__3079_,data_stage_1__3078_,data_stage_1__3077_,data_stage_1__3076_,
  data_stage_1__3075_,data_stage_1__3074_,data_stage_1__3073_,data_stage_1__3072_,
  data_stage_1__3071_,data_stage_1__3070_,data_stage_1__3069_,data_stage_1__3068_,
  data_stage_1__3067_,data_stage_1__3066_,data_stage_1__3065_,data_stage_1__3064_,
  data_stage_1__3063_,data_stage_1__3062_,data_stage_1__3061_,data_stage_1__3060_,
  data_stage_1__3059_,data_stage_1__3058_,data_stage_1__3057_,data_stage_1__3056_,
  data_stage_1__3055_,data_stage_1__3054_,data_stage_1__3053_,data_stage_1__3052_,
  data_stage_1__3051_,data_stage_1__3050_,data_stage_1__3049_,data_stage_1__3048_,
  data_stage_1__3047_,data_stage_1__3046_,data_stage_1__3045_,data_stage_1__3044_,
  data_stage_1__3043_,data_stage_1__3042_,data_stage_1__3041_,data_stage_1__3040_,
  data_stage_1__3039_,data_stage_1__3038_,data_stage_1__3037_,data_stage_1__3036_,
  data_stage_1__3035_,data_stage_1__3034_,data_stage_1__3033_,data_stage_1__3032_,
  data_stage_1__3031_,data_stage_1__3030_,data_stage_1__3029_,data_stage_1__3028_,
  data_stage_1__3027_,data_stage_1__3026_,data_stage_1__3025_,data_stage_1__3024_,
  data_stage_1__3023_,data_stage_1__3022_,data_stage_1__3021_,data_stage_1__3020_,
  data_stage_1__3019_,data_stage_1__3018_,data_stage_1__3017_,data_stage_1__3016_,
  data_stage_1__3015_,data_stage_1__3014_,data_stage_1__3013_,data_stage_1__3012_,
  data_stage_1__3011_,data_stage_1__3010_,data_stage_1__3009_,data_stage_1__3008_,
  data_stage_1__3007_,data_stage_1__3006_,data_stage_1__3005_,data_stage_1__3004_,
  data_stage_1__3003_,data_stage_1__3002_,data_stage_1__3001_,data_stage_1__3000_,
  data_stage_1__2999_,data_stage_1__2998_,data_stage_1__2997_,data_stage_1__2996_,
  data_stage_1__2995_,data_stage_1__2994_,data_stage_1__2993_,data_stage_1__2992_,
  data_stage_1__2991_,data_stage_1__2990_,data_stage_1__2989_,data_stage_1__2988_,
  data_stage_1__2987_,data_stage_1__2986_,data_stage_1__2985_,data_stage_1__2984_,
  data_stage_1__2983_,data_stage_1__2982_,data_stage_1__2981_,data_stage_1__2980_,
  data_stage_1__2979_,data_stage_1__2978_,data_stage_1__2977_,data_stage_1__2976_,
  data_stage_1__2975_,data_stage_1__2974_,data_stage_1__2973_,data_stage_1__2972_,
  data_stage_1__2971_,data_stage_1__2970_,data_stage_1__2969_,data_stage_1__2968_,
  data_stage_1__2967_,data_stage_1__2966_,data_stage_1__2965_,data_stage_1__2964_,
  data_stage_1__2963_,data_stage_1__2962_,data_stage_1__2961_,data_stage_1__2960_,
  data_stage_1__2959_,data_stage_1__2958_,data_stage_1__2957_,data_stage_1__2956_,
  data_stage_1__2955_,data_stage_1__2954_,data_stage_1__2953_,data_stage_1__2952_,
  data_stage_1__2951_,data_stage_1__2950_,data_stage_1__2949_,data_stage_1__2948_,
  data_stage_1__2947_,data_stage_1__2946_,data_stage_1__2945_,data_stage_1__2944_,
  data_stage_1__2943_,data_stage_1__2942_,data_stage_1__2941_,data_stage_1__2940_,
  data_stage_1__2939_,data_stage_1__2938_,data_stage_1__2937_,data_stage_1__2936_,
  data_stage_1__2935_,data_stage_1__2934_,data_stage_1__2933_,data_stage_1__2932_,
  data_stage_1__2931_,data_stage_1__2930_,data_stage_1__2929_,data_stage_1__2928_,
  data_stage_1__2927_,data_stage_1__2926_,data_stage_1__2925_,data_stage_1__2924_,
  data_stage_1__2923_,data_stage_1__2922_,data_stage_1__2921_,data_stage_1__2920_,
  data_stage_1__2919_,data_stage_1__2918_,data_stage_1__2917_,data_stage_1__2916_,
  data_stage_1__2915_,data_stage_1__2914_,data_stage_1__2913_,data_stage_1__2912_,
  data_stage_1__2911_,data_stage_1__2910_,data_stage_1__2909_,data_stage_1__2908_,
  data_stage_1__2907_,data_stage_1__2906_,data_stage_1__2905_,data_stage_1__2904_,
  data_stage_1__2903_,data_stage_1__2902_,data_stage_1__2901_,data_stage_1__2900_,
  data_stage_1__2899_,data_stage_1__2898_,data_stage_1__2897_,data_stage_1__2896_,
  data_stage_1__2895_,data_stage_1__2894_,data_stage_1__2893_,data_stage_1__2892_,
  data_stage_1__2891_,data_stage_1__2890_,data_stage_1__2889_,data_stage_1__2888_,
  data_stage_1__2887_,data_stage_1__2886_,data_stage_1__2885_,data_stage_1__2884_,
  data_stage_1__2883_,data_stage_1__2882_,data_stage_1__2881_,data_stage_1__2880_,
  data_stage_1__2879_,data_stage_1__2878_,data_stage_1__2877_,data_stage_1__2876_,
  data_stage_1__2875_,data_stage_1__2874_,data_stage_1__2873_,data_stage_1__2872_,
  data_stage_1__2871_,data_stage_1__2870_,data_stage_1__2869_,data_stage_1__2868_,
  data_stage_1__2867_,data_stage_1__2866_,data_stage_1__2865_,data_stage_1__2864_,
  data_stage_1__2863_,data_stage_1__2862_,data_stage_1__2861_,data_stage_1__2860_,
  data_stage_1__2859_,data_stage_1__2858_,data_stage_1__2857_,data_stage_1__2856_,
  data_stage_1__2855_,data_stage_1__2854_,data_stage_1__2853_,data_stage_1__2852_,
  data_stage_1__2851_,data_stage_1__2850_,data_stage_1__2849_,data_stage_1__2848_,
  data_stage_1__2847_,data_stage_1__2846_,data_stage_1__2845_,data_stage_1__2844_,
  data_stage_1__2843_,data_stage_1__2842_,data_stage_1__2841_,data_stage_1__2840_,
  data_stage_1__2839_,data_stage_1__2838_,data_stage_1__2837_,data_stage_1__2836_,
  data_stage_1__2835_,data_stage_1__2834_,data_stage_1__2833_,data_stage_1__2832_,
  data_stage_1__2831_,data_stage_1__2830_,data_stage_1__2829_,data_stage_1__2828_,
  data_stage_1__2827_,data_stage_1__2826_,data_stage_1__2825_,data_stage_1__2824_,
  data_stage_1__2823_,data_stage_1__2822_,data_stage_1__2821_,data_stage_1__2820_,
  data_stage_1__2819_,data_stage_1__2818_,data_stage_1__2817_,data_stage_1__2816_,
  data_stage_1__2815_,data_stage_1__2814_,data_stage_1__2813_,data_stage_1__2812_,
  data_stage_1__2811_,data_stage_1__2810_,data_stage_1__2809_,data_stage_1__2808_,
  data_stage_1__2807_,data_stage_1__2806_,data_stage_1__2805_,data_stage_1__2804_,
  data_stage_1__2803_,data_stage_1__2802_,data_stage_1__2801_,data_stage_1__2800_,
  data_stage_1__2799_,data_stage_1__2798_,data_stage_1__2797_,data_stage_1__2796_,
  data_stage_1__2795_,data_stage_1__2794_,data_stage_1__2793_,data_stage_1__2792_,
  data_stage_1__2791_,data_stage_1__2790_,data_stage_1__2789_,data_stage_1__2788_,
  data_stage_1__2787_,data_stage_1__2786_,data_stage_1__2785_,data_stage_1__2784_,
  data_stage_1__2783_,data_stage_1__2782_,data_stage_1__2781_,data_stage_1__2780_,
  data_stage_1__2779_,data_stage_1__2778_,data_stage_1__2777_,data_stage_1__2776_,
  data_stage_1__2775_,data_stage_1__2774_,data_stage_1__2773_,data_stage_1__2772_,
  data_stage_1__2771_,data_stage_1__2770_,data_stage_1__2769_,data_stage_1__2768_,
  data_stage_1__2767_,data_stage_1__2766_,data_stage_1__2765_,data_stage_1__2764_,
  data_stage_1__2763_,data_stage_1__2762_,data_stage_1__2761_,data_stage_1__2760_,
  data_stage_1__2759_,data_stage_1__2758_,data_stage_1__2757_,data_stage_1__2756_,
  data_stage_1__2755_,data_stage_1__2754_,data_stage_1__2753_,data_stage_1__2752_,
  data_stage_1__2751_,data_stage_1__2750_,data_stage_1__2749_,data_stage_1__2748_,
  data_stage_1__2747_,data_stage_1__2746_,data_stage_1__2745_,data_stage_1__2744_,
  data_stage_1__2743_,data_stage_1__2742_,data_stage_1__2741_,data_stage_1__2740_,
  data_stage_1__2739_,data_stage_1__2738_,data_stage_1__2737_,data_stage_1__2736_,
  data_stage_1__2735_,data_stage_1__2734_,data_stage_1__2733_,data_stage_1__2732_,
  data_stage_1__2731_,data_stage_1__2730_,data_stage_1__2729_,data_stage_1__2728_,
  data_stage_1__2727_,data_stage_1__2726_,data_stage_1__2725_,data_stage_1__2724_,
  data_stage_1__2723_,data_stage_1__2722_,data_stage_1__2721_,data_stage_1__2720_,
  data_stage_1__2719_,data_stage_1__2718_,data_stage_1__2717_,data_stage_1__2716_,
  data_stage_1__2715_,data_stage_1__2714_,data_stage_1__2713_,data_stage_1__2712_,
  data_stage_1__2711_,data_stage_1__2710_,data_stage_1__2709_,data_stage_1__2708_,
  data_stage_1__2707_,data_stage_1__2706_,data_stage_1__2705_,data_stage_1__2704_,
  data_stage_1__2703_,data_stage_1__2702_,data_stage_1__2701_,data_stage_1__2700_,
  data_stage_1__2699_,data_stage_1__2698_,data_stage_1__2697_,data_stage_1__2696_,
  data_stage_1__2695_,data_stage_1__2694_,data_stage_1__2693_,data_stage_1__2692_,
  data_stage_1__2691_,data_stage_1__2690_,data_stage_1__2689_,data_stage_1__2688_,
  data_stage_1__2687_,data_stage_1__2686_,data_stage_1__2685_,data_stage_1__2684_,
  data_stage_1__2683_,data_stage_1__2682_,data_stage_1__2681_,data_stage_1__2680_,
  data_stage_1__2679_,data_stage_1__2678_,data_stage_1__2677_,data_stage_1__2676_,
  data_stage_1__2675_,data_stage_1__2674_,data_stage_1__2673_,data_stage_1__2672_,
  data_stage_1__2671_,data_stage_1__2670_,data_stage_1__2669_,data_stage_1__2668_,
  data_stage_1__2667_,data_stage_1__2666_,data_stage_1__2665_,data_stage_1__2664_,
  data_stage_1__2663_,data_stage_1__2662_,data_stage_1__2661_,data_stage_1__2660_,
  data_stage_1__2659_,data_stage_1__2658_,data_stage_1__2657_,data_stage_1__2656_,
  data_stage_1__2655_,data_stage_1__2654_,data_stage_1__2653_,data_stage_1__2652_,
  data_stage_1__2651_,data_stage_1__2650_,data_stage_1__2649_,data_stage_1__2648_,
  data_stage_1__2647_,data_stage_1__2646_,data_stage_1__2645_,data_stage_1__2644_,
  data_stage_1__2643_,data_stage_1__2642_,data_stage_1__2641_,data_stage_1__2640_,
  data_stage_1__2639_,data_stage_1__2638_,data_stage_1__2637_,data_stage_1__2636_,
  data_stage_1__2635_,data_stage_1__2634_,data_stage_1__2633_,data_stage_1__2632_,
  data_stage_1__2631_,data_stage_1__2630_,data_stage_1__2629_,data_stage_1__2628_,
  data_stage_1__2627_,data_stage_1__2626_,data_stage_1__2625_,data_stage_1__2624_,
  data_stage_1__2623_,data_stage_1__2622_,data_stage_1__2621_,data_stage_1__2620_,
  data_stage_1__2619_,data_stage_1__2618_,data_stage_1__2617_,data_stage_1__2616_,
  data_stage_1__2615_,data_stage_1__2614_,data_stage_1__2613_,data_stage_1__2612_,
  data_stage_1__2611_,data_stage_1__2610_,data_stage_1__2609_,data_stage_1__2608_,
  data_stage_1__2607_,data_stage_1__2606_,data_stage_1__2605_,data_stage_1__2604_,
  data_stage_1__2603_,data_stage_1__2602_,data_stage_1__2601_,data_stage_1__2600_,
  data_stage_1__2599_,data_stage_1__2598_,data_stage_1__2597_,data_stage_1__2596_,
  data_stage_1__2595_,data_stage_1__2594_,data_stage_1__2593_,data_stage_1__2592_,
  data_stage_1__2591_,data_stage_1__2590_,data_stage_1__2589_,data_stage_1__2588_,
  data_stage_1__2587_,data_stage_1__2586_,data_stage_1__2585_,data_stage_1__2584_,
  data_stage_1__2583_,data_stage_1__2582_,data_stage_1__2581_,data_stage_1__2580_,
  data_stage_1__2579_,data_stage_1__2578_,data_stage_1__2577_,data_stage_1__2576_,
  data_stage_1__2575_,data_stage_1__2574_,data_stage_1__2573_,data_stage_1__2572_,
  data_stage_1__2571_,data_stage_1__2570_,data_stage_1__2569_,data_stage_1__2568_,
  data_stage_1__2567_,data_stage_1__2566_,data_stage_1__2565_,data_stage_1__2564_,
  data_stage_1__2563_,data_stage_1__2562_,data_stage_1__2561_,data_stage_1__2560_,
  data_stage_1__2559_,data_stage_1__2558_,data_stage_1__2557_,data_stage_1__2556_,
  data_stage_1__2555_,data_stage_1__2554_,data_stage_1__2553_,data_stage_1__2552_,
  data_stage_1__2551_,data_stage_1__2550_,data_stage_1__2549_,data_stage_1__2548_,
  data_stage_1__2547_,data_stage_1__2546_,data_stage_1__2545_,data_stage_1__2544_,
  data_stage_1__2543_,data_stage_1__2542_,data_stage_1__2541_,data_stage_1__2540_,
  data_stage_1__2539_,data_stage_1__2538_,data_stage_1__2537_,data_stage_1__2536_,
  data_stage_1__2535_,data_stage_1__2534_,data_stage_1__2533_,data_stage_1__2532_,
  data_stage_1__2531_,data_stage_1__2530_,data_stage_1__2529_,data_stage_1__2528_,
  data_stage_1__2527_,data_stage_1__2526_,data_stage_1__2525_,data_stage_1__2524_,
  data_stage_1__2523_,data_stage_1__2522_,data_stage_1__2521_,data_stage_1__2520_,
  data_stage_1__2519_,data_stage_1__2518_,data_stage_1__2517_,data_stage_1__2516_,
  data_stage_1__2515_,data_stage_1__2514_,data_stage_1__2513_,data_stage_1__2512_,
  data_stage_1__2511_,data_stage_1__2510_,data_stage_1__2509_,data_stage_1__2508_,
  data_stage_1__2507_,data_stage_1__2506_,data_stage_1__2505_,data_stage_1__2504_,
  data_stage_1__2503_,data_stage_1__2502_,data_stage_1__2501_,data_stage_1__2500_,
  data_stage_1__2499_,data_stage_1__2498_,data_stage_1__2497_,data_stage_1__2496_,
  data_stage_1__2495_,data_stage_1__2494_,data_stage_1__2493_,data_stage_1__2492_,
  data_stage_1__2491_,data_stage_1__2490_,data_stage_1__2489_,data_stage_1__2488_,
  data_stage_1__2487_,data_stage_1__2486_,data_stage_1__2485_,data_stage_1__2484_,
  data_stage_1__2483_,data_stage_1__2482_,data_stage_1__2481_,data_stage_1__2480_,
  data_stage_1__2479_,data_stage_1__2478_,data_stage_1__2477_,data_stage_1__2476_,
  data_stage_1__2475_,data_stage_1__2474_,data_stage_1__2473_,data_stage_1__2472_,
  data_stage_1__2471_,data_stage_1__2470_,data_stage_1__2469_,data_stage_1__2468_,
  data_stage_1__2467_,data_stage_1__2466_,data_stage_1__2465_,data_stage_1__2464_,
  data_stage_1__2463_,data_stage_1__2462_,data_stage_1__2461_,data_stage_1__2460_,
  data_stage_1__2459_,data_stage_1__2458_,data_stage_1__2457_,data_stage_1__2456_,
  data_stage_1__2455_,data_stage_1__2454_,data_stage_1__2453_,data_stage_1__2452_,
  data_stage_1__2451_,data_stage_1__2450_,data_stage_1__2449_,data_stage_1__2448_,
  data_stage_1__2447_,data_stage_1__2446_,data_stage_1__2445_,data_stage_1__2444_,
  data_stage_1__2443_,data_stage_1__2442_,data_stage_1__2441_,data_stage_1__2440_,
  data_stage_1__2439_,data_stage_1__2438_,data_stage_1__2437_,data_stage_1__2436_,
  data_stage_1__2435_,data_stage_1__2434_,data_stage_1__2433_,data_stage_1__2432_,
  data_stage_1__2431_,data_stage_1__2430_,data_stage_1__2429_,data_stage_1__2428_,
  data_stage_1__2427_,data_stage_1__2426_,data_stage_1__2425_,data_stage_1__2424_,
  data_stage_1__2423_,data_stage_1__2422_,data_stage_1__2421_,data_stage_1__2420_,
  data_stage_1__2419_,data_stage_1__2418_,data_stage_1__2417_,data_stage_1__2416_,
  data_stage_1__2415_,data_stage_1__2414_,data_stage_1__2413_,data_stage_1__2412_,
  data_stage_1__2411_,data_stage_1__2410_,data_stage_1__2409_,data_stage_1__2408_,
  data_stage_1__2407_,data_stage_1__2406_,data_stage_1__2405_,data_stage_1__2404_,
  data_stage_1__2403_,data_stage_1__2402_,data_stage_1__2401_,data_stage_1__2400_,
  data_stage_1__2399_,data_stage_1__2398_,data_stage_1__2397_,data_stage_1__2396_,
  data_stage_1__2395_,data_stage_1__2394_,data_stage_1__2393_,data_stage_1__2392_,
  data_stage_1__2391_,data_stage_1__2390_,data_stage_1__2389_,data_stage_1__2388_,
  data_stage_1__2387_,data_stage_1__2386_,data_stage_1__2385_,data_stage_1__2384_,
  data_stage_1__2383_,data_stage_1__2382_,data_stage_1__2381_,data_stage_1__2380_,
  data_stage_1__2379_,data_stage_1__2378_,data_stage_1__2377_,data_stage_1__2376_,
  data_stage_1__2375_,data_stage_1__2374_,data_stage_1__2373_,data_stage_1__2372_,
  data_stage_1__2371_,data_stage_1__2370_,data_stage_1__2369_,data_stage_1__2368_,
  data_stage_1__2367_,data_stage_1__2366_,data_stage_1__2365_,data_stage_1__2364_,
  data_stage_1__2363_,data_stage_1__2362_,data_stage_1__2361_,data_stage_1__2360_,
  data_stage_1__2359_,data_stage_1__2358_,data_stage_1__2357_,data_stage_1__2356_,
  data_stage_1__2355_,data_stage_1__2354_,data_stage_1__2353_,data_stage_1__2352_,
  data_stage_1__2351_,data_stage_1__2350_,data_stage_1__2349_,data_stage_1__2348_,
  data_stage_1__2347_,data_stage_1__2346_,data_stage_1__2345_,data_stage_1__2344_,
  data_stage_1__2343_,data_stage_1__2342_,data_stage_1__2341_,data_stage_1__2340_,
  data_stage_1__2339_,data_stage_1__2338_,data_stage_1__2337_,data_stage_1__2336_,
  data_stage_1__2335_,data_stage_1__2334_,data_stage_1__2333_,data_stage_1__2332_,
  data_stage_1__2331_,data_stage_1__2330_,data_stage_1__2329_,data_stage_1__2328_,
  data_stage_1__2327_,data_stage_1__2326_,data_stage_1__2325_,data_stage_1__2324_,
  data_stage_1__2323_,data_stage_1__2322_,data_stage_1__2321_,data_stage_1__2320_,
  data_stage_1__2319_,data_stage_1__2318_,data_stage_1__2317_,data_stage_1__2316_,
  data_stage_1__2315_,data_stage_1__2314_,data_stage_1__2313_,data_stage_1__2312_,
  data_stage_1__2311_,data_stage_1__2310_,data_stage_1__2309_,data_stage_1__2308_,
  data_stage_1__2307_,data_stage_1__2306_,data_stage_1__2305_,data_stage_1__2304_,
  data_stage_1__2303_,data_stage_1__2302_,data_stage_1__2301_,data_stage_1__2300_,
  data_stage_1__2299_,data_stage_1__2298_,data_stage_1__2297_,data_stage_1__2296_,
  data_stage_1__2295_,data_stage_1__2294_,data_stage_1__2293_,data_stage_1__2292_,
  data_stage_1__2291_,data_stage_1__2290_,data_stage_1__2289_,data_stage_1__2288_,
  data_stage_1__2287_,data_stage_1__2286_,data_stage_1__2285_,data_stage_1__2284_,
  data_stage_1__2283_,data_stage_1__2282_,data_stage_1__2281_,data_stage_1__2280_,
  data_stage_1__2279_,data_stage_1__2278_,data_stage_1__2277_,data_stage_1__2276_,
  data_stage_1__2275_,data_stage_1__2274_,data_stage_1__2273_,data_stage_1__2272_,
  data_stage_1__2271_,data_stage_1__2270_,data_stage_1__2269_,data_stage_1__2268_,
  data_stage_1__2267_,data_stage_1__2266_,data_stage_1__2265_,data_stage_1__2264_,
  data_stage_1__2263_,data_stage_1__2262_,data_stage_1__2261_,data_stage_1__2260_,
  data_stage_1__2259_,data_stage_1__2258_,data_stage_1__2257_,data_stage_1__2256_,
  data_stage_1__2255_,data_stage_1__2254_,data_stage_1__2253_,data_stage_1__2252_,
  data_stage_1__2251_,data_stage_1__2250_,data_stage_1__2249_,data_stage_1__2248_,
  data_stage_1__2247_,data_stage_1__2246_,data_stage_1__2245_,data_stage_1__2244_,
  data_stage_1__2243_,data_stage_1__2242_,data_stage_1__2241_,data_stage_1__2240_,
  data_stage_1__2239_,data_stage_1__2238_,data_stage_1__2237_,data_stage_1__2236_,
  data_stage_1__2235_,data_stage_1__2234_,data_stage_1__2233_,data_stage_1__2232_,
  data_stage_1__2231_,data_stage_1__2230_,data_stage_1__2229_,data_stage_1__2228_,
  data_stage_1__2227_,data_stage_1__2226_,data_stage_1__2225_,data_stage_1__2224_,
  data_stage_1__2223_,data_stage_1__2222_,data_stage_1__2221_,data_stage_1__2220_,
  data_stage_1__2219_,data_stage_1__2218_,data_stage_1__2217_,data_stage_1__2216_,
  data_stage_1__2215_,data_stage_1__2214_,data_stage_1__2213_,data_stage_1__2212_,
  data_stage_1__2211_,data_stage_1__2210_,data_stage_1__2209_,data_stage_1__2208_,
  data_stage_1__2207_,data_stage_1__2206_,data_stage_1__2205_,data_stage_1__2204_,
  data_stage_1__2203_,data_stage_1__2202_,data_stage_1__2201_,data_stage_1__2200_,
  data_stage_1__2199_,data_stage_1__2198_,data_stage_1__2197_,data_stage_1__2196_,
  data_stage_1__2195_,data_stage_1__2194_,data_stage_1__2193_,data_stage_1__2192_,
  data_stage_1__2191_,data_stage_1__2190_,data_stage_1__2189_,data_stage_1__2188_,
  data_stage_1__2187_,data_stage_1__2186_,data_stage_1__2185_,data_stage_1__2184_,
  data_stage_1__2183_,data_stage_1__2182_,data_stage_1__2181_,data_stage_1__2180_,
  data_stage_1__2179_,data_stage_1__2178_,data_stage_1__2177_,data_stage_1__2176_,
  data_stage_1__2175_,data_stage_1__2174_,data_stage_1__2173_,data_stage_1__2172_,
  data_stage_1__2171_,data_stage_1__2170_,data_stage_1__2169_,data_stage_1__2168_,
  data_stage_1__2167_,data_stage_1__2166_,data_stage_1__2165_,data_stage_1__2164_,
  data_stage_1__2163_,data_stage_1__2162_,data_stage_1__2161_,data_stage_1__2160_,
  data_stage_1__2159_,data_stage_1__2158_,data_stage_1__2157_,data_stage_1__2156_,
  data_stage_1__2155_,data_stage_1__2154_,data_stage_1__2153_,data_stage_1__2152_,
  data_stage_1__2151_,data_stage_1__2150_,data_stage_1__2149_,data_stage_1__2148_,
  data_stage_1__2147_,data_stage_1__2146_,data_stage_1__2145_,data_stage_1__2144_,
  data_stage_1__2143_,data_stage_1__2142_,data_stage_1__2141_,data_stage_1__2140_,
  data_stage_1__2139_,data_stage_1__2138_,data_stage_1__2137_,data_stage_1__2136_,
  data_stage_1__2135_,data_stage_1__2134_,data_stage_1__2133_,data_stage_1__2132_,
  data_stage_1__2131_,data_stage_1__2130_,data_stage_1__2129_,data_stage_1__2128_,
  data_stage_1__2127_,data_stage_1__2126_,data_stage_1__2125_,data_stage_1__2124_,
  data_stage_1__2123_,data_stage_1__2122_,data_stage_1__2121_,data_stage_1__2120_,
  data_stage_1__2119_,data_stage_1__2118_,data_stage_1__2117_,data_stage_1__2116_,
  data_stage_1__2115_,data_stage_1__2114_,data_stage_1__2113_,data_stage_1__2112_,
  data_stage_1__2111_,data_stage_1__2110_,data_stage_1__2109_,data_stage_1__2108_,
  data_stage_1__2107_,data_stage_1__2106_,data_stage_1__2105_,data_stage_1__2104_,
  data_stage_1__2103_,data_stage_1__2102_,data_stage_1__2101_,data_stage_1__2100_,
  data_stage_1__2099_,data_stage_1__2098_,data_stage_1__2097_,data_stage_1__2096_,
  data_stage_1__2095_,data_stage_1__2094_,data_stage_1__2093_,data_stage_1__2092_,
  data_stage_1__2091_,data_stage_1__2090_,data_stage_1__2089_,data_stage_1__2088_,
  data_stage_1__2087_,data_stage_1__2086_,data_stage_1__2085_,data_stage_1__2084_,
  data_stage_1__2083_,data_stage_1__2082_,data_stage_1__2081_,data_stage_1__2080_,
  data_stage_1__2079_,data_stage_1__2078_,data_stage_1__2077_,data_stage_1__2076_,
  data_stage_1__2075_,data_stage_1__2074_,data_stage_1__2073_,data_stage_1__2072_,
  data_stage_1__2071_,data_stage_1__2070_,data_stage_1__2069_,data_stage_1__2068_,
  data_stage_1__2067_,data_stage_1__2066_,data_stage_1__2065_,data_stage_1__2064_,
  data_stage_1__2063_,data_stage_1__2062_,data_stage_1__2061_,data_stage_1__2060_,
  data_stage_1__2059_,data_stage_1__2058_,data_stage_1__2057_,data_stage_1__2056_,
  data_stage_1__2055_,data_stage_1__2054_,data_stage_1__2053_,data_stage_1__2052_,
  data_stage_1__2051_,data_stage_1__2050_,data_stage_1__2049_,data_stage_1__2048_,
  data_stage_1__2047_,data_stage_1__2046_,data_stage_1__2045_,data_stage_1__2044_,
  data_stage_1__2043_,data_stage_1__2042_,data_stage_1__2041_,data_stage_1__2040_,
  data_stage_1__2039_,data_stage_1__2038_,data_stage_1__2037_,data_stage_1__2036_,
  data_stage_1__2035_,data_stage_1__2034_,data_stage_1__2033_,data_stage_1__2032_,
  data_stage_1__2031_,data_stage_1__2030_,data_stage_1__2029_,data_stage_1__2028_,
  data_stage_1__2027_,data_stage_1__2026_,data_stage_1__2025_,data_stage_1__2024_,
  data_stage_1__2023_,data_stage_1__2022_,data_stage_1__2021_,data_stage_1__2020_,
  data_stage_1__2019_,data_stage_1__2018_,data_stage_1__2017_,data_stage_1__2016_,
  data_stage_1__2015_,data_stage_1__2014_,data_stage_1__2013_,data_stage_1__2012_,
  data_stage_1__2011_,data_stage_1__2010_,data_stage_1__2009_,data_stage_1__2008_,
  data_stage_1__2007_,data_stage_1__2006_,data_stage_1__2005_,data_stage_1__2004_,
  data_stage_1__2003_,data_stage_1__2002_,data_stage_1__2001_,data_stage_1__2000_,
  data_stage_1__1999_,data_stage_1__1998_,data_stage_1__1997_,data_stage_1__1996_,
  data_stage_1__1995_,data_stage_1__1994_,data_stage_1__1993_,data_stage_1__1992_,
  data_stage_1__1991_,data_stage_1__1990_,data_stage_1__1989_,data_stage_1__1988_,
  data_stage_1__1987_,data_stage_1__1986_,data_stage_1__1985_,data_stage_1__1984_,
  data_stage_1__1983_,data_stage_1__1982_,data_stage_1__1981_,data_stage_1__1980_,
  data_stage_1__1979_,data_stage_1__1978_,data_stage_1__1977_,data_stage_1__1976_,
  data_stage_1__1975_,data_stage_1__1974_,data_stage_1__1973_,data_stage_1__1972_,
  data_stage_1__1971_,data_stage_1__1970_,data_stage_1__1969_,data_stage_1__1968_,
  data_stage_1__1967_,data_stage_1__1966_,data_stage_1__1965_,data_stage_1__1964_,
  data_stage_1__1963_,data_stage_1__1962_,data_stage_1__1961_,data_stage_1__1960_,
  data_stage_1__1959_,data_stage_1__1958_,data_stage_1__1957_,data_stage_1__1956_,
  data_stage_1__1955_,data_stage_1__1954_,data_stage_1__1953_,data_stage_1__1952_,
  data_stage_1__1951_,data_stage_1__1950_,data_stage_1__1949_,data_stage_1__1948_,
  data_stage_1__1947_,data_stage_1__1946_,data_stage_1__1945_,data_stage_1__1944_,
  data_stage_1__1943_,data_stage_1__1942_,data_stage_1__1941_,data_stage_1__1940_,
  data_stage_1__1939_,data_stage_1__1938_,data_stage_1__1937_,data_stage_1__1936_,
  data_stage_1__1935_,data_stage_1__1934_,data_stage_1__1933_,data_stage_1__1932_,
  data_stage_1__1931_,data_stage_1__1930_,data_stage_1__1929_,data_stage_1__1928_,
  data_stage_1__1927_,data_stage_1__1926_,data_stage_1__1925_,data_stage_1__1924_,
  data_stage_1__1923_,data_stage_1__1922_,data_stage_1__1921_,data_stage_1__1920_,
  data_stage_1__1919_,data_stage_1__1918_,data_stage_1__1917_,data_stage_1__1916_,
  data_stage_1__1915_,data_stage_1__1914_,data_stage_1__1913_,data_stage_1__1912_,
  data_stage_1__1911_,data_stage_1__1910_,data_stage_1__1909_,data_stage_1__1908_,
  data_stage_1__1907_,data_stage_1__1906_,data_stage_1__1905_,data_stage_1__1904_,
  data_stage_1__1903_,data_stage_1__1902_,data_stage_1__1901_,data_stage_1__1900_,
  data_stage_1__1899_,data_stage_1__1898_,data_stage_1__1897_,data_stage_1__1896_,
  data_stage_1__1895_,data_stage_1__1894_,data_stage_1__1893_,data_stage_1__1892_,
  data_stage_1__1891_,data_stage_1__1890_,data_stage_1__1889_,data_stage_1__1888_,
  data_stage_1__1887_,data_stage_1__1886_,data_stage_1__1885_,data_stage_1__1884_,
  data_stage_1__1883_,data_stage_1__1882_,data_stage_1__1881_,data_stage_1__1880_,
  data_stage_1__1879_,data_stage_1__1878_,data_stage_1__1877_,data_stage_1__1876_,
  data_stage_1__1875_,data_stage_1__1874_,data_stage_1__1873_,data_stage_1__1872_,
  data_stage_1__1871_,data_stage_1__1870_,data_stage_1__1869_,data_stage_1__1868_,
  data_stage_1__1867_,data_stage_1__1866_,data_stage_1__1865_,data_stage_1__1864_,
  data_stage_1__1863_,data_stage_1__1862_,data_stage_1__1861_,data_stage_1__1860_,
  data_stage_1__1859_,data_stage_1__1858_,data_stage_1__1857_,data_stage_1__1856_,
  data_stage_1__1855_,data_stage_1__1854_,data_stage_1__1853_,data_stage_1__1852_,
  data_stage_1__1851_,data_stage_1__1850_,data_stage_1__1849_,data_stage_1__1848_,
  data_stage_1__1847_,data_stage_1__1846_,data_stage_1__1845_,data_stage_1__1844_,
  data_stage_1__1843_,data_stage_1__1842_,data_stage_1__1841_,data_stage_1__1840_,
  data_stage_1__1839_,data_stage_1__1838_,data_stage_1__1837_,data_stage_1__1836_,
  data_stage_1__1835_,data_stage_1__1834_,data_stage_1__1833_,data_stage_1__1832_,
  data_stage_1__1831_,data_stage_1__1830_,data_stage_1__1829_,data_stage_1__1828_,
  data_stage_1__1827_,data_stage_1__1826_,data_stage_1__1825_,data_stage_1__1824_,
  data_stage_1__1823_,data_stage_1__1822_,data_stage_1__1821_,data_stage_1__1820_,
  data_stage_1__1819_,data_stage_1__1818_,data_stage_1__1817_,data_stage_1__1816_,
  data_stage_1__1815_,data_stage_1__1814_,data_stage_1__1813_,data_stage_1__1812_,
  data_stage_1__1811_,data_stage_1__1810_,data_stage_1__1809_,data_stage_1__1808_,
  data_stage_1__1807_,data_stage_1__1806_,data_stage_1__1805_,data_stage_1__1804_,
  data_stage_1__1803_,data_stage_1__1802_,data_stage_1__1801_,data_stage_1__1800_,
  data_stage_1__1799_,data_stage_1__1798_,data_stage_1__1797_,data_stage_1__1796_,
  data_stage_1__1795_,data_stage_1__1794_,data_stage_1__1793_,data_stage_1__1792_,
  data_stage_1__1791_,data_stage_1__1790_,data_stage_1__1789_,data_stage_1__1788_,
  data_stage_1__1787_,data_stage_1__1786_,data_stage_1__1785_,data_stage_1__1784_,
  data_stage_1__1783_,data_stage_1__1782_,data_stage_1__1781_,data_stage_1__1780_,
  data_stage_1__1779_,data_stage_1__1778_,data_stage_1__1777_,data_stage_1__1776_,
  data_stage_1__1775_,data_stage_1__1774_,data_stage_1__1773_,data_stage_1__1772_,
  data_stage_1__1771_,data_stage_1__1770_,data_stage_1__1769_,data_stage_1__1768_,
  data_stage_1__1767_,data_stage_1__1766_,data_stage_1__1765_,data_stage_1__1764_,
  data_stage_1__1763_,data_stage_1__1762_,data_stage_1__1761_,data_stage_1__1760_,
  data_stage_1__1759_,data_stage_1__1758_,data_stage_1__1757_,data_stage_1__1756_,
  data_stage_1__1755_,data_stage_1__1754_,data_stage_1__1753_,data_stage_1__1752_,
  data_stage_1__1751_,data_stage_1__1750_,data_stage_1__1749_,data_stage_1__1748_,
  data_stage_1__1747_,data_stage_1__1746_,data_stage_1__1745_,data_stage_1__1744_,
  data_stage_1__1743_,data_stage_1__1742_,data_stage_1__1741_,data_stage_1__1740_,
  data_stage_1__1739_,data_stage_1__1738_,data_stage_1__1737_,data_stage_1__1736_,
  data_stage_1__1735_,data_stage_1__1734_,data_stage_1__1733_,data_stage_1__1732_,
  data_stage_1__1731_,data_stage_1__1730_,data_stage_1__1729_,data_stage_1__1728_,
  data_stage_1__1727_,data_stage_1__1726_,data_stage_1__1725_,data_stage_1__1724_,
  data_stage_1__1723_,data_stage_1__1722_,data_stage_1__1721_,data_stage_1__1720_,
  data_stage_1__1719_,data_stage_1__1718_,data_stage_1__1717_,data_stage_1__1716_,
  data_stage_1__1715_,data_stage_1__1714_,data_stage_1__1713_,data_stage_1__1712_,
  data_stage_1__1711_,data_stage_1__1710_,data_stage_1__1709_,data_stage_1__1708_,
  data_stage_1__1707_,data_stage_1__1706_,data_stage_1__1705_,data_stage_1__1704_,
  data_stage_1__1703_,data_stage_1__1702_,data_stage_1__1701_,data_stage_1__1700_,
  data_stage_1__1699_,data_stage_1__1698_,data_stage_1__1697_,data_stage_1__1696_,
  data_stage_1__1695_,data_stage_1__1694_,data_stage_1__1693_,data_stage_1__1692_,
  data_stage_1__1691_,data_stage_1__1690_,data_stage_1__1689_,data_stage_1__1688_,
  data_stage_1__1687_,data_stage_1__1686_,data_stage_1__1685_,data_stage_1__1684_,
  data_stage_1__1683_,data_stage_1__1682_,data_stage_1__1681_,data_stage_1__1680_,
  data_stage_1__1679_,data_stage_1__1678_,data_stage_1__1677_,data_stage_1__1676_,
  data_stage_1__1675_,data_stage_1__1674_,data_stage_1__1673_,data_stage_1__1672_,
  data_stage_1__1671_,data_stage_1__1670_,data_stage_1__1669_,data_stage_1__1668_,
  data_stage_1__1667_,data_stage_1__1666_,data_stage_1__1665_,data_stage_1__1664_,
  data_stage_1__1663_,data_stage_1__1662_,data_stage_1__1661_,data_stage_1__1660_,
  data_stage_1__1659_,data_stage_1__1658_,data_stage_1__1657_,data_stage_1__1656_,
  data_stage_1__1655_,data_stage_1__1654_,data_stage_1__1653_,data_stage_1__1652_,
  data_stage_1__1651_,data_stage_1__1650_,data_stage_1__1649_,data_stage_1__1648_,
  data_stage_1__1647_,data_stage_1__1646_,data_stage_1__1645_,data_stage_1__1644_,
  data_stage_1__1643_,data_stage_1__1642_,data_stage_1__1641_,data_stage_1__1640_,
  data_stage_1__1639_,data_stage_1__1638_,data_stage_1__1637_,data_stage_1__1636_,
  data_stage_1__1635_,data_stage_1__1634_,data_stage_1__1633_,data_stage_1__1632_,
  data_stage_1__1631_,data_stage_1__1630_,data_stage_1__1629_,data_stage_1__1628_,
  data_stage_1__1627_,data_stage_1__1626_,data_stage_1__1625_,data_stage_1__1624_,
  data_stage_1__1623_,data_stage_1__1622_,data_stage_1__1621_,data_stage_1__1620_,
  data_stage_1__1619_,data_stage_1__1618_,data_stage_1__1617_,data_stage_1__1616_,
  data_stage_1__1615_,data_stage_1__1614_,data_stage_1__1613_,data_stage_1__1612_,
  data_stage_1__1611_,data_stage_1__1610_,data_stage_1__1609_,data_stage_1__1608_,
  data_stage_1__1607_,data_stage_1__1606_,data_stage_1__1605_,data_stage_1__1604_,
  data_stage_1__1603_,data_stage_1__1602_,data_stage_1__1601_,data_stage_1__1600_,
  data_stage_1__1599_,data_stage_1__1598_,data_stage_1__1597_,data_stage_1__1596_,
  data_stage_1__1595_,data_stage_1__1594_,data_stage_1__1593_,data_stage_1__1592_,
  data_stage_1__1591_,data_stage_1__1590_,data_stage_1__1589_,data_stage_1__1588_,
  data_stage_1__1587_,data_stage_1__1586_,data_stage_1__1585_,data_stage_1__1584_,
  data_stage_1__1583_,data_stage_1__1582_,data_stage_1__1581_,data_stage_1__1580_,
  data_stage_1__1579_,data_stage_1__1578_,data_stage_1__1577_,data_stage_1__1576_,
  data_stage_1__1575_,data_stage_1__1574_,data_stage_1__1573_,data_stage_1__1572_,
  data_stage_1__1571_,data_stage_1__1570_,data_stage_1__1569_,data_stage_1__1568_,
  data_stage_1__1567_,data_stage_1__1566_,data_stage_1__1565_,data_stage_1__1564_,
  data_stage_1__1563_,data_stage_1__1562_,data_stage_1__1561_,data_stage_1__1560_,
  data_stage_1__1559_,data_stage_1__1558_,data_stage_1__1557_,data_stage_1__1556_,
  data_stage_1__1555_,data_stage_1__1554_,data_stage_1__1553_,data_stage_1__1552_,
  data_stage_1__1551_,data_stage_1__1550_,data_stage_1__1549_,data_stage_1__1548_,
  data_stage_1__1547_,data_stage_1__1546_,data_stage_1__1545_,data_stage_1__1544_,
  data_stage_1__1543_,data_stage_1__1542_,data_stage_1__1541_,data_stage_1__1540_,
  data_stage_1__1539_,data_stage_1__1538_,data_stage_1__1537_,data_stage_1__1536_,
  data_stage_1__1535_,data_stage_1__1534_,data_stage_1__1533_,data_stage_1__1532_,
  data_stage_1__1531_,data_stage_1__1530_,data_stage_1__1529_,data_stage_1__1528_,
  data_stage_1__1527_,data_stage_1__1526_,data_stage_1__1525_,data_stage_1__1524_,
  data_stage_1__1523_,data_stage_1__1522_,data_stage_1__1521_,data_stage_1__1520_,
  data_stage_1__1519_,data_stage_1__1518_,data_stage_1__1517_,data_stage_1__1516_,
  data_stage_1__1515_,data_stage_1__1514_,data_stage_1__1513_,data_stage_1__1512_,
  data_stage_1__1511_,data_stage_1__1510_,data_stage_1__1509_,data_stage_1__1508_,
  data_stage_1__1507_,data_stage_1__1506_,data_stage_1__1505_,data_stage_1__1504_,
  data_stage_1__1503_,data_stage_1__1502_,data_stage_1__1501_,data_stage_1__1500_,
  data_stage_1__1499_,data_stage_1__1498_,data_stage_1__1497_,data_stage_1__1496_,
  data_stage_1__1495_,data_stage_1__1494_,data_stage_1__1493_,data_stage_1__1492_,
  data_stage_1__1491_,data_stage_1__1490_,data_stage_1__1489_,data_stage_1__1488_,
  data_stage_1__1487_,data_stage_1__1486_,data_stage_1__1485_,data_stage_1__1484_,
  data_stage_1__1483_,data_stage_1__1482_,data_stage_1__1481_,data_stage_1__1480_,
  data_stage_1__1479_,data_stage_1__1478_,data_stage_1__1477_,data_stage_1__1476_,
  data_stage_1__1475_,data_stage_1__1474_,data_stage_1__1473_,data_stage_1__1472_,
  data_stage_1__1471_,data_stage_1__1470_,data_stage_1__1469_,data_stage_1__1468_,
  data_stage_1__1467_,data_stage_1__1466_,data_stage_1__1465_,data_stage_1__1464_,
  data_stage_1__1463_,data_stage_1__1462_,data_stage_1__1461_,data_stage_1__1460_,
  data_stage_1__1459_,data_stage_1__1458_,data_stage_1__1457_,data_stage_1__1456_,
  data_stage_1__1455_,data_stage_1__1454_,data_stage_1__1453_,data_stage_1__1452_,
  data_stage_1__1451_,data_stage_1__1450_,data_stage_1__1449_,data_stage_1__1448_,
  data_stage_1__1447_,data_stage_1__1446_,data_stage_1__1445_,data_stage_1__1444_,
  data_stage_1__1443_,data_stage_1__1442_,data_stage_1__1441_,data_stage_1__1440_,
  data_stage_1__1439_,data_stage_1__1438_,data_stage_1__1437_,data_stage_1__1436_,
  data_stage_1__1435_,data_stage_1__1434_,data_stage_1__1433_,data_stage_1__1432_,
  data_stage_1__1431_,data_stage_1__1430_,data_stage_1__1429_,data_stage_1__1428_,
  data_stage_1__1427_,data_stage_1__1426_,data_stage_1__1425_,data_stage_1__1424_,
  data_stage_1__1423_,data_stage_1__1422_,data_stage_1__1421_,data_stage_1__1420_,
  data_stage_1__1419_,data_stage_1__1418_,data_stage_1__1417_,data_stage_1__1416_,
  data_stage_1__1415_,data_stage_1__1414_,data_stage_1__1413_,data_stage_1__1412_,
  data_stage_1__1411_,data_stage_1__1410_,data_stage_1__1409_,data_stage_1__1408_,
  data_stage_1__1407_,data_stage_1__1406_,data_stage_1__1405_,data_stage_1__1404_,
  data_stage_1__1403_,data_stage_1__1402_,data_stage_1__1401_,data_stage_1__1400_,
  data_stage_1__1399_,data_stage_1__1398_,data_stage_1__1397_,data_stage_1__1396_,
  data_stage_1__1395_,data_stage_1__1394_,data_stage_1__1393_,data_stage_1__1392_,
  data_stage_1__1391_,data_stage_1__1390_,data_stage_1__1389_,data_stage_1__1388_,
  data_stage_1__1387_,data_stage_1__1386_,data_stage_1__1385_,data_stage_1__1384_,
  data_stage_1__1383_,data_stage_1__1382_,data_stage_1__1381_,data_stage_1__1380_,
  data_stage_1__1379_,data_stage_1__1378_,data_stage_1__1377_,data_stage_1__1376_,
  data_stage_1__1375_,data_stage_1__1374_,data_stage_1__1373_,data_stage_1__1372_,
  data_stage_1__1371_,data_stage_1__1370_,data_stage_1__1369_,data_stage_1__1368_,
  data_stage_1__1367_,data_stage_1__1366_,data_stage_1__1365_,data_stage_1__1364_,
  data_stage_1__1363_,data_stage_1__1362_,data_stage_1__1361_,data_stage_1__1360_,
  data_stage_1__1359_,data_stage_1__1358_,data_stage_1__1357_,data_stage_1__1356_,
  data_stage_1__1355_,data_stage_1__1354_,data_stage_1__1353_,data_stage_1__1352_,
  data_stage_1__1351_,data_stage_1__1350_,data_stage_1__1349_,data_stage_1__1348_,
  data_stage_1__1347_,data_stage_1__1346_,data_stage_1__1345_,data_stage_1__1344_,
  data_stage_1__1343_,data_stage_1__1342_,data_stage_1__1341_,data_stage_1__1340_,
  data_stage_1__1339_,data_stage_1__1338_,data_stage_1__1337_,data_stage_1__1336_,
  data_stage_1__1335_,data_stage_1__1334_,data_stage_1__1333_,data_stage_1__1332_,
  data_stage_1__1331_,data_stage_1__1330_,data_stage_1__1329_,data_stage_1__1328_,
  data_stage_1__1327_,data_stage_1__1326_,data_stage_1__1325_,data_stage_1__1324_,
  data_stage_1__1323_,data_stage_1__1322_,data_stage_1__1321_,data_stage_1__1320_,
  data_stage_1__1319_,data_stage_1__1318_,data_stage_1__1317_,data_stage_1__1316_,
  data_stage_1__1315_,data_stage_1__1314_,data_stage_1__1313_,data_stage_1__1312_,
  data_stage_1__1311_,data_stage_1__1310_,data_stage_1__1309_,data_stage_1__1308_,
  data_stage_1__1307_,data_stage_1__1306_,data_stage_1__1305_,data_stage_1__1304_,
  data_stage_1__1303_,data_stage_1__1302_,data_stage_1__1301_,data_stage_1__1300_,
  data_stage_1__1299_,data_stage_1__1298_,data_stage_1__1297_,data_stage_1__1296_,
  data_stage_1__1295_,data_stage_1__1294_,data_stage_1__1293_,data_stage_1__1292_,
  data_stage_1__1291_,data_stage_1__1290_,data_stage_1__1289_,data_stage_1__1288_,
  data_stage_1__1287_,data_stage_1__1286_,data_stage_1__1285_,data_stage_1__1284_,
  data_stage_1__1283_,data_stage_1__1282_,data_stage_1__1281_,data_stage_1__1280_,
  data_stage_1__1279_,data_stage_1__1278_,data_stage_1__1277_,data_stage_1__1276_,
  data_stage_1__1275_,data_stage_1__1274_,data_stage_1__1273_,data_stage_1__1272_,
  data_stage_1__1271_,data_stage_1__1270_,data_stage_1__1269_,data_stage_1__1268_,
  data_stage_1__1267_,data_stage_1__1266_,data_stage_1__1265_,data_stage_1__1264_,
  data_stage_1__1263_,data_stage_1__1262_,data_stage_1__1261_,data_stage_1__1260_,
  data_stage_1__1259_,data_stage_1__1258_,data_stage_1__1257_,data_stage_1__1256_,
  data_stage_1__1255_,data_stage_1__1254_,data_stage_1__1253_,data_stage_1__1252_,
  data_stage_1__1251_,data_stage_1__1250_,data_stage_1__1249_,data_stage_1__1248_,
  data_stage_1__1247_,data_stage_1__1246_,data_stage_1__1245_,data_stage_1__1244_,
  data_stage_1__1243_,data_stage_1__1242_,data_stage_1__1241_,data_stage_1__1240_,
  data_stage_1__1239_,data_stage_1__1238_,data_stage_1__1237_,data_stage_1__1236_,
  data_stage_1__1235_,data_stage_1__1234_,data_stage_1__1233_,data_stage_1__1232_,
  data_stage_1__1231_,data_stage_1__1230_,data_stage_1__1229_,data_stage_1__1228_,
  data_stage_1__1227_,data_stage_1__1226_,data_stage_1__1225_,data_stage_1__1224_,
  data_stage_1__1223_,data_stage_1__1222_,data_stage_1__1221_,data_stage_1__1220_,
  data_stage_1__1219_,data_stage_1__1218_,data_stage_1__1217_,data_stage_1__1216_,
  data_stage_1__1215_,data_stage_1__1214_,data_stage_1__1213_,data_stage_1__1212_,
  data_stage_1__1211_,data_stage_1__1210_,data_stage_1__1209_,data_stage_1__1208_,
  data_stage_1__1207_,data_stage_1__1206_,data_stage_1__1205_,data_stage_1__1204_,
  data_stage_1__1203_,data_stage_1__1202_,data_stage_1__1201_,data_stage_1__1200_,
  data_stage_1__1199_,data_stage_1__1198_,data_stage_1__1197_,data_stage_1__1196_,
  data_stage_1__1195_,data_stage_1__1194_,data_stage_1__1193_,data_stage_1__1192_,
  data_stage_1__1191_,data_stage_1__1190_,data_stage_1__1189_,data_stage_1__1188_,
  data_stage_1__1187_,data_stage_1__1186_,data_stage_1__1185_,data_stage_1__1184_,
  data_stage_1__1183_,data_stage_1__1182_,data_stage_1__1181_,data_stage_1__1180_,
  data_stage_1__1179_,data_stage_1__1178_,data_stage_1__1177_,data_stage_1__1176_,
  data_stage_1__1175_,data_stage_1__1174_,data_stage_1__1173_,data_stage_1__1172_,
  data_stage_1__1171_,data_stage_1__1170_,data_stage_1__1169_,data_stage_1__1168_,
  data_stage_1__1167_,data_stage_1__1166_,data_stage_1__1165_,data_stage_1__1164_,
  data_stage_1__1163_,data_stage_1__1162_,data_stage_1__1161_,data_stage_1__1160_,
  data_stage_1__1159_,data_stage_1__1158_,data_stage_1__1157_,data_stage_1__1156_,
  data_stage_1__1155_,data_stage_1__1154_,data_stage_1__1153_,data_stage_1__1152_,
  data_stage_1__1151_,data_stage_1__1150_,data_stage_1__1149_,data_stage_1__1148_,
  data_stage_1__1147_,data_stage_1__1146_,data_stage_1__1145_,data_stage_1__1144_,
  data_stage_1__1143_,data_stage_1__1142_,data_stage_1__1141_,data_stage_1__1140_,
  data_stage_1__1139_,data_stage_1__1138_,data_stage_1__1137_,data_stage_1__1136_,
  data_stage_1__1135_,data_stage_1__1134_,data_stage_1__1133_,data_stage_1__1132_,
  data_stage_1__1131_,data_stage_1__1130_,data_stage_1__1129_,data_stage_1__1128_,
  data_stage_1__1127_,data_stage_1__1126_,data_stage_1__1125_,data_stage_1__1124_,
  data_stage_1__1123_,data_stage_1__1122_,data_stage_1__1121_,data_stage_1__1120_,
  data_stage_1__1119_,data_stage_1__1118_,data_stage_1__1117_,data_stage_1__1116_,
  data_stage_1__1115_,data_stage_1__1114_,data_stage_1__1113_,data_stage_1__1112_,
  data_stage_1__1111_,data_stage_1__1110_,data_stage_1__1109_,data_stage_1__1108_,
  data_stage_1__1107_,data_stage_1__1106_,data_stage_1__1105_,data_stage_1__1104_,
  data_stage_1__1103_,data_stage_1__1102_,data_stage_1__1101_,data_stage_1__1100_,
  data_stage_1__1099_,data_stage_1__1098_,data_stage_1__1097_,data_stage_1__1096_,
  data_stage_1__1095_,data_stage_1__1094_,data_stage_1__1093_,data_stage_1__1092_,
  data_stage_1__1091_,data_stage_1__1090_,data_stage_1__1089_,data_stage_1__1088_,
  data_stage_1__1087_,data_stage_1__1086_,data_stage_1__1085_,data_stage_1__1084_,
  data_stage_1__1083_,data_stage_1__1082_,data_stage_1__1081_,data_stage_1__1080_,
  data_stage_1__1079_,data_stage_1__1078_,data_stage_1__1077_,data_stage_1__1076_,
  data_stage_1__1075_,data_stage_1__1074_,data_stage_1__1073_,data_stage_1__1072_,
  data_stage_1__1071_,data_stage_1__1070_,data_stage_1__1069_,data_stage_1__1068_,
  data_stage_1__1067_,data_stage_1__1066_,data_stage_1__1065_,data_stage_1__1064_,
  data_stage_1__1063_,data_stage_1__1062_,data_stage_1__1061_,data_stage_1__1060_,
  data_stage_1__1059_,data_stage_1__1058_,data_stage_1__1057_,data_stage_1__1056_,
  data_stage_1__1055_,data_stage_1__1054_,data_stage_1__1053_,data_stage_1__1052_,
  data_stage_1__1051_,data_stage_1__1050_,data_stage_1__1049_,data_stage_1__1048_,
  data_stage_1__1047_,data_stage_1__1046_,data_stage_1__1045_,data_stage_1__1044_,
  data_stage_1__1043_,data_stage_1__1042_,data_stage_1__1041_,data_stage_1__1040_,
  data_stage_1__1039_,data_stage_1__1038_,data_stage_1__1037_,data_stage_1__1036_,
  data_stage_1__1035_,data_stage_1__1034_,data_stage_1__1033_,data_stage_1__1032_,
  data_stage_1__1031_,data_stage_1__1030_,data_stage_1__1029_,data_stage_1__1028_,
  data_stage_1__1027_,data_stage_1__1026_,data_stage_1__1025_,data_stage_1__1024_,
  data_stage_1__1023_,data_stage_1__1022_,data_stage_1__1021_,data_stage_1__1020_,
  data_stage_1__1019_,data_stage_1__1018_,data_stage_1__1017_,data_stage_1__1016_,
  data_stage_1__1015_,data_stage_1__1014_,data_stage_1__1013_,data_stage_1__1012_,
  data_stage_1__1011_,data_stage_1__1010_,data_stage_1__1009_,data_stage_1__1008_,
  data_stage_1__1007_,data_stage_1__1006_,data_stage_1__1005_,data_stage_1__1004_,
  data_stage_1__1003_,data_stage_1__1002_,data_stage_1__1001_,data_stage_1__1000_,
  data_stage_1__999_,data_stage_1__998_,data_stage_1__997_,data_stage_1__996_,
  data_stage_1__995_,data_stage_1__994_,data_stage_1__993_,data_stage_1__992_,
  data_stage_1__991_,data_stage_1__990_,data_stage_1__989_,data_stage_1__988_,
  data_stage_1__987_,data_stage_1__986_,data_stage_1__985_,data_stage_1__984_,
  data_stage_1__983_,data_stage_1__982_,data_stage_1__981_,data_stage_1__980_,data_stage_1__979_,
  data_stage_1__978_,data_stage_1__977_,data_stage_1__976_,data_stage_1__975_,
  data_stage_1__974_,data_stage_1__973_,data_stage_1__972_,data_stage_1__971_,
  data_stage_1__970_,data_stage_1__969_,data_stage_1__968_,data_stage_1__967_,
  data_stage_1__966_,data_stage_1__965_,data_stage_1__964_,data_stage_1__963_,
  data_stage_1__962_,data_stage_1__961_,data_stage_1__960_,data_stage_1__959_,data_stage_1__958_,
  data_stage_1__957_,data_stage_1__956_,data_stage_1__955_,data_stage_1__954_,
  data_stage_1__953_,data_stage_1__952_,data_stage_1__951_,data_stage_1__950_,
  data_stage_1__949_,data_stage_1__948_,data_stage_1__947_,data_stage_1__946_,
  data_stage_1__945_,data_stage_1__944_,data_stage_1__943_,data_stage_1__942_,
  data_stage_1__941_,data_stage_1__940_,data_stage_1__939_,data_stage_1__938_,data_stage_1__937_,
  data_stage_1__936_,data_stage_1__935_,data_stage_1__934_,data_stage_1__933_,
  data_stage_1__932_,data_stage_1__931_,data_stage_1__930_,data_stage_1__929_,
  data_stage_1__928_,data_stage_1__927_,data_stage_1__926_,data_stage_1__925_,
  data_stage_1__924_,data_stage_1__923_,data_stage_1__922_,data_stage_1__921_,data_stage_1__920_,
  data_stage_1__919_,data_stage_1__918_,data_stage_1__917_,data_stage_1__916_,
  data_stage_1__915_,data_stage_1__914_,data_stage_1__913_,data_stage_1__912_,
  data_stage_1__911_,data_stage_1__910_,data_stage_1__909_,data_stage_1__908_,
  data_stage_1__907_,data_stage_1__906_,data_stage_1__905_,data_stage_1__904_,
  data_stage_1__903_,data_stage_1__902_,data_stage_1__901_,data_stage_1__900_,data_stage_1__899_,
  data_stage_1__898_,data_stage_1__897_,data_stage_1__896_,data_stage_1__895_,
  data_stage_1__894_,data_stage_1__893_,data_stage_1__892_,data_stage_1__891_,
  data_stage_1__890_,data_stage_1__889_,data_stage_1__888_,data_stage_1__887_,
  data_stage_1__886_,data_stage_1__885_,data_stage_1__884_,data_stage_1__883_,
  data_stage_1__882_,data_stage_1__881_,data_stage_1__880_,data_stage_1__879_,data_stage_1__878_,
  data_stage_1__877_,data_stage_1__876_,data_stage_1__875_,data_stage_1__874_,
  data_stage_1__873_,data_stage_1__872_,data_stage_1__871_,data_stage_1__870_,
  data_stage_1__869_,data_stage_1__868_,data_stage_1__867_,data_stage_1__866_,
  data_stage_1__865_,data_stage_1__864_,data_stage_1__863_,data_stage_1__862_,
  data_stage_1__861_,data_stage_1__860_,data_stage_1__859_,data_stage_1__858_,data_stage_1__857_,
  data_stage_1__856_,data_stage_1__855_,data_stage_1__854_,data_stage_1__853_,
  data_stage_1__852_,data_stage_1__851_,data_stage_1__850_,data_stage_1__849_,
  data_stage_1__848_,data_stage_1__847_,data_stage_1__846_,data_stage_1__845_,
  data_stage_1__844_,data_stage_1__843_,data_stage_1__842_,data_stage_1__841_,data_stage_1__840_,
  data_stage_1__839_,data_stage_1__838_,data_stage_1__837_,data_stage_1__836_,
  data_stage_1__835_,data_stage_1__834_,data_stage_1__833_,data_stage_1__832_,
  data_stage_1__831_,data_stage_1__830_,data_stage_1__829_,data_stage_1__828_,
  data_stage_1__827_,data_stage_1__826_,data_stage_1__825_,data_stage_1__824_,
  data_stage_1__823_,data_stage_1__822_,data_stage_1__821_,data_stage_1__820_,data_stage_1__819_,
  data_stage_1__818_,data_stage_1__817_,data_stage_1__816_,data_stage_1__815_,
  data_stage_1__814_,data_stage_1__813_,data_stage_1__812_,data_stage_1__811_,
  data_stage_1__810_,data_stage_1__809_,data_stage_1__808_,data_stage_1__807_,
  data_stage_1__806_,data_stage_1__805_,data_stage_1__804_,data_stage_1__803_,
  data_stage_1__802_,data_stage_1__801_,data_stage_1__800_,data_stage_1__799_,data_stage_1__798_,
  data_stage_1__797_,data_stage_1__796_,data_stage_1__795_,data_stage_1__794_,
  data_stage_1__793_,data_stage_1__792_,data_stage_1__791_,data_stage_1__790_,
  data_stage_1__789_,data_stage_1__788_,data_stage_1__787_,data_stage_1__786_,
  data_stage_1__785_,data_stage_1__784_,data_stage_1__783_,data_stage_1__782_,
  data_stage_1__781_,data_stage_1__780_,data_stage_1__779_,data_stage_1__778_,data_stage_1__777_,
  data_stage_1__776_,data_stage_1__775_,data_stage_1__774_,data_stage_1__773_,
  data_stage_1__772_,data_stage_1__771_,data_stage_1__770_,data_stage_1__769_,
  data_stage_1__768_,data_stage_1__767_,data_stage_1__766_,data_stage_1__765_,
  data_stage_1__764_,data_stage_1__763_,data_stage_1__762_,data_stage_1__761_,data_stage_1__760_,
  data_stage_1__759_,data_stage_1__758_,data_stage_1__757_,data_stage_1__756_,
  data_stage_1__755_,data_stage_1__754_,data_stage_1__753_,data_stage_1__752_,
  data_stage_1__751_,data_stage_1__750_,data_stage_1__749_,data_stage_1__748_,
  data_stage_1__747_,data_stage_1__746_,data_stage_1__745_,data_stage_1__744_,
  data_stage_1__743_,data_stage_1__742_,data_stage_1__741_,data_stage_1__740_,data_stage_1__739_,
  data_stage_1__738_,data_stage_1__737_,data_stage_1__736_,data_stage_1__735_,
  data_stage_1__734_,data_stage_1__733_,data_stage_1__732_,data_stage_1__731_,
  data_stage_1__730_,data_stage_1__729_,data_stage_1__728_,data_stage_1__727_,
  data_stage_1__726_,data_stage_1__725_,data_stage_1__724_,data_stage_1__723_,
  data_stage_1__722_,data_stage_1__721_,data_stage_1__720_,data_stage_1__719_,data_stage_1__718_,
  data_stage_1__717_,data_stage_1__716_,data_stage_1__715_,data_stage_1__714_,
  data_stage_1__713_,data_stage_1__712_,data_stage_1__711_,data_stage_1__710_,
  data_stage_1__709_,data_stage_1__708_,data_stage_1__707_,data_stage_1__706_,
  data_stage_1__705_,data_stage_1__704_,data_stage_1__703_,data_stage_1__702_,
  data_stage_1__701_,data_stage_1__700_,data_stage_1__699_,data_stage_1__698_,data_stage_1__697_,
  data_stage_1__696_,data_stage_1__695_,data_stage_1__694_,data_stage_1__693_,
  data_stage_1__692_,data_stage_1__691_,data_stage_1__690_,data_stage_1__689_,
  data_stage_1__688_,data_stage_1__687_,data_stage_1__686_,data_stage_1__685_,
  data_stage_1__684_,data_stage_1__683_,data_stage_1__682_,data_stage_1__681_,data_stage_1__680_,
  data_stage_1__679_,data_stage_1__678_,data_stage_1__677_,data_stage_1__676_,
  data_stage_1__675_,data_stage_1__674_,data_stage_1__673_,data_stage_1__672_,
  data_stage_1__671_,data_stage_1__670_,data_stage_1__669_,data_stage_1__668_,
  data_stage_1__667_,data_stage_1__666_,data_stage_1__665_,data_stage_1__664_,
  data_stage_1__663_,data_stage_1__662_,data_stage_1__661_,data_stage_1__660_,data_stage_1__659_,
  data_stage_1__658_,data_stage_1__657_,data_stage_1__656_,data_stage_1__655_,
  data_stage_1__654_,data_stage_1__653_,data_stage_1__652_,data_stage_1__651_,
  data_stage_1__650_,data_stage_1__649_,data_stage_1__648_,data_stage_1__647_,
  data_stage_1__646_,data_stage_1__645_,data_stage_1__644_,data_stage_1__643_,
  data_stage_1__642_,data_stage_1__641_,data_stage_1__640_,data_stage_1__639_,data_stage_1__638_,
  data_stage_1__637_,data_stage_1__636_,data_stage_1__635_,data_stage_1__634_,
  data_stage_1__633_,data_stage_1__632_,data_stage_1__631_,data_stage_1__630_,
  data_stage_1__629_,data_stage_1__628_,data_stage_1__627_,data_stage_1__626_,
  data_stage_1__625_,data_stage_1__624_,data_stage_1__623_,data_stage_1__622_,
  data_stage_1__621_,data_stage_1__620_,data_stage_1__619_,data_stage_1__618_,data_stage_1__617_,
  data_stage_1__616_,data_stage_1__615_,data_stage_1__614_,data_stage_1__613_,
  data_stage_1__612_,data_stage_1__611_,data_stage_1__610_,data_stage_1__609_,
  data_stage_1__608_,data_stage_1__607_,data_stage_1__606_,data_stage_1__605_,
  data_stage_1__604_,data_stage_1__603_,data_stage_1__602_,data_stage_1__601_,data_stage_1__600_,
  data_stage_1__599_,data_stage_1__598_,data_stage_1__597_,data_stage_1__596_,
  data_stage_1__595_,data_stage_1__594_,data_stage_1__593_,data_stage_1__592_,
  data_stage_1__591_,data_stage_1__590_,data_stage_1__589_,data_stage_1__588_,
  data_stage_1__587_,data_stage_1__586_,data_stage_1__585_,data_stage_1__584_,
  data_stage_1__583_,data_stage_1__582_,data_stage_1__581_,data_stage_1__580_,data_stage_1__579_,
  data_stage_1__578_,data_stage_1__577_,data_stage_1__576_,data_stage_1__575_,
  data_stage_1__574_,data_stage_1__573_,data_stage_1__572_,data_stage_1__571_,
  data_stage_1__570_,data_stage_1__569_,data_stage_1__568_,data_stage_1__567_,
  data_stage_1__566_,data_stage_1__565_,data_stage_1__564_,data_stage_1__563_,
  data_stage_1__562_,data_stage_1__561_,data_stage_1__560_,data_stage_1__559_,data_stage_1__558_,
  data_stage_1__557_,data_stage_1__556_,data_stage_1__555_,data_stage_1__554_,
  data_stage_1__553_,data_stage_1__552_,data_stage_1__551_,data_stage_1__550_,
  data_stage_1__549_,data_stage_1__548_,data_stage_1__547_,data_stage_1__546_,
  data_stage_1__545_,data_stage_1__544_,data_stage_1__543_,data_stage_1__542_,
  data_stage_1__541_,data_stage_1__540_,data_stage_1__539_,data_stage_1__538_,data_stage_1__537_,
  data_stage_1__536_,data_stage_1__535_,data_stage_1__534_,data_stage_1__533_,
  data_stage_1__532_,data_stage_1__531_,data_stage_1__530_,data_stage_1__529_,
  data_stage_1__528_,data_stage_1__527_,data_stage_1__526_,data_stage_1__525_,
  data_stage_1__524_,data_stage_1__523_,data_stage_1__522_,data_stage_1__521_,data_stage_1__520_,
  data_stage_1__519_,data_stage_1__518_,data_stage_1__517_,data_stage_1__516_,
  data_stage_1__515_,data_stage_1__514_,data_stage_1__513_,data_stage_1__512_,
  data_stage_1__511_,data_stage_1__510_,data_stage_1__509_,data_stage_1__508_,
  data_stage_1__507_,data_stage_1__506_,data_stage_1__505_,data_stage_1__504_,
  data_stage_1__503_,data_stage_1__502_,data_stage_1__501_,data_stage_1__500_,data_stage_1__499_,
  data_stage_1__498_,data_stage_1__497_,data_stage_1__496_,data_stage_1__495_,
  data_stage_1__494_,data_stage_1__493_,data_stage_1__492_,data_stage_1__491_,
  data_stage_1__490_,data_stage_1__489_,data_stage_1__488_,data_stage_1__487_,
  data_stage_1__486_,data_stage_1__485_,data_stage_1__484_,data_stage_1__483_,
  data_stage_1__482_,data_stage_1__481_,data_stage_1__480_,data_stage_1__479_,data_stage_1__478_,
  data_stage_1__477_,data_stage_1__476_,data_stage_1__475_,data_stage_1__474_,
  data_stage_1__473_,data_stage_1__472_,data_stage_1__471_,data_stage_1__470_,
  data_stage_1__469_,data_stage_1__468_,data_stage_1__467_,data_stage_1__466_,
  data_stage_1__465_,data_stage_1__464_,data_stage_1__463_,data_stage_1__462_,
  data_stage_1__461_,data_stage_1__460_,data_stage_1__459_,data_stage_1__458_,data_stage_1__457_,
  data_stage_1__456_,data_stage_1__455_,data_stage_1__454_,data_stage_1__453_,
  data_stage_1__452_,data_stage_1__451_,data_stage_1__450_,data_stage_1__449_,
  data_stage_1__448_,data_stage_1__447_,data_stage_1__446_,data_stage_1__445_,
  data_stage_1__444_,data_stage_1__443_,data_stage_1__442_,data_stage_1__441_,data_stage_1__440_,
  data_stage_1__439_,data_stage_1__438_,data_stage_1__437_,data_stage_1__436_,
  data_stage_1__435_,data_stage_1__434_,data_stage_1__433_,data_stage_1__432_,
  data_stage_1__431_,data_stage_1__430_,data_stage_1__429_,data_stage_1__428_,
  data_stage_1__427_,data_stage_1__426_,data_stage_1__425_,data_stage_1__424_,
  data_stage_1__423_,data_stage_1__422_,data_stage_1__421_,data_stage_1__420_,data_stage_1__419_,
  data_stage_1__418_,data_stage_1__417_,data_stage_1__416_,data_stage_1__415_,
  data_stage_1__414_,data_stage_1__413_,data_stage_1__412_,data_stage_1__411_,
  data_stage_1__410_,data_stage_1__409_,data_stage_1__408_,data_stage_1__407_,
  data_stage_1__406_,data_stage_1__405_,data_stage_1__404_,data_stage_1__403_,
  data_stage_1__402_,data_stage_1__401_,data_stage_1__400_,data_stage_1__399_,data_stage_1__398_,
  data_stage_1__397_,data_stage_1__396_,data_stage_1__395_,data_stage_1__394_,
  data_stage_1__393_,data_stage_1__392_,data_stage_1__391_,data_stage_1__390_,
  data_stage_1__389_,data_stage_1__388_,data_stage_1__387_,data_stage_1__386_,
  data_stage_1__385_,data_stage_1__384_,data_stage_1__383_,data_stage_1__382_,
  data_stage_1__381_,data_stage_1__380_,data_stage_1__379_,data_stage_1__378_,data_stage_1__377_,
  data_stage_1__376_,data_stage_1__375_,data_stage_1__374_,data_stage_1__373_,
  data_stage_1__372_,data_stage_1__371_,data_stage_1__370_,data_stage_1__369_,
  data_stage_1__368_,data_stage_1__367_,data_stage_1__366_,data_stage_1__365_,
  data_stage_1__364_,data_stage_1__363_,data_stage_1__362_,data_stage_1__361_,data_stage_1__360_,
  data_stage_1__359_,data_stage_1__358_,data_stage_1__357_,data_stage_1__356_,
  data_stage_1__355_,data_stage_1__354_,data_stage_1__353_,data_stage_1__352_,
  data_stage_1__351_,data_stage_1__350_,data_stage_1__349_,data_stage_1__348_,
  data_stage_1__347_,data_stage_1__346_,data_stage_1__345_,data_stage_1__344_,
  data_stage_1__343_,data_stage_1__342_,data_stage_1__341_,data_stage_1__340_,data_stage_1__339_,
  data_stage_1__338_,data_stage_1__337_,data_stage_1__336_,data_stage_1__335_,
  data_stage_1__334_,data_stage_1__333_,data_stage_1__332_,data_stage_1__331_,
  data_stage_1__330_,data_stage_1__329_,data_stage_1__328_,data_stage_1__327_,
  data_stage_1__326_,data_stage_1__325_,data_stage_1__324_,data_stage_1__323_,
  data_stage_1__322_,data_stage_1__321_,data_stage_1__320_,data_stage_1__319_,data_stage_1__318_,
  data_stage_1__317_,data_stage_1__316_,data_stage_1__315_,data_stage_1__314_,
  data_stage_1__313_,data_stage_1__312_,data_stage_1__311_,data_stage_1__310_,
  data_stage_1__309_,data_stage_1__308_,data_stage_1__307_,data_stage_1__306_,
  data_stage_1__305_,data_stage_1__304_,data_stage_1__303_,data_stage_1__302_,
  data_stage_1__301_,data_stage_1__300_,data_stage_1__299_,data_stage_1__298_,data_stage_1__297_,
  data_stage_1__296_,data_stage_1__295_,data_stage_1__294_,data_stage_1__293_,
  data_stage_1__292_,data_stage_1__291_,data_stage_1__290_,data_stage_1__289_,
  data_stage_1__288_,data_stage_1__287_,data_stage_1__286_,data_stage_1__285_,
  data_stage_1__284_,data_stage_1__283_,data_stage_1__282_,data_stage_1__281_,data_stage_1__280_,
  data_stage_1__279_,data_stage_1__278_,data_stage_1__277_,data_stage_1__276_,
  data_stage_1__275_,data_stage_1__274_,data_stage_1__273_,data_stage_1__272_,
  data_stage_1__271_,data_stage_1__270_,data_stage_1__269_,data_stage_1__268_,
  data_stage_1__267_,data_stage_1__266_,data_stage_1__265_,data_stage_1__264_,
  data_stage_1__263_,data_stage_1__262_,data_stage_1__261_,data_stage_1__260_,data_stage_1__259_,
  data_stage_1__258_,data_stage_1__257_,data_stage_1__256_,data_stage_1__255_,
  data_stage_1__254_,data_stage_1__253_,data_stage_1__252_,data_stage_1__251_,
  data_stage_1__250_,data_stage_1__249_,data_stage_1__248_,data_stage_1__247_,
  data_stage_1__246_,data_stage_1__245_,data_stage_1__244_,data_stage_1__243_,
  data_stage_1__242_,data_stage_1__241_,data_stage_1__240_,data_stage_1__239_,data_stage_1__238_,
  data_stage_1__237_,data_stage_1__236_,data_stage_1__235_,data_stage_1__234_,
  data_stage_1__233_,data_stage_1__232_,data_stage_1__231_,data_stage_1__230_,
  data_stage_1__229_,data_stage_1__228_,data_stage_1__227_,data_stage_1__226_,
  data_stage_1__225_,data_stage_1__224_,data_stage_1__223_,data_stage_1__222_,
  data_stage_1__221_,data_stage_1__220_,data_stage_1__219_,data_stage_1__218_,data_stage_1__217_,
  data_stage_1__216_,data_stage_1__215_,data_stage_1__214_,data_stage_1__213_,
  data_stage_1__212_,data_stage_1__211_,data_stage_1__210_,data_stage_1__209_,
  data_stage_1__208_,data_stage_1__207_,data_stage_1__206_,data_stage_1__205_,
  data_stage_1__204_,data_stage_1__203_,data_stage_1__202_,data_stage_1__201_,data_stage_1__200_,
  data_stage_1__199_,data_stage_1__198_,data_stage_1__197_,data_stage_1__196_,
  data_stage_1__195_,data_stage_1__194_,data_stage_1__193_,data_stage_1__192_,
  data_stage_1__191_,data_stage_1__190_,data_stage_1__189_,data_stage_1__188_,
  data_stage_1__187_,data_stage_1__186_,data_stage_1__185_,data_stage_1__184_,
  data_stage_1__183_,data_stage_1__182_,data_stage_1__181_,data_stage_1__180_,data_stage_1__179_,
  data_stage_1__178_,data_stage_1__177_,data_stage_1__176_,data_stage_1__175_,
  data_stage_1__174_,data_stage_1__173_,data_stage_1__172_,data_stage_1__171_,
  data_stage_1__170_,data_stage_1__169_,data_stage_1__168_,data_stage_1__167_,
  data_stage_1__166_,data_stage_1__165_,data_stage_1__164_,data_stage_1__163_,
  data_stage_1__162_,data_stage_1__161_,data_stage_1__160_,data_stage_1__159_,data_stage_1__158_,
  data_stage_1__157_,data_stage_1__156_,data_stage_1__155_,data_stage_1__154_,
  data_stage_1__153_,data_stage_1__152_,data_stage_1__151_,data_stage_1__150_,
  data_stage_1__149_,data_stage_1__148_,data_stage_1__147_,data_stage_1__146_,
  data_stage_1__145_,data_stage_1__144_,data_stage_1__143_,data_stage_1__142_,
  data_stage_1__141_,data_stage_1__140_,data_stage_1__139_,data_stage_1__138_,data_stage_1__137_,
  data_stage_1__136_,data_stage_1__135_,data_stage_1__134_,data_stage_1__133_,
  data_stage_1__132_,data_stage_1__131_,data_stage_1__130_,data_stage_1__129_,
  data_stage_1__128_,data_stage_1__127_,data_stage_1__126_,data_stage_1__125_,
  data_stage_1__124_,data_stage_1__123_,data_stage_1__122_,data_stage_1__121_,data_stage_1__120_,
  data_stage_1__119_,data_stage_1__118_,data_stage_1__117_,data_stage_1__116_,
  data_stage_1__115_,data_stage_1__114_,data_stage_1__113_,data_stage_1__112_,
  data_stage_1__111_,data_stage_1__110_,data_stage_1__109_,data_stage_1__108_,
  data_stage_1__107_,data_stage_1__106_,data_stage_1__105_,data_stage_1__104_,
  data_stage_1__103_,data_stage_1__102_,data_stage_1__101_,data_stage_1__100_,data_stage_1__99_,
  data_stage_1__98_,data_stage_1__97_,data_stage_1__96_,data_stage_1__95_,
  data_stage_1__94_,data_stage_1__93_,data_stage_1__92_,data_stage_1__91_,data_stage_1__90_,
  data_stage_1__89_,data_stage_1__88_,data_stage_1__87_,data_stage_1__86_,
  data_stage_1__85_,data_stage_1__84_,data_stage_1__83_,data_stage_1__82_,
  data_stage_1__81_,data_stage_1__80_,data_stage_1__79_,data_stage_1__78_,data_stage_1__77_,
  data_stage_1__76_,data_stage_1__75_,data_stage_1__74_,data_stage_1__73_,
  data_stage_1__72_,data_stage_1__71_,data_stage_1__70_,data_stage_1__69_,data_stage_1__68_,
  data_stage_1__67_,data_stage_1__66_,data_stage_1__65_,data_stage_1__64_,
  data_stage_1__63_,data_stage_1__62_,data_stage_1__61_,data_stage_1__60_,data_stage_1__59_,
  data_stage_1__58_,data_stage_1__57_,data_stage_1__56_,data_stage_1__55_,
  data_stage_1__54_,data_stage_1__53_,data_stage_1__52_,data_stage_1__51_,data_stage_1__50_,
  data_stage_1__49_,data_stage_1__48_,data_stage_1__47_,data_stage_1__46_,
  data_stage_1__45_,data_stage_1__44_,data_stage_1__43_,data_stage_1__42_,
  data_stage_1__41_,data_stage_1__40_,data_stage_1__39_,data_stage_1__38_,data_stage_1__37_,
  data_stage_1__36_,data_stage_1__35_,data_stage_1__34_,data_stage_1__33_,
  data_stage_1__32_,data_stage_1__31_,data_stage_1__30_,data_stage_1__29_,data_stage_1__28_,
  data_stage_1__27_,data_stage_1__26_,data_stage_1__25_,data_stage_1__24_,
  data_stage_1__23_,data_stage_1__22_,data_stage_1__21_,data_stage_1__20_,data_stage_1__19_,
  data_stage_1__18_,data_stage_1__17_,data_stage_1__16_,data_stage_1__15_,
  data_stage_1__14_,data_stage_1__13_,data_stage_1__12_,data_stage_1__11_,data_stage_1__10_,
  data_stage_1__9_,data_stage_1__8_,data_stage_1__7_,data_stage_1__6_,
  data_stage_1__5_,data_stage_1__4_,data_stage_1__3_,data_stage_1__2_,data_stage_1__1_,
  data_stage_1__0_,data_stage_2__8191_,data_stage_2__8190_,data_stage_2__8189_,
  data_stage_2__8188_,data_stage_2__8187_,data_stage_2__8186_,data_stage_2__8185_,
  data_stage_2__8184_,data_stage_2__8183_,data_stage_2__8182_,data_stage_2__8181_,
  data_stage_2__8180_,data_stage_2__8179_,data_stage_2__8178_,data_stage_2__8177_,
  data_stage_2__8176_,data_stage_2__8175_,data_stage_2__8174_,data_stage_2__8173_,
  data_stage_2__8172_,data_stage_2__8171_,data_stage_2__8170_,data_stage_2__8169_,
  data_stage_2__8168_,data_stage_2__8167_,data_stage_2__8166_,data_stage_2__8165_,
  data_stage_2__8164_,data_stage_2__8163_,data_stage_2__8162_,data_stage_2__8161_,
  data_stage_2__8160_,data_stage_2__8159_,data_stage_2__8158_,data_stage_2__8157_,
  data_stage_2__8156_,data_stage_2__8155_,data_stage_2__8154_,data_stage_2__8153_,
  data_stage_2__8152_,data_stage_2__8151_,data_stage_2__8150_,data_stage_2__8149_,
  data_stage_2__8148_,data_stage_2__8147_,data_stage_2__8146_,data_stage_2__8145_,
  data_stage_2__8144_,data_stage_2__8143_,data_stage_2__8142_,data_stage_2__8141_,
  data_stage_2__8140_,data_stage_2__8139_,data_stage_2__8138_,data_stage_2__8137_,
  data_stage_2__8136_,data_stage_2__8135_,data_stage_2__8134_,data_stage_2__8133_,
  data_stage_2__8132_,data_stage_2__8131_,data_stage_2__8130_,data_stage_2__8129_,
  data_stage_2__8128_,data_stage_2__8127_,data_stage_2__8126_,data_stage_2__8125_,
  data_stage_2__8124_,data_stage_2__8123_,data_stage_2__8122_,data_stage_2__8121_,
  data_stage_2__8120_,data_stage_2__8119_,data_stage_2__8118_,data_stage_2__8117_,
  data_stage_2__8116_,data_stage_2__8115_,data_stage_2__8114_,data_stage_2__8113_,
  data_stage_2__8112_,data_stage_2__8111_,data_stage_2__8110_,data_stage_2__8109_,
  data_stage_2__8108_,data_stage_2__8107_,data_stage_2__8106_,data_stage_2__8105_,
  data_stage_2__8104_,data_stage_2__8103_,data_stage_2__8102_,data_stage_2__8101_,
  data_stage_2__8100_,data_stage_2__8099_,data_stage_2__8098_,data_stage_2__8097_,
  data_stage_2__8096_,data_stage_2__8095_,data_stage_2__8094_,data_stage_2__8093_,
  data_stage_2__8092_,data_stage_2__8091_,data_stage_2__8090_,data_stage_2__8089_,
  data_stage_2__8088_,data_stage_2__8087_,data_stage_2__8086_,data_stage_2__8085_,
  data_stage_2__8084_,data_stage_2__8083_,data_stage_2__8082_,data_stage_2__8081_,
  data_stage_2__8080_,data_stage_2__8079_,data_stage_2__8078_,data_stage_2__8077_,
  data_stage_2__8076_,data_stage_2__8075_,data_stage_2__8074_,data_stage_2__8073_,
  data_stage_2__8072_,data_stage_2__8071_,data_stage_2__8070_,data_stage_2__8069_,
  data_stage_2__8068_,data_stage_2__8067_,data_stage_2__8066_,data_stage_2__8065_,
  data_stage_2__8064_,data_stage_2__8063_,data_stage_2__8062_,data_stage_2__8061_,
  data_stage_2__8060_,data_stage_2__8059_,data_stage_2__8058_,data_stage_2__8057_,
  data_stage_2__8056_,data_stage_2__8055_,data_stage_2__8054_,data_stage_2__8053_,
  data_stage_2__8052_,data_stage_2__8051_,data_stage_2__8050_,data_stage_2__8049_,
  data_stage_2__8048_,data_stage_2__8047_,data_stage_2__8046_,data_stage_2__8045_,
  data_stage_2__8044_,data_stage_2__8043_,data_stage_2__8042_,data_stage_2__8041_,
  data_stage_2__8040_,data_stage_2__8039_,data_stage_2__8038_,data_stage_2__8037_,
  data_stage_2__8036_,data_stage_2__8035_,data_stage_2__8034_,data_stage_2__8033_,
  data_stage_2__8032_,data_stage_2__8031_,data_stage_2__8030_,data_stage_2__8029_,
  data_stage_2__8028_,data_stage_2__8027_,data_stage_2__8026_,data_stage_2__8025_,
  data_stage_2__8024_,data_stage_2__8023_,data_stage_2__8022_,data_stage_2__8021_,
  data_stage_2__8020_,data_stage_2__8019_,data_stage_2__8018_,data_stage_2__8017_,
  data_stage_2__8016_,data_stage_2__8015_,data_stage_2__8014_,data_stage_2__8013_,
  data_stage_2__8012_,data_stage_2__8011_,data_stage_2__8010_,data_stage_2__8009_,
  data_stage_2__8008_,data_stage_2__8007_,data_stage_2__8006_,data_stage_2__8005_,
  data_stage_2__8004_,data_stage_2__8003_,data_stage_2__8002_,data_stage_2__8001_,
  data_stage_2__8000_,data_stage_2__7999_,data_stage_2__7998_,data_stage_2__7997_,
  data_stage_2__7996_,data_stage_2__7995_,data_stage_2__7994_,data_stage_2__7993_,
  data_stage_2__7992_,data_stage_2__7991_,data_stage_2__7990_,data_stage_2__7989_,
  data_stage_2__7988_,data_stage_2__7987_,data_stage_2__7986_,data_stage_2__7985_,
  data_stage_2__7984_,data_stage_2__7983_,data_stage_2__7982_,data_stage_2__7981_,
  data_stage_2__7980_,data_stage_2__7979_,data_stage_2__7978_,data_stage_2__7977_,
  data_stage_2__7976_,data_stage_2__7975_,data_stage_2__7974_,data_stage_2__7973_,
  data_stage_2__7972_,data_stage_2__7971_,data_stage_2__7970_,data_stage_2__7969_,
  data_stage_2__7968_,data_stage_2__7967_,data_stage_2__7966_,data_stage_2__7965_,
  data_stage_2__7964_,data_stage_2__7963_,data_stage_2__7962_,data_stage_2__7961_,
  data_stage_2__7960_,data_stage_2__7959_,data_stage_2__7958_,data_stage_2__7957_,
  data_stage_2__7956_,data_stage_2__7955_,data_stage_2__7954_,data_stage_2__7953_,
  data_stage_2__7952_,data_stage_2__7951_,data_stage_2__7950_,data_stage_2__7949_,
  data_stage_2__7948_,data_stage_2__7947_,data_stage_2__7946_,data_stage_2__7945_,
  data_stage_2__7944_,data_stage_2__7943_,data_stage_2__7942_,data_stage_2__7941_,
  data_stage_2__7940_,data_stage_2__7939_,data_stage_2__7938_,data_stage_2__7937_,
  data_stage_2__7936_,data_stage_2__7935_,data_stage_2__7934_,data_stage_2__7933_,
  data_stage_2__7932_,data_stage_2__7931_,data_stage_2__7930_,data_stage_2__7929_,
  data_stage_2__7928_,data_stage_2__7927_,data_stage_2__7926_,data_stage_2__7925_,
  data_stage_2__7924_,data_stage_2__7923_,data_stage_2__7922_,data_stage_2__7921_,
  data_stage_2__7920_,data_stage_2__7919_,data_stage_2__7918_,data_stage_2__7917_,
  data_stage_2__7916_,data_stage_2__7915_,data_stage_2__7914_,data_stage_2__7913_,
  data_stage_2__7912_,data_stage_2__7911_,data_stage_2__7910_,data_stage_2__7909_,
  data_stage_2__7908_,data_stage_2__7907_,data_stage_2__7906_,data_stage_2__7905_,
  data_stage_2__7904_,data_stage_2__7903_,data_stage_2__7902_,data_stage_2__7901_,
  data_stage_2__7900_,data_stage_2__7899_,data_stage_2__7898_,data_stage_2__7897_,
  data_stage_2__7896_,data_stage_2__7895_,data_stage_2__7894_,data_stage_2__7893_,
  data_stage_2__7892_,data_stage_2__7891_,data_stage_2__7890_,data_stage_2__7889_,
  data_stage_2__7888_,data_stage_2__7887_,data_stage_2__7886_,data_stage_2__7885_,
  data_stage_2__7884_,data_stage_2__7883_,data_stage_2__7882_,data_stage_2__7881_,
  data_stage_2__7880_,data_stage_2__7879_,data_stage_2__7878_,data_stage_2__7877_,
  data_stage_2__7876_,data_stage_2__7875_,data_stage_2__7874_,data_stage_2__7873_,
  data_stage_2__7872_,data_stage_2__7871_,data_stage_2__7870_,data_stage_2__7869_,
  data_stage_2__7868_,data_stage_2__7867_,data_stage_2__7866_,data_stage_2__7865_,
  data_stage_2__7864_,data_stage_2__7863_,data_stage_2__7862_,data_stage_2__7861_,
  data_stage_2__7860_,data_stage_2__7859_,data_stage_2__7858_,data_stage_2__7857_,
  data_stage_2__7856_,data_stage_2__7855_,data_stage_2__7854_,data_stage_2__7853_,
  data_stage_2__7852_,data_stage_2__7851_,data_stage_2__7850_,data_stage_2__7849_,
  data_stage_2__7848_,data_stage_2__7847_,data_stage_2__7846_,data_stage_2__7845_,
  data_stage_2__7844_,data_stage_2__7843_,data_stage_2__7842_,data_stage_2__7841_,
  data_stage_2__7840_,data_stage_2__7839_,data_stage_2__7838_,data_stage_2__7837_,
  data_stage_2__7836_,data_stage_2__7835_,data_stage_2__7834_,data_stage_2__7833_,
  data_stage_2__7832_,data_stage_2__7831_,data_stage_2__7830_,data_stage_2__7829_,
  data_stage_2__7828_,data_stage_2__7827_,data_stage_2__7826_,data_stage_2__7825_,
  data_stage_2__7824_,data_stage_2__7823_,data_stage_2__7822_,data_stage_2__7821_,
  data_stage_2__7820_,data_stage_2__7819_,data_stage_2__7818_,data_stage_2__7817_,
  data_stage_2__7816_,data_stage_2__7815_,data_stage_2__7814_,data_stage_2__7813_,
  data_stage_2__7812_,data_stage_2__7811_,data_stage_2__7810_,data_stage_2__7809_,
  data_stage_2__7808_,data_stage_2__7807_,data_stage_2__7806_,data_stage_2__7805_,
  data_stage_2__7804_,data_stage_2__7803_,data_stage_2__7802_,data_stage_2__7801_,
  data_stage_2__7800_,data_stage_2__7799_,data_stage_2__7798_,data_stage_2__7797_,
  data_stage_2__7796_,data_stage_2__7795_,data_stage_2__7794_,data_stage_2__7793_,
  data_stage_2__7792_,data_stage_2__7791_,data_stage_2__7790_,data_stage_2__7789_,
  data_stage_2__7788_,data_stage_2__7787_,data_stage_2__7786_,data_stage_2__7785_,
  data_stage_2__7784_,data_stage_2__7783_,data_stage_2__7782_,data_stage_2__7781_,
  data_stage_2__7780_,data_stage_2__7779_,data_stage_2__7778_,data_stage_2__7777_,
  data_stage_2__7776_,data_stage_2__7775_,data_stage_2__7774_,data_stage_2__7773_,
  data_stage_2__7772_,data_stage_2__7771_,data_stage_2__7770_,data_stage_2__7769_,
  data_stage_2__7768_,data_stage_2__7767_,data_stage_2__7766_,data_stage_2__7765_,
  data_stage_2__7764_,data_stage_2__7763_,data_stage_2__7762_,data_stage_2__7761_,
  data_stage_2__7760_,data_stage_2__7759_,data_stage_2__7758_,data_stage_2__7757_,
  data_stage_2__7756_,data_stage_2__7755_,data_stage_2__7754_,data_stage_2__7753_,
  data_stage_2__7752_,data_stage_2__7751_,data_stage_2__7750_,data_stage_2__7749_,
  data_stage_2__7748_,data_stage_2__7747_,data_stage_2__7746_,data_stage_2__7745_,
  data_stage_2__7744_,data_stage_2__7743_,data_stage_2__7742_,data_stage_2__7741_,
  data_stage_2__7740_,data_stage_2__7739_,data_stage_2__7738_,data_stage_2__7737_,
  data_stage_2__7736_,data_stage_2__7735_,data_stage_2__7734_,data_stage_2__7733_,
  data_stage_2__7732_,data_stage_2__7731_,data_stage_2__7730_,data_stage_2__7729_,
  data_stage_2__7728_,data_stage_2__7727_,data_stage_2__7726_,data_stage_2__7725_,
  data_stage_2__7724_,data_stage_2__7723_,data_stage_2__7722_,data_stage_2__7721_,
  data_stage_2__7720_,data_stage_2__7719_,data_stage_2__7718_,data_stage_2__7717_,
  data_stage_2__7716_,data_stage_2__7715_,data_stage_2__7714_,data_stage_2__7713_,
  data_stage_2__7712_,data_stage_2__7711_,data_stage_2__7710_,data_stage_2__7709_,
  data_stage_2__7708_,data_stage_2__7707_,data_stage_2__7706_,data_stage_2__7705_,
  data_stage_2__7704_,data_stage_2__7703_,data_stage_2__7702_,data_stage_2__7701_,
  data_stage_2__7700_,data_stage_2__7699_,data_stage_2__7698_,data_stage_2__7697_,
  data_stage_2__7696_,data_stage_2__7695_,data_stage_2__7694_,data_stage_2__7693_,
  data_stage_2__7692_,data_stage_2__7691_,data_stage_2__7690_,data_stage_2__7689_,
  data_stage_2__7688_,data_stage_2__7687_,data_stage_2__7686_,data_stage_2__7685_,
  data_stage_2__7684_,data_stage_2__7683_,data_stage_2__7682_,data_stage_2__7681_,
  data_stage_2__7680_,data_stage_2__7679_,data_stage_2__7678_,data_stage_2__7677_,
  data_stage_2__7676_,data_stage_2__7675_,data_stage_2__7674_,data_stage_2__7673_,
  data_stage_2__7672_,data_stage_2__7671_,data_stage_2__7670_,data_stage_2__7669_,
  data_stage_2__7668_,data_stage_2__7667_,data_stage_2__7666_,data_stage_2__7665_,
  data_stage_2__7664_,data_stage_2__7663_,data_stage_2__7662_,data_stage_2__7661_,
  data_stage_2__7660_,data_stage_2__7659_,data_stage_2__7658_,data_stage_2__7657_,
  data_stage_2__7656_,data_stage_2__7655_,data_stage_2__7654_,data_stage_2__7653_,
  data_stage_2__7652_,data_stage_2__7651_,data_stage_2__7650_,data_stage_2__7649_,
  data_stage_2__7648_,data_stage_2__7647_,data_stage_2__7646_,data_stage_2__7645_,
  data_stage_2__7644_,data_stage_2__7643_,data_stage_2__7642_,data_stage_2__7641_,
  data_stage_2__7640_,data_stage_2__7639_,data_stage_2__7638_,data_stage_2__7637_,
  data_stage_2__7636_,data_stage_2__7635_,data_stage_2__7634_,data_stage_2__7633_,
  data_stage_2__7632_,data_stage_2__7631_,data_stage_2__7630_,data_stage_2__7629_,
  data_stage_2__7628_,data_stage_2__7627_,data_stage_2__7626_,data_stage_2__7625_,
  data_stage_2__7624_,data_stage_2__7623_,data_stage_2__7622_,data_stage_2__7621_,
  data_stage_2__7620_,data_stage_2__7619_,data_stage_2__7618_,data_stage_2__7617_,
  data_stage_2__7616_,data_stage_2__7615_,data_stage_2__7614_,data_stage_2__7613_,
  data_stage_2__7612_,data_stage_2__7611_,data_stage_2__7610_,data_stage_2__7609_,
  data_stage_2__7608_,data_stage_2__7607_,data_stage_2__7606_,data_stage_2__7605_,
  data_stage_2__7604_,data_stage_2__7603_,data_stage_2__7602_,data_stage_2__7601_,
  data_stage_2__7600_,data_stage_2__7599_,data_stage_2__7598_,data_stage_2__7597_,
  data_stage_2__7596_,data_stage_2__7595_,data_stage_2__7594_,data_stage_2__7593_,
  data_stage_2__7592_,data_stage_2__7591_,data_stage_2__7590_,data_stage_2__7589_,
  data_stage_2__7588_,data_stage_2__7587_,data_stage_2__7586_,data_stage_2__7585_,
  data_stage_2__7584_,data_stage_2__7583_,data_stage_2__7582_,data_stage_2__7581_,
  data_stage_2__7580_,data_stage_2__7579_,data_stage_2__7578_,data_stage_2__7577_,
  data_stage_2__7576_,data_stage_2__7575_,data_stage_2__7574_,data_stage_2__7573_,
  data_stage_2__7572_,data_stage_2__7571_,data_stage_2__7570_,data_stage_2__7569_,
  data_stage_2__7568_,data_stage_2__7567_,data_stage_2__7566_,data_stage_2__7565_,
  data_stage_2__7564_,data_stage_2__7563_,data_stage_2__7562_,data_stage_2__7561_,
  data_stage_2__7560_,data_stage_2__7559_,data_stage_2__7558_,data_stage_2__7557_,
  data_stage_2__7556_,data_stage_2__7555_,data_stage_2__7554_,data_stage_2__7553_,
  data_stage_2__7552_,data_stage_2__7551_,data_stage_2__7550_,data_stage_2__7549_,
  data_stage_2__7548_,data_stage_2__7547_,data_stage_2__7546_,data_stage_2__7545_,
  data_stage_2__7544_,data_stage_2__7543_,data_stage_2__7542_,data_stage_2__7541_,
  data_stage_2__7540_,data_stage_2__7539_,data_stage_2__7538_,data_stage_2__7537_,
  data_stage_2__7536_,data_stage_2__7535_,data_stage_2__7534_,data_stage_2__7533_,
  data_stage_2__7532_,data_stage_2__7531_,data_stage_2__7530_,data_stage_2__7529_,
  data_stage_2__7528_,data_stage_2__7527_,data_stage_2__7526_,data_stage_2__7525_,
  data_stage_2__7524_,data_stage_2__7523_,data_stage_2__7522_,data_stage_2__7521_,
  data_stage_2__7520_,data_stage_2__7519_,data_stage_2__7518_,data_stage_2__7517_,
  data_stage_2__7516_,data_stage_2__7515_,data_stage_2__7514_,data_stage_2__7513_,
  data_stage_2__7512_,data_stage_2__7511_,data_stage_2__7510_,data_stage_2__7509_,
  data_stage_2__7508_,data_stage_2__7507_,data_stage_2__7506_,data_stage_2__7505_,
  data_stage_2__7504_,data_stage_2__7503_,data_stage_2__7502_,data_stage_2__7501_,
  data_stage_2__7500_,data_stage_2__7499_,data_stage_2__7498_,data_stage_2__7497_,
  data_stage_2__7496_,data_stage_2__7495_,data_stage_2__7494_,data_stage_2__7493_,
  data_stage_2__7492_,data_stage_2__7491_,data_stage_2__7490_,data_stage_2__7489_,
  data_stage_2__7488_,data_stage_2__7487_,data_stage_2__7486_,data_stage_2__7485_,
  data_stage_2__7484_,data_stage_2__7483_,data_stage_2__7482_,data_stage_2__7481_,
  data_stage_2__7480_,data_stage_2__7479_,data_stage_2__7478_,data_stage_2__7477_,
  data_stage_2__7476_,data_stage_2__7475_,data_stage_2__7474_,data_stage_2__7473_,
  data_stage_2__7472_,data_stage_2__7471_,data_stage_2__7470_,data_stage_2__7469_,
  data_stage_2__7468_,data_stage_2__7467_,data_stage_2__7466_,data_stage_2__7465_,
  data_stage_2__7464_,data_stage_2__7463_,data_stage_2__7462_,data_stage_2__7461_,
  data_stage_2__7460_,data_stage_2__7459_,data_stage_2__7458_,data_stage_2__7457_,
  data_stage_2__7456_,data_stage_2__7455_,data_stage_2__7454_,data_stage_2__7453_,
  data_stage_2__7452_,data_stage_2__7451_,data_stage_2__7450_,data_stage_2__7449_,
  data_stage_2__7448_,data_stage_2__7447_,data_stage_2__7446_,data_stage_2__7445_,
  data_stage_2__7444_,data_stage_2__7443_,data_stage_2__7442_,data_stage_2__7441_,
  data_stage_2__7440_,data_stage_2__7439_,data_stage_2__7438_,data_stage_2__7437_,
  data_stage_2__7436_,data_stage_2__7435_,data_stage_2__7434_,data_stage_2__7433_,
  data_stage_2__7432_,data_stage_2__7431_,data_stage_2__7430_,data_stage_2__7429_,
  data_stage_2__7428_,data_stage_2__7427_,data_stage_2__7426_,data_stage_2__7425_,
  data_stage_2__7424_,data_stage_2__7423_,data_stage_2__7422_,data_stage_2__7421_,
  data_stage_2__7420_,data_stage_2__7419_,data_stage_2__7418_,data_stage_2__7417_,
  data_stage_2__7416_,data_stage_2__7415_,data_stage_2__7414_,data_stage_2__7413_,
  data_stage_2__7412_,data_stage_2__7411_,data_stage_2__7410_,data_stage_2__7409_,
  data_stage_2__7408_,data_stage_2__7407_,data_stage_2__7406_,data_stage_2__7405_,
  data_stage_2__7404_,data_stage_2__7403_,data_stage_2__7402_,data_stage_2__7401_,
  data_stage_2__7400_,data_stage_2__7399_,data_stage_2__7398_,data_stage_2__7397_,
  data_stage_2__7396_,data_stage_2__7395_,data_stage_2__7394_,data_stage_2__7393_,
  data_stage_2__7392_,data_stage_2__7391_,data_stage_2__7390_,data_stage_2__7389_,
  data_stage_2__7388_,data_stage_2__7387_,data_stage_2__7386_,data_stage_2__7385_,
  data_stage_2__7384_,data_stage_2__7383_,data_stage_2__7382_,data_stage_2__7381_,
  data_stage_2__7380_,data_stage_2__7379_,data_stage_2__7378_,data_stage_2__7377_,
  data_stage_2__7376_,data_stage_2__7375_,data_stage_2__7374_,data_stage_2__7373_,
  data_stage_2__7372_,data_stage_2__7371_,data_stage_2__7370_,data_stage_2__7369_,
  data_stage_2__7368_,data_stage_2__7367_,data_stage_2__7366_,data_stage_2__7365_,
  data_stage_2__7364_,data_stage_2__7363_,data_stage_2__7362_,data_stage_2__7361_,
  data_stage_2__7360_,data_stage_2__7359_,data_stage_2__7358_,data_stage_2__7357_,
  data_stage_2__7356_,data_stage_2__7355_,data_stage_2__7354_,data_stage_2__7353_,
  data_stage_2__7352_,data_stage_2__7351_,data_stage_2__7350_,data_stage_2__7349_,
  data_stage_2__7348_,data_stage_2__7347_,data_stage_2__7346_,data_stage_2__7345_,
  data_stage_2__7344_,data_stage_2__7343_,data_stage_2__7342_,data_stage_2__7341_,
  data_stage_2__7340_,data_stage_2__7339_,data_stage_2__7338_,data_stage_2__7337_,
  data_stage_2__7336_,data_stage_2__7335_,data_stage_2__7334_,data_stage_2__7333_,
  data_stage_2__7332_,data_stage_2__7331_,data_stage_2__7330_,data_stage_2__7329_,
  data_stage_2__7328_,data_stage_2__7327_,data_stage_2__7326_,data_stage_2__7325_,
  data_stage_2__7324_,data_stage_2__7323_,data_stage_2__7322_,data_stage_2__7321_,
  data_stage_2__7320_,data_stage_2__7319_,data_stage_2__7318_,data_stage_2__7317_,
  data_stage_2__7316_,data_stage_2__7315_,data_stage_2__7314_,data_stage_2__7313_,
  data_stage_2__7312_,data_stage_2__7311_,data_stage_2__7310_,data_stage_2__7309_,
  data_stage_2__7308_,data_stage_2__7307_,data_stage_2__7306_,data_stage_2__7305_,
  data_stage_2__7304_,data_stage_2__7303_,data_stage_2__7302_,data_stage_2__7301_,
  data_stage_2__7300_,data_stage_2__7299_,data_stage_2__7298_,data_stage_2__7297_,
  data_stage_2__7296_,data_stage_2__7295_,data_stage_2__7294_,data_stage_2__7293_,
  data_stage_2__7292_,data_stage_2__7291_,data_stage_2__7290_,data_stage_2__7289_,
  data_stage_2__7288_,data_stage_2__7287_,data_stage_2__7286_,data_stage_2__7285_,
  data_stage_2__7284_,data_stage_2__7283_,data_stage_2__7282_,data_stage_2__7281_,
  data_stage_2__7280_,data_stage_2__7279_,data_stage_2__7278_,data_stage_2__7277_,
  data_stage_2__7276_,data_stage_2__7275_,data_stage_2__7274_,data_stage_2__7273_,
  data_stage_2__7272_,data_stage_2__7271_,data_stage_2__7270_,data_stage_2__7269_,
  data_stage_2__7268_,data_stage_2__7267_,data_stage_2__7266_,data_stage_2__7265_,
  data_stage_2__7264_,data_stage_2__7263_,data_stage_2__7262_,data_stage_2__7261_,
  data_stage_2__7260_,data_stage_2__7259_,data_stage_2__7258_,data_stage_2__7257_,
  data_stage_2__7256_,data_stage_2__7255_,data_stage_2__7254_,data_stage_2__7253_,
  data_stage_2__7252_,data_stage_2__7251_,data_stage_2__7250_,data_stage_2__7249_,
  data_stage_2__7248_,data_stage_2__7247_,data_stage_2__7246_,data_stage_2__7245_,
  data_stage_2__7244_,data_stage_2__7243_,data_stage_2__7242_,data_stage_2__7241_,
  data_stage_2__7240_,data_stage_2__7239_,data_stage_2__7238_,data_stage_2__7237_,
  data_stage_2__7236_,data_stage_2__7235_,data_stage_2__7234_,data_stage_2__7233_,
  data_stage_2__7232_,data_stage_2__7231_,data_stage_2__7230_,data_stage_2__7229_,
  data_stage_2__7228_,data_stage_2__7227_,data_stage_2__7226_,data_stage_2__7225_,
  data_stage_2__7224_,data_stage_2__7223_,data_stage_2__7222_,data_stage_2__7221_,
  data_stage_2__7220_,data_stage_2__7219_,data_stage_2__7218_,data_stage_2__7217_,
  data_stage_2__7216_,data_stage_2__7215_,data_stage_2__7214_,data_stage_2__7213_,
  data_stage_2__7212_,data_stage_2__7211_,data_stage_2__7210_,data_stage_2__7209_,
  data_stage_2__7208_,data_stage_2__7207_,data_stage_2__7206_,data_stage_2__7205_,
  data_stage_2__7204_,data_stage_2__7203_,data_stage_2__7202_,data_stage_2__7201_,
  data_stage_2__7200_,data_stage_2__7199_,data_stage_2__7198_,data_stage_2__7197_,
  data_stage_2__7196_,data_stage_2__7195_,data_stage_2__7194_,data_stage_2__7193_,
  data_stage_2__7192_,data_stage_2__7191_,data_stage_2__7190_,data_stage_2__7189_,
  data_stage_2__7188_,data_stage_2__7187_,data_stage_2__7186_,data_stage_2__7185_,
  data_stage_2__7184_,data_stage_2__7183_,data_stage_2__7182_,data_stage_2__7181_,
  data_stage_2__7180_,data_stage_2__7179_,data_stage_2__7178_,data_stage_2__7177_,
  data_stage_2__7176_,data_stage_2__7175_,data_stage_2__7174_,data_stage_2__7173_,
  data_stage_2__7172_,data_stage_2__7171_,data_stage_2__7170_,data_stage_2__7169_,
  data_stage_2__7168_,data_stage_2__7167_,data_stage_2__7166_,data_stage_2__7165_,
  data_stage_2__7164_,data_stage_2__7163_,data_stage_2__7162_,data_stage_2__7161_,
  data_stage_2__7160_,data_stage_2__7159_,data_stage_2__7158_,data_stage_2__7157_,
  data_stage_2__7156_,data_stage_2__7155_,data_stage_2__7154_,data_stage_2__7153_,
  data_stage_2__7152_,data_stage_2__7151_,data_stage_2__7150_,data_stage_2__7149_,
  data_stage_2__7148_,data_stage_2__7147_,data_stage_2__7146_,data_stage_2__7145_,
  data_stage_2__7144_,data_stage_2__7143_,data_stage_2__7142_,data_stage_2__7141_,
  data_stage_2__7140_,data_stage_2__7139_,data_stage_2__7138_,data_stage_2__7137_,
  data_stage_2__7136_,data_stage_2__7135_,data_stage_2__7134_,data_stage_2__7133_,
  data_stage_2__7132_,data_stage_2__7131_,data_stage_2__7130_,data_stage_2__7129_,
  data_stage_2__7128_,data_stage_2__7127_,data_stage_2__7126_,data_stage_2__7125_,
  data_stage_2__7124_,data_stage_2__7123_,data_stage_2__7122_,data_stage_2__7121_,
  data_stage_2__7120_,data_stage_2__7119_,data_stage_2__7118_,data_stage_2__7117_,
  data_stage_2__7116_,data_stage_2__7115_,data_stage_2__7114_,data_stage_2__7113_,
  data_stage_2__7112_,data_stage_2__7111_,data_stage_2__7110_,data_stage_2__7109_,
  data_stage_2__7108_,data_stage_2__7107_,data_stage_2__7106_,data_stage_2__7105_,
  data_stage_2__7104_,data_stage_2__7103_,data_stage_2__7102_,data_stage_2__7101_,
  data_stage_2__7100_,data_stage_2__7099_,data_stage_2__7098_,data_stage_2__7097_,
  data_stage_2__7096_,data_stage_2__7095_,data_stage_2__7094_,data_stage_2__7093_,
  data_stage_2__7092_,data_stage_2__7091_,data_stage_2__7090_,data_stage_2__7089_,
  data_stage_2__7088_,data_stage_2__7087_,data_stage_2__7086_,data_stage_2__7085_,
  data_stage_2__7084_,data_stage_2__7083_,data_stage_2__7082_,data_stage_2__7081_,
  data_stage_2__7080_,data_stage_2__7079_,data_stage_2__7078_,data_stage_2__7077_,
  data_stage_2__7076_,data_stage_2__7075_,data_stage_2__7074_,data_stage_2__7073_,
  data_stage_2__7072_,data_stage_2__7071_,data_stage_2__7070_,data_stage_2__7069_,
  data_stage_2__7068_,data_stage_2__7067_,data_stage_2__7066_,data_stage_2__7065_,
  data_stage_2__7064_,data_stage_2__7063_,data_stage_2__7062_,data_stage_2__7061_,
  data_stage_2__7060_,data_stage_2__7059_,data_stage_2__7058_,data_stage_2__7057_,
  data_stage_2__7056_,data_stage_2__7055_,data_stage_2__7054_,data_stage_2__7053_,
  data_stage_2__7052_,data_stage_2__7051_,data_stage_2__7050_,data_stage_2__7049_,
  data_stage_2__7048_,data_stage_2__7047_,data_stage_2__7046_,data_stage_2__7045_,
  data_stage_2__7044_,data_stage_2__7043_,data_stage_2__7042_,data_stage_2__7041_,
  data_stage_2__7040_,data_stage_2__7039_,data_stage_2__7038_,data_stage_2__7037_,
  data_stage_2__7036_,data_stage_2__7035_,data_stage_2__7034_,data_stage_2__7033_,
  data_stage_2__7032_,data_stage_2__7031_,data_stage_2__7030_,data_stage_2__7029_,
  data_stage_2__7028_,data_stage_2__7027_,data_stage_2__7026_,data_stage_2__7025_,
  data_stage_2__7024_,data_stage_2__7023_,data_stage_2__7022_,data_stage_2__7021_,
  data_stage_2__7020_,data_stage_2__7019_,data_stage_2__7018_,data_stage_2__7017_,
  data_stage_2__7016_,data_stage_2__7015_,data_stage_2__7014_,data_stage_2__7013_,
  data_stage_2__7012_,data_stage_2__7011_,data_stage_2__7010_,data_stage_2__7009_,
  data_stage_2__7008_,data_stage_2__7007_,data_stage_2__7006_,data_stage_2__7005_,
  data_stage_2__7004_,data_stage_2__7003_,data_stage_2__7002_,data_stage_2__7001_,
  data_stage_2__7000_,data_stage_2__6999_,data_stage_2__6998_,data_stage_2__6997_,
  data_stage_2__6996_,data_stage_2__6995_,data_stage_2__6994_,data_stage_2__6993_,
  data_stage_2__6992_,data_stage_2__6991_,data_stage_2__6990_,data_stage_2__6989_,
  data_stage_2__6988_,data_stage_2__6987_,data_stage_2__6986_,data_stage_2__6985_,
  data_stage_2__6984_,data_stage_2__6983_,data_stage_2__6982_,data_stage_2__6981_,
  data_stage_2__6980_,data_stage_2__6979_,data_stage_2__6978_,data_stage_2__6977_,
  data_stage_2__6976_,data_stage_2__6975_,data_stage_2__6974_,data_stage_2__6973_,
  data_stage_2__6972_,data_stage_2__6971_,data_stage_2__6970_,data_stage_2__6969_,
  data_stage_2__6968_,data_stage_2__6967_,data_stage_2__6966_,data_stage_2__6965_,
  data_stage_2__6964_,data_stage_2__6963_,data_stage_2__6962_,data_stage_2__6961_,
  data_stage_2__6960_,data_stage_2__6959_,data_stage_2__6958_,data_stage_2__6957_,
  data_stage_2__6956_,data_stage_2__6955_,data_stage_2__6954_,data_stage_2__6953_,
  data_stage_2__6952_,data_stage_2__6951_,data_stage_2__6950_,data_stage_2__6949_,
  data_stage_2__6948_,data_stage_2__6947_,data_stage_2__6946_,data_stage_2__6945_,
  data_stage_2__6944_,data_stage_2__6943_,data_stage_2__6942_,data_stage_2__6941_,
  data_stage_2__6940_,data_stage_2__6939_,data_stage_2__6938_,data_stage_2__6937_,
  data_stage_2__6936_,data_stage_2__6935_,data_stage_2__6934_,data_stage_2__6933_,
  data_stage_2__6932_,data_stage_2__6931_,data_stage_2__6930_,data_stage_2__6929_,
  data_stage_2__6928_,data_stage_2__6927_,data_stage_2__6926_,data_stage_2__6925_,
  data_stage_2__6924_,data_stage_2__6923_,data_stage_2__6922_,data_stage_2__6921_,
  data_stage_2__6920_,data_stage_2__6919_,data_stage_2__6918_,data_stage_2__6917_,
  data_stage_2__6916_,data_stage_2__6915_,data_stage_2__6914_,data_stage_2__6913_,
  data_stage_2__6912_,data_stage_2__6911_,data_stage_2__6910_,data_stage_2__6909_,
  data_stage_2__6908_,data_stage_2__6907_,data_stage_2__6906_,data_stage_2__6905_,
  data_stage_2__6904_,data_stage_2__6903_,data_stage_2__6902_,data_stage_2__6901_,
  data_stage_2__6900_,data_stage_2__6899_,data_stage_2__6898_,data_stage_2__6897_,
  data_stage_2__6896_,data_stage_2__6895_,data_stage_2__6894_,data_stage_2__6893_,
  data_stage_2__6892_,data_stage_2__6891_,data_stage_2__6890_,data_stage_2__6889_,
  data_stage_2__6888_,data_stage_2__6887_,data_stage_2__6886_,data_stage_2__6885_,
  data_stage_2__6884_,data_stage_2__6883_,data_stage_2__6882_,data_stage_2__6881_,
  data_stage_2__6880_,data_stage_2__6879_,data_stage_2__6878_,data_stage_2__6877_,
  data_stage_2__6876_,data_stage_2__6875_,data_stage_2__6874_,data_stage_2__6873_,
  data_stage_2__6872_,data_stage_2__6871_,data_stage_2__6870_,data_stage_2__6869_,
  data_stage_2__6868_,data_stage_2__6867_,data_stage_2__6866_,data_stage_2__6865_,
  data_stage_2__6864_,data_stage_2__6863_,data_stage_2__6862_,data_stage_2__6861_,
  data_stage_2__6860_,data_stage_2__6859_,data_stage_2__6858_,data_stage_2__6857_,
  data_stage_2__6856_,data_stage_2__6855_,data_stage_2__6854_,data_stage_2__6853_,
  data_stage_2__6852_,data_stage_2__6851_,data_stage_2__6850_,data_stage_2__6849_,
  data_stage_2__6848_,data_stage_2__6847_,data_stage_2__6846_,data_stage_2__6845_,
  data_stage_2__6844_,data_stage_2__6843_,data_stage_2__6842_,data_stage_2__6841_,
  data_stage_2__6840_,data_stage_2__6839_,data_stage_2__6838_,data_stage_2__6837_,
  data_stage_2__6836_,data_stage_2__6835_,data_stage_2__6834_,data_stage_2__6833_,
  data_stage_2__6832_,data_stage_2__6831_,data_stage_2__6830_,data_stage_2__6829_,
  data_stage_2__6828_,data_stage_2__6827_,data_stage_2__6826_,data_stage_2__6825_,
  data_stage_2__6824_,data_stage_2__6823_,data_stage_2__6822_,data_stage_2__6821_,
  data_stage_2__6820_,data_stage_2__6819_,data_stage_2__6818_,data_stage_2__6817_,
  data_stage_2__6816_,data_stage_2__6815_,data_stage_2__6814_,data_stage_2__6813_,
  data_stage_2__6812_,data_stage_2__6811_,data_stage_2__6810_,data_stage_2__6809_,
  data_stage_2__6808_,data_stage_2__6807_,data_stage_2__6806_,data_stage_2__6805_,
  data_stage_2__6804_,data_stage_2__6803_,data_stage_2__6802_,data_stage_2__6801_,
  data_stage_2__6800_,data_stage_2__6799_,data_stage_2__6798_,data_stage_2__6797_,
  data_stage_2__6796_,data_stage_2__6795_,data_stage_2__6794_,data_stage_2__6793_,
  data_stage_2__6792_,data_stage_2__6791_,data_stage_2__6790_,data_stage_2__6789_,
  data_stage_2__6788_,data_stage_2__6787_,data_stage_2__6786_,data_stage_2__6785_,
  data_stage_2__6784_,data_stage_2__6783_,data_stage_2__6782_,data_stage_2__6781_,
  data_stage_2__6780_,data_stage_2__6779_,data_stage_2__6778_,data_stage_2__6777_,
  data_stage_2__6776_,data_stage_2__6775_,data_stage_2__6774_,data_stage_2__6773_,
  data_stage_2__6772_,data_stage_2__6771_,data_stage_2__6770_,data_stage_2__6769_,
  data_stage_2__6768_,data_stage_2__6767_,data_stage_2__6766_,data_stage_2__6765_,
  data_stage_2__6764_,data_stage_2__6763_,data_stage_2__6762_,data_stage_2__6761_,
  data_stage_2__6760_,data_stage_2__6759_,data_stage_2__6758_,data_stage_2__6757_,
  data_stage_2__6756_,data_stage_2__6755_,data_stage_2__6754_,data_stage_2__6753_,
  data_stage_2__6752_,data_stage_2__6751_,data_stage_2__6750_,data_stage_2__6749_,
  data_stage_2__6748_,data_stage_2__6747_,data_stage_2__6746_,data_stage_2__6745_,
  data_stage_2__6744_,data_stage_2__6743_,data_stage_2__6742_,data_stage_2__6741_,
  data_stage_2__6740_,data_stage_2__6739_,data_stage_2__6738_,data_stage_2__6737_,
  data_stage_2__6736_,data_stage_2__6735_,data_stage_2__6734_,data_stage_2__6733_,
  data_stage_2__6732_,data_stage_2__6731_,data_stage_2__6730_,data_stage_2__6729_,
  data_stage_2__6728_,data_stage_2__6727_,data_stage_2__6726_,data_stage_2__6725_,
  data_stage_2__6724_,data_stage_2__6723_,data_stage_2__6722_,data_stage_2__6721_,
  data_stage_2__6720_,data_stage_2__6719_,data_stage_2__6718_,data_stage_2__6717_,
  data_stage_2__6716_,data_stage_2__6715_,data_stage_2__6714_,data_stage_2__6713_,
  data_stage_2__6712_,data_stage_2__6711_,data_stage_2__6710_,data_stage_2__6709_,
  data_stage_2__6708_,data_stage_2__6707_,data_stage_2__6706_,data_stage_2__6705_,
  data_stage_2__6704_,data_stage_2__6703_,data_stage_2__6702_,data_stage_2__6701_,
  data_stage_2__6700_,data_stage_2__6699_,data_stage_2__6698_,data_stage_2__6697_,
  data_stage_2__6696_,data_stage_2__6695_,data_stage_2__6694_,data_stage_2__6693_,
  data_stage_2__6692_,data_stage_2__6691_,data_stage_2__6690_,data_stage_2__6689_,
  data_stage_2__6688_,data_stage_2__6687_,data_stage_2__6686_,data_stage_2__6685_,
  data_stage_2__6684_,data_stage_2__6683_,data_stage_2__6682_,data_stage_2__6681_,
  data_stage_2__6680_,data_stage_2__6679_,data_stage_2__6678_,data_stage_2__6677_,
  data_stage_2__6676_,data_stage_2__6675_,data_stage_2__6674_,data_stage_2__6673_,
  data_stage_2__6672_,data_stage_2__6671_,data_stage_2__6670_,data_stage_2__6669_,
  data_stage_2__6668_,data_stage_2__6667_,data_stage_2__6666_,data_stage_2__6665_,
  data_stage_2__6664_,data_stage_2__6663_,data_stage_2__6662_,data_stage_2__6661_,
  data_stage_2__6660_,data_stage_2__6659_,data_stage_2__6658_,data_stage_2__6657_,
  data_stage_2__6656_,data_stage_2__6655_,data_stage_2__6654_,data_stage_2__6653_,
  data_stage_2__6652_,data_stage_2__6651_,data_stage_2__6650_,data_stage_2__6649_,
  data_stage_2__6648_,data_stage_2__6647_,data_stage_2__6646_,data_stage_2__6645_,
  data_stage_2__6644_,data_stage_2__6643_,data_stage_2__6642_,data_stage_2__6641_,
  data_stage_2__6640_,data_stage_2__6639_,data_stage_2__6638_,data_stage_2__6637_,
  data_stage_2__6636_,data_stage_2__6635_,data_stage_2__6634_,data_stage_2__6633_,
  data_stage_2__6632_,data_stage_2__6631_,data_stage_2__6630_,data_stage_2__6629_,
  data_stage_2__6628_,data_stage_2__6627_,data_stage_2__6626_,data_stage_2__6625_,
  data_stage_2__6624_,data_stage_2__6623_,data_stage_2__6622_,data_stage_2__6621_,
  data_stage_2__6620_,data_stage_2__6619_,data_stage_2__6618_,data_stage_2__6617_,
  data_stage_2__6616_,data_stage_2__6615_,data_stage_2__6614_,data_stage_2__6613_,
  data_stage_2__6612_,data_stage_2__6611_,data_stage_2__6610_,data_stage_2__6609_,
  data_stage_2__6608_,data_stage_2__6607_,data_stage_2__6606_,data_stage_2__6605_,
  data_stage_2__6604_,data_stage_2__6603_,data_stage_2__6602_,data_stage_2__6601_,
  data_stage_2__6600_,data_stage_2__6599_,data_stage_2__6598_,data_stage_2__6597_,
  data_stage_2__6596_,data_stage_2__6595_,data_stage_2__6594_,data_stage_2__6593_,
  data_stage_2__6592_,data_stage_2__6591_,data_stage_2__6590_,data_stage_2__6589_,
  data_stage_2__6588_,data_stage_2__6587_,data_stage_2__6586_,data_stage_2__6585_,
  data_stage_2__6584_,data_stage_2__6583_,data_stage_2__6582_,data_stage_2__6581_,
  data_stage_2__6580_,data_stage_2__6579_,data_stage_2__6578_,data_stage_2__6577_,
  data_stage_2__6576_,data_stage_2__6575_,data_stage_2__6574_,data_stage_2__6573_,
  data_stage_2__6572_,data_stage_2__6571_,data_stage_2__6570_,data_stage_2__6569_,
  data_stage_2__6568_,data_stage_2__6567_,data_stage_2__6566_,data_stage_2__6565_,
  data_stage_2__6564_,data_stage_2__6563_,data_stage_2__6562_,data_stage_2__6561_,
  data_stage_2__6560_,data_stage_2__6559_,data_stage_2__6558_,data_stage_2__6557_,
  data_stage_2__6556_,data_stage_2__6555_,data_stage_2__6554_,data_stage_2__6553_,
  data_stage_2__6552_,data_stage_2__6551_,data_stage_2__6550_,data_stage_2__6549_,
  data_stage_2__6548_,data_stage_2__6547_,data_stage_2__6546_,data_stage_2__6545_,
  data_stage_2__6544_,data_stage_2__6543_,data_stage_2__6542_,data_stage_2__6541_,
  data_stage_2__6540_,data_stage_2__6539_,data_stage_2__6538_,data_stage_2__6537_,
  data_stage_2__6536_,data_stage_2__6535_,data_stage_2__6534_,data_stage_2__6533_,
  data_stage_2__6532_,data_stage_2__6531_,data_stage_2__6530_,data_stage_2__6529_,
  data_stage_2__6528_,data_stage_2__6527_,data_stage_2__6526_,data_stage_2__6525_,
  data_stage_2__6524_,data_stage_2__6523_,data_stage_2__6522_,data_stage_2__6521_,
  data_stage_2__6520_,data_stage_2__6519_,data_stage_2__6518_,data_stage_2__6517_,
  data_stage_2__6516_,data_stage_2__6515_,data_stage_2__6514_,data_stage_2__6513_,
  data_stage_2__6512_,data_stage_2__6511_,data_stage_2__6510_,data_stage_2__6509_,
  data_stage_2__6508_,data_stage_2__6507_,data_stage_2__6506_,data_stage_2__6505_,
  data_stage_2__6504_,data_stage_2__6503_,data_stage_2__6502_,data_stage_2__6501_,
  data_stage_2__6500_,data_stage_2__6499_,data_stage_2__6498_,data_stage_2__6497_,
  data_stage_2__6496_,data_stage_2__6495_,data_stage_2__6494_,data_stage_2__6493_,
  data_stage_2__6492_,data_stage_2__6491_,data_stage_2__6490_,data_stage_2__6489_,
  data_stage_2__6488_,data_stage_2__6487_,data_stage_2__6486_,data_stage_2__6485_,
  data_stage_2__6484_,data_stage_2__6483_,data_stage_2__6482_,data_stage_2__6481_,
  data_stage_2__6480_,data_stage_2__6479_,data_stage_2__6478_,data_stage_2__6477_,
  data_stage_2__6476_,data_stage_2__6475_,data_stage_2__6474_,data_stage_2__6473_,
  data_stage_2__6472_,data_stage_2__6471_,data_stage_2__6470_,data_stage_2__6469_,
  data_stage_2__6468_,data_stage_2__6467_,data_stage_2__6466_,data_stage_2__6465_,
  data_stage_2__6464_,data_stage_2__6463_,data_stage_2__6462_,data_stage_2__6461_,
  data_stage_2__6460_,data_stage_2__6459_,data_stage_2__6458_,data_stage_2__6457_,
  data_stage_2__6456_,data_stage_2__6455_,data_stage_2__6454_,data_stage_2__6453_,
  data_stage_2__6452_,data_stage_2__6451_,data_stage_2__6450_,data_stage_2__6449_,
  data_stage_2__6448_,data_stage_2__6447_,data_stage_2__6446_,data_stage_2__6445_,
  data_stage_2__6444_,data_stage_2__6443_,data_stage_2__6442_,data_stage_2__6441_,
  data_stage_2__6440_,data_stage_2__6439_,data_stage_2__6438_,data_stage_2__6437_,
  data_stage_2__6436_,data_stage_2__6435_,data_stage_2__6434_,data_stage_2__6433_,
  data_stage_2__6432_,data_stage_2__6431_,data_stage_2__6430_,data_stage_2__6429_,
  data_stage_2__6428_,data_stage_2__6427_,data_stage_2__6426_,data_stage_2__6425_,
  data_stage_2__6424_,data_stage_2__6423_,data_stage_2__6422_,data_stage_2__6421_,
  data_stage_2__6420_,data_stage_2__6419_,data_stage_2__6418_,data_stage_2__6417_,
  data_stage_2__6416_,data_stage_2__6415_,data_stage_2__6414_,data_stage_2__6413_,
  data_stage_2__6412_,data_stage_2__6411_,data_stage_2__6410_,data_stage_2__6409_,
  data_stage_2__6408_,data_stage_2__6407_,data_stage_2__6406_,data_stage_2__6405_,
  data_stage_2__6404_,data_stage_2__6403_,data_stage_2__6402_,data_stage_2__6401_,
  data_stage_2__6400_,data_stage_2__6399_,data_stage_2__6398_,data_stage_2__6397_,
  data_stage_2__6396_,data_stage_2__6395_,data_stage_2__6394_,data_stage_2__6393_,
  data_stage_2__6392_,data_stage_2__6391_,data_stage_2__6390_,data_stage_2__6389_,
  data_stage_2__6388_,data_stage_2__6387_,data_stage_2__6386_,data_stage_2__6385_,
  data_stage_2__6384_,data_stage_2__6383_,data_stage_2__6382_,data_stage_2__6381_,
  data_stage_2__6380_,data_stage_2__6379_,data_stage_2__6378_,data_stage_2__6377_,
  data_stage_2__6376_,data_stage_2__6375_,data_stage_2__6374_,data_stage_2__6373_,
  data_stage_2__6372_,data_stage_2__6371_,data_stage_2__6370_,data_stage_2__6369_,
  data_stage_2__6368_,data_stage_2__6367_,data_stage_2__6366_,data_stage_2__6365_,
  data_stage_2__6364_,data_stage_2__6363_,data_stage_2__6362_,data_stage_2__6361_,
  data_stage_2__6360_,data_stage_2__6359_,data_stage_2__6358_,data_stage_2__6357_,
  data_stage_2__6356_,data_stage_2__6355_,data_stage_2__6354_,data_stage_2__6353_,
  data_stage_2__6352_,data_stage_2__6351_,data_stage_2__6350_,data_stage_2__6349_,
  data_stage_2__6348_,data_stage_2__6347_,data_stage_2__6346_,data_stage_2__6345_,
  data_stage_2__6344_,data_stage_2__6343_,data_stage_2__6342_,data_stage_2__6341_,
  data_stage_2__6340_,data_stage_2__6339_,data_stage_2__6338_,data_stage_2__6337_,
  data_stage_2__6336_,data_stage_2__6335_,data_stage_2__6334_,data_stage_2__6333_,
  data_stage_2__6332_,data_stage_2__6331_,data_stage_2__6330_,data_stage_2__6329_,
  data_stage_2__6328_,data_stage_2__6327_,data_stage_2__6326_,data_stage_2__6325_,
  data_stage_2__6324_,data_stage_2__6323_,data_stage_2__6322_,data_stage_2__6321_,
  data_stage_2__6320_,data_stage_2__6319_,data_stage_2__6318_,data_stage_2__6317_,
  data_stage_2__6316_,data_stage_2__6315_,data_stage_2__6314_,data_stage_2__6313_,
  data_stage_2__6312_,data_stage_2__6311_,data_stage_2__6310_,data_stage_2__6309_,
  data_stage_2__6308_,data_stage_2__6307_,data_stage_2__6306_,data_stage_2__6305_,
  data_stage_2__6304_,data_stage_2__6303_,data_stage_2__6302_,data_stage_2__6301_,
  data_stage_2__6300_,data_stage_2__6299_,data_stage_2__6298_,data_stage_2__6297_,
  data_stage_2__6296_,data_stage_2__6295_,data_stage_2__6294_,data_stage_2__6293_,
  data_stage_2__6292_,data_stage_2__6291_,data_stage_2__6290_,data_stage_2__6289_,
  data_stage_2__6288_,data_stage_2__6287_,data_stage_2__6286_,data_stage_2__6285_,
  data_stage_2__6284_,data_stage_2__6283_,data_stage_2__6282_,data_stage_2__6281_,
  data_stage_2__6280_,data_stage_2__6279_,data_stage_2__6278_,data_stage_2__6277_,
  data_stage_2__6276_,data_stage_2__6275_,data_stage_2__6274_,data_stage_2__6273_,
  data_stage_2__6272_,data_stage_2__6271_,data_stage_2__6270_,data_stage_2__6269_,
  data_stage_2__6268_,data_stage_2__6267_,data_stage_2__6266_,data_stage_2__6265_,
  data_stage_2__6264_,data_stage_2__6263_,data_stage_2__6262_,data_stage_2__6261_,
  data_stage_2__6260_,data_stage_2__6259_,data_stage_2__6258_,data_stage_2__6257_,
  data_stage_2__6256_,data_stage_2__6255_,data_stage_2__6254_,data_stage_2__6253_,
  data_stage_2__6252_,data_stage_2__6251_,data_stage_2__6250_,data_stage_2__6249_,
  data_stage_2__6248_,data_stage_2__6247_,data_stage_2__6246_,data_stage_2__6245_,
  data_stage_2__6244_,data_stage_2__6243_,data_stage_2__6242_,data_stage_2__6241_,
  data_stage_2__6240_,data_stage_2__6239_,data_stage_2__6238_,data_stage_2__6237_,
  data_stage_2__6236_,data_stage_2__6235_,data_stage_2__6234_,data_stage_2__6233_,
  data_stage_2__6232_,data_stage_2__6231_,data_stage_2__6230_,data_stage_2__6229_,
  data_stage_2__6228_,data_stage_2__6227_,data_stage_2__6226_,data_stage_2__6225_,
  data_stage_2__6224_,data_stage_2__6223_,data_stage_2__6222_,data_stage_2__6221_,
  data_stage_2__6220_,data_stage_2__6219_,data_stage_2__6218_,data_stage_2__6217_,
  data_stage_2__6216_,data_stage_2__6215_,data_stage_2__6214_,data_stage_2__6213_,
  data_stage_2__6212_,data_stage_2__6211_,data_stage_2__6210_,data_stage_2__6209_,
  data_stage_2__6208_,data_stage_2__6207_,data_stage_2__6206_,data_stage_2__6205_,
  data_stage_2__6204_,data_stage_2__6203_,data_stage_2__6202_,data_stage_2__6201_,
  data_stage_2__6200_,data_stage_2__6199_,data_stage_2__6198_,data_stage_2__6197_,
  data_stage_2__6196_,data_stage_2__6195_,data_stage_2__6194_,data_stage_2__6193_,
  data_stage_2__6192_,data_stage_2__6191_,data_stage_2__6190_,data_stage_2__6189_,
  data_stage_2__6188_,data_stage_2__6187_,data_stage_2__6186_,data_stage_2__6185_,
  data_stage_2__6184_,data_stage_2__6183_,data_stage_2__6182_,data_stage_2__6181_,
  data_stage_2__6180_,data_stage_2__6179_,data_stage_2__6178_,data_stage_2__6177_,
  data_stage_2__6176_,data_stage_2__6175_,data_stage_2__6174_,data_stage_2__6173_,
  data_stage_2__6172_,data_stage_2__6171_,data_stage_2__6170_,data_stage_2__6169_,
  data_stage_2__6168_,data_stage_2__6167_,data_stage_2__6166_,data_stage_2__6165_,
  data_stage_2__6164_,data_stage_2__6163_,data_stage_2__6162_,data_stage_2__6161_,
  data_stage_2__6160_,data_stage_2__6159_,data_stage_2__6158_,data_stage_2__6157_,
  data_stage_2__6156_,data_stage_2__6155_,data_stage_2__6154_,data_stage_2__6153_,
  data_stage_2__6152_,data_stage_2__6151_,data_stage_2__6150_,data_stage_2__6149_,
  data_stage_2__6148_,data_stage_2__6147_,data_stage_2__6146_,data_stage_2__6145_,
  data_stage_2__6144_,data_stage_2__6143_,data_stage_2__6142_,data_stage_2__6141_,
  data_stage_2__6140_,data_stage_2__6139_,data_stage_2__6138_,data_stage_2__6137_,
  data_stage_2__6136_,data_stage_2__6135_,data_stage_2__6134_,data_stage_2__6133_,
  data_stage_2__6132_,data_stage_2__6131_,data_stage_2__6130_,data_stage_2__6129_,
  data_stage_2__6128_,data_stage_2__6127_,data_stage_2__6126_,data_stage_2__6125_,
  data_stage_2__6124_,data_stage_2__6123_,data_stage_2__6122_,data_stage_2__6121_,
  data_stage_2__6120_,data_stage_2__6119_,data_stage_2__6118_,data_stage_2__6117_,
  data_stage_2__6116_,data_stage_2__6115_,data_stage_2__6114_,data_stage_2__6113_,
  data_stage_2__6112_,data_stage_2__6111_,data_stage_2__6110_,data_stage_2__6109_,
  data_stage_2__6108_,data_stage_2__6107_,data_stage_2__6106_,data_stage_2__6105_,
  data_stage_2__6104_,data_stage_2__6103_,data_stage_2__6102_,data_stage_2__6101_,
  data_stage_2__6100_,data_stage_2__6099_,data_stage_2__6098_,data_stage_2__6097_,
  data_stage_2__6096_,data_stage_2__6095_,data_stage_2__6094_,data_stage_2__6093_,
  data_stage_2__6092_,data_stage_2__6091_,data_stage_2__6090_,data_stage_2__6089_,
  data_stage_2__6088_,data_stage_2__6087_,data_stage_2__6086_,data_stage_2__6085_,
  data_stage_2__6084_,data_stage_2__6083_,data_stage_2__6082_,data_stage_2__6081_,
  data_stage_2__6080_,data_stage_2__6079_,data_stage_2__6078_,data_stage_2__6077_,
  data_stage_2__6076_,data_stage_2__6075_,data_stage_2__6074_,data_stage_2__6073_,
  data_stage_2__6072_,data_stage_2__6071_,data_stage_2__6070_,data_stage_2__6069_,
  data_stage_2__6068_,data_stage_2__6067_,data_stage_2__6066_,data_stage_2__6065_,
  data_stage_2__6064_,data_stage_2__6063_,data_stage_2__6062_,data_stage_2__6061_,
  data_stage_2__6060_,data_stage_2__6059_,data_stage_2__6058_,data_stage_2__6057_,
  data_stage_2__6056_,data_stage_2__6055_,data_stage_2__6054_,data_stage_2__6053_,
  data_stage_2__6052_,data_stage_2__6051_,data_stage_2__6050_,data_stage_2__6049_,
  data_stage_2__6048_,data_stage_2__6047_,data_stage_2__6046_,data_stage_2__6045_,
  data_stage_2__6044_,data_stage_2__6043_,data_stage_2__6042_,data_stage_2__6041_,
  data_stage_2__6040_,data_stage_2__6039_,data_stage_2__6038_,data_stage_2__6037_,
  data_stage_2__6036_,data_stage_2__6035_,data_stage_2__6034_,data_stage_2__6033_,
  data_stage_2__6032_,data_stage_2__6031_,data_stage_2__6030_,data_stage_2__6029_,
  data_stage_2__6028_,data_stage_2__6027_,data_stage_2__6026_,data_stage_2__6025_,
  data_stage_2__6024_,data_stage_2__6023_,data_stage_2__6022_,data_stage_2__6021_,
  data_stage_2__6020_,data_stage_2__6019_,data_stage_2__6018_,data_stage_2__6017_,
  data_stage_2__6016_,data_stage_2__6015_,data_stage_2__6014_,data_stage_2__6013_,
  data_stage_2__6012_,data_stage_2__6011_,data_stage_2__6010_,data_stage_2__6009_,
  data_stage_2__6008_,data_stage_2__6007_,data_stage_2__6006_,data_stage_2__6005_,
  data_stage_2__6004_,data_stage_2__6003_,data_stage_2__6002_,data_stage_2__6001_,
  data_stage_2__6000_,data_stage_2__5999_,data_stage_2__5998_,data_stage_2__5997_,
  data_stage_2__5996_,data_stage_2__5995_,data_stage_2__5994_,data_stage_2__5993_,
  data_stage_2__5992_,data_stage_2__5991_,data_stage_2__5990_,data_stage_2__5989_,
  data_stage_2__5988_,data_stage_2__5987_,data_stage_2__5986_,data_stage_2__5985_,
  data_stage_2__5984_,data_stage_2__5983_,data_stage_2__5982_,data_stage_2__5981_,
  data_stage_2__5980_,data_stage_2__5979_,data_stage_2__5978_,data_stage_2__5977_,
  data_stage_2__5976_,data_stage_2__5975_,data_stage_2__5974_,data_stage_2__5973_,
  data_stage_2__5972_,data_stage_2__5971_,data_stage_2__5970_,data_stage_2__5969_,
  data_stage_2__5968_,data_stage_2__5967_,data_stage_2__5966_,data_stage_2__5965_,
  data_stage_2__5964_,data_stage_2__5963_,data_stage_2__5962_,data_stage_2__5961_,
  data_stage_2__5960_,data_stage_2__5959_,data_stage_2__5958_,data_stage_2__5957_,
  data_stage_2__5956_,data_stage_2__5955_,data_stage_2__5954_,data_stage_2__5953_,
  data_stage_2__5952_,data_stage_2__5951_,data_stage_2__5950_,data_stage_2__5949_,
  data_stage_2__5948_,data_stage_2__5947_,data_stage_2__5946_,data_stage_2__5945_,
  data_stage_2__5944_,data_stage_2__5943_,data_stage_2__5942_,data_stage_2__5941_,
  data_stage_2__5940_,data_stage_2__5939_,data_stage_2__5938_,data_stage_2__5937_,
  data_stage_2__5936_,data_stage_2__5935_,data_stage_2__5934_,data_stage_2__5933_,
  data_stage_2__5932_,data_stage_2__5931_,data_stage_2__5930_,data_stage_2__5929_,
  data_stage_2__5928_,data_stage_2__5927_,data_stage_2__5926_,data_stage_2__5925_,
  data_stage_2__5924_,data_stage_2__5923_,data_stage_2__5922_,data_stage_2__5921_,
  data_stage_2__5920_,data_stage_2__5919_,data_stage_2__5918_,data_stage_2__5917_,
  data_stage_2__5916_,data_stage_2__5915_,data_stage_2__5914_,data_stage_2__5913_,
  data_stage_2__5912_,data_stage_2__5911_,data_stage_2__5910_,data_stage_2__5909_,
  data_stage_2__5908_,data_stage_2__5907_,data_stage_2__5906_,data_stage_2__5905_,
  data_stage_2__5904_,data_stage_2__5903_,data_stage_2__5902_,data_stage_2__5901_,
  data_stage_2__5900_,data_stage_2__5899_,data_stage_2__5898_,data_stage_2__5897_,
  data_stage_2__5896_,data_stage_2__5895_,data_stage_2__5894_,data_stage_2__5893_,
  data_stage_2__5892_,data_stage_2__5891_,data_stage_2__5890_,data_stage_2__5889_,
  data_stage_2__5888_,data_stage_2__5887_,data_stage_2__5886_,data_stage_2__5885_,
  data_stage_2__5884_,data_stage_2__5883_,data_stage_2__5882_,data_stage_2__5881_,
  data_stage_2__5880_,data_stage_2__5879_,data_stage_2__5878_,data_stage_2__5877_,
  data_stage_2__5876_,data_stage_2__5875_,data_stage_2__5874_,data_stage_2__5873_,
  data_stage_2__5872_,data_stage_2__5871_,data_stage_2__5870_,data_stage_2__5869_,
  data_stage_2__5868_,data_stage_2__5867_,data_stage_2__5866_,data_stage_2__5865_,
  data_stage_2__5864_,data_stage_2__5863_,data_stage_2__5862_,data_stage_2__5861_,
  data_stage_2__5860_,data_stage_2__5859_,data_stage_2__5858_,data_stage_2__5857_,
  data_stage_2__5856_,data_stage_2__5855_,data_stage_2__5854_,data_stage_2__5853_,
  data_stage_2__5852_,data_stage_2__5851_,data_stage_2__5850_,data_stage_2__5849_,
  data_stage_2__5848_,data_stage_2__5847_,data_stage_2__5846_,data_stage_2__5845_,
  data_stage_2__5844_,data_stage_2__5843_,data_stage_2__5842_,data_stage_2__5841_,
  data_stage_2__5840_,data_stage_2__5839_,data_stage_2__5838_,data_stage_2__5837_,
  data_stage_2__5836_,data_stage_2__5835_,data_stage_2__5834_,data_stage_2__5833_,
  data_stage_2__5832_,data_stage_2__5831_,data_stage_2__5830_,data_stage_2__5829_,
  data_stage_2__5828_,data_stage_2__5827_,data_stage_2__5826_,data_stage_2__5825_,
  data_stage_2__5824_,data_stage_2__5823_,data_stage_2__5822_,data_stage_2__5821_,
  data_stage_2__5820_,data_stage_2__5819_,data_stage_2__5818_,data_stage_2__5817_,
  data_stage_2__5816_,data_stage_2__5815_,data_stage_2__5814_,data_stage_2__5813_,
  data_stage_2__5812_,data_stage_2__5811_,data_stage_2__5810_,data_stage_2__5809_,
  data_stage_2__5808_,data_stage_2__5807_,data_stage_2__5806_,data_stage_2__5805_,
  data_stage_2__5804_,data_stage_2__5803_,data_stage_2__5802_,data_stage_2__5801_,
  data_stage_2__5800_,data_stage_2__5799_,data_stage_2__5798_,data_stage_2__5797_,
  data_stage_2__5796_,data_stage_2__5795_,data_stage_2__5794_,data_stage_2__5793_,
  data_stage_2__5792_,data_stage_2__5791_,data_stage_2__5790_,data_stage_2__5789_,
  data_stage_2__5788_,data_stage_2__5787_,data_stage_2__5786_,data_stage_2__5785_,
  data_stage_2__5784_,data_stage_2__5783_,data_stage_2__5782_,data_stage_2__5781_,
  data_stage_2__5780_,data_stage_2__5779_,data_stage_2__5778_,data_stage_2__5777_,
  data_stage_2__5776_,data_stage_2__5775_,data_stage_2__5774_,data_stage_2__5773_,
  data_stage_2__5772_,data_stage_2__5771_,data_stage_2__5770_,data_stage_2__5769_,
  data_stage_2__5768_,data_stage_2__5767_,data_stage_2__5766_,data_stage_2__5765_,
  data_stage_2__5764_,data_stage_2__5763_,data_stage_2__5762_,data_stage_2__5761_,
  data_stage_2__5760_,data_stage_2__5759_,data_stage_2__5758_,data_stage_2__5757_,
  data_stage_2__5756_,data_stage_2__5755_,data_stage_2__5754_,data_stage_2__5753_,
  data_stage_2__5752_,data_stage_2__5751_,data_stage_2__5750_,data_stage_2__5749_,
  data_stage_2__5748_,data_stage_2__5747_,data_stage_2__5746_,data_stage_2__5745_,
  data_stage_2__5744_,data_stage_2__5743_,data_stage_2__5742_,data_stage_2__5741_,
  data_stage_2__5740_,data_stage_2__5739_,data_stage_2__5738_,data_stage_2__5737_,
  data_stage_2__5736_,data_stage_2__5735_,data_stage_2__5734_,data_stage_2__5733_,
  data_stage_2__5732_,data_stage_2__5731_,data_stage_2__5730_,data_stage_2__5729_,
  data_stage_2__5728_,data_stage_2__5727_,data_stage_2__5726_,data_stage_2__5725_,
  data_stage_2__5724_,data_stage_2__5723_,data_stage_2__5722_,data_stage_2__5721_,
  data_stage_2__5720_,data_stage_2__5719_,data_stage_2__5718_,data_stage_2__5717_,
  data_stage_2__5716_,data_stage_2__5715_,data_stage_2__5714_,data_stage_2__5713_,
  data_stage_2__5712_,data_stage_2__5711_,data_stage_2__5710_,data_stage_2__5709_,
  data_stage_2__5708_,data_stage_2__5707_,data_stage_2__5706_,data_stage_2__5705_,
  data_stage_2__5704_,data_stage_2__5703_,data_stage_2__5702_,data_stage_2__5701_,
  data_stage_2__5700_,data_stage_2__5699_,data_stage_2__5698_,data_stage_2__5697_,
  data_stage_2__5696_,data_stage_2__5695_,data_stage_2__5694_,data_stage_2__5693_,
  data_stage_2__5692_,data_stage_2__5691_,data_stage_2__5690_,data_stage_2__5689_,
  data_stage_2__5688_,data_stage_2__5687_,data_stage_2__5686_,data_stage_2__5685_,
  data_stage_2__5684_,data_stage_2__5683_,data_stage_2__5682_,data_stage_2__5681_,
  data_stage_2__5680_,data_stage_2__5679_,data_stage_2__5678_,data_stage_2__5677_,
  data_stage_2__5676_,data_stage_2__5675_,data_stage_2__5674_,data_stage_2__5673_,
  data_stage_2__5672_,data_stage_2__5671_,data_stage_2__5670_,data_stage_2__5669_,
  data_stage_2__5668_,data_stage_2__5667_,data_stage_2__5666_,data_stage_2__5665_,
  data_stage_2__5664_,data_stage_2__5663_,data_stage_2__5662_,data_stage_2__5661_,
  data_stage_2__5660_,data_stage_2__5659_,data_stage_2__5658_,data_stage_2__5657_,
  data_stage_2__5656_,data_stage_2__5655_,data_stage_2__5654_,data_stage_2__5653_,
  data_stage_2__5652_,data_stage_2__5651_,data_stage_2__5650_,data_stage_2__5649_,
  data_stage_2__5648_,data_stage_2__5647_,data_stage_2__5646_,data_stage_2__5645_,
  data_stage_2__5644_,data_stage_2__5643_,data_stage_2__5642_,data_stage_2__5641_,
  data_stage_2__5640_,data_stage_2__5639_,data_stage_2__5638_,data_stage_2__5637_,
  data_stage_2__5636_,data_stage_2__5635_,data_stage_2__5634_,data_stage_2__5633_,
  data_stage_2__5632_,data_stage_2__5631_,data_stage_2__5630_,data_stage_2__5629_,
  data_stage_2__5628_,data_stage_2__5627_,data_stage_2__5626_,data_stage_2__5625_,
  data_stage_2__5624_,data_stage_2__5623_,data_stage_2__5622_,data_stage_2__5621_,
  data_stage_2__5620_,data_stage_2__5619_,data_stage_2__5618_,data_stage_2__5617_,
  data_stage_2__5616_,data_stage_2__5615_,data_stage_2__5614_,data_stage_2__5613_,
  data_stage_2__5612_,data_stage_2__5611_,data_stage_2__5610_,data_stage_2__5609_,
  data_stage_2__5608_,data_stage_2__5607_,data_stage_2__5606_,data_stage_2__5605_,
  data_stage_2__5604_,data_stage_2__5603_,data_stage_2__5602_,data_stage_2__5601_,
  data_stage_2__5600_,data_stage_2__5599_,data_stage_2__5598_,data_stage_2__5597_,
  data_stage_2__5596_,data_stage_2__5595_,data_stage_2__5594_,data_stage_2__5593_,
  data_stage_2__5592_,data_stage_2__5591_,data_stage_2__5590_,data_stage_2__5589_,
  data_stage_2__5588_,data_stage_2__5587_,data_stage_2__5586_,data_stage_2__5585_,
  data_stage_2__5584_,data_stage_2__5583_,data_stage_2__5582_,data_stage_2__5581_,
  data_stage_2__5580_,data_stage_2__5579_,data_stage_2__5578_,data_stage_2__5577_,
  data_stage_2__5576_,data_stage_2__5575_,data_stage_2__5574_,data_stage_2__5573_,
  data_stage_2__5572_,data_stage_2__5571_,data_stage_2__5570_,data_stage_2__5569_,
  data_stage_2__5568_,data_stage_2__5567_,data_stage_2__5566_,data_stage_2__5565_,
  data_stage_2__5564_,data_stage_2__5563_,data_stage_2__5562_,data_stage_2__5561_,
  data_stage_2__5560_,data_stage_2__5559_,data_stage_2__5558_,data_stage_2__5557_,
  data_stage_2__5556_,data_stage_2__5555_,data_stage_2__5554_,data_stage_2__5553_,
  data_stage_2__5552_,data_stage_2__5551_,data_stage_2__5550_,data_stage_2__5549_,
  data_stage_2__5548_,data_stage_2__5547_,data_stage_2__5546_,data_stage_2__5545_,
  data_stage_2__5544_,data_stage_2__5543_,data_stage_2__5542_,data_stage_2__5541_,
  data_stage_2__5540_,data_stage_2__5539_,data_stage_2__5538_,data_stage_2__5537_,
  data_stage_2__5536_,data_stage_2__5535_,data_stage_2__5534_,data_stage_2__5533_,
  data_stage_2__5532_,data_stage_2__5531_,data_stage_2__5530_,data_stage_2__5529_,
  data_stage_2__5528_,data_stage_2__5527_,data_stage_2__5526_,data_stage_2__5525_,
  data_stage_2__5524_,data_stage_2__5523_,data_stage_2__5522_,data_stage_2__5521_,
  data_stage_2__5520_,data_stage_2__5519_,data_stage_2__5518_,data_stage_2__5517_,
  data_stage_2__5516_,data_stage_2__5515_,data_stage_2__5514_,data_stage_2__5513_,
  data_stage_2__5512_,data_stage_2__5511_,data_stage_2__5510_,data_stage_2__5509_,
  data_stage_2__5508_,data_stage_2__5507_,data_stage_2__5506_,data_stage_2__5505_,
  data_stage_2__5504_,data_stage_2__5503_,data_stage_2__5502_,data_stage_2__5501_,
  data_stage_2__5500_,data_stage_2__5499_,data_stage_2__5498_,data_stage_2__5497_,
  data_stage_2__5496_,data_stage_2__5495_,data_stage_2__5494_,data_stage_2__5493_,
  data_stage_2__5492_,data_stage_2__5491_,data_stage_2__5490_,data_stage_2__5489_,
  data_stage_2__5488_,data_stage_2__5487_,data_stage_2__5486_,data_stage_2__5485_,
  data_stage_2__5484_,data_stage_2__5483_,data_stage_2__5482_,data_stage_2__5481_,
  data_stage_2__5480_,data_stage_2__5479_,data_stage_2__5478_,data_stage_2__5477_,
  data_stage_2__5476_,data_stage_2__5475_,data_stage_2__5474_,data_stage_2__5473_,
  data_stage_2__5472_,data_stage_2__5471_,data_stage_2__5470_,data_stage_2__5469_,
  data_stage_2__5468_,data_stage_2__5467_,data_stage_2__5466_,data_stage_2__5465_,
  data_stage_2__5464_,data_stage_2__5463_,data_stage_2__5462_,data_stage_2__5461_,
  data_stage_2__5460_,data_stage_2__5459_,data_stage_2__5458_,data_stage_2__5457_,
  data_stage_2__5456_,data_stage_2__5455_,data_stage_2__5454_,data_stage_2__5453_,
  data_stage_2__5452_,data_stage_2__5451_,data_stage_2__5450_,data_stage_2__5449_,
  data_stage_2__5448_,data_stage_2__5447_,data_stage_2__5446_,data_stage_2__5445_,
  data_stage_2__5444_,data_stage_2__5443_,data_stage_2__5442_,data_stage_2__5441_,
  data_stage_2__5440_,data_stage_2__5439_,data_stage_2__5438_,data_stage_2__5437_,
  data_stage_2__5436_,data_stage_2__5435_,data_stage_2__5434_,data_stage_2__5433_,
  data_stage_2__5432_,data_stage_2__5431_,data_stage_2__5430_,data_stage_2__5429_,
  data_stage_2__5428_,data_stage_2__5427_,data_stage_2__5426_,data_stage_2__5425_,
  data_stage_2__5424_,data_stage_2__5423_,data_stage_2__5422_,data_stage_2__5421_,
  data_stage_2__5420_,data_stage_2__5419_,data_stage_2__5418_,data_stage_2__5417_,
  data_stage_2__5416_,data_stage_2__5415_,data_stage_2__5414_,data_stage_2__5413_,
  data_stage_2__5412_,data_stage_2__5411_,data_stage_2__5410_,data_stage_2__5409_,
  data_stage_2__5408_,data_stage_2__5407_,data_stage_2__5406_,data_stage_2__5405_,
  data_stage_2__5404_,data_stage_2__5403_,data_stage_2__5402_,data_stage_2__5401_,
  data_stage_2__5400_,data_stage_2__5399_,data_stage_2__5398_,data_stage_2__5397_,
  data_stage_2__5396_,data_stage_2__5395_,data_stage_2__5394_,data_stage_2__5393_,
  data_stage_2__5392_,data_stage_2__5391_,data_stage_2__5390_,data_stage_2__5389_,
  data_stage_2__5388_,data_stage_2__5387_,data_stage_2__5386_,data_stage_2__5385_,
  data_stage_2__5384_,data_stage_2__5383_,data_stage_2__5382_,data_stage_2__5381_,
  data_stage_2__5380_,data_stage_2__5379_,data_stage_2__5378_,data_stage_2__5377_,
  data_stage_2__5376_,data_stage_2__5375_,data_stage_2__5374_,data_stage_2__5373_,
  data_stage_2__5372_,data_stage_2__5371_,data_stage_2__5370_,data_stage_2__5369_,
  data_stage_2__5368_,data_stage_2__5367_,data_stage_2__5366_,data_stage_2__5365_,
  data_stage_2__5364_,data_stage_2__5363_,data_stage_2__5362_,data_stage_2__5361_,
  data_stage_2__5360_,data_stage_2__5359_,data_stage_2__5358_,data_stage_2__5357_,
  data_stage_2__5356_,data_stage_2__5355_,data_stage_2__5354_,data_stage_2__5353_,
  data_stage_2__5352_,data_stage_2__5351_,data_stage_2__5350_,data_stage_2__5349_,
  data_stage_2__5348_,data_stage_2__5347_,data_stage_2__5346_,data_stage_2__5345_,
  data_stage_2__5344_,data_stage_2__5343_,data_stage_2__5342_,data_stage_2__5341_,
  data_stage_2__5340_,data_stage_2__5339_,data_stage_2__5338_,data_stage_2__5337_,
  data_stage_2__5336_,data_stage_2__5335_,data_stage_2__5334_,data_stage_2__5333_,
  data_stage_2__5332_,data_stage_2__5331_,data_stage_2__5330_,data_stage_2__5329_,
  data_stage_2__5328_,data_stage_2__5327_,data_stage_2__5326_,data_stage_2__5325_,
  data_stage_2__5324_,data_stage_2__5323_,data_stage_2__5322_,data_stage_2__5321_,
  data_stage_2__5320_,data_stage_2__5319_,data_stage_2__5318_,data_stage_2__5317_,
  data_stage_2__5316_,data_stage_2__5315_,data_stage_2__5314_,data_stage_2__5313_,
  data_stage_2__5312_,data_stage_2__5311_,data_stage_2__5310_,data_stage_2__5309_,
  data_stage_2__5308_,data_stage_2__5307_,data_stage_2__5306_,data_stage_2__5305_,
  data_stage_2__5304_,data_stage_2__5303_,data_stage_2__5302_,data_stage_2__5301_,
  data_stage_2__5300_,data_stage_2__5299_,data_stage_2__5298_,data_stage_2__5297_,
  data_stage_2__5296_,data_stage_2__5295_,data_stage_2__5294_,data_stage_2__5293_,
  data_stage_2__5292_,data_stage_2__5291_,data_stage_2__5290_,data_stage_2__5289_,
  data_stage_2__5288_,data_stage_2__5287_,data_stage_2__5286_,data_stage_2__5285_,
  data_stage_2__5284_,data_stage_2__5283_,data_stage_2__5282_,data_stage_2__5281_,
  data_stage_2__5280_,data_stage_2__5279_,data_stage_2__5278_,data_stage_2__5277_,
  data_stage_2__5276_,data_stage_2__5275_,data_stage_2__5274_,data_stage_2__5273_,
  data_stage_2__5272_,data_stage_2__5271_,data_stage_2__5270_,data_stage_2__5269_,
  data_stage_2__5268_,data_stage_2__5267_,data_stage_2__5266_,data_stage_2__5265_,
  data_stage_2__5264_,data_stage_2__5263_,data_stage_2__5262_,data_stage_2__5261_,
  data_stage_2__5260_,data_stage_2__5259_,data_stage_2__5258_,data_stage_2__5257_,
  data_stage_2__5256_,data_stage_2__5255_,data_stage_2__5254_,data_stage_2__5253_,
  data_stage_2__5252_,data_stage_2__5251_,data_stage_2__5250_,data_stage_2__5249_,
  data_stage_2__5248_,data_stage_2__5247_,data_stage_2__5246_,data_stage_2__5245_,
  data_stage_2__5244_,data_stage_2__5243_,data_stage_2__5242_,data_stage_2__5241_,
  data_stage_2__5240_,data_stage_2__5239_,data_stage_2__5238_,data_stage_2__5237_,
  data_stage_2__5236_,data_stage_2__5235_,data_stage_2__5234_,data_stage_2__5233_,
  data_stage_2__5232_,data_stage_2__5231_,data_stage_2__5230_,data_stage_2__5229_,
  data_stage_2__5228_,data_stage_2__5227_,data_stage_2__5226_,data_stage_2__5225_,
  data_stage_2__5224_,data_stage_2__5223_,data_stage_2__5222_,data_stage_2__5221_,
  data_stage_2__5220_,data_stage_2__5219_,data_stage_2__5218_,data_stage_2__5217_,
  data_stage_2__5216_,data_stage_2__5215_,data_stage_2__5214_,data_stage_2__5213_,
  data_stage_2__5212_,data_stage_2__5211_,data_stage_2__5210_,data_stage_2__5209_,
  data_stage_2__5208_,data_stage_2__5207_,data_stage_2__5206_,data_stage_2__5205_,
  data_stage_2__5204_,data_stage_2__5203_,data_stage_2__5202_,data_stage_2__5201_,
  data_stage_2__5200_,data_stage_2__5199_,data_stage_2__5198_,data_stage_2__5197_,
  data_stage_2__5196_,data_stage_2__5195_,data_stage_2__5194_,data_stage_2__5193_,
  data_stage_2__5192_,data_stage_2__5191_,data_stage_2__5190_,data_stage_2__5189_,
  data_stage_2__5188_,data_stage_2__5187_,data_stage_2__5186_,data_stage_2__5185_,
  data_stage_2__5184_,data_stage_2__5183_,data_stage_2__5182_,data_stage_2__5181_,
  data_stage_2__5180_,data_stage_2__5179_,data_stage_2__5178_,data_stage_2__5177_,
  data_stage_2__5176_,data_stage_2__5175_,data_stage_2__5174_,data_stage_2__5173_,
  data_stage_2__5172_,data_stage_2__5171_,data_stage_2__5170_,data_stage_2__5169_,
  data_stage_2__5168_,data_stage_2__5167_,data_stage_2__5166_,data_stage_2__5165_,
  data_stage_2__5164_,data_stage_2__5163_,data_stage_2__5162_,data_stage_2__5161_,
  data_stage_2__5160_,data_stage_2__5159_,data_stage_2__5158_,data_stage_2__5157_,
  data_stage_2__5156_,data_stage_2__5155_,data_stage_2__5154_,data_stage_2__5153_,
  data_stage_2__5152_,data_stage_2__5151_,data_stage_2__5150_,data_stage_2__5149_,
  data_stage_2__5148_,data_stage_2__5147_,data_stage_2__5146_,data_stage_2__5145_,
  data_stage_2__5144_,data_stage_2__5143_,data_stage_2__5142_,data_stage_2__5141_,
  data_stage_2__5140_,data_stage_2__5139_,data_stage_2__5138_,data_stage_2__5137_,
  data_stage_2__5136_,data_stage_2__5135_,data_stage_2__5134_,data_stage_2__5133_,
  data_stage_2__5132_,data_stage_2__5131_,data_stage_2__5130_,data_stage_2__5129_,
  data_stage_2__5128_,data_stage_2__5127_,data_stage_2__5126_,data_stage_2__5125_,
  data_stage_2__5124_,data_stage_2__5123_,data_stage_2__5122_,data_stage_2__5121_,
  data_stage_2__5120_,data_stage_2__5119_,data_stage_2__5118_,data_stage_2__5117_,
  data_stage_2__5116_,data_stage_2__5115_,data_stage_2__5114_,data_stage_2__5113_,
  data_stage_2__5112_,data_stage_2__5111_,data_stage_2__5110_,data_stage_2__5109_,
  data_stage_2__5108_,data_stage_2__5107_,data_stage_2__5106_,data_stage_2__5105_,
  data_stage_2__5104_,data_stage_2__5103_,data_stage_2__5102_,data_stage_2__5101_,
  data_stage_2__5100_,data_stage_2__5099_,data_stage_2__5098_,data_stage_2__5097_,
  data_stage_2__5096_,data_stage_2__5095_,data_stage_2__5094_,data_stage_2__5093_,
  data_stage_2__5092_,data_stage_2__5091_,data_stage_2__5090_,data_stage_2__5089_,
  data_stage_2__5088_,data_stage_2__5087_,data_stage_2__5086_,data_stage_2__5085_,
  data_stage_2__5084_,data_stage_2__5083_,data_stage_2__5082_,data_stage_2__5081_,
  data_stage_2__5080_,data_stage_2__5079_,data_stage_2__5078_,data_stage_2__5077_,
  data_stage_2__5076_,data_stage_2__5075_,data_stage_2__5074_,data_stage_2__5073_,
  data_stage_2__5072_,data_stage_2__5071_,data_stage_2__5070_,data_stage_2__5069_,
  data_stage_2__5068_,data_stage_2__5067_,data_stage_2__5066_,data_stage_2__5065_,
  data_stage_2__5064_,data_stage_2__5063_,data_stage_2__5062_,data_stage_2__5061_,
  data_stage_2__5060_,data_stage_2__5059_,data_stage_2__5058_,data_stage_2__5057_,
  data_stage_2__5056_,data_stage_2__5055_,data_stage_2__5054_,data_stage_2__5053_,
  data_stage_2__5052_,data_stage_2__5051_,data_stage_2__5050_,data_stage_2__5049_,
  data_stage_2__5048_,data_stage_2__5047_,data_stage_2__5046_,data_stage_2__5045_,
  data_stage_2__5044_,data_stage_2__5043_,data_stage_2__5042_,data_stage_2__5041_,
  data_stage_2__5040_,data_stage_2__5039_,data_stage_2__5038_,data_stage_2__5037_,
  data_stage_2__5036_,data_stage_2__5035_,data_stage_2__5034_,data_stage_2__5033_,
  data_stage_2__5032_,data_stage_2__5031_,data_stage_2__5030_,data_stage_2__5029_,
  data_stage_2__5028_,data_stage_2__5027_,data_stage_2__5026_,data_stage_2__5025_,
  data_stage_2__5024_,data_stage_2__5023_,data_stage_2__5022_,data_stage_2__5021_,
  data_stage_2__5020_,data_stage_2__5019_,data_stage_2__5018_,data_stage_2__5017_,
  data_stage_2__5016_,data_stage_2__5015_,data_stage_2__5014_,data_stage_2__5013_,
  data_stage_2__5012_,data_stage_2__5011_,data_stage_2__5010_,data_stage_2__5009_,
  data_stage_2__5008_,data_stage_2__5007_,data_stage_2__5006_,data_stage_2__5005_,
  data_stage_2__5004_,data_stage_2__5003_,data_stage_2__5002_,data_stage_2__5001_,
  data_stage_2__5000_,data_stage_2__4999_,data_stage_2__4998_,data_stage_2__4997_,
  data_stage_2__4996_,data_stage_2__4995_,data_stage_2__4994_,data_stage_2__4993_,
  data_stage_2__4992_,data_stage_2__4991_,data_stage_2__4990_,data_stage_2__4989_,
  data_stage_2__4988_,data_stage_2__4987_,data_stage_2__4986_,data_stage_2__4985_,
  data_stage_2__4984_,data_stage_2__4983_,data_stage_2__4982_,data_stage_2__4981_,
  data_stage_2__4980_,data_stage_2__4979_,data_stage_2__4978_,data_stage_2__4977_,
  data_stage_2__4976_,data_stage_2__4975_,data_stage_2__4974_,data_stage_2__4973_,
  data_stage_2__4972_,data_stage_2__4971_,data_stage_2__4970_,data_stage_2__4969_,
  data_stage_2__4968_,data_stage_2__4967_,data_stage_2__4966_,data_stage_2__4965_,
  data_stage_2__4964_,data_stage_2__4963_,data_stage_2__4962_,data_stage_2__4961_,
  data_stage_2__4960_,data_stage_2__4959_,data_stage_2__4958_,data_stage_2__4957_,
  data_stage_2__4956_,data_stage_2__4955_,data_stage_2__4954_,data_stage_2__4953_,
  data_stage_2__4952_,data_stage_2__4951_,data_stage_2__4950_,data_stage_2__4949_,
  data_stage_2__4948_,data_stage_2__4947_,data_stage_2__4946_,data_stage_2__4945_,
  data_stage_2__4944_,data_stage_2__4943_,data_stage_2__4942_,data_stage_2__4941_,
  data_stage_2__4940_,data_stage_2__4939_,data_stage_2__4938_,data_stage_2__4937_,
  data_stage_2__4936_,data_stage_2__4935_,data_stage_2__4934_,data_stage_2__4933_,
  data_stage_2__4932_,data_stage_2__4931_,data_stage_2__4930_,data_stage_2__4929_,
  data_stage_2__4928_,data_stage_2__4927_,data_stage_2__4926_,data_stage_2__4925_,
  data_stage_2__4924_,data_stage_2__4923_,data_stage_2__4922_,data_stage_2__4921_,
  data_stage_2__4920_,data_stage_2__4919_,data_stage_2__4918_,data_stage_2__4917_,
  data_stage_2__4916_,data_stage_2__4915_,data_stage_2__4914_,data_stage_2__4913_,
  data_stage_2__4912_,data_stage_2__4911_,data_stage_2__4910_,data_stage_2__4909_,
  data_stage_2__4908_,data_stage_2__4907_,data_stage_2__4906_,data_stage_2__4905_,
  data_stage_2__4904_,data_stage_2__4903_,data_stage_2__4902_,data_stage_2__4901_,
  data_stage_2__4900_,data_stage_2__4899_,data_stage_2__4898_,data_stage_2__4897_,
  data_stage_2__4896_,data_stage_2__4895_,data_stage_2__4894_,data_stage_2__4893_,
  data_stage_2__4892_,data_stage_2__4891_,data_stage_2__4890_,data_stage_2__4889_,
  data_stage_2__4888_,data_stage_2__4887_,data_stage_2__4886_,data_stage_2__4885_,
  data_stage_2__4884_,data_stage_2__4883_,data_stage_2__4882_,data_stage_2__4881_,
  data_stage_2__4880_,data_stage_2__4879_,data_stage_2__4878_,data_stage_2__4877_,
  data_stage_2__4876_,data_stage_2__4875_,data_stage_2__4874_,data_stage_2__4873_,
  data_stage_2__4872_,data_stage_2__4871_,data_stage_2__4870_,data_stage_2__4869_,
  data_stage_2__4868_,data_stage_2__4867_,data_stage_2__4866_,data_stage_2__4865_,
  data_stage_2__4864_,data_stage_2__4863_,data_stage_2__4862_,data_stage_2__4861_,
  data_stage_2__4860_,data_stage_2__4859_,data_stage_2__4858_,data_stage_2__4857_,
  data_stage_2__4856_,data_stage_2__4855_,data_stage_2__4854_,data_stage_2__4853_,
  data_stage_2__4852_,data_stage_2__4851_,data_stage_2__4850_,data_stage_2__4849_,
  data_stage_2__4848_,data_stage_2__4847_,data_stage_2__4846_,data_stage_2__4845_,
  data_stage_2__4844_,data_stage_2__4843_,data_stage_2__4842_,data_stage_2__4841_,
  data_stage_2__4840_,data_stage_2__4839_,data_stage_2__4838_,data_stage_2__4837_,
  data_stage_2__4836_,data_stage_2__4835_,data_stage_2__4834_,data_stage_2__4833_,
  data_stage_2__4832_,data_stage_2__4831_,data_stage_2__4830_,data_stage_2__4829_,
  data_stage_2__4828_,data_stage_2__4827_,data_stage_2__4826_,data_stage_2__4825_,
  data_stage_2__4824_,data_stage_2__4823_,data_stage_2__4822_,data_stage_2__4821_,
  data_stage_2__4820_,data_stage_2__4819_,data_stage_2__4818_,data_stage_2__4817_,
  data_stage_2__4816_,data_stage_2__4815_,data_stage_2__4814_,data_stage_2__4813_,
  data_stage_2__4812_,data_stage_2__4811_,data_stage_2__4810_,data_stage_2__4809_,
  data_stage_2__4808_,data_stage_2__4807_,data_stage_2__4806_,data_stage_2__4805_,
  data_stage_2__4804_,data_stage_2__4803_,data_stage_2__4802_,data_stage_2__4801_,
  data_stage_2__4800_,data_stage_2__4799_,data_stage_2__4798_,data_stage_2__4797_,
  data_stage_2__4796_,data_stage_2__4795_,data_stage_2__4794_,data_stage_2__4793_,
  data_stage_2__4792_,data_stage_2__4791_,data_stage_2__4790_,data_stage_2__4789_,
  data_stage_2__4788_,data_stage_2__4787_,data_stage_2__4786_,data_stage_2__4785_,
  data_stage_2__4784_,data_stage_2__4783_,data_stage_2__4782_,data_stage_2__4781_,
  data_stage_2__4780_,data_stage_2__4779_,data_stage_2__4778_,data_stage_2__4777_,
  data_stage_2__4776_,data_stage_2__4775_,data_stage_2__4774_,data_stage_2__4773_,
  data_stage_2__4772_,data_stage_2__4771_,data_stage_2__4770_,data_stage_2__4769_,
  data_stage_2__4768_,data_stage_2__4767_,data_stage_2__4766_,data_stage_2__4765_,
  data_stage_2__4764_,data_stage_2__4763_,data_stage_2__4762_,data_stage_2__4761_,
  data_stage_2__4760_,data_stage_2__4759_,data_stage_2__4758_,data_stage_2__4757_,
  data_stage_2__4756_,data_stage_2__4755_,data_stage_2__4754_,data_stage_2__4753_,
  data_stage_2__4752_,data_stage_2__4751_,data_stage_2__4750_,data_stage_2__4749_,
  data_stage_2__4748_,data_stage_2__4747_,data_stage_2__4746_,data_stage_2__4745_,
  data_stage_2__4744_,data_stage_2__4743_,data_stage_2__4742_,data_stage_2__4741_,
  data_stage_2__4740_,data_stage_2__4739_,data_stage_2__4738_,data_stage_2__4737_,
  data_stage_2__4736_,data_stage_2__4735_,data_stage_2__4734_,data_stage_2__4733_,
  data_stage_2__4732_,data_stage_2__4731_,data_stage_2__4730_,data_stage_2__4729_,
  data_stage_2__4728_,data_stage_2__4727_,data_stage_2__4726_,data_stage_2__4725_,
  data_stage_2__4724_,data_stage_2__4723_,data_stage_2__4722_,data_stage_2__4721_,
  data_stage_2__4720_,data_stage_2__4719_,data_stage_2__4718_,data_stage_2__4717_,
  data_stage_2__4716_,data_stage_2__4715_,data_stage_2__4714_,data_stage_2__4713_,
  data_stage_2__4712_,data_stage_2__4711_,data_stage_2__4710_,data_stage_2__4709_,
  data_stage_2__4708_,data_stage_2__4707_,data_stage_2__4706_,data_stage_2__4705_,
  data_stage_2__4704_,data_stage_2__4703_,data_stage_2__4702_,data_stage_2__4701_,
  data_stage_2__4700_,data_stage_2__4699_,data_stage_2__4698_,data_stage_2__4697_,
  data_stage_2__4696_,data_stage_2__4695_,data_stage_2__4694_,data_stage_2__4693_,
  data_stage_2__4692_,data_stage_2__4691_,data_stage_2__4690_,data_stage_2__4689_,
  data_stage_2__4688_,data_stage_2__4687_,data_stage_2__4686_,data_stage_2__4685_,
  data_stage_2__4684_,data_stage_2__4683_,data_stage_2__4682_,data_stage_2__4681_,
  data_stage_2__4680_,data_stage_2__4679_,data_stage_2__4678_,data_stage_2__4677_,
  data_stage_2__4676_,data_stage_2__4675_,data_stage_2__4674_,data_stage_2__4673_,
  data_stage_2__4672_,data_stage_2__4671_,data_stage_2__4670_,data_stage_2__4669_,
  data_stage_2__4668_,data_stage_2__4667_,data_stage_2__4666_,data_stage_2__4665_,
  data_stage_2__4664_,data_stage_2__4663_,data_stage_2__4662_,data_stage_2__4661_,
  data_stage_2__4660_,data_stage_2__4659_,data_stage_2__4658_,data_stage_2__4657_,
  data_stage_2__4656_,data_stage_2__4655_,data_stage_2__4654_,data_stage_2__4653_,
  data_stage_2__4652_,data_stage_2__4651_,data_stage_2__4650_,data_stage_2__4649_,
  data_stage_2__4648_,data_stage_2__4647_,data_stage_2__4646_,data_stage_2__4645_,
  data_stage_2__4644_,data_stage_2__4643_,data_stage_2__4642_,data_stage_2__4641_,
  data_stage_2__4640_,data_stage_2__4639_,data_stage_2__4638_,data_stage_2__4637_,
  data_stage_2__4636_,data_stage_2__4635_,data_stage_2__4634_,data_stage_2__4633_,
  data_stage_2__4632_,data_stage_2__4631_,data_stage_2__4630_,data_stage_2__4629_,
  data_stage_2__4628_,data_stage_2__4627_,data_stage_2__4626_,data_stage_2__4625_,
  data_stage_2__4624_,data_stage_2__4623_,data_stage_2__4622_,data_stage_2__4621_,
  data_stage_2__4620_,data_stage_2__4619_,data_stage_2__4618_,data_stage_2__4617_,
  data_stage_2__4616_,data_stage_2__4615_,data_stage_2__4614_,data_stage_2__4613_,
  data_stage_2__4612_,data_stage_2__4611_,data_stage_2__4610_,data_stage_2__4609_,
  data_stage_2__4608_,data_stage_2__4607_,data_stage_2__4606_,data_stage_2__4605_,
  data_stage_2__4604_,data_stage_2__4603_,data_stage_2__4602_,data_stage_2__4601_,
  data_stage_2__4600_,data_stage_2__4599_,data_stage_2__4598_,data_stage_2__4597_,
  data_stage_2__4596_,data_stage_2__4595_,data_stage_2__4594_,data_stage_2__4593_,
  data_stage_2__4592_,data_stage_2__4591_,data_stage_2__4590_,data_stage_2__4589_,
  data_stage_2__4588_,data_stage_2__4587_,data_stage_2__4586_,data_stage_2__4585_,
  data_stage_2__4584_,data_stage_2__4583_,data_stage_2__4582_,data_stage_2__4581_,
  data_stage_2__4580_,data_stage_2__4579_,data_stage_2__4578_,data_stage_2__4577_,
  data_stage_2__4576_,data_stage_2__4575_,data_stage_2__4574_,data_stage_2__4573_,
  data_stage_2__4572_,data_stage_2__4571_,data_stage_2__4570_,data_stage_2__4569_,
  data_stage_2__4568_,data_stage_2__4567_,data_stage_2__4566_,data_stage_2__4565_,
  data_stage_2__4564_,data_stage_2__4563_,data_stage_2__4562_,data_stage_2__4561_,
  data_stage_2__4560_,data_stage_2__4559_,data_stage_2__4558_,data_stage_2__4557_,
  data_stage_2__4556_,data_stage_2__4555_,data_stage_2__4554_,data_stage_2__4553_,
  data_stage_2__4552_,data_stage_2__4551_,data_stage_2__4550_,data_stage_2__4549_,
  data_stage_2__4548_,data_stage_2__4547_,data_stage_2__4546_,data_stage_2__4545_,
  data_stage_2__4544_,data_stage_2__4543_,data_stage_2__4542_,data_stage_2__4541_,
  data_stage_2__4540_,data_stage_2__4539_,data_stage_2__4538_,data_stage_2__4537_,
  data_stage_2__4536_,data_stage_2__4535_,data_stage_2__4534_,data_stage_2__4533_,
  data_stage_2__4532_,data_stage_2__4531_,data_stage_2__4530_,data_stage_2__4529_,
  data_stage_2__4528_,data_stage_2__4527_,data_stage_2__4526_,data_stage_2__4525_,
  data_stage_2__4524_,data_stage_2__4523_,data_stage_2__4522_,data_stage_2__4521_,
  data_stage_2__4520_,data_stage_2__4519_,data_stage_2__4518_,data_stage_2__4517_,
  data_stage_2__4516_,data_stage_2__4515_,data_stage_2__4514_,data_stage_2__4513_,
  data_stage_2__4512_,data_stage_2__4511_,data_stage_2__4510_,data_stage_2__4509_,
  data_stage_2__4508_,data_stage_2__4507_,data_stage_2__4506_,data_stage_2__4505_,
  data_stage_2__4504_,data_stage_2__4503_,data_stage_2__4502_,data_stage_2__4501_,
  data_stage_2__4500_,data_stage_2__4499_,data_stage_2__4498_,data_stage_2__4497_,
  data_stage_2__4496_,data_stage_2__4495_,data_stage_2__4494_,data_stage_2__4493_,
  data_stage_2__4492_,data_stage_2__4491_,data_stage_2__4490_,data_stage_2__4489_,
  data_stage_2__4488_,data_stage_2__4487_,data_stage_2__4486_,data_stage_2__4485_,
  data_stage_2__4484_,data_stage_2__4483_,data_stage_2__4482_,data_stage_2__4481_,
  data_stage_2__4480_,data_stage_2__4479_,data_stage_2__4478_,data_stage_2__4477_,
  data_stage_2__4476_,data_stage_2__4475_,data_stage_2__4474_,data_stage_2__4473_,
  data_stage_2__4472_,data_stage_2__4471_,data_stage_2__4470_,data_stage_2__4469_,
  data_stage_2__4468_,data_stage_2__4467_,data_stage_2__4466_,data_stage_2__4465_,
  data_stage_2__4464_,data_stage_2__4463_,data_stage_2__4462_,data_stage_2__4461_,
  data_stage_2__4460_,data_stage_2__4459_,data_stage_2__4458_,data_stage_2__4457_,
  data_stage_2__4456_,data_stage_2__4455_,data_stage_2__4454_,data_stage_2__4453_,
  data_stage_2__4452_,data_stage_2__4451_,data_stage_2__4450_,data_stage_2__4449_,
  data_stage_2__4448_,data_stage_2__4447_,data_stage_2__4446_,data_stage_2__4445_,
  data_stage_2__4444_,data_stage_2__4443_,data_stage_2__4442_,data_stage_2__4441_,
  data_stage_2__4440_,data_stage_2__4439_,data_stage_2__4438_,data_stage_2__4437_,
  data_stage_2__4436_,data_stage_2__4435_,data_stage_2__4434_,data_stage_2__4433_,
  data_stage_2__4432_,data_stage_2__4431_,data_stage_2__4430_,data_stage_2__4429_,
  data_stage_2__4428_,data_stage_2__4427_,data_stage_2__4426_,data_stage_2__4425_,
  data_stage_2__4424_,data_stage_2__4423_,data_stage_2__4422_,data_stage_2__4421_,
  data_stage_2__4420_,data_stage_2__4419_,data_stage_2__4418_,data_stage_2__4417_,
  data_stage_2__4416_,data_stage_2__4415_,data_stage_2__4414_,data_stage_2__4413_,
  data_stage_2__4412_,data_stage_2__4411_,data_stage_2__4410_,data_stage_2__4409_,
  data_stage_2__4408_,data_stage_2__4407_,data_stage_2__4406_,data_stage_2__4405_,
  data_stage_2__4404_,data_stage_2__4403_,data_stage_2__4402_,data_stage_2__4401_,
  data_stage_2__4400_,data_stage_2__4399_,data_stage_2__4398_,data_stage_2__4397_,
  data_stage_2__4396_,data_stage_2__4395_,data_stage_2__4394_,data_stage_2__4393_,
  data_stage_2__4392_,data_stage_2__4391_,data_stage_2__4390_,data_stage_2__4389_,
  data_stage_2__4388_,data_stage_2__4387_,data_stage_2__4386_,data_stage_2__4385_,
  data_stage_2__4384_,data_stage_2__4383_,data_stage_2__4382_,data_stage_2__4381_,
  data_stage_2__4380_,data_stage_2__4379_,data_stage_2__4378_,data_stage_2__4377_,
  data_stage_2__4376_,data_stage_2__4375_,data_stage_2__4374_,data_stage_2__4373_,
  data_stage_2__4372_,data_stage_2__4371_,data_stage_2__4370_,data_stage_2__4369_,
  data_stage_2__4368_,data_stage_2__4367_,data_stage_2__4366_,data_stage_2__4365_,
  data_stage_2__4364_,data_stage_2__4363_,data_stage_2__4362_,data_stage_2__4361_,
  data_stage_2__4360_,data_stage_2__4359_,data_stage_2__4358_,data_stage_2__4357_,
  data_stage_2__4356_,data_stage_2__4355_,data_stage_2__4354_,data_stage_2__4353_,
  data_stage_2__4352_,data_stage_2__4351_,data_stage_2__4350_,data_stage_2__4349_,
  data_stage_2__4348_,data_stage_2__4347_,data_stage_2__4346_,data_stage_2__4345_,
  data_stage_2__4344_,data_stage_2__4343_,data_stage_2__4342_,data_stage_2__4341_,
  data_stage_2__4340_,data_stage_2__4339_,data_stage_2__4338_,data_stage_2__4337_,
  data_stage_2__4336_,data_stage_2__4335_,data_stage_2__4334_,data_stage_2__4333_,
  data_stage_2__4332_,data_stage_2__4331_,data_stage_2__4330_,data_stage_2__4329_,
  data_stage_2__4328_,data_stage_2__4327_,data_stage_2__4326_,data_stage_2__4325_,
  data_stage_2__4324_,data_stage_2__4323_,data_stage_2__4322_,data_stage_2__4321_,
  data_stage_2__4320_,data_stage_2__4319_,data_stage_2__4318_,data_stage_2__4317_,
  data_stage_2__4316_,data_stage_2__4315_,data_stage_2__4314_,data_stage_2__4313_,
  data_stage_2__4312_,data_stage_2__4311_,data_stage_2__4310_,data_stage_2__4309_,
  data_stage_2__4308_,data_stage_2__4307_,data_stage_2__4306_,data_stage_2__4305_,
  data_stage_2__4304_,data_stage_2__4303_,data_stage_2__4302_,data_stage_2__4301_,
  data_stage_2__4300_,data_stage_2__4299_,data_stage_2__4298_,data_stage_2__4297_,
  data_stage_2__4296_,data_stage_2__4295_,data_stage_2__4294_,data_stage_2__4293_,
  data_stage_2__4292_,data_stage_2__4291_,data_stage_2__4290_,data_stage_2__4289_,
  data_stage_2__4288_,data_stage_2__4287_,data_stage_2__4286_,data_stage_2__4285_,
  data_stage_2__4284_,data_stage_2__4283_,data_stage_2__4282_,data_stage_2__4281_,
  data_stage_2__4280_,data_stage_2__4279_,data_stage_2__4278_,data_stage_2__4277_,
  data_stage_2__4276_,data_stage_2__4275_,data_stage_2__4274_,data_stage_2__4273_,
  data_stage_2__4272_,data_stage_2__4271_,data_stage_2__4270_,data_stage_2__4269_,
  data_stage_2__4268_,data_stage_2__4267_,data_stage_2__4266_,data_stage_2__4265_,
  data_stage_2__4264_,data_stage_2__4263_,data_stage_2__4262_,data_stage_2__4261_,
  data_stage_2__4260_,data_stage_2__4259_,data_stage_2__4258_,data_stage_2__4257_,
  data_stage_2__4256_,data_stage_2__4255_,data_stage_2__4254_,data_stage_2__4253_,
  data_stage_2__4252_,data_stage_2__4251_,data_stage_2__4250_,data_stage_2__4249_,
  data_stage_2__4248_,data_stage_2__4247_,data_stage_2__4246_,data_stage_2__4245_,
  data_stage_2__4244_,data_stage_2__4243_,data_stage_2__4242_,data_stage_2__4241_,
  data_stage_2__4240_,data_stage_2__4239_,data_stage_2__4238_,data_stage_2__4237_,
  data_stage_2__4236_,data_stage_2__4235_,data_stage_2__4234_,data_stage_2__4233_,
  data_stage_2__4232_,data_stage_2__4231_,data_stage_2__4230_,data_stage_2__4229_,
  data_stage_2__4228_,data_stage_2__4227_,data_stage_2__4226_,data_stage_2__4225_,
  data_stage_2__4224_,data_stage_2__4223_,data_stage_2__4222_,data_stage_2__4221_,
  data_stage_2__4220_,data_stage_2__4219_,data_stage_2__4218_,data_stage_2__4217_,
  data_stage_2__4216_,data_stage_2__4215_,data_stage_2__4214_,data_stage_2__4213_,
  data_stage_2__4212_,data_stage_2__4211_,data_stage_2__4210_,data_stage_2__4209_,
  data_stage_2__4208_,data_stage_2__4207_,data_stage_2__4206_,data_stage_2__4205_,
  data_stage_2__4204_,data_stage_2__4203_,data_stage_2__4202_,data_stage_2__4201_,
  data_stage_2__4200_,data_stage_2__4199_,data_stage_2__4198_,data_stage_2__4197_,
  data_stage_2__4196_,data_stage_2__4195_,data_stage_2__4194_,data_stage_2__4193_,
  data_stage_2__4192_,data_stage_2__4191_,data_stage_2__4190_,data_stage_2__4189_,
  data_stage_2__4188_,data_stage_2__4187_,data_stage_2__4186_,data_stage_2__4185_,
  data_stage_2__4184_,data_stage_2__4183_,data_stage_2__4182_,data_stage_2__4181_,
  data_stage_2__4180_,data_stage_2__4179_,data_stage_2__4178_,data_stage_2__4177_,
  data_stage_2__4176_,data_stage_2__4175_,data_stage_2__4174_,data_stage_2__4173_,
  data_stage_2__4172_,data_stage_2__4171_,data_stage_2__4170_,data_stage_2__4169_,
  data_stage_2__4168_,data_stage_2__4167_,data_stage_2__4166_,data_stage_2__4165_,
  data_stage_2__4164_,data_stage_2__4163_,data_stage_2__4162_,data_stage_2__4161_,
  data_stage_2__4160_,data_stage_2__4159_,data_stage_2__4158_,data_stage_2__4157_,
  data_stage_2__4156_,data_stage_2__4155_,data_stage_2__4154_,data_stage_2__4153_,
  data_stage_2__4152_,data_stage_2__4151_,data_stage_2__4150_,data_stage_2__4149_,
  data_stage_2__4148_,data_stage_2__4147_,data_stage_2__4146_,data_stage_2__4145_,
  data_stage_2__4144_,data_stage_2__4143_,data_stage_2__4142_,data_stage_2__4141_,
  data_stage_2__4140_,data_stage_2__4139_,data_stage_2__4138_,data_stage_2__4137_,
  data_stage_2__4136_,data_stage_2__4135_,data_stage_2__4134_,data_stage_2__4133_,
  data_stage_2__4132_,data_stage_2__4131_,data_stage_2__4130_,data_stage_2__4129_,
  data_stage_2__4128_,data_stage_2__4127_,data_stage_2__4126_,data_stage_2__4125_,
  data_stage_2__4124_,data_stage_2__4123_,data_stage_2__4122_,data_stage_2__4121_,
  data_stage_2__4120_,data_stage_2__4119_,data_stage_2__4118_,data_stage_2__4117_,
  data_stage_2__4116_,data_stage_2__4115_,data_stage_2__4114_,data_stage_2__4113_,
  data_stage_2__4112_,data_stage_2__4111_,data_stage_2__4110_,data_stage_2__4109_,
  data_stage_2__4108_,data_stage_2__4107_,data_stage_2__4106_,data_stage_2__4105_,
  data_stage_2__4104_,data_stage_2__4103_,data_stage_2__4102_,data_stage_2__4101_,
  data_stage_2__4100_,data_stage_2__4099_,data_stage_2__4098_,data_stage_2__4097_,
  data_stage_2__4096_,data_stage_2__4095_,data_stage_2__4094_,data_stage_2__4093_,
  data_stage_2__4092_,data_stage_2__4091_,data_stage_2__4090_,data_stage_2__4089_,
  data_stage_2__4088_,data_stage_2__4087_,data_stage_2__4086_,data_stage_2__4085_,
  data_stage_2__4084_,data_stage_2__4083_,data_stage_2__4082_,data_stage_2__4081_,
  data_stage_2__4080_,data_stage_2__4079_,data_stage_2__4078_,data_stage_2__4077_,
  data_stage_2__4076_,data_stage_2__4075_,data_stage_2__4074_,data_stage_2__4073_,
  data_stage_2__4072_,data_stage_2__4071_,data_stage_2__4070_,data_stage_2__4069_,
  data_stage_2__4068_,data_stage_2__4067_,data_stage_2__4066_,data_stage_2__4065_,
  data_stage_2__4064_,data_stage_2__4063_,data_stage_2__4062_,data_stage_2__4061_,
  data_stage_2__4060_,data_stage_2__4059_,data_stage_2__4058_,data_stage_2__4057_,
  data_stage_2__4056_,data_stage_2__4055_,data_stage_2__4054_,data_stage_2__4053_,
  data_stage_2__4052_,data_stage_2__4051_,data_stage_2__4050_,data_stage_2__4049_,
  data_stage_2__4048_,data_stage_2__4047_,data_stage_2__4046_,data_stage_2__4045_,
  data_stage_2__4044_,data_stage_2__4043_,data_stage_2__4042_,data_stage_2__4041_,
  data_stage_2__4040_,data_stage_2__4039_,data_stage_2__4038_,data_stage_2__4037_,
  data_stage_2__4036_,data_stage_2__4035_,data_stage_2__4034_,data_stage_2__4033_,
  data_stage_2__4032_,data_stage_2__4031_,data_stage_2__4030_,data_stage_2__4029_,
  data_stage_2__4028_,data_stage_2__4027_,data_stage_2__4026_,data_stage_2__4025_,
  data_stage_2__4024_,data_stage_2__4023_,data_stage_2__4022_,data_stage_2__4021_,
  data_stage_2__4020_,data_stage_2__4019_,data_stage_2__4018_,data_stage_2__4017_,
  data_stage_2__4016_,data_stage_2__4015_,data_stage_2__4014_,data_stage_2__4013_,
  data_stage_2__4012_,data_stage_2__4011_,data_stage_2__4010_,data_stage_2__4009_,
  data_stage_2__4008_,data_stage_2__4007_,data_stage_2__4006_,data_stage_2__4005_,
  data_stage_2__4004_,data_stage_2__4003_,data_stage_2__4002_,data_stage_2__4001_,
  data_stage_2__4000_,data_stage_2__3999_,data_stage_2__3998_,data_stage_2__3997_,
  data_stage_2__3996_,data_stage_2__3995_,data_stage_2__3994_,data_stage_2__3993_,
  data_stage_2__3992_,data_stage_2__3991_,data_stage_2__3990_,data_stage_2__3989_,
  data_stage_2__3988_,data_stage_2__3987_,data_stage_2__3986_,data_stage_2__3985_,
  data_stage_2__3984_,data_stage_2__3983_,data_stage_2__3982_,data_stage_2__3981_,
  data_stage_2__3980_,data_stage_2__3979_,data_stage_2__3978_,data_stage_2__3977_,
  data_stage_2__3976_,data_stage_2__3975_,data_stage_2__3974_,data_stage_2__3973_,
  data_stage_2__3972_,data_stage_2__3971_,data_stage_2__3970_,data_stage_2__3969_,
  data_stage_2__3968_,data_stage_2__3967_,data_stage_2__3966_,data_stage_2__3965_,
  data_stage_2__3964_,data_stage_2__3963_,data_stage_2__3962_,data_stage_2__3961_,
  data_stage_2__3960_,data_stage_2__3959_,data_stage_2__3958_,data_stage_2__3957_,
  data_stage_2__3956_,data_stage_2__3955_,data_stage_2__3954_,data_stage_2__3953_,
  data_stage_2__3952_,data_stage_2__3951_,data_stage_2__3950_,data_stage_2__3949_,
  data_stage_2__3948_,data_stage_2__3947_,data_stage_2__3946_,data_stage_2__3945_,
  data_stage_2__3944_,data_stage_2__3943_,data_stage_2__3942_,data_stage_2__3941_,
  data_stage_2__3940_,data_stage_2__3939_,data_stage_2__3938_,data_stage_2__3937_,
  data_stage_2__3936_,data_stage_2__3935_,data_stage_2__3934_,data_stage_2__3933_,
  data_stage_2__3932_,data_stage_2__3931_,data_stage_2__3930_,data_stage_2__3929_,
  data_stage_2__3928_,data_stage_2__3927_,data_stage_2__3926_,data_stage_2__3925_,
  data_stage_2__3924_,data_stage_2__3923_,data_stage_2__3922_,data_stage_2__3921_,
  data_stage_2__3920_,data_stage_2__3919_,data_stage_2__3918_,data_stage_2__3917_,
  data_stage_2__3916_,data_stage_2__3915_,data_stage_2__3914_,data_stage_2__3913_,
  data_stage_2__3912_,data_stage_2__3911_,data_stage_2__3910_,data_stage_2__3909_,
  data_stage_2__3908_,data_stage_2__3907_,data_stage_2__3906_,data_stage_2__3905_,
  data_stage_2__3904_,data_stage_2__3903_,data_stage_2__3902_,data_stage_2__3901_,
  data_stage_2__3900_,data_stage_2__3899_,data_stage_2__3898_,data_stage_2__3897_,
  data_stage_2__3896_,data_stage_2__3895_,data_stage_2__3894_,data_stage_2__3893_,
  data_stage_2__3892_,data_stage_2__3891_,data_stage_2__3890_,data_stage_2__3889_,
  data_stage_2__3888_,data_stage_2__3887_,data_stage_2__3886_,data_stage_2__3885_,
  data_stage_2__3884_,data_stage_2__3883_,data_stage_2__3882_,data_stage_2__3881_,
  data_stage_2__3880_,data_stage_2__3879_,data_stage_2__3878_,data_stage_2__3877_,
  data_stage_2__3876_,data_stage_2__3875_,data_stage_2__3874_,data_stage_2__3873_,
  data_stage_2__3872_,data_stage_2__3871_,data_stage_2__3870_,data_stage_2__3869_,
  data_stage_2__3868_,data_stage_2__3867_,data_stage_2__3866_,data_stage_2__3865_,
  data_stage_2__3864_,data_stage_2__3863_,data_stage_2__3862_,data_stage_2__3861_,
  data_stage_2__3860_,data_stage_2__3859_,data_stage_2__3858_,data_stage_2__3857_,
  data_stage_2__3856_,data_stage_2__3855_,data_stage_2__3854_,data_stage_2__3853_,
  data_stage_2__3852_,data_stage_2__3851_,data_stage_2__3850_,data_stage_2__3849_,
  data_stage_2__3848_,data_stage_2__3847_,data_stage_2__3846_,data_stage_2__3845_,
  data_stage_2__3844_,data_stage_2__3843_,data_stage_2__3842_,data_stage_2__3841_,
  data_stage_2__3840_,data_stage_2__3839_,data_stage_2__3838_,data_stage_2__3837_,
  data_stage_2__3836_,data_stage_2__3835_,data_stage_2__3834_,data_stage_2__3833_,
  data_stage_2__3832_,data_stage_2__3831_,data_stage_2__3830_,data_stage_2__3829_,
  data_stage_2__3828_,data_stage_2__3827_,data_stage_2__3826_,data_stage_2__3825_,
  data_stage_2__3824_,data_stage_2__3823_,data_stage_2__3822_,data_stage_2__3821_,
  data_stage_2__3820_,data_stage_2__3819_,data_stage_2__3818_,data_stage_2__3817_,
  data_stage_2__3816_,data_stage_2__3815_,data_stage_2__3814_,data_stage_2__3813_,
  data_stage_2__3812_,data_stage_2__3811_,data_stage_2__3810_,data_stage_2__3809_,
  data_stage_2__3808_,data_stage_2__3807_,data_stage_2__3806_,data_stage_2__3805_,
  data_stage_2__3804_,data_stage_2__3803_,data_stage_2__3802_,data_stage_2__3801_,
  data_stage_2__3800_,data_stage_2__3799_,data_stage_2__3798_,data_stage_2__3797_,
  data_stage_2__3796_,data_stage_2__3795_,data_stage_2__3794_,data_stage_2__3793_,
  data_stage_2__3792_,data_stage_2__3791_,data_stage_2__3790_,data_stage_2__3789_,
  data_stage_2__3788_,data_stage_2__3787_,data_stage_2__3786_,data_stage_2__3785_,
  data_stage_2__3784_,data_stage_2__3783_,data_stage_2__3782_,data_stage_2__3781_,
  data_stage_2__3780_,data_stage_2__3779_,data_stage_2__3778_,data_stage_2__3777_,
  data_stage_2__3776_,data_stage_2__3775_,data_stage_2__3774_,data_stage_2__3773_,
  data_stage_2__3772_,data_stage_2__3771_,data_stage_2__3770_,data_stage_2__3769_,
  data_stage_2__3768_,data_stage_2__3767_,data_stage_2__3766_,data_stage_2__3765_,
  data_stage_2__3764_,data_stage_2__3763_,data_stage_2__3762_,data_stage_2__3761_,
  data_stage_2__3760_,data_stage_2__3759_,data_stage_2__3758_,data_stage_2__3757_,
  data_stage_2__3756_,data_stage_2__3755_,data_stage_2__3754_,data_stage_2__3753_,
  data_stage_2__3752_,data_stage_2__3751_,data_stage_2__3750_,data_stage_2__3749_,
  data_stage_2__3748_,data_stage_2__3747_,data_stage_2__3746_,data_stage_2__3745_,
  data_stage_2__3744_,data_stage_2__3743_,data_stage_2__3742_,data_stage_2__3741_,
  data_stage_2__3740_,data_stage_2__3739_,data_stage_2__3738_,data_stage_2__3737_,
  data_stage_2__3736_,data_stage_2__3735_,data_stage_2__3734_,data_stage_2__3733_,
  data_stage_2__3732_,data_stage_2__3731_,data_stage_2__3730_,data_stage_2__3729_,
  data_stage_2__3728_,data_stage_2__3727_,data_stage_2__3726_,data_stage_2__3725_,
  data_stage_2__3724_,data_stage_2__3723_,data_stage_2__3722_,data_stage_2__3721_,
  data_stage_2__3720_,data_stage_2__3719_,data_stage_2__3718_,data_stage_2__3717_,
  data_stage_2__3716_,data_stage_2__3715_,data_stage_2__3714_,data_stage_2__3713_,
  data_stage_2__3712_,data_stage_2__3711_,data_stage_2__3710_,data_stage_2__3709_,
  data_stage_2__3708_,data_stage_2__3707_,data_stage_2__3706_,data_stage_2__3705_,
  data_stage_2__3704_,data_stage_2__3703_,data_stage_2__3702_,data_stage_2__3701_,
  data_stage_2__3700_,data_stage_2__3699_,data_stage_2__3698_,data_stage_2__3697_,
  data_stage_2__3696_,data_stage_2__3695_,data_stage_2__3694_,data_stage_2__3693_,
  data_stage_2__3692_,data_stage_2__3691_,data_stage_2__3690_,data_stage_2__3689_,
  data_stage_2__3688_,data_stage_2__3687_,data_stage_2__3686_,data_stage_2__3685_,
  data_stage_2__3684_,data_stage_2__3683_,data_stage_2__3682_,data_stage_2__3681_,
  data_stage_2__3680_,data_stage_2__3679_,data_stage_2__3678_,data_stage_2__3677_,
  data_stage_2__3676_,data_stage_2__3675_,data_stage_2__3674_,data_stage_2__3673_,
  data_stage_2__3672_,data_stage_2__3671_,data_stage_2__3670_,data_stage_2__3669_,
  data_stage_2__3668_,data_stage_2__3667_,data_stage_2__3666_,data_stage_2__3665_,
  data_stage_2__3664_,data_stage_2__3663_,data_stage_2__3662_,data_stage_2__3661_,
  data_stage_2__3660_,data_stage_2__3659_,data_stage_2__3658_,data_stage_2__3657_,
  data_stage_2__3656_,data_stage_2__3655_,data_stage_2__3654_,data_stage_2__3653_,
  data_stage_2__3652_,data_stage_2__3651_,data_stage_2__3650_,data_stage_2__3649_,
  data_stage_2__3648_,data_stage_2__3647_,data_stage_2__3646_,data_stage_2__3645_,
  data_stage_2__3644_,data_stage_2__3643_,data_stage_2__3642_,data_stage_2__3641_,
  data_stage_2__3640_,data_stage_2__3639_,data_stage_2__3638_,data_stage_2__3637_,
  data_stage_2__3636_,data_stage_2__3635_,data_stage_2__3634_,data_stage_2__3633_,
  data_stage_2__3632_,data_stage_2__3631_,data_stage_2__3630_,data_stage_2__3629_,
  data_stage_2__3628_,data_stage_2__3627_,data_stage_2__3626_,data_stage_2__3625_,
  data_stage_2__3624_,data_stage_2__3623_,data_stage_2__3622_,data_stage_2__3621_,
  data_stage_2__3620_,data_stage_2__3619_,data_stage_2__3618_,data_stage_2__3617_,
  data_stage_2__3616_,data_stage_2__3615_,data_stage_2__3614_,data_stage_2__3613_,
  data_stage_2__3612_,data_stage_2__3611_,data_stage_2__3610_,data_stage_2__3609_,
  data_stage_2__3608_,data_stage_2__3607_,data_stage_2__3606_,data_stage_2__3605_,
  data_stage_2__3604_,data_stage_2__3603_,data_stage_2__3602_,data_stage_2__3601_,
  data_stage_2__3600_,data_stage_2__3599_,data_stage_2__3598_,data_stage_2__3597_,
  data_stage_2__3596_,data_stage_2__3595_,data_stage_2__3594_,data_stage_2__3593_,
  data_stage_2__3592_,data_stage_2__3591_,data_stage_2__3590_,data_stage_2__3589_,
  data_stage_2__3588_,data_stage_2__3587_,data_stage_2__3586_,data_stage_2__3585_,
  data_stage_2__3584_,data_stage_2__3583_,data_stage_2__3582_,data_stage_2__3581_,
  data_stage_2__3580_,data_stage_2__3579_,data_stage_2__3578_,data_stage_2__3577_,
  data_stage_2__3576_,data_stage_2__3575_,data_stage_2__3574_,data_stage_2__3573_,
  data_stage_2__3572_,data_stage_2__3571_,data_stage_2__3570_,data_stage_2__3569_,
  data_stage_2__3568_,data_stage_2__3567_,data_stage_2__3566_,data_stage_2__3565_,
  data_stage_2__3564_,data_stage_2__3563_,data_stage_2__3562_,data_stage_2__3561_,
  data_stage_2__3560_,data_stage_2__3559_,data_stage_2__3558_,data_stage_2__3557_,
  data_stage_2__3556_,data_stage_2__3555_,data_stage_2__3554_,data_stage_2__3553_,
  data_stage_2__3552_,data_stage_2__3551_,data_stage_2__3550_,data_stage_2__3549_,
  data_stage_2__3548_,data_stage_2__3547_,data_stage_2__3546_,data_stage_2__3545_,
  data_stage_2__3544_,data_stage_2__3543_,data_stage_2__3542_,data_stage_2__3541_,
  data_stage_2__3540_,data_stage_2__3539_,data_stage_2__3538_,data_stage_2__3537_,
  data_stage_2__3536_,data_stage_2__3535_,data_stage_2__3534_,data_stage_2__3533_,
  data_stage_2__3532_,data_stage_2__3531_,data_stage_2__3530_,data_stage_2__3529_,
  data_stage_2__3528_,data_stage_2__3527_,data_stage_2__3526_,data_stage_2__3525_,
  data_stage_2__3524_,data_stage_2__3523_,data_stage_2__3522_,data_stage_2__3521_,
  data_stage_2__3520_,data_stage_2__3519_,data_stage_2__3518_,data_stage_2__3517_,
  data_stage_2__3516_,data_stage_2__3515_,data_stage_2__3514_,data_stage_2__3513_,
  data_stage_2__3512_,data_stage_2__3511_,data_stage_2__3510_,data_stage_2__3509_,
  data_stage_2__3508_,data_stage_2__3507_,data_stage_2__3506_,data_stage_2__3505_,
  data_stage_2__3504_,data_stage_2__3503_,data_stage_2__3502_,data_stage_2__3501_,
  data_stage_2__3500_,data_stage_2__3499_,data_stage_2__3498_,data_stage_2__3497_,
  data_stage_2__3496_,data_stage_2__3495_,data_stage_2__3494_,data_stage_2__3493_,
  data_stage_2__3492_,data_stage_2__3491_,data_stage_2__3490_,data_stage_2__3489_,
  data_stage_2__3488_,data_stage_2__3487_,data_stage_2__3486_,data_stage_2__3485_,
  data_stage_2__3484_,data_stage_2__3483_,data_stage_2__3482_,data_stage_2__3481_,
  data_stage_2__3480_,data_stage_2__3479_,data_stage_2__3478_,data_stage_2__3477_,
  data_stage_2__3476_,data_stage_2__3475_,data_stage_2__3474_,data_stage_2__3473_,
  data_stage_2__3472_,data_stage_2__3471_,data_stage_2__3470_,data_stage_2__3469_,
  data_stage_2__3468_,data_stage_2__3467_,data_stage_2__3466_,data_stage_2__3465_,
  data_stage_2__3464_,data_stage_2__3463_,data_stage_2__3462_,data_stage_2__3461_,
  data_stage_2__3460_,data_stage_2__3459_,data_stage_2__3458_,data_stage_2__3457_,
  data_stage_2__3456_,data_stage_2__3455_,data_stage_2__3454_,data_stage_2__3453_,
  data_stage_2__3452_,data_stage_2__3451_,data_stage_2__3450_,data_stage_2__3449_,
  data_stage_2__3448_,data_stage_2__3447_,data_stage_2__3446_,data_stage_2__3445_,
  data_stage_2__3444_,data_stage_2__3443_,data_stage_2__3442_,data_stage_2__3441_,
  data_stage_2__3440_,data_stage_2__3439_,data_stage_2__3438_,data_stage_2__3437_,
  data_stage_2__3436_,data_stage_2__3435_,data_stage_2__3434_,data_stage_2__3433_,
  data_stage_2__3432_,data_stage_2__3431_,data_stage_2__3430_,data_stage_2__3429_,
  data_stage_2__3428_,data_stage_2__3427_,data_stage_2__3426_,data_stage_2__3425_,
  data_stage_2__3424_,data_stage_2__3423_,data_stage_2__3422_,data_stage_2__3421_,
  data_stage_2__3420_,data_stage_2__3419_,data_stage_2__3418_,data_stage_2__3417_,
  data_stage_2__3416_,data_stage_2__3415_,data_stage_2__3414_,data_stage_2__3413_,
  data_stage_2__3412_,data_stage_2__3411_,data_stage_2__3410_,data_stage_2__3409_,
  data_stage_2__3408_,data_stage_2__3407_,data_stage_2__3406_,data_stage_2__3405_,
  data_stage_2__3404_,data_stage_2__3403_,data_stage_2__3402_,data_stage_2__3401_,
  data_stage_2__3400_,data_stage_2__3399_,data_stage_2__3398_,data_stage_2__3397_,
  data_stage_2__3396_,data_stage_2__3395_,data_stage_2__3394_,data_stage_2__3393_,
  data_stage_2__3392_,data_stage_2__3391_,data_stage_2__3390_,data_stage_2__3389_,
  data_stage_2__3388_,data_stage_2__3387_,data_stage_2__3386_,data_stage_2__3385_,
  data_stage_2__3384_,data_stage_2__3383_,data_stage_2__3382_,data_stage_2__3381_,
  data_stage_2__3380_,data_stage_2__3379_,data_stage_2__3378_,data_stage_2__3377_,
  data_stage_2__3376_,data_stage_2__3375_,data_stage_2__3374_,data_stage_2__3373_,
  data_stage_2__3372_,data_stage_2__3371_,data_stage_2__3370_,data_stage_2__3369_,
  data_stage_2__3368_,data_stage_2__3367_,data_stage_2__3366_,data_stage_2__3365_,
  data_stage_2__3364_,data_stage_2__3363_,data_stage_2__3362_,data_stage_2__3361_,
  data_stage_2__3360_,data_stage_2__3359_,data_stage_2__3358_,data_stage_2__3357_,
  data_stage_2__3356_,data_stage_2__3355_,data_stage_2__3354_,data_stage_2__3353_,
  data_stage_2__3352_,data_stage_2__3351_,data_stage_2__3350_,data_stage_2__3349_,
  data_stage_2__3348_,data_stage_2__3347_,data_stage_2__3346_,data_stage_2__3345_,
  data_stage_2__3344_,data_stage_2__3343_,data_stage_2__3342_,data_stage_2__3341_,
  data_stage_2__3340_,data_stage_2__3339_,data_stage_2__3338_,data_stage_2__3337_,
  data_stage_2__3336_,data_stage_2__3335_,data_stage_2__3334_,data_stage_2__3333_,
  data_stage_2__3332_,data_stage_2__3331_,data_stage_2__3330_,data_stage_2__3329_,
  data_stage_2__3328_,data_stage_2__3327_,data_stage_2__3326_,data_stage_2__3325_,
  data_stage_2__3324_,data_stage_2__3323_,data_stage_2__3322_,data_stage_2__3321_,
  data_stage_2__3320_,data_stage_2__3319_,data_stage_2__3318_,data_stage_2__3317_,
  data_stage_2__3316_,data_stage_2__3315_,data_stage_2__3314_,data_stage_2__3313_,
  data_stage_2__3312_,data_stage_2__3311_,data_stage_2__3310_,data_stage_2__3309_,
  data_stage_2__3308_,data_stage_2__3307_,data_stage_2__3306_,data_stage_2__3305_,
  data_stage_2__3304_,data_stage_2__3303_,data_stage_2__3302_,data_stage_2__3301_,
  data_stage_2__3300_,data_stage_2__3299_,data_stage_2__3298_,data_stage_2__3297_,
  data_stage_2__3296_,data_stage_2__3295_,data_stage_2__3294_,data_stage_2__3293_,
  data_stage_2__3292_,data_stage_2__3291_,data_stage_2__3290_,data_stage_2__3289_,
  data_stage_2__3288_,data_stage_2__3287_,data_stage_2__3286_,data_stage_2__3285_,
  data_stage_2__3284_,data_stage_2__3283_,data_stage_2__3282_,data_stage_2__3281_,
  data_stage_2__3280_,data_stage_2__3279_,data_stage_2__3278_,data_stage_2__3277_,
  data_stage_2__3276_,data_stage_2__3275_,data_stage_2__3274_,data_stage_2__3273_,
  data_stage_2__3272_,data_stage_2__3271_,data_stage_2__3270_,data_stage_2__3269_,
  data_stage_2__3268_,data_stage_2__3267_,data_stage_2__3266_,data_stage_2__3265_,
  data_stage_2__3264_,data_stage_2__3263_,data_stage_2__3262_,data_stage_2__3261_,
  data_stage_2__3260_,data_stage_2__3259_,data_stage_2__3258_,data_stage_2__3257_,
  data_stage_2__3256_,data_stage_2__3255_,data_stage_2__3254_,data_stage_2__3253_,
  data_stage_2__3252_,data_stage_2__3251_,data_stage_2__3250_,data_stage_2__3249_,
  data_stage_2__3248_,data_stage_2__3247_,data_stage_2__3246_,data_stage_2__3245_,
  data_stage_2__3244_,data_stage_2__3243_,data_stage_2__3242_,data_stage_2__3241_,
  data_stage_2__3240_,data_stage_2__3239_,data_stage_2__3238_,data_stage_2__3237_,
  data_stage_2__3236_,data_stage_2__3235_,data_stage_2__3234_,data_stage_2__3233_,
  data_stage_2__3232_,data_stage_2__3231_,data_stage_2__3230_,data_stage_2__3229_,
  data_stage_2__3228_,data_stage_2__3227_,data_stage_2__3226_,data_stage_2__3225_,
  data_stage_2__3224_,data_stage_2__3223_,data_stage_2__3222_,data_stage_2__3221_,
  data_stage_2__3220_,data_stage_2__3219_,data_stage_2__3218_,data_stage_2__3217_,
  data_stage_2__3216_,data_stage_2__3215_,data_stage_2__3214_,data_stage_2__3213_,
  data_stage_2__3212_,data_stage_2__3211_,data_stage_2__3210_,data_stage_2__3209_,
  data_stage_2__3208_,data_stage_2__3207_,data_stage_2__3206_,data_stage_2__3205_,
  data_stage_2__3204_,data_stage_2__3203_,data_stage_2__3202_,data_stage_2__3201_,
  data_stage_2__3200_,data_stage_2__3199_,data_stage_2__3198_,data_stage_2__3197_,
  data_stage_2__3196_,data_stage_2__3195_,data_stage_2__3194_,data_stage_2__3193_,
  data_stage_2__3192_,data_stage_2__3191_,data_stage_2__3190_,data_stage_2__3189_,
  data_stage_2__3188_,data_stage_2__3187_,data_stage_2__3186_,data_stage_2__3185_,
  data_stage_2__3184_,data_stage_2__3183_,data_stage_2__3182_,data_stage_2__3181_,
  data_stage_2__3180_,data_stage_2__3179_,data_stage_2__3178_,data_stage_2__3177_,
  data_stage_2__3176_,data_stage_2__3175_,data_stage_2__3174_,data_stage_2__3173_,
  data_stage_2__3172_,data_stage_2__3171_,data_stage_2__3170_,data_stage_2__3169_,
  data_stage_2__3168_,data_stage_2__3167_,data_stage_2__3166_,data_stage_2__3165_,
  data_stage_2__3164_,data_stage_2__3163_,data_stage_2__3162_,data_stage_2__3161_,
  data_stage_2__3160_,data_stage_2__3159_,data_stage_2__3158_,data_stage_2__3157_,
  data_stage_2__3156_,data_stage_2__3155_,data_stage_2__3154_,data_stage_2__3153_,
  data_stage_2__3152_,data_stage_2__3151_,data_stage_2__3150_,data_stage_2__3149_,
  data_stage_2__3148_,data_stage_2__3147_,data_stage_2__3146_,data_stage_2__3145_,
  data_stage_2__3144_,data_stage_2__3143_,data_stage_2__3142_,data_stage_2__3141_,
  data_stage_2__3140_,data_stage_2__3139_,data_stage_2__3138_,data_stage_2__3137_,
  data_stage_2__3136_,data_stage_2__3135_,data_stage_2__3134_,data_stage_2__3133_,
  data_stage_2__3132_,data_stage_2__3131_,data_stage_2__3130_,data_stage_2__3129_,
  data_stage_2__3128_,data_stage_2__3127_,data_stage_2__3126_,data_stage_2__3125_,
  data_stage_2__3124_,data_stage_2__3123_,data_stage_2__3122_,data_stage_2__3121_,
  data_stage_2__3120_,data_stage_2__3119_,data_stage_2__3118_,data_stage_2__3117_,
  data_stage_2__3116_,data_stage_2__3115_,data_stage_2__3114_,data_stage_2__3113_,
  data_stage_2__3112_,data_stage_2__3111_,data_stage_2__3110_,data_stage_2__3109_,
  data_stage_2__3108_,data_stage_2__3107_,data_stage_2__3106_,data_stage_2__3105_,
  data_stage_2__3104_,data_stage_2__3103_,data_stage_2__3102_,data_stage_2__3101_,
  data_stage_2__3100_,data_stage_2__3099_,data_stage_2__3098_,data_stage_2__3097_,
  data_stage_2__3096_,data_stage_2__3095_,data_stage_2__3094_,data_stage_2__3093_,
  data_stage_2__3092_,data_stage_2__3091_,data_stage_2__3090_,data_stage_2__3089_,
  data_stage_2__3088_,data_stage_2__3087_,data_stage_2__3086_,data_stage_2__3085_,
  data_stage_2__3084_,data_stage_2__3083_,data_stage_2__3082_,data_stage_2__3081_,
  data_stage_2__3080_,data_stage_2__3079_,data_stage_2__3078_,data_stage_2__3077_,
  data_stage_2__3076_,data_stage_2__3075_,data_stage_2__3074_,data_stage_2__3073_,
  data_stage_2__3072_,data_stage_2__3071_,data_stage_2__3070_,data_stage_2__3069_,
  data_stage_2__3068_,data_stage_2__3067_,data_stage_2__3066_,data_stage_2__3065_,
  data_stage_2__3064_,data_stage_2__3063_,data_stage_2__3062_,data_stage_2__3061_,
  data_stage_2__3060_,data_stage_2__3059_,data_stage_2__3058_,data_stage_2__3057_,
  data_stage_2__3056_,data_stage_2__3055_,data_stage_2__3054_,data_stage_2__3053_,
  data_stage_2__3052_,data_stage_2__3051_,data_stage_2__3050_,data_stage_2__3049_,
  data_stage_2__3048_,data_stage_2__3047_,data_stage_2__3046_,data_stage_2__3045_,
  data_stage_2__3044_,data_stage_2__3043_,data_stage_2__3042_,data_stage_2__3041_,
  data_stage_2__3040_,data_stage_2__3039_,data_stage_2__3038_,data_stage_2__3037_,
  data_stage_2__3036_,data_stage_2__3035_,data_stage_2__3034_,data_stage_2__3033_,
  data_stage_2__3032_,data_stage_2__3031_,data_stage_2__3030_,data_stage_2__3029_,
  data_stage_2__3028_,data_stage_2__3027_,data_stage_2__3026_,data_stage_2__3025_,
  data_stage_2__3024_,data_stage_2__3023_,data_stage_2__3022_,data_stage_2__3021_,
  data_stage_2__3020_,data_stage_2__3019_,data_stage_2__3018_,data_stage_2__3017_,
  data_stage_2__3016_,data_stage_2__3015_,data_stage_2__3014_,data_stage_2__3013_,
  data_stage_2__3012_,data_stage_2__3011_,data_stage_2__3010_,data_stage_2__3009_,
  data_stage_2__3008_,data_stage_2__3007_,data_stage_2__3006_,data_stage_2__3005_,
  data_stage_2__3004_,data_stage_2__3003_,data_stage_2__3002_,data_stage_2__3001_,
  data_stage_2__3000_,data_stage_2__2999_,data_stage_2__2998_,data_stage_2__2997_,
  data_stage_2__2996_,data_stage_2__2995_,data_stage_2__2994_,data_stage_2__2993_,
  data_stage_2__2992_,data_stage_2__2991_,data_stage_2__2990_,data_stage_2__2989_,
  data_stage_2__2988_,data_stage_2__2987_,data_stage_2__2986_,data_stage_2__2985_,
  data_stage_2__2984_,data_stage_2__2983_,data_stage_2__2982_,data_stage_2__2981_,
  data_stage_2__2980_,data_stage_2__2979_,data_stage_2__2978_,data_stage_2__2977_,
  data_stage_2__2976_,data_stage_2__2975_,data_stage_2__2974_,data_stage_2__2973_,
  data_stage_2__2972_,data_stage_2__2971_,data_stage_2__2970_,data_stage_2__2969_,
  data_stage_2__2968_,data_stage_2__2967_,data_stage_2__2966_,data_stage_2__2965_,
  data_stage_2__2964_,data_stage_2__2963_,data_stage_2__2962_,data_stage_2__2961_,
  data_stage_2__2960_,data_stage_2__2959_,data_stage_2__2958_,data_stage_2__2957_,
  data_stage_2__2956_,data_stage_2__2955_,data_stage_2__2954_,data_stage_2__2953_,
  data_stage_2__2952_,data_stage_2__2951_,data_stage_2__2950_,data_stage_2__2949_,
  data_stage_2__2948_,data_stage_2__2947_,data_stage_2__2946_,data_stage_2__2945_,
  data_stage_2__2944_,data_stage_2__2943_,data_stage_2__2942_,data_stage_2__2941_,
  data_stage_2__2940_,data_stage_2__2939_,data_stage_2__2938_,data_stage_2__2937_,
  data_stage_2__2936_,data_stage_2__2935_,data_stage_2__2934_,data_stage_2__2933_,
  data_stage_2__2932_,data_stage_2__2931_,data_stage_2__2930_,data_stage_2__2929_,
  data_stage_2__2928_,data_stage_2__2927_,data_stage_2__2926_,data_stage_2__2925_,
  data_stage_2__2924_,data_stage_2__2923_,data_stage_2__2922_,data_stage_2__2921_,
  data_stage_2__2920_,data_stage_2__2919_,data_stage_2__2918_,data_stage_2__2917_,
  data_stage_2__2916_,data_stage_2__2915_,data_stage_2__2914_,data_stage_2__2913_,
  data_stage_2__2912_,data_stage_2__2911_,data_stage_2__2910_,data_stage_2__2909_,
  data_stage_2__2908_,data_stage_2__2907_,data_stage_2__2906_,data_stage_2__2905_,
  data_stage_2__2904_,data_stage_2__2903_,data_stage_2__2902_,data_stage_2__2901_,
  data_stage_2__2900_,data_stage_2__2899_,data_stage_2__2898_,data_stage_2__2897_,
  data_stage_2__2896_,data_stage_2__2895_,data_stage_2__2894_,data_stage_2__2893_,
  data_stage_2__2892_,data_stage_2__2891_,data_stage_2__2890_,data_stage_2__2889_,
  data_stage_2__2888_,data_stage_2__2887_,data_stage_2__2886_,data_stage_2__2885_,
  data_stage_2__2884_,data_stage_2__2883_,data_stage_2__2882_,data_stage_2__2881_,
  data_stage_2__2880_,data_stage_2__2879_,data_stage_2__2878_,data_stage_2__2877_,
  data_stage_2__2876_,data_stage_2__2875_,data_stage_2__2874_,data_stage_2__2873_,
  data_stage_2__2872_,data_stage_2__2871_,data_stage_2__2870_,data_stage_2__2869_,
  data_stage_2__2868_,data_stage_2__2867_,data_stage_2__2866_,data_stage_2__2865_,
  data_stage_2__2864_,data_stage_2__2863_,data_stage_2__2862_,data_stage_2__2861_,
  data_stage_2__2860_,data_stage_2__2859_,data_stage_2__2858_,data_stage_2__2857_,
  data_stage_2__2856_,data_stage_2__2855_,data_stage_2__2854_,data_stage_2__2853_,
  data_stage_2__2852_,data_stage_2__2851_,data_stage_2__2850_,data_stage_2__2849_,
  data_stage_2__2848_,data_stage_2__2847_,data_stage_2__2846_,data_stage_2__2845_,
  data_stage_2__2844_,data_stage_2__2843_,data_stage_2__2842_,data_stage_2__2841_,
  data_stage_2__2840_,data_stage_2__2839_,data_stage_2__2838_,data_stage_2__2837_,
  data_stage_2__2836_,data_stage_2__2835_,data_stage_2__2834_,data_stage_2__2833_,
  data_stage_2__2832_,data_stage_2__2831_,data_stage_2__2830_,data_stage_2__2829_,
  data_stage_2__2828_,data_stage_2__2827_,data_stage_2__2826_,data_stage_2__2825_,
  data_stage_2__2824_,data_stage_2__2823_,data_stage_2__2822_,data_stage_2__2821_,
  data_stage_2__2820_,data_stage_2__2819_,data_stage_2__2818_,data_stage_2__2817_,
  data_stage_2__2816_,data_stage_2__2815_,data_stage_2__2814_,data_stage_2__2813_,
  data_stage_2__2812_,data_stage_2__2811_,data_stage_2__2810_,data_stage_2__2809_,
  data_stage_2__2808_,data_stage_2__2807_,data_stage_2__2806_,data_stage_2__2805_,
  data_stage_2__2804_,data_stage_2__2803_,data_stage_2__2802_,data_stage_2__2801_,
  data_stage_2__2800_,data_stage_2__2799_,data_stage_2__2798_,data_stage_2__2797_,
  data_stage_2__2796_,data_stage_2__2795_,data_stage_2__2794_,data_stage_2__2793_,
  data_stage_2__2792_,data_stage_2__2791_,data_stage_2__2790_,data_stage_2__2789_,
  data_stage_2__2788_,data_stage_2__2787_,data_stage_2__2786_,data_stage_2__2785_,
  data_stage_2__2784_,data_stage_2__2783_,data_stage_2__2782_,data_stage_2__2781_,
  data_stage_2__2780_,data_stage_2__2779_,data_stage_2__2778_,data_stage_2__2777_,
  data_stage_2__2776_,data_stage_2__2775_,data_stage_2__2774_,data_stage_2__2773_,
  data_stage_2__2772_,data_stage_2__2771_,data_stage_2__2770_,data_stage_2__2769_,
  data_stage_2__2768_,data_stage_2__2767_,data_stage_2__2766_,data_stage_2__2765_,
  data_stage_2__2764_,data_stage_2__2763_,data_stage_2__2762_,data_stage_2__2761_,
  data_stage_2__2760_,data_stage_2__2759_,data_stage_2__2758_,data_stage_2__2757_,
  data_stage_2__2756_,data_stage_2__2755_,data_stage_2__2754_,data_stage_2__2753_,
  data_stage_2__2752_,data_stage_2__2751_,data_stage_2__2750_,data_stage_2__2749_,
  data_stage_2__2748_,data_stage_2__2747_,data_stage_2__2746_,data_stage_2__2745_,
  data_stage_2__2744_,data_stage_2__2743_,data_stage_2__2742_,data_stage_2__2741_,
  data_stage_2__2740_,data_stage_2__2739_,data_stage_2__2738_,data_stage_2__2737_,
  data_stage_2__2736_,data_stage_2__2735_,data_stage_2__2734_,data_stage_2__2733_,
  data_stage_2__2732_,data_stage_2__2731_,data_stage_2__2730_,data_stage_2__2729_,
  data_stage_2__2728_,data_stage_2__2727_,data_stage_2__2726_,data_stage_2__2725_,
  data_stage_2__2724_,data_stage_2__2723_,data_stage_2__2722_,data_stage_2__2721_,
  data_stage_2__2720_,data_stage_2__2719_,data_stage_2__2718_,data_stage_2__2717_,
  data_stage_2__2716_,data_stage_2__2715_,data_stage_2__2714_,data_stage_2__2713_,
  data_stage_2__2712_,data_stage_2__2711_,data_stage_2__2710_,data_stage_2__2709_,
  data_stage_2__2708_,data_stage_2__2707_,data_stage_2__2706_,data_stage_2__2705_,
  data_stage_2__2704_,data_stage_2__2703_,data_stage_2__2702_,data_stage_2__2701_,
  data_stage_2__2700_,data_stage_2__2699_,data_stage_2__2698_,data_stage_2__2697_,
  data_stage_2__2696_,data_stage_2__2695_,data_stage_2__2694_,data_stage_2__2693_,
  data_stage_2__2692_,data_stage_2__2691_,data_stage_2__2690_,data_stage_2__2689_,
  data_stage_2__2688_,data_stage_2__2687_,data_stage_2__2686_,data_stage_2__2685_,
  data_stage_2__2684_,data_stage_2__2683_,data_stage_2__2682_,data_stage_2__2681_,
  data_stage_2__2680_,data_stage_2__2679_,data_stage_2__2678_,data_stage_2__2677_,
  data_stage_2__2676_,data_stage_2__2675_,data_stage_2__2674_,data_stage_2__2673_,
  data_stage_2__2672_,data_stage_2__2671_,data_stage_2__2670_,data_stage_2__2669_,
  data_stage_2__2668_,data_stage_2__2667_,data_stage_2__2666_,data_stage_2__2665_,
  data_stage_2__2664_,data_stage_2__2663_,data_stage_2__2662_,data_stage_2__2661_,
  data_stage_2__2660_,data_stage_2__2659_,data_stage_2__2658_,data_stage_2__2657_,
  data_stage_2__2656_,data_stage_2__2655_,data_stage_2__2654_,data_stage_2__2653_,
  data_stage_2__2652_,data_stage_2__2651_,data_stage_2__2650_,data_stage_2__2649_,
  data_stage_2__2648_,data_stage_2__2647_,data_stage_2__2646_,data_stage_2__2645_,
  data_stage_2__2644_,data_stage_2__2643_,data_stage_2__2642_,data_stage_2__2641_,
  data_stage_2__2640_,data_stage_2__2639_,data_stage_2__2638_,data_stage_2__2637_,
  data_stage_2__2636_,data_stage_2__2635_,data_stage_2__2634_,data_stage_2__2633_,
  data_stage_2__2632_,data_stage_2__2631_,data_stage_2__2630_,data_stage_2__2629_,
  data_stage_2__2628_,data_stage_2__2627_,data_stage_2__2626_,data_stage_2__2625_,
  data_stage_2__2624_,data_stage_2__2623_,data_stage_2__2622_,data_stage_2__2621_,
  data_stage_2__2620_,data_stage_2__2619_,data_stage_2__2618_,data_stage_2__2617_,
  data_stage_2__2616_,data_stage_2__2615_,data_stage_2__2614_,data_stage_2__2613_,
  data_stage_2__2612_,data_stage_2__2611_,data_stage_2__2610_,data_stage_2__2609_,
  data_stage_2__2608_,data_stage_2__2607_,data_stage_2__2606_,data_stage_2__2605_,
  data_stage_2__2604_,data_stage_2__2603_,data_stage_2__2602_,data_stage_2__2601_,
  data_stage_2__2600_,data_stage_2__2599_,data_stage_2__2598_,data_stage_2__2597_,
  data_stage_2__2596_,data_stage_2__2595_,data_stage_2__2594_,data_stage_2__2593_,
  data_stage_2__2592_,data_stage_2__2591_,data_stage_2__2590_,data_stage_2__2589_,
  data_stage_2__2588_,data_stage_2__2587_,data_stage_2__2586_,data_stage_2__2585_,
  data_stage_2__2584_,data_stage_2__2583_,data_stage_2__2582_,data_stage_2__2581_,
  data_stage_2__2580_,data_stage_2__2579_,data_stage_2__2578_,data_stage_2__2577_,
  data_stage_2__2576_,data_stage_2__2575_,data_stage_2__2574_,data_stage_2__2573_,
  data_stage_2__2572_,data_stage_2__2571_,data_stage_2__2570_,data_stage_2__2569_,
  data_stage_2__2568_,data_stage_2__2567_,data_stage_2__2566_,data_stage_2__2565_,
  data_stage_2__2564_,data_stage_2__2563_,data_stage_2__2562_,data_stage_2__2561_,
  data_stage_2__2560_,data_stage_2__2559_,data_stage_2__2558_,data_stage_2__2557_,
  data_stage_2__2556_,data_stage_2__2555_,data_stage_2__2554_,data_stage_2__2553_,
  data_stage_2__2552_,data_stage_2__2551_,data_stage_2__2550_,data_stage_2__2549_,
  data_stage_2__2548_,data_stage_2__2547_,data_stage_2__2546_,data_stage_2__2545_,
  data_stage_2__2544_,data_stage_2__2543_,data_stage_2__2542_,data_stage_2__2541_,
  data_stage_2__2540_,data_stage_2__2539_,data_stage_2__2538_,data_stage_2__2537_,
  data_stage_2__2536_,data_stage_2__2535_,data_stage_2__2534_,data_stage_2__2533_,
  data_stage_2__2532_,data_stage_2__2531_,data_stage_2__2530_,data_stage_2__2529_,
  data_stage_2__2528_,data_stage_2__2527_,data_stage_2__2526_,data_stage_2__2525_,
  data_stage_2__2524_,data_stage_2__2523_,data_stage_2__2522_,data_stage_2__2521_,
  data_stage_2__2520_,data_stage_2__2519_,data_stage_2__2518_,data_stage_2__2517_,
  data_stage_2__2516_,data_stage_2__2515_,data_stage_2__2514_,data_stage_2__2513_,
  data_stage_2__2512_,data_stage_2__2511_,data_stage_2__2510_,data_stage_2__2509_,
  data_stage_2__2508_,data_stage_2__2507_,data_stage_2__2506_,data_stage_2__2505_,
  data_stage_2__2504_,data_stage_2__2503_,data_stage_2__2502_,data_stage_2__2501_,
  data_stage_2__2500_,data_stage_2__2499_,data_stage_2__2498_,data_stage_2__2497_,
  data_stage_2__2496_,data_stage_2__2495_,data_stage_2__2494_,data_stage_2__2493_,
  data_stage_2__2492_,data_stage_2__2491_,data_stage_2__2490_,data_stage_2__2489_,
  data_stage_2__2488_,data_stage_2__2487_,data_stage_2__2486_,data_stage_2__2485_,
  data_stage_2__2484_,data_stage_2__2483_,data_stage_2__2482_,data_stage_2__2481_,
  data_stage_2__2480_,data_stage_2__2479_,data_stage_2__2478_,data_stage_2__2477_,
  data_stage_2__2476_,data_stage_2__2475_,data_stage_2__2474_,data_stage_2__2473_,
  data_stage_2__2472_,data_stage_2__2471_,data_stage_2__2470_,data_stage_2__2469_,
  data_stage_2__2468_,data_stage_2__2467_,data_stage_2__2466_,data_stage_2__2465_,
  data_stage_2__2464_,data_stage_2__2463_,data_stage_2__2462_,data_stage_2__2461_,
  data_stage_2__2460_,data_stage_2__2459_,data_stage_2__2458_,data_stage_2__2457_,
  data_stage_2__2456_,data_stage_2__2455_,data_stage_2__2454_,data_stage_2__2453_,
  data_stage_2__2452_,data_stage_2__2451_,data_stage_2__2450_,data_stage_2__2449_,
  data_stage_2__2448_,data_stage_2__2447_,data_stage_2__2446_,data_stage_2__2445_,
  data_stage_2__2444_,data_stage_2__2443_,data_stage_2__2442_,data_stage_2__2441_,
  data_stage_2__2440_,data_stage_2__2439_,data_stage_2__2438_,data_stage_2__2437_,
  data_stage_2__2436_,data_stage_2__2435_,data_stage_2__2434_,data_stage_2__2433_,
  data_stage_2__2432_,data_stage_2__2431_,data_stage_2__2430_,data_stage_2__2429_,
  data_stage_2__2428_,data_stage_2__2427_,data_stage_2__2426_,data_stage_2__2425_,
  data_stage_2__2424_,data_stage_2__2423_,data_stage_2__2422_,data_stage_2__2421_,
  data_stage_2__2420_,data_stage_2__2419_,data_stage_2__2418_,data_stage_2__2417_,
  data_stage_2__2416_,data_stage_2__2415_,data_stage_2__2414_,data_stage_2__2413_,
  data_stage_2__2412_,data_stage_2__2411_,data_stage_2__2410_,data_stage_2__2409_,
  data_stage_2__2408_,data_stage_2__2407_,data_stage_2__2406_,data_stage_2__2405_,
  data_stage_2__2404_,data_stage_2__2403_,data_stage_2__2402_,data_stage_2__2401_,
  data_stage_2__2400_,data_stage_2__2399_,data_stage_2__2398_,data_stage_2__2397_,
  data_stage_2__2396_,data_stage_2__2395_,data_stage_2__2394_,data_stage_2__2393_,
  data_stage_2__2392_,data_stage_2__2391_,data_stage_2__2390_,data_stage_2__2389_,
  data_stage_2__2388_,data_stage_2__2387_,data_stage_2__2386_,data_stage_2__2385_,
  data_stage_2__2384_,data_stage_2__2383_,data_stage_2__2382_,data_stage_2__2381_,
  data_stage_2__2380_,data_stage_2__2379_,data_stage_2__2378_,data_stage_2__2377_,
  data_stage_2__2376_,data_stage_2__2375_,data_stage_2__2374_,data_stage_2__2373_,
  data_stage_2__2372_,data_stage_2__2371_,data_stage_2__2370_,data_stage_2__2369_,
  data_stage_2__2368_,data_stage_2__2367_,data_stage_2__2366_,data_stage_2__2365_,
  data_stage_2__2364_,data_stage_2__2363_,data_stage_2__2362_,data_stage_2__2361_,
  data_stage_2__2360_,data_stage_2__2359_,data_stage_2__2358_,data_stage_2__2357_,
  data_stage_2__2356_,data_stage_2__2355_,data_stage_2__2354_,data_stage_2__2353_,
  data_stage_2__2352_,data_stage_2__2351_,data_stage_2__2350_,data_stage_2__2349_,
  data_stage_2__2348_,data_stage_2__2347_,data_stage_2__2346_,data_stage_2__2345_,
  data_stage_2__2344_,data_stage_2__2343_,data_stage_2__2342_,data_stage_2__2341_,
  data_stage_2__2340_,data_stage_2__2339_,data_stage_2__2338_,data_stage_2__2337_,
  data_stage_2__2336_,data_stage_2__2335_,data_stage_2__2334_,data_stage_2__2333_,
  data_stage_2__2332_,data_stage_2__2331_,data_stage_2__2330_,data_stage_2__2329_,
  data_stage_2__2328_,data_stage_2__2327_,data_stage_2__2326_,data_stage_2__2325_,
  data_stage_2__2324_,data_stage_2__2323_,data_stage_2__2322_,data_stage_2__2321_,
  data_stage_2__2320_,data_stage_2__2319_,data_stage_2__2318_,data_stage_2__2317_,
  data_stage_2__2316_,data_stage_2__2315_,data_stage_2__2314_,data_stage_2__2313_,
  data_stage_2__2312_,data_stage_2__2311_,data_stage_2__2310_,data_stage_2__2309_,
  data_stage_2__2308_,data_stage_2__2307_,data_stage_2__2306_,data_stage_2__2305_,
  data_stage_2__2304_,data_stage_2__2303_,data_stage_2__2302_,data_stage_2__2301_,
  data_stage_2__2300_,data_stage_2__2299_,data_stage_2__2298_,data_stage_2__2297_,
  data_stage_2__2296_,data_stage_2__2295_,data_stage_2__2294_,data_stage_2__2293_,
  data_stage_2__2292_,data_stage_2__2291_,data_stage_2__2290_,data_stage_2__2289_,
  data_stage_2__2288_,data_stage_2__2287_,data_stage_2__2286_,data_stage_2__2285_,
  data_stage_2__2284_,data_stage_2__2283_,data_stage_2__2282_,data_stage_2__2281_,
  data_stage_2__2280_,data_stage_2__2279_,data_stage_2__2278_,data_stage_2__2277_,
  data_stage_2__2276_,data_stage_2__2275_,data_stage_2__2274_,data_stage_2__2273_,
  data_stage_2__2272_,data_stage_2__2271_,data_stage_2__2270_,data_stage_2__2269_,
  data_stage_2__2268_,data_stage_2__2267_,data_stage_2__2266_,data_stage_2__2265_,
  data_stage_2__2264_,data_stage_2__2263_,data_stage_2__2262_,data_stage_2__2261_,
  data_stage_2__2260_,data_stage_2__2259_,data_stage_2__2258_,data_stage_2__2257_,
  data_stage_2__2256_,data_stage_2__2255_,data_stage_2__2254_,data_stage_2__2253_,
  data_stage_2__2252_,data_stage_2__2251_,data_stage_2__2250_,data_stage_2__2249_,
  data_stage_2__2248_,data_stage_2__2247_,data_stage_2__2246_,data_stage_2__2245_,
  data_stage_2__2244_,data_stage_2__2243_,data_stage_2__2242_,data_stage_2__2241_,
  data_stage_2__2240_,data_stage_2__2239_,data_stage_2__2238_,data_stage_2__2237_,
  data_stage_2__2236_,data_stage_2__2235_,data_stage_2__2234_,data_stage_2__2233_,
  data_stage_2__2232_,data_stage_2__2231_,data_stage_2__2230_,data_stage_2__2229_,
  data_stage_2__2228_,data_stage_2__2227_,data_stage_2__2226_,data_stage_2__2225_,
  data_stage_2__2224_,data_stage_2__2223_,data_stage_2__2222_,data_stage_2__2221_,
  data_stage_2__2220_,data_stage_2__2219_,data_stage_2__2218_,data_stage_2__2217_,
  data_stage_2__2216_,data_stage_2__2215_,data_stage_2__2214_,data_stage_2__2213_,
  data_stage_2__2212_,data_stage_2__2211_,data_stage_2__2210_,data_stage_2__2209_,
  data_stage_2__2208_,data_stage_2__2207_,data_stage_2__2206_,data_stage_2__2205_,
  data_stage_2__2204_,data_stage_2__2203_,data_stage_2__2202_,data_stage_2__2201_,
  data_stage_2__2200_,data_stage_2__2199_,data_stage_2__2198_,data_stage_2__2197_,
  data_stage_2__2196_,data_stage_2__2195_,data_stage_2__2194_,data_stage_2__2193_,
  data_stage_2__2192_,data_stage_2__2191_,data_stage_2__2190_,data_stage_2__2189_,
  data_stage_2__2188_,data_stage_2__2187_,data_stage_2__2186_,data_stage_2__2185_,
  data_stage_2__2184_,data_stage_2__2183_,data_stage_2__2182_,data_stage_2__2181_,
  data_stage_2__2180_,data_stage_2__2179_,data_stage_2__2178_,data_stage_2__2177_,
  data_stage_2__2176_,data_stage_2__2175_,data_stage_2__2174_,data_stage_2__2173_,
  data_stage_2__2172_,data_stage_2__2171_,data_stage_2__2170_,data_stage_2__2169_,
  data_stage_2__2168_,data_stage_2__2167_,data_stage_2__2166_,data_stage_2__2165_,
  data_stage_2__2164_,data_stage_2__2163_,data_stage_2__2162_,data_stage_2__2161_,
  data_stage_2__2160_,data_stage_2__2159_,data_stage_2__2158_,data_stage_2__2157_,
  data_stage_2__2156_,data_stage_2__2155_,data_stage_2__2154_,data_stage_2__2153_,
  data_stage_2__2152_,data_stage_2__2151_,data_stage_2__2150_,data_stage_2__2149_,
  data_stage_2__2148_,data_stage_2__2147_,data_stage_2__2146_,data_stage_2__2145_,
  data_stage_2__2144_,data_stage_2__2143_,data_stage_2__2142_,data_stage_2__2141_,
  data_stage_2__2140_,data_stage_2__2139_,data_stage_2__2138_,data_stage_2__2137_,
  data_stage_2__2136_,data_stage_2__2135_,data_stage_2__2134_,data_stage_2__2133_,
  data_stage_2__2132_,data_stage_2__2131_,data_stage_2__2130_,data_stage_2__2129_,
  data_stage_2__2128_,data_stage_2__2127_,data_stage_2__2126_,data_stage_2__2125_,
  data_stage_2__2124_,data_stage_2__2123_,data_stage_2__2122_,data_stage_2__2121_,
  data_stage_2__2120_,data_stage_2__2119_,data_stage_2__2118_,data_stage_2__2117_,
  data_stage_2__2116_,data_stage_2__2115_,data_stage_2__2114_,data_stage_2__2113_,
  data_stage_2__2112_,data_stage_2__2111_,data_stage_2__2110_,data_stage_2__2109_,
  data_stage_2__2108_,data_stage_2__2107_,data_stage_2__2106_,data_stage_2__2105_,
  data_stage_2__2104_,data_stage_2__2103_,data_stage_2__2102_,data_stage_2__2101_,
  data_stage_2__2100_,data_stage_2__2099_,data_stage_2__2098_,data_stage_2__2097_,
  data_stage_2__2096_,data_stage_2__2095_,data_stage_2__2094_,data_stage_2__2093_,
  data_stage_2__2092_,data_stage_2__2091_,data_stage_2__2090_,data_stage_2__2089_,
  data_stage_2__2088_,data_stage_2__2087_,data_stage_2__2086_,data_stage_2__2085_,
  data_stage_2__2084_,data_stage_2__2083_,data_stage_2__2082_,data_stage_2__2081_,
  data_stage_2__2080_,data_stage_2__2079_,data_stage_2__2078_,data_stage_2__2077_,
  data_stage_2__2076_,data_stage_2__2075_,data_stage_2__2074_,data_stage_2__2073_,
  data_stage_2__2072_,data_stage_2__2071_,data_stage_2__2070_,data_stage_2__2069_,
  data_stage_2__2068_,data_stage_2__2067_,data_stage_2__2066_,data_stage_2__2065_,
  data_stage_2__2064_,data_stage_2__2063_,data_stage_2__2062_,data_stage_2__2061_,
  data_stage_2__2060_,data_stage_2__2059_,data_stage_2__2058_,data_stage_2__2057_,
  data_stage_2__2056_,data_stage_2__2055_,data_stage_2__2054_,data_stage_2__2053_,
  data_stage_2__2052_,data_stage_2__2051_,data_stage_2__2050_,data_stage_2__2049_,
  data_stage_2__2048_,data_stage_2__2047_,data_stage_2__2046_,data_stage_2__2045_,
  data_stage_2__2044_,data_stage_2__2043_,data_stage_2__2042_,data_stage_2__2041_,
  data_stage_2__2040_,data_stage_2__2039_,data_stage_2__2038_,data_stage_2__2037_,
  data_stage_2__2036_,data_stage_2__2035_,data_stage_2__2034_,data_stage_2__2033_,
  data_stage_2__2032_,data_stage_2__2031_,data_stage_2__2030_,data_stage_2__2029_,
  data_stage_2__2028_,data_stage_2__2027_,data_stage_2__2026_,data_stage_2__2025_,
  data_stage_2__2024_,data_stage_2__2023_,data_stage_2__2022_,data_stage_2__2021_,
  data_stage_2__2020_,data_stage_2__2019_,data_stage_2__2018_,data_stage_2__2017_,
  data_stage_2__2016_,data_stage_2__2015_,data_stage_2__2014_,data_stage_2__2013_,
  data_stage_2__2012_,data_stage_2__2011_,data_stage_2__2010_,data_stage_2__2009_,
  data_stage_2__2008_,data_stage_2__2007_,data_stage_2__2006_,data_stage_2__2005_,
  data_stage_2__2004_,data_stage_2__2003_,data_stage_2__2002_,data_stage_2__2001_,
  data_stage_2__2000_,data_stage_2__1999_,data_stage_2__1998_,data_stage_2__1997_,
  data_stage_2__1996_,data_stage_2__1995_,data_stage_2__1994_,data_stage_2__1993_,
  data_stage_2__1992_,data_stage_2__1991_,data_stage_2__1990_,data_stage_2__1989_,
  data_stage_2__1988_,data_stage_2__1987_,data_stage_2__1986_,data_stage_2__1985_,
  data_stage_2__1984_,data_stage_2__1983_,data_stage_2__1982_,data_stage_2__1981_,
  data_stage_2__1980_,data_stage_2__1979_,data_stage_2__1978_,data_stage_2__1977_,
  data_stage_2__1976_,data_stage_2__1975_,data_stage_2__1974_,data_stage_2__1973_,
  data_stage_2__1972_,data_stage_2__1971_,data_stage_2__1970_,data_stage_2__1969_,
  data_stage_2__1968_,data_stage_2__1967_,data_stage_2__1966_,data_stage_2__1965_,
  data_stage_2__1964_,data_stage_2__1963_,data_stage_2__1962_,data_stage_2__1961_,
  data_stage_2__1960_,data_stage_2__1959_,data_stage_2__1958_,data_stage_2__1957_,
  data_stage_2__1956_,data_stage_2__1955_,data_stage_2__1954_,data_stage_2__1953_,
  data_stage_2__1952_,data_stage_2__1951_,data_stage_2__1950_,data_stage_2__1949_,
  data_stage_2__1948_,data_stage_2__1947_,data_stage_2__1946_,data_stage_2__1945_,
  data_stage_2__1944_,data_stage_2__1943_,data_stage_2__1942_,data_stage_2__1941_,
  data_stage_2__1940_,data_stage_2__1939_,data_stage_2__1938_,data_stage_2__1937_,
  data_stage_2__1936_,data_stage_2__1935_,data_stage_2__1934_,data_stage_2__1933_,
  data_stage_2__1932_,data_stage_2__1931_,data_stage_2__1930_,data_stage_2__1929_,
  data_stage_2__1928_,data_stage_2__1927_,data_stage_2__1926_,data_stage_2__1925_,
  data_stage_2__1924_,data_stage_2__1923_,data_stage_2__1922_,data_stage_2__1921_,
  data_stage_2__1920_,data_stage_2__1919_,data_stage_2__1918_,data_stage_2__1917_,
  data_stage_2__1916_,data_stage_2__1915_,data_stage_2__1914_,data_stage_2__1913_,
  data_stage_2__1912_,data_stage_2__1911_,data_stage_2__1910_,data_stage_2__1909_,
  data_stage_2__1908_,data_stage_2__1907_,data_stage_2__1906_,data_stage_2__1905_,
  data_stage_2__1904_,data_stage_2__1903_,data_stage_2__1902_,data_stage_2__1901_,
  data_stage_2__1900_,data_stage_2__1899_,data_stage_2__1898_,data_stage_2__1897_,
  data_stage_2__1896_,data_stage_2__1895_,data_stage_2__1894_,data_stage_2__1893_,
  data_stage_2__1892_,data_stage_2__1891_,data_stage_2__1890_,data_stage_2__1889_,
  data_stage_2__1888_,data_stage_2__1887_,data_stage_2__1886_,data_stage_2__1885_,
  data_stage_2__1884_,data_stage_2__1883_,data_stage_2__1882_,data_stage_2__1881_,
  data_stage_2__1880_,data_stage_2__1879_,data_stage_2__1878_,data_stage_2__1877_,
  data_stage_2__1876_,data_stage_2__1875_,data_stage_2__1874_,data_stage_2__1873_,
  data_stage_2__1872_,data_stage_2__1871_,data_stage_2__1870_,data_stage_2__1869_,
  data_stage_2__1868_,data_stage_2__1867_,data_stage_2__1866_,data_stage_2__1865_,
  data_stage_2__1864_,data_stage_2__1863_,data_stage_2__1862_,data_stage_2__1861_,
  data_stage_2__1860_,data_stage_2__1859_,data_stage_2__1858_,data_stage_2__1857_,
  data_stage_2__1856_,data_stage_2__1855_,data_stage_2__1854_,data_stage_2__1853_,
  data_stage_2__1852_,data_stage_2__1851_,data_stage_2__1850_,data_stage_2__1849_,
  data_stage_2__1848_,data_stage_2__1847_,data_stage_2__1846_,data_stage_2__1845_,
  data_stage_2__1844_,data_stage_2__1843_,data_stage_2__1842_,data_stage_2__1841_,
  data_stage_2__1840_,data_stage_2__1839_,data_stage_2__1838_,data_stage_2__1837_,
  data_stage_2__1836_,data_stage_2__1835_,data_stage_2__1834_,data_stage_2__1833_,
  data_stage_2__1832_,data_stage_2__1831_,data_stage_2__1830_,data_stage_2__1829_,
  data_stage_2__1828_,data_stage_2__1827_,data_stage_2__1826_,data_stage_2__1825_,
  data_stage_2__1824_,data_stage_2__1823_,data_stage_2__1822_,data_stage_2__1821_,
  data_stage_2__1820_,data_stage_2__1819_,data_stage_2__1818_,data_stage_2__1817_,
  data_stage_2__1816_,data_stage_2__1815_,data_stage_2__1814_,data_stage_2__1813_,
  data_stage_2__1812_,data_stage_2__1811_,data_stage_2__1810_,data_stage_2__1809_,
  data_stage_2__1808_,data_stage_2__1807_,data_stage_2__1806_,data_stage_2__1805_,
  data_stage_2__1804_,data_stage_2__1803_,data_stage_2__1802_,data_stage_2__1801_,
  data_stage_2__1800_,data_stage_2__1799_,data_stage_2__1798_,data_stage_2__1797_,
  data_stage_2__1796_,data_stage_2__1795_,data_stage_2__1794_,data_stage_2__1793_,
  data_stage_2__1792_,data_stage_2__1791_,data_stage_2__1790_,data_stage_2__1789_,
  data_stage_2__1788_,data_stage_2__1787_,data_stage_2__1786_,data_stage_2__1785_,
  data_stage_2__1784_,data_stage_2__1783_,data_stage_2__1782_,data_stage_2__1781_,
  data_stage_2__1780_,data_stage_2__1779_,data_stage_2__1778_,data_stage_2__1777_,
  data_stage_2__1776_,data_stage_2__1775_,data_stage_2__1774_,data_stage_2__1773_,
  data_stage_2__1772_,data_stage_2__1771_,data_stage_2__1770_,data_stage_2__1769_,
  data_stage_2__1768_,data_stage_2__1767_,data_stage_2__1766_,data_stage_2__1765_,
  data_stage_2__1764_,data_stage_2__1763_,data_stage_2__1762_,data_stage_2__1761_,
  data_stage_2__1760_,data_stage_2__1759_,data_stage_2__1758_,data_stage_2__1757_,
  data_stage_2__1756_,data_stage_2__1755_,data_stage_2__1754_,data_stage_2__1753_,
  data_stage_2__1752_,data_stage_2__1751_,data_stage_2__1750_,data_stage_2__1749_,
  data_stage_2__1748_,data_stage_2__1747_,data_stage_2__1746_,data_stage_2__1745_,
  data_stage_2__1744_,data_stage_2__1743_,data_stage_2__1742_,data_stage_2__1741_,
  data_stage_2__1740_,data_stage_2__1739_,data_stage_2__1738_,data_stage_2__1737_,
  data_stage_2__1736_,data_stage_2__1735_,data_stage_2__1734_,data_stage_2__1733_,
  data_stage_2__1732_,data_stage_2__1731_,data_stage_2__1730_,data_stage_2__1729_,
  data_stage_2__1728_,data_stage_2__1727_,data_stage_2__1726_,data_stage_2__1725_,
  data_stage_2__1724_,data_stage_2__1723_,data_stage_2__1722_,data_stage_2__1721_,
  data_stage_2__1720_,data_stage_2__1719_,data_stage_2__1718_,data_stage_2__1717_,
  data_stage_2__1716_,data_stage_2__1715_,data_stage_2__1714_,data_stage_2__1713_,
  data_stage_2__1712_,data_stage_2__1711_,data_stage_2__1710_,data_stage_2__1709_,
  data_stage_2__1708_,data_stage_2__1707_,data_stage_2__1706_,data_stage_2__1705_,
  data_stage_2__1704_,data_stage_2__1703_,data_stage_2__1702_,data_stage_2__1701_,
  data_stage_2__1700_,data_stage_2__1699_,data_stage_2__1698_,data_stage_2__1697_,
  data_stage_2__1696_,data_stage_2__1695_,data_stage_2__1694_,data_stage_2__1693_,
  data_stage_2__1692_,data_stage_2__1691_,data_stage_2__1690_,data_stage_2__1689_,
  data_stage_2__1688_,data_stage_2__1687_,data_stage_2__1686_,data_stage_2__1685_,
  data_stage_2__1684_,data_stage_2__1683_,data_stage_2__1682_,data_stage_2__1681_,
  data_stage_2__1680_,data_stage_2__1679_,data_stage_2__1678_,data_stage_2__1677_,
  data_stage_2__1676_,data_stage_2__1675_,data_stage_2__1674_,data_stage_2__1673_,
  data_stage_2__1672_,data_stage_2__1671_,data_stage_2__1670_,data_stage_2__1669_,
  data_stage_2__1668_,data_stage_2__1667_,data_stage_2__1666_,data_stage_2__1665_,
  data_stage_2__1664_,data_stage_2__1663_,data_stage_2__1662_,data_stage_2__1661_,
  data_stage_2__1660_,data_stage_2__1659_,data_stage_2__1658_,data_stage_2__1657_,
  data_stage_2__1656_,data_stage_2__1655_,data_stage_2__1654_,data_stage_2__1653_,
  data_stage_2__1652_,data_stage_2__1651_,data_stage_2__1650_,data_stage_2__1649_,
  data_stage_2__1648_,data_stage_2__1647_,data_stage_2__1646_,data_stage_2__1645_,
  data_stage_2__1644_,data_stage_2__1643_,data_stage_2__1642_,data_stage_2__1641_,
  data_stage_2__1640_,data_stage_2__1639_,data_stage_2__1638_,data_stage_2__1637_,
  data_stage_2__1636_,data_stage_2__1635_,data_stage_2__1634_,data_stage_2__1633_,
  data_stage_2__1632_,data_stage_2__1631_,data_stage_2__1630_,data_stage_2__1629_,
  data_stage_2__1628_,data_stage_2__1627_,data_stage_2__1626_,data_stage_2__1625_,
  data_stage_2__1624_,data_stage_2__1623_,data_stage_2__1622_,data_stage_2__1621_,
  data_stage_2__1620_,data_stage_2__1619_,data_stage_2__1618_,data_stage_2__1617_,
  data_stage_2__1616_,data_stage_2__1615_,data_stage_2__1614_,data_stage_2__1613_,
  data_stage_2__1612_,data_stage_2__1611_,data_stage_2__1610_,data_stage_2__1609_,
  data_stage_2__1608_,data_stage_2__1607_,data_stage_2__1606_,data_stage_2__1605_,
  data_stage_2__1604_,data_stage_2__1603_,data_stage_2__1602_,data_stage_2__1601_,
  data_stage_2__1600_,data_stage_2__1599_,data_stage_2__1598_,data_stage_2__1597_,
  data_stage_2__1596_,data_stage_2__1595_,data_stage_2__1594_,data_stage_2__1593_,
  data_stage_2__1592_,data_stage_2__1591_,data_stage_2__1590_,data_stage_2__1589_,
  data_stage_2__1588_,data_stage_2__1587_,data_stage_2__1586_,data_stage_2__1585_,
  data_stage_2__1584_,data_stage_2__1583_,data_stage_2__1582_,data_stage_2__1581_,
  data_stage_2__1580_,data_stage_2__1579_,data_stage_2__1578_,data_stage_2__1577_,
  data_stage_2__1576_,data_stage_2__1575_,data_stage_2__1574_,data_stage_2__1573_,
  data_stage_2__1572_,data_stage_2__1571_,data_stage_2__1570_,data_stage_2__1569_,
  data_stage_2__1568_,data_stage_2__1567_,data_stage_2__1566_,data_stage_2__1565_,
  data_stage_2__1564_,data_stage_2__1563_,data_stage_2__1562_,data_stage_2__1561_,
  data_stage_2__1560_,data_stage_2__1559_,data_stage_2__1558_,data_stage_2__1557_,
  data_stage_2__1556_,data_stage_2__1555_,data_stage_2__1554_,data_stage_2__1553_,
  data_stage_2__1552_,data_stage_2__1551_,data_stage_2__1550_,data_stage_2__1549_,
  data_stage_2__1548_,data_stage_2__1547_,data_stage_2__1546_,data_stage_2__1545_,
  data_stage_2__1544_,data_stage_2__1543_,data_stage_2__1542_,data_stage_2__1541_,
  data_stage_2__1540_,data_stage_2__1539_,data_stage_2__1538_,data_stage_2__1537_,
  data_stage_2__1536_,data_stage_2__1535_,data_stage_2__1534_,data_stage_2__1533_,
  data_stage_2__1532_,data_stage_2__1531_,data_stage_2__1530_,data_stage_2__1529_,
  data_stage_2__1528_,data_stage_2__1527_,data_stage_2__1526_,data_stage_2__1525_,
  data_stage_2__1524_,data_stage_2__1523_,data_stage_2__1522_,data_stage_2__1521_,
  data_stage_2__1520_,data_stage_2__1519_,data_stage_2__1518_,data_stage_2__1517_,
  data_stage_2__1516_,data_stage_2__1515_,data_stage_2__1514_,data_stage_2__1513_,
  data_stage_2__1512_,data_stage_2__1511_,data_stage_2__1510_,data_stage_2__1509_,
  data_stage_2__1508_,data_stage_2__1507_,data_stage_2__1506_,data_stage_2__1505_,
  data_stage_2__1504_,data_stage_2__1503_,data_stage_2__1502_,data_stage_2__1501_,
  data_stage_2__1500_,data_stage_2__1499_,data_stage_2__1498_,data_stage_2__1497_,
  data_stage_2__1496_,data_stage_2__1495_,data_stage_2__1494_,data_stage_2__1493_,
  data_stage_2__1492_,data_stage_2__1491_,data_stage_2__1490_,data_stage_2__1489_,
  data_stage_2__1488_,data_stage_2__1487_,data_stage_2__1486_,data_stage_2__1485_,
  data_stage_2__1484_,data_stage_2__1483_,data_stage_2__1482_,data_stage_2__1481_,
  data_stage_2__1480_,data_stage_2__1479_,data_stage_2__1478_,data_stage_2__1477_,
  data_stage_2__1476_,data_stage_2__1475_,data_stage_2__1474_,data_stage_2__1473_,
  data_stage_2__1472_,data_stage_2__1471_,data_stage_2__1470_,data_stage_2__1469_,
  data_stage_2__1468_,data_stage_2__1467_,data_stage_2__1466_,data_stage_2__1465_,
  data_stage_2__1464_,data_stage_2__1463_,data_stage_2__1462_,data_stage_2__1461_,
  data_stage_2__1460_,data_stage_2__1459_,data_stage_2__1458_,data_stage_2__1457_,
  data_stage_2__1456_,data_stage_2__1455_,data_stage_2__1454_,data_stage_2__1453_,
  data_stage_2__1452_,data_stage_2__1451_,data_stage_2__1450_,data_stage_2__1449_,
  data_stage_2__1448_,data_stage_2__1447_,data_stage_2__1446_,data_stage_2__1445_,
  data_stage_2__1444_,data_stage_2__1443_,data_stage_2__1442_,data_stage_2__1441_,
  data_stage_2__1440_,data_stage_2__1439_,data_stage_2__1438_,data_stage_2__1437_,
  data_stage_2__1436_,data_stage_2__1435_,data_stage_2__1434_,data_stage_2__1433_,
  data_stage_2__1432_,data_stage_2__1431_,data_stage_2__1430_,data_stage_2__1429_,
  data_stage_2__1428_,data_stage_2__1427_,data_stage_2__1426_,data_stage_2__1425_,
  data_stage_2__1424_,data_stage_2__1423_,data_stage_2__1422_,data_stage_2__1421_,
  data_stage_2__1420_,data_stage_2__1419_,data_stage_2__1418_,data_stage_2__1417_,
  data_stage_2__1416_,data_stage_2__1415_,data_stage_2__1414_,data_stage_2__1413_,
  data_stage_2__1412_,data_stage_2__1411_,data_stage_2__1410_,data_stage_2__1409_,
  data_stage_2__1408_,data_stage_2__1407_,data_stage_2__1406_,data_stage_2__1405_,
  data_stage_2__1404_,data_stage_2__1403_,data_stage_2__1402_,data_stage_2__1401_,
  data_stage_2__1400_,data_stage_2__1399_,data_stage_2__1398_,data_stage_2__1397_,
  data_stage_2__1396_,data_stage_2__1395_,data_stage_2__1394_,data_stage_2__1393_,
  data_stage_2__1392_,data_stage_2__1391_,data_stage_2__1390_,data_stage_2__1389_,
  data_stage_2__1388_,data_stage_2__1387_,data_stage_2__1386_,data_stage_2__1385_,
  data_stage_2__1384_,data_stage_2__1383_,data_stage_2__1382_,data_stage_2__1381_,
  data_stage_2__1380_,data_stage_2__1379_,data_stage_2__1378_,data_stage_2__1377_,
  data_stage_2__1376_,data_stage_2__1375_,data_stage_2__1374_,data_stage_2__1373_,
  data_stage_2__1372_,data_stage_2__1371_,data_stage_2__1370_,data_stage_2__1369_,
  data_stage_2__1368_,data_stage_2__1367_,data_stage_2__1366_,data_stage_2__1365_,
  data_stage_2__1364_,data_stage_2__1363_,data_stage_2__1362_,data_stage_2__1361_,
  data_stage_2__1360_,data_stage_2__1359_,data_stage_2__1358_,data_stage_2__1357_,
  data_stage_2__1356_,data_stage_2__1355_,data_stage_2__1354_,data_stage_2__1353_,
  data_stage_2__1352_,data_stage_2__1351_,data_stage_2__1350_,data_stage_2__1349_,
  data_stage_2__1348_,data_stage_2__1347_,data_stage_2__1346_,data_stage_2__1345_,
  data_stage_2__1344_,data_stage_2__1343_,data_stage_2__1342_,data_stage_2__1341_,
  data_stage_2__1340_,data_stage_2__1339_,data_stage_2__1338_,data_stage_2__1337_,
  data_stage_2__1336_,data_stage_2__1335_,data_stage_2__1334_,data_stage_2__1333_,
  data_stage_2__1332_,data_stage_2__1331_,data_stage_2__1330_,data_stage_2__1329_,
  data_stage_2__1328_,data_stage_2__1327_,data_stage_2__1326_,data_stage_2__1325_,
  data_stage_2__1324_,data_stage_2__1323_,data_stage_2__1322_,data_stage_2__1321_,
  data_stage_2__1320_,data_stage_2__1319_,data_stage_2__1318_,data_stage_2__1317_,
  data_stage_2__1316_,data_stage_2__1315_,data_stage_2__1314_,data_stage_2__1313_,
  data_stage_2__1312_,data_stage_2__1311_,data_stage_2__1310_,data_stage_2__1309_,
  data_stage_2__1308_,data_stage_2__1307_,data_stage_2__1306_,data_stage_2__1305_,
  data_stage_2__1304_,data_stage_2__1303_,data_stage_2__1302_,data_stage_2__1301_,
  data_stage_2__1300_,data_stage_2__1299_,data_stage_2__1298_,data_stage_2__1297_,
  data_stage_2__1296_,data_stage_2__1295_,data_stage_2__1294_,data_stage_2__1293_,
  data_stage_2__1292_,data_stage_2__1291_,data_stage_2__1290_,data_stage_2__1289_,
  data_stage_2__1288_,data_stage_2__1287_,data_stage_2__1286_,data_stage_2__1285_,
  data_stage_2__1284_,data_stage_2__1283_,data_stage_2__1282_,data_stage_2__1281_,
  data_stage_2__1280_,data_stage_2__1279_,data_stage_2__1278_,data_stage_2__1277_,
  data_stage_2__1276_,data_stage_2__1275_,data_stage_2__1274_,data_stage_2__1273_,
  data_stage_2__1272_,data_stage_2__1271_,data_stage_2__1270_,data_stage_2__1269_,
  data_stage_2__1268_,data_stage_2__1267_,data_stage_2__1266_,data_stage_2__1265_,
  data_stage_2__1264_,data_stage_2__1263_,data_stage_2__1262_,data_stage_2__1261_,
  data_stage_2__1260_,data_stage_2__1259_,data_stage_2__1258_,data_stage_2__1257_,
  data_stage_2__1256_,data_stage_2__1255_,data_stage_2__1254_,data_stage_2__1253_,
  data_stage_2__1252_,data_stage_2__1251_,data_stage_2__1250_,data_stage_2__1249_,
  data_stage_2__1248_,data_stage_2__1247_,data_stage_2__1246_,data_stage_2__1245_,
  data_stage_2__1244_,data_stage_2__1243_,data_stage_2__1242_,data_stage_2__1241_,
  data_stage_2__1240_,data_stage_2__1239_,data_stage_2__1238_,data_stage_2__1237_,
  data_stage_2__1236_,data_stage_2__1235_,data_stage_2__1234_,data_stage_2__1233_,
  data_stage_2__1232_,data_stage_2__1231_,data_stage_2__1230_,data_stage_2__1229_,
  data_stage_2__1228_,data_stage_2__1227_,data_stage_2__1226_,data_stage_2__1225_,
  data_stage_2__1224_,data_stage_2__1223_,data_stage_2__1222_,data_stage_2__1221_,
  data_stage_2__1220_,data_stage_2__1219_,data_stage_2__1218_,data_stage_2__1217_,
  data_stage_2__1216_,data_stage_2__1215_,data_stage_2__1214_,data_stage_2__1213_,
  data_stage_2__1212_,data_stage_2__1211_,data_stage_2__1210_,data_stage_2__1209_,
  data_stage_2__1208_,data_stage_2__1207_,data_stage_2__1206_,data_stage_2__1205_,
  data_stage_2__1204_,data_stage_2__1203_,data_stage_2__1202_,data_stage_2__1201_,
  data_stage_2__1200_,data_stage_2__1199_,data_stage_2__1198_,data_stage_2__1197_,
  data_stage_2__1196_,data_stage_2__1195_,data_stage_2__1194_,data_stage_2__1193_,
  data_stage_2__1192_,data_stage_2__1191_,data_stage_2__1190_,data_stage_2__1189_,
  data_stage_2__1188_,data_stage_2__1187_,data_stage_2__1186_,data_stage_2__1185_,
  data_stage_2__1184_,data_stage_2__1183_,data_stage_2__1182_,data_stage_2__1181_,
  data_stage_2__1180_,data_stage_2__1179_,data_stage_2__1178_,data_stage_2__1177_,
  data_stage_2__1176_,data_stage_2__1175_,data_stage_2__1174_,data_stage_2__1173_,
  data_stage_2__1172_,data_stage_2__1171_,data_stage_2__1170_,data_stage_2__1169_,
  data_stage_2__1168_,data_stage_2__1167_,data_stage_2__1166_,data_stage_2__1165_,
  data_stage_2__1164_,data_stage_2__1163_,data_stage_2__1162_,data_stage_2__1161_,
  data_stage_2__1160_,data_stage_2__1159_,data_stage_2__1158_,data_stage_2__1157_,
  data_stage_2__1156_,data_stage_2__1155_,data_stage_2__1154_,data_stage_2__1153_,
  data_stage_2__1152_,data_stage_2__1151_,data_stage_2__1150_,data_stage_2__1149_,
  data_stage_2__1148_,data_stage_2__1147_,data_stage_2__1146_,data_stage_2__1145_,
  data_stage_2__1144_,data_stage_2__1143_,data_stage_2__1142_,data_stage_2__1141_,
  data_stage_2__1140_,data_stage_2__1139_,data_stage_2__1138_,data_stage_2__1137_,
  data_stage_2__1136_,data_stage_2__1135_,data_stage_2__1134_,data_stage_2__1133_,
  data_stage_2__1132_,data_stage_2__1131_,data_stage_2__1130_,data_stage_2__1129_,
  data_stage_2__1128_,data_stage_2__1127_,data_stage_2__1126_,data_stage_2__1125_,
  data_stage_2__1124_,data_stage_2__1123_,data_stage_2__1122_,data_stage_2__1121_,
  data_stage_2__1120_,data_stage_2__1119_,data_stage_2__1118_,data_stage_2__1117_,
  data_stage_2__1116_,data_stage_2__1115_,data_stage_2__1114_,data_stage_2__1113_,
  data_stage_2__1112_,data_stage_2__1111_,data_stage_2__1110_,data_stage_2__1109_,
  data_stage_2__1108_,data_stage_2__1107_,data_stage_2__1106_,data_stage_2__1105_,
  data_stage_2__1104_,data_stage_2__1103_,data_stage_2__1102_,data_stage_2__1101_,
  data_stage_2__1100_,data_stage_2__1099_,data_stage_2__1098_,data_stage_2__1097_,
  data_stage_2__1096_,data_stage_2__1095_,data_stage_2__1094_,data_stage_2__1093_,
  data_stage_2__1092_,data_stage_2__1091_,data_stage_2__1090_,data_stage_2__1089_,
  data_stage_2__1088_,data_stage_2__1087_,data_stage_2__1086_,data_stage_2__1085_,
  data_stage_2__1084_,data_stage_2__1083_,data_stage_2__1082_,data_stage_2__1081_,
  data_stage_2__1080_,data_stage_2__1079_,data_stage_2__1078_,data_stage_2__1077_,
  data_stage_2__1076_,data_stage_2__1075_,data_stage_2__1074_,data_stage_2__1073_,
  data_stage_2__1072_,data_stage_2__1071_,data_stage_2__1070_,data_stage_2__1069_,
  data_stage_2__1068_,data_stage_2__1067_,data_stage_2__1066_,data_stage_2__1065_,
  data_stage_2__1064_,data_stage_2__1063_,data_stage_2__1062_,data_stage_2__1061_,
  data_stage_2__1060_,data_stage_2__1059_,data_stage_2__1058_,data_stage_2__1057_,
  data_stage_2__1056_,data_stage_2__1055_,data_stage_2__1054_,data_stage_2__1053_,
  data_stage_2__1052_,data_stage_2__1051_,data_stage_2__1050_,data_stage_2__1049_,
  data_stage_2__1048_,data_stage_2__1047_,data_stage_2__1046_,data_stage_2__1045_,
  data_stage_2__1044_,data_stage_2__1043_,data_stage_2__1042_,data_stage_2__1041_,
  data_stage_2__1040_,data_stage_2__1039_,data_stage_2__1038_,data_stage_2__1037_,
  data_stage_2__1036_,data_stage_2__1035_,data_stage_2__1034_,data_stage_2__1033_,
  data_stage_2__1032_,data_stage_2__1031_,data_stage_2__1030_,data_stage_2__1029_,
  data_stage_2__1028_,data_stage_2__1027_,data_stage_2__1026_,data_stage_2__1025_,
  data_stage_2__1024_,data_stage_2__1023_,data_stage_2__1022_,data_stage_2__1021_,
  data_stage_2__1020_,data_stage_2__1019_,data_stage_2__1018_,data_stage_2__1017_,
  data_stage_2__1016_,data_stage_2__1015_,data_stage_2__1014_,data_stage_2__1013_,
  data_stage_2__1012_,data_stage_2__1011_,data_stage_2__1010_,data_stage_2__1009_,
  data_stage_2__1008_,data_stage_2__1007_,data_stage_2__1006_,data_stage_2__1005_,
  data_stage_2__1004_,data_stage_2__1003_,data_stage_2__1002_,data_stage_2__1001_,
  data_stage_2__1000_,data_stage_2__999_,data_stage_2__998_,data_stage_2__997_,
  data_stage_2__996_,data_stage_2__995_,data_stage_2__994_,data_stage_2__993_,
  data_stage_2__992_,data_stage_2__991_,data_stage_2__990_,data_stage_2__989_,data_stage_2__988_,
  data_stage_2__987_,data_stage_2__986_,data_stage_2__985_,data_stage_2__984_,
  data_stage_2__983_,data_stage_2__982_,data_stage_2__981_,data_stage_2__980_,
  data_stage_2__979_,data_stage_2__978_,data_stage_2__977_,data_stage_2__976_,
  data_stage_2__975_,data_stage_2__974_,data_stage_2__973_,data_stage_2__972_,
  data_stage_2__971_,data_stage_2__970_,data_stage_2__969_,data_stage_2__968_,data_stage_2__967_,
  data_stage_2__966_,data_stage_2__965_,data_stage_2__964_,data_stage_2__963_,
  data_stage_2__962_,data_stage_2__961_,data_stage_2__960_,data_stage_2__959_,
  data_stage_2__958_,data_stage_2__957_,data_stage_2__956_,data_stage_2__955_,
  data_stage_2__954_,data_stage_2__953_,data_stage_2__952_,data_stage_2__951_,data_stage_2__950_,
  data_stage_2__949_,data_stage_2__948_,data_stage_2__947_,data_stage_2__946_,
  data_stage_2__945_,data_stage_2__944_,data_stage_2__943_,data_stage_2__942_,
  data_stage_2__941_,data_stage_2__940_,data_stage_2__939_,data_stage_2__938_,
  data_stage_2__937_,data_stage_2__936_,data_stage_2__935_,data_stage_2__934_,
  data_stage_2__933_,data_stage_2__932_,data_stage_2__931_,data_stage_2__930_,data_stage_2__929_,
  data_stage_2__928_,data_stage_2__927_,data_stage_2__926_,data_stage_2__925_,
  data_stage_2__924_,data_stage_2__923_,data_stage_2__922_,data_stage_2__921_,
  data_stage_2__920_,data_stage_2__919_,data_stage_2__918_,data_stage_2__917_,
  data_stage_2__916_,data_stage_2__915_,data_stage_2__914_,data_stage_2__913_,
  data_stage_2__912_,data_stage_2__911_,data_stage_2__910_,data_stage_2__909_,data_stage_2__908_,
  data_stage_2__907_,data_stage_2__906_,data_stage_2__905_,data_stage_2__904_,
  data_stage_2__903_,data_stage_2__902_,data_stage_2__901_,data_stage_2__900_,
  data_stage_2__899_,data_stage_2__898_,data_stage_2__897_,data_stage_2__896_,
  data_stage_2__895_,data_stage_2__894_,data_stage_2__893_,data_stage_2__892_,
  data_stage_2__891_,data_stage_2__890_,data_stage_2__889_,data_stage_2__888_,data_stage_2__887_,
  data_stage_2__886_,data_stage_2__885_,data_stage_2__884_,data_stage_2__883_,
  data_stage_2__882_,data_stage_2__881_,data_stage_2__880_,data_stage_2__879_,
  data_stage_2__878_,data_stage_2__877_,data_stage_2__876_,data_stage_2__875_,
  data_stage_2__874_,data_stage_2__873_,data_stage_2__872_,data_stage_2__871_,data_stage_2__870_,
  data_stage_2__869_,data_stage_2__868_,data_stage_2__867_,data_stage_2__866_,
  data_stage_2__865_,data_stage_2__864_,data_stage_2__863_,data_stage_2__862_,
  data_stage_2__861_,data_stage_2__860_,data_stage_2__859_,data_stage_2__858_,
  data_stage_2__857_,data_stage_2__856_,data_stage_2__855_,data_stage_2__854_,
  data_stage_2__853_,data_stage_2__852_,data_stage_2__851_,data_stage_2__850_,data_stage_2__849_,
  data_stage_2__848_,data_stage_2__847_,data_stage_2__846_,data_stage_2__845_,
  data_stage_2__844_,data_stage_2__843_,data_stage_2__842_,data_stage_2__841_,
  data_stage_2__840_,data_stage_2__839_,data_stage_2__838_,data_stage_2__837_,
  data_stage_2__836_,data_stage_2__835_,data_stage_2__834_,data_stage_2__833_,
  data_stage_2__832_,data_stage_2__831_,data_stage_2__830_,data_stage_2__829_,data_stage_2__828_,
  data_stage_2__827_,data_stage_2__826_,data_stage_2__825_,data_stage_2__824_,
  data_stage_2__823_,data_stage_2__822_,data_stage_2__821_,data_stage_2__820_,
  data_stage_2__819_,data_stage_2__818_,data_stage_2__817_,data_stage_2__816_,
  data_stage_2__815_,data_stage_2__814_,data_stage_2__813_,data_stage_2__812_,
  data_stage_2__811_,data_stage_2__810_,data_stage_2__809_,data_stage_2__808_,data_stage_2__807_,
  data_stage_2__806_,data_stage_2__805_,data_stage_2__804_,data_stage_2__803_,
  data_stage_2__802_,data_stage_2__801_,data_stage_2__800_,data_stage_2__799_,
  data_stage_2__798_,data_stage_2__797_,data_stage_2__796_,data_stage_2__795_,
  data_stage_2__794_,data_stage_2__793_,data_stage_2__792_,data_stage_2__791_,data_stage_2__790_,
  data_stage_2__789_,data_stage_2__788_,data_stage_2__787_,data_stage_2__786_,
  data_stage_2__785_,data_stage_2__784_,data_stage_2__783_,data_stage_2__782_,
  data_stage_2__781_,data_stage_2__780_,data_stage_2__779_,data_stage_2__778_,
  data_stage_2__777_,data_stage_2__776_,data_stage_2__775_,data_stage_2__774_,
  data_stage_2__773_,data_stage_2__772_,data_stage_2__771_,data_stage_2__770_,data_stage_2__769_,
  data_stage_2__768_,data_stage_2__767_,data_stage_2__766_,data_stage_2__765_,
  data_stage_2__764_,data_stage_2__763_,data_stage_2__762_,data_stage_2__761_,
  data_stage_2__760_,data_stage_2__759_,data_stage_2__758_,data_stage_2__757_,
  data_stage_2__756_,data_stage_2__755_,data_stage_2__754_,data_stage_2__753_,
  data_stage_2__752_,data_stage_2__751_,data_stage_2__750_,data_stage_2__749_,data_stage_2__748_,
  data_stage_2__747_,data_stage_2__746_,data_stage_2__745_,data_stage_2__744_,
  data_stage_2__743_,data_stage_2__742_,data_stage_2__741_,data_stage_2__740_,
  data_stage_2__739_,data_stage_2__738_,data_stage_2__737_,data_stage_2__736_,
  data_stage_2__735_,data_stage_2__734_,data_stage_2__733_,data_stage_2__732_,
  data_stage_2__731_,data_stage_2__730_,data_stage_2__729_,data_stage_2__728_,data_stage_2__727_,
  data_stage_2__726_,data_stage_2__725_,data_stage_2__724_,data_stage_2__723_,
  data_stage_2__722_,data_stage_2__721_,data_stage_2__720_,data_stage_2__719_,
  data_stage_2__718_,data_stage_2__717_,data_stage_2__716_,data_stage_2__715_,
  data_stage_2__714_,data_stage_2__713_,data_stage_2__712_,data_stage_2__711_,data_stage_2__710_,
  data_stage_2__709_,data_stage_2__708_,data_stage_2__707_,data_stage_2__706_,
  data_stage_2__705_,data_stage_2__704_,data_stage_2__703_,data_stage_2__702_,
  data_stage_2__701_,data_stage_2__700_,data_stage_2__699_,data_stage_2__698_,
  data_stage_2__697_,data_stage_2__696_,data_stage_2__695_,data_stage_2__694_,
  data_stage_2__693_,data_stage_2__692_,data_stage_2__691_,data_stage_2__690_,data_stage_2__689_,
  data_stage_2__688_,data_stage_2__687_,data_stage_2__686_,data_stage_2__685_,
  data_stage_2__684_,data_stage_2__683_,data_stage_2__682_,data_stage_2__681_,
  data_stage_2__680_,data_stage_2__679_,data_stage_2__678_,data_stage_2__677_,
  data_stage_2__676_,data_stage_2__675_,data_stage_2__674_,data_stage_2__673_,
  data_stage_2__672_,data_stage_2__671_,data_stage_2__670_,data_stage_2__669_,data_stage_2__668_,
  data_stage_2__667_,data_stage_2__666_,data_stage_2__665_,data_stage_2__664_,
  data_stage_2__663_,data_stage_2__662_,data_stage_2__661_,data_stage_2__660_,
  data_stage_2__659_,data_stage_2__658_,data_stage_2__657_,data_stage_2__656_,
  data_stage_2__655_,data_stage_2__654_,data_stage_2__653_,data_stage_2__652_,
  data_stage_2__651_,data_stage_2__650_,data_stage_2__649_,data_stage_2__648_,data_stage_2__647_,
  data_stage_2__646_,data_stage_2__645_,data_stage_2__644_,data_stage_2__643_,
  data_stage_2__642_,data_stage_2__641_,data_stage_2__640_,data_stage_2__639_,
  data_stage_2__638_,data_stage_2__637_,data_stage_2__636_,data_stage_2__635_,
  data_stage_2__634_,data_stage_2__633_,data_stage_2__632_,data_stage_2__631_,data_stage_2__630_,
  data_stage_2__629_,data_stage_2__628_,data_stage_2__627_,data_stage_2__626_,
  data_stage_2__625_,data_stage_2__624_,data_stage_2__623_,data_stage_2__622_,
  data_stage_2__621_,data_stage_2__620_,data_stage_2__619_,data_stage_2__618_,
  data_stage_2__617_,data_stage_2__616_,data_stage_2__615_,data_stage_2__614_,
  data_stage_2__613_,data_stage_2__612_,data_stage_2__611_,data_stage_2__610_,data_stage_2__609_,
  data_stage_2__608_,data_stage_2__607_,data_stage_2__606_,data_stage_2__605_,
  data_stage_2__604_,data_stage_2__603_,data_stage_2__602_,data_stage_2__601_,
  data_stage_2__600_,data_stage_2__599_,data_stage_2__598_,data_stage_2__597_,
  data_stage_2__596_,data_stage_2__595_,data_stage_2__594_,data_stage_2__593_,
  data_stage_2__592_,data_stage_2__591_,data_stage_2__590_,data_stage_2__589_,data_stage_2__588_,
  data_stage_2__587_,data_stage_2__586_,data_stage_2__585_,data_stage_2__584_,
  data_stage_2__583_,data_stage_2__582_,data_stage_2__581_,data_stage_2__580_,
  data_stage_2__579_,data_stage_2__578_,data_stage_2__577_,data_stage_2__576_,
  data_stage_2__575_,data_stage_2__574_,data_stage_2__573_,data_stage_2__572_,
  data_stage_2__571_,data_stage_2__570_,data_stage_2__569_,data_stage_2__568_,data_stage_2__567_,
  data_stage_2__566_,data_stage_2__565_,data_stage_2__564_,data_stage_2__563_,
  data_stage_2__562_,data_stage_2__561_,data_stage_2__560_,data_stage_2__559_,
  data_stage_2__558_,data_stage_2__557_,data_stage_2__556_,data_stage_2__555_,
  data_stage_2__554_,data_stage_2__553_,data_stage_2__552_,data_stage_2__551_,data_stage_2__550_,
  data_stage_2__549_,data_stage_2__548_,data_stage_2__547_,data_stage_2__546_,
  data_stage_2__545_,data_stage_2__544_,data_stage_2__543_,data_stage_2__542_,
  data_stage_2__541_,data_stage_2__540_,data_stage_2__539_,data_stage_2__538_,
  data_stage_2__537_,data_stage_2__536_,data_stage_2__535_,data_stage_2__534_,
  data_stage_2__533_,data_stage_2__532_,data_stage_2__531_,data_stage_2__530_,data_stage_2__529_,
  data_stage_2__528_,data_stage_2__527_,data_stage_2__526_,data_stage_2__525_,
  data_stage_2__524_,data_stage_2__523_,data_stage_2__522_,data_stage_2__521_,
  data_stage_2__520_,data_stage_2__519_,data_stage_2__518_,data_stage_2__517_,
  data_stage_2__516_,data_stage_2__515_,data_stage_2__514_,data_stage_2__513_,
  data_stage_2__512_,data_stage_2__511_,data_stage_2__510_,data_stage_2__509_,data_stage_2__508_,
  data_stage_2__507_,data_stage_2__506_,data_stage_2__505_,data_stage_2__504_,
  data_stage_2__503_,data_stage_2__502_,data_stage_2__501_,data_stage_2__500_,
  data_stage_2__499_,data_stage_2__498_,data_stage_2__497_,data_stage_2__496_,
  data_stage_2__495_,data_stage_2__494_,data_stage_2__493_,data_stage_2__492_,
  data_stage_2__491_,data_stage_2__490_,data_stage_2__489_,data_stage_2__488_,data_stage_2__487_,
  data_stage_2__486_,data_stage_2__485_,data_stage_2__484_,data_stage_2__483_,
  data_stage_2__482_,data_stage_2__481_,data_stage_2__480_,data_stage_2__479_,
  data_stage_2__478_,data_stage_2__477_,data_stage_2__476_,data_stage_2__475_,
  data_stage_2__474_,data_stage_2__473_,data_stage_2__472_,data_stage_2__471_,data_stage_2__470_,
  data_stage_2__469_,data_stage_2__468_,data_stage_2__467_,data_stage_2__466_,
  data_stage_2__465_,data_stage_2__464_,data_stage_2__463_,data_stage_2__462_,
  data_stage_2__461_,data_stage_2__460_,data_stage_2__459_,data_stage_2__458_,
  data_stage_2__457_,data_stage_2__456_,data_stage_2__455_,data_stage_2__454_,
  data_stage_2__453_,data_stage_2__452_,data_stage_2__451_,data_stage_2__450_,data_stage_2__449_,
  data_stage_2__448_,data_stage_2__447_,data_stage_2__446_,data_stage_2__445_,
  data_stage_2__444_,data_stage_2__443_,data_stage_2__442_,data_stage_2__441_,
  data_stage_2__440_,data_stage_2__439_,data_stage_2__438_,data_stage_2__437_,
  data_stage_2__436_,data_stage_2__435_,data_stage_2__434_,data_stage_2__433_,
  data_stage_2__432_,data_stage_2__431_,data_stage_2__430_,data_stage_2__429_,data_stage_2__428_,
  data_stage_2__427_,data_stage_2__426_,data_stage_2__425_,data_stage_2__424_,
  data_stage_2__423_,data_stage_2__422_,data_stage_2__421_,data_stage_2__420_,
  data_stage_2__419_,data_stage_2__418_,data_stage_2__417_,data_stage_2__416_,
  data_stage_2__415_,data_stage_2__414_,data_stage_2__413_,data_stage_2__412_,
  data_stage_2__411_,data_stage_2__410_,data_stage_2__409_,data_stage_2__408_,data_stage_2__407_,
  data_stage_2__406_,data_stage_2__405_,data_stage_2__404_,data_stage_2__403_,
  data_stage_2__402_,data_stage_2__401_,data_stage_2__400_,data_stage_2__399_,
  data_stage_2__398_,data_stage_2__397_,data_stage_2__396_,data_stage_2__395_,
  data_stage_2__394_,data_stage_2__393_,data_stage_2__392_,data_stage_2__391_,data_stage_2__390_,
  data_stage_2__389_,data_stage_2__388_,data_stage_2__387_,data_stage_2__386_,
  data_stage_2__385_,data_stage_2__384_,data_stage_2__383_,data_stage_2__382_,
  data_stage_2__381_,data_stage_2__380_,data_stage_2__379_,data_stage_2__378_,
  data_stage_2__377_,data_stage_2__376_,data_stage_2__375_,data_stage_2__374_,
  data_stage_2__373_,data_stage_2__372_,data_stage_2__371_,data_stage_2__370_,data_stage_2__369_,
  data_stage_2__368_,data_stage_2__367_,data_stage_2__366_,data_stage_2__365_,
  data_stage_2__364_,data_stage_2__363_,data_stage_2__362_,data_stage_2__361_,
  data_stage_2__360_,data_stage_2__359_,data_stage_2__358_,data_stage_2__357_,
  data_stage_2__356_,data_stage_2__355_,data_stage_2__354_,data_stage_2__353_,
  data_stage_2__352_,data_stage_2__351_,data_stage_2__350_,data_stage_2__349_,data_stage_2__348_,
  data_stage_2__347_,data_stage_2__346_,data_stage_2__345_,data_stage_2__344_,
  data_stage_2__343_,data_stage_2__342_,data_stage_2__341_,data_stage_2__340_,
  data_stage_2__339_,data_stage_2__338_,data_stage_2__337_,data_stage_2__336_,
  data_stage_2__335_,data_stage_2__334_,data_stage_2__333_,data_stage_2__332_,
  data_stage_2__331_,data_stage_2__330_,data_stage_2__329_,data_stage_2__328_,data_stage_2__327_,
  data_stage_2__326_,data_stage_2__325_,data_stage_2__324_,data_stage_2__323_,
  data_stage_2__322_,data_stage_2__321_,data_stage_2__320_,data_stage_2__319_,
  data_stage_2__318_,data_stage_2__317_,data_stage_2__316_,data_stage_2__315_,
  data_stage_2__314_,data_stage_2__313_,data_stage_2__312_,data_stage_2__311_,data_stage_2__310_,
  data_stage_2__309_,data_stage_2__308_,data_stage_2__307_,data_stage_2__306_,
  data_stage_2__305_,data_stage_2__304_,data_stage_2__303_,data_stage_2__302_,
  data_stage_2__301_,data_stage_2__300_,data_stage_2__299_,data_stage_2__298_,
  data_stage_2__297_,data_stage_2__296_,data_stage_2__295_,data_stage_2__294_,
  data_stage_2__293_,data_stage_2__292_,data_stage_2__291_,data_stage_2__290_,data_stage_2__289_,
  data_stage_2__288_,data_stage_2__287_,data_stage_2__286_,data_stage_2__285_,
  data_stage_2__284_,data_stage_2__283_,data_stage_2__282_,data_stage_2__281_,
  data_stage_2__280_,data_stage_2__279_,data_stage_2__278_,data_stage_2__277_,
  data_stage_2__276_,data_stage_2__275_,data_stage_2__274_,data_stage_2__273_,
  data_stage_2__272_,data_stage_2__271_,data_stage_2__270_,data_stage_2__269_,data_stage_2__268_,
  data_stage_2__267_,data_stage_2__266_,data_stage_2__265_,data_stage_2__264_,
  data_stage_2__263_,data_stage_2__262_,data_stage_2__261_,data_stage_2__260_,
  data_stage_2__259_,data_stage_2__258_,data_stage_2__257_,data_stage_2__256_,
  data_stage_2__255_,data_stage_2__254_,data_stage_2__253_,data_stage_2__252_,
  data_stage_2__251_,data_stage_2__250_,data_stage_2__249_,data_stage_2__248_,data_stage_2__247_,
  data_stage_2__246_,data_stage_2__245_,data_stage_2__244_,data_stage_2__243_,
  data_stage_2__242_,data_stage_2__241_,data_stage_2__240_,data_stage_2__239_,
  data_stage_2__238_,data_stage_2__237_,data_stage_2__236_,data_stage_2__235_,
  data_stage_2__234_,data_stage_2__233_,data_stage_2__232_,data_stage_2__231_,data_stage_2__230_,
  data_stage_2__229_,data_stage_2__228_,data_stage_2__227_,data_stage_2__226_,
  data_stage_2__225_,data_stage_2__224_,data_stage_2__223_,data_stage_2__222_,
  data_stage_2__221_,data_stage_2__220_,data_stage_2__219_,data_stage_2__218_,
  data_stage_2__217_,data_stage_2__216_,data_stage_2__215_,data_stage_2__214_,
  data_stage_2__213_,data_stage_2__212_,data_stage_2__211_,data_stage_2__210_,data_stage_2__209_,
  data_stage_2__208_,data_stage_2__207_,data_stage_2__206_,data_stage_2__205_,
  data_stage_2__204_,data_stage_2__203_,data_stage_2__202_,data_stage_2__201_,
  data_stage_2__200_,data_stage_2__199_,data_stage_2__198_,data_stage_2__197_,
  data_stage_2__196_,data_stage_2__195_,data_stage_2__194_,data_stage_2__193_,
  data_stage_2__192_,data_stage_2__191_,data_stage_2__190_,data_stage_2__189_,data_stage_2__188_,
  data_stage_2__187_,data_stage_2__186_,data_stage_2__185_,data_stage_2__184_,
  data_stage_2__183_,data_stage_2__182_,data_stage_2__181_,data_stage_2__180_,
  data_stage_2__179_,data_stage_2__178_,data_stage_2__177_,data_stage_2__176_,
  data_stage_2__175_,data_stage_2__174_,data_stage_2__173_,data_stage_2__172_,
  data_stage_2__171_,data_stage_2__170_,data_stage_2__169_,data_stage_2__168_,data_stage_2__167_,
  data_stage_2__166_,data_stage_2__165_,data_stage_2__164_,data_stage_2__163_,
  data_stage_2__162_,data_stage_2__161_,data_stage_2__160_,data_stage_2__159_,
  data_stage_2__158_,data_stage_2__157_,data_stage_2__156_,data_stage_2__155_,
  data_stage_2__154_,data_stage_2__153_,data_stage_2__152_,data_stage_2__151_,data_stage_2__150_,
  data_stage_2__149_,data_stage_2__148_,data_stage_2__147_,data_stage_2__146_,
  data_stage_2__145_,data_stage_2__144_,data_stage_2__143_,data_stage_2__142_,
  data_stage_2__141_,data_stage_2__140_,data_stage_2__139_,data_stage_2__138_,
  data_stage_2__137_,data_stage_2__136_,data_stage_2__135_,data_stage_2__134_,
  data_stage_2__133_,data_stage_2__132_,data_stage_2__131_,data_stage_2__130_,data_stage_2__129_,
  data_stage_2__128_,data_stage_2__127_,data_stage_2__126_,data_stage_2__125_,
  data_stage_2__124_,data_stage_2__123_,data_stage_2__122_,data_stage_2__121_,
  data_stage_2__120_,data_stage_2__119_,data_stage_2__118_,data_stage_2__117_,
  data_stage_2__116_,data_stage_2__115_,data_stage_2__114_,data_stage_2__113_,
  data_stage_2__112_,data_stage_2__111_,data_stage_2__110_,data_stage_2__109_,data_stage_2__108_,
  data_stage_2__107_,data_stage_2__106_,data_stage_2__105_,data_stage_2__104_,
  data_stage_2__103_,data_stage_2__102_,data_stage_2__101_,data_stage_2__100_,
  data_stage_2__99_,data_stage_2__98_,data_stage_2__97_,data_stage_2__96_,data_stage_2__95_,
  data_stage_2__94_,data_stage_2__93_,data_stage_2__92_,data_stage_2__91_,
  data_stage_2__90_,data_stage_2__89_,data_stage_2__88_,data_stage_2__87_,
  data_stage_2__86_,data_stage_2__85_,data_stage_2__84_,data_stage_2__83_,data_stage_2__82_,
  data_stage_2__81_,data_stage_2__80_,data_stage_2__79_,data_stage_2__78_,
  data_stage_2__77_,data_stage_2__76_,data_stage_2__75_,data_stage_2__74_,data_stage_2__73_,
  data_stage_2__72_,data_stage_2__71_,data_stage_2__70_,data_stage_2__69_,
  data_stage_2__68_,data_stage_2__67_,data_stage_2__66_,data_stage_2__65_,data_stage_2__64_,
  data_stage_2__63_,data_stage_2__62_,data_stage_2__61_,data_stage_2__60_,
  data_stage_2__59_,data_stage_2__58_,data_stage_2__57_,data_stage_2__56_,data_stage_2__55_,
  data_stage_2__54_,data_stage_2__53_,data_stage_2__52_,data_stage_2__51_,
  data_stage_2__50_,data_stage_2__49_,data_stage_2__48_,data_stage_2__47_,
  data_stage_2__46_,data_stage_2__45_,data_stage_2__44_,data_stage_2__43_,data_stage_2__42_,
  data_stage_2__41_,data_stage_2__40_,data_stage_2__39_,data_stage_2__38_,
  data_stage_2__37_,data_stage_2__36_,data_stage_2__35_,data_stage_2__34_,data_stage_2__33_,
  data_stage_2__32_,data_stage_2__31_,data_stage_2__30_,data_stage_2__29_,
  data_stage_2__28_,data_stage_2__27_,data_stage_2__26_,data_stage_2__25_,data_stage_2__24_,
  data_stage_2__23_,data_stage_2__22_,data_stage_2__21_,data_stage_2__20_,
  data_stage_2__19_,data_stage_2__18_,data_stage_2__17_,data_stage_2__16_,data_stage_2__15_,
  data_stage_2__14_,data_stage_2__13_,data_stage_2__12_,data_stage_2__11_,
  data_stage_2__10_,data_stage_2__9_,data_stage_2__8_,data_stage_2__7_,data_stage_2__6_,
  data_stage_2__5_,data_stage_2__4_,data_stage_2__3_,data_stage_2__2_,
  data_stage_2__1_,data_stage_2__0_,data_stage_3__8191_,data_stage_3__8190_,data_stage_3__8189_,
  data_stage_3__8188_,data_stage_3__8187_,data_stage_3__8186_,data_stage_3__8185_,
  data_stage_3__8184_,data_stage_3__8183_,data_stage_3__8182_,data_stage_3__8181_,
  data_stage_3__8180_,data_stage_3__8179_,data_stage_3__8178_,data_stage_3__8177_,
  data_stage_3__8176_,data_stage_3__8175_,data_stage_3__8174_,data_stage_3__8173_,
  data_stage_3__8172_,data_stage_3__8171_,data_stage_3__8170_,data_stage_3__8169_,
  data_stage_3__8168_,data_stage_3__8167_,data_stage_3__8166_,data_stage_3__8165_,
  data_stage_3__8164_,data_stage_3__8163_,data_stage_3__8162_,data_stage_3__8161_,
  data_stage_3__8160_,data_stage_3__8159_,data_stage_3__8158_,data_stage_3__8157_,
  data_stage_3__8156_,data_stage_3__8155_,data_stage_3__8154_,data_stage_3__8153_,
  data_stage_3__8152_,data_stage_3__8151_,data_stage_3__8150_,data_stage_3__8149_,
  data_stage_3__8148_,data_stage_3__8147_,data_stage_3__8146_,data_stage_3__8145_,
  data_stage_3__8144_,data_stage_3__8143_,data_stage_3__8142_,data_stage_3__8141_,
  data_stage_3__8140_,data_stage_3__8139_,data_stage_3__8138_,data_stage_3__8137_,
  data_stage_3__8136_,data_stage_3__8135_,data_stage_3__8134_,data_stage_3__8133_,
  data_stage_3__8132_,data_stage_3__8131_,data_stage_3__8130_,data_stage_3__8129_,
  data_stage_3__8128_,data_stage_3__8127_,data_stage_3__8126_,data_stage_3__8125_,
  data_stage_3__8124_,data_stage_3__8123_,data_stage_3__8122_,data_stage_3__8121_,
  data_stage_3__8120_,data_stage_3__8119_,data_stage_3__8118_,data_stage_3__8117_,
  data_stage_3__8116_,data_stage_3__8115_,data_stage_3__8114_,data_stage_3__8113_,
  data_stage_3__8112_,data_stage_3__8111_,data_stage_3__8110_,data_stage_3__8109_,
  data_stage_3__8108_,data_stage_3__8107_,data_stage_3__8106_,data_stage_3__8105_,
  data_stage_3__8104_,data_stage_3__8103_,data_stage_3__8102_,data_stage_3__8101_,
  data_stage_3__8100_,data_stage_3__8099_,data_stage_3__8098_,data_stage_3__8097_,
  data_stage_3__8096_,data_stage_3__8095_,data_stage_3__8094_,data_stage_3__8093_,
  data_stage_3__8092_,data_stage_3__8091_,data_stage_3__8090_,data_stage_3__8089_,
  data_stage_3__8088_,data_stage_3__8087_,data_stage_3__8086_,data_stage_3__8085_,
  data_stage_3__8084_,data_stage_3__8083_,data_stage_3__8082_,data_stage_3__8081_,
  data_stage_3__8080_,data_stage_3__8079_,data_stage_3__8078_,data_stage_3__8077_,
  data_stage_3__8076_,data_stage_3__8075_,data_stage_3__8074_,data_stage_3__8073_,
  data_stage_3__8072_,data_stage_3__8071_,data_stage_3__8070_,data_stage_3__8069_,
  data_stage_3__8068_,data_stage_3__8067_,data_stage_3__8066_,data_stage_3__8065_,
  data_stage_3__8064_,data_stage_3__8063_,data_stage_3__8062_,data_stage_3__8061_,
  data_stage_3__8060_,data_stage_3__8059_,data_stage_3__8058_,data_stage_3__8057_,
  data_stage_3__8056_,data_stage_3__8055_,data_stage_3__8054_,data_stage_3__8053_,
  data_stage_3__8052_,data_stage_3__8051_,data_stage_3__8050_,data_stage_3__8049_,
  data_stage_3__8048_,data_stage_3__8047_,data_stage_3__8046_,data_stage_3__8045_,
  data_stage_3__8044_,data_stage_3__8043_,data_stage_3__8042_,data_stage_3__8041_,
  data_stage_3__8040_,data_stage_3__8039_,data_stage_3__8038_,data_stage_3__8037_,
  data_stage_3__8036_,data_stage_3__8035_,data_stage_3__8034_,data_stage_3__8033_,
  data_stage_3__8032_,data_stage_3__8031_,data_stage_3__8030_,data_stage_3__8029_,
  data_stage_3__8028_,data_stage_3__8027_,data_stage_3__8026_,data_stage_3__8025_,
  data_stage_3__8024_,data_stage_3__8023_,data_stage_3__8022_,data_stage_3__8021_,
  data_stage_3__8020_,data_stage_3__8019_,data_stage_3__8018_,data_stage_3__8017_,
  data_stage_3__8016_,data_stage_3__8015_,data_stage_3__8014_,data_stage_3__8013_,
  data_stage_3__8012_,data_stage_3__8011_,data_stage_3__8010_,data_stage_3__8009_,
  data_stage_3__8008_,data_stage_3__8007_,data_stage_3__8006_,data_stage_3__8005_,
  data_stage_3__8004_,data_stage_3__8003_,data_stage_3__8002_,data_stage_3__8001_,
  data_stage_3__8000_,data_stage_3__7999_,data_stage_3__7998_,data_stage_3__7997_,
  data_stage_3__7996_,data_stage_3__7995_,data_stage_3__7994_,data_stage_3__7993_,
  data_stage_3__7992_,data_stage_3__7991_,data_stage_3__7990_,data_stage_3__7989_,
  data_stage_3__7988_,data_stage_3__7987_,data_stage_3__7986_,data_stage_3__7985_,
  data_stage_3__7984_,data_stage_3__7983_,data_stage_3__7982_,data_stage_3__7981_,
  data_stage_3__7980_,data_stage_3__7979_,data_stage_3__7978_,data_stage_3__7977_,
  data_stage_3__7976_,data_stage_3__7975_,data_stage_3__7974_,data_stage_3__7973_,
  data_stage_3__7972_,data_stage_3__7971_,data_stage_3__7970_,data_stage_3__7969_,
  data_stage_3__7968_,data_stage_3__7967_,data_stage_3__7966_,data_stage_3__7965_,
  data_stage_3__7964_,data_stage_3__7963_,data_stage_3__7962_,data_stage_3__7961_,
  data_stage_3__7960_,data_stage_3__7959_,data_stage_3__7958_,data_stage_3__7957_,
  data_stage_3__7956_,data_stage_3__7955_,data_stage_3__7954_,data_stage_3__7953_,
  data_stage_3__7952_,data_stage_3__7951_,data_stage_3__7950_,data_stage_3__7949_,
  data_stage_3__7948_,data_stage_3__7947_,data_stage_3__7946_,data_stage_3__7945_,
  data_stage_3__7944_,data_stage_3__7943_,data_stage_3__7942_,data_stage_3__7941_,
  data_stage_3__7940_,data_stage_3__7939_,data_stage_3__7938_,data_stage_3__7937_,
  data_stage_3__7936_,data_stage_3__7935_,data_stage_3__7934_,data_stage_3__7933_,
  data_stage_3__7932_,data_stage_3__7931_,data_stage_3__7930_,data_stage_3__7929_,
  data_stage_3__7928_,data_stage_3__7927_,data_stage_3__7926_,data_stage_3__7925_,
  data_stage_3__7924_,data_stage_3__7923_,data_stage_3__7922_,data_stage_3__7921_,
  data_stage_3__7920_,data_stage_3__7919_,data_stage_3__7918_,data_stage_3__7917_,
  data_stage_3__7916_,data_stage_3__7915_,data_stage_3__7914_,data_stage_3__7913_,
  data_stage_3__7912_,data_stage_3__7911_,data_stage_3__7910_,data_stage_3__7909_,
  data_stage_3__7908_,data_stage_3__7907_,data_stage_3__7906_,data_stage_3__7905_,
  data_stage_3__7904_,data_stage_3__7903_,data_stage_3__7902_,data_stage_3__7901_,
  data_stage_3__7900_,data_stage_3__7899_,data_stage_3__7898_,data_stage_3__7897_,
  data_stage_3__7896_,data_stage_3__7895_,data_stage_3__7894_,data_stage_3__7893_,
  data_stage_3__7892_,data_stage_3__7891_,data_stage_3__7890_,data_stage_3__7889_,
  data_stage_3__7888_,data_stage_3__7887_,data_stage_3__7886_,data_stage_3__7885_,
  data_stage_3__7884_,data_stage_3__7883_,data_stage_3__7882_,data_stage_3__7881_,
  data_stage_3__7880_,data_stage_3__7879_,data_stage_3__7878_,data_stage_3__7877_,
  data_stage_3__7876_,data_stage_3__7875_,data_stage_3__7874_,data_stage_3__7873_,
  data_stage_3__7872_,data_stage_3__7871_,data_stage_3__7870_,data_stage_3__7869_,
  data_stage_3__7868_,data_stage_3__7867_,data_stage_3__7866_,data_stage_3__7865_,
  data_stage_3__7864_,data_stage_3__7863_,data_stage_3__7862_,data_stage_3__7861_,
  data_stage_3__7860_,data_stage_3__7859_,data_stage_3__7858_,data_stage_3__7857_,
  data_stage_3__7856_,data_stage_3__7855_,data_stage_3__7854_,data_stage_3__7853_,
  data_stage_3__7852_,data_stage_3__7851_,data_stage_3__7850_,data_stage_3__7849_,
  data_stage_3__7848_,data_stage_3__7847_,data_stage_3__7846_,data_stage_3__7845_,
  data_stage_3__7844_,data_stage_3__7843_,data_stage_3__7842_,data_stage_3__7841_,
  data_stage_3__7840_,data_stage_3__7839_,data_stage_3__7838_,data_stage_3__7837_,
  data_stage_3__7836_,data_stage_3__7835_,data_stage_3__7834_,data_stage_3__7833_,
  data_stage_3__7832_,data_stage_3__7831_,data_stage_3__7830_,data_stage_3__7829_,
  data_stage_3__7828_,data_stage_3__7827_,data_stage_3__7826_,data_stage_3__7825_,
  data_stage_3__7824_,data_stage_3__7823_,data_stage_3__7822_,data_stage_3__7821_,
  data_stage_3__7820_,data_stage_3__7819_,data_stage_3__7818_,data_stage_3__7817_,
  data_stage_3__7816_,data_stage_3__7815_,data_stage_3__7814_,data_stage_3__7813_,
  data_stage_3__7812_,data_stage_3__7811_,data_stage_3__7810_,data_stage_3__7809_,
  data_stage_3__7808_,data_stage_3__7807_,data_stage_3__7806_,data_stage_3__7805_,
  data_stage_3__7804_,data_stage_3__7803_,data_stage_3__7802_,data_stage_3__7801_,
  data_stage_3__7800_,data_stage_3__7799_,data_stage_3__7798_,data_stage_3__7797_,
  data_stage_3__7796_,data_stage_3__7795_,data_stage_3__7794_,data_stage_3__7793_,
  data_stage_3__7792_,data_stage_3__7791_,data_stage_3__7790_,data_stage_3__7789_,
  data_stage_3__7788_,data_stage_3__7787_,data_stage_3__7786_,data_stage_3__7785_,
  data_stage_3__7784_,data_stage_3__7783_,data_stage_3__7782_,data_stage_3__7781_,
  data_stage_3__7780_,data_stage_3__7779_,data_stage_3__7778_,data_stage_3__7777_,
  data_stage_3__7776_,data_stage_3__7775_,data_stage_3__7774_,data_stage_3__7773_,
  data_stage_3__7772_,data_stage_3__7771_,data_stage_3__7770_,data_stage_3__7769_,
  data_stage_3__7768_,data_stage_3__7767_,data_stage_3__7766_,data_stage_3__7765_,
  data_stage_3__7764_,data_stage_3__7763_,data_stage_3__7762_,data_stage_3__7761_,
  data_stage_3__7760_,data_stage_3__7759_,data_stage_3__7758_,data_stage_3__7757_,
  data_stage_3__7756_,data_stage_3__7755_,data_stage_3__7754_,data_stage_3__7753_,
  data_stage_3__7752_,data_stage_3__7751_,data_stage_3__7750_,data_stage_3__7749_,
  data_stage_3__7748_,data_stage_3__7747_,data_stage_3__7746_,data_stage_3__7745_,
  data_stage_3__7744_,data_stage_3__7743_,data_stage_3__7742_,data_stage_3__7741_,
  data_stage_3__7740_,data_stage_3__7739_,data_stage_3__7738_,data_stage_3__7737_,
  data_stage_3__7736_,data_stage_3__7735_,data_stage_3__7734_,data_stage_3__7733_,
  data_stage_3__7732_,data_stage_3__7731_,data_stage_3__7730_,data_stage_3__7729_,
  data_stage_3__7728_,data_stage_3__7727_,data_stage_3__7726_,data_stage_3__7725_,
  data_stage_3__7724_,data_stage_3__7723_,data_stage_3__7722_,data_stage_3__7721_,
  data_stage_3__7720_,data_stage_3__7719_,data_stage_3__7718_,data_stage_3__7717_,
  data_stage_3__7716_,data_stage_3__7715_,data_stage_3__7714_,data_stage_3__7713_,
  data_stage_3__7712_,data_stage_3__7711_,data_stage_3__7710_,data_stage_3__7709_,
  data_stage_3__7708_,data_stage_3__7707_,data_stage_3__7706_,data_stage_3__7705_,
  data_stage_3__7704_,data_stage_3__7703_,data_stage_3__7702_,data_stage_3__7701_,
  data_stage_3__7700_,data_stage_3__7699_,data_stage_3__7698_,data_stage_3__7697_,
  data_stage_3__7696_,data_stage_3__7695_,data_stage_3__7694_,data_stage_3__7693_,
  data_stage_3__7692_,data_stage_3__7691_,data_stage_3__7690_,data_stage_3__7689_,
  data_stage_3__7688_,data_stage_3__7687_,data_stage_3__7686_,data_stage_3__7685_,
  data_stage_3__7684_,data_stage_3__7683_,data_stage_3__7682_,data_stage_3__7681_,
  data_stage_3__7680_,data_stage_3__7679_,data_stage_3__7678_,data_stage_3__7677_,
  data_stage_3__7676_,data_stage_3__7675_,data_stage_3__7674_,data_stage_3__7673_,
  data_stage_3__7672_,data_stage_3__7671_,data_stage_3__7670_,data_stage_3__7669_,
  data_stage_3__7668_,data_stage_3__7667_,data_stage_3__7666_,data_stage_3__7665_,
  data_stage_3__7664_,data_stage_3__7663_,data_stage_3__7662_,data_stage_3__7661_,
  data_stage_3__7660_,data_stage_3__7659_,data_stage_3__7658_,data_stage_3__7657_,
  data_stage_3__7656_,data_stage_3__7655_,data_stage_3__7654_,data_stage_3__7653_,
  data_stage_3__7652_,data_stage_3__7651_,data_stage_3__7650_,data_stage_3__7649_,
  data_stage_3__7648_,data_stage_3__7647_,data_stage_3__7646_,data_stage_3__7645_,
  data_stage_3__7644_,data_stage_3__7643_,data_stage_3__7642_,data_stage_3__7641_,
  data_stage_3__7640_,data_stage_3__7639_,data_stage_3__7638_,data_stage_3__7637_,
  data_stage_3__7636_,data_stage_3__7635_,data_stage_3__7634_,data_stage_3__7633_,
  data_stage_3__7632_,data_stage_3__7631_,data_stage_3__7630_,data_stage_3__7629_,
  data_stage_3__7628_,data_stage_3__7627_,data_stage_3__7626_,data_stage_3__7625_,
  data_stage_3__7624_,data_stage_3__7623_,data_stage_3__7622_,data_stage_3__7621_,
  data_stage_3__7620_,data_stage_3__7619_,data_stage_3__7618_,data_stage_3__7617_,
  data_stage_3__7616_,data_stage_3__7615_,data_stage_3__7614_,data_stage_3__7613_,
  data_stage_3__7612_,data_stage_3__7611_,data_stage_3__7610_,data_stage_3__7609_,
  data_stage_3__7608_,data_stage_3__7607_,data_stage_3__7606_,data_stage_3__7605_,
  data_stage_3__7604_,data_stage_3__7603_,data_stage_3__7602_,data_stage_3__7601_,
  data_stage_3__7600_,data_stage_3__7599_,data_stage_3__7598_,data_stage_3__7597_,
  data_stage_3__7596_,data_stage_3__7595_,data_stage_3__7594_,data_stage_3__7593_,
  data_stage_3__7592_,data_stage_3__7591_,data_stage_3__7590_,data_stage_3__7589_,
  data_stage_3__7588_,data_stage_3__7587_,data_stage_3__7586_,data_stage_3__7585_,
  data_stage_3__7584_,data_stage_3__7583_,data_stage_3__7582_,data_stage_3__7581_,
  data_stage_3__7580_,data_stage_3__7579_,data_stage_3__7578_,data_stage_3__7577_,
  data_stage_3__7576_,data_stage_3__7575_,data_stage_3__7574_,data_stage_3__7573_,
  data_stage_3__7572_,data_stage_3__7571_,data_stage_3__7570_,data_stage_3__7569_,
  data_stage_3__7568_,data_stage_3__7567_,data_stage_3__7566_,data_stage_3__7565_,
  data_stage_3__7564_,data_stage_3__7563_,data_stage_3__7562_,data_stage_3__7561_,
  data_stage_3__7560_,data_stage_3__7559_,data_stage_3__7558_,data_stage_3__7557_,
  data_stage_3__7556_,data_stage_3__7555_,data_stage_3__7554_,data_stage_3__7553_,
  data_stage_3__7552_,data_stage_3__7551_,data_stage_3__7550_,data_stage_3__7549_,
  data_stage_3__7548_,data_stage_3__7547_,data_stage_3__7546_,data_stage_3__7545_,
  data_stage_3__7544_,data_stage_3__7543_,data_stage_3__7542_,data_stage_3__7541_,
  data_stage_3__7540_,data_stage_3__7539_,data_stage_3__7538_,data_stage_3__7537_,
  data_stage_3__7536_,data_stage_3__7535_,data_stage_3__7534_,data_stage_3__7533_,
  data_stage_3__7532_,data_stage_3__7531_,data_stage_3__7530_,data_stage_3__7529_,
  data_stage_3__7528_,data_stage_3__7527_,data_stage_3__7526_,data_stage_3__7525_,
  data_stage_3__7524_,data_stage_3__7523_,data_stage_3__7522_,data_stage_3__7521_,
  data_stage_3__7520_,data_stage_3__7519_,data_stage_3__7518_,data_stage_3__7517_,
  data_stage_3__7516_,data_stage_3__7515_,data_stage_3__7514_,data_stage_3__7513_,
  data_stage_3__7512_,data_stage_3__7511_,data_stage_3__7510_,data_stage_3__7509_,
  data_stage_3__7508_,data_stage_3__7507_,data_stage_3__7506_,data_stage_3__7505_,
  data_stage_3__7504_,data_stage_3__7503_,data_stage_3__7502_,data_stage_3__7501_,
  data_stage_3__7500_,data_stage_3__7499_,data_stage_3__7498_,data_stage_3__7497_,
  data_stage_3__7496_,data_stage_3__7495_,data_stage_3__7494_,data_stage_3__7493_,
  data_stage_3__7492_,data_stage_3__7491_,data_stage_3__7490_,data_stage_3__7489_,
  data_stage_3__7488_,data_stage_3__7487_,data_stage_3__7486_,data_stage_3__7485_,
  data_stage_3__7484_,data_stage_3__7483_,data_stage_3__7482_,data_stage_3__7481_,
  data_stage_3__7480_,data_stage_3__7479_,data_stage_3__7478_,data_stage_3__7477_,
  data_stage_3__7476_,data_stage_3__7475_,data_stage_3__7474_,data_stage_3__7473_,
  data_stage_3__7472_,data_stage_3__7471_,data_stage_3__7470_,data_stage_3__7469_,
  data_stage_3__7468_,data_stage_3__7467_,data_stage_3__7466_,data_stage_3__7465_,
  data_stage_3__7464_,data_stage_3__7463_,data_stage_3__7462_,data_stage_3__7461_,
  data_stage_3__7460_,data_stage_3__7459_,data_stage_3__7458_,data_stage_3__7457_,
  data_stage_3__7456_,data_stage_3__7455_,data_stage_3__7454_,data_stage_3__7453_,
  data_stage_3__7452_,data_stage_3__7451_,data_stage_3__7450_,data_stage_3__7449_,
  data_stage_3__7448_,data_stage_3__7447_,data_stage_3__7446_,data_stage_3__7445_,
  data_stage_3__7444_,data_stage_3__7443_,data_stage_3__7442_,data_stage_3__7441_,
  data_stage_3__7440_,data_stage_3__7439_,data_stage_3__7438_,data_stage_3__7437_,
  data_stage_3__7436_,data_stage_3__7435_,data_stage_3__7434_,data_stage_3__7433_,
  data_stage_3__7432_,data_stage_3__7431_,data_stage_3__7430_,data_stage_3__7429_,
  data_stage_3__7428_,data_stage_3__7427_,data_stage_3__7426_,data_stage_3__7425_,
  data_stage_3__7424_,data_stage_3__7423_,data_stage_3__7422_,data_stage_3__7421_,
  data_stage_3__7420_,data_stage_3__7419_,data_stage_3__7418_,data_stage_3__7417_,
  data_stage_3__7416_,data_stage_3__7415_,data_stage_3__7414_,data_stage_3__7413_,
  data_stage_3__7412_,data_stage_3__7411_,data_stage_3__7410_,data_stage_3__7409_,
  data_stage_3__7408_,data_stage_3__7407_,data_stage_3__7406_,data_stage_3__7405_,
  data_stage_3__7404_,data_stage_3__7403_,data_stage_3__7402_,data_stage_3__7401_,
  data_stage_3__7400_,data_stage_3__7399_,data_stage_3__7398_,data_stage_3__7397_,
  data_stage_3__7396_,data_stage_3__7395_,data_stage_3__7394_,data_stage_3__7393_,
  data_stage_3__7392_,data_stage_3__7391_,data_stage_3__7390_,data_stage_3__7389_,
  data_stage_3__7388_,data_stage_3__7387_,data_stage_3__7386_,data_stage_3__7385_,
  data_stage_3__7384_,data_stage_3__7383_,data_stage_3__7382_,data_stage_3__7381_,
  data_stage_3__7380_,data_stage_3__7379_,data_stage_3__7378_,data_stage_3__7377_,
  data_stage_3__7376_,data_stage_3__7375_,data_stage_3__7374_,data_stage_3__7373_,
  data_stage_3__7372_,data_stage_3__7371_,data_stage_3__7370_,data_stage_3__7369_,
  data_stage_3__7368_,data_stage_3__7367_,data_stage_3__7366_,data_stage_3__7365_,
  data_stage_3__7364_,data_stage_3__7363_,data_stage_3__7362_,data_stage_3__7361_,
  data_stage_3__7360_,data_stage_3__7359_,data_stage_3__7358_,data_stage_3__7357_,
  data_stage_3__7356_,data_stage_3__7355_,data_stage_3__7354_,data_stage_3__7353_,
  data_stage_3__7352_,data_stage_3__7351_,data_stage_3__7350_,data_stage_3__7349_,
  data_stage_3__7348_,data_stage_3__7347_,data_stage_3__7346_,data_stage_3__7345_,
  data_stage_3__7344_,data_stage_3__7343_,data_stage_3__7342_,data_stage_3__7341_,
  data_stage_3__7340_,data_stage_3__7339_,data_stage_3__7338_,data_stage_3__7337_,
  data_stage_3__7336_,data_stage_3__7335_,data_stage_3__7334_,data_stage_3__7333_,
  data_stage_3__7332_,data_stage_3__7331_,data_stage_3__7330_,data_stage_3__7329_,
  data_stage_3__7328_,data_stage_3__7327_,data_stage_3__7326_,data_stage_3__7325_,
  data_stage_3__7324_,data_stage_3__7323_,data_stage_3__7322_,data_stage_3__7321_,
  data_stage_3__7320_,data_stage_3__7319_,data_stage_3__7318_,data_stage_3__7317_,
  data_stage_3__7316_,data_stage_3__7315_,data_stage_3__7314_,data_stage_3__7313_,
  data_stage_3__7312_,data_stage_3__7311_,data_stage_3__7310_,data_stage_3__7309_,
  data_stage_3__7308_,data_stage_3__7307_,data_stage_3__7306_,data_stage_3__7305_,
  data_stage_3__7304_,data_stage_3__7303_,data_stage_3__7302_,data_stage_3__7301_,
  data_stage_3__7300_,data_stage_3__7299_,data_stage_3__7298_,data_stage_3__7297_,
  data_stage_3__7296_,data_stage_3__7295_,data_stage_3__7294_,data_stage_3__7293_,
  data_stage_3__7292_,data_stage_3__7291_,data_stage_3__7290_,data_stage_3__7289_,
  data_stage_3__7288_,data_stage_3__7287_,data_stage_3__7286_,data_stage_3__7285_,
  data_stage_3__7284_,data_stage_3__7283_,data_stage_3__7282_,data_stage_3__7281_,
  data_stage_3__7280_,data_stage_3__7279_,data_stage_3__7278_,data_stage_3__7277_,
  data_stage_3__7276_,data_stage_3__7275_,data_stage_3__7274_,data_stage_3__7273_,
  data_stage_3__7272_,data_stage_3__7271_,data_stage_3__7270_,data_stage_3__7269_,
  data_stage_3__7268_,data_stage_3__7267_,data_stage_3__7266_,data_stage_3__7265_,
  data_stage_3__7264_,data_stage_3__7263_,data_stage_3__7262_,data_stage_3__7261_,
  data_stage_3__7260_,data_stage_3__7259_,data_stage_3__7258_,data_stage_3__7257_,
  data_stage_3__7256_,data_stage_3__7255_,data_stage_3__7254_,data_stage_3__7253_,
  data_stage_3__7252_,data_stage_3__7251_,data_stage_3__7250_,data_stage_3__7249_,
  data_stage_3__7248_,data_stage_3__7247_,data_stage_3__7246_,data_stage_3__7245_,
  data_stage_3__7244_,data_stage_3__7243_,data_stage_3__7242_,data_stage_3__7241_,
  data_stage_3__7240_,data_stage_3__7239_,data_stage_3__7238_,data_stage_3__7237_,
  data_stage_3__7236_,data_stage_3__7235_,data_stage_3__7234_,data_stage_3__7233_,
  data_stage_3__7232_,data_stage_3__7231_,data_stage_3__7230_,data_stage_3__7229_,
  data_stage_3__7228_,data_stage_3__7227_,data_stage_3__7226_,data_stage_3__7225_,
  data_stage_3__7224_,data_stage_3__7223_,data_stage_3__7222_,data_stage_3__7221_,
  data_stage_3__7220_,data_stage_3__7219_,data_stage_3__7218_,data_stage_3__7217_,
  data_stage_3__7216_,data_stage_3__7215_,data_stage_3__7214_,data_stage_3__7213_,
  data_stage_3__7212_,data_stage_3__7211_,data_stage_3__7210_,data_stage_3__7209_,
  data_stage_3__7208_,data_stage_3__7207_,data_stage_3__7206_,data_stage_3__7205_,
  data_stage_3__7204_,data_stage_3__7203_,data_stage_3__7202_,data_stage_3__7201_,
  data_stage_3__7200_,data_stage_3__7199_,data_stage_3__7198_,data_stage_3__7197_,
  data_stage_3__7196_,data_stage_3__7195_,data_stage_3__7194_,data_stage_3__7193_,
  data_stage_3__7192_,data_stage_3__7191_,data_stage_3__7190_,data_stage_3__7189_,
  data_stage_3__7188_,data_stage_3__7187_,data_stage_3__7186_,data_stage_3__7185_,
  data_stage_3__7184_,data_stage_3__7183_,data_stage_3__7182_,data_stage_3__7181_,
  data_stage_3__7180_,data_stage_3__7179_,data_stage_3__7178_,data_stage_3__7177_,
  data_stage_3__7176_,data_stage_3__7175_,data_stage_3__7174_,data_stage_3__7173_,
  data_stage_3__7172_,data_stage_3__7171_,data_stage_3__7170_,data_stage_3__7169_,
  data_stage_3__7168_,data_stage_3__7167_,data_stage_3__7166_,data_stage_3__7165_,
  data_stage_3__7164_,data_stage_3__7163_,data_stage_3__7162_,data_stage_3__7161_,
  data_stage_3__7160_,data_stage_3__7159_,data_stage_3__7158_,data_stage_3__7157_,
  data_stage_3__7156_,data_stage_3__7155_,data_stage_3__7154_,data_stage_3__7153_,
  data_stage_3__7152_,data_stage_3__7151_,data_stage_3__7150_,data_stage_3__7149_,
  data_stage_3__7148_,data_stage_3__7147_,data_stage_3__7146_,data_stage_3__7145_,
  data_stage_3__7144_,data_stage_3__7143_,data_stage_3__7142_,data_stage_3__7141_,
  data_stage_3__7140_,data_stage_3__7139_,data_stage_3__7138_,data_stage_3__7137_,
  data_stage_3__7136_,data_stage_3__7135_,data_stage_3__7134_,data_stage_3__7133_,
  data_stage_3__7132_,data_stage_3__7131_,data_stage_3__7130_,data_stage_3__7129_,
  data_stage_3__7128_,data_stage_3__7127_,data_stage_3__7126_,data_stage_3__7125_,
  data_stage_3__7124_,data_stage_3__7123_,data_stage_3__7122_,data_stage_3__7121_,
  data_stage_3__7120_,data_stage_3__7119_,data_stage_3__7118_,data_stage_3__7117_,
  data_stage_3__7116_,data_stage_3__7115_,data_stage_3__7114_,data_stage_3__7113_,
  data_stage_3__7112_,data_stage_3__7111_,data_stage_3__7110_,data_stage_3__7109_,
  data_stage_3__7108_,data_stage_3__7107_,data_stage_3__7106_,data_stage_3__7105_,
  data_stage_3__7104_,data_stage_3__7103_,data_stage_3__7102_,data_stage_3__7101_,
  data_stage_3__7100_,data_stage_3__7099_,data_stage_3__7098_,data_stage_3__7097_,
  data_stage_3__7096_,data_stage_3__7095_,data_stage_3__7094_,data_stage_3__7093_,
  data_stage_3__7092_,data_stage_3__7091_,data_stage_3__7090_,data_stage_3__7089_,
  data_stage_3__7088_,data_stage_3__7087_,data_stage_3__7086_,data_stage_3__7085_,
  data_stage_3__7084_,data_stage_3__7083_,data_stage_3__7082_,data_stage_3__7081_,
  data_stage_3__7080_,data_stage_3__7079_,data_stage_3__7078_,data_stage_3__7077_,
  data_stage_3__7076_,data_stage_3__7075_,data_stage_3__7074_,data_stage_3__7073_,
  data_stage_3__7072_,data_stage_3__7071_,data_stage_3__7070_,data_stage_3__7069_,
  data_stage_3__7068_,data_stage_3__7067_,data_stage_3__7066_,data_stage_3__7065_,
  data_stage_3__7064_,data_stage_3__7063_,data_stage_3__7062_,data_stage_3__7061_,
  data_stage_3__7060_,data_stage_3__7059_,data_stage_3__7058_,data_stage_3__7057_,
  data_stage_3__7056_,data_stage_3__7055_,data_stage_3__7054_,data_stage_3__7053_,
  data_stage_3__7052_,data_stage_3__7051_,data_stage_3__7050_,data_stage_3__7049_,
  data_stage_3__7048_,data_stage_3__7047_,data_stage_3__7046_,data_stage_3__7045_,
  data_stage_3__7044_,data_stage_3__7043_,data_stage_3__7042_,data_stage_3__7041_,
  data_stage_3__7040_,data_stage_3__7039_,data_stage_3__7038_,data_stage_3__7037_,
  data_stage_3__7036_,data_stage_3__7035_,data_stage_3__7034_,data_stage_3__7033_,
  data_stage_3__7032_,data_stage_3__7031_,data_stage_3__7030_,data_stage_3__7029_,
  data_stage_3__7028_,data_stage_3__7027_,data_stage_3__7026_,data_stage_3__7025_,
  data_stage_3__7024_,data_stage_3__7023_,data_stage_3__7022_,data_stage_3__7021_,
  data_stage_3__7020_,data_stage_3__7019_,data_stage_3__7018_,data_stage_3__7017_,
  data_stage_3__7016_,data_stage_3__7015_,data_stage_3__7014_,data_stage_3__7013_,
  data_stage_3__7012_,data_stage_3__7011_,data_stage_3__7010_,data_stage_3__7009_,
  data_stage_3__7008_,data_stage_3__7007_,data_stage_3__7006_,data_stage_3__7005_,
  data_stage_3__7004_,data_stage_3__7003_,data_stage_3__7002_,data_stage_3__7001_,
  data_stage_3__7000_,data_stage_3__6999_,data_stage_3__6998_,data_stage_3__6997_,
  data_stage_3__6996_,data_stage_3__6995_,data_stage_3__6994_,data_stage_3__6993_,
  data_stage_3__6992_,data_stage_3__6991_,data_stage_3__6990_,data_stage_3__6989_,
  data_stage_3__6988_,data_stage_3__6987_,data_stage_3__6986_,data_stage_3__6985_,
  data_stage_3__6984_,data_stage_3__6983_,data_stage_3__6982_,data_stage_3__6981_,
  data_stage_3__6980_,data_stage_3__6979_,data_stage_3__6978_,data_stage_3__6977_,
  data_stage_3__6976_,data_stage_3__6975_,data_stage_3__6974_,data_stage_3__6973_,
  data_stage_3__6972_,data_stage_3__6971_,data_stage_3__6970_,data_stage_3__6969_,
  data_stage_3__6968_,data_stage_3__6967_,data_stage_3__6966_,data_stage_3__6965_,
  data_stage_3__6964_,data_stage_3__6963_,data_stage_3__6962_,data_stage_3__6961_,
  data_stage_3__6960_,data_stage_3__6959_,data_stage_3__6958_,data_stage_3__6957_,
  data_stage_3__6956_,data_stage_3__6955_,data_stage_3__6954_,data_stage_3__6953_,
  data_stage_3__6952_,data_stage_3__6951_,data_stage_3__6950_,data_stage_3__6949_,
  data_stage_3__6948_,data_stage_3__6947_,data_stage_3__6946_,data_stage_3__6945_,
  data_stage_3__6944_,data_stage_3__6943_,data_stage_3__6942_,data_stage_3__6941_,
  data_stage_3__6940_,data_stage_3__6939_,data_stage_3__6938_,data_stage_3__6937_,
  data_stage_3__6936_,data_stage_3__6935_,data_stage_3__6934_,data_stage_3__6933_,
  data_stage_3__6932_,data_stage_3__6931_,data_stage_3__6930_,data_stage_3__6929_,
  data_stage_3__6928_,data_stage_3__6927_,data_stage_3__6926_,data_stage_3__6925_,
  data_stage_3__6924_,data_stage_3__6923_,data_stage_3__6922_,data_stage_3__6921_,
  data_stage_3__6920_,data_stage_3__6919_,data_stage_3__6918_,data_stage_3__6917_,
  data_stage_3__6916_,data_stage_3__6915_,data_stage_3__6914_,data_stage_3__6913_,
  data_stage_3__6912_,data_stage_3__6911_,data_stage_3__6910_,data_stage_3__6909_,
  data_stage_3__6908_,data_stage_3__6907_,data_stage_3__6906_,data_stage_3__6905_,
  data_stage_3__6904_,data_stage_3__6903_,data_stage_3__6902_,data_stage_3__6901_,
  data_stage_3__6900_,data_stage_3__6899_,data_stage_3__6898_,data_stage_3__6897_,
  data_stage_3__6896_,data_stage_3__6895_,data_stage_3__6894_,data_stage_3__6893_,
  data_stage_3__6892_,data_stage_3__6891_,data_stage_3__6890_,data_stage_3__6889_,
  data_stage_3__6888_,data_stage_3__6887_,data_stage_3__6886_,data_stage_3__6885_,
  data_stage_3__6884_,data_stage_3__6883_,data_stage_3__6882_,data_stage_3__6881_,
  data_stage_3__6880_,data_stage_3__6879_,data_stage_3__6878_,data_stage_3__6877_,
  data_stage_3__6876_,data_stage_3__6875_,data_stage_3__6874_,data_stage_3__6873_,
  data_stage_3__6872_,data_stage_3__6871_,data_stage_3__6870_,data_stage_3__6869_,
  data_stage_3__6868_,data_stage_3__6867_,data_stage_3__6866_,data_stage_3__6865_,
  data_stage_3__6864_,data_stage_3__6863_,data_stage_3__6862_,data_stage_3__6861_,
  data_stage_3__6860_,data_stage_3__6859_,data_stage_3__6858_,data_stage_3__6857_,
  data_stage_3__6856_,data_stage_3__6855_,data_stage_3__6854_,data_stage_3__6853_,
  data_stage_3__6852_,data_stage_3__6851_,data_stage_3__6850_,data_stage_3__6849_,
  data_stage_3__6848_,data_stage_3__6847_,data_stage_3__6846_,data_stage_3__6845_,
  data_stage_3__6844_,data_stage_3__6843_,data_stage_3__6842_,data_stage_3__6841_,
  data_stage_3__6840_,data_stage_3__6839_,data_stage_3__6838_,data_stage_3__6837_,
  data_stage_3__6836_,data_stage_3__6835_,data_stage_3__6834_,data_stage_3__6833_,
  data_stage_3__6832_,data_stage_3__6831_,data_stage_3__6830_,data_stage_3__6829_,
  data_stage_3__6828_,data_stage_3__6827_,data_stage_3__6826_,data_stage_3__6825_,
  data_stage_3__6824_,data_stage_3__6823_,data_stage_3__6822_,data_stage_3__6821_,
  data_stage_3__6820_,data_stage_3__6819_,data_stage_3__6818_,data_stage_3__6817_,
  data_stage_3__6816_,data_stage_3__6815_,data_stage_3__6814_,data_stage_3__6813_,
  data_stage_3__6812_,data_stage_3__6811_,data_stage_3__6810_,data_stage_3__6809_,
  data_stage_3__6808_,data_stage_3__6807_,data_stage_3__6806_,data_stage_3__6805_,
  data_stage_3__6804_,data_stage_3__6803_,data_stage_3__6802_,data_stage_3__6801_,
  data_stage_3__6800_,data_stage_3__6799_,data_stage_3__6798_,data_stage_3__6797_,
  data_stage_3__6796_,data_stage_3__6795_,data_stage_3__6794_,data_stage_3__6793_,
  data_stage_3__6792_,data_stage_3__6791_,data_stage_3__6790_,data_stage_3__6789_,
  data_stage_3__6788_,data_stage_3__6787_,data_stage_3__6786_,data_stage_3__6785_,
  data_stage_3__6784_,data_stage_3__6783_,data_stage_3__6782_,data_stage_3__6781_,
  data_stage_3__6780_,data_stage_3__6779_,data_stage_3__6778_,data_stage_3__6777_,
  data_stage_3__6776_,data_stage_3__6775_,data_stage_3__6774_,data_stage_3__6773_,
  data_stage_3__6772_,data_stage_3__6771_,data_stage_3__6770_,data_stage_3__6769_,
  data_stage_3__6768_,data_stage_3__6767_,data_stage_3__6766_,data_stage_3__6765_,
  data_stage_3__6764_,data_stage_3__6763_,data_stage_3__6762_,data_stage_3__6761_,
  data_stage_3__6760_,data_stage_3__6759_,data_stage_3__6758_,data_stage_3__6757_,
  data_stage_3__6756_,data_stage_3__6755_,data_stage_3__6754_,data_stage_3__6753_,
  data_stage_3__6752_,data_stage_3__6751_,data_stage_3__6750_,data_stage_3__6749_,
  data_stage_3__6748_,data_stage_3__6747_,data_stage_3__6746_,data_stage_3__6745_,
  data_stage_3__6744_,data_stage_3__6743_,data_stage_3__6742_,data_stage_3__6741_,
  data_stage_3__6740_,data_stage_3__6739_,data_stage_3__6738_,data_stage_3__6737_,
  data_stage_3__6736_,data_stage_3__6735_,data_stage_3__6734_,data_stage_3__6733_,
  data_stage_3__6732_,data_stage_3__6731_,data_stage_3__6730_,data_stage_3__6729_,
  data_stage_3__6728_,data_stage_3__6727_,data_stage_3__6726_,data_stage_3__6725_,
  data_stage_3__6724_,data_stage_3__6723_,data_stage_3__6722_,data_stage_3__6721_,
  data_stage_3__6720_,data_stage_3__6719_,data_stage_3__6718_,data_stage_3__6717_,
  data_stage_3__6716_,data_stage_3__6715_,data_stage_3__6714_,data_stage_3__6713_,
  data_stage_3__6712_,data_stage_3__6711_,data_stage_3__6710_,data_stage_3__6709_,
  data_stage_3__6708_,data_stage_3__6707_,data_stage_3__6706_,data_stage_3__6705_,
  data_stage_3__6704_,data_stage_3__6703_,data_stage_3__6702_,data_stage_3__6701_,
  data_stage_3__6700_,data_stage_3__6699_,data_stage_3__6698_,data_stage_3__6697_,
  data_stage_3__6696_,data_stage_3__6695_,data_stage_3__6694_,data_stage_3__6693_,
  data_stage_3__6692_,data_stage_3__6691_,data_stage_3__6690_,data_stage_3__6689_,
  data_stage_3__6688_,data_stage_3__6687_,data_stage_3__6686_,data_stage_3__6685_,
  data_stage_3__6684_,data_stage_3__6683_,data_stage_3__6682_,data_stage_3__6681_,
  data_stage_3__6680_,data_stage_3__6679_,data_stage_3__6678_,data_stage_3__6677_,
  data_stage_3__6676_,data_stage_3__6675_,data_stage_3__6674_,data_stage_3__6673_,
  data_stage_3__6672_,data_stage_3__6671_,data_stage_3__6670_,data_stage_3__6669_,
  data_stage_3__6668_,data_stage_3__6667_,data_stage_3__6666_,data_stage_3__6665_,
  data_stage_3__6664_,data_stage_3__6663_,data_stage_3__6662_,data_stage_3__6661_,
  data_stage_3__6660_,data_stage_3__6659_,data_stage_3__6658_,data_stage_3__6657_,
  data_stage_3__6656_,data_stage_3__6655_,data_stage_3__6654_,data_stage_3__6653_,
  data_stage_3__6652_,data_stage_3__6651_,data_stage_3__6650_,data_stage_3__6649_,
  data_stage_3__6648_,data_stage_3__6647_,data_stage_3__6646_,data_stage_3__6645_,
  data_stage_3__6644_,data_stage_3__6643_,data_stage_3__6642_,data_stage_3__6641_,
  data_stage_3__6640_,data_stage_3__6639_,data_stage_3__6638_,data_stage_3__6637_,
  data_stage_3__6636_,data_stage_3__6635_,data_stage_3__6634_,data_stage_3__6633_,
  data_stage_3__6632_,data_stage_3__6631_,data_stage_3__6630_,data_stage_3__6629_,
  data_stage_3__6628_,data_stage_3__6627_,data_stage_3__6626_,data_stage_3__6625_,
  data_stage_3__6624_,data_stage_3__6623_,data_stage_3__6622_,data_stage_3__6621_,
  data_stage_3__6620_,data_stage_3__6619_,data_stage_3__6618_,data_stage_3__6617_,
  data_stage_3__6616_,data_stage_3__6615_,data_stage_3__6614_,data_stage_3__6613_,
  data_stage_3__6612_,data_stage_3__6611_,data_stage_3__6610_,data_stage_3__6609_,
  data_stage_3__6608_,data_stage_3__6607_,data_stage_3__6606_,data_stage_3__6605_,
  data_stage_3__6604_,data_stage_3__6603_,data_stage_3__6602_,data_stage_3__6601_,
  data_stage_3__6600_,data_stage_3__6599_,data_stage_3__6598_,data_stage_3__6597_,
  data_stage_3__6596_,data_stage_3__6595_,data_stage_3__6594_,data_stage_3__6593_,
  data_stage_3__6592_,data_stage_3__6591_,data_stage_3__6590_,data_stage_3__6589_,
  data_stage_3__6588_,data_stage_3__6587_,data_stage_3__6586_,data_stage_3__6585_,
  data_stage_3__6584_,data_stage_3__6583_,data_stage_3__6582_,data_stage_3__6581_,
  data_stage_3__6580_,data_stage_3__6579_,data_stage_3__6578_,data_stage_3__6577_,
  data_stage_3__6576_,data_stage_3__6575_,data_stage_3__6574_,data_stage_3__6573_,
  data_stage_3__6572_,data_stage_3__6571_,data_stage_3__6570_,data_stage_3__6569_,
  data_stage_3__6568_,data_stage_3__6567_,data_stage_3__6566_,data_stage_3__6565_,
  data_stage_3__6564_,data_stage_3__6563_,data_stage_3__6562_,data_stage_3__6561_,
  data_stage_3__6560_,data_stage_3__6559_,data_stage_3__6558_,data_stage_3__6557_,
  data_stage_3__6556_,data_stage_3__6555_,data_stage_3__6554_,data_stage_3__6553_,
  data_stage_3__6552_,data_stage_3__6551_,data_stage_3__6550_,data_stage_3__6549_,
  data_stage_3__6548_,data_stage_3__6547_,data_stage_3__6546_,data_stage_3__6545_,
  data_stage_3__6544_,data_stage_3__6543_,data_stage_3__6542_,data_stage_3__6541_,
  data_stage_3__6540_,data_stage_3__6539_,data_stage_3__6538_,data_stage_3__6537_,
  data_stage_3__6536_,data_stage_3__6535_,data_stage_3__6534_,data_stage_3__6533_,
  data_stage_3__6532_,data_stage_3__6531_,data_stage_3__6530_,data_stage_3__6529_,
  data_stage_3__6528_,data_stage_3__6527_,data_stage_3__6526_,data_stage_3__6525_,
  data_stage_3__6524_,data_stage_3__6523_,data_stage_3__6522_,data_stage_3__6521_,
  data_stage_3__6520_,data_stage_3__6519_,data_stage_3__6518_,data_stage_3__6517_,
  data_stage_3__6516_,data_stage_3__6515_,data_stage_3__6514_,data_stage_3__6513_,
  data_stage_3__6512_,data_stage_3__6511_,data_stage_3__6510_,data_stage_3__6509_,
  data_stage_3__6508_,data_stage_3__6507_,data_stage_3__6506_,data_stage_3__6505_,
  data_stage_3__6504_,data_stage_3__6503_,data_stage_3__6502_,data_stage_3__6501_,
  data_stage_3__6500_,data_stage_3__6499_,data_stage_3__6498_,data_stage_3__6497_,
  data_stage_3__6496_,data_stage_3__6495_,data_stage_3__6494_,data_stage_3__6493_,
  data_stage_3__6492_,data_stage_3__6491_,data_stage_3__6490_,data_stage_3__6489_,
  data_stage_3__6488_,data_stage_3__6487_,data_stage_3__6486_,data_stage_3__6485_,
  data_stage_3__6484_,data_stage_3__6483_,data_stage_3__6482_,data_stage_3__6481_,
  data_stage_3__6480_,data_stage_3__6479_,data_stage_3__6478_,data_stage_3__6477_,
  data_stage_3__6476_,data_stage_3__6475_,data_stage_3__6474_,data_stage_3__6473_,
  data_stage_3__6472_,data_stage_3__6471_,data_stage_3__6470_,data_stage_3__6469_,
  data_stage_3__6468_,data_stage_3__6467_,data_stage_3__6466_,data_stage_3__6465_,
  data_stage_3__6464_,data_stage_3__6463_,data_stage_3__6462_,data_stage_3__6461_,
  data_stage_3__6460_,data_stage_3__6459_,data_stage_3__6458_,data_stage_3__6457_,
  data_stage_3__6456_,data_stage_3__6455_,data_stage_3__6454_,data_stage_3__6453_,
  data_stage_3__6452_,data_stage_3__6451_,data_stage_3__6450_,data_stage_3__6449_,
  data_stage_3__6448_,data_stage_3__6447_,data_stage_3__6446_,data_stage_3__6445_,
  data_stage_3__6444_,data_stage_3__6443_,data_stage_3__6442_,data_stage_3__6441_,
  data_stage_3__6440_,data_stage_3__6439_,data_stage_3__6438_,data_stage_3__6437_,
  data_stage_3__6436_,data_stage_3__6435_,data_stage_3__6434_,data_stage_3__6433_,
  data_stage_3__6432_,data_stage_3__6431_,data_stage_3__6430_,data_stage_3__6429_,
  data_stage_3__6428_,data_stage_3__6427_,data_stage_3__6426_,data_stage_3__6425_,
  data_stage_3__6424_,data_stage_3__6423_,data_stage_3__6422_,data_stage_3__6421_,
  data_stage_3__6420_,data_stage_3__6419_,data_stage_3__6418_,data_stage_3__6417_,
  data_stage_3__6416_,data_stage_3__6415_,data_stage_3__6414_,data_stage_3__6413_,
  data_stage_3__6412_,data_stage_3__6411_,data_stage_3__6410_,data_stage_3__6409_,
  data_stage_3__6408_,data_stage_3__6407_,data_stage_3__6406_,data_stage_3__6405_,
  data_stage_3__6404_,data_stage_3__6403_,data_stage_3__6402_,data_stage_3__6401_,
  data_stage_3__6400_,data_stage_3__6399_,data_stage_3__6398_,data_stage_3__6397_,
  data_stage_3__6396_,data_stage_3__6395_,data_stage_3__6394_,data_stage_3__6393_,
  data_stage_3__6392_,data_stage_3__6391_,data_stage_3__6390_,data_stage_3__6389_,
  data_stage_3__6388_,data_stage_3__6387_,data_stage_3__6386_,data_stage_3__6385_,
  data_stage_3__6384_,data_stage_3__6383_,data_stage_3__6382_,data_stage_3__6381_,
  data_stage_3__6380_,data_stage_3__6379_,data_stage_3__6378_,data_stage_3__6377_,
  data_stage_3__6376_,data_stage_3__6375_,data_stage_3__6374_,data_stage_3__6373_,
  data_stage_3__6372_,data_stage_3__6371_,data_stage_3__6370_,data_stage_3__6369_,
  data_stage_3__6368_,data_stage_3__6367_,data_stage_3__6366_,data_stage_3__6365_,
  data_stage_3__6364_,data_stage_3__6363_,data_stage_3__6362_,data_stage_3__6361_,
  data_stage_3__6360_,data_stage_3__6359_,data_stage_3__6358_,data_stage_3__6357_,
  data_stage_3__6356_,data_stage_3__6355_,data_stage_3__6354_,data_stage_3__6353_,
  data_stage_3__6352_,data_stage_3__6351_,data_stage_3__6350_,data_stage_3__6349_,
  data_stage_3__6348_,data_stage_3__6347_,data_stage_3__6346_,data_stage_3__6345_,
  data_stage_3__6344_,data_stage_3__6343_,data_stage_3__6342_,data_stage_3__6341_,
  data_stage_3__6340_,data_stage_3__6339_,data_stage_3__6338_,data_stage_3__6337_,
  data_stage_3__6336_,data_stage_3__6335_,data_stage_3__6334_,data_stage_3__6333_,
  data_stage_3__6332_,data_stage_3__6331_,data_stage_3__6330_,data_stage_3__6329_,
  data_stage_3__6328_,data_stage_3__6327_,data_stage_3__6326_,data_stage_3__6325_,
  data_stage_3__6324_,data_stage_3__6323_,data_stage_3__6322_,data_stage_3__6321_,
  data_stage_3__6320_,data_stage_3__6319_,data_stage_3__6318_,data_stage_3__6317_,
  data_stage_3__6316_,data_stage_3__6315_,data_stage_3__6314_,data_stage_3__6313_,
  data_stage_3__6312_,data_stage_3__6311_,data_stage_3__6310_,data_stage_3__6309_,
  data_stage_3__6308_,data_stage_3__6307_,data_stage_3__6306_,data_stage_3__6305_,
  data_stage_3__6304_,data_stage_3__6303_,data_stage_3__6302_,data_stage_3__6301_,
  data_stage_3__6300_,data_stage_3__6299_,data_stage_3__6298_,data_stage_3__6297_,
  data_stage_3__6296_,data_stage_3__6295_,data_stage_3__6294_,data_stage_3__6293_,
  data_stage_3__6292_,data_stage_3__6291_,data_stage_3__6290_,data_stage_3__6289_,
  data_stage_3__6288_,data_stage_3__6287_,data_stage_3__6286_,data_stage_3__6285_,
  data_stage_3__6284_,data_stage_3__6283_,data_stage_3__6282_,data_stage_3__6281_,
  data_stage_3__6280_,data_stage_3__6279_,data_stage_3__6278_,data_stage_3__6277_,
  data_stage_3__6276_,data_stage_3__6275_,data_stage_3__6274_,data_stage_3__6273_,
  data_stage_3__6272_,data_stage_3__6271_,data_stage_3__6270_,data_stage_3__6269_,
  data_stage_3__6268_,data_stage_3__6267_,data_stage_3__6266_,data_stage_3__6265_,
  data_stage_3__6264_,data_stage_3__6263_,data_stage_3__6262_,data_stage_3__6261_,
  data_stage_3__6260_,data_stage_3__6259_,data_stage_3__6258_,data_stage_3__6257_,
  data_stage_3__6256_,data_stage_3__6255_,data_stage_3__6254_,data_stage_3__6253_,
  data_stage_3__6252_,data_stage_3__6251_,data_stage_3__6250_,data_stage_3__6249_,
  data_stage_3__6248_,data_stage_3__6247_,data_stage_3__6246_,data_stage_3__6245_,
  data_stage_3__6244_,data_stage_3__6243_,data_stage_3__6242_,data_stage_3__6241_,
  data_stage_3__6240_,data_stage_3__6239_,data_stage_3__6238_,data_stage_3__6237_,
  data_stage_3__6236_,data_stage_3__6235_,data_stage_3__6234_,data_stage_3__6233_,
  data_stage_3__6232_,data_stage_3__6231_,data_stage_3__6230_,data_stage_3__6229_,
  data_stage_3__6228_,data_stage_3__6227_,data_stage_3__6226_,data_stage_3__6225_,
  data_stage_3__6224_,data_stage_3__6223_,data_stage_3__6222_,data_stage_3__6221_,
  data_stage_3__6220_,data_stage_3__6219_,data_stage_3__6218_,data_stage_3__6217_,
  data_stage_3__6216_,data_stage_3__6215_,data_stage_3__6214_,data_stage_3__6213_,
  data_stage_3__6212_,data_stage_3__6211_,data_stage_3__6210_,data_stage_3__6209_,
  data_stage_3__6208_,data_stage_3__6207_,data_stage_3__6206_,data_stage_3__6205_,
  data_stage_3__6204_,data_stage_3__6203_,data_stage_3__6202_,data_stage_3__6201_,
  data_stage_3__6200_,data_stage_3__6199_,data_stage_3__6198_,data_stage_3__6197_,
  data_stage_3__6196_,data_stage_3__6195_,data_stage_3__6194_,data_stage_3__6193_,
  data_stage_3__6192_,data_stage_3__6191_,data_stage_3__6190_,data_stage_3__6189_,
  data_stage_3__6188_,data_stage_3__6187_,data_stage_3__6186_,data_stage_3__6185_,
  data_stage_3__6184_,data_stage_3__6183_,data_stage_3__6182_,data_stage_3__6181_,
  data_stage_3__6180_,data_stage_3__6179_,data_stage_3__6178_,data_stage_3__6177_,
  data_stage_3__6176_,data_stage_3__6175_,data_stage_3__6174_,data_stage_3__6173_,
  data_stage_3__6172_,data_stage_3__6171_,data_stage_3__6170_,data_stage_3__6169_,
  data_stage_3__6168_,data_stage_3__6167_,data_stage_3__6166_,data_stage_3__6165_,
  data_stage_3__6164_,data_stage_3__6163_,data_stage_3__6162_,data_stage_3__6161_,
  data_stage_3__6160_,data_stage_3__6159_,data_stage_3__6158_,data_stage_3__6157_,
  data_stage_3__6156_,data_stage_3__6155_,data_stage_3__6154_,data_stage_3__6153_,
  data_stage_3__6152_,data_stage_3__6151_,data_stage_3__6150_,data_stage_3__6149_,
  data_stage_3__6148_,data_stage_3__6147_,data_stage_3__6146_,data_stage_3__6145_,
  data_stage_3__6144_,data_stage_3__6143_,data_stage_3__6142_,data_stage_3__6141_,
  data_stage_3__6140_,data_stage_3__6139_,data_stage_3__6138_,data_stage_3__6137_,
  data_stage_3__6136_,data_stage_3__6135_,data_stage_3__6134_,data_stage_3__6133_,
  data_stage_3__6132_,data_stage_3__6131_,data_stage_3__6130_,data_stage_3__6129_,
  data_stage_3__6128_,data_stage_3__6127_,data_stage_3__6126_,data_stage_3__6125_,
  data_stage_3__6124_,data_stage_3__6123_,data_stage_3__6122_,data_stage_3__6121_,
  data_stage_3__6120_,data_stage_3__6119_,data_stage_3__6118_,data_stage_3__6117_,
  data_stage_3__6116_,data_stage_3__6115_,data_stage_3__6114_,data_stage_3__6113_,
  data_stage_3__6112_,data_stage_3__6111_,data_stage_3__6110_,data_stage_3__6109_,
  data_stage_3__6108_,data_stage_3__6107_,data_stage_3__6106_,data_stage_3__6105_,
  data_stage_3__6104_,data_stage_3__6103_,data_stage_3__6102_,data_stage_3__6101_,
  data_stage_3__6100_,data_stage_3__6099_,data_stage_3__6098_,data_stage_3__6097_,
  data_stage_3__6096_,data_stage_3__6095_,data_stage_3__6094_,data_stage_3__6093_,
  data_stage_3__6092_,data_stage_3__6091_,data_stage_3__6090_,data_stage_3__6089_,
  data_stage_3__6088_,data_stage_3__6087_,data_stage_3__6086_,data_stage_3__6085_,
  data_stage_3__6084_,data_stage_3__6083_,data_stage_3__6082_,data_stage_3__6081_,
  data_stage_3__6080_,data_stage_3__6079_,data_stage_3__6078_,data_stage_3__6077_,
  data_stage_3__6076_,data_stage_3__6075_,data_stage_3__6074_,data_stage_3__6073_,
  data_stage_3__6072_,data_stage_3__6071_,data_stage_3__6070_,data_stage_3__6069_,
  data_stage_3__6068_,data_stage_3__6067_,data_stage_3__6066_,data_stage_3__6065_,
  data_stage_3__6064_,data_stage_3__6063_,data_stage_3__6062_,data_stage_3__6061_,
  data_stage_3__6060_,data_stage_3__6059_,data_stage_3__6058_,data_stage_3__6057_,
  data_stage_3__6056_,data_stage_3__6055_,data_stage_3__6054_,data_stage_3__6053_,
  data_stage_3__6052_,data_stage_3__6051_,data_stage_3__6050_,data_stage_3__6049_,
  data_stage_3__6048_,data_stage_3__6047_,data_stage_3__6046_,data_stage_3__6045_,
  data_stage_3__6044_,data_stage_3__6043_,data_stage_3__6042_,data_stage_3__6041_,
  data_stage_3__6040_,data_stage_3__6039_,data_stage_3__6038_,data_stage_3__6037_,
  data_stage_3__6036_,data_stage_3__6035_,data_stage_3__6034_,data_stage_3__6033_,
  data_stage_3__6032_,data_stage_3__6031_,data_stage_3__6030_,data_stage_3__6029_,
  data_stage_3__6028_,data_stage_3__6027_,data_stage_3__6026_,data_stage_3__6025_,
  data_stage_3__6024_,data_stage_3__6023_,data_stage_3__6022_,data_stage_3__6021_,
  data_stage_3__6020_,data_stage_3__6019_,data_stage_3__6018_,data_stage_3__6017_,
  data_stage_3__6016_,data_stage_3__6015_,data_stage_3__6014_,data_stage_3__6013_,
  data_stage_3__6012_,data_stage_3__6011_,data_stage_3__6010_,data_stage_3__6009_,
  data_stage_3__6008_,data_stage_3__6007_,data_stage_3__6006_,data_stage_3__6005_,
  data_stage_3__6004_,data_stage_3__6003_,data_stage_3__6002_,data_stage_3__6001_,
  data_stage_3__6000_,data_stage_3__5999_,data_stage_3__5998_,data_stage_3__5997_,
  data_stage_3__5996_,data_stage_3__5995_,data_stage_3__5994_,data_stage_3__5993_,
  data_stage_3__5992_,data_stage_3__5991_,data_stage_3__5990_,data_stage_3__5989_,
  data_stage_3__5988_,data_stage_3__5987_,data_stage_3__5986_,data_stage_3__5985_,
  data_stage_3__5984_,data_stage_3__5983_,data_stage_3__5982_,data_stage_3__5981_,
  data_stage_3__5980_,data_stage_3__5979_,data_stage_3__5978_,data_stage_3__5977_,
  data_stage_3__5976_,data_stage_3__5975_,data_stage_3__5974_,data_stage_3__5973_,
  data_stage_3__5972_,data_stage_3__5971_,data_stage_3__5970_,data_stage_3__5969_,
  data_stage_3__5968_,data_stage_3__5967_,data_stage_3__5966_,data_stage_3__5965_,
  data_stage_3__5964_,data_stage_3__5963_,data_stage_3__5962_,data_stage_3__5961_,
  data_stage_3__5960_,data_stage_3__5959_,data_stage_3__5958_,data_stage_3__5957_,
  data_stage_3__5956_,data_stage_3__5955_,data_stage_3__5954_,data_stage_3__5953_,
  data_stage_3__5952_,data_stage_3__5951_,data_stage_3__5950_,data_stage_3__5949_,
  data_stage_3__5948_,data_stage_3__5947_,data_stage_3__5946_,data_stage_3__5945_,
  data_stage_3__5944_,data_stage_3__5943_,data_stage_3__5942_,data_stage_3__5941_,
  data_stage_3__5940_,data_stage_3__5939_,data_stage_3__5938_,data_stage_3__5937_,
  data_stage_3__5936_,data_stage_3__5935_,data_stage_3__5934_,data_stage_3__5933_,
  data_stage_3__5932_,data_stage_3__5931_,data_stage_3__5930_,data_stage_3__5929_,
  data_stage_3__5928_,data_stage_3__5927_,data_stage_3__5926_,data_stage_3__5925_,
  data_stage_3__5924_,data_stage_3__5923_,data_stage_3__5922_,data_stage_3__5921_,
  data_stage_3__5920_,data_stage_3__5919_,data_stage_3__5918_,data_stage_3__5917_,
  data_stage_3__5916_,data_stage_3__5915_,data_stage_3__5914_,data_stage_3__5913_,
  data_stage_3__5912_,data_stage_3__5911_,data_stage_3__5910_,data_stage_3__5909_,
  data_stage_3__5908_,data_stage_3__5907_,data_stage_3__5906_,data_stage_3__5905_,
  data_stage_3__5904_,data_stage_3__5903_,data_stage_3__5902_,data_stage_3__5901_,
  data_stage_3__5900_,data_stage_3__5899_,data_stage_3__5898_,data_stage_3__5897_,
  data_stage_3__5896_,data_stage_3__5895_,data_stage_3__5894_,data_stage_3__5893_,
  data_stage_3__5892_,data_stage_3__5891_,data_stage_3__5890_,data_stage_3__5889_,
  data_stage_3__5888_,data_stage_3__5887_,data_stage_3__5886_,data_stage_3__5885_,
  data_stage_3__5884_,data_stage_3__5883_,data_stage_3__5882_,data_stage_3__5881_,
  data_stage_3__5880_,data_stage_3__5879_,data_stage_3__5878_,data_stage_3__5877_,
  data_stage_3__5876_,data_stage_3__5875_,data_stage_3__5874_,data_stage_3__5873_,
  data_stage_3__5872_,data_stage_3__5871_,data_stage_3__5870_,data_stage_3__5869_,
  data_stage_3__5868_,data_stage_3__5867_,data_stage_3__5866_,data_stage_3__5865_,
  data_stage_3__5864_,data_stage_3__5863_,data_stage_3__5862_,data_stage_3__5861_,
  data_stage_3__5860_,data_stage_3__5859_,data_stage_3__5858_,data_stage_3__5857_,
  data_stage_3__5856_,data_stage_3__5855_,data_stage_3__5854_,data_stage_3__5853_,
  data_stage_3__5852_,data_stage_3__5851_,data_stage_3__5850_,data_stage_3__5849_,
  data_stage_3__5848_,data_stage_3__5847_,data_stage_3__5846_,data_stage_3__5845_,
  data_stage_3__5844_,data_stage_3__5843_,data_stage_3__5842_,data_stage_3__5841_,
  data_stage_3__5840_,data_stage_3__5839_,data_stage_3__5838_,data_stage_3__5837_,
  data_stage_3__5836_,data_stage_3__5835_,data_stage_3__5834_,data_stage_3__5833_,
  data_stage_3__5832_,data_stage_3__5831_,data_stage_3__5830_,data_stage_3__5829_,
  data_stage_3__5828_,data_stage_3__5827_,data_stage_3__5826_,data_stage_3__5825_,
  data_stage_3__5824_,data_stage_3__5823_,data_stage_3__5822_,data_stage_3__5821_,
  data_stage_3__5820_,data_stage_3__5819_,data_stage_3__5818_,data_stage_3__5817_,
  data_stage_3__5816_,data_stage_3__5815_,data_stage_3__5814_,data_stage_3__5813_,
  data_stage_3__5812_,data_stage_3__5811_,data_stage_3__5810_,data_stage_3__5809_,
  data_stage_3__5808_,data_stage_3__5807_,data_stage_3__5806_,data_stage_3__5805_,
  data_stage_3__5804_,data_stage_3__5803_,data_stage_3__5802_,data_stage_3__5801_,
  data_stage_3__5800_,data_stage_3__5799_,data_stage_3__5798_,data_stage_3__5797_,
  data_stage_3__5796_,data_stage_3__5795_,data_stage_3__5794_,data_stage_3__5793_,
  data_stage_3__5792_,data_stage_3__5791_,data_stage_3__5790_,data_stage_3__5789_,
  data_stage_3__5788_,data_stage_3__5787_,data_stage_3__5786_,data_stage_3__5785_,
  data_stage_3__5784_,data_stage_3__5783_,data_stage_3__5782_,data_stage_3__5781_,
  data_stage_3__5780_,data_stage_3__5779_,data_stage_3__5778_,data_stage_3__5777_,
  data_stage_3__5776_,data_stage_3__5775_,data_stage_3__5774_,data_stage_3__5773_,
  data_stage_3__5772_,data_stage_3__5771_,data_stage_3__5770_,data_stage_3__5769_,
  data_stage_3__5768_,data_stage_3__5767_,data_stage_3__5766_,data_stage_3__5765_,
  data_stage_3__5764_,data_stage_3__5763_,data_stage_3__5762_,data_stage_3__5761_,
  data_stage_3__5760_,data_stage_3__5759_,data_stage_3__5758_,data_stage_3__5757_,
  data_stage_3__5756_,data_stage_3__5755_,data_stage_3__5754_,data_stage_3__5753_,
  data_stage_3__5752_,data_stage_3__5751_,data_stage_3__5750_,data_stage_3__5749_,
  data_stage_3__5748_,data_stage_3__5747_,data_stage_3__5746_,data_stage_3__5745_,
  data_stage_3__5744_,data_stage_3__5743_,data_stage_3__5742_,data_stage_3__5741_,
  data_stage_3__5740_,data_stage_3__5739_,data_stage_3__5738_,data_stage_3__5737_,
  data_stage_3__5736_,data_stage_3__5735_,data_stage_3__5734_,data_stage_3__5733_,
  data_stage_3__5732_,data_stage_3__5731_,data_stage_3__5730_,data_stage_3__5729_,
  data_stage_3__5728_,data_stage_3__5727_,data_stage_3__5726_,data_stage_3__5725_,
  data_stage_3__5724_,data_stage_3__5723_,data_stage_3__5722_,data_stage_3__5721_,
  data_stage_3__5720_,data_stage_3__5719_,data_stage_3__5718_,data_stage_3__5717_,
  data_stage_3__5716_,data_stage_3__5715_,data_stage_3__5714_,data_stage_3__5713_,
  data_stage_3__5712_,data_stage_3__5711_,data_stage_3__5710_,data_stage_3__5709_,
  data_stage_3__5708_,data_stage_3__5707_,data_stage_3__5706_,data_stage_3__5705_,
  data_stage_3__5704_,data_stage_3__5703_,data_stage_3__5702_,data_stage_3__5701_,
  data_stage_3__5700_,data_stage_3__5699_,data_stage_3__5698_,data_stage_3__5697_,
  data_stage_3__5696_,data_stage_3__5695_,data_stage_3__5694_,data_stage_3__5693_,
  data_stage_3__5692_,data_stage_3__5691_,data_stage_3__5690_,data_stage_3__5689_,
  data_stage_3__5688_,data_stage_3__5687_,data_stage_3__5686_,data_stage_3__5685_,
  data_stage_3__5684_,data_stage_3__5683_,data_stage_3__5682_,data_stage_3__5681_,
  data_stage_3__5680_,data_stage_3__5679_,data_stage_3__5678_,data_stage_3__5677_,
  data_stage_3__5676_,data_stage_3__5675_,data_stage_3__5674_,data_stage_3__5673_,
  data_stage_3__5672_,data_stage_3__5671_,data_stage_3__5670_,data_stage_3__5669_,
  data_stage_3__5668_,data_stage_3__5667_,data_stage_3__5666_,data_stage_3__5665_,
  data_stage_3__5664_,data_stage_3__5663_,data_stage_3__5662_,data_stage_3__5661_,
  data_stage_3__5660_,data_stage_3__5659_,data_stage_3__5658_,data_stage_3__5657_,
  data_stage_3__5656_,data_stage_3__5655_,data_stage_3__5654_,data_stage_3__5653_,
  data_stage_3__5652_,data_stage_3__5651_,data_stage_3__5650_,data_stage_3__5649_,
  data_stage_3__5648_,data_stage_3__5647_,data_stage_3__5646_,data_stage_3__5645_,
  data_stage_3__5644_,data_stage_3__5643_,data_stage_3__5642_,data_stage_3__5641_,
  data_stage_3__5640_,data_stage_3__5639_,data_stage_3__5638_,data_stage_3__5637_,
  data_stage_3__5636_,data_stage_3__5635_,data_stage_3__5634_,data_stage_3__5633_,
  data_stage_3__5632_,data_stage_3__5631_,data_stage_3__5630_,data_stage_3__5629_,
  data_stage_3__5628_,data_stage_3__5627_,data_stage_3__5626_,data_stage_3__5625_,
  data_stage_3__5624_,data_stage_3__5623_,data_stage_3__5622_,data_stage_3__5621_,
  data_stage_3__5620_,data_stage_3__5619_,data_stage_3__5618_,data_stage_3__5617_,
  data_stage_3__5616_,data_stage_3__5615_,data_stage_3__5614_,data_stage_3__5613_,
  data_stage_3__5612_,data_stage_3__5611_,data_stage_3__5610_,data_stage_3__5609_,
  data_stage_3__5608_,data_stage_3__5607_,data_stage_3__5606_,data_stage_3__5605_,
  data_stage_3__5604_,data_stage_3__5603_,data_stage_3__5602_,data_stage_3__5601_,
  data_stage_3__5600_,data_stage_3__5599_,data_stage_3__5598_,data_stage_3__5597_,
  data_stage_3__5596_,data_stage_3__5595_,data_stage_3__5594_,data_stage_3__5593_,
  data_stage_3__5592_,data_stage_3__5591_,data_stage_3__5590_,data_stage_3__5589_,
  data_stage_3__5588_,data_stage_3__5587_,data_stage_3__5586_,data_stage_3__5585_,
  data_stage_3__5584_,data_stage_3__5583_,data_stage_3__5582_,data_stage_3__5581_,
  data_stage_3__5580_,data_stage_3__5579_,data_stage_3__5578_,data_stage_3__5577_,
  data_stage_3__5576_,data_stage_3__5575_,data_stage_3__5574_,data_stage_3__5573_,
  data_stage_3__5572_,data_stage_3__5571_,data_stage_3__5570_,data_stage_3__5569_,
  data_stage_3__5568_,data_stage_3__5567_,data_stage_3__5566_,data_stage_3__5565_,
  data_stage_3__5564_,data_stage_3__5563_,data_stage_3__5562_,data_stage_3__5561_,
  data_stage_3__5560_,data_stage_3__5559_,data_stage_3__5558_,data_stage_3__5557_,
  data_stage_3__5556_,data_stage_3__5555_,data_stage_3__5554_,data_stage_3__5553_,
  data_stage_3__5552_,data_stage_3__5551_,data_stage_3__5550_,data_stage_3__5549_,
  data_stage_3__5548_,data_stage_3__5547_,data_stage_3__5546_,data_stage_3__5545_,
  data_stage_3__5544_,data_stage_3__5543_,data_stage_3__5542_,data_stage_3__5541_,
  data_stage_3__5540_,data_stage_3__5539_,data_stage_3__5538_,data_stage_3__5537_,
  data_stage_3__5536_,data_stage_3__5535_,data_stage_3__5534_,data_stage_3__5533_,
  data_stage_3__5532_,data_stage_3__5531_,data_stage_3__5530_,data_stage_3__5529_,
  data_stage_3__5528_,data_stage_3__5527_,data_stage_3__5526_,data_stage_3__5525_,
  data_stage_3__5524_,data_stage_3__5523_,data_stage_3__5522_,data_stage_3__5521_,
  data_stage_3__5520_,data_stage_3__5519_,data_stage_3__5518_,data_stage_3__5517_,
  data_stage_3__5516_,data_stage_3__5515_,data_stage_3__5514_,data_stage_3__5513_,
  data_stage_3__5512_,data_stage_3__5511_,data_stage_3__5510_,data_stage_3__5509_,
  data_stage_3__5508_,data_stage_3__5507_,data_stage_3__5506_,data_stage_3__5505_,
  data_stage_3__5504_,data_stage_3__5503_,data_stage_3__5502_,data_stage_3__5501_,
  data_stage_3__5500_,data_stage_3__5499_,data_stage_3__5498_,data_stage_3__5497_,
  data_stage_3__5496_,data_stage_3__5495_,data_stage_3__5494_,data_stage_3__5493_,
  data_stage_3__5492_,data_stage_3__5491_,data_stage_3__5490_,data_stage_3__5489_,
  data_stage_3__5488_,data_stage_3__5487_,data_stage_3__5486_,data_stage_3__5485_,
  data_stage_3__5484_,data_stage_3__5483_,data_stage_3__5482_,data_stage_3__5481_,
  data_stage_3__5480_,data_stage_3__5479_,data_stage_3__5478_,data_stage_3__5477_,
  data_stage_3__5476_,data_stage_3__5475_,data_stage_3__5474_,data_stage_3__5473_,
  data_stage_3__5472_,data_stage_3__5471_,data_stage_3__5470_,data_stage_3__5469_,
  data_stage_3__5468_,data_stage_3__5467_,data_stage_3__5466_,data_stage_3__5465_,
  data_stage_3__5464_,data_stage_3__5463_,data_stage_3__5462_,data_stage_3__5461_,
  data_stage_3__5460_,data_stage_3__5459_,data_stage_3__5458_,data_stage_3__5457_,
  data_stage_3__5456_,data_stage_3__5455_,data_stage_3__5454_,data_stage_3__5453_,
  data_stage_3__5452_,data_stage_3__5451_,data_stage_3__5450_,data_stage_3__5449_,
  data_stage_3__5448_,data_stage_3__5447_,data_stage_3__5446_,data_stage_3__5445_,
  data_stage_3__5444_,data_stage_3__5443_,data_stage_3__5442_,data_stage_3__5441_,
  data_stage_3__5440_,data_stage_3__5439_,data_stage_3__5438_,data_stage_3__5437_,
  data_stage_3__5436_,data_stage_3__5435_,data_stage_3__5434_,data_stage_3__5433_,
  data_stage_3__5432_,data_stage_3__5431_,data_stage_3__5430_,data_stage_3__5429_,
  data_stage_3__5428_,data_stage_3__5427_,data_stage_3__5426_,data_stage_3__5425_,
  data_stage_3__5424_,data_stage_3__5423_,data_stage_3__5422_,data_stage_3__5421_,
  data_stage_3__5420_,data_stage_3__5419_,data_stage_3__5418_,data_stage_3__5417_,
  data_stage_3__5416_,data_stage_3__5415_,data_stage_3__5414_,data_stage_3__5413_,
  data_stage_3__5412_,data_stage_3__5411_,data_stage_3__5410_,data_stage_3__5409_,
  data_stage_3__5408_,data_stage_3__5407_,data_stage_3__5406_,data_stage_3__5405_,
  data_stage_3__5404_,data_stage_3__5403_,data_stage_3__5402_,data_stage_3__5401_,
  data_stage_3__5400_,data_stage_3__5399_,data_stage_3__5398_,data_stage_3__5397_,
  data_stage_3__5396_,data_stage_3__5395_,data_stage_3__5394_,data_stage_3__5393_,
  data_stage_3__5392_,data_stage_3__5391_,data_stage_3__5390_,data_stage_3__5389_,
  data_stage_3__5388_,data_stage_3__5387_,data_stage_3__5386_,data_stage_3__5385_,
  data_stage_3__5384_,data_stage_3__5383_,data_stage_3__5382_,data_stage_3__5381_,
  data_stage_3__5380_,data_stage_3__5379_,data_stage_3__5378_,data_stage_3__5377_,
  data_stage_3__5376_,data_stage_3__5375_,data_stage_3__5374_,data_stage_3__5373_,
  data_stage_3__5372_,data_stage_3__5371_,data_stage_3__5370_,data_stage_3__5369_,
  data_stage_3__5368_,data_stage_3__5367_,data_stage_3__5366_,data_stage_3__5365_,
  data_stage_3__5364_,data_stage_3__5363_,data_stage_3__5362_,data_stage_3__5361_,
  data_stage_3__5360_,data_stage_3__5359_,data_stage_3__5358_,data_stage_3__5357_,
  data_stage_3__5356_,data_stage_3__5355_,data_stage_3__5354_,data_stage_3__5353_,
  data_stage_3__5352_,data_stage_3__5351_,data_stage_3__5350_,data_stage_3__5349_,
  data_stage_3__5348_,data_stage_3__5347_,data_stage_3__5346_,data_stage_3__5345_,
  data_stage_3__5344_,data_stage_3__5343_,data_stage_3__5342_,data_stage_3__5341_,
  data_stage_3__5340_,data_stage_3__5339_,data_stage_3__5338_,data_stage_3__5337_,
  data_stage_3__5336_,data_stage_3__5335_,data_stage_3__5334_,data_stage_3__5333_,
  data_stage_3__5332_,data_stage_3__5331_,data_stage_3__5330_,data_stage_3__5329_,
  data_stage_3__5328_,data_stage_3__5327_,data_stage_3__5326_,data_stage_3__5325_,
  data_stage_3__5324_,data_stage_3__5323_,data_stage_3__5322_,data_stage_3__5321_,
  data_stage_3__5320_,data_stage_3__5319_,data_stage_3__5318_,data_stage_3__5317_,
  data_stage_3__5316_,data_stage_3__5315_,data_stage_3__5314_,data_stage_3__5313_,
  data_stage_3__5312_,data_stage_3__5311_,data_stage_3__5310_,data_stage_3__5309_,
  data_stage_3__5308_,data_stage_3__5307_,data_stage_3__5306_,data_stage_3__5305_,
  data_stage_3__5304_,data_stage_3__5303_,data_stage_3__5302_,data_stage_3__5301_,
  data_stage_3__5300_,data_stage_3__5299_,data_stage_3__5298_,data_stage_3__5297_,
  data_stage_3__5296_,data_stage_3__5295_,data_stage_3__5294_,data_stage_3__5293_,
  data_stage_3__5292_,data_stage_3__5291_,data_stage_3__5290_,data_stage_3__5289_,
  data_stage_3__5288_,data_stage_3__5287_,data_stage_3__5286_,data_stage_3__5285_,
  data_stage_3__5284_,data_stage_3__5283_,data_stage_3__5282_,data_stage_3__5281_,
  data_stage_3__5280_,data_stage_3__5279_,data_stage_3__5278_,data_stage_3__5277_,
  data_stage_3__5276_,data_stage_3__5275_,data_stage_3__5274_,data_stage_3__5273_,
  data_stage_3__5272_,data_stage_3__5271_,data_stage_3__5270_,data_stage_3__5269_,
  data_stage_3__5268_,data_stage_3__5267_,data_stage_3__5266_,data_stage_3__5265_,
  data_stage_3__5264_,data_stage_3__5263_,data_stage_3__5262_,data_stage_3__5261_,
  data_stage_3__5260_,data_stage_3__5259_,data_stage_3__5258_,data_stage_3__5257_,
  data_stage_3__5256_,data_stage_3__5255_,data_stage_3__5254_,data_stage_3__5253_,
  data_stage_3__5252_,data_stage_3__5251_,data_stage_3__5250_,data_stage_3__5249_,
  data_stage_3__5248_,data_stage_3__5247_,data_stage_3__5246_,data_stage_3__5245_,
  data_stage_3__5244_,data_stage_3__5243_,data_stage_3__5242_,data_stage_3__5241_,
  data_stage_3__5240_,data_stage_3__5239_,data_stage_3__5238_,data_stage_3__5237_,
  data_stage_3__5236_,data_stage_3__5235_,data_stage_3__5234_,data_stage_3__5233_,
  data_stage_3__5232_,data_stage_3__5231_,data_stage_3__5230_,data_stage_3__5229_,
  data_stage_3__5228_,data_stage_3__5227_,data_stage_3__5226_,data_stage_3__5225_,
  data_stage_3__5224_,data_stage_3__5223_,data_stage_3__5222_,data_stage_3__5221_,
  data_stage_3__5220_,data_stage_3__5219_,data_stage_3__5218_,data_stage_3__5217_,
  data_stage_3__5216_,data_stage_3__5215_,data_stage_3__5214_,data_stage_3__5213_,
  data_stage_3__5212_,data_stage_3__5211_,data_stage_3__5210_,data_stage_3__5209_,
  data_stage_3__5208_,data_stage_3__5207_,data_stage_3__5206_,data_stage_3__5205_,
  data_stage_3__5204_,data_stage_3__5203_,data_stage_3__5202_,data_stage_3__5201_,
  data_stage_3__5200_,data_stage_3__5199_,data_stage_3__5198_,data_stage_3__5197_,
  data_stage_3__5196_,data_stage_3__5195_,data_stage_3__5194_,data_stage_3__5193_,
  data_stage_3__5192_,data_stage_3__5191_,data_stage_3__5190_,data_stage_3__5189_,
  data_stage_3__5188_,data_stage_3__5187_,data_stage_3__5186_,data_stage_3__5185_,
  data_stage_3__5184_,data_stage_3__5183_,data_stage_3__5182_,data_stage_3__5181_,
  data_stage_3__5180_,data_stage_3__5179_,data_stage_3__5178_,data_stage_3__5177_,
  data_stage_3__5176_,data_stage_3__5175_,data_stage_3__5174_,data_stage_3__5173_,
  data_stage_3__5172_,data_stage_3__5171_,data_stage_3__5170_,data_stage_3__5169_,
  data_stage_3__5168_,data_stage_3__5167_,data_stage_3__5166_,data_stage_3__5165_,
  data_stage_3__5164_,data_stage_3__5163_,data_stage_3__5162_,data_stage_3__5161_,
  data_stage_3__5160_,data_stage_3__5159_,data_stage_3__5158_,data_stage_3__5157_,
  data_stage_3__5156_,data_stage_3__5155_,data_stage_3__5154_,data_stage_3__5153_,
  data_stage_3__5152_,data_stage_3__5151_,data_stage_3__5150_,data_stage_3__5149_,
  data_stage_3__5148_,data_stage_3__5147_,data_stage_3__5146_,data_stage_3__5145_,
  data_stage_3__5144_,data_stage_3__5143_,data_stage_3__5142_,data_stage_3__5141_,
  data_stage_3__5140_,data_stage_3__5139_,data_stage_3__5138_,data_stage_3__5137_,
  data_stage_3__5136_,data_stage_3__5135_,data_stage_3__5134_,data_stage_3__5133_,
  data_stage_3__5132_,data_stage_3__5131_,data_stage_3__5130_,data_stage_3__5129_,
  data_stage_3__5128_,data_stage_3__5127_,data_stage_3__5126_,data_stage_3__5125_,
  data_stage_3__5124_,data_stage_3__5123_,data_stage_3__5122_,data_stage_3__5121_,
  data_stage_3__5120_,data_stage_3__5119_,data_stage_3__5118_,data_stage_3__5117_,
  data_stage_3__5116_,data_stage_3__5115_,data_stage_3__5114_,data_stage_3__5113_,
  data_stage_3__5112_,data_stage_3__5111_,data_stage_3__5110_,data_stage_3__5109_,
  data_stage_3__5108_,data_stage_3__5107_,data_stage_3__5106_,data_stage_3__5105_,
  data_stage_3__5104_,data_stage_3__5103_,data_stage_3__5102_,data_stage_3__5101_,
  data_stage_3__5100_,data_stage_3__5099_,data_stage_3__5098_,data_stage_3__5097_,
  data_stage_3__5096_,data_stage_3__5095_,data_stage_3__5094_,data_stage_3__5093_,
  data_stage_3__5092_,data_stage_3__5091_,data_stage_3__5090_,data_stage_3__5089_,
  data_stage_3__5088_,data_stage_3__5087_,data_stage_3__5086_,data_stage_3__5085_,
  data_stage_3__5084_,data_stage_3__5083_,data_stage_3__5082_,data_stage_3__5081_,
  data_stage_3__5080_,data_stage_3__5079_,data_stage_3__5078_,data_stage_3__5077_,
  data_stage_3__5076_,data_stage_3__5075_,data_stage_3__5074_,data_stage_3__5073_,
  data_stage_3__5072_,data_stage_3__5071_,data_stage_3__5070_,data_stage_3__5069_,
  data_stage_3__5068_,data_stage_3__5067_,data_stage_3__5066_,data_stage_3__5065_,
  data_stage_3__5064_,data_stage_3__5063_,data_stage_3__5062_,data_stage_3__5061_,
  data_stage_3__5060_,data_stage_3__5059_,data_stage_3__5058_,data_stage_3__5057_,
  data_stage_3__5056_,data_stage_3__5055_,data_stage_3__5054_,data_stage_3__5053_,
  data_stage_3__5052_,data_stage_3__5051_,data_stage_3__5050_,data_stage_3__5049_,
  data_stage_3__5048_,data_stage_3__5047_,data_stage_3__5046_,data_stage_3__5045_,
  data_stage_3__5044_,data_stage_3__5043_,data_stage_3__5042_,data_stage_3__5041_,
  data_stage_3__5040_,data_stage_3__5039_,data_stage_3__5038_,data_stage_3__5037_,
  data_stage_3__5036_,data_stage_3__5035_,data_stage_3__5034_,data_stage_3__5033_,
  data_stage_3__5032_,data_stage_3__5031_,data_stage_3__5030_,data_stage_3__5029_,
  data_stage_3__5028_,data_stage_3__5027_,data_stage_3__5026_,data_stage_3__5025_,
  data_stage_3__5024_,data_stage_3__5023_,data_stage_3__5022_,data_stage_3__5021_,
  data_stage_3__5020_,data_stage_3__5019_,data_stage_3__5018_,data_stage_3__5017_,
  data_stage_3__5016_,data_stage_3__5015_,data_stage_3__5014_,data_stage_3__5013_,
  data_stage_3__5012_,data_stage_3__5011_,data_stage_3__5010_,data_stage_3__5009_,
  data_stage_3__5008_,data_stage_3__5007_,data_stage_3__5006_,data_stage_3__5005_,
  data_stage_3__5004_,data_stage_3__5003_,data_stage_3__5002_,data_stage_3__5001_,
  data_stage_3__5000_,data_stage_3__4999_,data_stage_3__4998_,data_stage_3__4997_,
  data_stage_3__4996_,data_stage_3__4995_,data_stage_3__4994_,data_stage_3__4993_,
  data_stage_3__4992_,data_stage_3__4991_,data_stage_3__4990_,data_stage_3__4989_,
  data_stage_3__4988_,data_stage_3__4987_,data_stage_3__4986_,data_stage_3__4985_,
  data_stage_3__4984_,data_stage_3__4983_,data_stage_3__4982_,data_stage_3__4981_,
  data_stage_3__4980_,data_stage_3__4979_,data_stage_3__4978_,data_stage_3__4977_,
  data_stage_3__4976_,data_stage_3__4975_,data_stage_3__4974_,data_stage_3__4973_,
  data_stage_3__4972_,data_stage_3__4971_,data_stage_3__4970_,data_stage_3__4969_,
  data_stage_3__4968_,data_stage_3__4967_,data_stage_3__4966_,data_stage_3__4965_,
  data_stage_3__4964_,data_stage_3__4963_,data_stage_3__4962_,data_stage_3__4961_,
  data_stage_3__4960_,data_stage_3__4959_,data_stage_3__4958_,data_stage_3__4957_,
  data_stage_3__4956_,data_stage_3__4955_,data_stage_3__4954_,data_stage_3__4953_,
  data_stage_3__4952_,data_stage_3__4951_,data_stage_3__4950_,data_stage_3__4949_,
  data_stage_3__4948_,data_stage_3__4947_,data_stage_3__4946_,data_stage_3__4945_,
  data_stage_3__4944_,data_stage_3__4943_,data_stage_3__4942_,data_stage_3__4941_,
  data_stage_3__4940_,data_stage_3__4939_,data_stage_3__4938_,data_stage_3__4937_,
  data_stage_3__4936_,data_stage_3__4935_,data_stage_3__4934_,data_stage_3__4933_,
  data_stage_3__4932_,data_stage_3__4931_,data_stage_3__4930_,data_stage_3__4929_,
  data_stage_3__4928_,data_stage_3__4927_,data_stage_3__4926_,data_stage_3__4925_,
  data_stage_3__4924_,data_stage_3__4923_,data_stage_3__4922_,data_stage_3__4921_,
  data_stage_3__4920_,data_stage_3__4919_,data_stage_3__4918_,data_stage_3__4917_,
  data_stage_3__4916_,data_stage_3__4915_,data_stage_3__4914_,data_stage_3__4913_,
  data_stage_3__4912_,data_stage_3__4911_,data_stage_3__4910_,data_stage_3__4909_,
  data_stage_3__4908_,data_stage_3__4907_,data_stage_3__4906_,data_stage_3__4905_,
  data_stage_3__4904_,data_stage_3__4903_,data_stage_3__4902_,data_stage_3__4901_,
  data_stage_3__4900_,data_stage_3__4899_,data_stage_3__4898_,data_stage_3__4897_,
  data_stage_3__4896_,data_stage_3__4895_,data_stage_3__4894_,data_stage_3__4893_,
  data_stage_3__4892_,data_stage_3__4891_,data_stage_3__4890_,data_stage_3__4889_,
  data_stage_3__4888_,data_stage_3__4887_,data_stage_3__4886_,data_stage_3__4885_,
  data_stage_3__4884_,data_stage_3__4883_,data_stage_3__4882_,data_stage_3__4881_,
  data_stage_3__4880_,data_stage_3__4879_,data_stage_3__4878_,data_stage_3__4877_,
  data_stage_3__4876_,data_stage_3__4875_,data_stage_3__4874_,data_stage_3__4873_,
  data_stage_3__4872_,data_stage_3__4871_,data_stage_3__4870_,data_stage_3__4869_,
  data_stage_3__4868_,data_stage_3__4867_,data_stage_3__4866_,data_stage_3__4865_,
  data_stage_3__4864_,data_stage_3__4863_,data_stage_3__4862_,data_stage_3__4861_,
  data_stage_3__4860_,data_stage_3__4859_,data_stage_3__4858_,data_stage_3__4857_,
  data_stage_3__4856_,data_stage_3__4855_,data_stage_3__4854_,data_stage_3__4853_,
  data_stage_3__4852_,data_stage_3__4851_,data_stage_3__4850_,data_stage_3__4849_,
  data_stage_3__4848_,data_stage_3__4847_,data_stage_3__4846_,data_stage_3__4845_,
  data_stage_3__4844_,data_stage_3__4843_,data_stage_3__4842_,data_stage_3__4841_,
  data_stage_3__4840_,data_stage_3__4839_,data_stage_3__4838_,data_stage_3__4837_,
  data_stage_3__4836_,data_stage_3__4835_,data_stage_3__4834_,data_stage_3__4833_,
  data_stage_3__4832_,data_stage_3__4831_,data_stage_3__4830_,data_stage_3__4829_,
  data_stage_3__4828_,data_stage_3__4827_,data_stage_3__4826_,data_stage_3__4825_,
  data_stage_3__4824_,data_stage_3__4823_,data_stage_3__4822_,data_stage_3__4821_,
  data_stage_3__4820_,data_stage_3__4819_,data_stage_3__4818_,data_stage_3__4817_,
  data_stage_3__4816_,data_stage_3__4815_,data_stage_3__4814_,data_stage_3__4813_,
  data_stage_3__4812_,data_stage_3__4811_,data_stage_3__4810_,data_stage_3__4809_,
  data_stage_3__4808_,data_stage_3__4807_,data_stage_3__4806_,data_stage_3__4805_,
  data_stage_3__4804_,data_stage_3__4803_,data_stage_3__4802_,data_stage_3__4801_,
  data_stage_3__4800_,data_stage_3__4799_,data_stage_3__4798_,data_stage_3__4797_,
  data_stage_3__4796_,data_stage_3__4795_,data_stage_3__4794_,data_stage_3__4793_,
  data_stage_3__4792_,data_stage_3__4791_,data_stage_3__4790_,data_stage_3__4789_,
  data_stage_3__4788_,data_stage_3__4787_,data_stage_3__4786_,data_stage_3__4785_,
  data_stage_3__4784_,data_stage_3__4783_,data_stage_3__4782_,data_stage_3__4781_,
  data_stage_3__4780_,data_stage_3__4779_,data_stage_3__4778_,data_stage_3__4777_,
  data_stage_3__4776_,data_stage_3__4775_,data_stage_3__4774_,data_stage_3__4773_,
  data_stage_3__4772_,data_stage_3__4771_,data_stage_3__4770_,data_stage_3__4769_,
  data_stage_3__4768_,data_stage_3__4767_,data_stage_3__4766_,data_stage_3__4765_,
  data_stage_3__4764_,data_stage_3__4763_,data_stage_3__4762_,data_stage_3__4761_,
  data_stage_3__4760_,data_stage_3__4759_,data_stage_3__4758_,data_stage_3__4757_,
  data_stage_3__4756_,data_stage_3__4755_,data_stage_3__4754_,data_stage_3__4753_,
  data_stage_3__4752_,data_stage_3__4751_,data_stage_3__4750_,data_stage_3__4749_,
  data_stage_3__4748_,data_stage_3__4747_,data_stage_3__4746_,data_stage_3__4745_,
  data_stage_3__4744_,data_stage_3__4743_,data_stage_3__4742_,data_stage_3__4741_,
  data_stage_3__4740_,data_stage_3__4739_,data_stage_3__4738_,data_stage_3__4737_,
  data_stage_3__4736_,data_stage_3__4735_,data_stage_3__4734_,data_stage_3__4733_,
  data_stage_3__4732_,data_stage_3__4731_,data_stage_3__4730_,data_stage_3__4729_,
  data_stage_3__4728_,data_stage_3__4727_,data_stage_3__4726_,data_stage_3__4725_,
  data_stage_3__4724_,data_stage_3__4723_,data_stage_3__4722_,data_stage_3__4721_,
  data_stage_3__4720_,data_stage_3__4719_,data_stage_3__4718_,data_stage_3__4717_,
  data_stage_3__4716_,data_stage_3__4715_,data_stage_3__4714_,data_stage_3__4713_,
  data_stage_3__4712_,data_stage_3__4711_,data_stage_3__4710_,data_stage_3__4709_,
  data_stage_3__4708_,data_stage_3__4707_,data_stage_3__4706_,data_stage_3__4705_,
  data_stage_3__4704_,data_stage_3__4703_,data_stage_3__4702_,data_stage_3__4701_,
  data_stage_3__4700_,data_stage_3__4699_,data_stage_3__4698_,data_stage_3__4697_,
  data_stage_3__4696_,data_stage_3__4695_,data_stage_3__4694_,data_stage_3__4693_,
  data_stage_3__4692_,data_stage_3__4691_,data_stage_3__4690_,data_stage_3__4689_,
  data_stage_3__4688_,data_stage_3__4687_,data_stage_3__4686_,data_stage_3__4685_,
  data_stage_3__4684_,data_stage_3__4683_,data_stage_3__4682_,data_stage_3__4681_,
  data_stage_3__4680_,data_stage_3__4679_,data_stage_3__4678_,data_stage_3__4677_,
  data_stage_3__4676_,data_stage_3__4675_,data_stage_3__4674_,data_stage_3__4673_,
  data_stage_3__4672_,data_stage_3__4671_,data_stage_3__4670_,data_stage_3__4669_,
  data_stage_3__4668_,data_stage_3__4667_,data_stage_3__4666_,data_stage_3__4665_,
  data_stage_3__4664_,data_stage_3__4663_,data_stage_3__4662_,data_stage_3__4661_,
  data_stage_3__4660_,data_stage_3__4659_,data_stage_3__4658_,data_stage_3__4657_,
  data_stage_3__4656_,data_stage_3__4655_,data_stage_3__4654_,data_stage_3__4653_,
  data_stage_3__4652_,data_stage_3__4651_,data_stage_3__4650_,data_stage_3__4649_,
  data_stage_3__4648_,data_stage_3__4647_,data_stage_3__4646_,data_stage_3__4645_,
  data_stage_3__4644_,data_stage_3__4643_,data_stage_3__4642_,data_stage_3__4641_,
  data_stage_3__4640_,data_stage_3__4639_,data_stage_3__4638_,data_stage_3__4637_,
  data_stage_3__4636_,data_stage_3__4635_,data_stage_3__4634_,data_stage_3__4633_,
  data_stage_3__4632_,data_stage_3__4631_,data_stage_3__4630_,data_stage_3__4629_,
  data_stage_3__4628_,data_stage_3__4627_,data_stage_3__4626_,data_stage_3__4625_,
  data_stage_3__4624_,data_stage_3__4623_,data_stage_3__4622_,data_stage_3__4621_,
  data_stage_3__4620_,data_stage_3__4619_,data_stage_3__4618_,data_stage_3__4617_,
  data_stage_3__4616_,data_stage_3__4615_,data_stage_3__4614_,data_stage_3__4613_,
  data_stage_3__4612_,data_stage_3__4611_,data_stage_3__4610_,data_stage_3__4609_,
  data_stage_3__4608_,data_stage_3__4607_,data_stage_3__4606_,data_stage_3__4605_,
  data_stage_3__4604_,data_stage_3__4603_,data_stage_3__4602_,data_stage_3__4601_,
  data_stage_3__4600_,data_stage_3__4599_,data_stage_3__4598_,data_stage_3__4597_,
  data_stage_3__4596_,data_stage_3__4595_,data_stage_3__4594_,data_stage_3__4593_,
  data_stage_3__4592_,data_stage_3__4591_,data_stage_3__4590_,data_stage_3__4589_,
  data_stage_3__4588_,data_stage_3__4587_,data_stage_3__4586_,data_stage_3__4585_,
  data_stage_3__4584_,data_stage_3__4583_,data_stage_3__4582_,data_stage_3__4581_,
  data_stage_3__4580_,data_stage_3__4579_,data_stage_3__4578_,data_stage_3__4577_,
  data_stage_3__4576_,data_stage_3__4575_,data_stage_3__4574_,data_stage_3__4573_,
  data_stage_3__4572_,data_stage_3__4571_,data_stage_3__4570_,data_stage_3__4569_,
  data_stage_3__4568_,data_stage_3__4567_,data_stage_3__4566_,data_stage_3__4565_,
  data_stage_3__4564_,data_stage_3__4563_,data_stage_3__4562_,data_stage_3__4561_,
  data_stage_3__4560_,data_stage_3__4559_,data_stage_3__4558_,data_stage_3__4557_,
  data_stage_3__4556_,data_stage_3__4555_,data_stage_3__4554_,data_stage_3__4553_,
  data_stage_3__4552_,data_stage_3__4551_,data_stage_3__4550_,data_stage_3__4549_,
  data_stage_3__4548_,data_stage_3__4547_,data_stage_3__4546_,data_stage_3__4545_,
  data_stage_3__4544_,data_stage_3__4543_,data_stage_3__4542_,data_stage_3__4541_,
  data_stage_3__4540_,data_stage_3__4539_,data_stage_3__4538_,data_stage_3__4537_,
  data_stage_3__4536_,data_stage_3__4535_,data_stage_3__4534_,data_stage_3__4533_,
  data_stage_3__4532_,data_stage_3__4531_,data_stage_3__4530_,data_stage_3__4529_,
  data_stage_3__4528_,data_stage_3__4527_,data_stage_3__4526_,data_stage_3__4525_,
  data_stage_3__4524_,data_stage_3__4523_,data_stage_3__4522_,data_stage_3__4521_,
  data_stage_3__4520_,data_stage_3__4519_,data_stage_3__4518_,data_stage_3__4517_,
  data_stage_3__4516_,data_stage_3__4515_,data_stage_3__4514_,data_stage_3__4513_,
  data_stage_3__4512_,data_stage_3__4511_,data_stage_3__4510_,data_stage_3__4509_,
  data_stage_3__4508_,data_stage_3__4507_,data_stage_3__4506_,data_stage_3__4505_,
  data_stage_3__4504_,data_stage_3__4503_,data_stage_3__4502_,data_stage_3__4501_,
  data_stage_3__4500_,data_stage_3__4499_,data_stage_3__4498_,data_stage_3__4497_,
  data_stage_3__4496_,data_stage_3__4495_,data_stage_3__4494_,data_stage_3__4493_,
  data_stage_3__4492_,data_stage_3__4491_,data_stage_3__4490_,data_stage_3__4489_,
  data_stage_3__4488_,data_stage_3__4487_,data_stage_3__4486_,data_stage_3__4485_,
  data_stage_3__4484_,data_stage_3__4483_,data_stage_3__4482_,data_stage_3__4481_,
  data_stage_3__4480_,data_stage_3__4479_,data_stage_3__4478_,data_stage_3__4477_,
  data_stage_3__4476_,data_stage_3__4475_,data_stage_3__4474_,data_stage_3__4473_,
  data_stage_3__4472_,data_stage_3__4471_,data_stage_3__4470_,data_stage_3__4469_,
  data_stage_3__4468_,data_stage_3__4467_,data_stage_3__4466_,data_stage_3__4465_,
  data_stage_3__4464_,data_stage_3__4463_,data_stage_3__4462_,data_stage_3__4461_,
  data_stage_3__4460_,data_stage_3__4459_,data_stage_3__4458_,data_stage_3__4457_,
  data_stage_3__4456_,data_stage_3__4455_,data_stage_3__4454_,data_stage_3__4453_,
  data_stage_3__4452_,data_stage_3__4451_,data_stage_3__4450_,data_stage_3__4449_,
  data_stage_3__4448_,data_stage_3__4447_,data_stage_3__4446_,data_stage_3__4445_,
  data_stage_3__4444_,data_stage_3__4443_,data_stage_3__4442_,data_stage_3__4441_,
  data_stage_3__4440_,data_stage_3__4439_,data_stage_3__4438_,data_stage_3__4437_,
  data_stage_3__4436_,data_stage_3__4435_,data_stage_3__4434_,data_stage_3__4433_,
  data_stage_3__4432_,data_stage_3__4431_,data_stage_3__4430_,data_stage_3__4429_,
  data_stage_3__4428_,data_stage_3__4427_,data_stage_3__4426_,data_stage_3__4425_,
  data_stage_3__4424_,data_stage_3__4423_,data_stage_3__4422_,data_stage_3__4421_,
  data_stage_3__4420_,data_stage_3__4419_,data_stage_3__4418_,data_stage_3__4417_,
  data_stage_3__4416_,data_stage_3__4415_,data_stage_3__4414_,data_stage_3__4413_,
  data_stage_3__4412_,data_stage_3__4411_,data_stage_3__4410_,data_stage_3__4409_,
  data_stage_3__4408_,data_stage_3__4407_,data_stage_3__4406_,data_stage_3__4405_,
  data_stage_3__4404_,data_stage_3__4403_,data_stage_3__4402_,data_stage_3__4401_,
  data_stage_3__4400_,data_stage_3__4399_,data_stage_3__4398_,data_stage_3__4397_,
  data_stage_3__4396_,data_stage_3__4395_,data_stage_3__4394_,data_stage_3__4393_,
  data_stage_3__4392_,data_stage_3__4391_,data_stage_3__4390_,data_stage_3__4389_,
  data_stage_3__4388_,data_stage_3__4387_,data_stage_3__4386_,data_stage_3__4385_,
  data_stage_3__4384_,data_stage_3__4383_,data_stage_3__4382_,data_stage_3__4381_,
  data_stage_3__4380_,data_stage_3__4379_,data_stage_3__4378_,data_stage_3__4377_,
  data_stage_3__4376_,data_stage_3__4375_,data_stage_3__4374_,data_stage_3__4373_,
  data_stage_3__4372_,data_stage_3__4371_,data_stage_3__4370_,data_stage_3__4369_,
  data_stage_3__4368_,data_stage_3__4367_,data_stage_3__4366_,data_stage_3__4365_,
  data_stage_3__4364_,data_stage_3__4363_,data_stage_3__4362_,data_stage_3__4361_,
  data_stage_3__4360_,data_stage_3__4359_,data_stage_3__4358_,data_stage_3__4357_,
  data_stage_3__4356_,data_stage_3__4355_,data_stage_3__4354_,data_stage_3__4353_,
  data_stage_3__4352_,data_stage_3__4351_,data_stage_3__4350_,data_stage_3__4349_,
  data_stage_3__4348_,data_stage_3__4347_,data_stage_3__4346_,data_stage_3__4345_,
  data_stage_3__4344_,data_stage_3__4343_,data_stage_3__4342_,data_stage_3__4341_,
  data_stage_3__4340_,data_stage_3__4339_,data_stage_3__4338_,data_stage_3__4337_,
  data_stage_3__4336_,data_stage_3__4335_,data_stage_3__4334_,data_stage_3__4333_,
  data_stage_3__4332_,data_stage_3__4331_,data_stage_3__4330_,data_stage_3__4329_,
  data_stage_3__4328_,data_stage_3__4327_,data_stage_3__4326_,data_stage_3__4325_,
  data_stage_3__4324_,data_stage_3__4323_,data_stage_3__4322_,data_stage_3__4321_,
  data_stage_3__4320_,data_stage_3__4319_,data_stage_3__4318_,data_stage_3__4317_,
  data_stage_3__4316_,data_stage_3__4315_,data_stage_3__4314_,data_stage_3__4313_,
  data_stage_3__4312_,data_stage_3__4311_,data_stage_3__4310_,data_stage_3__4309_,
  data_stage_3__4308_,data_stage_3__4307_,data_stage_3__4306_,data_stage_3__4305_,
  data_stage_3__4304_,data_stage_3__4303_,data_stage_3__4302_,data_stage_3__4301_,
  data_stage_3__4300_,data_stage_3__4299_,data_stage_3__4298_,data_stage_3__4297_,
  data_stage_3__4296_,data_stage_3__4295_,data_stage_3__4294_,data_stage_3__4293_,
  data_stage_3__4292_,data_stage_3__4291_,data_stage_3__4290_,data_stage_3__4289_,
  data_stage_3__4288_,data_stage_3__4287_,data_stage_3__4286_,data_stage_3__4285_,
  data_stage_3__4284_,data_stage_3__4283_,data_stage_3__4282_,data_stage_3__4281_,
  data_stage_3__4280_,data_stage_3__4279_,data_stage_3__4278_,data_stage_3__4277_,
  data_stage_3__4276_,data_stage_3__4275_,data_stage_3__4274_,data_stage_3__4273_,
  data_stage_3__4272_,data_stage_3__4271_,data_stage_3__4270_,data_stage_3__4269_,
  data_stage_3__4268_,data_stage_3__4267_,data_stage_3__4266_,data_stage_3__4265_,
  data_stage_3__4264_,data_stage_3__4263_,data_stage_3__4262_,data_stage_3__4261_,
  data_stage_3__4260_,data_stage_3__4259_,data_stage_3__4258_,data_stage_3__4257_,
  data_stage_3__4256_,data_stage_3__4255_,data_stage_3__4254_,data_stage_3__4253_,
  data_stage_3__4252_,data_stage_3__4251_,data_stage_3__4250_,data_stage_3__4249_,
  data_stage_3__4248_,data_stage_3__4247_,data_stage_3__4246_,data_stage_3__4245_,
  data_stage_3__4244_,data_stage_3__4243_,data_stage_3__4242_,data_stage_3__4241_,
  data_stage_3__4240_,data_stage_3__4239_,data_stage_3__4238_,data_stage_3__4237_,
  data_stage_3__4236_,data_stage_3__4235_,data_stage_3__4234_,data_stage_3__4233_,
  data_stage_3__4232_,data_stage_3__4231_,data_stage_3__4230_,data_stage_3__4229_,
  data_stage_3__4228_,data_stage_3__4227_,data_stage_3__4226_,data_stage_3__4225_,
  data_stage_3__4224_,data_stage_3__4223_,data_stage_3__4222_,data_stage_3__4221_,
  data_stage_3__4220_,data_stage_3__4219_,data_stage_3__4218_,data_stage_3__4217_,
  data_stage_3__4216_,data_stage_3__4215_,data_stage_3__4214_,data_stage_3__4213_,
  data_stage_3__4212_,data_stage_3__4211_,data_stage_3__4210_,data_stage_3__4209_,
  data_stage_3__4208_,data_stage_3__4207_,data_stage_3__4206_,data_stage_3__4205_,
  data_stage_3__4204_,data_stage_3__4203_,data_stage_3__4202_,data_stage_3__4201_,
  data_stage_3__4200_,data_stage_3__4199_,data_stage_3__4198_,data_stage_3__4197_,
  data_stage_3__4196_,data_stage_3__4195_,data_stage_3__4194_,data_stage_3__4193_,
  data_stage_3__4192_,data_stage_3__4191_,data_stage_3__4190_,data_stage_3__4189_,
  data_stage_3__4188_,data_stage_3__4187_,data_stage_3__4186_,data_stage_3__4185_,
  data_stage_3__4184_,data_stage_3__4183_,data_stage_3__4182_,data_stage_3__4181_,
  data_stage_3__4180_,data_stage_3__4179_,data_stage_3__4178_,data_stage_3__4177_,
  data_stage_3__4176_,data_stage_3__4175_,data_stage_3__4174_,data_stage_3__4173_,
  data_stage_3__4172_,data_stage_3__4171_,data_stage_3__4170_,data_stage_3__4169_,
  data_stage_3__4168_,data_stage_3__4167_,data_stage_3__4166_,data_stage_3__4165_,
  data_stage_3__4164_,data_stage_3__4163_,data_stage_3__4162_,data_stage_3__4161_,
  data_stage_3__4160_,data_stage_3__4159_,data_stage_3__4158_,data_stage_3__4157_,
  data_stage_3__4156_,data_stage_3__4155_,data_stage_3__4154_,data_stage_3__4153_,
  data_stage_3__4152_,data_stage_3__4151_,data_stage_3__4150_,data_stage_3__4149_,
  data_stage_3__4148_,data_stage_3__4147_,data_stage_3__4146_,data_stage_3__4145_,
  data_stage_3__4144_,data_stage_3__4143_,data_stage_3__4142_,data_stage_3__4141_,
  data_stage_3__4140_,data_stage_3__4139_,data_stage_3__4138_,data_stage_3__4137_,
  data_stage_3__4136_,data_stage_3__4135_,data_stage_3__4134_,data_stage_3__4133_,
  data_stage_3__4132_,data_stage_3__4131_,data_stage_3__4130_,data_stage_3__4129_,
  data_stage_3__4128_,data_stage_3__4127_,data_stage_3__4126_,data_stage_3__4125_,
  data_stage_3__4124_,data_stage_3__4123_,data_stage_3__4122_,data_stage_3__4121_,
  data_stage_3__4120_,data_stage_3__4119_,data_stage_3__4118_,data_stage_3__4117_,
  data_stage_3__4116_,data_stage_3__4115_,data_stage_3__4114_,data_stage_3__4113_,
  data_stage_3__4112_,data_stage_3__4111_,data_stage_3__4110_,data_stage_3__4109_,
  data_stage_3__4108_,data_stage_3__4107_,data_stage_3__4106_,data_stage_3__4105_,
  data_stage_3__4104_,data_stage_3__4103_,data_stage_3__4102_,data_stage_3__4101_,
  data_stage_3__4100_,data_stage_3__4099_,data_stage_3__4098_,data_stage_3__4097_,
  data_stage_3__4096_,data_stage_3__4095_,data_stage_3__4094_,data_stage_3__4093_,
  data_stage_3__4092_,data_stage_3__4091_,data_stage_3__4090_,data_stage_3__4089_,
  data_stage_3__4088_,data_stage_3__4087_,data_stage_3__4086_,data_stage_3__4085_,
  data_stage_3__4084_,data_stage_3__4083_,data_stage_3__4082_,data_stage_3__4081_,
  data_stage_3__4080_,data_stage_3__4079_,data_stage_3__4078_,data_stage_3__4077_,
  data_stage_3__4076_,data_stage_3__4075_,data_stage_3__4074_,data_stage_3__4073_,
  data_stage_3__4072_,data_stage_3__4071_,data_stage_3__4070_,data_stage_3__4069_,
  data_stage_3__4068_,data_stage_3__4067_,data_stage_3__4066_,data_stage_3__4065_,
  data_stage_3__4064_,data_stage_3__4063_,data_stage_3__4062_,data_stage_3__4061_,
  data_stage_3__4060_,data_stage_3__4059_,data_stage_3__4058_,data_stage_3__4057_,
  data_stage_3__4056_,data_stage_3__4055_,data_stage_3__4054_,data_stage_3__4053_,
  data_stage_3__4052_,data_stage_3__4051_,data_stage_3__4050_,data_stage_3__4049_,
  data_stage_3__4048_,data_stage_3__4047_,data_stage_3__4046_,data_stage_3__4045_,
  data_stage_3__4044_,data_stage_3__4043_,data_stage_3__4042_,data_stage_3__4041_,
  data_stage_3__4040_,data_stage_3__4039_,data_stage_3__4038_,data_stage_3__4037_,
  data_stage_3__4036_,data_stage_3__4035_,data_stage_3__4034_,data_stage_3__4033_,
  data_stage_3__4032_,data_stage_3__4031_,data_stage_3__4030_,data_stage_3__4029_,
  data_stage_3__4028_,data_stage_3__4027_,data_stage_3__4026_,data_stage_3__4025_,
  data_stage_3__4024_,data_stage_3__4023_,data_stage_3__4022_,data_stage_3__4021_,
  data_stage_3__4020_,data_stage_3__4019_,data_stage_3__4018_,data_stage_3__4017_,
  data_stage_3__4016_,data_stage_3__4015_,data_stage_3__4014_,data_stage_3__4013_,
  data_stage_3__4012_,data_stage_3__4011_,data_stage_3__4010_,data_stage_3__4009_,
  data_stage_3__4008_,data_stage_3__4007_,data_stage_3__4006_,data_stage_3__4005_,
  data_stage_3__4004_,data_stage_3__4003_,data_stage_3__4002_,data_stage_3__4001_,
  data_stage_3__4000_,data_stage_3__3999_,data_stage_3__3998_,data_stage_3__3997_,
  data_stage_3__3996_,data_stage_3__3995_,data_stage_3__3994_,data_stage_3__3993_,
  data_stage_3__3992_,data_stage_3__3991_,data_stage_3__3990_,data_stage_3__3989_,
  data_stage_3__3988_,data_stage_3__3987_,data_stage_3__3986_,data_stage_3__3985_,
  data_stage_3__3984_,data_stage_3__3983_,data_stage_3__3982_,data_stage_3__3981_,
  data_stage_3__3980_,data_stage_3__3979_,data_stage_3__3978_,data_stage_3__3977_,
  data_stage_3__3976_,data_stage_3__3975_,data_stage_3__3974_,data_stage_3__3973_,
  data_stage_3__3972_,data_stage_3__3971_,data_stage_3__3970_,data_stage_3__3969_,
  data_stage_3__3968_,data_stage_3__3967_,data_stage_3__3966_,data_stage_3__3965_,
  data_stage_3__3964_,data_stage_3__3963_,data_stage_3__3962_,data_stage_3__3961_,
  data_stage_3__3960_,data_stage_3__3959_,data_stage_3__3958_,data_stage_3__3957_,
  data_stage_3__3956_,data_stage_3__3955_,data_stage_3__3954_,data_stage_3__3953_,
  data_stage_3__3952_,data_stage_3__3951_,data_stage_3__3950_,data_stage_3__3949_,
  data_stage_3__3948_,data_stage_3__3947_,data_stage_3__3946_,data_stage_3__3945_,
  data_stage_3__3944_,data_stage_3__3943_,data_stage_3__3942_,data_stage_3__3941_,
  data_stage_3__3940_,data_stage_3__3939_,data_stage_3__3938_,data_stage_3__3937_,
  data_stage_3__3936_,data_stage_3__3935_,data_stage_3__3934_,data_stage_3__3933_,
  data_stage_3__3932_,data_stage_3__3931_,data_stage_3__3930_,data_stage_3__3929_,
  data_stage_3__3928_,data_stage_3__3927_,data_stage_3__3926_,data_stage_3__3925_,
  data_stage_3__3924_,data_stage_3__3923_,data_stage_3__3922_,data_stage_3__3921_,
  data_stage_3__3920_,data_stage_3__3919_,data_stage_3__3918_,data_stage_3__3917_,
  data_stage_3__3916_,data_stage_3__3915_,data_stage_3__3914_,data_stage_3__3913_,
  data_stage_3__3912_,data_stage_3__3911_,data_stage_3__3910_,data_stage_3__3909_,
  data_stage_3__3908_,data_stage_3__3907_,data_stage_3__3906_,data_stage_3__3905_,
  data_stage_3__3904_,data_stage_3__3903_,data_stage_3__3902_,data_stage_3__3901_,
  data_stage_3__3900_,data_stage_3__3899_,data_stage_3__3898_,data_stage_3__3897_,
  data_stage_3__3896_,data_stage_3__3895_,data_stage_3__3894_,data_stage_3__3893_,
  data_stage_3__3892_,data_stage_3__3891_,data_stage_3__3890_,data_stage_3__3889_,
  data_stage_3__3888_,data_stage_3__3887_,data_stage_3__3886_,data_stage_3__3885_,
  data_stage_3__3884_,data_stage_3__3883_,data_stage_3__3882_,data_stage_3__3881_,
  data_stage_3__3880_,data_stage_3__3879_,data_stage_3__3878_,data_stage_3__3877_,
  data_stage_3__3876_,data_stage_3__3875_,data_stage_3__3874_,data_stage_3__3873_,
  data_stage_3__3872_,data_stage_3__3871_,data_stage_3__3870_,data_stage_3__3869_,
  data_stage_3__3868_,data_stage_3__3867_,data_stage_3__3866_,data_stage_3__3865_,
  data_stage_3__3864_,data_stage_3__3863_,data_stage_3__3862_,data_stage_3__3861_,
  data_stage_3__3860_,data_stage_3__3859_,data_stage_3__3858_,data_stage_3__3857_,
  data_stage_3__3856_,data_stage_3__3855_,data_stage_3__3854_,data_stage_3__3853_,
  data_stage_3__3852_,data_stage_3__3851_,data_stage_3__3850_,data_stage_3__3849_,
  data_stage_3__3848_,data_stage_3__3847_,data_stage_3__3846_,data_stage_3__3845_,
  data_stage_3__3844_,data_stage_3__3843_,data_stage_3__3842_,data_stage_3__3841_,
  data_stage_3__3840_,data_stage_3__3839_,data_stage_3__3838_,data_stage_3__3837_,
  data_stage_3__3836_,data_stage_3__3835_,data_stage_3__3834_,data_stage_3__3833_,
  data_stage_3__3832_,data_stage_3__3831_,data_stage_3__3830_,data_stage_3__3829_,
  data_stage_3__3828_,data_stage_3__3827_,data_stage_3__3826_,data_stage_3__3825_,
  data_stage_3__3824_,data_stage_3__3823_,data_stage_3__3822_,data_stage_3__3821_,
  data_stage_3__3820_,data_stage_3__3819_,data_stage_3__3818_,data_stage_3__3817_,
  data_stage_3__3816_,data_stage_3__3815_,data_stage_3__3814_,data_stage_3__3813_,
  data_stage_3__3812_,data_stage_3__3811_,data_stage_3__3810_,data_stage_3__3809_,
  data_stage_3__3808_,data_stage_3__3807_,data_stage_3__3806_,data_stage_3__3805_,
  data_stage_3__3804_,data_stage_3__3803_,data_stage_3__3802_,data_stage_3__3801_,
  data_stage_3__3800_,data_stage_3__3799_,data_stage_3__3798_,data_stage_3__3797_,
  data_stage_3__3796_,data_stage_3__3795_,data_stage_3__3794_,data_stage_3__3793_,
  data_stage_3__3792_,data_stage_3__3791_,data_stage_3__3790_,data_stage_3__3789_,
  data_stage_3__3788_,data_stage_3__3787_,data_stage_3__3786_,data_stage_3__3785_,
  data_stage_3__3784_,data_stage_3__3783_,data_stage_3__3782_,data_stage_3__3781_,
  data_stage_3__3780_,data_stage_3__3779_,data_stage_3__3778_,data_stage_3__3777_,
  data_stage_3__3776_,data_stage_3__3775_,data_stage_3__3774_,data_stage_3__3773_,
  data_stage_3__3772_,data_stage_3__3771_,data_stage_3__3770_,data_stage_3__3769_,
  data_stage_3__3768_,data_stage_3__3767_,data_stage_3__3766_,data_stage_3__3765_,
  data_stage_3__3764_,data_stage_3__3763_,data_stage_3__3762_,data_stage_3__3761_,
  data_stage_3__3760_,data_stage_3__3759_,data_stage_3__3758_,data_stage_3__3757_,
  data_stage_3__3756_,data_stage_3__3755_,data_stage_3__3754_,data_stage_3__3753_,
  data_stage_3__3752_,data_stage_3__3751_,data_stage_3__3750_,data_stage_3__3749_,
  data_stage_3__3748_,data_stage_3__3747_,data_stage_3__3746_,data_stage_3__3745_,
  data_stage_3__3744_,data_stage_3__3743_,data_stage_3__3742_,data_stage_3__3741_,
  data_stage_3__3740_,data_stage_3__3739_,data_stage_3__3738_,data_stage_3__3737_,
  data_stage_3__3736_,data_stage_3__3735_,data_stage_3__3734_,data_stage_3__3733_,
  data_stage_3__3732_,data_stage_3__3731_,data_stage_3__3730_,data_stage_3__3729_,
  data_stage_3__3728_,data_stage_3__3727_,data_stage_3__3726_,data_stage_3__3725_,
  data_stage_3__3724_,data_stage_3__3723_,data_stage_3__3722_,data_stage_3__3721_,
  data_stage_3__3720_,data_stage_3__3719_,data_stage_3__3718_,data_stage_3__3717_,
  data_stage_3__3716_,data_stage_3__3715_,data_stage_3__3714_,data_stage_3__3713_,
  data_stage_3__3712_,data_stage_3__3711_,data_stage_3__3710_,data_stage_3__3709_,
  data_stage_3__3708_,data_stage_3__3707_,data_stage_3__3706_,data_stage_3__3705_,
  data_stage_3__3704_,data_stage_3__3703_,data_stage_3__3702_,data_stage_3__3701_,
  data_stage_3__3700_,data_stage_3__3699_,data_stage_3__3698_,data_stage_3__3697_,
  data_stage_3__3696_,data_stage_3__3695_,data_stage_3__3694_,data_stage_3__3693_,
  data_stage_3__3692_,data_stage_3__3691_,data_stage_3__3690_,data_stage_3__3689_,
  data_stage_3__3688_,data_stage_3__3687_,data_stage_3__3686_,data_stage_3__3685_,
  data_stage_3__3684_,data_stage_3__3683_,data_stage_3__3682_,data_stage_3__3681_,
  data_stage_3__3680_,data_stage_3__3679_,data_stage_3__3678_,data_stage_3__3677_,
  data_stage_3__3676_,data_stage_3__3675_,data_stage_3__3674_,data_stage_3__3673_,
  data_stage_3__3672_,data_stage_3__3671_,data_stage_3__3670_,data_stage_3__3669_,
  data_stage_3__3668_,data_stage_3__3667_,data_stage_3__3666_,data_stage_3__3665_,
  data_stage_3__3664_,data_stage_3__3663_,data_stage_3__3662_,data_stage_3__3661_,
  data_stage_3__3660_,data_stage_3__3659_,data_stage_3__3658_,data_stage_3__3657_,
  data_stage_3__3656_,data_stage_3__3655_,data_stage_3__3654_,data_stage_3__3653_,
  data_stage_3__3652_,data_stage_3__3651_,data_stage_3__3650_,data_stage_3__3649_,
  data_stage_3__3648_,data_stage_3__3647_,data_stage_3__3646_,data_stage_3__3645_,
  data_stage_3__3644_,data_stage_3__3643_,data_stage_3__3642_,data_stage_3__3641_,
  data_stage_3__3640_,data_stage_3__3639_,data_stage_3__3638_,data_stage_3__3637_,
  data_stage_3__3636_,data_stage_3__3635_,data_stage_3__3634_,data_stage_3__3633_,
  data_stage_3__3632_,data_stage_3__3631_,data_stage_3__3630_,data_stage_3__3629_,
  data_stage_3__3628_,data_stage_3__3627_,data_stage_3__3626_,data_stage_3__3625_,
  data_stage_3__3624_,data_stage_3__3623_,data_stage_3__3622_,data_stage_3__3621_,
  data_stage_3__3620_,data_stage_3__3619_,data_stage_3__3618_,data_stage_3__3617_,
  data_stage_3__3616_,data_stage_3__3615_,data_stage_3__3614_,data_stage_3__3613_,
  data_stage_3__3612_,data_stage_3__3611_,data_stage_3__3610_,data_stage_3__3609_,
  data_stage_3__3608_,data_stage_3__3607_,data_stage_3__3606_,data_stage_3__3605_,
  data_stage_3__3604_,data_stage_3__3603_,data_stage_3__3602_,data_stage_3__3601_,
  data_stage_3__3600_,data_stage_3__3599_,data_stage_3__3598_,data_stage_3__3597_,
  data_stage_3__3596_,data_stage_3__3595_,data_stage_3__3594_,data_stage_3__3593_,
  data_stage_3__3592_,data_stage_3__3591_,data_stage_3__3590_,data_stage_3__3589_,
  data_stage_3__3588_,data_stage_3__3587_,data_stage_3__3586_,data_stage_3__3585_,
  data_stage_3__3584_,data_stage_3__3583_,data_stage_3__3582_,data_stage_3__3581_,
  data_stage_3__3580_,data_stage_3__3579_,data_stage_3__3578_,data_stage_3__3577_,
  data_stage_3__3576_,data_stage_3__3575_,data_stage_3__3574_,data_stage_3__3573_,
  data_stage_3__3572_,data_stage_3__3571_,data_stage_3__3570_,data_stage_3__3569_,
  data_stage_3__3568_,data_stage_3__3567_,data_stage_3__3566_,data_stage_3__3565_,
  data_stage_3__3564_,data_stage_3__3563_,data_stage_3__3562_,data_stage_3__3561_,
  data_stage_3__3560_,data_stage_3__3559_,data_stage_3__3558_,data_stage_3__3557_,
  data_stage_3__3556_,data_stage_3__3555_,data_stage_3__3554_,data_stage_3__3553_,
  data_stage_3__3552_,data_stage_3__3551_,data_stage_3__3550_,data_stage_3__3549_,
  data_stage_3__3548_,data_stage_3__3547_,data_stage_3__3546_,data_stage_3__3545_,
  data_stage_3__3544_,data_stage_3__3543_,data_stage_3__3542_,data_stage_3__3541_,
  data_stage_3__3540_,data_stage_3__3539_,data_stage_3__3538_,data_stage_3__3537_,
  data_stage_3__3536_,data_stage_3__3535_,data_stage_3__3534_,data_stage_3__3533_,
  data_stage_3__3532_,data_stage_3__3531_,data_stage_3__3530_,data_stage_3__3529_,
  data_stage_3__3528_,data_stage_3__3527_,data_stage_3__3526_,data_stage_3__3525_,
  data_stage_3__3524_,data_stage_3__3523_,data_stage_3__3522_,data_stage_3__3521_,
  data_stage_3__3520_,data_stage_3__3519_,data_stage_3__3518_,data_stage_3__3517_,
  data_stage_3__3516_,data_stage_3__3515_,data_stage_3__3514_,data_stage_3__3513_,
  data_stage_3__3512_,data_stage_3__3511_,data_stage_3__3510_,data_stage_3__3509_,
  data_stage_3__3508_,data_stage_3__3507_,data_stage_3__3506_,data_stage_3__3505_,
  data_stage_3__3504_,data_stage_3__3503_,data_stage_3__3502_,data_stage_3__3501_,
  data_stage_3__3500_,data_stage_3__3499_,data_stage_3__3498_,data_stage_3__3497_,
  data_stage_3__3496_,data_stage_3__3495_,data_stage_3__3494_,data_stage_3__3493_,
  data_stage_3__3492_,data_stage_3__3491_,data_stage_3__3490_,data_stage_3__3489_,
  data_stage_3__3488_,data_stage_3__3487_,data_stage_3__3486_,data_stage_3__3485_,
  data_stage_3__3484_,data_stage_3__3483_,data_stage_3__3482_,data_stage_3__3481_,
  data_stage_3__3480_,data_stage_3__3479_,data_stage_3__3478_,data_stage_3__3477_,
  data_stage_3__3476_,data_stage_3__3475_,data_stage_3__3474_,data_stage_3__3473_,
  data_stage_3__3472_,data_stage_3__3471_,data_stage_3__3470_,data_stage_3__3469_,
  data_stage_3__3468_,data_stage_3__3467_,data_stage_3__3466_,data_stage_3__3465_,
  data_stage_3__3464_,data_stage_3__3463_,data_stage_3__3462_,data_stage_3__3461_,
  data_stage_3__3460_,data_stage_3__3459_,data_stage_3__3458_,data_stage_3__3457_,
  data_stage_3__3456_,data_stage_3__3455_,data_stage_3__3454_,data_stage_3__3453_,
  data_stage_3__3452_,data_stage_3__3451_,data_stage_3__3450_,data_stage_3__3449_,
  data_stage_3__3448_,data_stage_3__3447_,data_stage_3__3446_,data_stage_3__3445_,
  data_stage_3__3444_,data_stage_3__3443_,data_stage_3__3442_,data_stage_3__3441_,
  data_stage_3__3440_,data_stage_3__3439_,data_stage_3__3438_,data_stage_3__3437_,
  data_stage_3__3436_,data_stage_3__3435_,data_stage_3__3434_,data_stage_3__3433_,
  data_stage_3__3432_,data_stage_3__3431_,data_stage_3__3430_,data_stage_3__3429_,
  data_stage_3__3428_,data_stage_3__3427_,data_stage_3__3426_,data_stage_3__3425_,
  data_stage_3__3424_,data_stage_3__3423_,data_stage_3__3422_,data_stage_3__3421_,
  data_stage_3__3420_,data_stage_3__3419_,data_stage_3__3418_,data_stage_3__3417_,
  data_stage_3__3416_,data_stage_3__3415_,data_stage_3__3414_,data_stage_3__3413_,
  data_stage_3__3412_,data_stage_3__3411_,data_stage_3__3410_,data_stage_3__3409_,
  data_stage_3__3408_,data_stage_3__3407_,data_stage_3__3406_,data_stage_3__3405_,
  data_stage_3__3404_,data_stage_3__3403_,data_stage_3__3402_,data_stage_3__3401_,
  data_stage_3__3400_,data_stage_3__3399_,data_stage_3__3398_,data_stage_3__3397_,
  data_stage_3__3396_,data_stage_3__3395_,data_stage_3__3394_,data_stage_3__3393_,
  data_stage_3__3392_,data_stage_3__3391_,data_stage_3__3390_,data_stage_3__3389_,
  data_stage_3__3388_,data_stage_3__3387_,data_stage_3__3386_,data_stage_3__3385_,
  data_stage_3__3384_,data_stage_3__3383_,data_stage_3__3382_,data_stage_3__3381_,
  data_stage_3__3380_,data_stage_3__3379_,data_stage_3__3378_,data_stage_3__3377_,
  data_stage_3__3376_,data_stage_3__3375_,data_stage_3__3374_,data_stage_3__3373_,
  data_stage_3__3372_,data_stage_3__3371_,data_stage_3__3370_,data_stage_3__3369_,
  data_stage_3__3368_,data_stage_3__3367_,data_stage_3__3366_,data_stage_3__3365_,
  data_stage_3__3364_,data_stage_3__3363_,data_stage_3__3362_,data_stage_3__3361_,
  data_stage_3__3360_,data_stage_3__3359_,data_stage_3__3358_,data_stage_3__3357_,
  data_stage_3__3356_,data_stage_3__3355_,data_stage_3__3354_,data_stage_3__3353_,
  data_stage_3__3352_,data_stage_3__3351_,data_stage_3__3350_,data_stage_3__3349_,
  data_stage_3__3348_,data_stage_3__3347_,data_stage_3__3346_,data_stage_3__3345_,
  data_stage_3__3344_,data_stage_3__3343_,data_stage_3__3342_,data_stage_3__3341_,
  data_stage_3__3340_,data_stage_3__3339_,data_stage_3__3338_,data_stage_3__3337_,
  data_stage_3__3336_,data_stage_3__3335_,data_stage_3__3334_,data_stage_3__3333_,
  data_stage_3__3332_,data_stage_3__3331_,data_stage_3__3330_,data_stage_3__3329_,
  data_stage_3__3328_,data_stage_3__3327_,data_stage_3__3326_,data_stage_3__3325_,
  data_stage_3__3324_,data_stage_3__3323_,data_stage_3__3322_,data_stage_3__3321_,
  data_stage_3__3320_,data_stage_3__3319_,data_stage_3__3318_,data_stage_3__3317_,
  data_stage_3__3316_,data_stage_3__3315_,data_stage_3__3314_,data_stage_3__3313_,
  data_stage_3__3312_,data_stage_3__3311_,data_stage_3__3310_,data_stage_3__3309_,
  data_stage_3__3308_,data_stage_3__3307_,data_stage_3__3306_,data_stage_3__3305_,
  data_stage_3__3304_,data_stage_3__3303_,data_stage_3__3302_,data_stage_3__3301_,
  data_stage_3__3300_,data_stage_3__3299_,data_stage_3__3298_,data_stage_3__3297_,
  data_stage_3__3296_,data_stage_3__3295_,data_stage_3__3294_,data_stage_3__3293_,
  data_stage_3__3292_,data_stage_3__3291_,data_stage_3__3290_,data_stage_3__3289_,
  data_stage_3__3288_,data_stage_3__3287_,data_stage_3__3286_,data_stage_3__3285_,
  data_stage_3__3284_,data_stage_3__3283_,data_stage_3__3282_,data_stage_3__3281_,
  data_stage_3__3280_,data_stage_3__3279_,data_stage_3__3278_,data_stage_3__3277_,
  data_stage_3__3276_,data_stage_3__3275_,data_stage_3__3274_,data_stage_3__3273_,
  data_stage_3__3272_,data_stage_3__3271_,data_stage_3__3270_,data_stage_3__3269_,
  data_stage_3__3268_,data_stage_3__3267_,data_stage_3__3266_,data_stage_3__3265_,
  data_stage_3__3264_,data_stage_3__3263_,data_stage_3__3262_,data_stage_3__3261_,
  data_stage_3__3260_,data_stage_3__3259_,data_stage_3__3258_,data_stage_3__3257_,
  data_stage_3__3256_,data_stage_3__3255_,data_stage_3__3254_,data_stage_3__3253_,
  data_stage_3__3252_,data_stage_3__3251_,data_stage_3__3250_,data_stage_3__3249_,
  data_stage_3__3248_,data_stage_3__3247_,data_stage_3__3246_,data_stage_3__3245_,
  data_stage_3__3244_,data_stage_3__3243_,data_stage_3__3242_,data_stage_3__3241_,
  data_stage_3__3240_,data_stage_3__3239_,data_stage_3__3238_,data_stage_3__3237_,
  data_stage_3__3236_,data_stage_3__3235_,data_stage_3__3234_,data_stage_3__3233_,
  data_stage_3__3232_,data_stage_3__3231_,data_stage_3__3230_,data_stage_3__3229_,
  data_stage_3__3228_,data_stage_3__3227_,data_stage_3__3226_,data_stage_3__3225_,
  data_stage_3__3224_,data_stage_3__3223_,data_stage_3__3222_,data_stage_3__3221_,
  data_stage_3__3220_,data_stage_3__3219_,data_stage_3__3218_,data_stage_3__3217_,
  data_stage_3__3216_,data_stage_3__3215_,data_stage_3__3214_,data_stage_3__3213_,
  data_stage_3__3212_,data_stage_3__3211_,data_stage_3__3210_,data_stage_3__3209_,
  data_stage_3__3208_,data_stage_3__3207_,data_stage_3__3206_,data_stage_3__3205_,
  data_stage_3__3204_,data_stage_3__3203_,data_stage_3__3202_,data_stage_3__3201_,
  data_stage_3__3200_,data_stage_3__3199_,data_stage_3__3198_,data_stage_3__3197_,
  data_stage_3__3196_,data_stage_3__3195_,data_stage_3__3194_,data_stage_3__3193_,
  data_stage_3__3192_,data_stage_3__3191_,data_stage_3__3190_,data_stage_3__3189_,
  data_stage_3__3188_,data_stage_3__3187_,data_stage_3__3186_,data_stage_3__3185_,
  data_stage_3__3184_,data_stage_3__3183_,data_stage_3__3182_,data_stage_3__3181_,
  data_stage_3__3180_,data_stage_3__3179_,data_stage_3__3178_,data_stage_3__3177_,
  data_stage_3__3176_,data_stage_3__3175_,data_stage_3__3174_,data_stage_3__3173_,
  data_stage_3__3172_,data_stage_3__3171_,data_stage_3__3170_,data_stage_3__3169_,
  data_stage_3__3168_,data_stage_3__3167_,data_stage_3__3166_,data_stage_3__3165_,
  data_stage_3__3164_,data_stage_3__3163_,data_stage_3__3162_,data_stage_3__3161_,
  data_stage_3__3160_,data_stage_3__3159_,data_stage_3__3158_,data_stage_3__3157_,
  data_stage_3__3156_,data_stage_3__3155_,data_stage_3__3154_,data_stage_3__3153_,
  data_stage_3__3152_,data_stage_3__3151_,data_stage_3__3150_,data_stage_3__3149_,
  data_stage_3__3148_,data_stage_3__3147_,data_stage_3__3146_,data_stage_3__3145_,
  data_stage_3__3144_,data_stage_3__3143_,data_stage_3__3142_,data_stage_3__3141_,
  data_stage_3__3140_,data_stage_3__3139_,data_stage_3__3138_,data_stage_3__3137_,
  data_stage_3__3136_,data_stage_3__3135_,data_stage_3__3134_,data_stage_3__3133_,
  data_stage_3__3132_,data_stage_3__3131_,data_stage_3__3130_,data_stage_3__3129_,
  data_stage_3__3128_,data_stage_3__3127_,data_stage_3__3126_,data_stage_3__3125_,
  data_stage_3__3124_,data_stage_3__3123_,data_stage_3__3122_,data_stage_3__3121_,
  data_stage_3__3120_,data_stage_3__3119_,data_stage_3__3118_,data_stage_3__3117_,
  data_stage_3__3116_,data_stage_3__3115_,data_stage_3__3114_,data_stage_3__3113_,
  data_stage_3__3112_,data_stage_3__3111_,data_stage_3__3110_,data_stage_3__3109_,
  data_stage_3__3108_,data_stage_3__3107_,data_stage_3__3106_,data_stage_3__3105_,
  data_stage_3__3104_,data_stage_3__3103_,data_stage_3__3102_,data_stage_3__3101_,
  data_stage_3__3100_,data_stage_3__3099_,data_stage_3__3098_,data_stage_3__3097_,
  data_stage_3__3096_,data_stage_3__3095_,data_stage_3__3094_,data_stage_3__3093_,
  data_stage_3__3092_,data_stage_3__3091_,data_stage_3__3090_,data_stage_3__3089_,
  data_stage_3__3088_,data_stage_3__3087_,data_stage_3__3086_,data_stage_3__3085_,
  data_stage_3__3084_,data_stage_3__3083_,data_stage_3__3082_,data_stage_3__3081_,
  data_stage_3__3080_,data_stage_3__3079_,data_stage_3__3078_,data_stage_3__3077_,
  data_stage_3__3076_,data_stage_3__3075_,data_stage_3__3074_,data_stage_3__3073_,
  data_stage_3__3072_,data_stage_3__3071_,data_stage_3__3070_,data_stage_3__3069_,
  data_stage_3__3068_,data_stage_3__3067_,data_stage_3__3066_,data_stage_3__3065_,
  data_stage_3__3064_,data_stage_3__3063_,data_stage_3__3062_,data_stage_3__3061_,
  data_stage_3__3060_,data_stage_3__3059_,data_stage_3__3058_,data_stage_3__3057_,
  data_stage_3__3056_,data_stage_3__3055_,data_stage_3__3054_,data_stage_3__3053_,
  data_stage_3__3052_,data_stage_3__3051_,data_stage_3__3050_,data_stage_3__3049_,
  data_stage_3__3048_,data_stage_3__3047_,data_stage_3__3046_,data_stage_3__3045_,
  data_stage_3__3044_,data_stage_3__3043_,data_stage_3__3042_,data_stage_3__3041_,
  data_stage_3__3040_,data_stage_3__3039_,data_stage_3__3038_,data_stage_3__3037_,
  data_stage_3__3036_,data_stage_3__3035_,data_stage_3__3034_,data_stage_3__3033_,
  data_stage_3__3032_,data_stage_3__3031_,data_stage_3__3030_,data_stage_3__3029_,
  data_stage_3__3028_,data_stage_3__3027_,data_stage_3__3026_,data_stage_3__3025_,
  data_stage_3__3024_,data_stage_3__3023_,data_stage_3__3022_,data_stage_3__3021_,
  data_stage_3__3020_,data_stage_3__3019_,data_stage_3__3018_,data_stage_3__3017_,
  data_stage_3__3016_,data_stage_3__3015_,data_stage_3__3014_,data_stage_3__3013_,
  data_stage_3__3012_,data_stage_3__3011_,data_stage_3__3010_,data_stage_3__3009_,
  data_stage_3__3008_,data_stage_3__3007_,data_stage_3__3006_,data_stage_3__3005_,
  data_stage_3__3004_,data_stage_3__3003_,data_stage_3__3002_,data_stage_3__3001_,
  data_stage_3__3000_,data_stage_3__2999_,data_stage_3__2998_,data_stage_3__2997_,
  data_stage_3__2996_,data_stage_3__2995_,data_stage_3__2994_,data_stage_3__2993_,
  data_stage_3__2992_,data_stage_3__2991_,data_stage_3__2990_,data_stage_3__2989_,
  data_stage_3__2988_,data_stage_3__2987_,data_stage_3__2986_,data_stage_3__2985_,
  data_stage_3__2984_,data_stage_3__2983_,data_stage_3__2982_,data_stage_3__2981_,
  data_stage_3__2980_,data_stage_3__2979_,data_stage_3__2978_,data_stage_3__2977_,
  data_stage_3__2976_,data_stage_3__2975_,data_stage_3__2974_,data_stage_3__2973_,
  data_stage_3__2972_,data_stage_3__2971_,data_stage_3__2970_,data_stage_3__2969_,
  data_stage_3__2968_,data_stage_3__2967_,data_stage_3__2966_,data_stage_3__2965_,
  data_stage_3__2964_,data_stage_3__2963_,data_stage_3__2962_,data_stage_3__2961_,
  data_stage_3__2960_,data_stage_3__2959_,data_stage_3__2958_,data_stage_3__2957_,
  data_stage_3__2956_,data_stage_3__2955_,data_stage_3__2954_,data_stage_3__2953_,
  data_stage_3__2952_,data_stage_3__2951_,data_stage_3__2950_,data_stage_3__2949_,
  data_stage_3__2948_,data_stage_3__2947_,data_stage_3__2946_,data_stage_3__2945_,
  data_stage_3__2944_,data_stage_3__2943_,data_stage_3__2942_,data_stage_3__2941_,
  data_stage_3__2940_,data_stage_3__2939_,data_stage_3__2938_,data_stage_3__2937_,
  data_stage_3__2936_,data_stage_3__2935_,data_stage_3__2934_,data_stage_3__2933_,
  data_stage_3__2932_,data_stage_3__2931_,data_stage_3__2930_,data_stage_3__2929_,
  data_stage_3__2928_,data_stage_3__2927_,data_stage_3__2926_,data_stage_3__2925_,
  data_stage_3__2924_,data_stage_3__2923_,data_stage_3__2922_,data_stage_3__2921_,
  data_stage_3__2920_,data_stage_3__2919_,data_stage_3__2918_,data_stage_3__2917_,
  data_stage_3__2916_,data_stage_3__2915_,data_stage_3__2914_,data_stage_3__2913_,
  data_stage_3__2912_,data_stage_3__2911_,data_stage_3__2910_,data_stage_3__2909_,
  data_stage_3__2908_,data_stage_3__2907_,data_stage_3__2906_,data_stage_3__2905_,
  data_stage_3__2904_,data_stage_3__2903_,data_stage_3__2902_,data_stage_3__2901_,
  data_stage_3__2900_,data_stage_3__2899_,data_stage_3__2898_,data_stage_3__2897_,
  data_stage_3__2896_,data_stage_3__2895_,data_stage_3__2894_,data_stage_3__2893_,
  data_stage_3__2892_,data_stage_3__2891_,data_stage_3__2890_,data_stage_3__2889_,
  data_stage_3__2888_,data_stage_3__2887_,data_stage_3__2886_,data_stage_3__2885_,
  data_stage_3__2884_,data_stage_3__2883_,data_stage_3__2882_,data_stage_3__2881_,
  data_stage_3__2880_,data_stage_3__2879_,data_stage_3__2878_,data_stage_3__2877_,
  data_stage_3__2876_,data_stage_3__2875_,data_stage_3__2874_,data_stage_3__2873_,
  data_stage_3__2872_,data_stage_3__2871_,data_stage_3__2870_,data_stage_3__2869_,
  data_stage_3__2868_,data_stage_3__2867_,data_stage_3__2866_,data_stage_3__2865_,
  data_stage_3__2864_,data_stage_3__2863_,data_stage_3__2862_,data_stage_3__2861_,
  data_stage_3__2860_,data_stage_3__2859_,data_stage_3__2858_,data_stage_3__2857_,
  data_stage_3__2856_,data_stage_3__2855_,data_stage_3__2854_,data_stage_3__2853_,
  data_stage_3__2852_,data_stage_3__2851_,data_stage_3__2850_,data_stage_3__2849_,
  data_stage_3__2848_,data_stage_3__2847_,data_stage_3__2846_,data_stage_3__2845_,
  data_stage_3__2844_,data_stage_3__2843_,data_stage_3__2842_,data_stage_3__2841_,
  data_stage_3__2840_,data_stage_3__2839_,data_stage_3__2838_,data_stage_3__2837_,
  data_stage_3__2836_,data_stage_3__2835_,data_stage_3__2834_,data_stage_3__2833_,
  data_stage_3__2832_,data_stage_3__2831_,data_stage_3__2830_,data_stage_3__2829_,
  data_stage_3__2828_,data_stage_3__2827_,data_stage_3__2826_,data_stage_3__2825_,
  data_stage_3__2824_,data_stage_3__2823_,data_stage_3__2822_,data_stage_3__2821_,
  data_stage_3__2820_,data_stage_3__2819_,data_stage_3__2818_,data_stage_3__2817_,
  data_stage_3__2816_,data_stage_3__2815_,data_stage_3__2814_,data_stage_3__2813_,
  data_stage_3__2812_,data_stage_3__2811_,data_stage_3__2810_,data_stage_3__2809_,
  data_stage_3__2808_,data_stage_3__2807_,data_stage_3__2806_,data_stage_3__2805_,
  data_stage_3__2804_,data_stage_3__2803_,data_stage_3__2802_,data_stage_3__2801_,
  data_stage_3__2800_,data_stage_3__2799_,data_stage_3__2798_,data_stage_3__2797_,
  data_stage_3__2796_,data_stage_3__2795_,data_stage_3__2794_,data_stage_3__2793_,
  data_stage_3__2792_,data_stage_3__2791_,data_stage_3__2790_,data_stage_3__2789_,
  data_stage_3__2788_,data_stage_3__2787_,data_stage_3__2786_,data_stage_3__2785_,
  data_stage_3__2784_,data_stage_3__2783_,data_stage_3__2782_,data_stage_3__2781_,
  data_stage_3__2780_,data_stage_3__2779_,data_stage_3__2778_,data_stage_3__2777_,
  data_stage_3__2776_,data_stage_3__2775_,data_stage_3__2774_,data_stage_3__2773_,
  data_stage_3__2772_,data_stage_3__2771_,data_stage_3__2770_,data_stage_3__2769_,
  data_stage_3__2768_,data_stage_3__2767_,data_stage_3__2766_,data_stage_3__2765_,
  data_stage_3__2764_,data_stage_3__2763_,data_stage_3__2762_,data_stage_3__2761_,
  data_stage_3__2760_,data_stage_3__2759_,data_stage_3__2758_,data_stage_3__2757_,
  data_stage_3__2756_,data_stage_3__2755_,data_stage_3__2754_,data_stage_3__2753_,
  data_stage_3__2752_,data_stage_3__2751_,data_stage_3__2750_,data_stage_3__2749_,
  data_stage_3__2748_,data_stage_3__2747_,data_stage_3__2746_,data_stage_3__2745_,
  data_stage_3__2744_,data_stage_3__2743_,data_stage_3__2742_,data_stage_3__2741_,
  data_stage_3__2740_,data_stage_3__2739_,data_stage_3__2738_,data_stage_3__2737_,
  data_stage_3__2736_,data_stage_3__2735_,data_stage_3__2734_,data_stage_3__2733_,
  data_stage_3__2732_,data_stage_3__2731_,data_stage_3__2730_,data_stage_3__2729_,
  data_stage_3__2728_,data_stage_3__2727_,data_stage_3__2726_,data_stage_3__2725_,
  data_stage_3__2724_,data_stage_3__2723_,data_stage_3__2722_,data_stage_3__2721_,
  data_stage_3__2720_,data_stage_3__2719_,data_stage_3__2718_,data_stage_3__2717_,
  data_stage_3__2716_,data_stage_3__2715_,data_stage_3__2714_,data_stage_3__2713_,
  data_stage_3__2712_,data_stage_3__2711_,data_stage_3__2710_,data_stage_3__2709_,
  data_stage_3__2708_,data_stage_3__2707_,data_stage_3__2706_,data_stage_3__2705_,
  data_stage_3__2704_,data_stage_3__2703_,data_stage_3__2702_,data_stage_3__2701_,
  data_stage_3__2700_,data_stage_3__2699_,data_stage_3__2698_,data_stage_3__2697_,
  data_stage_3__2696_,data_stage_3__2695_,data_stage_3__2694_,data_stage_3__2693_,
  data_stage_3__2692_,data_stage_3__2691_,data_stage_3__2690_,data_stage_3__2689_,
  data_stage_3__2688_,data_stage_3__2687_,data_stage_3__2686_,data_stage_3__2685_,
  data_stage_3__2684_,data_stage_3__2683_,data_stage_3__2682_,data_stage_3__2681_,
  data_stage_3__2680_,data_stage_3__2679_,data_stage_3__2678_,data_stage_3__2677_,
  data_stage_3__2676_,data_stage_3__2675_,data_stage_3__2674_,data_stage_3__2673_,
  data_stage_3__2672_,data_stage_3__2671_,data_stage_3__2670_,data_stage_3__2669_,
  data_stage_3__2668_,data_stage_3__2667_,data_stage_3__2666_,data_stage_3__2665_,
  data_stage_3__2664_,data_stage_3__2663_,data_stage_3__2662_,data_stage_3__2661_,
  data_stage_3__2660_,data_stage_3__2659_,data_stage_3__2658_,data_stage_3__2657_,
  data_stage_3__2656_,data_stage_3__2655_,data_stage_3__2654_,data_stage_3__2653_,
  data_stage_3__2652_,data_stage_3__2651_,data_stage_3__2650_,data_stage_3__2649_,
  data_stage_3__2648_,data_stage_3__2647_,data_stage_3__2646_,data_stage_3__2645_,
  data_stage_3__2644_,data_stage_3__2643_,data_stage_3__2642_,data_stage_3__2641_,
  data_stage_3__2640_,data_stage_3__2639_,data_stage_3__2638_,data_stage_3__2637_,
  data_stage_3__2636_,data_stage_3__2635_,data_stage_3__2634_,data_stage_3__2633_,
  data_stage_3__2632_,data_stage_3__2631_,data_stage_3__2630_,data_stage_3__2629_,
  data_stage_3__2628_,data_stage_3__2627_,data_stage_3__2626_,data_stage_3__2625_,
  data_stage_3__2624_,data_stage_3__2623_,data_stage_3__2622_,data_stage_3__2621_,
  data_stage_3__2620_,data_stage_3__2619_,data_stage_3__2618_,data_stage_3__2617_,
  data_stage_3__2616_,data_stage_3__2615_,data_stage_3__2614_,data_stage_3__2613_,
  data_stage_3__2612_,data_stage_3__2611_,data_stage_3__2610_,data_stage_3__2609_,
  data_stage_3__2608_,data_stage_3__2607_,data_stage_3__2606_,data_stage_3__2605_,
  data_stage_3__2604_,data_stage_3__2603_,data_stage_3__2602_,data_stage_3__2601_,
  data_stage_3__2600_,data_stage_3__2599_,data_stage_3__2598_,data_stage_3__2597_,
  data_stage_3__2596_,data_stage_3__2595_,data_stage_3__2594_,data_stage_3__2593_,
  data_stage_3__2592_,data_stage_3__2591_,data_stage_3__2590_,data_stage_3__2589_,
  data_stage_3__2588_,data_stage_3__2587_,data_stage_3__2586_,data_stage_3__2585_,
  data_stage_3__2584_,data_stage_3__2583_,data_stage_3__2582_,data_stage_3__2581_,
  data_stage_3__2580_,data_stage_3__2579_,data_stage_3__2578_,data_stage_3__2577_,
  data_stage_3__2576_,data_stage_3__2575_,data_stage_3__2574_,data_stage_3__2573_,
  data_stage_3__2572_,data_stage_3__2571_,data_stage_3__2570_,data_stage_3__2569_,
  data_stage_3__2568_,data_stage_3__2567_,data_stage_3__2566_,data_stage_3__2565_,
  data_stage_3__2564_,data_stage_3__2563_,data_stage_3__2562_,data_stage_3__2561_,
  data_stage_3__2560_,data_stage_3__2559_,data_stage_3__2558_,data_stage_3__2557_,
  data_stage_3__2556_,data_stage_3__2555_,data_stage_3__2554_,data_stage_3__2553_,
  data_stage_3__2552_,data_stage_3__2551_,data_stage_3__2550_,data_stage_3__2549_,
  data_stage_3__2548_,data_stage_3__2547_,data_stage_3__2546_,data_stage_3__2545_,
  data_stage_3__2544_,data_stage_3__2543_,data_stage_3__2542_,data_stage_3__2541_,
  data_stage_3__2540_,data_stage_3__2539_,data_stage_3__2538_,data_stage_3__2537_,
  data_stage_3__2536_,data_stage_3__2535_,data_stage_3__2534_,data_stage_3__2533_,
  data_stage_3__2532_,data_stage_3__2531_,data_stage_3__2530_,data_stage_3__2529_,
  data_stage_3__2528_,data_stage_3__2527_,data_stage_3__2526_,data_stage_3__2525_,
  data_stage_3__2524_,data_stage_3__2523_,data_stage_3__2522_,data_stage_3__2521_,
  data_stage_3__2520_,data_stage_3__2519_,data_stage_3__2518_,data_stage_3__2517_,
  data_stage_3__2516_,data_stage_3__2515_,data_stage_3__2514_,data_stage_3__2513_,
  data_stage_3__2512_,data_stage_3__2511_,data_stage_3__2510_,data_stage_3__2509_,
  data_stage_3__2508_,data_stage_3__2507_,data_stage_3__2506_,data_stage_3__2505_,
  data_stage_3__2504_,data_stage_3__2503_,data_stage_3__2502_,data_stage_3__2501_,
  data_stage_3__2500_,data_stage_3__2499_,data_stage_3__2498_,data_stage_3__2497_,
  data_stage_3__2496_,data_stage_3__2495_,data_stage_3__2494_,data_stage_3__2493_,
  data_stage_3__2492_,data_stage_3__2491_,data_stage_3__2490_,data_stage_3__2489_,
  data_stage_3__2488_,data_stage_3__2487_,data_stage_3__2486_,data_stage_3__2485_,
  data_stage_3__2484_,data_stage_3__2483_,data_stage_3__2482_,data_stage_3__2481_,
  data_stage_3__2480_,data_stage_3__2479_,data_stage_3__2478_,data_stage_3__2477_,
  data_stage_3__2476_,data_stage_3__2475_,data_stage_3__2474_,data_stage_3__2473_,
  data_stage_3__2472_,data_stage_3__2471_,data_stage_3__2470_,data_stage_3__2469_,
  data_stage_3__2468_,data_stage_3__2467_,data_stage_3__2466_,data_stage_3__2465_,
  data_stage_3__2464_,data_stage_3__2463_,data_stage_3__2462_,data_stage_3__2461_,
  data_stage_3__2460_,data_stage_3__2459_,data_stage_3__2458_,data_stage_3__2457_,
  data_stage_3__2456_,data_stage_3__2455_,data_stage_3__2454_,data_stage_3__2453_,
  data_stage_3__2452_,data_stage_3__2451_,data_stage_3__2450_,data_stage_3__2449_,
  data_stage_3__2448_,data_stage_3__2447_,data_stage_3__2446_,data_stage_3__2445_,
  data_stage_3__2444_,data_stage_3__2443_,data_stage_3__2442_,data_stage_3__2441_,
  data_stage_3__2440_,data_stage_3__2439_,data_stage_3__2438_,data_stage_3__2437_,
  data_stage_3__2436_,data_stage_3__2435_,data_stage_3__2434_,data_stage_3__2433_,
  data_stage_3__2432_,data_stage_3__2431_,data_stage_3__2430_,data_stage_3__2429_,
  data_stage_3__2428_,data_stage_3__2427_,data_stage_3__2426_,data_stage_3__2425_,
  data_stage_3__2424_,data_stage_3__2423_,data_stage_3__2422_,data_stage_3__2421_,
  data_stage_3__2420_,data_stage_3__2419_,data_stage_3__2418_,data_stage_3__2417_,
  data_stage_3__2416_,data_stage_3__2415_,data_stage_3__2414_,data_stage_3__2413_,
  data_stage_3__2412_,data_stage_3__2411_,data_stage_3__2410_,data_stage_3__2409_,
  data_stage_3__2408_,data_stage_3__2407_,data_stage_3__2406_,data_stage_3__2405_,
  data_stage_3__2404_,data_stage_3__2403_,data_stage_3__2402_,data_stage_3__2401_,
  data_stage_3__2400_,data_stage_3__2399_,data_stage_3__2398_,data_stage_3__2397_,
  data_stage_3__2396_,data_stage_3__2395_,data_stage_3__2394_,data_stage_3__2393_,
  data_stage_3__2392_,data_stage_3__2391_,data_stage_3__2390_,data_stage_3__2389_,
  data_stage_3__2388_,data_stage_3__2387_,data_stage_3__2386_,data_stage_3__2385_,
  data_stage_3__2384_,data_stage_3__2383_,data_stage_3__2382_,data_stage_3__2381_,
  data_stage_3__2380_,data_stage_3__2379_,data_stage_3__2378_,data_stage_3__2377_,
  data_stage_3__2376_,data_stage_3__2375_,data_stage_3__2374_,data_stage_3__2373_,
  data_stage_3__2372_,data_stage_3__2371_,data_stage_3__2370_,data_stage_3__2369_,
  data_stage_3__2368_,data_stage_3__2367_,data_stage_3__2366_,data_stage_3__2365_,
  data_stage_3__2364_,data_stage_3__2363_,data_stage_3__2362_,data_stage_3__2361_,
  data_stage_3__2360_,data_stage_3__2359_,data_stage_3__2358_,data_stage_3__2357_,
  data_stage_3__2356_,data_stage_3__2355_,data_stage_3__2354_,data_stage_3__2353_,
  data_stage_3__2352_,data_stage_3__2351_,data_stage_3__2350_,data_stage_3__2349_,
  data_stage_3__2348_,data_stage_3__2347_,data_stage_3__2346_,data_stage_3__2345_,
  data_stage_3__2344_,data_stage_3__2343_,data_stage_3__2342_,data_stage_3__2341_,
  data_stage_3__2340_,data_stage_3__2339_,data_stage_3__2338_,data_stage_3__2337_,
  data_stage_3__2336_,data_stage_3__2335_,data_stage_3__2334_,data_stage_3__2333_,
  data_stage_3__2332_,data_stage_3__2331_,data_stage_3__2330_,data_stage_3__2329_,
  data_stage_3__2328_,data_stage_3__2327_,data_stage_3__2326_,data_stage_3__2325_,
  data_stage_3__2324_,data_stage_3__2323_,data_stage_3__2322_,data_stage_3__2321_,
  data_stage_3__2320_,data_stage_3__2319_,data_stage_3__2318_,data_stage_3__2317_,
  data_stage_3__2316_,data_stage_3__2315_,data_stage_3__2314_,data_stage_3__2313_,
  data_stage_3__2312_,data_stage_3__2311_,data_stage_3__2310_,data_stage_3__2309_,
  data_stage_3__2308_,data_stage_3__2307_,data_stage_3__2306_,data_stage_3__2305_,
  data_stage_3__2304_,data_stage_3__2303_,data_stage_3__2302_,data_stage_3__2301_,
  data_stage_3__2300_,data_stage_3__2299_,data_stage_3__2298_,data_stage_3__2297_,
  data_stage_3__2296_,data_stage_3__2295_,data_stage_3__2294_,data_stage_3__2293_,
  data_stage_3__2292_,data_stage_3__2291_,data_stage_3__2290_,data_stage_3__2289_,
  data_stage_3__2288_,data_stage_3__2287_,data_stage_3__2286_,data_stage_3__2285_,
  data_stage_3__2284_,data_stage_3__2283_,data_stage_3__2282_,data_stage_3__2281_,
  data_stage_3__2280_,data_stage_3__2279_,data_stage_3__2278_,data_stage_3__2277_,
  data_stage_3__2276_,data_stage_3__2275_,data_stage_3__2274_,data_stage_3__2273_,
  data_stage_3__2272_,data_stage_3__2271_,data_stage_3__2270_,data_stage_3__2269_,
  data_stage_3__2268_,data_stage_3__2267_,data_stage_3__2266_,data_stage_3__2265_,
  data_stage_3__2264_,data_stage_3__2263_,data_stage_3__2262_,data_stage_3__2261_,
  data_stage_3__2260_,data_stage_3__2259_,data_stage_3__2258_,data_stage_3__2257_,
  data_stage_3__2256_,data_stage_3__2255_,data_stage_3__2254_,data_stage_3__2253_,
  data_stage_3__2252_,data_stage_3__2251_,data_stage_3__2250_,data_stage_3__2249_,
  data_stage_3__2248_,data_stage_3__2247_,data_stage_3__2246_,data_stage_3__2245_,
  data_stage_3__2244_,data_stage_3__2243_,data_stage_3__2242_,data_stage_3__2241_,
  data_stage_3__2240_,data_stage_3__2239_,data_stage_3__2238_,data_stage_3__2237_,
  data_stage_3__2236_,data_stage_3__2235_,data_stage_3__2234_,data_stage_3__2233_,
  data_stage_3__2232_,data_stage_3__2231_,data_stage_3__2230_,data_stage_3__2229_,
  data_stage_3__2228_,data_stage_3__2227_,data_stage_3__2226_,data_stage_3__2225_,
  data_stage_3__2224_,data_stage_3__2223_,data_stage_3__2222_,data_stage_3__2221_,
  data_stage_3__2220_,data_stage_3__2219_,data_stage_3__2218_,data_stage_3__2217_,
  data_stage_3__2216_,data_stage_3__2215_,data_stage_3__2214_,data_stage_3__2213_,
  data_stage_3__2212_,data_stage_3__2211_,data_stage_3__2210_,data_stage_3__2209_,
  data_stage_3__2208_,data_stage_3__2207_,data_stage_3__2206_,data_stage_3__2205_,
  data_stage_3__2204_,data_stage_3__2203_,data_stage_3__2202_,data_stage_3__2201_,
  data_stage_3__2200_,data_stage_3__2199_,data_stage_3__2198_,data_stage_3__2197_,
  data_stage_3__2196_,data_stage_3__2195_,data_stage_3__2194_,data_stage_3__2193_,
  data_stage_3__2192_,data_stage_3__2191_,data_stage_3__2190_,data_stage_3__2189_,
  data_stage_3__2188_,data_stage_3__2187_,data_stage_3__2186_,data_stage_3__2185_,
  data_stage_3__2184_,data_stage_3__2183_,data_stage_3__2182_,data_stage_3__2181_,
  data_stage_3__2180_,data_stage_3__2179_,data_stage_3__2178_,data_stage_3__2177_,
  data_stage_3__2176_,data_stage_3__2175_,data_stage_3__2174_,data_stage_3__2173_,
  data_stage_3__2172_,data_stage_3__2171_,data_stage_3__2170_,data_stage_3__2169_,
  data_stage_3__2168_,data_stage_3__2167_,data_stage_3__2166_,data_stage_3__2165_,
  data_stage_3__2164_,data_stage_3__2163_,data_stage_3__2162_,data_stage_3__2161_,
  data_stage_3__2160_,data_stage_3__2159_,data_stage_3__2158_,data_stage_3__2157_,
  data_stage_3__2156_,data_stage_3__2155_,data_stage_3__2154_,data_stage_3__2153_,
  data_stage_3__2152_,data_stage_3__2151_,data_stage_3__2150_,data_stage_3__2149_,
  data_stage_3__2148_,data_stage_3__2147_,data_stage_3__2146_,data_stage_3__2145_,
  data_stage_3__2144_,data_stage_3__2143_,data_stage_3__2142_,data_stage_3__2141_,
  data_stage_3__2140_,data_stage_3__2139_,data_stage_3__2138_,data_stage_3__2137_,
  data_stage_3__2136_,data_stage_3__2135_,data_stage_3__2134_,data_stage_3__2133_,
  data_stage_3__2132_,data_stage_3__2131_,data_stage_3__2130_,data_stage_3__2129_,
  data_stage_3__2128_,data_stage_3__2127_,data_stage_3__2126_,data_stage_3__2125_,
  data_stage_3__2124_,data_stage_3__2123_,data_stage_3__2122_,data_stage_3__2121_,
  data_stage_3__2120_,data_stage_3__2119_,data_stage_3__2118_,data_stage_3__2117_,
  data_stage_3__2116_,data_stage_3__2115_,data_stage_3__2114_,data_stage_3__2113_,
  data_stage_3__2112_,data_stage_3__2111_,data_stage_3__2110_,data_stage_3__2109_,
  data_stage_3__2108_,data_stage_3__2107_,data_stage_3__2106_,data_stage_3__2105_,
  data_stage_3__2104_,data_stage_3__2103_,data_stage_3__2102_,data_stage_3__2101_,
  data_stage_3__2100_,data_stage_3__2099_,data_stage_3__2098_,data_stage_3__2097_,
  data_stage_3__2096_,data_stage_3__2095_,data_stage_3__2094_,data_stage_3__2093_,
  data_stage_3__2092_,data_stage_3__2091_,data_stage_3__2090_,data_stage_3__2089_,
  data_stage_3__2088_,data_stage_3__2087_,data_stage_3__2086_,data_stage_3__2085_,
  data_stage_3__2084_,data_stage_3__2083_,data_stage_3__2082_,data_stage_3__2081_,
  data_stage_3__2080_,data_stage_3__2079_,data_stage_3__2078_,data_stage_3__2077_,
  data_stage_3__2076_,data_stage_3__2075_,data_stage_3__2074_,data_stage_3__2073_,
  data_stage_3__2072_,data_stage_3__2071_,data_stage_3__2070_,data_stage_3__2069_,
  data_stage_3__2068_,data_stage_3__2067_,data_stage_3__2066_,data_stage_3__2065_,
  data_stage_3__2064_,data_stage_3__2063_,data_stage_3__2062_,data_stage_3__2061_,
  data_stage_3__2060_,data_stage_3__2059_,data_stage_3__2058_,data_stage_3__2057_,
  data_stage_3__2056_,data_stage_3__2055_,data_stage_3__2054_,data_stage_3__2053_,
  data_stage_3__2052_,data_stage_3__2051_,data_stage_3__2050_,data_stage_3__2049_,
  data_stage_3__2048_,data_stage_3__2047_,data_stage_3__2046_,data_stage_3__2045_,
  data_stage_3__2044_,data_stage_3__2043_,data_stage_3__2042_,data_stage_3__2041_,
  data_stage_3__2040_,data_stage_3__2039_,data_stage_3__2038_,data_stage_3__2037_,
  data_stage_3__2036_,data_stage_3__2035_,data_stage_3__2034_,data_stage_3__2033_,
  data_stage_3__2032_,data_stage_3__2031_,data_stage_3__2030_,data_stage_3__2029_,
  data_stage_3__2028_,data_stage_3__2027_,data_stage_3__2026_,data_stage_3__2025_,
  data_stage_3__2024_,data_stage_3__2023_,data_stage_3__2022_,data_stage_3__2021_,
  data_stage_3__2020_,data_stage_3__2019_,data_stage_3__2018_,data_stage_3__2017_,
  data_stage_3__2016_,data_stage_3__2015_,data_stage_3__2014_,data_stage_3__2013_,
  data_stage_3__2012_,data_stage_3__2011_,data_stage_3__2010_,data_stage_3__2009_,
  data_stage_3__2008_,data_stage_3__2007_,data_stage_3__2006_,data_stage_3__2005_,
  data_stage_3__2004_,data_stage_3__2003_,data_stage_3__2002_,data_stage_3__2001_,
  data_stage_3__2000_,data_stage_3__1999_,data_stage_3__1998_,data_stage_3__1997_,
  data_stage_3__1996_,data_stage_3__1995_,data_stage_3__1994_,data_stage_3__1993_,
  data_stage_3__1992_,data_stage_3__1991_,data_stage_3__1990_,data_stage_3__1989_,
  data_stage_3__1988_,data_stage_3__1987_,data_stage_3__1986_,data_stage_3__1985_,
  data_stage_3__1984_,data_stage_3__1983_,data_stage_3__1982_,data_stage_3__1981_,
  data_stage_3__1980_,data_stage_3__1979_,data_stage_3__1978_,data_stage_3__1977_,
  data_stage_3__1976_,data_stage_3__1975_,data_stage_3__1974_,data_stage_3__1973_,
  data_stage_3__1972_,data_stage_3__1971_,data_stage_3__1970_,data_stage_3__1969_,
  data_stage_3__1968_,data_stage_3__1967_,data_stage_3__1966_,data_stage_3__1965_,
  data_stage_3__1964_,data_stage_3__1963_,data_stage_3__1962_,data_stage_3__1961_,
  data_stage_3__1960_,data_stage_3__1959_,data_stage_3__1958_,data_stage_3__1957_,
  data_stage_3__1956_,data_stage_3__1955_,data_stage_3__1954_,data_stage_3__1953_,
  data_stage_3__1952_,data_stage_3__1951_,data_stage_3__1950_,data_stage_3__1949_,
  data_stage_3__1948_,data_stage_3__1947_,data_stage_3__1946_,data_stage_3__1945_,
  data_stage_3__1944_,data_stage_3__1943_,data_stage_3__1942_,data_stage_3__1941_,
  data_stage_3__1940_,data_stage_3__1939_,data_stage_3__1938_,data_stage_3__1937_,
  data_stage_3__1936_,data_stage_3__1935_,data_stage_3__1934_,data_stage_3__1933_,
  data_stage_3__1932_,data_stage_3__1931_,data_stage_3__1930_,data_stage_3__1929_,
  data_stage_3__1928_,data_stage_3__1927_,data_stage_3__1926_,data_stage_3__1925_,
  data_stage_3__1924_,data_stage_3__1923_,data_stage_3__1922_,data_stage_3__1921_,
  data_stage_3__1920_,data_stage_3__1919_,data_stage_3__1918_,data_stage_3__1917_,
  data_stage_3__1916_,data_stage_3__1915_,data_stage_3__1914_,data_stage_3__1913_,
  data_stage_3__1912_,data_stage_3__1911_,data_stage_3__1910_,data_stage_3__1909_,
  data_stage_3__1908_,data_stage_3__1907_,data_stage_3__1906_,data_stage_3__1905_,
  data_stage_3__1904_,data_stage_3__1903_,data_stage_3__1902_,data_stage_3__1901_,
  data_stage_3__1900_,data_stage_3__1899_,data_stage_3__1898_,data_stage_3__1897_,
  data_stage_3__1896_,data_stage_3__1895_,data_stage_3__1894_,data_stage_3__1893_,
  data_stage_3__1892_,data_stage_3__1891_,data_stage_3__1890_,data_stage_3__1889_,
  data_stage_3__1888_,data_stage_3__1887_,data_stage_3__1886_,data_stage_3__1885_,
  data_stage_3__1884_,data_stage_3__1883_,data_stage_3__1882_,data_stage_3__1881_,
  data_stage_3__1880_,data_stage_3__1879_,data_stage_3__1878_,data_stage_3__1877_,
  data_stage_3__1876_,data_stage_3__1875_,data_stage_3__1874_,data_stage_3__1873_,
  data_stage_3__1872_,data_stage_3__1871_,data_stage_3__1870_,data_stage_3__1869_,
  data_stage_3__1868_,data_stage_3__1867_,data_stage_3__1866_,data_stage_3__1865_,
  data_stage_3__1864_,data_stage_3__1863_,data_stage_3__1862_,data_stage_3__1861_,
  data_stage_3__1860_,data_stage_3__1859_,data_stage_3__1858_,data_stage_3__1857_,
  data_stage_3__1856_,data_stage_3__1855_,data_stage_3__1854_,data_stage_3__1853_,
  data_stage_3__1852_,data_stage_3__1851_,data_stage_3__1850_,data_stage_3__1849_,
  data_stage_3__1848_,data_stage_3__1847_,data_stage_3__1846_,data_stage_3__1845_,
  data_stage_3__1844_,data_stage_3__1843_,data_stage_3__1842_,data_stage_3__1841_,
  data_stage_3__1840_,data_stage_3__1839_,data_stage_3__1838_,data_stage_3__1837_,
  data_stage_3__1836_,data_stage_3__1835_,data_stage_3__1834_,data_stage_3__1833_,
  data_stage_3__1832_,data_stage_3__1831_,data_stage_3__1830_,data_stage_3__1829_,
  data_stage_3__1828_,data_stage_3__1827_,data_stage_3__1826_,data_stage_3__1825_,
  data_stage_3__1824_,data_stage_3__1823_,data_stage_3__1822_,data_stage_3__1821_,
  data_stage_3__1820_,data_stage_3__1819_,data_stage_3__1818_,data_stage_3__1817_,
  data_stage_3__1816_,data_stage_3__1815_,data_stage_3__1814_,data_stage_3__1813_,
  data_stage_3__1812_,data_stage_3__1811_,data_stage_3__1810_,data_stage_3__1809_,
  data_stage_3__1808_,data_stage_3__1807_,data_stage_3__1806_,data_stage_3__1805_,
  data_stage_3__1804_,data_stage_3__1803_,data_stage_3__1802_,data_stage_3__1801_,
  data_stage_3__1800_,data_stage_3__1799_,data_stage_3__1798_,data_stage_3__1797_,
  data_stage_3__1796_,data_stage_3__1795_,data_stage_3__1794_,data_stage_3__1793_,
  data_stage_3__1792_,data_stage_3__1791_,data_stage_3__1790_,data_stage_3__1789_,
  data_stage_3__1788_,data_stage_3__1787_,data_stage_3__1786_,data_stage_3__1785_,
  data_stage_3__1784_,data_stage_3__1783_,data_stage_3__1782_,data_stage_3__1781_,
  data_stage_3__1780_,data_stage_3__1779_,data_stage_3__1778_,data_stage_3__1777_,
  data_stage_3__1776_,data_stage_3__1775_,data_stage_3__1774_,data_stage_3__1773_,
  data_stage_3__1772_,data_stage_3__1771_,data_stage_3__1770_,data_stage_3__1769_,
  data_stage_3__1768_,data_stage_3__1767_,data_stage_3__1766_,data_stage_3__1765_,
  data_stage_3__1764_,data_stage_3__1763_,data_stage_3__1762_,data_stage_3__1761_,
  data_stage_3__1760_,data_stage_3__1759_,data_stage_3__1758_,data_stage_3__1757_,
  data_stage_3__1756_,data_stage_3__1755_,data_stage_3__1754_,data_stage_3__1753_,
  data_stage_3__1752_,data_stage_3__1751_,data_stage_3__1750_,data_stage_3__1749_,
  data_stage_3__1748_,data_stage_3__1747_,data_stage_3__1746_,data_stage_3__1745_,
  data_stage_3__1744_,data_stage_3__1743_,data_stage_3__1742_,data_stage_3__1741_,
  data_stage_3__1740_,data_stage_3__1739_,data_stage_3__1738_,data_stage_3__1737_,
  data_stage_3__1736_,data_stage_3__1735_,data_stage_3__1734_,data_stage_3__1733_,
  data_stage_3__1732_,data_stage_3__1731_,data_stage_3__1730_,data_stage_3__1729_,
  data_stage_3__1728_,data_stage_3__1727_,data_stage_3__1726_,data_stage_3__1725_,
  data_stage_3__1724_,data_stage_3__1723_,data_stage_3__1722_,data_stage_3__1721_,
  data_stage_3__1720_,data_stage_3__1719_,data_stage_3__1718_,data_stage_3__1717_,
  data_stage_3__1716_,data_stage_3__1715_,data_stage_3__1714_,data_stage_3__1713_,
  data_stage_3__1712_,data_stage_3__1711_,data_stage_3__1710_,data_stage_3__1709_,
  data_stage_3__1708_,data_stage_3__1707_,data_stage_3__1706_,data_stage_3__1705_,
  data_stage_3__1704_,data_stage_3__1703_,data_stage_3__1702_,data_stage_3__1701_,
  data_stage_3__1700_,data_stage_3__1699_,data_stage_3__1698_,data_stage_3__1697_,
  data_stage_3__1696_,data_stage_3__1695_,data_stage_3__1694_,data_stage_3__1693_,
  data_stage_3__1692_,data_stage_3__1691_,data_stage_3__1690_,data_stage_3__1689_,
  data_stage_3__1688_,data_stage_3__1687_,data_stage_3__1686_,data_stage_3__1685_,
  data_stage_3__1684_,data_stage_3__1683_,data_stage_3__1682_,data_stage_3__1681_,
  data_stage_3__1680_,data_stage_3__1679_,data_stage_3__1678_,data_stage_3__1677_,
  data_stage_3__1676_,data_stage_3__1675_,data_stage_3__1674_,data_stage_3__1673_,
  data_stage_3__1672_,data_stage_3__1671_,data_stage_3__1670_,data_stage_3__1669_,
  data_stage_3__1668_,data_stage_3__1667_,data_stage_3__1666_,data_stage_3__1665_,
  data_stage_3__1664_,data_stage_3__1663_,data_stage_3__1662_,data_stage_3__1661_,
  data_stage_3__1660_,data_stage_3__1659_,data_stage_3__1658_,data_stage_3__1657_,
  data_stage_3__1656_,data_stage_3__1655_,data_stage_3__1654_,data_stage_3__1653_,
  data_stage_3__1652_,data_stage_3__1651_,data_stage_3__1650_,data_stage_3__1649_,
  data_stage_3__1648_,data_stage_3__1647_,data_stage_3__1646_,data_stage_3__1645_,
  data_stage_3__1644_,data_stage_3__1643_,data_stage_3__1642_,data_stage_3__1641_,
  data_stage_3__1640_,data_stage_3__1639_,data_stage_3__1638_,data_stage_3__1637_,
  data_stage_3__1636_,data_stage_3__1635_,data_stage_3__1634_,data_stage_3__1633_,
  data_stage_3__1632_,data_stage_3__1631_,data_stage_3__1630_,data_stage_3__1629_,
  data_stage_3__1628_,data_stage_3__1627_,data_stage_3__1626_,data_stage_3__1625_,
  data_stage_3__1624_,data_stage_3__1623_,data_stage_3__1622_,data_stage_3__1621_,
  data_stage_3__1620_,data_stage_3__1619_,data_stage_3__1618_,data_stage_3__1617_,
  data_stage_3__1616_,data_stage_3__1615_,data_stage_3__1614_,data_stage_3__1613_,
  data_stage_3__1612_,data_stage_3__1611_,data_stage_3__1610_,data_stage_3__1609_,
  data_stage_3__1608_,data_stage_3__1607_,data_stage_3__1606_,data_stage_3__1605_,
  data_stage_3__1604_,data_stage_3__1603_,data_stage_3__1602_,data_stage_3__1601_,
  data_stage_3__1600_,data_stage_3__1599_,data_stage_3__1598_,data_stage_3__1597_,
  data_stage_3__1596_,data_stage_3__1595_,data_stage_3__1594_,data_stage_3__1593_,
  data_stage_3__1592_,data_stage_3__1591_,data_stage_3__1590_,data_stage_3__1589_,
  data_stage_3__1588_,data_stage_3__1587_,data_stage_3__1586_,data_stage_3__1585_,
  data_stage_3__1584_,data_stage_3__1583_,data_stage_3__1582_,data_stage_3__1581_,
  data_stage_3__1580_,data_stage_3__1579_,data_stage_3__1578_,data_stage_3__1577_,
  data_stage_3__1576_,data_stage_3__1575_,data_stage_3__1574_,data_stage_3__1573_,
  data_stage_3__1572_,data_stage_3__1571_,data_stage_3__1570_,data_stage_3__1569_,
  data_stage_3__1568_,data_stage_3__1567_,data_stage_3__1566_,data_stage_3__1565_,
  data_stage_3__1564_,data_stage_3__1563_,data_stage_3__1562_,data_stage_3__1561_,
  data_stage_3__1560_,data_stage_3__1559_,data_stage_3__1558_,data_stage_3__1557_,
  data_stage_3__1556_,data_stage_3__1555_,data_stage_3__1554_,data_stage_3__1553_,
  data_stage_3__1552_,data_stage_3__1551_,data_stage_3__1550_,data_stage_3__1549_,
  data_stage_3__1548_,data_stage_3__1547_,data_stage_3__1546_,data_stage_3__1545_,
  data_stage_3__1544_,data_stage_3__1543_,data_stage_3__1542_,data_stage_3__1541_,
  data_stage_3__1540_,data_stage_3__1539_,data_stage_3__1538_,data_stage_3__1537_,
  data_stage_3__1536_,data_stage_3__1535_,data_stage_3__1534_,data_stage_3__1533_,
  data_stage_3__1532_,data_stage_3__1531_,data_stage_3__1530_,data_stage_3__1529_,
  data_stage_3__1528_,data_stage_3__1527_,data_stage_3__1526_,data_stage_3__1525_,
  data_stage_3__1524_,data_stage_3__1523_,data_stage_3__1522_,data_stage_3__1521_,
  data_stage_3__1520_,data_stage_3__1519_,data_stage_3__1518_,data_stage_3__1517_,
  data_stage_3__1516_,data_stage_3__1515_,data_stage_3__1514_,data_stage_3__1513_,
  data_stage_3__1512_,data_stage_3__1511_,data_stage_3__1510_,data_stage_3__1509_,
  data_stage_3__1508_,data_stage_3__1507_,data_stage_3__1506_,data_stage_3__1505_,
  data_stage_3__1504_,data_stage_3__1503_,data_stage_3__1502_,data_stage_3__1501_,
  data_stage_3__1500_,data_stage_3__1499_,data_stage_3__1498_,data_stage_3__1497_,
  data_stage_3__1496_,data_stage_3__1495_,data_stage_3__1494_,data_stage_3__1493_,
  data_stage_3__1492_,data_stage_3__1491_,data_stage_3__1490_,data_stage_3__1489_,
  data_stage_3__1488_,data_stage_3__1487_,data_stage_3__1486_,data_stage_3__1485_,
  data_stage_3__1484_,data_stage_3__1483_,data_stage_3__1482_,data_stage_3__1481_,
  data_stage_3__1480_,data_stage_3__1479_,data_stage_3__1478_,data_stage_3__1477_,
  data_stage_3__1476_,data_stage_3__1475_,data_stage_3__1474_,data_stage_3__1473_,
  data_stage_3__1472_,data_stage_3__1471_,data_stage_3__1470_,data_stage_3__1469_,
  data_stage_3__1468_,data_stage_3__1467_,data_stage_3__1466_,data_stage_3__1465_,
  data_stage_3__1464_,data_stage_3__1463_,data_stage_3__1462_,data_stage_3__1461_,
  data_stage_3__1460_,data_stage_3__1459_,data_stage_3__1458_,data_stage_3__1457_,
  data_stage_3__1456_,data_stage_3__1455_,data_stage_3__1454_,data_stage_3__1453_,
  data_stage_3__1452_,data_stage_3__1451_,data_stage_3__1450_,data_stage_3__1449_,
  data_stage_3__1448_,data_stage_3__1447_,data_stage_3__1446_,data_stage_3__1445_,
  data_stage_3__1444_,data_stage_3__1443_,data_stage_3__1442_,data_stage_3__1441_,
  data_stage_3__1440_,data_stage_3__1439_,data_stage_3__1438_,data_stage_3__1437_,
  data_stage_3__1436_,data_stage_3__1435_,data_stage_3__1434_,data_stage_3__1433_,
  data_stage_3__1432_,data_stage_3__1431_,data_stage_3__1430_,data_stage_3__1429_,
  data_stage_3__1428_,data_stage_3__1427_,data_stage_3__1426_,data_stage_3__1425_,
  data_stage_3__1424_,data_stage_3__1423_,data_stage_3__1422_,data_stage_3__1421_,
  data_stage_3__1420_,data_stage_3__1419_,data_stage_3__1418_,data_stage_3__1417_,
  data_stage_3__1416_,data_stage_3__1415_,data_stage_3__1414_,data_stage_3__1413_,
  data_stage_3__1412_,data_stage_3__1411_,data_stage_3__1410_,data_stage_3__1409_,
  data_stage_3__1408_,data_stage_3__1407_,data_stage_3__1406_,data_stage_3__1405_,
  data_stage_3__1404_,data_stage_3__1403_,data_stage_3__1402_,data_stage_3__1401_,
  data_stage_3__1400_,data_stage_3__1399_,data_stage_3__1398_,data_stage_3__1397_,
  data_stage_3__1396_,data_stage_3__1395_,data_stage_3__1394_,data_stage_3__1393_,
  data_stage_3__1392_,data_stage_3__1391_,data_stage_3__1390_,data_stage_3__1389_,
  data_stage_3__1388_,data_stage_3__1387_,data_stage_3__1386_,data_stage_3__1385_,
  data_stage_3__1384_,data_stage_3__1383_,data_stage_3__1382_,data_stage_3__1381_,
  data_stage_3__1380_,data_stage_3__1379_,data_stage_3__1378_,data_stage_3__1377_,
  data_stage_3__1376_,data_stage_3__1375_,data_stage_3__1374_,data_stage_3__1373_,
  data_stage_3__1372_,data_stage_3__1371_,data_stage_3__1370_,data_stage_3__1369_,
  data_stage_3__1368_,data_stage_3__1367_,data_stage_3__1366_,data_stage_3__1365_,
  data_stage_3__1364_,data_stage_3__1363_,data_stage_3__1362_,data_stage_3__1361_,
  data_stage_3__1360_,data_stage_3__1359_,data_stage_3__1358_,data_stage_3__1357_,
  data_stage_3__1356_,data_stage_3__1355_,data_stage_3__1354_,data_stage_3__1353_,
  data_stage_3__1352_,data_stage_3__1351_,data_stage_3__1350_,data_stage_3__1349_,
  data_stage_3__1348_,data_stage_3__1347_,data_stage_3__1346_,data_stage_3__1345_,
  data_stage_3__1344_,data_stage_3__1343_,data_stage_3__1342_,data_stage_3__1341_,
  data_stage_3__1340_,data_stage_3__1339_,data_stage_3__1338_,data_stage_3__1337_,
  data_stage_3__1336_,data_stage_3__1335_,data_stage_3__1334_,data_stage_3__1333_,
  data_stage_3__1332_,data_stage_3__1331_,data_stage_3__1330_,data_stage_3__1329_,
  data_stage_3__1328_,data_stage_3__1327_,data_stage_3__1326_,data_stage_3__1325_,
  data_stage_3__1324_,data_stage_3__1323_,data_stage_3__1322_,data_stage_3__1321_,
  data_stage_3__1320_,data_stage_3__1319_,data_stage_3__1318_,data_stage_3__1317_,
  data_stage_3__1316_,data_stage_3__1315_,data_stage_3__1314_,data_stage_3__1313_,
  data_stage_3__1312_,data_stage_3__1311_,data_stage_3__1310_,data_stage_3__1309_,
  data_stage_3__1308_,data_stage_3__1307_,data_stage_3__1306_,data_stage_3__1305_,
  data_stage_3__1304_,data_stage_3__1303_,data_stage_3__1302_,data_stage_3__1301_,
  data_stage_3__1300_,data_stage_3__1299_,data_stage_3__1298_,data_stage_3__1297_,
  data_stage_3__1296_,data_stage_3__1295_,data_stage_3__1294_,data_stage_3__1293_,
  data_stage_3__1292_,data_stage_3__1291_,data_stage_3__1290_,data_stage_3__1289_,
  data_stage_3__1288_,data_stage_3__1287_,data_stage_3__1286_,data_stage_3__1285_,
  data_stage_3__1284_,data_stage_3__1283_,data_stage_3__1282_,data_stage_3__1281_,
  data_stage_3__1280_,data_stage_3__1279_,data_stage_3__1278_,data_stage_3__1277_,
  data_stage_3__1276_,data_stage_3__1275_,data_stage_3__1274_,data_stage_3__1273_,
  data_stage_3__1272_,data_stage_3__1271_,data_stage_3__1270_,data_stage_3__1269_,
  data_stage_3__1268_,data_stage_3__1267_,data_stage_3__1266_,data_stage_3__1265_,
  data_stage_3__1264_,data_stage_3__1263_,data_stage_3__1262_,data_stage_3__1261_,
  data_stage_3__1260_,data_stage_3__1259_,data_stage_3__1258_,data_stage_3__1257_,
  data_stage_3__1256_,data_stage_3__1255_,data_stage_3__1254_,data_stage_3__1253_,
  data_stage_3__1252_,data_stage_3__1251_,data_stage_3__1250_,data_stage_3__1249_,
  data_stage_3__1248_,data_stage_3__1247_,data_stage_3__1246_,data_stage_3__1245_,
  data_stage_3__1244_,data_stage_3__1243_,data_stage_3__1242_,data_stage_3__1241_,
  data_stage_3__1240_,data_stage_3__1239_,data_stage_3__1238_,data_stage_3__1237_,
  data_stage_3__1236_,data_stage_3__1235_,data_stage_3__1234_,data_stage_3__1233_,
  data_stage_3__1232_,data_stage_3__1231_,data_stage_3__1230_,data_stage_3__1229_,
  data_stage_3__1228_,data_stage_3__1227_,data_stage_3__1226_,data_stage_3__1225_,
  data_stage_3__1224_,data_stage_3__1223_,data_stage_3__1222_,data_stage_3__1221_,
  data_stage_3__1220_,data_stage_3__1219_,data_stage_3__1218_,data_stage_3__1217_,
  data_stage_3__1216_,data_stage_3__1215_,data_stage_3__1214_,data_stage_3__1213_,
  data_stage_3__1212_,data_stage_3__1211_,data_stage_3__1210_,data_stage_3__1209_,
  data_stage_3__1208_,data_stage_3__1207_,data_stage_3__1206_,data_stage_3__1205_,
  data_stage_3__1204_,data_stage_3__1203_,data_stage_3__1202_,data_stage_3__1201_,
  data_stage_3__1200_,data_stage_3__1199_,data_stage_3__1198_,data_stage_3__1197_,
  data_stage_3__1196_,data_stage_3__1195_,data_stage_3__1194_,data_stage_3__1193_,
  data_stage_3__1192_,data_stage_3__1191_,data_stage_3__1190_,data_stage_3__1189_,
  data_stage_3__1188_,data_stage_3__1187_,data_stage_3__1186_,data_stage_3__1185_,
  data_stage_3__1184_,data_stage_3__1183_,data_stage_3__1182_,data_stage_3__1181_,
  data_stage_3__1180_,data_stage_3__1179_,data_stage_3__1178_,data_stage_3__1177_,
  data_stage_3__1176_,data_stage_3__1175_,data_stage_3__1174_,data_stage_3__1173_,
  data_stage_3__1172_,data_stage_3__1171_,data_stage_3__1170_,data_stage_3__1169_,
  data_stage_3__1168_,data_stage_3__1167_,data_stage_3__1166_,data_stage_3__1165_,
  data_stage_3__1164_,data_stage_3__1163_,data_stage_3__1162_,data_stage_3__1161_,
  data_stage_3__1160_,data_stage_3__1159_,data_stage_3__1158_,data_stage_3__1157_,
  data_stage_3__1156_,data_stage_3__1155_,data_stage_3__1154_,data_stage_3__1153_,
  data_stage_3__1152_,data_stage_3__1151_,data_stage_3__1150_,data_stage_3__1149_,
  data_stage_3__1148_,data_stage_3__1147_,data_stage_3__1146_,data_stage_3__1145_,
  data_stage_3__1144_,data_stage_3__1143_,data_stage_3__1142_,data_stage_3__1141_,
  data_stage_3__1140_,data_stage_3__1139_,data_stage_3__1138_,data_stage_3__1137_,
  data_stage_3__1136_,data_stage_3__1135_,data_stage_3__1134_,data_stage_3__1133_,
  data_stage_3__1132_,data_stage_3__1131_,data_stage_3__1130_,data_stage_3__1129_,
  data_stage_3__1128_,data_stage_3__1127_,data_stage_3__1126_,data_stage_3__1125_,
  data_stage_3__1124_,data_stage_3__1123_,data_stage_3__1122_,data_stage_3__1121_,
  data_stage_3__1120_,data_stage_3__1119_,data_stage_3__1118_,data_stage_3__1117_,
  data_stage_3__1116_,data_stage_3__1115_,data_stage_3__1114_,data_stage_3__1113_,
  data_stage_3__1112_,data_stage_3__1111_,data_stage_3__1110_,data_stage_3__1109_,
  data_stage_3__1108_,data_stage_3__1107_,data_stage_3__1106_,data_stage_3__1105_,
  data_stage_3__1104_,data_stage_3__1103_,data_stage_3__1102_,data_stage_3__1101_,
  data_stage_3__1100_,data_stage_3__1099_,data_stage_3__1098_,data_stage_3__1097_,
  data_stage_3__1096_,data_stage_3__1095_,data_stage_3__1094_,data_stage_3__1093_,
  data_stage_3__1092_,data_stage_3__1091_,data_stage_3__1090_,data_stage_3__1089_,
  data_stage_3__1088_,data_stage_3__1087_,data_stage_3__1086_,data_stage_3__1085_,
  data_stage_3__1084_,data_stage_3__1083_,data_stage_3__1082_,data_stage_3__1081_,
  data_stage_3__1080_,data_stage_3__1079_,data_stage_3__1078_,data_stage_3__1077_,
  data_stage_3__1076_,data_stage_3__1075_,data_stage_3__1074_,data_stage_3__1073_,
  data_stage_3__1072_,data_stage_3__1071_,data_stage_3__1070_,data_stage_3__1069_,
  data_stage_3__1068_,data_stage_3__1067_,data_stage_3__1066_,data_stage_3__1065_,
  data_stage_3__1064_,data_stage_3__1063_,data_stage_3__1062_,data_stage_3__1061_,
  data_stage_3__1060_,data_stage_3__1059_,data_stage_3__1058_,data_stage_3__1057_,
  data_stage_3__1056_,data_stage_3__1055_,data_stage_3__1054_,data_stage_3__1053_,
  data_stage_3__1052_,data_stage_3__1051_,data_stage_3__1050_,data_stage_3__1049_,
  data_stage_3__1048_,data_stage_3__1047_,data_stage_3__1046_,data_stage_3__1045_,
  data_stage_3__1044_,data_stage_3__1043_,data_stage_3__1042_,data_stage_3__1041_,
  data_stage_3__1040_,data_stage_3__1039_,data_stage_3__1038_,data_stage_3__1037_,
  data_stage_3__1036_,data_stage_3__1035_,data_stage_3__1034_,data_stage_3__1033_,
  data_stage_3__1032_,data_stage_3__1031_,data_stage_3__1030_,data_stage_3__1029_,
  data_stage_3__1028_,data_stage_3__1027_,data_stage_3__1026_,data_stage_3__1025_,
  data_stage_3__1024_,data_stage_3__1023_,data_stage_3__1022_,data_stage_3__1021_,
  data_stage_3__1020_,data_stage_3__1019_,data_stage_3__1018_,data_stage_3__1017_,
  data_stage_3__1016_,data_stage_3__1015_,data_stage_3__1014_,data_stage_3__1013_,
  data_stage_3__1012_,data_stage_3__1011_,data_stage_3__1010_,data_stage_3__1009_,
  data_stage_3__1008_,data_stage_3__1007_,data_stage_3__1006_,data_stage_3__1005_,
  data_stage_3__1004_,data_stage_3__1003_,data_stage_3__1002_,data_stage_3__1001_,
  data_stage_3__1000_,data_stage_3__999_,data_stage_3__998_,data_stage_3__997_,
  data_stage_3__996_,data_stage_3__995_,data_stage_3__994_,data_stage_3__993_,
  data_stage_3__992_,data_stage_3__991_,data_stage_3__990_,data_stage_3__989_,
  data_stage_3__988_,data_stage_3__987_,data_stage_3__986_,data_stage_3__985_,
  data_stage_3__984_,data_stage_3__983_,data_stage_3__982_,data_stage_3__981_,data_stage_3__980_,
  data_stage_3__979_,data_stage_3__978_,data_stage_3__977_,data_stage_3__976_,
  data_stage_3__975_,data_stage_3__974_,data_stage_3__973_,data_stage_3__972_,
  data_stage_3__971_,data_stage_3__970_,data_stage_3__969_,data_stage_3__968_,
  data_stage_3__967_,data_stage_3__966_,data_stage_3__965_,data_stage_3__964_,
  data_stage_3__963_,data_stage_3__962_,data_stage_3__961_,data_stage_3__960_,data_stage_3__959_,
  data_stage_3__958_,data_stage_3__957_,data_stage_3__956_,data_stage_3__955_,
  data_stage_3__954_,data_stage_3__953_,data_stage_3__952_,data_stage_3__951_,
  data_stage_3__950_,data_stage_3__949_,data_stage_3__948_,data_stage_3__947_,
  data_stage_3__946_,data_stage_3__945_,data_stage_3__944_,data_stage_3__943_,
  data_stage_3__942_,data_stage_3__941_,data_stage_3__940_,data_stage_3__939_,data_stage_3__938_,
  data_stage_3__937_,data_stage_3__936_,data_stage_3__935_,data_stage_3__934_,
  data_stage_3__933_,data_stage_3__932_,data_stage_3__931_,data_stage_3__930_,
  data_stage_3__929_,data_stage_3__928_,data_stage_3__927_,data_stage_3__926_,
  data_stage_3__925_,data_stage_3__924_,data_stage_3__923_,data_stage_3__922_,
  data_stage_3__921_,data_stage_3__920_,data_stage_3__919_,data_stage_3__918_,data_stage_3__917_,
  data_stage_3__916_,data_stage_3__915_,data_stage_3__914_,data_stage_3__913_,
  data_stage_3__912_,data_stage_3__911_,data_stage_3__910_,data_stage_3__909_,
  data_stage_3__908_,data_stage_3__907_,data_stage_3__906_,data_stage_3__905_,
  data_stage_3__904_,data_stage_3__903_,data_stage_3__902_,data_stage_3__901_,data_stage_3__900_,
  data_stage_3__899_,data_stage_3__898_,data_stage_3__897_,data_stage_3__896_,
  data_stage_3__895_,data_stage_3__894_,data_stage_3__893_,data_stage_3__892_,
  data_stage_3__891_,data_stage_3__890_,data_stage_3__889_,data_stage_3__888_,
  data_stage_3__887_,data_stage_3__886_,data_stage_3__885_,data_stage_3__884_,
  data_stage_3__883_,data_stage_3__882_,data_stage_3__881_,data_stage_3__880_,data_stage_3__879_,
  data_stage_3__878_,data_stage_3__877_,data_stage_3__876_,data_stage_3__875_,
  data_stage_3__874_,data_stage_3__873_,data_stage_3__872_,data_stage_3__871_,
  data_stage_3__870_,data_stage_3__869_,data_stage_3__868_,data_stage_3__867_,
  data_stage_3__866_,data_stage_3__865_,data_stage_3__864_,data_stage_3__863_,
  data_stage_3__862_,data_stage_3__861_,data_stage_3__860_,data_stage_3__859_,data_stage_3__858_,
  data_stage_3__857_,data_stage_3__856_,data_stage_3__855_,data_stage_3__854_,
  data_stage_3__853_,data_stage_3__852_,data_stage_3__851_,data_stage_3__850_,
  data_stage_3__849_,data_stage_3__848_,data_stage_3__847_,data_stage_3__846_,
  data_stage_3__845_,data_stage_3__844_,data_stage_3__843_,data_stage_3__842_,
  data_stage_3__841_,data_stage_3__840_,data_stage_3__839_,data_stage_3__838_,data_stage_3__837_,
  data_stage_3__836_,data_stage_3__835_,data_stage_3__834_,data_stage_3__833_,
  data_stage_3__832_,data_stage_3__831_,data_stage_3__830_,data_stage_3__829_,
  data_stage_3__828_,data_stage_3__827_,data_stage_3__826_,data_stage_3__825_,
  data_stage_3__824_,data_stage_3__823_,data_stage_3__822_,data_stage_3__821_,data_stage_3__820_,
  data_stage_3__819_,data_stage_3__818_,data_stage_3__817_,data_stage_3__816_,
  data_stage_3__815_,data_stage_3__814_,data_stage_3__813_,data_stage_3__812_,
  data_stage_3__811_,data_stage_3__810_,data_stage_3__809_,data_stage_3__808_,
  data_stage_3__807_,data_stage_3__806_,data_stage_3__805_,data_stage_3__804_,
  data_stage_3__803_,data_stage_3__802_,data_stage_3__801_,data_stage_3__800_,data_stage_3__799_,
  data_stage_3__798_,data_stage_3__797_,data_stage_3__796_,data_stage_3__795_,
  data_stage_3__794_,data_stage_3__793_,data_stage_3__792_,data_stage_3__791_,
  data_stage_3__790_,data_stage_3__789_,data_stage_3__788_,data_stage_3__787_,
  data_stage_3__786_,data_stage_3__785_,data_stage_3__784_,data_stage_3__783_,
  data_stage_3__782_,data_stage_3__781_,data_stage_3__780_,data_stage_3__779_,data_stage_3__778_,
  data_stage_3__777_,data_stage_3__776_,data_stage_3__775_,data_stage_3__774_,
  data_stage_3__773_,data_stage_3__772_,data_stage_3__771_,data_stage_3__770_,
  data_stage_3__769_,data_stage_3__768_,data_stage_3__767_,data_stage_3__766_,
  data_stage_3__765_,data_stage_3__764_,data_stage_3__763_,data_stage_3__762_,
  data_stage_3__761_,data_stage_3__760_,data_stage_3__759_,data_stage_3__758_,data_stage_3__757_,
  data_stage_3__756_,data_stage_3__755_,data_stage_3__754_,data_stage_3__753_,
  data_stage_3__752_,data_stage_3__751_,data_stage_3__750_,data_stage_3__749_,
  data_stage_3__748_,data_stage_3__747_,data_stage_3__746_,data_stage_3__745_,
  data_stage_3__744_,data_stage_3__743_,data_stage_3__742_,data_stage_3__741_,data_stage_3__740_,
  data_stage_3__739_,data_stage_3__738_,data_stage_3__737_,data_stage_3__736_,
  data_stage_3__735_,data_stage_3__734_,data_stage_3__733_,data_stage_3__732_,
  data_stage_3__731_,data_stage_3__730_,data_stage_3__729_,data_stage_3__728_,
  data_stage_3__727_,data_stage_3__726_,data_stage_3__725_,data_stage_3__724_,
  data_stage_3__723_,data_stage_3__722_,data_stage_3__721_,data_stage_3__720_,data_stage_3__719_,
  data_stage_3__718_,data_stage_3__717_,data_stage_3__716_,data_stage_3__715_,
  data_stage_3__714_,data_stage_3__713_,data_stage_3__712_,data_stage_3__711_,
  data_stage_3__710_,data_stage_3__709_,data_stage_3__708_,data_stage_3__707_,
  data_stage_3__706_,data_stage_3__705_,data_stage_3__704_,data_stage_3__703_,
  data_stage_3__702_,data_stage_3__701_,data_stage_3__700_,data_stage_3__699_,data_stage_3__698_,
  data_stage_3__697_,data_stage_3__696_,data_stage_3__695_,data_stage_3__694_,
  data_stage_3__693_,data_stage_3__692_,data_stage_3__691_,data_stage_3__690_,
  data_stage_3__689_,data_stage_3__688_,data_stage_3__687_,data_stage_3__686_,
  data_stage_3__685_,data_stage_3__684_,data_stage_3__683_,data_stage_3__682_,
  data_stage_3__681_,data_stage_3__680_,data_stage_3__679_,data_stage_3__678_,data_stage_3__677_,
  data_stage_3__676_,data_stage_3__675_,data_stage_3__674_,data_stage_3__673_,
  data_stage_3__672_,data_stage_3__671_,data_stage_3__670_,data_stage_3__669_,
  data_stage_3__668_,data_stage_3__667_,data_stage_3__666_,data_stage_3__665_,
  data_stage_3__664_,data_stage_3__663_,data_stage_3__662_,data_stage_3__661_,data_stage_3__660_,
  data_stage_3__659_,data_stage_3__658_,data_stage_3__657_,data_stage_3__656_,
  data_stage_3__655_,data_stage_3__654_,data_stage_3__653_,data_stage_3__652_,
  data_stage_3__651_,data_stage_3__650_,data_stage_3__649_,data_stage_3__648_,
  data_stage_3__647_,data_stage_3__646_,data_stage_3__645_,data_stage_3__644_,
  data_stage_3__643_,data_stage_3__642_,data_stage_3__641_,data_stage_3__640_,data_stage_3__639_,
  data_stage_3__638_,data_stage_3__637_,data_stage_3__636_,data_stage_3__635_,
  data_stage_3__634_,data_stage_3__633_,data_stage_3__632_,data_stage_3__631_,
  data_stage_3__630_,data_stage_3__629_,data_stage_3__628_,data_stage_3__627_,
  data_stage_3__626_,data_stage_3__625_,data_stage_3__624_,data_stage_3__623_,
  data_stage_3__622_,data_stage_3__621_,data_stage_3__620_,data_stage_3__619_,data_stage_3__618_,
  data_stage_3__617_,data_stage_3__616_,data_stage_3__615_,data_stage_3__614_,
  data_stage_3__613_,data_stage_3__612_,data_stage_3__611_,data_stage_3__610_,
  data_stage_3__609_,data_stage_3__608_,data_stage_3__607_,data_stage_3__606_,
  data_stage_3__605_,data_stage_3__604_,data_stage_3__603_,data_stage_3__602_,
  data_stage_3__601_,data_stage_3__600_,data_stage_3__599_,data_stage_3__598_,data_stage_3__597_,
  data_stage_3__596_,data_stage_3__595_,data_stage_3__594_,data_stage_3__593_,
  data_stage_3__592_,data_stage_3__591_,data_stage_3__590_,data_stage_3__589_,
  data_stage_3__588_,data_stage_3__587_,data_stage_3__586_,data_stage_3__585_,
  data_stage_3__584_,data_stage_3__583_,data_stage_3__582_,data_stage_3__581_,data_stage_3__580_,
  data_stage_3__579_,data_stage_3__578_,data_stage_3__577_,data_stage_3__576_,
  data_stage_3__575_,data_stage_3__574_,data_stage_3__573_,data_stage_3__572_,
  data_stage_3__571_,data_stage_3__570_,data_stage_3__569_,data_stage_3__568_,
  data_stage_3__567_,data_stage_3__566_,data_stage_3__565_,data_stage_3__564_,
  data_stage_3__563_,data_stage_3__562_,data_stage_3__561_,data_stage_3__560_,data_stage_3__559_,
  data_stage_3__558_,data_stage_3__557_,data_stage_3__556_,data_stage_3__555_,
  data_stage_3__554_,data_stage_3__553_,data_stage_3__552_,data_stage_3__551_,
  data_stage_3__550_,data_stage_3__549_,data_stage_3__548_,data_stage_3__547_,
  data_stage_3__546_,data_stage_3__545_,data_stage_3__544_,data_stage_3__543_,
  data_stage_3__542_,data_stage_3__541_,data_stage_3__540_,data_stage_3__539_,data_stage_3__538_,
  data_stage_3__537_,data_stage_3__536_,data_stage_3__535_,data_stage_3__534_,
  data_stage_3__533_,data_stage_3__532_,data_stage_3__531_,data_stage_3__530_,
  data_stage_3__529_,data_stage_3__528_,data_stage_3__527_,data_stage_3__526_,
  data_stage_3__525_,data_stage_3__524_,data_stage_3__523_,data_stage_3__522_,
  data_stage_3__521_,data_stage_3__520_,data_stage_3__519_,data_stage_3__518_,data_stage_3__517_,
  data_stage_3__516_,data_stage_3__515_,data_stage_3__514_,data_stage_3__513_,
  data_stage_3__512_,data_stage_3__511_,data_stage_3__510_,data_stage_3__509_,
  data_stage_3__508_,data_stage_3__507_,data_stage_3__506_,data_stage_3__505_,
  data_stage_3__504_,data_stage_3__503_,data_stage_3__502_,data_stage_3__501_,data_stage_3__500_,
  data_stage_3__499_,data_stage_3__498_,data_stage_3__497_,data_stage_3__496_,
  data_stage_3__495_,data_stage_3__494_,data_stage_3__493_,data_stage_3__492_,
  data_stage_3__491_,data_stage_3__490_,data_stage_3__489_,data_stage_3__488_,
  data_stage_3__487_,data_stage_3__486_,data_stage_3__485_,data_stage_3__484_,
  data_stage_3__483_,data_stage_3__482_,data_stage_3__481_,data_stage_3__480_,data_stage_3__479_,
  data_stage_3__478_,data_stage_3__477_,data_stage_3__476_,data_stage_3__475_,
  data_stage_3__474_,data_stage_3__473_,data_stage_3__472_,data_stage_3__471_,
  data_stage_3__470_,data_stage_3__469_,data_stage_3__468_,data_stage_3__467_,
  data_stage_3__466_,data_stage_3__465_,data_stage_3__464_,data_stage_3__463_,
  data_stage_3__462_,data_stage_3__461_,data_stage_3__460_,data_stage_3__459_,data_stage_3__458_,
  data_stage_3__457_,data_stage_3__456_,data_stage_3__455_,data_stage_3__454_,
  data_stage_3__453_,data_stage_3__452_,data_stage_3__451_,data_stage_3__450_,
  data_stage_3__449_,data_stage_3__448_,data_stage_3__447_,data_stage_3__446_,
  data_stage_3__445_,data_stage_3__444_,data_stage_3__443_,data_stage_3__442_,
  data_stage_3__441_,data_stage_3__440_,data_stage_3__439_,data_stage_3__438_,data_stage_3__437_,
  data_stage_3__436_,data_stage_3__435_,data_stage_3__434_,data_stage_3__433_,
  data_stage_3__432_,data_stage_3__431_,data_stage_3__430_,data_stage_3__429_,
  data_stage_3__428_,data_stage_3__427_,data_stage_3__426_,data_stage_3__425_,
  data_stage_3__424_,data_stage_3__423_,data_stage_3__422_,data_stage_3__421_,data_stage_3__420_,
  data_stage_3__419_,data_stage_3__418_,data_stage_3__417_,data_stage_3__416_,
  data_stage_3__415_,data_stage_3__414_,data_stage_3__413_,data_stage_3__412_,
  data_stage_3__411_,data_stage_3__410_,data_stage_3__409_,data_stage_3__408_,
  data_stage_3__407_,data_stage_3__406_,data_stage_3__405_,data_stage_3__404_,
  data_stage_3__403_,data_stage_3__402_,data_stage_3__401_,data_stage_3__400_,data_stage_3__399_,
  data_stage_3__398_,data_stage_3__397_,data_stage_3__396_,data_stage_3__395_,
  data_stage_3__394_,data_stage_3__393_,data_stage_3__392_,data_stage_3__391_,
  data_stage_3__390_,data_stage_3__389_,data_stage_3__388_,data_stage_3__387_,
  data_stage_3__386_,data_stage_3__385_,data_stage_3__384_,data_stage_3__383_,
  data_stage_3__382_,data_stage_3__381_,data_stage_3__380_,data_stage_3__379_,data_stage_3__378_,
  data_stage_3__377_,data_stage_3__376_,data_stage_3__375_,data_stage_3__374_,
  data_stage_3__373_,data_stage_3__372_,data_stage_3__371_,data_stage_3__370_,
  data_stage_3__369_,data_stage_3__368_,data_stage_3__367_,data_stage_3__366_,
  data_stage_3__365_,data_stage_3__364_,data_stage_3__363_,data_stage_3__362_,
  data_stage_3__361_,data_stage_3__360_,data_stage_3__359_,data_stage_3__358_,data_stage_3__357_,
  data_stage_3__356_,data_stage_3__355_,data_stage_3__354_,data_stage_3__353_,
  data_stage_3__352_,data_stage_3__351_,data_stage_3__350_,data_stage_3__349_,
  data_stage_3__348_,data_stage_3__347_,data_stage_3__346_,data_stage_3__345_,
  data_stage_3__344_,data_stage_3__343_,data_stage_3__342_,data_stage_3__341_,data_stage_3__340_,
  data_stage_3__339_,data_stage_3__338_,data_stage_3__337_,data_stage_3__336_,
  data_stage_3__335_,data_stage_3__334_,data_stage_3__333_,data_stage_3__332_,
  data_stage_3__331_,data_stage_3__330_,data_stage_3__329_,data_stage_3__328_,
  data_stage_3__327_,data_stage_3__326_,data_stage_3__325_,data_stage_3__324_,
  data_stage_3__323_,data_stage_3__322_,data_stage_3__321_,data_stage_3__320_,data_stage_3__319_,
  data_stage_3__318_,data_stage_3__317_,data_stage_3__316_,data_stage_3__315_,
  data_stage_3__314_,data_stage_3__313_,data_stage_3__312_,data_stage_3__311_,
  data_stage_3__310_,data_stage_3__309_,data_stage_3__308_,data_stage_3__307_,
  data_stage_3__306_,data_stage_3__305_,data_stage_3__304_,data_stage_3__303_,
  data_stage_3__302_,data_stage_3__301_,data_stage_3__300_,data_stage_3__299_,data_stage_3__298_,
  data_stage_3__297_,data_stage_3__296_,data_stage_3__295_,data_stage_3__294_,
  data_stage_3__293_,data_stage_3__292_,data_stage_3__291_,data_stage_3__290_,
  data_stage_3__289_,data_stage_3__288_,data_stage_3__287_,data_stage_3__286_,
  data_stage_3__285_,data_stage_3__284_,data_stage_3__283_,data_stage_3__282_,
  data_stage_3__281_,data_stage_3__280_,data_stage_3__279_,data_stage_3__278_,data_stage_3__277_,
  data_stage_3__276_,data_stage_3__275_,data_stage_3__274_,data_stage_3__273_,
  data_stage_3__272_,data_stage_3__271_,data_stage_3__270_,data_stage_3__269_,
  data_stage_3__268_,data_stage_3__267_,data_stage_3__266_,data_stage_3__265_,
  data_stage_3__264_,data_stage_3__263_,data_stage_3__262_,data_stage_3__261_,data_stage_3__260_,
  data_stage_3__259_,data_stage_3__258_,data_stage_3__257_,data_stage_3__256_,
  data_stage_3__255_,data_stage_3__254_,data_stage_3__253_,data_stage_3__252_,
  data_stage_3__251_,data_stage_3__250_,data_stage_3__249_,data_stage_3__248_,
  data_stage_3__247_,data_stage_3__246_,data_stage_3__245_,data_stage_3__244_,
  data_stage_3__243_,data_stage_3__242_,data_stage_3__241_,data_stage_3__240_,data_stage_3__239_,
  data_stage_3__238_,data_stage_3__237_,data_stage_3__236_,data_stage_3__235_,
  data_stage_3__234_,data_stage_3__233_,data_stage_3__232_,data_stage_3__231_,
  data_stage_3__230_,data_stage_3__229_,data_stage_3__228_,data_stage_3__227_,
  data_stage_3__226_,data_stage_3__225_,data_stage_3__224_,data_stage_3__223_,
  data_stage_3__222_,data_stage_3__221_,data_stage_3__220_,data_stage_3__219_,data_stage_3__218_,
  data_stage_3__217_,data_stage_3__216_,data_stage_3__215_,data_stage_3__214_,
  data_stage_3__213_,data_stage_3__212_,data_stage_3__211_,data_stage_3__210_,
  data_stage_3__209_,data_stage_3__208_,data_stage_3__207_,data_stage_3__206_,
  data_stage_3__205_,data_stage_3__204_,data_stage_3__203_,data_stage_3__202_,
  data_stage_3__201_,data_stage_3__200_,data_stage_3__199_,data_stage_3__198_,data_stage_3__197_,
  data_stage_3__196_,data_stage_3__195_,data_stage_3__194_,data_stage_3__193_,
  data_stage_3__192_,data_stage_3__191_,data_stage_3__190_,data_stage_3__189_,
  data_stage_3__188_,data_stage_3__187_,data_stage_3__186_,data_stage_3__185_,
  data_stage_3__184_,data_stage_3__183_,data_stage_3__182_,data_stage_3__181_,data_stage_3__180_,
  data_stage_3__179_,data_stage_3__178_,data_stage_3__177_,data_stage_3__176_,
  data_stage_3__175_,data_stage_3__174_,data_stage_3__173_,data_stage_3__172_,
  data_stage_3__171_,data_stage_3__170_,data_stage_3__169_,data_stage_3__168_,
  data_stage_3__167_,data_stage_3__166_,data_stage_3__165_,data_stage_3__164_,
  data_stage_3__163_,data_stage_3__162_,data_stage_3__161_,data_stage_3__160_,data_stage_3__159_,
  data_stage_3__158_,data_stage_3__157_,data_stage_3__156_,data_stage_3__155_,
  data_stage_3__154_,data_stage_3__153_,data_stage_3__152_,data_stage_3__151_,
  data_stage_3__150_,data_stage_3__149_,data_stage_3__148_,data_stage_3__147_,
  data_stage_3__146_,data_stage_3__145_,data_stage_3__144_,data_stage_3__143_,
  data_stage_3__142_,data_stage_3__141_,data_stage_3__140_,data_stage_3__139_,data_stage_3__138_,
  data_stage_3__137_,data_stage_3__136_,data_stage_3__135_,data_stage_3__134_,
  data_stage_3__133_,data_stage_3__132_,data_stage_3__131_,data_stage_3__130_,
  data_stage_3__129_,data_stage_3__128_,data_stage_3__127_,data_stage_3__126_,
  data_stage_3__125_,data_stage_3__124_,data_stage_3__123_,data_stage_3__122_,
  data_stage_3__121_,data_stage_3__120_,data_stage_3__119_,data_stage_3__118_,data_stage_3__117_,
  data_stage_3__116_,data_stage_3__115_,data_stage_3__114_,data_stage_3__113_,
  data_stage_3__112_,data_stage_3__111_,data_stage_3__110_,data_stage_3__109_,
  data_stage_3__108_,data_stage_3__107_,data_stage_3__106_,data_stage_3__105_,
  data_stage_3__104_,data_stage_3__103_,data_stage_3__102_,data_stage_3__101_,data_stage_3__100_,
  data_stage_3__99_,data_stage_3__98_,data_stage_3__97_,data_stage_3__96_,
  data_stage_3__95_,data_stage_3__94_,data_stage_3__93_,data_stage_3__92_,
  data_stage_3__91_,data_stage_3__90_,data_stage_3__89_,data_stage_3__88_,data_stage_3__87_,
  data_stage_3__86_,data_stage_3__85_,data_stage_3__84_,data_stage_3__83_,
  data_stage_3__82_,data_stage_3__81_,data_stage_3__80_,data_stage_3__79_,data_stage_3__78_,
  data_stage_3__77_,data_stage_3__76_,data_stage_3__75_,data_stage_3__74_,
  data_stage_3__73_,data_stage_3__72_,data_stage_3__71_,data_stage_3__70_,data_stage_3__69_,
  data_stage_3__68_,data_stage_3__67_,data_stage_3__66_,data_stage_3__65_,
  data_stage_3__64_,data_stage_3__63_,data_stage_3__62_,data_stage_3__61_,data_stage_3__60_,
  data_stage_3__59_,data_stage_3__58_,data_stage_3__57_,data_stage_3__56_,
  data_stage_3__55_,data_stage_3__54_,data_stage_3__53_,data_stage_3__52_,
  data_stage_3__51_,data_stage_3__50_,data_stage_3__49_,data_stage_3__48_,data_stage_3__47_,
  data_stage_3__46_,data_stage_3__45_,data_stage_3__44_,data_stage_3__43_,
  data_stage_3__42_,data_stage_3__41_,data_stage_3__40_,data_stage_3__39_,data_stage_3__38_,
  data_stage_3__37_,data_stage_3__36_,data_stage_3__35_,data_stage_3__34_,
  data_stage_3__33_,data_stage_3__32_,data_stage_3__31_,data_stage_3__30_,data_stage_3__29_,
  data_stage_3__28_,data_stage_3__27_,data_stage_3__26_,data_stage_3__25_,
  data_stage_3__24_,data_stage_3__23_,data_stage_3__22_,data_stage_3__21_,data_stage_3__20_,
  data_stage_3__19_,data_stage_3__18_,data_stage_3__17_,data_stage_3__16_,
  data_stage_3__15_,data_stage_3__14_,data_stage_3__13_,data_stage_3__12_,
  data_stage_3__11_,data_stage_3__10_,data_stage_3__9_,data_stage_3__8_,data_stage_3__7_,
  data_stage_3__6_,data_stage_3__5_,data_stage_3__4_,data_stage_3__3_,data_stage_3__2_,
  data_stage_3__1_,data_stage_3__0_,data_stage_4__8191_,data_stage_4__8190_,
  data_stage_4__8189_,data_stage_4__8188_,data_stage_4__8187_,data_stage_4__8186_,
  data_stage_4__8185_,data_stage_4__8184_,data_stage_4__8183_,data_stage_4__8182_,
  data_stage_4__8181_,data_stage_4__8180_,data_stage_4__8179_,data_stage_4__8178_,
  data_stage_4__8177_,data_stage_4__8176_,data_stage_4__8175_,data_stage_4__8174_,
  data_stage_4__8173_,data_stage_4__8172_,data_stage_4__8171_,data_stage_4__8170_,
  data_stage_4__8169_,data_stage_4__8168_,data_stage_4__8167_,data_stage_4__8166_,
  data_stage_4__8165_,data_stage_4__8164_,data_stage_4__8163_,data_stage_4__8162_,
  data_stage_4__8161_,data_stage_4__8160_,data_stage_4__8159_,data_stage_4__8158_,
  data_stage_4__8157_,data_stage_4__8156_,data_stage_4__8155_,data_stage_4__8154_,
  data_stage_4__8153_,data_stage_4__8152_,data_stage_4__8151_,data_stage_4__8150_,
  data_stage_4__8149_,data_stage_4__8148_,data_stage_4__8147_,data_stage_4__8146_,
  data_stage_4__8145_,data_stage_4__8144_,data_stage_4__8143_,data_stage_4__8142_,
  data_stage_4__8141_,data_stage_4__8140_,data_stage_4__8139_,data_stage_4__8138_,
  data_stage_4__8137_,data_stage_4__8136_,data_stage_4__8135_,data_stage_4__8134_,
  data_stage_4__8133_,data_stage_4__8132_,data_stage_4__8131_,data_stage_4__8130_,
  data_stage_4__8129_,data_stage_4__8128_,data_stage_4__8127_,data_stage_4__8126_,
  data_stage_4__8125_,data_stage_4__8124_,data_stage_4__8123_,data_stage_4__8122_,
  data_stage_4__8121_,data_stage_4__8120_,data_stage_4__8119_,data_stage_4__8118_,
  data_stage_4__8117_,data_stage_4__8116_,data_stage_4__8115_,data_stage_4__8114_,
  data_stage_4__8113_,data_stage_4__8112_,data_stage_4__8111_,data_stage_4__8110_,
  data_stage_4__8109_,data_stage_4__8108_,data_stage_4__8107_,data_stage_4__8106_,
  data_stage_4__8105_,data_stage_4__8104_,data_stage_4__8103_,data_stage_4__8102_,
  data_stage_4__8101_,data_stage_4__8100_,data_stage_4__8099_,data_stage_4__8098_,
  data_stage_4__8097_,data_stage_4__8096_,data_stage_4__8095_,data_stage_4__8094_,
  data_stage_4__8093_,data_stage_4__8092_,data_stage_4__8091_,data_stage_4__8090_,
  data_stage_4__8089_,data_stage_4__8088_,data_stage_4__8087_,data_stage_4__8086_,
  data_stage_4__8085_,data_stage_4__8084_,data_stage_4__8083_,data_stage_4__8082_,
  data_stage_4__8081_,data_stage_4__8080_,data_stage_4__8079_,data_stage_4__8078_,
  data_stage_4__8077_,data_stage_4__8076_,data_stage_4__8075_,data_stage_4__8074_,
  data_stage_4__8073_,data_stage_4__8072_,data_stage_4__8071_,data_stage_4__8070_,
  data_stage_4__8069_,data_stage_4__8068_,data_stage_4__8067_,data_stage_4__8066_,
  data_stage_4__8065_,data_stage_4__8064_,data_stage_4__8063_,data_stage_4__8062_,
  data_stage_4__8061_,data_stage_4__8060_,data_stage_4__8059_,data_stage_4__8058_,
  data_stage_4__8057_,data_stage_4__8056_,data_stage_4__8055_,data_stage_4__8054_,
  data_stage_4__8053_,data_stage_4__8052_,data_stage_4__8051_,data_stage_4__8050_,
  data_stage_4__8049_,data_stage_4__8048_,data_stage_4__8047_,data_stage_4__8046_,
  data_stage_4__8045_,data_stage_4__8044_,data_stage_4__8043_,data_stage_4__8042_,
  data_stage_4__8041_,data_stage_4__8040_,data_stage_4__8039_,data_stage_4__8038_,
  data_stage_4__8037_,data_stage_4__8036_,data_stage_4__8035_,data_stage_4__8034_,
  data_stage_4__8033_,data_stage_4__8032_,data_stage_4__8031_,data_stage_4__8030_,
  data_stage_4__8029_,data_stage_4__8028_,data_stage_4__8027_,data_stage_4__8026_,
  data_stage_4__8025_,data_stage_4__8024_,data_stage_4__8023_,data_stage_4__8022_,
  data_stage_4__8021_,data_stage_4__8020_,data_stage_4__8019_,data_stage_4__8018_,
  data_stage_4__8017_,data_stage_4__8016_,data_stage_4__8015_,data_stage_4__8014_,
  data_stage_4__8013_,data_stage_4__8012_,data_stage_4__8011_,data_stage_4__8010_,
  data_stage_4__8009_,data_stage_4__8008_,data_stage_4__8007_,data_stage_4__8006_,
  data_stage_4__8005_,data_stage_4__8004_,data_stage_4__8003_,data_stage_4__8002_,
  data_stage_4__8001_,data_stage_4__8000_,data_stage_4__7999_,data_stage_4__7998_,
  data_stage_4__7997_,data_stage_4__7996_,data_stage_4__7995_,data_stage_4__7994_,
  data_stage_4__7993_,data_stage_4__7992_,data_stage_4__7991_,data_stage_4__7990_,
  data_stage_4__7989_,data_stage_4__7988_,data_stage_4__7987_,data_stage_4__7986_,
  data_stage_4__7985_,data_stage_4__7984_,data_stage_4__7983_,data_stage_4__7982_,
  data_stage_4__7981_,data_stage_4__7980_,data_stage_4__7979_,data_stage_4__7978_,
  data_stage_4__7977_,data_stage_4__7976_,data_stage_4__7975_,data_stage_4__7974_,
  data_stage_4__7973_,data_stage_4__7972_,data_stage_4__7971_,data_stage_4__7970_,
  data_stage_4__7969_,data_stage_4__7968_,data_stage_4__7967_,data_stage_4__7966_,
  data_stage_4__7965_,data_stage_4__7964_,data_stage_4__7963_,data_stage_4__7962_,
  data_stage_4__7961_,data_stage_4__7960_,data_stage_4__7959_,data_stage_4__7958_,
  data_stage_4__7957_,data_stage_4__7956_,data_stage_4__7955_,data_stage_4__7954_,
  data_stage_4__7953_,data_stage_4__7952_,data_stage_4__7951_,data_stage_4__7950_,
  data_stage_4__7949_,data_stage_4__7948_,data_stage_4__7947_,data_stage_4__7946_,
  data_stage_4__7945_,data_stage_4__7944_,data_stage_4__7943_,data_stage_4__7942_,
  data_stage_4__7941_,data_stage_4__7940_,data_stage_4__7939_,data_stage_4__7938_,
  data_stage_4__7937_,data_stage_4__7936_,data_stage_4__7935_,data_stage_4__7934_,
  data_stage_4__7933_,data_stage_4__7932_,data_stage_4__7931_,data_stage_4__7930_,
  data_stage_4__7929_,data_stage_4__7928_,data_stage_4__7927_,data_stage_4__7926_,
  data_stage_4__7925_,data_stage_4__7924_,data_stage_4__7923_,data_stage_4__7922_,
  data_stage_4__7921_,data_stage_4__7920_,data_stage_4__7919_,data_stage_4__7918_,
  data_stage_4__7917_,data_stage_4__7916_,data_stage_4__7915_,data_stage_4__7914_,
  data_stage_4__7913_,data_stage_4__7912_,data_stage_4__7911_,data_stage_4__7910_,
  data_stage_4__7909_,data_stage_4__7908_,data_stage_4__7907_,data_stage_4__7906_,
  data_stage_4__7905_,data_stage_4__7904_,data_stage_4__7903_,data_stage_4__7902_,
  data_stage_4__7901_,data_stage_4__7900_,data_stage_4__7899_,data_stage_4__7898_,
  data_stage_4__7897_,data_stage_4__7896_,data_stage_4__7895_,data_stage_4__7894_,
  data_stage_4__7893_,data_stage_4__7892_,data_stage_4__7891_,data_stage_4__7890_,
  data_stage_4__7889_,data_stage_4__7888_,data_stage_4__7887_,data_stage_4__7886_,
  data_stage_4__7885_,data_stage_4__7884_,data_stage_4__7883_,data_stage_4__7882_,
  data_stage_4__7881_,data_stage_4__7880_,data_stage_4__7879_,data_stage_4__7878_,
  data_stage_4__7877_,data_stage_4__7876_,data_stage_4__7875_,data_stage_4__7874_,
  data_stage_4__7873_,data_stage_4__7872_,data_stage_4__7871_,data_stage_4__7870_,
  data_stage_4__7869_,data_stage_4__7868_,data_stage_4__7867_,data_stage_4__7866_,
  data_stage_4__7865_,data_stage_4__7864_,data_stage_4__7863_,data_stage_4__7862_,
  data_stage_4__7861_,data_stage_4__7860_,data_stage_4__7859_,data_stage_4__7858_,
  data_stage_4__7857_,data_stage_4__7856_,data_stage_4__7855_,data_stage_4__7854_,
  data_stage_4__7853_,data_stage_4__7852_,data_stage_4__7851_,data_stage_4__7850_,
  data_stage_4__7849_,data_stage_4__7848_,data_stage_4__7847_,data_stage_4__7846_,
  data_stage_4__7845_,data_stage_4__7844_,data_stage_4__7843_,data_stage_4__7842_,
  data_stage_4__7841_,data_stage_4__7840_,data_stage_4__7839_,data_stage_4__7838_,
  data_stage_4__7837_,data_stage_4__7836_,data_stage_4__7835_,data_stage_4__7834_,
  data_stage_4__7833_,data_stage_4__7832_,data_stage_4__7831_,data_stage_4__7830_,
  data_stage_4__7829_,data_stage_4__7828_,data_stage_4__7827_,data_stage_4__7826_,
  data_stage_4__7825_,data_stage_4__7824_,data_stage_4__7823_,data_stage_4__7822_,
  data_stage_4__7821_,data_stage_4__7820_,data_stage_4__7819_,data_stage_4__7818_,
  data_stage_4__7817_,data_stage_4__7816_,data_stage_4__7815_,data_stage_4__7814_,
  data_stage_4__7813_,data_stage_4__7812_,data_stage_4__7811_,data_stage_4__7810_,
  data_stage_4__7809_,data_stage_4__7808_,data_stage_4__7807_,data_stage_4__7806_,
  data_stage_4__7805_,data_stage_4__7804_,data_stage_4__7803_,data_stage_4__7802_,
  data_stage_4__7801_,data_stage_4__7800_,data_stage_4__7799_,data_stage_4__7798_,
  data_stage_4__7797_,data_stage_4__7796_,data_stage_4__7795_,data_stage_4__7794_,
  data_stage_4__7793_,data_stage_4__7792_,data_stage_4__7791_,data_stage_4__7790_,
  data_stage_4__7789_,data_stage_4__7788_,data_stage_4__7787_,data_stage_4__7786_,
  data_stage_4__7785_,data_stage_4__7784_,data_stage_4__7783_,data_stage_4__7782_,
  data_stage_4__7781_,data_stage_4__7780_,data_stage_4__7779_,data_stage_4__7778_,
  data_stage_4__7777_,data_stage_4__7776_,data_stage_4__7775_,data_stage_4__7774_,
  data_stage_4__7773_,data_stage_4__7772_,data_stage_4__7771_,data_stage_4__7770_,
  data_stage_4__7769_,data_stage_4__7768_,data_stage_4__7767_,data_stage_4__7766_,
  data_stage_4__7765_,data_stage_4__7764_,data_stage_4__7763_,data_stage_4__7762_,
  data_stage_4__7761_,data_stage_4__7760_,data_stage_4__7759_,data_stage_4__7758_,
  data_stage_4__7757_,data_stage_4__7756_,data_stage_4__7755_,data_stage_4__7754_,
  data_stage_4__7753_,data_stage_4__7752_,data_stage_4__7751_,data_stage_4__7750_,
  data_stage_4__7749_,data_stage_4__7748_,data_stage_4__7747_,data_stage_4__7746_,
  data_stage_4__7745_,data_stage_4__7744_,data_stage_4__7743_,data_stage_4__7742_,
  data_stage_4__7741_,data_stage_4__7740_,data_stage_4__7739_,data_stage_4__7738_,
  data_stage_4__7737_,data_stage_4__7736_,data_stage_4__7735_,data_stage_4__7734_,
  data_stage_4__7733_,data_stage_4__7732_,data_stage_4__7731_,data_stage_4__7730_,
  data_stage_4__7729_,data_stage_4__7728_,data_stage_4__7727_,data_stage_4__7726_,
  data_stage_4__7725_,data_stage_4__7724_,data_stage_4__7723_,data_stage_4__7722_,
  data_stage_4__7721_,data_stage_4__7720_,data_stage_4__7719_,data_stage_4__7718_,
  data_stage_4__7717_,data_stage_4__7716_,data_stage_4__7715_,data_stage_4__7714_,
  data_stage_4__7713_,data_stage_4__7712_,data_stage_4__7711_,data_stage_4__7710_,
  data_stage_4__7709_,data_stage_4__7708_,data_stage_4__7707_,data_stage_4__7706_,
  data_stage_4__7705_,data_stage_4__7704_,data_stage_4__7703_,data_stage_4__7702_,
  data_stage_4__7701_,data_stage_4__7700_,data_stage_4__7699_,data_stage_4__7698_,
  data_stage_4__7697_,data_stage_4__7696_,data_stage_4__7695_,data_stage_4__7694_,
  data_stage_4__7693_,data_stage_4__7692_,data_stage_4__7691_,data_stage_4__7690_,
  data_stage_4__7689_,data_stage_4__7688_,data_stage_4__7687_,data_stage_4__7686_,
  data_stage_4__7685_,data_stage_4__7684_,data_stage_4__7683_,data_stage_4__7682_,
  data_stage_4__7681_,data_stage_4__7680_,data_stage_4__7679_,data_stage_4__7678_,
  data_stage_4__7677_,data_stage_4__7676_,data_stage_4__7675_,data_stage_4__7674_,
  data_stage_4__7673_,data_stage_4__7672_,data_stage_4__7671_,data_stage_4__7670_,
  data_stage_4__7669_,data_stage_4__7668_,data_stage_4__7667_,data_stage_4__7666_,
  data_stage_4__7665_,data_stage_4__7664_,data_stage_4__7663_,data_stage_4__7662_,
  data_stage_4__7661_,data_stage_4__7660_,data_stage_4__7659_,data_stage_4__7658_,
  data_stage_4__7657_,data_stage_4__7656_,data_stage_4__7655_,data_stage_4__7654_,
  data_stage_4__7653_,data_stage_4__7652_,data_stage_4__7651_,data_stage_4__7650_,
  data_stage_4__7649_,data_stage_4__7648_,data_stage_4__7647_,data_stage_4__7646_,
  data_stage_4__7645_,data_stage_4__7644_,data_stage_4__7643_,data_stage_4__7642_,
  data_stage_4__7641_,data_stage_4__7640_,data_stage_4__7639_,data_stage_4__7638_,
  data_stage_4__7637_,data_stage_4__7636_,data_stage_4__7635_,data_stage_4__7634_,
  data_stage_4__7633_,data_stage_4__7632_,data_stage_4__7631_,data_stage_4__7630_,
  data_stage_4__7629_,data_stage_4__7628_,data_stage_4__7627_,data_stage_4__7626_,
  data_stage_4__7625_,data_stage_4__7624_,data_stage_4__7623_,data_stage_4__7622_,
  data_stage_4__7621_,data_stage_4__7620_,data_stage_4__7619_,data_stage_4__7618_,
  data_stage_4__7617_,data_stage_4__7616_,data_stage_4__7615_,data_stage_4__7614_,
  data_stage_4__7613_,data_stage_4__7612_,data_stage_4__7611_,data_stage_4__7610_,
  data_stage_4__7609_,data_stage_4__7608_,data_stage_4__7607_,data_stage_4__7606_,
  data_stage_4__7605_,data_stage_4__7604_,data_stage_4__7603_,data_stage_4__7602_,
  data_stage_4__7601_,data_stage_4__7600_,data_stage_4__7599_,data_stage_4__7598_,
  data_stage_4__7597_,data_stage_4__7596_,data_stage_4__7595_,data_stage_4__7594_,
  data_stage_4__7593_,data_stage_4__7592_,data_stage_4__7591_,data_stage_4__7590_,
  data_stage_4__7589_,data_stage_4__7588_,data_stage_4__7587_,data_stage_4__7586_,
  data_stage_4__7585_,data_stage_4__7584_,data_stage_4__7583_,data_stage_4__7582_,
  data_stage_4__7581_,data_stage_4__7580_,data_stage_4__7579_,data_stage_4__7578_,
  data_stage_4__7577_,data_stage_4__7576_,data_stage_4__7575_,data_stage_4__7574_,
  data_stage_4__7573_,data_stage_4__7572_,data_stage_4__7571_,data_stage_4__7570_,
  data_stage_4__7569_,data_stage_4__7568_,data_stage_4__7567_,data_stage_4__7566_,
  data_stage_4__7565_,data_stage_4__7564_,data_stage_4__7563_,data_stage_4__7562_,
  data_stage_4__7561_,data_stage_4__7560_,data_stage_4__7559_,data_stage_4__7558_,
  data_stage_4__7557_,data_stage_4__7556_,data_stage_4__7555_,data_stage_4__7554_,
  data_stage_4__7553_,data_stage_4__7552_,data_stage_4__7551_,data_stage_4__7550_,
  data_stage_4__7549_,data_stage_4__7548_,data_stage_4__7547_,data_stage_4__7546_,
  data_stage_4__7545_,data_stage_4__7544_,data_stage_4__7543_,data_stage_4__7542_,
  data_stage_4__7541_,data_stage_4__7540_,data_stage_4__7539_,data_stage_4__7538_,
  data_stage_4__7537_,data_stage_4__7536_,data_stage_4__7535_,data_stage_4__7534_,
  data_stage_4__7533_,data_stage_4__7532_,data_stage_4__7531_,data_stage_4__7530_,
  data_stage_4__7529_,data_stage_4__7528_,data_stage_4__7527_,data_stage_4__7526_,
  data_stage_4__7525_,data_stage_4__7524_,data_stage_4__7523_,data_stage_4__7522_,
  data_stage_4__7521_,data_stage_4__7520_,data_stage_4__7519_,data_stage_4__7518_,
  data_stage_4__7517_,data_stage_4__7516_,data_stage_4__7515_,data_stage_4__7514_,
  data_stage_4__7513_,data_stage_4__7512_,data_stage_4__7511_,data_stage_4__7510_,
  data_stage_4__7509_,data_stage_4__7508_,data_stage_4__7507_,data_stage_4__7506_,
  data_stage_4__7505_,data_stage_4__7504_,data_stage_4__7503_,data_stage_4__7502_,
  data_stage_4__7501_,data_stage_4__7500_,data_stage_4__7499_,data_stage_4__7498_,
  data_stage_4__7497_,data_stage_4__7496_,data_stage_4__7495_,data_stage_4__7494_,
  data_stage_4__7493_,data_stage_4__7492_,data_stage_4__7491_,data_stage_4__7490_,
  data_stage_4__7489_,data_stage_4__7488_,data_stage_4__7487_,data_stage_4__7486_,
  data_stage_4__7485_,data_stage_4__7484_,data_stage_4__7483_,data_stage_4__7482_,
  data_stage_4__7481_,data_stage_4__7480_,data_stage_4__7479_,data_stage_4__7478_,
  data_stage_4__7477_,data_stage_4__7476_,data_stage_4__7475_,data_stage_4__7474_,
  data_stage_4__7473_,data_stage_4__7472_,data_stage_4__7471_,data_stage_4__7470_,
  data_stage_4__7469_,data_stage_4__7468_,data_stage_4__7467_,data_stage_4__7466_,
  data_stage_4__7465_,data_stage_4__7464_,data_stage_4__7463_,data_stage_4__7462_,
  data_stage_4__7461_,data_stage_4__7460_,data_stage_4__7459_,data_stage_4__7458_,
  data_stage_4__7457_,data_stage_4__7456_,data_stage_4__7455_,data_stage_4__7454_,
  data_stage_4__7453_,data_stage_4__7452_,data_stage_4__7451_,data_stage_4__7450_,
  data_stage_4__7449_,data_stage_4__7448_,data_stage_4__7447_,data_stage_4__7446_,
  data_stage_4__7445_,data_stage_4__7444_,data_stage_4__7443_,data_stage_4__7442_,
  data_stage_4__7441_,data_stage_4__7440_,data_stage_4__7439_,data_stage_4__7438_,
  data_stage_4__7437_,data_stage_4__7436_,data_stage_4__7435_,data_stage_4__7434_,
  data_stage_4__7433_,data_stage_4__7432_,data_stage_4__7431_,data_stage_4__7430_,
  data_stage_4__7429_,data_stage_4__7428_,data_stage_4__7427_,data_stage_4__7426_,
  data_stage_4__7425_,data_stage_4__7424_,data_stage_4__7423_,data_stage_4__7422_,
  data_stage_4__7421_,data_stage_4__7420_,data_stage_4__7419_,data_stage_4__7418_,
  data_stage_4__7417_,data_stage_4__7416_,data_stage_4__7415_,data_stage_4__7414_,
  data_stage_4__7413_,data_stage_4__7412_,data_stage_4__7411_,data_stage_4__7410_,
  data_stage_4__7409_,data_stage_4__7408_,data_stage_4__7407_,data_stage_4__7406_,
  data_stage_4__7405_,data_stage_4__7404_,data_stage_4__7403_,data_stage_4__7402_,
  data_stage_4__7401_,data_stage_4__7400_,data_stage_4__7399_,data_stage_4__7398_,
  data_stage_4__7397_,data_stage_4__7396_,data_stage_4__7395_,data_stage_4__7394_,
  data_stage_4__7393_,data_stage_4__7392_,data_stage_4__7391_,data_stage_4__7390_,
  data_stage_4__7389_,data_stage_4__7388_,data_stage_4__7387_,data_stage_4__7386_,
  data_stage_4__7385_,data_stage_4__7384_,data_stage_4__7383_,data_stage_4__7382_,
  data_stage_4__7381_,data_stage_4__7380_,data_stage_4__7379_,data_stage_4__7378_,
  data_stage_4__7377_,data_stage_4__7376_,data_stage_4__7375_,data_stage_4__7374_,
  data_stage_4__7373_,data_stage_4__7372_,data_stage_4__7371_,data_stage_4__7370_,
  data_stage_4__7369_,data_stage_4__7368_,data_stage_4__7367_,data_stage_4__7366_,
  data_stage_4__7365_,data_stage_4__7364_,data_stage_4__7363_,data_stage_4__7362_,
  data_stage_4__7361_,data_stage_4__7360_,data_stage_4__7359_,data_stage_4__7358_,
  data_stage_4__7357_,data_stage_4__7356_,data_stage_4__7355_,data_stage_4__7354_,
  data_stage_4__7353_,data_stage_4__7352_,data_stage_4__7351_,data_stage_4__7350_,
  data_stage_4__7349_,data_stage_4__7348_,data_stage_4__7347_,data_stage_4__7346_,
  data_stage_4__7345_,data_stage_4__7344_,data_stage_4__7343_,data_stage_4__7342_,
  data_stage_4__7341_,data_stage_4__7340_,data_stage_4__7339_,data_stage_4__7338_,
  data_stage_4__7337_,data_stage_4__7336_,data_stage_4__7335_,data_stage_4__7334_,
  data_stage_4__7333_,data_stage_4__7332_,data_stage_4__7331_,data_stage_4__7330_,
  data_stage_4__7329_,data_stage_4__7328_,data_stage_4__7327_,data_stage_4__7326_,
  data_stage_4__7325_,data_stage_4__7324_,data_stage_4__7323_,data_stage_4__7322_,
  data_stage_4__7321_,data_stage_4__7320_,data_stage_4__7319_,data_stage_4__7318_,
  data_stage_4__7317_,data_stage_4__7316_,data_stage_4__7315_,data_stage_4__7314_,
  data_stage_4__7313_,data_stage_4__7312_,data_stage_4__7311_,data_stage_4__7310_,
  data_stage_4__7309_,data_stage_4__7308_,data_stage_4__7307_,data_stage_4__7306_,
  data_stage_4__7305_,data_stage_4__7304_,data_stage_4__7303_,data_stage_4__7302_,
  data_stage_4__7301_,data_stage_4__7300_,data_stage_4__7299_,data_stage_4__7298_,
  data_stage_4__7297_,data_stage_4__7296_,data_stage_4__7295_,data_stage_4__7294_,
  data_stage_4__7293_,data_stage_4__7292_,data_stage_4__7291_,data_stage_4__7290_,
  data_stage_4__7289_,data_stage_4__7288_,data_stage_4__7287_,data_stage_4__7286_,
  data_stage_4__7285_,data_stage_4__7284_,data_stage_4__7283_,data_stage_4__7282_,
  data_stage_4__7281_,data_stage_4__7280_,data_stage_4__7279_,data_stage_4__7278_,
  data_stage_4__7277_,data_stage_4__7276_,data_stage_4__7275_,data_stage_4__7274_,
  data_stage_4__7273_,data_stage_4__7272_,data_stage_4__7271_,data_stage_4__7270_,
  data_stage_4__7269_,data_stage_4__7268_,data_stage_4__7267_,data_stage_4__7266_,
  data_stage_4__7265_,data_stage_4__7264_,data_stage_4__7263_,data_stage_4__7262_,
  data_stage_4__7261_,data_stage_4__7260_,data_stage_4__7259_,data_stage_4__7258_,
  data_stage_4__7257_,data_stage_4__7256_,data_stage_4__7255_,data_stage_4__7254_,
  data_stage_4__7253_,data_stage_4__7252_,data_stage_4__7251_,data_stage_4__7250_,
  data_stage_4__7249_,data_stage_4__7248_,data_stage_4__7247_,data_stage_4__7246_,
  data_stage_4__7245_,data_stage_4__7244_,data_stage_4__7243_,data_stage_4__7242_,
  data_stage_4__7241_,data_stage_4__7240_,data_stage_4__7239_,data_stage_4__7238_,
  data_stage_4__7237_,data_stage_4__7236_,data_stage_4__7235_,data_stage_4__7234_,
  data_stage_4__7233_,data_stage_4__7232_,data_stage_4__7231_,data_stage_4__7230_,
  data_stage_4__7229_,data_stage_4__7228_,data_stage_4__7227_,data_stage_4__7226_,
  data_stage_4__7225_,data_stage_4__7224_,data_stage_4__7223_,data_stage_4__7222_,
  data_stage_4__7221_,data_stage_4__7220_,data_stage_4__7219_,data_stage_4__7218_,
  data_stage_4__7217_,data_stage_4__7216_,data_stage_4__7215_,data_stage_4__7214_,
  data_stage_4__7213_,data_stage_4__7212_,data_stage_4__7211_,data_stage_4__7210_,
  data_stage_4__7209_,data_stage_4__7208_,data_stage_4__7207_,data_stage_4__7206_,
  data_stage_4__7205_,data_stage_4__7204_,data_stage_4__7203_,data_stage_4__7202_,
  data_stage_4__7201_,data_stage_4__7200_,data_stage_4__7199_,data_stage_4__7198_,
  data_stage_4__7197_,data_stage_4__7196_,data_stage_4__7195_,data_stage_4__7194_,
  data_stage_4__7193_,data_stage_4__7192_,data_stage_4__7191_,data_stage_4__7190_,
  data_stage_4__7189_,data_stage_4__7188_,data_stage_4__7187_,data_stage_4__7186_,
  data_stage_4__7185_,data_stage_4__7184_,data_stage_4__7183_,data_stage_4__7182_,
  data_stage_4__7181_,data_stage_4__7180_,data_stage_4__7179_,data_stage_4__7178_,
  data_stage_4__7177_,data_stage_4__7176_,data_stage_4__7175_,data_stage_4__7174_,
  data_stage_4__7173_,data_stage_4__7172_,data_stage_4__7171_,data_stage_4__7170_,
  data_stage_4__7169_,data_stage_4__7168_,data_stage_4__7167_,data_stage_4__7166_,
  data_stage_4__7165_,data_stage_4__7164_,data_stage_4__7163_,data_stage_4__7162_,
  data_stage_4__7161_,data_stage_4__7160_,data_stage_4__7159_,data_stage_4__7158_,
  data_stage_4__7157_,data_stage_4__7156_,data_stage_4__7155_,data_stage_4__7154_,
  data_stage_4__7153_,data_stage_4__7152_,data_stage_4__7151_,data_stage_4__7150_,
  data_stage_4__7149_,data_stage_4__7148_,data_stage_4__7147_,data_stage_4__7146_,
  data_stage_4__7145_,data_stage_4__7144_,data_stage_4__7143_,data_stage_4__7142_,
  data_stage_4__7141_,data_stage_4__7140_,data_stage_4__7139_,data_stage_4__7138_,
  data_stage_4__7137_,data_stage_4__7136_,data_stage_4__7135_,data_stage_4__7134_,
  data_stage_4__7133_,data_stage_4__7132_,data_stage_4__7131_,data_stage_4__7130_,
  data_stage_4__7129_,data_stage_4__7128_,data_stage_4__7127_,data_stage_4__7126_,
  data_stage_4__7125_,data_stage_4__7124_,data_stage_4__7123_,data_stage_4__7122_,
  data_stage_4__7121_,data_stage_4__7120_,data_stage_4__7119_,data_stage_4__7118_,
  data_stage_4__7117_,data_stage_4__7116_,data_stage_4__7115_,data_stage_4__7114_,
  data_stage_4__7113_,data_stage_4__7112_,data_stage_4__7111_,data_stage_4__7110_,
  data_stage_4__7109_,data_stage_4__7108_,data_stage_4__7107_,data_stage_4__7106_,
  data_stage_4__7105_,data_stage_4__7104_,data_stage_4__7103_,data_stage_4__7102_,
  data_stage_4__7101_,data_stage_4__7100_,data_stage_4__7099_,data_stage_4__7098_,
  data_stage_4__7097_,data_stage_4__7096_,data_stage_4__7095_,data_stage_4__7094_,
  data_stage_4__7093_,data_stage_4__7092_,data_stage_4__7091_,data_stage_4__7090_,
  data_stage_4__7089_,data_stage_4__7088_,data_stage_4__7087_,data_stage_4__7086_,
  data_stage_4__7085_,data_stage_4__7084_,data_stage_4__7083_,data_stage_4__7082_,
  data_stage_4__7081_,data_stage_4__7080_,data_stage_4__7079_,data_stage_4__7078_,
  data_stage_4__7077_,data_stage_4__7076_,data_stage_4__7075_,data_stage_4__7074_,
  data_stage_4__7073_,data_stage_4__7072_,data_stage_4__7071_,data_stage_4__7070_,
  data_stage_4__7069_,data_stage_4__7068_,data_stage_4__7067_,data_stage_4__7066_,
  data_stage_4__7065_,data_stage_4__7064_,data_stage_4__7063_,data_stage_4__7062_,
  data_stage_4__7061_,data_stage_4__7060_,data_stage_4__7059_,data_stage_4__7058_,
  data_stage_4__7057_,data_stage_4__7056_,data_stage_4__7055_,data_stage_4__7054_,
  data_stage_4__7053_,data_stage_4__7052_,data_stage_4__7051_,data_stage_4__7050_,
  data_stage_4__7049_,data_stage_4__7048_,data_stage_4__7047_,data_stage_4__7046_,
  data_stage_4__7045_,data_stage_4__7044_,data_stage_4__7043_,data_stage_4__7042_,
  data_stage_4__7041_,data_stage_4__7040_,data_stage_4__7039_,data_stage_4__7038_,
  data_stage_4__7037_,data_stage_4__7036_,data_stage_4__7035_,data_stage_4__7034_,
  data_stage_4__7033_,data_stage_4__7032_,data_stage_4__7031_,data_stage_4__7030_,
  data_stage_4__7029_,data_stage_4__7028_,data_stage_4__7027_,data_stage_4__7026_,
  data_stage_4__7025_,data_stage_4__7024_,data_stage_4__7023_,data_stage_4__7022_,
  data_stage_4__7021_,data_stage_4__7020_,data_stage_4__7019_,data_stage_4__7018_,
  data_stage_4__7017_,data_stage_4__7016_,data_stage_4__7015_,data_stage_4__7014_,
  data_stage_4__7013_,data_stage_4__7012_,data_stage_4__7011_,data_stage_4__7010_,
  data_stage_4__7009_,data_stage_4__7008_,data_stage_4__7007_,data_stage_4__7006_,
  data_stage_4__7005_,data_stage_4__7004_,data_stage_4__7003_,data_stage_4__7002_,
  data_stage_4__7001_,data_stage_4__7000_,data_stage_4__6999_,data_stage_4__6998_,
  data_stage_4__6997_,data_stage_4__6996_,data_stage_4__6995_,data_stage_4__6994_,
  data_stage_4__6993_,data_stage_4__6992_,data_stage_4__6991_,data_stage_4__6990_,
  data_stage_4__6989_,data_stage_4__6988_,data_stage_4__6987_,data_stage_4__6986_,
  data_stage_4__6985_,data_stage_4__6984_,data_stage_4__6983_,data_stage_4__6982_,
  data_stage_4__6981_,data_stage_4__6980_,data_stage_4__6979_,data_stage_4__6978_,
  data_stage_4__6977_,data_stage_4__6976_,data_stage_4__6975_,data_stage_4__6974_,
  data_stage_4__6973_,data_stage_4__6972_,data_stage_4__6971_,data_stage_4__6970_,
  data_stage_4__6969_,data_stage_4__6968_,data_stage_4__6967_,data_stage_4__6966_,
  data_stage_4__6965_,data_stage_4__6964_,data_stage_4__6963_,data_stage_4__6962_,
  data_stage_4__6961_,data_stage_4__6960_,data_stage_4__6959_,data_stage_4__6958_,
  data_stage_4__6957_,data_stage_4__6956_,data_stage_4__6955_,data_stage_4__6954_,
  data_stage_4__6953_,data_stage_4__6952_,data_stage_4__6951_,data_stage_4__6950_,
  data_stage_4__6949_,data_stage_4__6948_,data_stage_4__6947_,data_stage_4__6946_,
  data_stage_4__6945_,data_stage_4__6944_,data_stage_4__6943_,data_stage_4__6942_,
  data_stage_4__6941_,data_stage_4__6940_,data_stage_4__6939_,data_stage_4__6938_,
  data_stage_4__6937_,data_stage_4__6936_,data_stage_4__6935_,data_stage_4__6934_,
  data_stage_4__6933_,data_stage_4__6932_,data_stage_4__6931_,data_stage_4__6930_,
  data_stage_4__6929_,data_stage_4__6928_,data_stage_4__6927_,data_stage_4__6926_,
  data_stage_4__6925_,data_stage_4__6924_,data_stage_4__6923_,data_stage_4__6922_,
  data_stage_4__6921_,data_stage_4__6920_,data_stage_4__6919_,data_stage_4__6918_,
  data_stage_4__6917_,data_stage_4__6916_,data_stage_4__6915_,data_stage_4__6914_,
  data_stage_4__6913_,data_stage_4__6912_,data_stage_4__6911_,data_stage_4__6910_,
  data_stage_4__6909_,data_stage_4__6908_,data_stage_4__6907_,data_stage_4__6906_,
  data_stage_4__6905_,data_stage_4__6904_,data_stage_4__6903_,data_stage_4__6902_,
  data_stage_4__6901_,data_stage_4__6900_,data_stage_4__6899_,data_stage_4__6898_,
  data_stage_4__6897_,data_stage_4__6896_,data_stage_4__6895_,data_stage_4__6894_,
  data_stage_4__6893_,data_stage_4__6892_,data_stage_4__6891_,data_stage_4__6890_,
  data_stage_4__6889_,data_stage_4__6888_,data_stage_4__6887_,data_stage_4__6886_,
  data_stage_4__6885_,data_stage_4__6884_,data_stage_4__6883_,data_stage_4__6882_,
  data_stage_4__6881_,data_stage_4__6880_,data_stage_4__6879_,data_stage_4__6878_,
  data_stage_4__6877_,data_stage_4__6876_,data_stage_4__6875_,data_stage_4__6874_,
  data_stage_4__6873_,data_stage_4__6872_,data_stage_4__6871_,data_stage_4__6870_,
  data_stage_4__6869_,data_stage_4__6868_,data_stage_4__6867_,data_stage_4__6866_,
  data_stage_4__6865_,data_stage_4__6864_,data_stage_4__6863_,data_stage_4__6862_,
  data_stage_4__6861_,data_stage_4__6860_,data_stage_4__6859_,data_stage_4__6858_,
  data_stage_4__6857_,data_stage_4__6856_,data_stage_4__6855_,data_stage_4__6854_,
  data_stage_4__6853_,data_stage_4__6852_,data_stage_4__6851_,data_stage_4__6850_,
  data_stage_4__6849_,data_stage_4__6848_,data_stage_4__6847_,data_stage_4__6846_,
  data_stage_4__6845_,data_stage_4__6844_,data_stage_4__6843_,data_stage_4__6842_,
  data_stage_4__6841_,data_stage_4__6840_,data_stage_4__6839_,data_stage_4__6838_,
  data_stage_4__6837_,data_stage_4__6836_,data_stage_4__6835_,data_stage_4__6834_,
  data_stage_4__6833_,data_stage_4__6832_,data_stage_4__6831_,data_stage_4__6830_,
  data_stage_4__6829_,data_stage_4__6828_,data_stage_4__6827_,data_stage_4__6826_,
  data_stage_4__6825_,data_stage_4__6824_,data_stage_4__6823_,data_stage_4__6822_,
  data_stage_4__6821_,data_stage_4__6820_,data_stage_4__6819_,data_stage_4__6818_,
  data_stage_4__6817_,data_stage_4__6816_,data_stage_4__6815_,data_stage_4__6814_,
  data_stage_4__6813_,data_stage_4__6812_,data_stage_4__6811_,data_stage_4__6810_,
  data_stage_4__6809_,data_stage_4__6808_,data_stage_4__6807_,data_stage_4__6806_,
  data_stage_4__6805_,data_stage_4__6804_,data_stage_4__6803_,data_stage_4__6802_,
  data_stage_4__6801_,data_stage_4__6800_,data_stage_4__6799_,data_stage_4__6798_,
  data_stage_4__6797_,data_stage_4__6796_,data_stage_4__6795_,data_stage_4__6794_,
  data_stage_4__6793_,data_stage_4__6792_,data_stage_4__6791_,data_stage_4__6790_,
  data_stage_4__6789_,data_stage_4__6788_,data_stage_4__6787_,data_stage_4__6786_,
  data_stage_4__6785_,data_stage_4__6784_,data_stage_4__6783_,data_stage_4__6782_,
  data_stage_4__6781_,data_stage_4__6780_,data_stage_4__6779_,data_stage_4__6778_,
  data_stage_4__6777_,data_stage_4__6776_,data_stage_4__6775_,data_stage_4__6774_,
  data_stage_4__6773_,data_stage_4__6772_,data_stage_4__6771_,data_stage_4__6770_,
  data_stage_4__6769_,data_stage_4__6768_,data_stage_4__6767_,data_stage_4__6766_,
  data_stage_4__6765_,data_stage_4__6764_,data_stage_4__6763_,data_stage_4__6762_,
  data_stage_4__6761_,data_stage_4__6760_,data_stage_4__6759_,data_stage_4__6758_,
  data_stage_4__6757_,data_stage_4__6756_,data_stage_4__6755_,data_stage_4__6754_,
  data_stage_4__6753_,data_stage_4__6752_,data_stage_4__6751_,data_stage_4__6750_,
  data_stage_4__6749_,data_stage_4__6748_,data_stage_4__6747_,data_stage_4__6746_,
  data_stage_4__6745_,data_stage_4__6744_,data_stage_4__6743_,data_stage_4__6742_,
  data_stage_4__6741_,data_stage_4__6740_,data_stage_4__6739_,data_stage_4__6738_,
  data_stage_4__6737_,data_stage_4__6736_,data_stage_4__6735_,data_stage_4__6734_,
  data_stage_4__6733_,data_stage_4__6732_,data_stage_4__6731_,data_stage_4__6730_,
  data_stage_4__6729_,data_stage_4__6728_,data_stage_4__6727_,data_stage_4__6726_,
  data_stage_4__6725_,data_stage_4__6724_,data_stage_4__6723_,data_stage_4__6722_,
  data_stage_4__6721_,data_stage_4__6720_,data_stage_4__6719_,data_stage_4__6718_,
  data_stage_4__6717_,data_stage_4__6716_,data_stage_4__6715_,data_stage_4__6714_,
  data_stage_4__6713_,data_stage_4__6712_,data_stage_4__6711_,data_stage_4__6710_,
  data_stage_4__6709_,data_stage_4__6708_,data_stage_4__6707_,data_stage_4__6706_,
  data_stage_4__6705_,data_stage_4__6704_,data_stage_4__6703_,data_stage_4__6702_,
  data_stage_4__6701_,data_stage_4__6700_,data_stage_4__6699_,data_stage_4__6698_,
  data_stage_4__6697_,data_stage_4__6696_,data_stage_4__6695_,data_stage_4__6694_,
  data_stage_4__6693_,data_stage_4__6692_,data_stage_4__6691_,data_stage_4__6690_,
  data_stage_4__6689_,data_stage_4__6688_,data_stage_4__6687_,data_stage_4__6686_,
  data_stage_4__6685_,data_stage_4__6684_,data_stage_4__6683_,data_stage_4__6682_,
  data_stage_4__6681_,data_stage_4__6680_,data_stage_4__6679_,data_stage_4__6678_,
  data_stage_4__6677_,data_stage_4__6676_,data_stage_4__6675_,data_stage_4__6674_,
  data_stage_4__6673_,data_stage_4__6672_,data_stage_4__6671_,data_stage_4__6670_,
  data_stage_4__6669_,data_stage_4__6668_,data_stage_4__6667_,data_stage_4__6666_,
  data_stage_4__6665_,data_stage_4__6664_,data_stage_4__6663_,data_stage_4__6662_,
  data_stage_4__6661_,data_stage_4__6660_,data_stage_4__6659_,data_stage_4__6658_,
  data_stage_4__6657_,data_stage_4__6656_,data_stage_4__6655_,data_stage_4__6654_,
  data_stage_4__6653_,data_stage_4__6652_,data_stage_4__6651_,data_stage_4__6650_,
  data_stage_4__6649_,data_stage_4__6648_,data_stage_4__6647_,data_stage_4__6646_,
  data_stage_4__6645_,data_stage_4__6644_,data_stage_4__6643_,data_stage_4__6642_,
  data_stage_4__6641_,data_stage_4__6640_,data_stage_4__6639_,data_stage_4__6638_,
  data_stage_4__6637_,data_stage_4__6636_,data_stage_4__6635_,data_stage_4__6634_,
  data_stage_4__6633_,data_stage_4__6632_,data_stage_4__6631_,data_stage_4__6630_,
  data_stage_4__6629_,data_stage_4__6628_,data_stage_4__6627_,data_stage_4__6626_,
  data_stage_4__6625_,data_stage_4__6624_,data_stage_4__6623_,data_stage_4__6622_,
  data_stage_4__6621_,data_stage_4__6620_,data_stage_4__6619_,data_stage_4__6618_,
  data_stage_4__6617_,data_stage_4__6616_,data_stage_4__6615_,data_stage_4__6614_,
  data_stage_4__6613_,data_stage_4__6612_,data_stage_4__6611_,data_stage_4__6610_,
  data_stage_4__6609_,data_stage_4__6608_,data_stage_4__6607_,data_stage_4__6606_,
  data_stage_4__6605_,data_stage_4__6604_,data_stage_4__6603_,data_stage_4__6602_,
  data_stage_4__6601_,data_stage_4__6600_,data_stage_4__6599_,data_stage_4__6598_,
  data_stage_4__6597_,data_stage_4__6596_,data_stage_4__6595_,data_stage_4__6594_,
  data_stage_4__6593_,data_stage_4__6592_,data_stage_4__6591_,data_stage_4__6590_,
  data_stage_4__6589_,data_stage_4__6588_,data_stage_4__6587_,data_stage_4__6586_,
  data_stage_4__6585_,data_stage_4__6584_,data_stage_4__6583_,data_stage_4__6582_,
  data_stage_4__6581_,data_stage_4__6580_,data_stage_4__6579_,data_stage_4__6578_,
  data_stage_4__6577_,data_stage_4__6576_,data_stage_4__6575_,data_stage_4__6574_,
  data_stage_4__6573_,data_stage_4__6572_,data_stage_4__6571_,data_stage_4__6570_,
  data_stage_4__6569_,data_stage_4__6568_,data_stage_4__6567_,data_stage_4__6566_,
  data_stage_4__6565_,data_stage_4__6564_,data_stage_4__6563_,data_stage_4__6562_,
  data_stage_4__6561_,data_stage_4__6560_,data_stage_4__6559_,data_stage_4__6558_,
  data_stage_4__6557_,data_stage_4__6556_,data_stage_4__6555_,data_stage_4__6554_,
  data_stage_4__6553_,data_stage_4__6552_,data_stage_4__6551_,data_stage_4__6550_,
  data_stage_4__6549_,data_stage_4__6548_,data_stage_4__6547_,data_stage_4__6546_,
  data_stage_4__6545_,data_stage_4__6544_,data_stage_4__6543_,data_stage_4__6542_,
  data_stage_4__6541_,data_stage_4__6540_,data_stage_4__6539_,data_stage_4__6538_,
  data_stage_4__6537_,data_stage_4__6536_,data_stage_4__6535_,data_stage_4__6534_,
  data_stage_4__6533_,data_stage_4__6532_,data_stage_4__6531_,data_stage_4__6530_,
  data_stage_4__6529_,data_stage_4__6528_,data_stage_4__6527_,data_stage_4__6526_,
  data_stage_4__6525_,data_stage_4__6524_,data_stage_4__6523_,data_stage_4__6522_,
  data_stage_4__6521_,data_stage_4__6520_,data_stage_4__6519_,data_stage_4__6518_,
  data_stage_4__6517_,data_stage_4__6516_,data_stage_4__6515_,data_stage_4__6514_,
  data_stage_4__6513_,data_stage_4__6512_,data_stage_4__6511_,data_stage_4__6510_,
  data_stage_4__6509_,data_stage_4__6508_,data_stage_4__6507_,data_stage_4__6506_,
  data_stage_4__6505_,data_stage_4__6504_,data_stage_4__6503_,data_stage_4__6502_,
  data_stage_4__6501_,data_stage_4__6500_,data_stage_4__6499_,data_stage_4__6498_,
  data_stage_4__6497_,data_stage_4__6496_,data_stage_4__6495_,data_stage_4__6494_,
  data_stage_4__6493_,data_stage_4__6492_,data_stage_4__6491_,data_stage_4__6490_,
  data_stage_4__6489_,data_stage_4__6488_,data_stage_4__6487_,data_stage_4__6486_,
  data_stage_4__6485_,data_stage_4__6484_,data_stage_4__6483_,data_stage_4__6482_,
  data_stage_4__6481_,data_stage_4__6480_,data_stage_4__6479_,data_stage_4__6478_,
  data_stage_4__6477_,data_stage_4__6476_,data_stage_4__6475_,data_stage_4__6474_,
  data_stage_4__6473_,data_stage_4__6472_,data_stage_4__6471_,data_stage_4__6470_,
  data_stage_4__6469_,data_stage_4__6468_,data_stage_4__6467_,data_stage_4__6466_,
  data_stage_4__6465_,data_stage_4__6464_,data_stage_4__6463_,data_stage_4__6462_,
  data_stage_4__6461_,data_stage_4__6460_,data_stage_4__6459_,data_stage_4__6458_,
  data_stage_4__6457_,data_stage_4__6456_,data_stage_4__6455_,data_stage_4__6454_,
  data_stage_4__6453_,data_stage_4__6452_,data_stage_4__6451_,data_stage_4__6450_,
  data_stage_4__6449_,data_stage_4__6448_,data_stage_4__6447_,data_stage_4__6446_,
  data_stage_4__6445_,data_stage_4__6444_,data_stage_4__6443_,data_stage_4__6442_,
  data_stage_4__6441_,data_stage_4__6440_,data_stage_4__6439_,data_stage_4__6438_,
  data_stage_4__6437_,data_stage_4__6436_,data_stage_4__6435_,data_stage_4__6434_,
  data_stage_4__6433_,data_stage_4__6432_,data_stage_4__6431_,data_stage_4__6430_,
  data_stage_4__6429_,data_stage_4__6428_,data_stage_4__6427_,data_stage_4__6426_,
  data_stage_4__6425_,data_stage_4__6424_,data_stage_4__6423_,data_stage_4__6422_,
  data_stage_4__6421_,data_stage_4__6420_,data_stage_4__6419_,data_stage_4__6418_,
  data_stage_4__6417_,data_stage_4__6416_,data_stage_4__6415_,data_stage_4__6414_,
  data_stage_4__6413_,data_stage_4__6412_,data_stage_4__6411_,data_stage_4__6410_,
  data_stage_4__6409_,data_stage_4__6408_,data_stage_4__6407_,data_stage_4__6406_,
  data_stage_4__6405_,data_stage_4__6404_,data_stage_4__6403_,data_stage_4__6402_,
  data_stage_4__6401_,data_stage_4__6400_,data_stage_4__6399_,data_stage_4__6398_,
  data_stage_4__6397_,data_stage_4__6396_,data_stage_4__6395_,data_stage_4__6394_,
  data_stage_4__6393_,data_stage_4__6392_,data_stage_4__6391_,data_stage_4__6390_,
  data_stage_4__6389_,data_stage_4__6388_,data_stage_4__6387_,data_stage_4__6386_,
  data_stage_4__6385_,data_stage_4__6384_,data_stage_4__6383_,data_stage_4__6382_,
  data_stage_4__6381_,data_stage_4__6380_,data_stage_4__6379_,data_stage_4__6378_,
  data_stage_4__6377_,data_stage_4__6376_,data_stage_4__6375_,data_stage_4__6374_,
  data_stage_4__6373_,data_stage_4__6372_,data_stage_4__6371_,data_stage_4__6370_,
  data_stage_4__6369_,data_stage_4__6368_,data_stage_4__6367_,data_stage_4__6366_,
  data_stage_4__6365_,data_stage_4__6364_,data_stage_4__6363_,data_stage_4__6362_,
  data_stage_4__6361_,data_stage_4__6360_,data_stage_4__6359_,data_stage_4__6358_,
  data_stage_4__6357_,data_stage_4__6356_,data_stage_4__6355_,data_stage_4__6354_,
  data_stage_4__6353_,data_stage_4__6352_,data_stage_4__6351_,data_stage_4__6350_,
  data_stage_4__6349_,data_stage_4__6348_,data_stage_4__6347_,data_stage_4__6346_,
  data_stage_4__6345_,data_stage_4__6344_,data_stage_4__6343_,data_stage_4__6342_,
  data_stage_4__6341_,data_stage_4__6340_,data_stage_4__6339_,data_stage_4__6338_,
  data_stage_4__6337_,data_stage_4__6336_,data_stage_4__6335_,data_stage_4__6334_,
  data_stage_4__6333_,data_stage_4__6332_,data_stage_4__6331_,data_stage_4__6330_,
  data_stage_4__6329_,data_stage_4__6328_,data_stage_4__6327_,data_stage_4__6326_,
  data_stage_4__6325_,data_stage_4__6324_,data_stage_4__6323_,data_stage_4__6322_,
  data_stage_4__6321_,data_stage_4__6320_,data_stage_4__6319_,data_stage_4__6318_,
  data_stage_4__6317_,data_stage_4__6316_,data_stage_4__6315_,data_stage_4__6314_,
  data_stage_4__6313_,data_stage_4__6312_,data_stage_4__6311_,data_stage_4__6310_,
  data_stage_4__6309_,data_stage_4__6308_,data_stage_4__6307_,data_stage_4__6306_,
  data_stage_4__6305_,data_stage_4__6304_,data_stage_4__6303_,data_stage_4__6302_,
  data_stage_4__6301_,data_stage_4__6300_,data_stage_4__6299_,data_stage_4__6298_,
  data_stage_4__6297_,data_stage_4__6296_,data_stage_4__6295_,data_stage_4__6294_,
  data_stage_4__6293_,data_stage_4__6292_,data_stage_4__6291_,data_stage_4__6290_,
  data_stage_4__6289_,data_stage_4__6288_,data_stage_4__6287_,data_stage_4__6286_,
  data_stage_4__6285_,data_stage_4__6284_,data_stage_4__6283_,data_stage_4__6282_,
  data_stage_4__6281_,data_stage_4__6280_,data_stage_4__6279_,data_stage_4__6278_,
  data_stage_4__6277_,data_stage_4__6276_,data_stage_4__6275_,data_stage_4__6274_,
  data_stage_4__6273_,data_stage_4__6272_,data_stage_4__6271_,data_stage_4__6270_,
  data_stage_4__6269_,data_stage_4__6268_,data_stage_4__6267_,data_stage_4__6266_,
  data_stage_4__6265_,data_stage_4__6264_,data_stage_4__6263_,data_stage_4__6262_,
  data_stage_4__6261_,data_stage_4__6260_,data_stage_4__6259_,data_stage_4__6258_,
  data_stage_4__6257_,data_stage_4__6256_,data_stage_4__6255_,data_stage_4__6254_,
  data_stage_4__6253_,data_stage_4__6252_,data_stage_4__6251_,data_stage_4__6250_,
  data_stage_4__6249_,data_stage_4__6248_,data_stage_4__6247_,data_stage_4__6246_,
  data_stage_4__6245_,data_stage_4__6244_,data_stage_4__6243_,data_stage_4__6242_,
  data_stage_4__6241_,data_stage_4__6240_,data_stage_4__6239_,data_stage_4__6238_,
  data_stage_4__6237_,data_stage_4__6236_,data_stage_4__6235_,data_stage_4__6234_,
  data_stage_4__6233_,data_stage_4__6232_,data_stage_4__6231_,data_stage_4__6230_,
  data_stage_4__6229_,data_stage_4__6228_,data_stage_4__6227_,data_stage_4__6226_,
  data_stage_4__6225_,data_stage_4__6224_,data_stage_4__6223_,data_stage_4__6222_,
  data_stage_4__6221_,data_stage_4__6220_,data_stage_4__6219_,data_stage_4__6218_,
  data_stage_4__6217_,data_stage_4__6216_,data_stage_4__6215_,data_stage_4__6214_,
  data_stage_4__6213_,data_stage_4__6212_,data_stage_4__6211_,data_stage_4__6210_,
  data_stage_4__6209_,data_stage_4__6208_,data_stage_4__6207_,data_stage_4__6206_,
  data_stage_4__6205_,data_stage_4__6204_,data_stage_4__6203_,data_stage_4__6202_,
  data_stage_4__6201_,data_stage_4__6200_,data_stage_4__6199_,data_stage_4__6198_,
  data_stage_4__6197_,data_stage_4__6196_,data_stage_4__6195_,data_stage_4__6194_,
  data_stage_4__6193_,data_stage_4__6192_,data_stage_4__6191_,data_stage_4__6190_,
  data_stage_4__6189_,data_stage_4__6188_,data_stage_4__6187_,data_stage_4__6186_,
  data_stage_4__6185_,data_stage_4__6184_,data_stage_4__6183_,data_stage_4__6182_,
  data_stage_4__6181_,data_stage_4__6180_,data_stage_4__6179_,data_stage_4__6178_,
  data_stage_4__6177_,data_stage_4__6176_,data_stage_4__6175_,data_stage_4__6174_,
  data_stage_4__6173_,data_stage_4__6172_,data_stage_4__6171_,data_stage_4__6170_,
  data_stage_4__6169_,data_stage_4__6168_,data_stage_4__6167_,data_stage_4__6166_,
  data_stage_4__6165_,data_stage_4__6164_,data_stage_4__6163_,data_stage_4__6162_,
  data_stage_4__6161_,data_stage_4__6160_,data_stage_4__6159_,data_stage_4__6158_,
  data_stage_4__6157_,data_stage_4__6156_,data_stage_4__6155_,data_stage_4__6154_,
  data_stage_4__6153_,data_stage_4__6152_,data_stage_4__6151_,data_stage_4__6150_,
  data_stage_4__6149_,data_stage_4__6148_,data_stage_4__6147_,data_stage_4__6146_,
  data_stage_4__6145_,data_stage_4__6144_,data_stage_4__6143_,data_stage_4__6142_,
  data_stage_4__6141_,data_stage_4__6140_,data_stage_4__6139_,data_stage_4__6138_,
  data_stage_4__6137_,data_stage_4__6136_,data_stage_4__6135_,data_stage_4__6134_,
  data_stage_4__6133_,data_stage_4__6132_,data_stage_4__6131_,data_stage_4__6130_,
  data_stage_4__6129_,data_stage_4__6128_,data_stage_4__6127_,data_stage_4__6126_,
  data_stage_4__6125_,data_stage_4__6124_,data_stage_4__6123_,data_stage_4__6122_,
  data_stage_4__6121_,data_stage_4__6120_,data_stage_4__6119_,data_stage_4__6118_,
  data_stage_4__6117_,data_stage_4__6116_,data_stage_4__6115_,data_stage_4__6114_,
  data_stage_4__6113_,data_stage_4__6112_,data_stage_4__6111_,data_stage_4__6110_,
  data_stage_4__6109_,data_stage_4__6108_,data_stage_4__6107_,data_stage_4__6106_,
  data_stage_4__6105_,data_stage_4__6104_,data_stage_4__6103_,data_stage_4__6102_,
  data_stage_4__6101_,data_stage_4__6100_,data_stage_4__6099_,data_stage_4__6098_,
  data_stage_4__6097_,data_stage_4__6096_,data_stage_4__6095_,data_stage_4__6094_,
  data_stage_4__6093_,data_stage_4__6092_,data_stage_4__6091_,data_stage_4__6090_,
  data_stage_4__6089_,data_stage_4__6088_,data_stage_4__6087_,data_stage_4__6086_,
  data_stage_4__6085_,data_stage_4__6084_,data_stage_4__6083_,data_stage_4__6082_,
  data_stage_4__6081_,data_stage_4__6080_,data_stage_4__6079_,data_stage_4__6078_,
  data_stage_4__6077_,data_stage_4__6076_,data_stage_4__6075_,data_stage_4__6074_,
  data_stage_4__6073_,data_stage_4__6072_,data_stage_4__6071_,data_stage_4__6070_,
  data_stage_4__6069_,data_stage_4__6068_,data_stage_4__6067_,data_stage_4__6066_,
  data_stage_4__6065_,data_stage_4__6064_,data_stage_4__6063_,data_stage_4__6062_,
  data_stage_4__6061_,data_stage_4__6060_,data_stage_4__6059_,data_stage_4__6058_,
  data_stage_4__6057_,data_stage_4__6056_,data_stage_4__6055_,data_stage_4__6054_,
  data_stage_4__6053_,data_stage_4__6052_,data_stage_4__6051_,data_stage_4__6050_,
  data_stage_4__6049_,data_stage_4__6048_,data_stage_4__6047_,data_stage_4__6046_,
  data_stage_4__6045_,data_stage_4__6044_,data_stage_4__6043_,data_stage_4__6042_,
  data_stage_4__6041_,data_stage_4__6040_,data_stage_4__6039_,data_stage_4__6038_,
  data_stage_4__6037_,data_stage_4__6036_,data_stage_4__6035_,data_stage_4__6034_,
  data_stage_4__6033_,data_stage_4__6032_,data_stage_4__6031_,data_stage_4__6030_,
  data_stage_4__6029_,data_stage_4__6028_,data_stage_4__6027_,data_stage_4__6026_,
  data_stage_4__6025_,data_stage_4__6024_,data_stage_4__6023_,data_stage_4__6022_,
  data_stage_4__6021_,data_stage_4__6020_,data_stage_4__6019_,data_stage_4__6018_,
  data_stage_4__6017_,data_stage_4__6016_,data_stage_4__6015_,data_stage_4__6014_,
  data_stage_4__6013_,data_stage_4__6012_,data_stage_4__6011_,data_stage_4__6010_,
  data_stage_4__6009_,data_stage_4__6008_,data_stage_4__6007_,data_stage_4__6006_,
  data_stage_4__6005_,data_stage_4__6004_,data_stage_4__6003_,data_stage_4__6002_,
  data_stage_4__6001_,data_stage_4__6000_,data_stage_4__5999_,data_stage_4__5998_,
  data_stage_4__5997_,data_stage_4__5996_,data_stage_4__5995_,data_stage_4__5994_,
  data_stage_4__5993_,data_stage_4__5992_,data_stage_4__5991_,data_stage_4__5990_,
  data_stage_4__5989_,data_stage_4__5988_,data_stage_4__5987_,data_stage_4__5986_,
  data_stage_4__5985_,data_stage_4__5984_,data_stage_4__5983_,data_stage_4__5982_,
  data_stage_4__5981_,data_stage_4__5980_,data_stage_4__5979_,data_stage_4__5978_,
  data_stage_4__5977_,data_stage_4__5976_,data_stage_4__5975_,data_stage_4__5974_,
  data_stage_4__5973_,data_stage_4__5972_,data_stage_4__5971_,data_stage_4__5970_,
  data_stage_4__5969_,data_stage_4__5968_,data_stage_4__5967_,data_stage_4__5966_,
  data_stage_4__5965_,data_stage_4__5964_,data_stage_4__5963_,data_stage_4__5962_,
  data_stage_4__5961_,data_stage_4__5960_,data_stage_4__5959_,data_stage_4__5958_,
  data_stage_4__5957_,data_stage_4__5956_,data_stage_4__5955_,data_stage_4__5954_,
  data_stage_4__5953_,data_stage_4__5952_,data_stage_4__5951_,data_stage_4__5950_,
  data_stage_4__5949_,data_stage_4__5948_,data_stage_4__5947_,data_stage_4__5946_,
  data_stage_4__5945_,data_stage_4__5944_,data_stage_4__5943_,data_stage_4__5942_,
  data_stage_4__5941_,data_stage_4__5940_,data_stage_4__5939_,data_stage_4__5938_,
  data_stage_4__5937_,data_stage_4__5936_,data_stage_4__5935_,data_stage_4__5934_,
  data_stage_4__5933_,data_stage_4__5932_,data_stage_4__5931_,data_stage_4__5930_,
  data_stage_4__5929_,data_stage_4__5928_,data_stage_4__5927_,data_stage_4__5926_,
  data_stage_4__5925_,data_stage_4__5924_,data_stage_4__5923_,data_stage_4__5922_,
  data_stage_4__5921_,data_stage_4__5920_,data_stage_4__5919_,data_stage_4__5918_,
  data_stage_4__5917_,data_stage_4__5916_,data_stage_4__5915_,data_stage_4__5914_,
  data_stage_4__5913_,data_stage_4__5912_,data_stage_4__5911_,data_stage_4__5910_,
  data_stage_4__5909_,data_stage_4__5908_,data_stage_4__5907_,data_stage_4__5906_,
  data_stage_4__5905_,data_stage_4__5904_,data_stage_4__5903_,data_stage_4__5902_,
  data_stage_4__5901_,data_stage_4__5900_,data_stage_4__5899_,data_stage_4__5898_,
  data_stage_4__5897_,data_stage_4__5896_,data_stage_4__5895_,data_stage_4__5894_,
  data_stage_4__5893_,data_stage_4__5892_,data_stage_4__5891_,data_stage_4__5890_,
  data_stage_4__5889_,data_stage_4__5888_,data_stage_4__5887_,data_stage_4__5886_,
  data_stage_4__5885_,data_stage_4__5884_,data_stage_4__5883_,data_stage_4__5882_,
  data_stage_4__5881_,data_stage_4__5880_,data_stage_4__5879_,data_stage_4__5878_,
  data_stage_4__5877_,data_stage_4__5876_,data_stage_4__5875_,data_stage_4__5874_,
  data_stage_4__5873_,data_stage_4__5872_,data_stage_4__5871_,data_stage_4__5870_,
  data_stage_4__5869_,data_stage_4__5868_,data_stage_4__5867_,data_stage_4__5866_,
  data_stage_4__5865_,data_stage_4__5864_,data_stage_4__5863_,data_stage_4__5862_,
  data_stage_4__5861_,data_stage_4__5860_,data_stage_4__5859_,data_stage_4__5858_,
  data_stage_4__5857_,data_stage_4__5856_,data_stage_4__5855_,data_stage_4__5854_,
  data_stage_4__5853_,data_stage_4__5852_,data_stage_4__5851_,data_stage_4__5850_,
  data_stage_4__5849_,data_stage_4__5848_,data_stage_4__5847_,data_stage_4__5846_,
  data_stage_4__5845_,data_stage_4__5844_,data_stage_4__5843_,data_stage_4__5842_,
  data_stage_4__5841_,data_stage_4__5840_,data_stage_4__5839_,data_stage_4__5838_,
  data_stage_4__5837_,data_stage_4__5836_,data_stage_4__5835_,data_stage_4__5834_,
  data_stage_4__5833_,data_stage_4__5832_,data_stage_4__5831_,data_stage_4__5830_,
  data_stage_4__5829_,data_stage_4__5828_,data_stage_4__5827_,data_stage_4__5826_,
  data_stage_4__5825_,data_stage_4__5824_,data_stage_4__5823_,data_stage_4__5822_,
  data_stage_4__5821_,data_stage_4__5820_,data_stage_4__5819_,data_stage_4__5818_,
  data_stage_4__5817_,data_stage_4__5816_,data_stage_4__5815_,data_stage_4__5814_,
  data_stage_4__5813_,data_stage_4__5812_,data_stage_4__5811_,data_stage_4__5810_,
  data_stage_4__5809_,data_stage_4__5808_,data_stage_4__5807_,data_stage_4__5806_,
  data_stage_4__5805_,data_stage_4__5804_,data_stage_4__5803_,data_stage_4__5802_,
  data_stage_4__5801_,data_stage_4__5800_,data_stage_4__5799_,data_stage_4__5798_,
  data_stage_4__5797_,data_stage_4__5796_,data_stage_4__5795_,data_stage_4__5794_,
  data_stage_4__5793_,data_stage_4__5792_,data_stage_4__5791_,data_stage_4__5790_,
  data_stage_4__5789_,data_stage_4__5788_,data_stage_4__5787_,data_stage_4__5786_,
  data_stage_4__5785_,data_stage_4__5784_,data_stage_4__5783_,data_stage_4__5782_,
  data_stage_4__5781_,data_stage_4__5780_,data_stage_4__5779_,data_stage_4__5778_,
  data_stage_4__5777_,data_stage_4__5776_,data_stage_4__5775_,data_stage_4__5774_,
  data_stage_4__5773_,data_stage_4__5772_,data_stage_4__5771_,data_stage_4__5770_,
  data_stage_4__5769_,data_stage_4__5768_,data_stage_4__5767_,data_stage_4__5766_,
  data_stage_4__5765_,data_stage_4__5764_,data_stage_4__5763_,data_stage_4__5762_,
  data_stage_4__5761_,data_stage_4__5760_,data_stage_4__5759_,data_stage_4__5758_,
  data_stage_4__5757_,data_stage_4__5756_,data_stage_4__5755_,data_stage_4__5754_,
  data_stage_4__5753_,data_stage_4__5752_,data_stage_4__5751_,data_stage_4__5750_,
  data_stage_4__5749_,data_stage_4__5748_,data_stage_4__5747_,data_stage_4__5746_,
  data_stage_4__5745_,data_stage_4__5744_,data_stage_4__5743_,data_stage_4__5742_,
  data_stage_4__5741_,data_stage_4__5740_,data_stage_4__5739_,data_stage_4__5738_,
  data_stage_4__5737_,data_stage_4__5736_,data_stage_4__5735_,data_stage_4__5734_,
  data_stage_4__5733_,data_stage_4__5732_,data_stage_4__5731_,data_stage_4__5730_,
  data_stage_4__5729_,data_stage_4__5728_,data_stage_4__5727_,data_stage_4__5726_,
  data_stage_4__5725_,data_stage_4__5724_,data_stage_4__5723_,data_stage_4__5722_,
  data_stage_4__5721_,data_stage_4__5720_,data_stage_4__5719_,data_stage_4__5718_,
  data_stage_4__5717_,data_stage_4__5716_,data_stage_4__5715_,data_stage_4__5714_,
  data_stage_4__5713_,data_stage_4__5712_,data_stage_4__5711_,data_stage_4__5710_,
  data_stage_4__5709_,data_stage_4__5708_,data_stage_4__5707_,data_stage_4__5706_,
  data_stage_4__5705_,data_stage_4__5704_,data_stage_4__5703_,data_stage_4__5702_,
  data_stage_4__5701_,data_stage_4__5700_,data_stage_4__5699_,data_stage_4__5698_,
  data_stage_4__5697_,data_stage_4__5696_,data_stage_4__5695_,data_stage_4__5694_,
  data_stage_4__5693_,data_stage_4__5692_,data_stage_4__5691_,data_stage_4__5690_,
  data_stage_4__5689_,data_stage_4__5688_,data_stage_4__5687_,data_stage_4__5686_,
  data_stage_4__5685_,data_stage_4__5684_,data_stage_4__5683_,data_stage_4__5682_,
  data_stage_4__5681_,data_stage_4__5680_,data_stage_4__5679_,data_stage_4__5678_,
  data_stage_4__5677_,data_stage_4__5676_,data_stage_4__5675_,data_stage_4__5674_,
  data_stage_4__5673_,data_stage_4__5672_,data_stage_4__5671_,data_stage_4__5670_,
  data_stage_4__5669_,data_stage_4__5668_,data_stage_4__5667_,data_stage_4__5666_,
  data_stage_4__5665_,data_stage_4__5664_,data_stage_4__5663_,data_stage_4__5662_,
  data_stage_4__5661_,data_stage_4__5660_,data_stage_4__5659_,data_stage_4__5658_,
  data_stage_4__5657_,data_stage_4__5656_,data_stage_4__5655_,data_stage_4__5654_,
  data_stage_4__5653_,data_stage_4__5652_,data_stage_4__5651_,data_stage_4__5650_,
  data_stage_4__5649_,data_stage_4__5648_,data_stage_4__5647_,data_stage_4__5646_,
  data_stage_4__5645_,data_stage_4__5644_,data_stage_4__5643_,data_stage_4__5642_,
  data_stage_4__5641_,data_stage_4__5640_,data_stage_4__5639_,data_stage_4__5638_,
  data_stage_4__5637_,data_stage_4__5636_,data_stage_4__5635_,data_stage_4__5634_,
  data_stage_4__5633_,data_stage_4__5632_,data_stage_4__5631_,data_stage_4__5630_,
  data_stage_4__5629_,data_stage_4__5628_,data_stage_4__5627_,data_stage_4__5626_,
  data_stage_4__5625_,data_stage_4__5624_,data_stage_4__5623_,data_stage_4__5622_,
  data_stage_4__5621_,data_stage_4__5620_,data_stage_4__5619_,data_stage_4__5618_,
  data_stage_4__5617_,data_stage_4__5616_,data_stage_4__5615_,data_stage_4__5614_,
  data_stage_4__5613_,data_stage_4__5612_,data_stage_4__5611_,data_stage_4__5610_,
  data_stage_4__5609_,data_stage_4__5608_,data_stage_4__5607_,data_stage_4__5606_,
  data_stage_4__5605_,data_stage_4__5604_,data_stage_4__5603_,data_stage_4__5602_,
  data_stage_4__5601_,data_stage_4__5600_,data_stage_4__5599_,data_stage_4__5598_,
  data_stage_4__5597_,data_stage_4__5596_,data_stage_4__5595_,data_stage_4__5594_,
  data_stage_4__5593_,data_stage_4__5592_,data_stage_4__5591_,data_stage_4__5590_,
  data_stage_4__5589_,data_stage_4__5588_,data_stage_4__5587_,data_stage_4__5586_,
  data_stage_4__5585_,data_stage_4__5584_,data_stage_4__5583_,data_stage_4__5582_,
  data_stage_4__5581_,data_stage_4__5580_,data_stage_4__5579_,data_stage_4__5578_,
  data_stage_4__5577_,data_stage_4__5576_,data_stage_4__5575_,data_stage_4__5574_,
  data_stage_4__5573_,data_stage_4__5572_,data_stage_4__5571_,data_stage_4__5570_,
  data_stage_4__5569_,data_stage_4__5568_,data_stage_4__5567_,data_stage_4__5566_,
  data_stage_4__5565_,data_stage_4__5564_,data_stage_4__5563_,data_stage_4__5562_,
  data_stage_4__5561_,data_stage_4__5560_,data_stage_4__5559_,data_stage_4__5558_,
  data_stage_4__5557_,data_stage_4__5556_,data_stage_4__5555_,data_stage_4__5554_,
  data_stage_4__5553_,data_stage_4__5552_,data_stage_4__5551_,data_stage_4__5550_,
  data_stage_4__5549_,data_stage_4__5548_,data_stage_4__5547_,data_stage_4__5546_,
  data_stage_4__5545_,data_stage_4__5544_,data_stage_4__5543_,data_stage_4__5542_,
  data_stage_4__5541_,data_stage_4__5540_,data_stage_4__5539_,data_stage_4__5538_,
  data_stage_4__5537_,data_stage_4__5536_,data_stage_4__5535_,data_stage_4__5534_,
  data_stage_4__5533_,data_stage_4__5532_,data_stage_4__5531_,data_stage_4__5530_,
  data_stage_4__5529_,data_stage_4__5528_,data_stage_4__5527_,data_stage_4__5526_,
  data_stage_4__5525_,data_stage_4__5524_,data_stage_4__5523_,data_stage_4__5522_,
  data_stage_4__5521_,data_stage_4__5520_,data_stage_4__5519_,data_stage_4__5518_,
  data_stage_4__5517_,data_stage_4__5516_,data_stage_4__5515_,data_stage_4__5514_,
  data_stage_4__5513_,data_stage_4__5512_,data_stage_4__5511_,data_stage_4__5510_,
  data_stage_4__5509_,data_stage_4__5508_,data_stage_4__5507_,data_stage_4__5506_,
  data_stage_4__5505_,data_stage_4__5504_,data_stage_4__5503_,data_stage_4__5502_,
  data_stage_4__5501_,data_stage_4__5500_,data_stage_4__5499_,data_stage_4__5498_,
  data_stage_4__5497_,data_stage_4__5496_,data_stage_4__5495_,data_stage_4__5494_,
  data_stage_4__5493_,data_stage_4__5492_,data_stage_4__5491_,data_stage_4__5490_,
  data_stage_4__5489_,data_stage_4__5488_,data_stage_4__5487_,data_stage_4__5486_,
  data_stage_4__5485_,data_stage_4__5484_,data_stage_4__5483_,data_stage_4__5482_,
  data_stage_4__5481_,data_stage_4__5480_,data_stage_4__5479_,data_stage_4__5478_,
  data_stage_4__5477_,data_stage_4__5476_,data_stage_4__5475_,data_stage_4__5474_,
  data_stage_4__5473_,data_stage_4__5472_,data_stage_4__5471_,data_stage_4__5470_,
  data_stage_4__5469_,data_stage_4__5468_,data_stage_4__5467_,data_stage_4__5466_,
  data_stage_4__5465_,data_stage_4__5464_,data_stage_4__5463_,data_stage_4__5462_,
  data_stage_4__5461_,data_stage_4__5460_,data_stage_4__5459_,data_stage_4__5458_,
  data_stage_4__5457_,data_stage_4__5456_,data_stage_4__5455_,data_stage_4__5454_,
  data_stage_4__5453_,data_stage_4__5452_,data_stage_4__5451_,data_stage_4__5450_,
  data_stage_4__5449_,data_stage_4__5448_,data_stage_4__5447_,data_stage_4__5446_,
  data_stage_4__5445_,data_stage_4__5444_,data_stage_4__5443_,data_stage_4__5442_,
  data_stage_4__5441_,data_stage_4__5440_,data_stage_4__5439_,data_stage_4__5438_,
  data_stage_4__5437_,data_stage_4__5436_,data_stage_4__5435_,data_stage_4__5434_,
  data_stage_4__5433_,data_stage_4__5432_,data_stage_4__5431_,data_stage_4__5430_,
  data_stage_4__5429_,data_stage_4__5428_,data_stage_4__5427_,data_stage_4__5426_,
  data_stage_4__5425_,data_stage_4__5424_,data_stage_4__5423_,data_stage_4__5422_,
  data_stage_4__5421_,data_stage_4__5420_,data_stage_4__5419_,data_stage_4__5418_,
  data_stage_4__5417_,data_stage_4__5416_,data_stage_4__5415_,data_stage_4__5414_,
  data_stage_4__5413_,data_stage_4__5412_,data_stage_4__5411_,data_stage_4__5410_,
  data_stage_4__5409_,data_stage_4__5408_,data_stage_4__5407_,data_stage_4__5406_,
  data_stage_4__5405_,data_stage_4__5404_,data_stage_4__5403_,data_stage_4__5402_,
  data_stage_4__5401_,data_stage_4__5400_,data_stage_4__5399_,data_stage_4__5398_,
  data_stage_4__5397_,data_stage_4__5396_,data_stage_4__5395_,data_stage_4__5394_,
  data_stage_4__5393_,data_stage_4__5392_,data_stage_4__5391_,data_stage_4__5390_,
  data_stage_4__5389_,data_stage_4__5388_,data_stage_4__5387_,data_stage_4__5386_,
  data_stage_4__5385_,data_stage_4__5384_,data_stage_4__5383_,data_stage_4__5382_,
  data_stage_4__5381_,data_stage_4__5380_,data_stage_4__5379_,data_stage_4__5378_,
  data_stage_4__5377_,data_stage_4__5376_,data_stage_4__5375_,data_stage_4__5374_,
  data_stage_4__5373_,data_stage_4__5372_,data_stage_4__5371_,data_stage_4__5370_,
  data_stage_4__5369_,data_stage_4__5368_,data_stage_4__5367_,data_stage_4__5366_,
  data_stage_4__5365_,data_stage_4__5364_,data_stage_4__5363_,data_stage_4__5362_,
  data_stage_4__5361_,data_stage_4__5360_,data_stage_4__5359_,data_stage_4__5358_,
  data_stage_4__5357_,data_stage_4__5356_,data_stage_4__5355_,data_stage_4__5354_,
  data_stage_4__5353_,data_stage_4__5352_,data_stage_4__5351_,data_stage_4__5350_,
  data_stage_4__5349_,data_stage_4__5348_,data_stage_4__5347_,data_stage_4__5346_,
  data_stage_4__5345_,data_stage_4__5344_,data_stage_4__5343_,data_stage_4__5342_,
  data_stage_4__5341_,data_stage_4__5340_,data_stage_4__5339_,data_stage_4__5338_,
  data_stage_4__5337_,data_stage_4__5336_,data_stage_4__5335_,data_stage_4__5334_,
  data_stage_4__5333_,data_stage_4__5332_,data_stage_4__5331_,data_stage_4__5330_,
  data_stage_4__5329_,data_stage_4__5328_,data_stage_4__5327_,data_stage_4__5326_,
  data_stage_4__5325_,data_stage_4__5324_,data_stage_4__5323_,data_stage_4__5322_,
  data_stage_4__5321_,data_stage_4__5320_,data_stage_4__5319_,data_stage_4__5318_,
  data_stage_4__5317_,data_stage_4__5316_,data_stage_4__5315_,data_stage_4__5314_,
  data_stage_4__5313_,data_stage_4__5312_,data_stage_4__5311_,data_stage_4__5310_,
  data_stage_4__5309_,data_stage_4__5308_,data_stage_4__5307_,data_stage_4__5306_,
  data_stage_4__5305_,data_stage_4__5304_,data_stage_4__5303_,data_stage_4__5302_,
  data_stage_4__5301_,data_stage_4__5300_,data_stage_4__5299_,data_stage_4__5298_,
  data_stage_4__5297_,data_stage_4__5296_,data_stage_4__5295_,data_stage_4__5294_,
  data_stage_4__5293_,data_stage_4__5292_,data_stage_4__5291_,data_stage_4__5290_,
  data_stage_4__5289_,data_stage_4__5288_,data_stage_4__5287_,data_stage_4__5286_,
  data_stage_4__5285_,data_stage_4__5284_,data_stage_4__5283_,data_stage_4__5282_,
  data_stage_4__5281_,data_stage_4__5280_,data_stage_4__5279_,data_stage_4__5278_,
  data_stage_4__5277_,data_stage_4__5276_,data_stage_4__5275_,data_stage_4__5274_,
  data_stage_4__5273_,data_stage_4__5272_,data_stage_4__5271_,data_stage_4__5270_,
  data_stage_4__5269_,data_stage_4__5268_,data_stage_4__5267_,data_stage_4__5266_,
  data_stage_4__5265_,data_stage_4__5264_,data_stage_4__5263_,data_stage_4__5262_,
  data_stage_4__5261_,data_stage_4__5260_,data_stage_4__5259_,data_stage_4__5258_,
  data_stage_4__5257_,data_stage_4__5256_,data_stage_4__5255_,data_stage_4__5254_,
  data_stage_4__5253_,data_stage_4__5252_,data_stage_4__5251_,data_stage_4__5250_,
  data_stage_4__5249_,data_stage_4__5248_,data_stage_4__5247_,data_stage_4__5246_,
  data_stage_4__5245_,data_stage_4__5244_,data_stage_4__5243_,data_stage_4__5242_,
  data_stage_4__5241_,data_stage_4__5240_,data_stage_4__5239_,data_stage_4__5238_,
  data_stage_4__5237_,data_stage_4__5236_,data_stage_4__5235_,data_stage_4__5234_,
  data_stage_4__5233_,data_stage_4__5232_,data_stage_4__5231_,data_stage_4__5230_,
  data_stage_4__5229_,data_stage_4__5228_,data_stage_4__5227_,data_stage_4__5226_,
  data_stage_4__5225_,data_stage_4__5224_,data_stage_4__5223_,data_stage_4__5222_,
  data_stage_4__5221_,data_stage_4__5220_,data_stage_4__5219_,data_stage_4__5218_,
  data_stage_4__5217_,data_stage_4__5216_,data_stage_4__5215_,data_stage_4__5214_,
  data_stage_4__5213_,data_stage_4__5212_,data_stage_4__5211_,data_stage_4__5210_,
  data_stage_4__5209_,data_stage_4__5208_,data_stage_4__5207_,data_stage_4__5206_,
  data_stage_4__5205_,data_stage_4__5204_,data_stage_4__5203_,data_stage_4__5202_,
  data_stage_4__5201_,data_stage_4__5200_,data_stage_4__5199_,data_stage_4__5198_,
  data_stage_4__5197_,data_stage_4__5196_,data_stage_4__5195_,data_stage_4__5194_,
  data_stage_4__5193_,data_stage_4__5192_,data_stage_4__5191_,data_stage_4__5190_,
  data_stage_4__5189_,data_stage_4__5188_,data_stage_4__5187_,data_stage_4__5186_,
  data_stage_4__5185_,data_stage_4__5184_,data_stage_4__5183_,data_stage_4__5182_,
  data_stage_4__5181_,data_stage_4__5180_,data_stage_4__5179_,data_stage_4__5178_,
  data_stage_4__5177_,data_stage_4__5176_,data_stage_4__5175_,data_stage_4__5174_,
  data_stage_4__5173_,data_stage_4__5172_,data_stage_4__5171_,data_stage_4__5170_,
  data_stage_4__5169_,data_stage_4__5168_,data_stage_4__5167_,data_stage_4__5166_,
  data_stage_4__5165_,data_stage_4__5164_,data_stage_4__5163_,data_stage_4__5162_,
  data_stage_4__5161_,data_stage_4__5160_,data_stage_4__5159_,data_stage_4__5158_,
  data_stage_4__5157_,data_stage_4__5156_,data_stage_4__5155_,data_stage_4__5154_,
  data_stage_4__5153_,data_stage_4__5152_,data_stage_4__5151_,data_stage_4__5150_,
  data_stage_4__5149_,data_stage_4__5148_,data_stage_4__5147_,data_stage_4__5146_,
  data_stage_4__5145_,data_stage_4__5144_,data_stage_4__5143_,data_stage_4__5142_,
  data_stage_4__5141_,data_stage_4__5140_,data_stage_4__5139_,data_stage_4__5138_,
  data_stage_4__5137_,data_stage_4__5136_,data_stage_4__5135_,data_stage_4__5134_,
  data_stage_4__5133_,data_stage_4__5132_,data_stage_4__5131_,data_stage_4__5130_,
  data_stage_4__5129_,data_stage_4__5128_,data_stage_4__5127_,data_stage_4__5126_,
  data_stage_4__5125_,data_stage_4__5124_,data_stage_4__5123_,data_stage_4__5122_,
  data_stage_4__5121_,data_stage_4__5120_,data_stage_4__5119_,data_stage_4__5118_,
  data_stage_4__5117_,data_stage_4__5116_,data_stage_4__5115_,data_stage_4__5114_,
  data_stage_4__5113_,data_stage_4__5112_,data_stage_4__5111_,data_stage_4__5110_,
  data_stage_4__5109_,data_stage_4__5108_,data_stage_4__5107_,data_stage_4__5106_,
  data_stage_4__5105_,data_stage_4__5104_,data_stage_4__5103_,data_stage_4__5102_,
  data_stage_4__5101_,data_stage_4__5100_,data_stage_4__5099_,data_stage_4__5098_,
  data_stage_4__5097_,data_stage_4__5096_,data_stage_4__5095_,data_stage_4__5094_,
  data_stage_4__5093_,data_stage_4__5092_,data_stage_4__5091_,data_stage_4__5090_,
  data_stage_4__5089_,data_stage_4__5088_,data_stage_4__5087_,data_stage_4__5086_,
  data_stage_4__5085_,data_stage_4__5084_,data_stage_4__5083_,data_stage_4__5082_,
  data_stage_4__5081_,data_stage_4__5080_,data_stage_4__5079_,data_stage_4__5078_,
  data_stage_4__5077_,data_stage_4__5076_,data_stage_4__5075_,data_stage_4__5074_,
  data_stage_4__5073_,data_stage_4__5072_,data_stage_4__5071_,data_stage_4__5070_,
  data_stage_4__5069_,data_stage_4__5068_,data_stage_4__5067_,data_stage_4__5066_,
  data_stage_4__5065_,data_stage_4__5064_,data_stage_4__5063_,data_stage_4__5062_,
  data_stage_4__5061_,data_stage_4__5060_,data_stage_4__5059_,data_stage_4__5058_,
  data_stage_4__5057_,data_stage_4__5056_,data_stage_4__5055_,data_stage_4__5054_,
  data_stage_4__5053_,data_stage_4__5052_,data_stage_4__5051_,data_stage_4__5050_,
  data_stage_4__5049_,data_stage_4__5048_,data_stage_4__5047_,data_stage_4__5046_,
  data_stage_4__5045_,data_stage_4__5044_,data_stage_4__5043_,data_stage_4__5042_,
  data_stage_4__5041_,data_stage_4__5040_,data_stage_4__5039_,data_stage_4__5038_,
  data_stage_4__5037_,data_stage_4__5036_,data_stage_4__5035_,data_stage_4__5034_,
  data_stage_4__5033_,data_stage_4__5032_,data_stage_4__5031_,data_stage_4__5030_,
  data_stage_4__5029_,data_stage_4__5028_,data_stage_4__5027_,data_stage_4__5026_,
  data_stage_4__5025_,data_stage_4__5024_,data_stage_4__5023_,data_stage_4__5022_,
  data_stage_4__5021_,data_stage_4__5020_,data_stage_4__5019_,data_stage_4__5018_,
  data_stage_4__5017_,data_stage_4__5016_,data_stage_4__5015_,data_stage_4__5014_,
  data_stage_4__5013_,data_stage_4__5012_,data_stage_4__5011_,data_stage_4__5010_,
  data_stage_4__5009_,data_stage_4__5008_,data_stage_4__5007_,data_stage_4__5006_,
  data_stage_4__5005_,data_stage_4__5004_,data_stage_4__5003_,data_stage_4__5002_,
  data_stage_4__5001_,data_stage_4__5000_,data_stage_4__4999_,data_stage_4__4998_,
  data_stage_4__4997_,data_stage_4__4996_,data_stage_4__4995_,data_stage_4__4994_,
  data_stage_4__4993_,data_stage_4__4992_,data_stage_4__4991_,data_stage_4__4990_,
  data_stage_4__4989_,data_stage_4__4988_,data_stage_4__4987_,data_stage_4__4986_,
  data_stage_4__4985_,data_stage_4__4984_,data_stage_4__4983_,data_stage_4__4982_,
  data_stage_4__4981_,data_stage_4__4980_,data_stage_4__4979_,data_stage_4__4978_,
  data_stage_4__4977_,data_stage_4__4976_,data_stage_4__4975_,data_stage_4__4974_,
  data_stage_4__4973_,data_stage_4__4972_,data_stage_4__4971_,data_stage_4__4970_,
  data_stage_4__4969_,data_stage_4__4968_,data_stage_4__4967_,data_stage_4__4966_,
  data_stage_4__4965_,data_stage_4__4964_,data_stage_4__4963_,data_stage_4__4962_,
  data_stage_4__4961_,data_stage_4__4960_,data_stage_4__4959_,data_stage_4__4958_,
  data_stage_4__4957_,data_stage_4__4956_,data_stage_4__4955_,data_stage_4__4954_,
  data_stage_4__4953_,data_stage_4__4952_,data_stage_4__4951_,data_stage_4__4950_,
  data_stage_4__4949_,data_stage_4__4948_,data_stage_4__4947_,data_stage_4__4946_,
  data_stage_4__4945_,data_stage_4__4944_,data_stage_4__4943_,data_stage_4__4942_,
  data_stage_4__4941_,data_stage_4__4940_,data_stage_4__4939_,data_stage_4__4938_,
  data_stage_4__4937_,data_stage_4__4936_,data_stage_4__4935_,data_stage_4__4934_,
  data_stage_4__4933_,data_stage_4__4932_,data_stage_4__4931_,data_stage_4__4930_,
  data_stage_4__4929_,data_stage_4__4928_,data_stage_4__4927_,data_stage_4__4926_,
  data_stage_4__4925_,data_stage_4__4924_,data_stage_4__4923_,data_stage_4__4922_,
  data_stage_4__4921_,data_stage_4__4920_,data_stage_4__4919_,data_stage_4__4918_,
  data_stage_4__4917_,data_stage_4__4916_,data_stage_4__4915_,data_stage_4__4914_,
  data_stage_4__4913_,data_stage_4__4912_,data_stage_4__4911_,data_stage_4__4910_,
  data_stage_4__4909_,data_stage_4__4908_,data_stage_4__4907_,data_stage_4__4906_,
  data_stage_4__4905_,data_stage_4__4904_,data_stage_4__4903_,data_stage_4__4902_,
  data_stage_4__4901_,data_stage_4__4900_,data_stage_4__4899_,data_stage_4__4898_,
  data_stage_4__4897_,data_stage_4__4896_,data_stage_4__4895_,data_stage_4__4894_,
  data_stage_4__4893_,data_stage_4__4892_,data_stage_4__4891_,data_stage_4__4890_,
  data_stage_4__4889_,data_stage_4__4888_,data_stage_4__4887_,data_stage_4__4886_,
  data_stage_4__4885_,data_stage_4__4884_,data_stage_4__4883_,data_stage_4__4882_,
  data_stage_4__4881_,data_stage_4__4880_,data_stage_4__4879_,data_stage_4__4878_,
  data_stage_4__4877_,data_stage_4__4876_,data_stage_4__4875_,data_stage_4__4874_,
  data_stage_4__4873_,data_stage_4__4872_,data_stage_4__4871_,data_stage_4__4870_,
  data_stage_4__4869_,data_stage_4__4868_,data_stage_4__4867_,data_stage_4__4866_,
  data_stage_4__4865_,data_stage_4__4864_,data_stage_4__4863_,data_stage_4__4862_,
  data_stage_4__4861_,data_stage_4__4860_,data_stage_4__4859_,data_stage_4__4858_,
  data_stage_4__4857_,data_stage_4__4856_,data_stage_4__4855_,data_stage_4__4854_,
  data_stage_4__4853_,data_stage_4__4852_,data_stage_4__4851_,data_stage_4__4850_,
  data_stage_4__4849_,data_stage_4__4848_,data_stage_4__4847_,data_stage_4__4846_,
  data_stage_4__4845_,data_stage_4__4844_,data_stage_4__4843_,data_stage_4__4842_,
  data_stage_4__4841_,data_stage_4__4840_,data_stage_4__4839_,data_stage_4__4838_,
  data_stage_4__4837_,data_stage_4__4836_,data_stage_4__4835_,data_stage_4__4834_,
  data_stage_4__4833_,data_stage_4__4832_,data_stage_4__4831_,data_stage_4__4830_,
  data_stage_4__4829_,data_stage_4__4828_,data_stage_4__4827_,data_stage_4__4826_,
  data_stage_4__4825_,data_stage_4__4824_,data_stage_4__4823_,data_stage_4__4822_,
  data_stage_4__4821_,data_stage_4__4820_,data_stage_4__4819_,data_stage_4__4818_,
  data_stage_4__4817_,data_stage_4__4816_,data_stage_4__4815_,data_stage_4__4814_,
  data_stage_4__4813_,data_stage_4__4812_,data_stage_4__4811_,data_stage_4__4810_,
  data_stage_4__4809_,data_stage_4__4808_,data_stage_4__4807_,data_stage_4__4806_,
  data_stage_4__4805_,data_stage_4__4804_,data_stage_4__4803_,data_stage_4__4802_,
  data_stage_4__4801_,data_stage_4__4800_,data_stage_4__4799_,data_stage_4__4798_,
  data_stage_4__4797_,data_stage_4__4796_,data_stage_4__4795_,data_stage_4__4794_,
  data_stage_4__4793_,data_stage_4__4792_,data_stage_4__4791_,data_stage_4__4790_,
  data_stage_4__4789_,data_stage_4__4788_,data_stage_4__4787_,data_stage_4__4786_,
  data_stage_4__4785_,data_stage_4__4784_,data_stage_4__4783_,data_stage_4__4782_,
  data_stage_4__4781_,data_stage_4__4780_,data_stage_4__4779_,data_stage_4__4778_,
  data_stage_4__4777_,data_stage_4__4776_,data_stage_4__4775_,data_stage_4__4774_,
  data_stage_4__4773_,data_stage_4__4772_,data_stage_4__4771_,data_stage_4__4770_,
  data_stage_4__4769_,data_stage_4__4768_,data_stage_4__4767_,data_stage_4__4766_,
  data_stage_4__4765_,data_stage_4__4764_,data_stage_4__4763_,data_stage_4__4762_,
  data_stage_4__4761_,data_stage_4__4760_,data_stage_4__4759_,data_stage_4__4758_,
  data_stage_4__4757_,data_stage_4__4756_,data_stage_4__4755_,data_stage_4__4754_,
  data_stage_4__4753_,data_stage_4__4752_,data_stage_4__4751_,data_stage_4__4750_,
  data_stage_4__4749_,data_stage_4__4748_,data_stage_4__4747_,data_stage_4__4746_,
  data_stage_4__4745_,data_stage_4__4744_,data_stage_4__4743_,data_stage_4__4742_,
  data_stage_4__4741_,data_stage_4__4740_,data_stage_4__4739_,data_stage_4__4738_,
  data_stage_4__4737_,data_stage_4__4736_,data_stage_4__4735_,data_stage_4__4734_,
  data_stage_4__4733_,data_stage_4__4732_,data_stage_4__4731_,data_stage_4__4730_,
  data_stage_4__4729_,data_stage_4__4728_,data_stage_4__4727_,data_stage_4__4726_,
  data_stage_4__4725_,data_stage_4__4724_,data_stage_4__4723_,data_stage_4__4722_,
  data_stage_4__4721_,data_stage_4__4720_,data_stage_4__4719_,data_stage_4__4718_,
  data_stage_4__4717_,data_stage_4__4716_,data_stage_4__4715_,data_stage_4__4714_,
  data_stage_4__4713_,data_stage_4__4712_,data_stage_4__4711_,data_stage_4__4710_,
  data_stage_4__4709_,data_stage_4__4708_,data_stage_4__4707_,data_stage_4__4706_,
  data_stage_4__4705_,data_stage_4__4704_,data_stage_4__4703_,data_stage_4__4702_,
  data_stage_4__4701_,data_stage_4__4700_,data_stage_4__4699_,data_stage_4__4698_,
  data_stage_4__4697_,data_stage_4__4696_,data_stage_4__4695_,data_stage_4__4694_,
  data_stage_4__4693_,data_stage_4__4692_,data_stage_4__4691_,data_stage_4__4690_,
  data_stage_4__4689_,data_stage_4__4688_,data_stage_4__4687_,data_stage_4__4686_,
  data_stage_4__4685_,data_stage_4__4684_,data_stage_4__4683_,data_stage_4__4682_,
  data_stage_4__4681_,data_stage_4__4680_,data_stage_4__4679_,data_stage_4__4678_,
  data_stage_4__4677_,data_stage_4__4676_,data_stage_4__4675_,data_stage_4__4674_,
  data_stage_4__4673_,data_stage_4__4672_,data_stage_4__4671_,data_stage_4__4670_,
  data_stage_4__4669_,data_stage_4__4668_,data_stage_4__4667_,data_stage_4__4666_,
  data_stage_4__4665_,data_stage_4__4664_,data_stage_4__4663_,data_stage_4__4662_,
  data_stage_4__4661_,data_stage_4__4660_,data_stage_4__4659_,data_stage_4__4658_,
  data_stage_4__4657_,data_stage_4__4656_,data_stage_4__4655_,data_stage_4__4654_,
  data_stage_4__4653_,data_stage_4__4652_,data_stage_4__4651_,data_stage_4__4650_,
  data_stage_4__4649_,data_stage_4__4648_,data_stage_4__4647_,data_stage_4__4646_,
  data_stage_4__4645_,data_stage_4__4644_,data_stage_4__4643_,data_stage_4__4642_,
  data_stage_4__4641_,data_stage_4__4640_,data_stage_4__4639_,data_stage_4__4638_,
  data_stage_4__4637_,data_stage_4__4636_,data_stage_4__4635_,data_stage_4__4634_,
  data_stage_4__4633_,data_stage_4__4632_,data_stage_4__4631_,data_stage_4__4630_,
  data_stage_4__4629_,data_stage_4__4628_,data_stage_4__4627_,data_stage_4__4626_,
  data_stage_4__4625_,data_stage_4__4624_,data_stage_4__4623_,data_stage_4__4622_,
  data_stage_4__4621_,data_stage_4__4620_,data_stage_4__4619_,data_stage_4__4618_,
  data_stage_4__4617_,data_stage_4__4616_,data_stage_4__4615_,data_stage_4__4614_,
  data_stage_4__4613_,data_stage_4__4612_,data_stage_4__4611_,data_stage_4__4610_,
  data_stage_4__4609_,data_stage_4__4608_,data_stage_4__4607_,data_stage_4__4606_,
  data_stage_4__4605_,data_stage_4__4604_,data_stage_4__4603_,data_stage_4__4602_,
  data_stage_4__4601_,data_stage_4__4600_,data_stage_4__4599_,data_stage_4__4598_,
  data_stage_4__4597_,data_stage_4__4596_,data_stage_4__4595_,data_stage_4__4594_,
  data_stage_4__4593_,data_stage_4__4592_,data_stage_4__4591_,data_stage_4__4590_,
  data_stage_4__4589_,data_stage_4__4588_,data_stage_4__4587_,data_stage_4__4586_,
  data_stage_4__4585_,data_stage_4__4584_,data_stage_4__4583_,data_stage_4__4582_,
  data_stage_4__4581_,data_stage_4__4580_,data_stage_4__4579_,data_stage_4__4578_,
  data_stage_4__4577_,data_stage_4__4576_,data_stage_4__4575_,data_stage_4__4574_,
  data_stage_4__4573_,data_stage_4__4572_,data_stage_4__4571_,data_stage_4__4570_,
  data_stage_4__4569_,data_stage_4__4568_,data_stage_4__4567_,data_stage_4__4566_,
  data_stage_4__4565_,data_stage_4__4564_,data_stage_4__4563_,data_stage_4__4562_,
  data_stage_4__4561_,data_stage_4__4560_,data_stage_4__4559_,data_stage_4__4558_,
  data_stage_4__4557_,data_stage_4__4556_,data_stage_4__4555_,data_stage_4__4554_,
  data_stage_4__4553_,data_stage_4__4552_,data_stage_4__4551_,data_stage_4__4550_,
  data_stage_4__4549_,data_stage_4__4548_,data_stage_4__4547_,data_stage_4__4546_,
  data_stage_4__4545_,data_stage_4__4544_,data_stage_4__4543_,data_stage_4__4542_,
  data_stage_4__4541_,data_stage_4__4540_,data_stage_4__4539_,data_stage_4__4538_,
  data_stage_4__4537_,data_stage_4__4536_,data_stage_4__4535_,data_stage_4__4534_,
  data_stage_4__4533_,data_stage_4__4532_,data_stage_4__4531_,data_stage_4__4530_,
  data_stage_4__4529_,data_stage_4__4528_,data_stage_4__4527_,data_stage_4__4526_,
  data_stage_4__4525_,data_stage_4__4524_,data_stage_4__4523_,data_stage_4__4522_,
  data_stage_4__4521_,data_stage_4__4520_,data_stage_4__4519_,data_stage_4__4518_,
  data_stage_4__4517_,data_stage_4__4516_,data_stage_4__4515_,data_stage_4__4514_,
  data_stage_4__4513_,data_stage_4__4512_,data_stage_4__4511_,data_stage_4__4510_,
  data_stage_4__4509_,data_stage_4__4508_,data_stage_4__4507_,data_stage_4__4506_,
  data_stage_4__4505_,data_stage_4__4504_,data_stage_4__4503_,data_stage_4__4502_,
  data_stage_4__4501_,data_stage_4__4500_,data_stage_4__4499_,data_stage_4__4498_,
  data_stage_4__4497_,data_stage_4__4496_,data_stage_4__4495_,data_stage_4__4494_,
  data_stage_4__4493_,data_stage_4__4492_,data_stage_4__4491_,data_stage_4__4490_,
  data_stage_4__4489_,data_stage_4__4488_,data_stage_4__4487_,data_stage_4__4486_,
  data_stage_4__4485_,data_stage_4__4484_,data_stage_4__4483_,data_stage_4__4482_,
  data_stage_4__4481_,data_stage_4__4480_,data_stage_4__4479_,data_stage_4__4478_,
  data_stage_4__4477_,data_stage_4__4476_,data_stage_4__4475_,data_stage_4__4474_,
  data_stage_4__4473_,data_stage_4__4472_,data_stage_4__4471_,data_stage_4__4470_,
  data_stage_4__4469_,data_stage_4__4468_,data_stage_4__4467_,data_stage_4__4466_,
  data_stage_4__4465_,data_stage_4__4464_,data_stage_4__4463_,data_stage_4__4462_,
  data_stage_4__4461_,data_stage_4__4460_,data_stage_4__4459_,data_stage_4__4458_,
  data_stage_4__4457_,data_stage_4__4456_,data_stage_4__4455_,data_stage_4__4454_,
  data_stage_4__4453_,data_stage_4__4452_,data_stage_4__4451_,data_stage_4__4450_,
  data_stage_4__4449_,data_stage_4__4448_,data_stage_4__4447_,data_stage_4__4446_,
  data_stage_4__4445_,data_stage_4__4444_,data_stage_4__4443_,data_stage_4__4442_,
  data_stage_4__4441_,data_stage_4__4440_,data_stage_4__4439_,data_stage_4__4438_,
  data_stage_4__4437_,data_stage_4__4436_,data_stage_4__4435_,data_stage_4__4434_,
  data_stage_4__4433_,data_stage_4__4432_,data_stage_4__4431_,data_stage_4__4430_,
  data_stage_4__4429_,data_stage_4__4428_,data_stage_4__4427_,data_stage_4__4426_,
  data_stage_4__4425_,data_stage_4__4424_,data_stage_4__4423_,data_stage_4__4422_,
  data_stage_4__4421_,data_stage_4__4420_,data_stage_4__4419_,data_stage_4__4418_,
  data_stage_4__4417_,data_stage_4__4416_,data_stage_4__4415_,data_stage_4__4414_,
  data_stage_4__4413_,data_stage_4__4412_,data_stage_4__4411_,data_stage_4__4410_,
  data_stage_4__4409_,data_stage_4__4408_,data_stage_4__4407_,data_stage_4__4406_,
  data_stage_4__4405_,data_stage_4__4404_,data_stage_4__4403_,data_stage_4__4402_,
  data_stage_4__4401_,data_stage_4__4400_,data_stage_4__4399_,data_stage_4__4398_,
  data_stage_4__4397_,data_stage_4__4396_,data_stage_4__4395_,data_stage_4__4394_,
  data_stage_4__4393_,data_stage_4__4392_,data_stage_4__4391_,data_stage_4__4390_,
  data_stage_4__4389_,data_stage_4__4388_,data_stage_4__4387_,data_stage_4__4386_,
  data_stage_4__4385_,data_stage_4__4384_,data_stage_4__4383_,data_stage_4__4382_,
  data_stage_4__4381_,data_stage_4__4380_,data_stage_4__4379_,data_stage_4__4378_,
  data_stage_4__4377_,data_stage_4__4376_,data_stage_4__4375_,data_stage_4__4374_,
  data_stage_4__4373_,data_stage_4__4372_,data_stage_4__4371_,data_stage_4__4370_,
  data_stage_4__4369_,data_stage_4__4368_,data_stage_4__4367_,data_stage_4__4366_,
  data_stage_4__4365_,data_stage_4__4364_,data_stage_4__4363_,data_stage_4__4362_,
  data_stage_4__4361_,data_stage_4__4360_,data_stage_4__4359_,data_stage_4__4358_,
  data_stage_4__4357_,data_stage_4__4356_,data_stage_4__4355_,data_stage_4__4354_,
  data_stage_4__4353_,data_stage_4__4352_,data_stage_4__4351_,data_stage_4__4350_,
  data_stage_4__4349_,data_stage_4__4348_,data_stage_4__4347_,data_stage_4__4346_,
  data_stage_4__4345_,data_stage_4__4344_,data_stage_4__4343_,data_stage_4__4342_,
  data_stage_4__4341_,data_stage_4__4340_,data_stage_4__4339_,data_stage_4__4338_,
  data_stage_4__4337_,data_stage_4__4336_,data_stage_4__4335_,data_stage_4__4334_,
  data_stage_4__4333_,data_stage_4__4332_,data_stage_4__4331_,data_stage_4__4330_,
  data_stage_4__4329_,data_stage_4__4328_,data_stage_4__4327_,data_stage_4__4326_,
  data_stage_4__4325_,data_stage_4__4324_,data_stage_4__4323_,data_stage_4__4322_,
  data_stage_4__4321_,data_stage_4__4320_,data_stage_4__4319_,data_stage_4__4318_,
  data_stage_4__4317_,data_stage_4__4316_,data_stage_4__4315_,data_stage_4__4314_,
  data_stage_4__4313_,data_stage_4__4312_,data_stage_4__4311_,data_stage_4__4310_,
  data_stage_4__4309_,data_stage_4__4308_,data_stage_4__4307_,data_stage_4__4306_,
  data_stage_4__4305_,data_stage_4__4304_,data_stage_4__4303_,data_stage_4__4302_,
  data_stage_4__4301_,data_stage_4__4300_,data_stage_4__4299_,data_stage_4__4298_,
  data_stage_4__4297_,data_stage_4__4296_,data_stage_4__4295_,data_stage_4__4294_,
  data_stage_4__4293_,data_stage_4__4292_,data_stage_4__4291_,data_stage_4__4290_,
  data_stage_4__4289_,data_stage_4__4288_,data_stage_4__4287_,data_stage_4__4286_,
  data_stage_4__4285_,data_stage_4__4284_,data_stage_4__4283_,data_stage_4__4282_,
  data_stage_4__4281_,data_stage_4__4280_,data_stage_4__4279_,data_stage_4__4278_,
  data_stage_4__4277_,data_stage_4__4276_,data_stage_4__4275_,data_stage_4__4274_,
  data_stage_4__4273_,data_stage_4__4272_,data_stage_4__4271_,data_stage_4__4270_,
  data_stage_4__4269_,data_stage_4__4268_,data_stage_4__4267_,data_stage_4__4266_,
  data_stage_4__4265_,data_stage_4__4264_,data_stage_4__4263_,data_stage_4__4262_,
  data_stage_4__4261_,data_stage_4__4260_,data_stage_4__4259_,data_stage_4__4258_,
  data_stage_4__4257_,data_stage_4__4256_,data_stage_4__4255_,data_stage_4__4254_,
  data_stage_4__4253_,data_stage_4__4252_,data_stage_4__4251_,data_stage_4__4250_,
  data_stage_4__4249_,data_stage_4__4248_,data_stage_4__4247_,data_stage_4__4246_,
  data_stage_4__4245_,data_stage_4__4244_,data_stage_4__4243_,data_stage_4__4242_,
  data_stage_4__4241_,data_stage_4__4240_,data_stage_4__4239_,data_stage_4__4238_,
  data_stage_4__4237_,data_stage_4__4236_,data_stage_4__4235_,data_stage_4__4234_,
  data_stage_4__4233_,data_stage_4__4232_,data_stage_4__4231_,data_stage_4__4230_,
  data_stage_4__4229_,data_stage_4__4228_,data_stage_4__4227_,data_stage_4__4226_,
  data_stage_4__4225_,data_stage_4__4224_,data_stage_4__4223_,data_stage_4__4222_,
  data_stage_4__4221_,data_stage_4__4220_,data_stage_4__4219_,data_stage_4__4218_,
  data_stage_4__4217_,data_stage_4__4216_,data_stage_4__4215_,data_stage_4__4214_,
  data_stage_4__4213_,data_stage_4__4212_,data_stage_4__4211_,data_stage_4__4210_,
  data_stage_4__4209_,data_stage_4__4208_,data_stage_4__4207_,data_stage_4__4206_,
  data_stage_4__4205_,data_stage_4__4204_,data_stage_4__4203_,data_stage_4__4202_,
  data_stage_4__4201_,data_stage_4__4200_,data_stage_4__4199_,data_stage_4__4198_,
  data_stage_4__4197_,data_stage_4__4196_,data_stage_4__4195_,data_stage_4__4194_,
  data_stage_4__4193_,data_stage_4__4192_,data_stage_4__4191_,data_stage_4__4190_,
  data_stage_4__4189_,data_stage_4__4188_,data_stage_4__4187_,data_stage_4__4186_,
  data_stage_4__4185_,data_stage_4__4184_,data_stage_4__4183_,data_stage_4__4182_,
  data_stage_4__4181_,data_stage_4__4180_,data_stage_4__4179_,data_stage_4__4178_,
  data_stage_4__4177_,data_stage_4__4176_,data_stage_4__4175_,data_stage_4__4174_,
  data_stage_4__4173_,data_stage_4__4172_,data_stage_4__4171_,data_stage_4__4170_,
  data_stage_4__4169_,data_stage_4__4168_,data_stage_4__4167_,data_stage_4__4166_,
  data_stage_4__4165_,data_stage_4__4164_,data_stage_4__4163_,data_stage_4__4162_,
  data_stage_4__4161_,data_stage_4__4160_,data_stage_4__4159_,data_stage_4__4158_,
  data_stage_4__4157_,data_stage_4__4156_,data_stage_4__4155_,data_stage_4__4154_,
  data_stage_4__4153_,data_stage_4__4152_,data_stage_4__4151_,data_stage_4__4150_,
  data_stage_4__4149_,data_stage_4__4148_,data_stage_4__4147_,data_stage_4__4146_,
  data_stage_4__4145_,data_stage_4__4144_,data_stage_4__4143_,data_stage_4__4142_,
  data_stage_4__4141_,data_stage_4__4140_,data_stage_4__4139_,data_stage_4__4138_,
  data_stage_4__4137_,data_stage_4__4136_,data_stage_4__4135_,data_stage_4__4134_,
  data_stage_4__4133_,data_stage_4__4132_,data_stage_4__4131_,data_stage_4__4130_,
  data_stage_4__4129_,data_stage_4__4128_,data_stage_4__4127_,data_stage_4__4126_,
  data_stage_4__4125_,data_stage_4__4124_,data_stage_4__4123_,data_stage_4__4122_,
  data_stage_4__4121_,data_stage_4__4120_,data_stage_4__4119_,data_stage_4__4118_,
  data_stage_4__4117_,data_stage_4__4116_,data_stage_4__4115_,data_stage_4__4114_,
  data_stage_4__4113_,data_stage_4__4112_,data_stage_4__4111_,data_stage_4__4110_,
  data_stage_4__4109_,data_stage_4__4108_,data_stage_4__4107_,data_stage_4__4106_,
  data_stage_4__4105_,data_stage_4__4104_,data_stage_4__4103_,data_stage_4__4102_,
  data_stage_4__4101_,data_stage_4__4100_,data_stage_4__4099_,data_stage_4__4098_,
  data_stage_4__4097_,data_stage_4__4096_,data_stage_4__4095_,data_stage_4__4094_,
  data_stage_4__4093_,data_stage_4__4092_,data_stage_4__4091_,data_stage_4__4090_,
  data_stage_4__4089_,data_stage_4__4088_,data_stage_4__4087_,data_stage_4__4086_,
  data_stage_4__4085_,data_stage_4__4084_,data_stage_4__4083_,data_stage_4__4082_,
  data_stage_4__4081_,data_stage_4__4080_,data_stage_4__4079_,data_stage_4__4078_,
  data_stage_4__4077_,data_stage_4__4076_,data_stage_4__4075_,data_stage_4__4074_,
  data_stage_4__4073_,data_stage_4__4072_,data_stage_4__4071_,data_stage_4__4070_,
  data_stage_4__4069_,data_stage_4__4068_,data_stage_4__4067_,data_stage_4__4066_,
  data_stage_4__4065_,data_stage_4__4064_,data_stage_4__4063_,data_stage_4__4062_,
  data_stage_4__4061_,data_stage_4__4060_,data_stage_4__4059_,data_stage_4__4058_,
  data_stage_4__4057_,data_stage_4__4056_,data_stage_4__4055_,data_stage_4__4054_,
  data_stage_4__4053_,data_stage_4__4052_,data_stage_4__4051_,data_stage_4__4050_,
  data_stage_4__4049_,data_stage_4__4048_,data_stage_4__4047_,data_stage_4__4046_,
  data_stage_4__4045_,data_stage_4__4044_,data_stage_4__4043_,data_stage_4__4042_,
  data_stage_4__4041_,data_stage_4__4040_,data_stage_4__4039_,data_stage_4__4038_,
  data_stage_4__4037_,data_stage_4__4036_,data_stage_4__4035_,data_stage_4__4034_,
  data_stage_4__4033_,data_stage_4__4032_,data_stage_4__4031_,data_stage_4__4030_,
  data_stage_4__4029_,data_stage_4__4028_,data_stage_4__4027_,data_stage_4__4026_,
  data_stage_4__4025_,data_stage_4__4024_,data_stage_4__4023_,data_stage_4__4022_,
  data_stage_4__4021_,data_stage_4__4020_,data_stage_4__4019_,data_stage_4__4018_,
  data_stage_4__4017_,data_stage_4__4016_,data_stage_4__4015_,data_stage_4__4014_,
  data_stage_4__4013_,data_stage_4__4012_,data_stage_4__4011_,data_stage_4__4010_,
  data_stage_4__4009_,data_stage_4__4008_,data_stage_4__4007_,data_stage_4__4006_,
  data_stage_4__4005_,data_stage_4__4004_,data_stage_4__4003_,data_stage_4__4002_,
  data_stage_4__4001_,data_stage_4__4000_,data_stage_4__3999_,data_stage_4__3998_,
  data_stage_4__3997_,data_stage_4__3996_,data_stage_4__3995_,data_stage_4__3994_,
  data_stage_4__3993_,data_stage_4__3992_,data_stage_4__3991_,data_stage_4__3990_,
  data_stage_4__3989_,data_stage_4__3988_,data_stage_4__3987_,data_stage_4__3986_,
  data_stage_4__3985_,data_stage_4__3984_,data_stage_4__3983_,data_stage_4__3982_,
  data_stage_4__3981_,data_stage_4__3980_,data_stage_4__3979_,data_stage_4__3978_,
  data_stage_4__3977_,data_stage_4__3976_,data_stage_4__3975_,data_stage_4__3974_,
  data_stage_4__3973_,data_stage_4__3972_,data_stage_4__3971_,data_stage_4__3970_,
  data_stage_4__3969_,data_stage_4__3968_,data_stage_4__3967_,data_stage_4__3966_,
  data_stage_4__3965_,data_stage_4__3964_,data_stage_4__3963_,data_stage_4__3962_,
  data_stage_4__3961_,data_stage_4__3960_,data_stage_4__3959_,data_stage_4__3958_,
  data_stage_4__3957_,data_stage_4__3956_,data_stage_4__3955_,data_stage_4__3954_,
  data_stage_4__3953_,data_stage_4__3952_,data_stage_4__3951_,data_stage_4__3950_,
  data_stage_4__3949_,data_stage_4__3948_,data_stage_4__3947_,data_stage_4__3946_,
  data_stage_4__3945_,data_stage_4__3944_,data_stage_4__3943_,data_stage_4__3942_,
  data_stage_4__3941_,data_stage_4__3940_,data_stage_4__3939_,data_stage_4__3938_,
  data_stage_4__3937_,data_stage_4__3936_,data_stage_4__3935_,data_stage_4__3934_,
  data_stage_4__3933_,data_stage_4__3932_,data_stage_4__3931_,data_stage_4__3930_,
  data_stage_4__3929_,data_stage_4__3928_,data_stage_4__3927_,data_stage_4__3926_,
  data_stage_4__3925_,data_stage_4__3924_,data_stage_4__3923_,data_stage_4__3922_,
  data_stage_4__3921_,data_stage_4__3920_,data_stage_4__3919_,data_stage_4__3918_,
  data_stage_4__3917_,data_stage_4__3916_,data_stage_4__3915_,data_stage_4__3914_,
  data_stage_4__3913_,data_stage_4__3912_,data_stage_4__3911_,data_stage_4__3910_,
  data_stage_4__3909_,data_stage_4__3908_,data_stage_4__3907_,data_stage_4__3906_,
  data_stage_4__3905_,data_stage_4__3904_,data_stage_4__3903_,data_stage_4__3902_,
  data_stage_4__3901_,data_stage_4__3900_,data_stage_4__3899_,data_stage_4__3898_,
  data_stage_4__3897_,data_stage_4__3896_,data_stage_4__3895_,data_stage_4__3894_,
  data_stage_4__3893_,data_stage_4__3892_,data_stage_4__3891_,data_stage_4__3890_,
  data_stage_4__3889_,data_stage_4__3888_,data_stage_4__3887_,data_stage_4__3886_,
  data_stage_4__3885_,data_stage_4__3884_,data_stage_4__3883_,data_stage_4__3882_,
  data_stage_4__3881_,data_stage_4__3880_,data_stage_4__3879_,data_stage_4__3878_,
  data_stage_4__3877_,data_stage_4__3876_,data_stage_4__3875_,data_stage_4__3874_,
  data_stage_4__3873_,data_stage_4__3872_,data_stage_4__3871_,data_stage_4__3870_,
  data_stage_4__3869_,data_stage_4__3868_,data_stage_4__3867_,data_stage_4__3866_,
  data_stage_4__3865_,data_stage_4__3864_,data_stage_4__3863_,data_stage_4__3862_,
  data_stage_4__3861_,data_stage_4__3860_,data_stage_4__3859_,data_stage_4__3858_,
  data_stage_4__3857_,data_stage_4__3856_,data_stage_4__3855_,data_stage_4__3854_,
  data_stage_4__3853_,data_stage_4__3852_,data_stage_4__3851_,data_stage_4__3850_,
  data_stage_4__3849_,data_stage_4__3848_,data_stage_4__3847_,data_stage_4__3846_,
  data_stage_4__3845_,data_stage_4__3844_,data_stage_4__3843_,data_stage_4__3842_,
  data_stage_4__3841_,data_stage_4__3840_,data_stage_4__3839_,data_stage_4__3838_,
  data_stage_4__3837_,data_stage_4__3836_,data_stage_4__3835_,data_stage_4__3834_,
  data_stage_4__3833_,data_stage_4__3832_,data_stage_4__3831_,data_stage_4__3830_,
  data_stage_4__3829_,data_stage_4__3828_,data_stage_4__3827_,data_stage_4__3826_,
  data_stage_4__3825_,data_stage_4__3824_,data_stage_4__3823_,data_stage_4__3822_,
  data_stage_4__3821_,data_stage_4__3820_,data_stage_4__3819_,data_stage_4__3818_,
  data_stage_4__3817_,data_stage_4__3816_,data_stage_4__3815_,data_stage_4__3814_,
  data_stage_4__3813_,data_stage_4__3812_,data_stage_4__3811_,data_stage_4__3810_,
  data_stage_4__3809_,data_stage_4__3808_,data_stage_4__3807_,data_stage_4__3806_,
  data_stage_4__3805_,data_stage_4__3804_,data_stage_4__3803_,data_stage_4__3802_,
  data_stage_4__3801_,data_stage_4__3800_,data_stage_4__3799_,data_stage_4__3798_,
  data_stage_4__3797_,data_stage_4__3796_,data_stage_4__3795_,data_stage_4__3794_,
  data_stage_4__3793_,data_stage_4__3792_,data_stage_4__3791_,data_stage_4__3790_,
  data_stage_4__3789_,data_stage_4__3788_,data_stage_4__3787_,data_stage_4__3786_,
  data_stage_4__3785_,data_stage_4__3784_,data_stage_4__3783_,data_stage_4__3782_,
  data_stage_4__3781_,data_stage_4__3780_,data_stage_4__3779_,data_stage_4__3778_,
  data_stage_4__3777_,data_stage_4__3776_,data_stage_4__3775_,data_stage_4__3774_,
  data_stage_4__3773_,data_stage_4__3772_,data_stage_4__3771_,data_stage_4__3770_,
  data_stage_4__3769_,data_stage_4__3768_,data_stage_4__3767_,data_stage_4__3766_,
  data_stage_4__3765_,data_stage_4__3764_,data_stage_4__3763_,data_stage_4__3762_,
  data_stage_4__3761_,data_stage_4__3760_,data_stage_4__3759_,data_stage_4__3758_,
  data_stage_4__3757_,data_stage_4__3756_,data_stage_4__3755_,data_stage_4__3754_,
  data_stage_4__3753_,data_stage_4__3752_,data_stage_4__3751_,data_stage_4__3750_,
  data_stage_4__3749_,data_stage_4__3748_,data_stage_4__3747_,data_stage_4__3746_,
  data_stage_4__3745_,data_stage_4__3744_,data_stage_4__3743_,data_stage_4__3742_,
  data_stage_4__3741_,data_stage_4__3740_,data_stage_4__3739_,data_stage_4__3738_,
  data_stage_4__3737_,data_stage_4__3736_,data_stage_4__3735_,data_stage_4__3734_,
  data_stage_4__3733_,data_stage_4__3732_,data_stage_4__3731_,data_stage_4__3730_,
  data_stage_4__3729_,data_stage_4__3728_,data_stage_4__3727_,data_stage_4__3726_,
  data_stage_4__3725_,data_stage_4__3724_,data_stage_4__3723_,data_stage_4__3722_,
  data_stage_4__3721_,data_stage_4__3720_,data_stage_4__3719_,data_stage_4__3718_,
  data_stage_4__3717_,data_stage_4__3716_,data_stage_4__3715_,data_stage_4__3714_,
  data_stage_4__3713_,data_stage_4__3712_,data_stage_4__3711_,data_stage_4__3710_,
  data_stage_4__3709_,data_stage_4__3708_,data_stage_4__3707_,data_stage_4__3706_,
  data_stage_4__3705_,data_stage_4__3704_,data_stage_4__3703_,data_stage_4__3702_,
  data_stage_4__3701_,data_stage_4__3700_,data_stage_4__3699_,data_stage_4__3698_,
  data_stage_4__3697_,data_stage_4__3696_,data_stage_4__3695_,data_stage_4__3694_,
  data_stage_4__3693_,data_stage_4__3692_,data_stage_4__3691_,data_stage_4__3690_,
  data_stage_4__3689_,data_stage_4__3688_,data_stage_4__3687_,data_stage_4__3686_,
  data_stage_4__3685_,data_stage_4__3684_,data_stage_4__3683_,data_stage_4__3682_,
  data_stage_4__3681_,data_stage_4__3680_,data_stage_4__3679_,data_stage_4__3678_,
  data_stage_4__3677_,data_stage_4__3676_,data_stage_4__3675_,data_stage_4__3674_,
  data_stage_4__3673_,data_stage_4__3672_,data_stage_4__3671_,data_stage_4__3670_,
  data_stage_4__3669_,data_stage_4__3668_,data_stage_4__3667_,data_stage_4__3666_,
  data_stage_4__3665_,data_stage_4__3664_,data_stage_4__3663_,data_stage_4__3662_,
  data_stage_4__3661_,data_stage_4__3660_,data_stage_4__3659_,data_stage_4__3658_,
  data_stage_4__3657_,data_stage_4__3656_,data_stage_4__3655_,data_stage_4__3654_,
  data_stage_4__3653_,data_stage_4__3652_,data_stage_4__3651_,data_stage_4__3650_,
  data_stage_4__3649_,data_stage_4__3648_,data_stage_4__3647_,data_stage_4__3646_,
  data_stage_4__3645_,data_stage_4__3644_,data_stage_4__3643_,data_stage_4__3642_,
  data_stage_4__3641_,data_stage_4__3640_,data_stage_4__3639_,data_stage_4__3638_,
  data_stage_4__3637_,data_stage_4__3636_,data_stage_4__3635_,data_stage_4__3634_,
  data_stage_4__3633_,data_stage_4__3632_,data_stage_4__3631_,data_stage_4__3630_,
  data_stage_4__3629_,data_stage_4__3628_,data_stage_4__3627_,data_stage_4__3626_,
  data_stage_4__3625_,data_stage_4__3624_,data_stage_4__3623_,data_stage_4__3622_,
  data_stage_4__3621_,data_stage_4__3620_,data_stage_4__3619_,data_stage_4__3618_,
  data_stage_4__3617_,data_stage_4__3616_,data_stage_4__3615_,data_stage_4__3614_,
  data_stage_4__3613_,data_stage_4__3612_,data_stage_4__3611_,data_stage_4__3610_,
  data_stage_4__3609_,data_stage_4__3608_,data_stage_4__3607_,data_stage_4__3606_,
  data_stage_4__3605_,data_stage_4__3604_,data_stage_4__3603_,data_stage_4__3602_,
  data_stage_4__3601_,data_stage_4__3600_,data_stage_4__3599_,data_stage_4__3598_,
  data_stage_4__3597_,data_stage_4__3596_,data_stage_4__3595_,data_stage_4__3594_,
  data_stage_4__3593_,data_stage_4__3592_,data_stage_4__3591_,data_stage_4__3590_,
  data_stage_4__3589_,data_stage_4__3588_,data_stage_4__3587_,data_stage_4__3586_,
  data_stage_4__3585_,data_stage_4__3584_,data_stage_4__3583_,data_stage_4__3582_,
  data_stage_4__3581_,data_stage_4__3580_,data_stage_4__3579_,data_stage_4__3578_,
  data_stage_4__3577_,data_stage_4__3576_,data_stage_4__3575_,data_stage_4__3574_,
  data_stage_4__3573_,data_stage_4__3572_,data_stage_4__3571_,data_stage_4__3570_,
  data_stage_4__3569_,data_stage_4__3568_,data_stage_4__3567_,data_stage_4__3566_,
  data_stage_4__3565_,data_stage_4__3564_,data_stage_4__3563_,data_stage_4__3562_,
  data_stage_4__3561_,data_stage_4__3560_,data_stage_4__3559_,data_stage_4__3558_,
  data_stage_4__3557_,data_stage_4__3556_,data_stage_4__3555_,data_stage_4__3554_,
  data_stage_4__3553_,data_stage_4__3552_,data_stage_4__3551_,data_stage_4__3550_,
  data_stage_4__3549_,data_stage_4__3548_,data_stage_4__3547_,data_stage_4__3546_,
  data_stage_4__3545_,data_stage_4__3544_,data_stage_4__3543_,data_stage_4__3542_,
  data_stage_4__3541_,data_stage_4__3540_,data_stage_4__3539_,data_stage_4__3538_,
  data_stage_4__3537_,data_stage_4__3536_,data_stage_4__3535_,data_stage_4__3534_,
  data_stage_4__3533_,data_stage_4__3532_,data_stage_4__3531_,data_stage_4__3530_,
  data_stage_4__3529_,data_stage_4__3528_,data_stage_4__3527_,data_stage_4__3526_,
  data_stage_4__3525_,data_stage_4__3524_,data_stage_4__3523_,data_stage_4__3522_,
  data_stage_4__3521_,data_stage_4__3520_,data_stage_4__3519_,data_stage_4__3518_,
  data_stage_4__3517_,data_stage_4__3516_,data_stage_4__3515_,data_stage_4__3514_,
  data_stage_4__3513_,data_stage_4__3512_,data_stage_4__3511_,data_stage_4__3510_,
  data_stage_4__3509_,data_stage_4__3508_,data_stage_4__3507_,data_stage_4__3506_,
  data_stage_4__3505_,data_stage_4__3504_,data_stage_4__3503_,data_stage_4__3502_,
  data_stage_4__3501_,data_stage_4__3500_,data_stage_4__3499_,data_stage_4__3498_,
  data_stage_4__3497_,data_stage_4__3496_,data_stage_4__3495_,data_stage_4__3494_,
  data_stage_4__3493_,data_stage_4__3492_,data_stage_4__3491_,data_stage_4__3490_,
  data_stage_4__3489_,data_stage_4__3488_,data_stage_4__3487_,data_stage_4__3486_,
  data_stage_4__3485_,data_stage_4__3484_,data_stage_4__3483_,data_stage_4__3482_,
  data_stage_4__3481_,data_stage_4__3480_,data_stage_4__3479_,data_stage_4__3478_,
  data_stage_4__3477_,data_stage_4__3476_,data_stage_4__3475_,data_stage_4__3474_,
  data_stage_4__3473_,data_stage_4__3472_,data_stage_4__3471_,data_stage_4__3470_,
  data_stage_4__3469_,data_stage_4__3468_,data_stage_4__3467_,data_stage_4__3466_,
  data_stage_4__3465_,data_stage_4__3464_,data_stage_4__3463_,data_stage_4__3462_,
  data_stage_4__3461_,data_stage_4__3460_,data_stage_4__3459_,data_stage_4__3458_,
  data_stage_4__3457_,data_stage_4__3456_,data_stage_4__3455_,data_stage_4__3454_,
  data_stage_4__3453_,data_stage_4__3452_,data_stage_4__3451_,data_stage_4__3450_,
  data_stage_4__3449_,data_stage_4__3448_,data_stage_4__3447_,data_stage_4__3446_,
  data_stage_4__3445_,data_stage_4__3444_,data_stage_4__3443_,data_stage_4__3442_,
  data_stage_4__3441_,data_stage_4__3440_,data_stage_4__3439_,data_stage_4__3438_,
  data_stage_4__3437_,data_stage_4__3436_,data_stage_4__3435_,data_stage_4__3434_,
  data_stage_4__3433_,data_stage_4__3432_,data_stage_4__3431_,data_stage_4__3430_,
  data_stage_4__3429_,data_stage_4__3428_,data_stage_4__3427_,data_stage_4__3426_,
  data_stage_4__3425_,data_stage_4__3424_,data_stage_4__3423_,data_stage_4__3422_,
  data_stage_4__3421_,data_stage_4__3420_,data_stage_4__3419_,data_stage_4__3418_,
  data_stage_4__3417_,data_stage_4__3416_,data_stage_4__3415_,data_stage_4__3414_,
  data_stage_4__3413_,data_stage_4__3412_,data_stage_4__3411_,data_stage_4__3410_,
  data_stage_4__3409_,data_stage_4__3408_,data_stage_4__3407_,data_stage_4__3406_,
  data_stage_4__3405_,data_stage_4__3404_,data_stage_4__3403_,data_stage_4__3402_,
  data_stage_4__3401_,data_stage_4__3400_,data_stage_4__3399_,data_stage_4__3398_,
  data_stage_4__3397_,data_stage_4__3396_,data_stage_4__3395_,data_stage_4__3394_,
  data_stage_4__3393_,data_stage_4__3392_,data_stage_4__3391_,data_stage_4__3390_,
  data_stage_4__3389_,data_stage_4__3388_,data_stage_4__3387_,data_stage_4__3386_,
  data_stage_4__3385_,data_stage_4__3384_,data_stage_4__3383_,data_stage_4__3382_,
  data_stage_4__3381_,data_stage_4__3380_,data_stage_4__3379_,data_stage_4__3378_,
  data_stage_4__3377_,data_stage_4__3376_,data_stage_4__3375_,data_stage_4__3374_,
  data_stage_4__3373_,data_stage_4__3372_,data_stage_4__3371_,data_stage_4__3370_,
  data_stage_4__3369_,data_stage_4__3368_,data_stage_4__3367_,data_stage_4__3366_,
  data_stage_4__3365_,data_stage_4__3364_,data_stage_4__3363_,data_stage_4__3362_,
  data_stage_4__3361_,data_stage_4__3360_,data_stage_4__3359_,data_stage_4__3358_,
  data_stage_4__3357_,data_stage_4__3356_,data_stage_4__3355_,data_stage_4__3354_,
  data_stage_4__3353_,data_stage_4__3352_,data_stage_4__3351_,data_stage_4__3350_,
  data_stage_4__3349_,data_stage_4__3348_,data_stage_4__3347_,data_stage_4__3346_,
  data_stage_4__3345_,data_stage_4__3344_,data_stage_4__3343_,data_stage_4__3342_,
  data_stage_4__3341_,data_stage_4__3340_,data_stage_4__3339_,data_stage_4__3338_,
  data_stage_4__3337_,data_stage_4__3336_,data_stage_4__3335_,data_stage_4__3334_,
  data_stage_4__3333_,data_stage_4__3332_,data_stage_4__3331_,data_stage_4__3330_,
  data_stage_4__3329_,data_stage_4__3328_,data_stage_4__3327_,data_stage_4__3326_,
  data_stage_4__3325_,data_stage_4__3324_,data_stage_4__3323_,data_stage_4__3322_,
  data_stage_4__3321_,data_stage_4__3320_,data_stage_4__3319_,data_stage_4__3318_,
  data_stage_4__3317_,data_stage_4__3316_,data_stage_4__3315_,data_stage_4__3314_,
  data_stage_4__3313_,data_stage_4__3312_,data_stage_4__3311_,data_stage_4__3310_,
  data_stage_4__3309_,data_stage_4__3308_,data_stage_4__3307_,data_stage_4__3306_,
  data_stage_4__3305_,data_stage_4__3304_,data_stage_4__3303_,data_stage_4__3302_,
  data_stage_4__3301_,data_stage_4__3300_,data_stage_4__3299_,data_stage_4__3298_,
  data_stage_4__3297_,data_stage_4__3296_,data_stage_4__3295_,data_stage_4__3294_,
  data_stage_4__3293_,data_stage_4__3292_,data_stage_4__3291_,data_stage_4__3290_,
  data_stage_4__3289_,data_stage_4__3288_,data_stage_4__3287_,data_stage_4__3286_,
  data_stage_4__3285_,data_stage_4__3284_,data_stage_4__3283_,data_stage_4__3282_,
  data_stage_4__3281_,data_stage_4__3280_,data_stage_4__3279_,data_stage_4__3278_,
  data_stage_4__3277_,data_stage_4__3276_,data_stage_4__3275_,data_stage_4__3274_,
  data_stage_4__3273_,data_stage_4__3272_,data_stage_4__3271_,data_stage_4__3270_,
  data_stage_4__3269_,data_stage_4__3268_,data_stage_4__3267_,data_stage_4__3266_,
  data_stage_4__3265_,data_stage_4__3264_,data_stage_4__3263_,data_stage_4__3262_,
  data_stage_4__3261_,data_stage_4__3260_,data_stage_4__3259_,data_stage_4__3258_,
  data_stage_4__3257_,data_stage_4__3256_,data_stage_4__3255_,data_stage_4__3254_,
  data_stage_4__3253_,data_stage_4__3252_,data_stage_4__3251_,data_stage_4__3250_,
  data_stage_4__3249_,data_stage_4__3248_,data_stage_4__3247_,data_stage_4__3246_,
  data_stage_4__3245_,data_stage_4__3244_,data_stage_4__3243_,data_stage_4__3242_,
  data_stage_4__3241_,data_stage_4__3240_,data_stage_4__3239_,data_stage_4__3238_,
  data_stage_4__3237_,data_stage_4__3236_,data_stage_4__3235_,data_stage_4__3234_,
  data_stage_4__3233_,data_stage_4__3232_,data_stage_4__3231_,data_stage_4__3230_,
  data_stage_4__3229_,data_stage_4__3228_,data_stage_4__3227_,data_stage_4__3226_,
  data_stage_4__3225_,data_stage_4__3224_,data_stage_4__3223_,data_stage_4__3222_,
  data_stage_4__3221_,data_stage_4__3220_,data_stage_4__3219_,data_stage_4__3218_,
  data_stage_4__3217_,data_stage_4__3216_,data_stage_4__3215_,data_stage_4__3214_,
  data_stage_4__3213_,data_stage_4__3212_,data_stage_4__3211_,data_stage_4__3210_,
  data_stage_4__3209_,data_stage_4__3208_,data_stage_4__3207_,data_stage_4__3206_,
  data_stage_4__3205_,data_stage_4__3204_,data_stage_4__3203_,data_stage_4__3202_,
  data_stage_4__3201_,data_stage_4__3200_,data_stage_4__3199_,data_stage_4__3198_,
  data_stage_4__3197_,data_stage_4__3196_,data_stage_4__3195_,data_stage_4__3194_,
  data_stage_4__3193_,data_stage_4__3192_,data_stage_4__3191_,data_stage_4__3190_,
  data_stage_4__3189_,data_stage_4__3188_,data_stage_4__3187_,data_stage_4__3186_,
  data_stage_4__3185_,data_stage_4__3184_,data_stage_4__3183_,data_stage_4__3182_,
  data_stage_4__3181_,data_stage_4__3180_,data_stage_4__3179_,data_stage_4__3178_,
  data_stage_4__3177_,data_stage_4__3176_,data_stage_4__3175_,data_stage_4__3174_,
  data_stage_4__3173_,data_stage_4__3172_,data_stage_4__3171_,data_stage_4__3170_,
  data_stage_4__3169_,data_stage_4__3168_,data_stage_4__3167_,data_stage_4__3166_,
  data_stage_4__3165_,data_stage_4__3164_,data_stage_4__3163_,data_stage_4__3162_,
  data_stage_4__3161_,data_stage_4__3160_,data_stage_4__3159_,data_stage_4__3158_,
  data_stage_4__3157_,data_stage_4__3156_,data_stage_4__3155_,data_stage_4__3154_,
  data_stage_4__3153_,data_stage_4__3152_,data_stage_4__3151_,data_stage_4__3150_,
  data_stage_4__3149_,data_stage_4__3148_,data_stage_4__3147_,data_stage_4__3146_,
  data_stage_4__3145_,data_stage_4__3144_,data_stage_4__3143_,data_stage_4__3142_,
  data_stage_4__3141_,data_stage_4__3140_,data_stage_4__3139_,data_stage_4__3138_,
  data_stage_4__3137_,data_stage_4__3136_,data_stage_4__3135_,data_stage_4__3134_,
  data_stage_4__3133_,data_stage_4__3132_,data_stage_4__3131_,data_stage_4__3130_,
  data_stage_4__3129_,data_stage_4__3128_,data_stage_4__3127_,data_stage_4__3126_,
  data_stage_4__3125_,data_stage_4__3124_,data_stage_4__3123_,data_stage_4__3122_,
  data_stage_4__3121_,data_stage_4__3120_,data_stage_4__3119_,data_stage_4__3118_,
  data_stage_4__3117_,data_stage_4__3116_,data_stage_4__3115_,data_stage_4__3114_,
  data_stage_4__3113_,data_stage_4__3112_,data_stage_4__3111_,data_stage_4__3110_,
  data_stage_4__3109_,data_stage_4__3108_,data_stage_4__3107_,data_stage_4__3106_,
  data_stage_4__3105_,data_stage_4__3104_,data_stage_4__3103_,data_stage_4__3102_,
  data_stage_4__3101_,data_stage_4__3100_,data_stage_4__3099_,data_stage_4__3098_,
  data_stage_4__3097_,data_stage_4__3096_,data_stage_4__3095_,data_stage_4__3094_,
  data_stage_4__3093_,data_stage_4__3092_,data_stage_4__3091_,data_stage_4__3090_,
  data_stage_4__3089_,data_stage_4__3088_,data_stage_4__3087_,data_stage_4__3086_,
  data_stage_4__3085_,data_stage_4__3084_,data_stage_4__3083_,data_stage_4__3082_,
  data_stage_4__3081_,data_stage_4__3080_,data_stage_4__3079_,data_stage_4__3078_,
  data_stage_4__3077_,data_stage_4__3076_,data_stage_4__3075_,data_stage_4__3074_,
  data_stage_4__3073_,data_stage_4__3072_,data_stage_4__3071_,data_stage_4__3070_,
  data_stage_4__3069_,data_stage_4__3068_,data_stage_4__3067_,data_stage_4__3066_,
  data_stage_4__3065_,data_stage_4__3064_,data_stage_4__3063_,data_stage_4__3062_,
  data_stage_4__3061_,data_stage_4__3060_,data_stage_4__3059_,data_stage_4__3058_,
  data_stage_4__3057_,data_stage_4__3056_,data_stage_4__3055_,data_stage_4__3054_,
  data_stage_4__3053_,data_stage_4__3052_,data_stage_4__3051_,data_stage_4__3050_,
  data_stage_4__3049_,data_stage_4__3048_,data_stage_4__3047_,data_stage_4__3046_,
  data_stage_4__3045_,data_stage_4__3044_,data_stage_4__3043_,data_stage_4__3042_,
  data_stage_4__3041_,data_stage_4__3040_,data_stage_4__3039_,data_stage_4__3038_,
  data_stage_4__3037_,data_stage_4__3036_,data_stage_4__3035_,data_stage_4__3034_,
  data_stage_4__3033_,data_stage_4__3032_,data_stage_4__3031_,data_stage_4__3030_,
  data_stage_4__3029_,data_stage_4__3028_,data_stage_4__3027_,data_stage_4__3026_,
  data_stage_4__3025_,data_stage_4__3024_,data_stage_4__3023_,data_stage_4__3022_,
  data_stage_4__3021_,data_stage_4__3020_,data_stage_4__3019_,data_stage_4__3018_,
  data_stage_4__3017_,data_stage_4__3016_,data_stage_4__3015_,data_stage_4__3014_,
  data_stage_4__3013_,data_stage_4__3012_,data_stage_4__3011_,data_stage_4__3010_,
  data_stage_4__3009_,data_stage_4__3008_,data_stage_4__3007_,data_stage_4__3006_,
  data_stage_4__3005_,data_stage_4__3004_,data_stage_4__3003_,data_stage_4__3002_,
  data_stage_4__3001_,data_stage_4__3000_,data_stage_4__2999_,data_stage_4__2998_,
  data_stage_4__2997_,data_stage_4__2996_,data_stage_4__2995_,data_stage_4__2994_,
  data_stage_4__2993_,data_stage_4__2992_,data_stage_4__2991_,data_stage_4__2990_,
  data_stage_4__2989_,data_stage_4__2988_,data_stage_4__2987_,data_stage_4__2986_,
  data_stage_4__2985_,data_stage_4__2984_,data_stage_4__2983_,data_stage_4__2982_,
  data_stage_4__2981_,data_stage_4__2980_,data_stage_4__2979_,data_stage_4__2978_,
  data_stage_4__2977_,data_stage_4__2976_,data_stage_4__2975_,data_stage_4__2974_,
  data_stage_4__2973_,data_stage_4__2972_,data_stage_4__2971_,data_stage_4__2970_,
  data_stage_4__2969_,data_stage_4__2968_,data_stage_4__2967_,data_stage_4__2966_,
  data_stage_4__2965_,data_stage_4__2964_,data_stage_4__2963_,data_stage_4__2962_,
  data_stage_4__2961_,data_stage_4__2960_,data_stage_4__2959_,data_stage_4__2958_,
  data_stage_4__2957_,data_stage_4__2956_,data_stage_4__2955_,data_stage_4__2954_,
  data_stage_4__2953_,data_stage_4__2952_,data_stage_4__2951_,data_stage_4__2950_,
  data_stage_4__2949_,data_stage_4__2948_,data_stage_4__2947_,data_stage_4__2946_,
  data_stage_4__2945_,data_stage_4__2944_,data_stage_4__2943_,data_stage_4__2942_,
  data_stage_4__2941_,data_stage_4__2940_,data_stage_4__2939_,data_stage_4__2938_,
  data_stage_4__2937_,data_stage_4__2936_,data_stage_4__2935_,data_stage_4__2934_,
  data_stage_4__2933_,data_stage_4__2932_,data_stage_4__2931_,data_stage_4__2930_,
  data_stage_4__2929_,data_stage_4__2928_,data_stage_4__2927_,data_stage_4__2926_,
  data_stage_4__2925_,data_stage_4__2924_,data_stage_4__2923_,data_stage_4__2922_,
  data_stage_4__2921_,data_stage_4__2920_,data_stage_4__2919_,data_stage_4__2918_,
  data_stage_4__2917_,data_stage_4__2916_,data_stage_4__2915_,data_stage_4__2914_,
  data_stage_4__2913_,data_stage_4__2912_,data_stage_4__2911_,data_stage_4__2910_,
  data_stage_4__2909_,data_stage_4__2908_,data_stage_4__2907_,data_stage_4__2906_,
  data_stage_4__2905_,data_stage_4__2904_,data_stage_4__2903_,data_stage_4__2902_,
  data_stage_4__2901_,data_stage_4__2900_,data_stage_4__2899_,data_stage_4__2898_,
  data_stage_4__2897_,data_stage_4__2896_,data_stage_4__2895_,data_stage_4__2894_,
  data_stage_4__2893_,data_stage_4__2892_,data_stage_4__2891_,data_stage_4__2890_,
  data_stage_4__2889_,data_stage_4__2888_,data_stage_4__2887_,data_stage_4__2886_,
  data_stage_4__2885_,data_stage_4__2884_,data_stage_4__2883_,data_stage_4__2882_,
  data_stage_4__2881_,data_stage_4__2880_,data_stage_4__2879_,data_stage_4__2878_,
  data_stage_4__2877_,data_stage_4__2876_,data_stage_4__2875_,data_stage_4__2874_,
  data_stage_4__2873_,data_stage_4__2872_,data_stage_4__2871_,data_stage_4__2870_,
  data_stage_4__2869_,data_stage_4__2868_,data_stage_4__2867_,data_stage_4__2866_,
  data_stage_4__2865_,data_stage_4__2864_,data_stage_4__2863_,data_stage_4__2862_,
  data_stage_4__2861_,data_stage_4__2860_,data_stage_4__2859_,data_stage_4__2858_,
  data_stage_4__2857_,data_stage_4__2856_,data_stage_4__2855_,data_stage_4__2854_,
  data_stage_4__2853_,data_stage_4__2852_,data_stage_4__2851_,data_stage_4__2850_,
  data_stage_4__2849_,data_stage_4__2848_,data_stage_4__2847_,data_stage_4__2846_,
  data_stage_4__2845_,data_stage_4__2844_,data_stage_4__2843_,data_stage_4__2842_,
  data_stage_4__2841_,data_stage_4__2840_,data_stage_4__2839_,data_stage_4__2838_,
  data_stage_4__2837_,data_stage_4__2836_,data_stage_4__2835_,data_stage_4__2834_,
  data_stage_4__2833_,data_stage_4__2832_,data_stage_4__2831_,data_stage_4__2830_,
  data_stage_4__2829_,data_stage_4__2828_,data_stage_4__2827_,data_stage_4__2826_,
  data_stage_4__2825_,data_stage_4__2824_,data_stage_4__2823_,data_stage_4__2822_,
  data_stage_4__2821_,data_stage_4__2820_,data_stage_4__2819_,data_stage_4__2818_,
  data_stage_4__2817_,data_stage_4__2816_,data_stage_4__2815_,data_stage_4__2814_,
  data_stage_4__2813_,data_stage_4__2812_,data_stage_4__2811_,data_stage_4__2810_,
  data_stage_4__2809_,data_stage_4__2808_,data_stage_4__2807_,data_stage_4__2806_,
  data_stage_4__2805_,data_stage_4__2804_,data_stage_4__2803_,data_stage_4__2802_,
  data_stage_4__2801_,data_stage_4__2800_,data_stage_4__2799_,data_stage_4__2798_,
  data_stage_4__2797_,data_stage_4__2796_,data_stage_4__2795_,data_stage_4__2794_,
  data_stage_4__2793_,data_stage_4__2792_,data_stage_4__2791_,data_stage_4__2790_,
  data_stage_4__2789_,data_stage_4__2788_,data_stage_4__2787_,data_stage_4__2786_,
  data_stage_4__2785_,data_stage_4__2784_,data_stage_4__2783_,data_stage_4__2782_,
  data_stage_4__2781_,data_stage_4__2780_,data_stage_4__2779_,data_stage_4__2778_,
  data_stage_4__2777_,data_stage_4__2776_,data_stage_4__2775_,data_stage_4__2774_,
  data_stage_4__2773_,data_stage_4__2772_,data_stage_4__2771_,data_stage_4__2770_,
  data_stage_4__2769_,data_stage_4__2768_,data_stage_4__2767_,data_stage_4__2766_,
  data_stage_4__2765_,data_stage_4__2764_,data_stage_4__2763_,data_stage_4__2762_,
  data_stage_4__2761_,data_stage_4__2760_,data_stage_4__2759_,data_stage_4__2758_,
  data_stage_4__2757_,data_stage_4__2756_,data_stage_4__2755_,data_stage_4__2754_,
  data_stage_4__2753_,data_stage_4__2752_,data_stage_4__2751_,data_stage_4__2750_,
  data_stage_4__2749_,data_stage_4__2748_,data_stage_4__2747_,data_stage_4__2746_,
  data_stage_4__2745_,data_stage_4__2744_,data_stage_4__2743_,data_stage_4__2742_,
  data_stage_4__2741_,data_stage_4__2740_,data_stage_4__2739_,data_stage_4__2738_,
  data_stage_4__2737_,data_stage_4__2736_,data_stage_4__2735_,data_stage_4__2734_,
  data_stage_4__2733_,data_stage_4__2732_,data_stage_4__2731_,data_stage_4__2730_,
  data_stage_4__2729_,data_stage_4__2728_,data_stage_4__2727_,data_stage_4__2726_,
  data_stage_4__2725_,data_stage_4__2724_,data_stage_4__2723_,data_stage_4__2722_,
  data_stage_4__2721_,data_stage_4__2720_,data_stage_4__2719_,data_stage_4__2718_,
  data_stage_4__2717_,data_stage_4__2716_,data_stage_4__2715_,data_stage_4__2714_,
  data_stage_4__2713_,data_stage_4__2712_,data_stage_4__2711_,data_stage_4__2710_,
  data_stage_4__2709_,data_stage_4__2708_,data_stage_4__2707_,data_stage_4__2706_,
  data_stage_4__2705_,data_stage_4__2704_,data_stage_4__2703_,data_stage_4__2702_,
  data_stage_4__2701_,data_stage_4__2700_,data_stage_4__2699_,data_stage_4__2698_,
  data_stage_4__2697_,data_stage_4__2696_,data_stage_4__2695_,data_stage_4__2694_,
  data_stage_4__2693_,data_stage_4__2692_,data_stage_4__2691_,data_stage_4__2690_,
  data_stage_4__2689_,data_stage_4__2688_,data_stage_4__2687_,data_stage_4__2686_,
  data_stage_4__2685_,data_stage_4__2684_,data_stage_4__2683_,data_stage_4__2682_,
  data_stage_4__2681_,data_stage_4__2680_,data_stage_4__2679_,data_stage_4__2678_,
  data_stage_4__2677_,data_stage_4__2676_,data_stage_4__2675_,data_stage_4__2674_,
  data_stage_4__2673_,data_stage_4__2672_,data_stage_4__2671_,data_stage_4__2670_,
  data_stage_4__2669_,data_stage_4__2668_,data_stage_4__2667_,data_stage_4__2666_,
  data_stage_4__2665_,data_stage_4__2664_,data_stage_4__2663_,data_stage_4__2662_,
  data_stage_4__2661_,data_stage_4__2660_,data_stage_4__2659_,data_stage_4__2658_,
  data_stage_4__2657_,data_stage_4__2656_,data_stage_4__2655_,data_stage_4__2654_,
  data_stage_4__2653_,data_stage_4__2652_,data_stage_4__2651_,data_stage_4__2650_,
  data_stage_4__2649_,data_stage_4__2648_,data_stage_4__2647_,data_stage_4__2646_,
  data_stage_4__2645_,data_stage_4__2644_,data_stage_4__2643_,data_stage_4__2642_,
  data_stage_4__2641_,data_stage_4__2640_,data_stage_4__2639_,data_stage_4__2638_,
  data_stage_4__2637_,data_stage_4__2636_,data_stage_4__2635_,data_stage_4__2634_,
  data_stage_4__2633_,data_stage_4__2632_,data_stage_4__2631_,data_stage_4__2630_,
  data_stage_4__2629_,data_stage_4__2628_,data_stage_4__2627_,data_stage_4__2626_,
  data_stage_4__2625_,data_stage_4__2624_,data_stage_4__2623_,data_stage_4__2622_,
  data_stage_4__2621_,data_stage_4__2620_,data_stage_4__2619_,data_stage_4__2618_,
  data_stage_4__2617_,data_stage_4__2616_,data_stage_4__2615_,data_stage_4__2614_,
  data_stage_4__2613_,data_stage_4__2612_,data_stage_4__2611_,data_stage_4__2610_,
  data_stage_4__2609_,data_stage_4__2608_,data_stage_4__2607_,data_stage_4__2606_,
  data_stage_4__2605_,data_stage_4__2604_,data_stage_4__2603_,data_stage_4__2602_,
  data_stage_4__2601_,data_stage_4__2600_,data_stage_4__2599_,data_stage_4__2598_,
  data_stage_4__2597_,data_stage_4__2596_,data_stage_4__2595_,data_stage_4__2594_,
  data_stage_4__2593_,data_stage_4__2592_,data_stage_4__2591_,data_stage_4__2590_,
  data_stage_4__2589_,data_stage_4__2588_,data_stage_4__2587_,data_stage_4__2586_,
  data_stage_4__2585_,data_stage_4__2584_,data_stage_4__2583_,data_stage_4__2582_,
  data_stage_4__2581_,data_stage_4__2580_,data_stage_4__2579_,data_stage_4__2578_,
  data_stage_4__2577_,data_stage_4__2576_,data_stage_4__2575_,data_stage_4__2574_,
  data_stage_4__2573_,data_stage_4__2572_,data_stage_4__2571_,data_stage_4__2570_,
  data_stage_4__2569_,data_stage_4__2568_,data_stage_4__2567_,data_stage_4__2566_,
  data_stage_4__2565_,data_stage_4__2564_,data_stage_4__2563_,data_stage_4__2562_,
  data_stage_4__2561_,data_stage_4__2560_,data_stage_4__2559_,data_stage_4__2558_,
  data_stage_4__2557_,data_stage_4__2556_,data_stage_4__2555_,data_stage_4__2554_,
  data_stage_4__2553_,data_stage_4__2552_,data_stage_4__2551_,data_stage_4__2550_,
  data_stage_4__2549_,data_stage_4__2548_,data_stage_4__2547_,data_stage_4__2546_,
  data_stage_4__2545_,data_stage_4__2544_,data_stage_4__2543_,data_stage_4__2542_,
  data_stage_4__2541_,data_stage_4__2540_,data_stage_4__2539_,data_stage_4__2538_,
  data_stage_4__2537_,data_stage_4__2536_,data_stage_4__2535_,data_stage_4__2534_,
  data_stage_4__2533_,data_stage_4__2532_,data_stage_4__2531_,data_stage_4__2530_,
  data_stage_4__2529_,data_stage_4__2528_,data_stage_4__2527_,data_stage_4__2526_,
  data_stage_4__2525_,data_stage_4__2524_,data_stage_4__2523_,data_stage_4__2522_,
  data_stage_4__2521_,data_stage_4__2520_,data_stage_4__2519_,data_stage_4__2518_,
  data_stage_4__2517_,data_stage_4__2516_,data_stage_4__2515_,data_stage_4__2514_,
  data_stage_4__2513_,data_stage_4__2512_,data_stage_4__2511_,data_stage_4__2510_,
  data_stage_4__2509_,data_stage_4__2508_,data_stage_4__2507_,data_stage_4__2506_,
  data_stage_4__2505_,data_stage_4__2504_,data_stage_4__2503_,data_stage_4__2502_,
  data_stage_4__2501_,data_stage_4__2500_,data_stage_4__2499_,data_stage_4__2498_,
  data_stage_4__2497_,data_stage_4__2496_,data_stage_4__2495_,data_stage_4__2494_,
  data_stage_4__2493_,data_stage_4__2492_,data_stage_4__2491_,data_stage_4__2490_,
  data_stage_4__2489_,data_stage_4__2488_,data_stage_4__2487_,data_stage_4__2486_,
  data_stage_4__2485_,data_stage_4__2484_,data_stage_4__2483_,data_stage_4__2482_,
  data_stage_4__2481_,data_stage_4__2480_,data_stage_4__2479_,data_stage_4__2478_,
  data_stage_4__2477_,data_stage_4__2476_,data_stage_4__2475_,data_stage_4__2474_,
  data_stage_4__2473_,data_stage_4__2472_,data_stage_4__2471_,data_stage_4__2470_,
  data_stage_4__2469_,data_stage_4__2468_,data_stage_4__2467_,data_stage_4__2466_,
  data_stage_4__2465_,data_stage_4__2464_,data_stage_4__2463_,data_stage_4__2462_,
  data_stage_4__2461_,data_stage_4__2460_,data_stage_4__2459_,data_stage_4__2458_,
  data_stage_4__2457_,data_stage_4__2456_,data_stage_4__2455_,data_stage_4__2454_,
  data_stage_4__2453_,data_stage_4__2452_,data_stage_4__2451_,data_stage_4__2450_,
  data_stage_4__2449_,data_stage_4__2448_,data_stage_4__2447_,data_stage_4__2446_,
  data_stage_4__2445_,data_stage_4__2444_,data_stage_4__2443_,data_stage_4__2442_,
  data_stage_4__2441_,data_stage_4__2440_,data_stage_4__2439_,data_stage_4__2438_,
  data_stage_4__2437_,data_stage_4__2436_,data_stage_4__2435_,data_stage_4__2434_,
  data_stage_4__2433_,data_stage_4__2432_,data_stage_4__2431_,data_stage_4__2430_,
  data_stage_4__2429_,data_stage_4__2428_,data_stage_4__2427_,data_stage_4__2426_,
  data_stage_4__2425_,data_stage_4__2424_,data_stage_4__2423_,data_stage_4__2422_,
  data_stage_4__2421_,data_stage_4__2420_,data_stage_4__2419_,data_stage_4__2418_,
  data_stage_4__2417_,data_stage_4__2416_,data_stage_4__2415_,data_stage_4__2414_,
  data_stage_4__2413_,data_stage_4__2412_,data_stage_4__2411_,data_stage_4__2410_,
  data_stage_4__2409_,data_stage_4__2408_,data_stage_4__2407_,data_stage_4__2406_,
  data_stage_4__2405_,data_stage_4__2404_,data_stage_4__2403_,data_stage_4__2402_,
  data_stage_4__2401_,data_stage_4__2400_,data_stage_4__2399_,data_stage_4__2398_,
  data_stage_4__2397_,data_stage_4__2396_,data_stage_4__2395_,data_stage_4__2394_,
  data_stage_4__2393_,data_stage_4__2392_,data_stage_4__2391_,data_stage_4__2390_,
  data_stage_4__2389_,data_stage_4__2388_,data_stage_4__2387_,data_stage_4__2386_,
  data_stage_4__2385_,data_stage_4__2384_,data_stage_4__2383_,data_stage_4__2382_,
  data_stage_4__2381_,data_stage_4__2380_,data_stage_4__2379_,data_stage_4__2378_,
  data_stage_4__2377_,data_stage_4__2376_,data_stage_4__2375_,data_stage_4__2374_,
  data_stage_4__2373_,data_stage_4__2372_,data_stage_4__2371_,data_stage_4__2370_,
  data_stage_4__2369_,data_stage_4__2368_,data_stage_4__2367_,data_stage_4__2366_,
  data_stage_4__2365_,data_stage_4__2364_,data_stage_4__2363_,data_stage_4__2362_,
  data_stage_4__2361_,data_stage_4__2360_,data_stage_4__2359_,data_stage_4__2358_,
  data_stage_4__2357_,data_stage_4__2356_,data_stage_4__2355_,data_stage_4__2354_,
  data_stage_4__2353_,data_stage_4__2352_,data_stage_4__2351_,data_stage_4__2350_,
  data_stage_4__2349_,data_stage_4__2348_,data_stage_4__2347_,data_stage_4__2346_,
  data_stage_4__2345_,data_stage_4__2344_,data_stage_4__2343_,data_stage_4__2342_,
  data_stage_4__2341_,data_stage_4__2340_,data_stage_4__2339_,data_stage_4__2338_,
  data_stage_4__2337_,data_stage_4__2336_,data_stage_4__2335_,data_stage_4__2334_,
  data_stage_4__2333_,data_stage_4__2332_,data_stage_4__2331_,data_stage_4__2330_,
  data_stage_4__2329_,data_stage_4__2328_,data_stage_4__2327_,data_stage_4__2326_,
  data_stage_4__2325_,data_stage_4__2324_,data_stage_4__2323_,data_stage_4__2322_,
  data_stage_4__2321_,data_stage_4__2320_,data_stage_4__2319_,data_stage_4__2318_,
  data_stage_4__2317_,data_stage_4__2316_,data_stage_4__2315_,data_stage_4__2314_,
  data_stage_4__2313_,data_stage_4__2312_,data_stage_4__2311_,data_stage_4__2310_,
  data_stage_4__2309_,data_stage_4__2308_,data_stage_4__2307_,data_stage_4__2306_,
  data_stage_4__2305_,data_stage_4__2304_,data_stage_4__2303_,data_stage_4__2302_,
  data_stage_4__2301_,data_stage_4__2300_,data_stage_4__2299_,data_stage_4__2298_,
  data_stage_4__2297_,data_stage_4__2296_,data_stage_4__2295_,data_stage_4__2294_,
  data_stage_4__2293_,data_stage_4__2292_,data_stage_4__2291_,data_stage_4__2290_,
  data_stage_4__2289_,data_stage_4__2288_,data_stage_4__2287_,data_stage_4__2286_,
  data_stage_4__2285_,data_stage_4__2284_,data_stage_4__2283_,data_stage_4__2282_,
  data_stage_4__2281_,data_stage_4__2280_,data_stage_4__2279_,data_stage_4__2278_,
  data_stage_4__2277_,data_stage_4__2276_,data_stage_4__2275_,data_stage_4__2274_,
  data_stage_4__2273_,data_stage_4__2272_,data_stage_4__2271_,data_stage_4__2270_,
  data_stage_4__2269_,data_stage_4__2268_,data_stage_4__2267_,data_stage_4__2266_,
  data_stage_4__2265_,data_stage_4__2264_,data_stage_4__2263_,data_stage_4__2262_,
  data_stage_4__2261_,data_stage_4__2260_,data_stage_4__2259_,data_stage_4__2258_,
  data_stage_4__2257_,data_stage_4__2256_,data_stage_4__2255_,data_stage_4__2254_,
  data_stage_4__2253_,data_stage_4__2252_,data_stage_4__2251_,data_stage_4__2250_,
  data_stage_4__2249_,data_stage_4__2248_,data_stage_4__2247_,data_stage_4__2246_,
  data_stage_4__2245_,data_stage_4__2244_,data_stage_4__2243_,data_stage_4__2242_,
  data_stage_4__2241_,data_stage_4__2240_,data_stage_4__2239_,data_stage_4__2238_,
  data_stage_4__2237_,data_stage_4__2236_,data_stage_4__2235_,data_stage_4__2234_,
  data_stage_4__2233_,data_stage_4__2232_,data_stage_4__2231_,data_stage_4__2230_,
  data_stage_4__2229_,data_stage_4__2228_,data_stage_4__2227_,data_stage_4__2226_,
  data_stage_4__2225_,data_stage_4__2224_,data_stage_4__2223_,data_stage_4__2222_,
  data_stage_4__2221_,data_stage_4__2220_,data_stage_4__2219_,data_stage_4__2218_,
  data_stage_4__2217_,data_stage_4__2216_,data_stage_4__2215_,data_stage_4__2214_,
  data_stage_4__2213_,data_stage_4__2212_,data_stage_4__2211_,data_stage_4__2210_,
  data_stage_4__2209_,data_stage_4__2208_,data_stage_4__2207_,data_stage_4__2206_,
  data_stage_4__2205_,data_stage_4__2204_,data_stage_4__2203_,data_stage_4__2202_,
  data_stage_4__2201_,data_stage_4__2200_,data_stage_4__2199_,data_stage_4__2198_,
  data_stage_4__2197_,data_stage_4__2196_,data_stage_4__2195_,data_stage_4__2194_,
  data_stage_4__2193_,data_stage_4__2192_,data_stage_4__2191_,data_stage_4__2190_,
  data_stage_4__2189_,data_stage_4__2188_,data_stage_4__2187_,data_stage_4__2186_,
  data_stage_4__2185_,data_stage_4__2184_,data_stage_4__2183_,data_stage_4__2182_,
  data_stage_4__2181_,data_stage_4__2180_,data_stage_4__2179_,data_stage_4__2178_,
  data_stage_4__2177_,data_stage_4__2176_,data_stage_4__2175_,data_stage_4__2174_,
  data_stage_4__2173_,data_stage_4__2172_,data_stage_4__2171_,data_stage_4__2170_,
  data_stage_4__2169_,data_stage_4__2168_,data_stage_4__2167_,data_stage_4__2166_,
  data_stage_4__2165_,data_stage_4__2164_,data_stage_4__2163_,data_stage_4__2162_,
  data_stage_4__2161_,data_stage_4__2160_,data_stage_4__2159_,data_stage_4__2158_,
  data_stage_4__2157_,data_stage_4__2156_,data_stage_4__2155_,data_stage_4__2154_,
  data_stage_4__2153_,data_stage_4__2152_,data_stage_4__2151_,data_stage_4__2150_,
  data_stage_4__2149_,data_stage_4__2148_,data_stage_4__2147_,data_stage_4__2146_,
  data_stage_4__2145_,data_stage_4__2144_,data_stage_4__2143_,data_stage_4__2142_,
  data_stage_4__2141_,data_stage_4__2140_,data_stage_4__2139_,data_stage_4__2138_,
  data_stage_4__2137_,data_stage_4__2136_,data_stage_4__2135_,data_stage_4__2134_,
  data_stage_4__2133_,data_stage_4__2132_,data_stage_4__2131_,data_stage_4__2130_,
  data_stage_4__2129_,data_stage_4__2128_,data_stage_4__2127_,data_stage_4__2126_,
  data_stage_4__2125_,data_stage_4__2124_,data_stage_4__2123_,data_stage_4__2122_,
  data_stage_4__2121_,data_stage_4__2120_,data_stage_4__2119_,data_stage_4__2118_,
  data_stage_4__2117_,data_stage_4__2116_,data_stage_4__2115_,data_stage_4__2114_,
  data_stage_4__2113_,data_stage_4__2112_,data_stage_4__2111_,data_stage_4__2110_,
  data_stage_4__2109_,data_stage_4__2108_,data_stage_4__2107_,data_stage_4__2106_,
  data_stage_4__2105_,data_stage_4__2104_,data_stage_4__2103_,data_stage_4__2102_,
  data_stage_4__2101_,data_stage_4__2100_,data_stage_4__2099_,data_stage_4__2098_,
  data_stage_4__2097_,data_stage_4__2096_,data_stage_4__2095_,data_stage_4__2094_,
  data_stage_4__2093_,data_stage_4__2092_,data_stage_4__2091_,data_stage_4__2090_,
  data_stage_4__2089_,data_stage_4__2088_,data_stage_4__2087_,data_stage_4__2086_,
  data_stage_4__2085_,data_stage_4__2084_,data_stage_4__2083_,data_stage_4__2082_,
  data_stage_4__2081_,data_stage_4__2080_,data_stage_4__2079_,data_stage_4__2078_,
  data_stage_4__2077_,data_stage_4__2076_,data_stage_4__2075_,data_stage_4__2074_,
  data_stage_4__2073_,data_stage_4__2072_,data_stage_4__2071_,data_stage_4__2070_,
  data_stage_4__2069_,data_stage_4__2068_,data_stage_4__2067_,data_stage_4__2066_,
  data_stage_4__2065_,data_stage_4__2064_,data_stage_4__2063_,data_stage_4__2062_,
  data_stage_4__2061_,data_stage_4__2060_,data_stage_4__2059_,data_stage_4__2058_,
  data_stage_4__2057_,data_stage_4__2056_,data_stage_4__2055_,data_stage_4__2054_,
  data_stage_4__2053_,data_stage_4__2052_,data_stage_4__2051_,data_stage_4__2050_,
  data_stage_4__2049_,data_stage_4__2048_,data_stage_4__2047_,data_stage_4__2046_,
  data_stage_4__2045_,data_stage_4__2044_,data_stage_4__2043_,data_stage_4__2042_,
  data_stage_4__2041_,data_stage_4__2040_,data_stage_4__2039_,data_stage_4__2038_,
  data_stage_4__2037_,data_stage_4__2036_,data_stage_4__2035_,data_stage_4__2034_,
  data_stage_4__2033_,data_stage_4__2032_,data_stage_4__2031_,data_stage_4__2030_,
  data_stage_4__2029_,data_stage_4__2028_,data_stage_4__2027_,data_stage_4__2026_,
  data_stage_4__2025_,data_stage_4__2024_,data_stage_4__2023_,data_stage_4__2022_,
  data_stage_4__2021_,data_stage_4__2020_,data_stage_4__2019_,data_stage_4__2018_,
  data_stage_4__2017_,data_stage_4__2016_,data_stage_4__2015_,data_stage_4__2014_,
  data_stage_4__2013_,data_stage_4__2012_,data_stage_4__2011_,data_stage_4__2010_,
  data_stage_4__2009_,data_stage_4__2008_,data_stage_4__2007_,data_stage_4__2006_,
  data_stage_4__2005_,data_stage_4__2004_,data_stage_4__2003_,data_stage_4__2002_,
  data_stage_4__2001_,data_stage_4__2000_,data_stage_4__1999_,data_stage_4__1998_,
  data_stage_4__1997_,data_stage_4__1996_,data_stage_4__1995_,data_stage_4__1994_,
  data_stage_4__1993_,data_stage_4__1992_,data_stage_4__1991_,data_stage_4__1990_,
  data_stage_4__1989_,data_stage_4__1988_,data_stage_4__1987_,data_stage_4__1986_,
  data_stage_4__1985_,data_stage_4__1984_,data_stage_4__1983_,data_stage_4__1982_,
  data_stage_4__1981_,data_stage_4__1980_,data_stage_4__1979_,data_stage_4__1978_,
  data_stage_4__1977_,data_stage_4__1976_,data_stage_4__1975_,data_stage_4__1974_,
  data_stage_4__1973_,data_stage_4__1972_,data_stage_4__1971_,data_stage_4__1970_,
  data_stage_4__1969_,data_stage_4__1968_,data_stage_4__1967_,data_stage_4__1966_,
  data_stage_4__1965_,data_stage_4__1964_,data_stage_4__1963_,data_stage_4__1962_,
  data_stage_4__1961_,data_stage_4__1960_,data_stage_4__1959_,data_stage_4__1958_,
  data_stage_4__1957_,data_stage_4__1956_,data_stage_4__1955_,data_stage_4__1954_,
  data_stage_4__1953_,data_stage_4__1952_,data_stage_4__1951_,data_stage_4__1950_,
  data_stage_4__1949_,data_stage_4__1948_,data_stage_4__1947_,data_stage_4__1946_,
  data_stage_4__1945_,data_stage_4__1944_,data_stage_4__1943_,data_stage_4__1942_,
  data_stage_4__1941_,data_stage_4__1940_,data_stage_4__1939_,data_stage_4__1938_,
  data_stage_4__1937_,data_stage_4__1936_,data_stage_4__1935_,data_stage_4__1934_,
  data_stage_4__1933_,data_stage_4__1932_,data_stage_4__1931_,data_stage_4__1930_,
  data_stage_4__1929_,data_stage_4__1928_,data_stage_4__1927_,data_stage_4__1926_,
  data_stage_4__1925_,data_stage_4__1924_,data_stage_4__1923_,data_stage_4__1922_,
  data_stage_4__1921_,data_stage_4__1920_,data_stage_4__1919_,data_stage_4__1918_,
  data_stage_4__1917_,data_stage_4__1916_,data_stage_4__1915_,data_stage_4__1914_,
  data_stage_4__1913_,data_stage_4__1912_,data_stage_4__1911_,data_stage_4__1910_,
  data_stage_4__1909_,data_stage_4__1908_,data_stage_4__1907_,data_stage_4__1906_,
  data_stage_4__1905_,data_stage_4__1904_,data_stage_4__1903_,data_stage_4__1902_,
  data_stage_4__1901_,data_stage_4__1900_,data_stage_4__1899_,data_stage_4__1898_,
  data_stage_4__1897_,data_stage_4__1896_,data_stage_4__1895_,data_stage_4__1894_,
  data_stage_4__1893_,data_stage_4__1892_,data_stage_4__1891_,data_stage_4__1890_,
  data_stage_4__1889_,data_stage_4__1888_,data_stage_4__1887_,data_stage_4__1886_,
  data_stage_4__1885_,data_stage_4__1884_,data_stage_4__1883_,data_stage_4__1882_,
  data_stage_4__1881_,data_stage_4__1880_,data_stage_4__1879_,data_stage_4__1878_,
  data_stage_4__1877_,data_stage_4__1876_,data_stage_4__1875_,data_stage_4__1874_,
  data_stage_4__1873_,data_stage_4__1872_,data_stage_4__1871_,data_stage_4__1870_,
  data_stage_4__1869_,data_stage_4__1868_,data_stage_4__1867_,data_stage_4__1866_,
  data_stage_4__1865_,data_stage_4__1864_,data_stage_4__1863_,data_stage_4__1862_,
  data_stage_4__1861_,data_stage_4__1860_,data_stage_4__1859_,data_stage_4__1858_,
  data_stage_4__1857_,data_stage_4__1856_,data_stage_4__1855_,data_stage_4__1854_,
  data_stage_4__1853_,data_stage_4__1852_,data_stage_4__1851_,data_stage_4__1850_,
  data_stage_4__1849_,data_stage_4__1848_,data_stage_4__1847_,data_stage_4__1846_,
  data_stage_4__1845_,data_stage_4__1844_,data_stage_4__1843_,data_stage_4__1842_,
  data_stage_4__1841_,data_stage_4__1840_,data_stage_4__1839_,data_stage_4__1838_,
  data_stage_4__1837_,data_stage_4__1836_,data_stage_4__1835_,data_stage_4__1834_,
  data_stage_4__1833_,data_stage_4__1832_,data_stage_4__1831_,data_stage_4__1830_,
  data_stage_4__1829_,data_stage_4__1828_,data_stage_4__1827_,data_stage_4__1826_,
  data_stage_4__1825_,data_stage_4__1824_,data_stage_4__1823_,data_stage_4__1822_,
  data_stage_4__1821_,data_stage_4__1820_,data_stage_4__1819_,data_stage_4__1818_,
  data_stage_4__1817_,data_stage_4__1816_,data_stage_4__1815_,data_stage_4__1814_,
  data_stage_4__1813_,data_stage_4__1812_,data_stage_4__1811_,data_stage_4__1810_,
  data_stage_4__1809_,data_stage_4__1808_,data_stage_4__1807_,data_stage_4__1806_,
  data_stage_4__1805_,data_stage_4__1804_,data_stage_4__1803_,data_stage_4__1802_,
  data_stage_4__1801_,data_stage_4__1800_,data_stage_4__1799_,data_stage_4__1798_,
  data_stage_4__1797_,data_stage_4__1796_,data_stage_4__1795_,data_stage_4__1794_,
  data_stage_4__1793_,data_stage_4__1792_,data_stage_4__1791_,data_stage_4__1790_,
  data_stage_4__1789_,data_stage_4__1788_,data_stage_4__1787_,data_stage_4__1786_,
  data_stage_4__1785_,data_stage_4__1784_,data_stage_4__1783_,data_stage_4__1782_,
  data_stage_4__1781_,data_stage_4__1780_,data_stage_4__1779_,data_stage_4__1778_,
  data_stage_4__1777_,data_stage_4__1776_,data_stage_4__1775_,data_stage_4__1774_,
  data_stage_4__1773_,data_stage_4__1772_,data_stage_4__1771_,data_stage_4__1770_,
  data_stage_4__1769_,data_stage_4__1768_,data_stage_4__1767_,data_stage_4__1766_,
  data_stage_4__1765_,data_stage_4__1764_,data_stage_4__1763_,data_stage_4__1762_,
  data_stage_4__1761_,data_stage_4__1760_,data_stage_4__1759_,data_stage_4__1758_,
  data_stage_4__1757_,data_stage_4__1756_,data_stage_4__1755_,data_stage_4__1754_,
  data_stage_4__1753_,data_stage_4__1752_,data_stage_4__1751_,data_stage_4__1750_,
  data_stage_4__1749_,data_stage_4__1748_,data_stage_4__1747_,data_stage_4__1746_,
  data_stage_4__1745_,data_stage_4__1744_,data_stage_4__1743_,data_stage_4__1742_,
  data_stage_4__1741_,data_stage_4__1740_,data_stage_4__1739_,data_stage_4__1738_,
  data_stage_4__1737_,data_stage_4__1736_,data_stage_4__1735_,data_stage_4__1734_,
  data_stage_4__1733_,data_stage_4__1732_,data_stage_4__1731_,data_stage_4__1730_,
  data_stage_4__1729_,data_stage_4__1728_,data_stage_4__1727_,data_stage_4__1726_,
  data_stage_4__1725_,data_stage_4__1724_,data_stage_4__1723_,data_stage_4__1722_,
  data_stage_4__1721_,data_stage_4__1720_,data_stage_4__1719_,data_stage_4__1718_,
  data_stage_4__1717_,data_stage_4__1716_,data_stage_4__1715_,data_stage_4__1714_,
  data_stage_4__1713_,data_stage_4__1712_,data_stage_4__1711_,data_stage_4__1710_,
  data_stage_4__1709_,data_stage_4__1708_,data_stage_4__1707_,data_stage_4__1706_,
  data_stage_4__1705_,data_stage_4__1704_,data_stage_4__1703_,data_stage_4__1702_,
  data_stage_4__1701_,data_stage_4__1700_,data_stage_4__1699_,data_stage_4__1698_,
  data_stage_4__1697_,data_stage_4__1696_,data_stage_4__1695_,data_stage_4__1694_,
  data_stage_4__1693_,data_stage_4__1692_,data_stage_4__1691_,data_stage_4__1690_,
  data_stage_4__1689_,data_stage_4__1688_,data_stage_4__1687_,data_stage_4__1686_,
  data_stage_4__1685_,data_stage_4__1684_,data_stage_4__1683_,data_stage_4__1682_,
  data_stage_4__1681_,data_stage_4__1680_,data_stage_4__1679_,data_stage_4__1678_,
  data_stage_4__1677_,data_stage_4__1676_,data_stage_4__1675_,data_stage_4__1674_,
  data_stage_4__1673_,data_stage_4__1672_,data_stage_4__1671_,data_stage_4__1670_,
  data_stage_4__1669_,data_stage_4__1668_,data_stage_4__1667_,data_stage_4__1666_,
  data_stage_4__1665_,data_stage_4__1664_,data_stage_4__1663_,data_stage_4__1662_,
  data_stage_4__1661_,data_stage_4__1660_,data_stage_4__1659_,data_stage_4__1658_,
  data_stage_4__1657_,data_stage_4__1656_,data_stage_4__1655_,data_stage_4__1654_,
  data_stage_4__1653_,data_stage_4__1652_,data_stage_4__1651_,data_stage_4__1650_,
  data_stage_4__1649_,data_stage_4__1648_,data_stage_4__1647_,data_stage_4__1646_,
  data_stage_4__1645_,data_stage_4__1644_,data_stage_4__1643_,data_stage_4__1642_,
  data_stage_4__1641_,data_stage_4__1640_,data_stage_4__1639_,data_stage_4__1638_,
  data_stage_4__1637_,data_stage_4__1636_,data_stage_4__1635_,data_stage_4__1634_,
  data_stage_4__1633_,data_stage_4__1632_,data_stage_4__1631_,data_stage_4__1630_,
  data_stage_4__1629_,data_stage_4__1628_,data_stage_4__1627_,data_stage_4__1626_,
  data_stage_4__1625_,data_stage_4__1624_,data_stage_4__1623_,data_stage_4__1622_,
  data_stage_4__1621_,data_stage_4__1620_,data_stage_4__1619_,data_stage_4__1618_,
  data_stage_4__1617_,data_stage_4__1616_,data_stage_4__1615_,data_stage_4__1614_,
  data_stage_4__1613_,data_stage_4__1612_,data_stage_4__1611_,data_stage_4__1610_,
  data_stage_4__1609_,data_stage_4__1608_,data_stage_4__1607_,data_stage_4__1606_,
  data_stage_4__1605_,data_stage_4__1604_,data_stage_4__1603_,data_stage_4__1602_,
  data_stage_4__1601_,data_stage_4__1600_,data_stage_4__1599_,data_stage_4__1598_,
  data_stage_4__1597_,data_stage_4__1596_,data_stage_4__1595_,data_stage_4__1594_,
  data_stage_4__1593_,data_stage_4__1592_,data_stage_4__1591_,data_stage_4__1590_,
  data_stage_4__1589_,data_stage_4__1588_,data_stage_4__1587_,data_stage_4__1586_,
  data_stage_4__1585_,data_stage_4__1584_,data_stage_4__1583_,data_stage_4__1582_,
  data_stage_4__1581_,data_stage_4__1580_,data_stage_4__1579_,data_stage_4__1578_,
  data_stage_4__1577_,data_stage_4__1576_,data_stage_4__1575_,data_stage_4__1574_,
  data_stage_4__1573_,data_stage_4__1572_,data_stage_4__1571_,data_stage_4__1570_,
  data_stage_4__1569_,data_stage_4__1568_,data_stage_4__1567_,data_stage_4__1566_,
  data_stage_4__1565_,data_stage_4__1564_,data_stage_4__1563_,data_stage_4__1562_,
  data_stage_4__1561_,data_stage_4__1560_,data_stage_4__1559_,data_stage_4__1558_,
  data_stage_4__1557_,data_stage_4__1556_,data_stage_4__1555_,data_stage_4__1554_,
  data_stage_4__1553_,data_stage_4__1552_,data_stage_4__1551_,data_stage_4__1550_,
  data_stage_4__1549_,data_stage_4__1548_,data_stage_4__1547_,data_stage_4__1546_,
  data_stage_4__1545_,data_stage_4__1544_,data_stage_4__1543_,data_stage_4__1542_,
  data_stage_4__1541_,data_stage_4__1540_,data_stage_4__1539_,data_stage_4__1538_,
  data_stage_4__1537_,data_stage_4__1536_,data_stage_4__1535_,data_stage_4__1534_,
  data_stage_4__1533_,data_stage_4__1532_,data_stage_4__1531_,data_stage_4__1530_,
  data_stage_4__1529_,data_stage_4__1528_,data_stage_4__1527_,data_stage_4__1526_,
  data_stage_4__1525_,data_stage_4__1524_,data_stage_4__1523_,data_stage_4__1522_,
  data_stage_4__1521_,data_stage_4__1520_,data_stage_4__1519_,data_stage_4__1518_,
  data_stage_4__1517_,data_stage_4__1516_,data_stage_4__1515_,data_stage_4__1514_,
  data_stage_4__1513_,data_stage_4__1512_,data_stage_4__1511_,data_stage_4__1510_,
  data_stage_4__1509_,data_stage_4__1508_,data_stage_4__1507_,data_stage_4__1506_,
  data_stage_4__1505_,data_stage_4__1504_,data_stage_4__1503_,data_stage_4__1502_,
  data_stage_4__1501_,data_stage_4__1500_,data_stage_4__1499_,data_stage_4__1498_,
  data_stage_4__1497_,data_stage_4__1496_,data_stage_4__1495_,data_stage_4__1494_,
  data_stage_4__1493_,data_stage_4__1492_,data_stage_4__1491_,data_stage_4__1490_,
  data_stage_4__1489_,data_stage_4__1488_,data_stage_4__1487_,data_stage_4__1486_,
  data_stage_4__1485_,data_stage_4__1484_,data_stage_4__1483_,data_stage_4__1482_,
  data_stage_4__1481_,data_stage_4__1480_,data_stage_4__1479_,data_stage_4__1478_,
  data_stage_4__1477_,data_stage_4__1476_,data_stage_4__1475_,data_stage_4__1474_,
  data_stage_4__1473_,data_stage_4__1472_,data_stage_4__1471_,data_stage_4__1470_,
  data_stage_4__1469_,data_stage_4__1468_,data_stage_4__1467_,data_stage_4__1466_,
  data_stage_4__1465_,data_stage_4__1464_,data_stage_4__1463_,data_stage_4__1462_,
  data_stage_4__1461_,data_stage_4__1460_,data_stage_4__1459_,data_stage_4__1458_,
  data_stage_4__1457_,data_stage_4__1456_,data_stage_4__1455_,data_stage_4__1454_,
  data_stage_4__1453_,data_stage_4__1452_,data_stage_4__1451_,data_stage_4__1450_,
  data_stage_4__1449_,data_stage_4__1448_,data_stage_4__1447_,data_stage_4__1446_,
  data_stage_4__1445_,data_stage_4__1444_,data_stage_4__1443_,data_stage_4__1442_,
  data_stage_4__1441_,data_stage_4__1440_,data_stage_4__1439_,data_stage_4__1438_,
  data_stage_4__1437_,data_stage_4__1436_,data_stage_4__1435_,data_stage_4__1434_,
  data_stage_4__1433_,data_stage_4__1432_,data_stage_4__1431_,data_stage_4__1430_,
  data_stage_4__1429_,data_stage_4__1428_,data_stage_4__1427_,data_stage_4__1426_,
  data_stage_4__1425_,data_stage_4__1424_,data_stage_4__1423_,data_stage_4__1422_,
  data_stage_4__1421_,data_stage_4__1420_,data_stage_4__1419_,data_stage_4__1418_,
  data_stage_4__1417_,data_stage_4__1416_,data_stage_4__1415_,data_stage_4__1414_,
  data_stage_4__1413_,data_stage_4__1412_,data_stage_4__1411_,data_stage_4__1410_,
  data_stage_4__1409_,data_stage_4__1408_,data_stage_4__1407_,data_stage_4__1406_,
  data_stage_4__1405_,data_stage_4__1404_,data_stage_4__1403_,data_stage_4__1402_,
  data_stage_4__1401_,data_stage_4__1400_,data_stage_4__1399_,data_stage_4__1398_,
  data_stage_4__1397_,data_stage_4__1396_,data_stage_4__1395_,data_stage_4__1394_,
  data_stage_4__1393_,data_stage_4__1392_,data_stage_4__1391_,data_stage_4__1390_,
  data_stage_4__1389_,data_stage_4__1388_,data_stage_4__1387_,data_stage_4__1386_,
  data_stage_4__1385_,data_stage_4__1384_,data_stage_4__1383_,data_stage_4__1382_,
  data_stage_4__1381_,data_stage_4__1380_,data_stage_4__1379_,data_stage_4__1378_,
  data_stage_4__1377_,data_stage_4__1376_,data_stage_4__1375_,data_stage_4__1374_,
  data_stage_4__1373_,data_stage_4__1372_,data_stage_4__1371_,data_stage_4__1370_,
  data_stage_4__1369_,data_stage_4__1368_,data_stage_4__1367_,data_stage_4__1366_,
  data_stage_4__1365_,data_stage_4__1364_,data_stage_4__1363_,data_stage_4__1362_,
  data_stage_4__1361_,data_stage_4__1360_,data_stage_4__1359_,data_stage_4__1358_,
  data_stage_4__1357_,data_stage_4__1356_,data_stage_4__1355_,data_stage_4__1354_,
  data_stage_4__1353_,data_stage_4__1352_,data_stage_4__1351_,data_stage_4__1350_,
  data_stage_4__1349_,data_stage_4__1348_,data_stage_4__1347_,data_stage_4__1346_,
  data_stage_4__1345_,data_stage_4__1344_,data_stage_4__1343_,data_stage_4__1342_,
  data_stage_4__1341_,data_stage_4__1340_,data_stage_4__1339_,data_stage_4__1338_,
  data_stage_4__1337_,data_stage_4__1336_,data_stage_4__1335_,data_stage_4__1334_,
  data_stage_4__1333_,data_stage_4__1332_,data_stage_4__1331_,data_stage_4__1330_,
  data_stage_4__1329_,data_stage_4__1328_,data_stage_4__1327_,data_stage_4__1326_,
  data_stage_4__1325_,data_stage_4__1324_,data_stage_4__1323_,data_stage_4__1322_,
  data_stage_4__1321_,data_stage_4__1320_,data_stage_4__1319_,data_stage_4__1318_,
  data_stage_4__1317_,data_stage_4__1316_,data_stage_4__1315_,data_stage_4__1314_,
  data_stage_4__1313_,data_stage_4__1312_,data_stage_4__1311_,data_stage_4__1310_,
  data_stage_4__1309_,data_stage_4__1308_,data_stage_4__1307_,data_stage_4__1306_,
  data_stage_4__1305_,data_stage_4__1304_,data_stage_4__1303_,data_stage_4__1302_,
  data_stage_4__1301_,data_stage_4__1300_,data_stage_4__1299_,data_stage_4__1298_,
  data_stage_4__1297_,data_stage_4__1296_,data_stage_4__1295_,data_stage_4__1294_,
  data_stage_4__1293_,data_stage_4__1292_,data_stage_4__1291_,data_stage_4__1290_,
  data_stage_4__1289_,data_stage_4__1288_,data_stage_4__1287_,data_stage_4__1286_,
  data_stage_4__1285_,data_stage_4__1284_,data_stage_4__1283_,data_stage_4__1282_,
  data_stage_4__1281_,data_stage_4__1280_,data_stage_4__1279_,data_stage_4__1278_,
  data_stage_4__1277_,data_stage_4__1276_,data_stage_4__1275_,data_stage_4__1274_,
  data_stage_4__1273_,data_stage_4__1272_,data_stage_4__1271_,data_stage_4__1270_,
  data_stage_4__1269_,data_stage_4__1268_,data_stage_4__1267_,data_stage_4__1266_,
  data_stage_4__1265_,data_stage_4__1264_,data_stage_4__1263_,data_stage_4__1262_,
  data_stage_4__1261_,data_stage_4__1260_,data_stage_4__1259_,data_stage_4__1258_,
  data_stage_4__1257_,data_stage_4__1256_,data_stage_4__1255_,data_stage_4__1254_,
  data_stage_4__1253_,data_stage_4__1252_,data_stage_4__1251_,data_stage_4__1250_,
  data_stage_4__1249_,data_stage_4__1248_,data_stage_4__1247_,data_stage_4__1246_,
  data_stage_4__1245_,data_stage_4__1244_,data_stage_4__1243_,data_stage_4__1242_,
  data_stage_4__1241_,data_stage_4__1240_,data_stage_4__1239_,data_stage_4__1238_,
  data_stage_4__1237_,data_stage_4__1236_,data_stage_4__1235_,data_stage_4__1234_,
  data_stage_4__1233_,data_stage_4__1232_,data_stage_4__1231_,data_stage_4__1230_,
  data_stage_4__1229_,data_stage_4__1228_,data_stage_4__1227_,data_stage_4__1226_,
  data_stage_4__1225_,data_stage_4__1224_,data_stage_4__1223_,data_stage_4__1222_,
  data_stage_4__1221_,data_stage_4__1220_,data_stage_4__1219_,data_stage_4__1218_,
  data_stage_4__1217_,data_stage_4__1216_,data_stage_4__1215_,data_stage_4__1214_,
  data_stage_4__1213_,data_stage_4__1212_,data_stage_4__1211_,data_stage_4__1210_,
  data_stage_4__1209_,data_stage_4__1208_,data_stage_4__1207_,data_stage_4__1206_,
  data_stage_4__1205_,data_stage_4__1204_,data_stage_4__1203_,data_stage_4__1202_,
  data_stage_4__1201_,data_stage_4__1200_,data_stage_4__1199_,data_stage_4__1198_,
  data_stage_4__1197_,data_stage_4__1196_,data_stage_4__1195_,data_stage_4__1194_,
  data_stage_4__1193_,data_stage_4__1192_,data_stage_4__1191_,data_stage_4__1190_,
  data_stage_4__1189_,data_stage_4__1188_,data_stage_4__1187_,data_stage_4__1186_,
  data_stage_4__1185_,data_stage_4__1184_,data_stage_4__1183_,data_stage_4__1182_,
  data_stage_4__1181_,data_stage_4__1180_,data_stage_4__1179_,data_stage_4__1178_,
  data_stage_4__1177_,data_stage_4__1176_,data_stage_4__1175_,data_stage_4__1174_,
  data_stage_4__1173_,data_stage_4__1172_,data_stage_4__1171_,data_stage_4__1170_,
  data_stage_4__1169_,data_stage_4__1168_,data_stage_4__1167_,data_stage_4__1166_,
  data_stage_4__1165_,data_stage_4__1164_,data_stage_4__1163_,data_stage_4__1162_,
  data_stage_4__1161_,data_stage_4__1160_,data_stage_4__1159_,data_stage_4__1158_,
  data_stage_4__1157_,data_stage_4__1156_,data_stage_4__1155_,data_stage_4__1154_,
  data_stage_4__1153_,data_stage_4__1152_,data_stage_4__1151_,data_stage_4__1150_,
  data_stage_4__1149_,data_stage_4__1148_,data_stage_4__1147_,data_stage_4__1146_,
  data_stage_4__1145_,data_stage_4__1144_,data_stage_4__1143_,data_stage_4__1142_,
  data_stage_4__1141_,data_stage_4__1140_,data_stage_4__1139_,data_stage_4__1138_,
  data_stage_4__1137_,data_stage_4__1136_,data_stage_4__1135_,data_stage_4__1134_,
  data_stage_4__1133_,data_stage_4__1132_,data_stage_4__1131_,data_stage_4__1130_,
  data_stage_4__1129_,data_stage_4__1128_,data_stage_4__1127_,data_stage_4__1126_,
  data_stage_4__1125_,data_stage_4__1124_,data_stage_4__1123_,data_stage_4__1122_,
  data_stage_4__1121_,data_stage_4__1120_,data_stage_4__1119_,data_stage_4__1118_,
  data_stage_4__1117_,data_stage_4__1116_,data_stage_4__1115_,data_stage_4__1114_,
  data_stage_4__1113_,data_stage_4__1112_,data_stage_4__1111_,data_stage_4__1110_,
  data_stage_4__1109_,data_stage_4__1108_,data_stage_4__1107_,data_stage_4__1106_,
  data_stage_4__1105_,data_stage_4__1104_,data_stage_4__1103_,data_stage_4__1102_,
  data_stage_4__1101_,data_stage_4__1100_,data_stage_4__1099_,data_stage_4__1098_,
  data_stage_4__1097_,data_stage_4__1096_,data_stage_4__1095_,data_stage_4__1094_,
  data_stage_4__1093_,data_stage_4__1092_,data_stage_4__1091_,data_stage_4__1090_,
  data_stage_4__1089_,data_stage_4__1088_,data_stage_4__1087_,data_stage_4__1086_,
  data_stage_4__1085_,data_stage_4__1084_,data_stage_4__1083_,data_stage_4__1082_,
  data_stage_4__1081_,data_stage_4__1080_,data_stage_4__1079_,data_stage_4__1078_,
  data_stage_4__1077_,data_stage_4__1076_,data_stage_4__1075_,data_stage_4__1074_,
  data_stage_4__1073_,data_stage_4__1072_,data_stage_4__1071_,data_stage_4__1070_,
  data_stage_4__1069_,data_stage_4__1068_,data_stage_4__1067_,data_stage_4__1066_,
  data_stage_4__1065_,data_stage_4__1064_,data_stage_4__1063_,data_stage_4__1062_,
  data_stage_4__1061_,data_stage_4__1060_,data_stage_4__1059_,data_stage_4__1058_,
  data_stage_4__1057_,data_stage_4__1056_,data_stage_4__1055_,data_stage_4__1054_,
  data_stage_4__1053_,data_stage_4__1052_,data_stage_4__1051_,data_stage_4__1050_,
  data_stage_4__1049_,data_stage_4__1048_,data_stage_4__1047_,data_stage_4__1046_,
  data_stage_4__1045_,data_stage_4__1044_,data_stage_4__1043_,data_stage_4__1042_,
  data_stage_4__1041_,data_stage_4__1040_,data_stage_4__1039_,data_stage_4__1038_,
  data_stage_4__1037_,data_stage_4__1036_,data_stage_4__1035_,data_stage_4__1034_,
  data_stage_4__1033_,data_stage_4__1032_,data_stage_4__1031_,data_stage_4__1030_,
  data_stage_4__1029_,data_stage_4__1028_,data_stage_4__1027_,data_stage_4__1026_,
  data_stage_4__1025_,data_stage_4__1024_,data_stage_4__1023_,data_stage_4__1022_,
  data_stage_4__1021_,data_stage_4__1020_,data_stage_4__1019_,data_stage_4__1018_,
  data_stage_4__1017_,data_stage_4__1016_,data_stage_4__1015_,data_stage_4__1014_,
  data_stage_4__1013_,data_stage_4__1012_,data_stage_4__1011_,data_stage_4__1010_,
  data_stage_4__1009_,data_stage_4__1008_,data_stage_4__1007_,data_stage_4__1006_,
  data_stage_4__1005_,data_stage_4__1004_,data_stage_4__1003_,data_stage_4__1002_,
  data_stage_4__1001_,data_stage_4__1000_,data_stage_4__999_,data_stage_4__998_,
  data_stage_4__997_,data_stage_4__996_,data_stage_4__995_,data_stage_4__994_,
  data_stage_4__993_,data_stage_4__992_,data_stage_4__991_,data_stage_4__990_,data_stage_4__989_,
  data_stage_4__988_,data_stage_4__987_,data_stage_4__986_,data_stage_4__985_,
  data_stage_4__984_,data_stage_4__983_,data_stage_4__982_,data_stage_4__981_,
  data_stage_4__980_,data_stage_4__979_,data_stage_4__978_,data_stage_4__977_,
  data_stage_4__976_,data_stage_4__975_,data_stage_4__974_,data_stage_4__973_,
  data_stage_4__972_,data_stage_4__971_,data_stage_4__970_,data_stage_4__969_,data_stage_4__968_,
  data_stage_4__967_,data_stage_4__966_,data_stage_4__965_,data_stage_4__964_,
  data_stage_4__963_,data_stage_4__962_,data_stage_4__961_,data_stage_4__960_,
  data_stage_4__959_,data_stage_4__958_,data_stage_4__957_,data_stage_4__956_,
  data_stage_4__955_,data_stage_4__954_,data_stage_4__953_,data_stage_4__952_,
  data_stage_4__951_,data_stage_4__950_,data_stage_4__949_,data_stage_4__948_,data_stage_4__947_,
  data_stage_4__946_,data_stage_4__945_,data_stage_4__944_,data_stage_4__943_,
  data_stage_4__942_,data_stage_4__941_,data_stage_4__940_,data_stage_4__939_,
  data_stage_4__938_,data_stage_4__937_,data_stage_4__936_,data_stage_4__935_,
  data_stage_4__934_,data_stage_4__933_,data_stage_4__932_,data_stage_4__931_,data_stage_4__930_,
  data_stage_4__929_,data_stage_4__928_,data_stage_4__927_,data_stage_4__926_,
  data_stage_4__925_,data_stage_4__924_,data_stage_4__923_,data_stage_4__922_,
  data_stage_4__921_,data_stage_4__920_,data_stage_4__919_,data_stage_4__918_,
  data_stage_4__917_,data_stage_4__916_,data_stage_4__915_,data_stage_4__914_,
  data_stage_4__913_,data_stage_4__912_,data_stage_4__911_,data_stage_4__910_,data_stage_4__909_,
  data_stage_4__908_,data_stage_4__907_,data_stage_4__906_,data_stage_4__905_,
  data_stage_4__904_,data_stage_4__903_,data_stage_4__902_,data_stage_4__901_,
  data_stage_4__900_,data_stage_4__899_,data_stage_4__898_,data_stage_4__897_,
  data_stage_4__896_,data_stage_4__895_,data_stage_4__894_,data_stage_4__893_,
  data_stage_4__892_,data_stage_4__891_,data_stage_4__890_,data_stage_4__889_,data_stage_4__888_,
  data_stage_4__887_,data_stage_4__886_,data_stage_4__885_,data_stage_4__884_,
  data_stage_4__883_,data_stage_4__882_,data_stage_4__881_,data_stage_4__880_,
  data_stage_4__879_,data_stage_4__878_,data_stage_4__877_,data_stage_4__876_,
  data_stage_4__875_,data_stage_4__874_,data_stage_4__873_,data_stage_4__872_,
  data_stage_4__871_,data_stage_4__870_,data_stage_4__869_,data_stage_4__868_,data_stage_4__867_,
  data_stage_4__866_,data_stage_4__865_,data_stage_4__864_,data_stage_4__863_,
  data_stage_4__862_,data_stage_4__861_,data_stage_4__860_,data_stage_4__859_,
  data_stage_4__858_,data_stage_4__857_,data_stage_4__856_,data_stage_4__855_,
  data_stage_4__854_,data_stage_4__853_,data_stage_4__852_,data_stage_4__851_,data_stage_4__850_,
  data_stage_4__849_,data_stage_4__848_,data_stage_4__847_,data_stage_4__846_,
  data_stage_4__845_,data_stage_4__844_,data_stage_4__843_,data_stage_4__842_,
  data_stage_4__841_,data_stage_4__840_,data_stage_4__839_,data_stage_4__838_,
  data_stage_4__837_,data_stage_4__836_,data_stage_4__835_,data_stage_4__834_,
  data_stage_4__833_,data_stage_4__832_,data_stage_4__831_,data_stage_4__830_,data_stage_4__829_,
  data_stage_4__828_,data_stage_4__827_,data_stage_4__826_,data_stage_4__825_,
  data_stage_4__824_,data_stage_4__823_,data_stage_4__822_,data_stage_4__821_,
  data_stage_4__820_,data_stage_4__819_,data_stage_4__818_,data_stage_4__817_,
  data_stage_4__816_,data_stage_4__815_,data_stage_4__814_,data_stage_4__813_,
  data_stage_4__812_,data_stage_4__811_,data_stage_4__810_,data_stage_4__809_,data_stage_4__808_,
  data_stage_4__807_,data_stage_4__806_,data_stage_4__805_,data_stage_4__804_,
  data_stage_4__803_,data_stage_4__802_,data_stage_4__801_,data_stage_4__800_,
  data_stage_4__799_,data_stage_4__798_,data_stage_4__797_,data_stage_4__796_,
  data_stage_4__795_,data_stage_4__794_,data_stage_4__793_,data_stage_4__792_,
  data_stage_4__791_,data_stage_4__790_,data_stage_4__789_,data_stage_4__788_,data_stage_4__787_,
  data_stage_4__786_,data_stage_4__785_,data_stage_4__784_,data_stage_4__783_,
  data_stage_4__782_,data_stage_4__781_,data_stage_4__780_,data_stage_4__779_,
  data_stage_4__778_,data_stage_4__777_,data_stage_4__776_,data_stage_4__775_,
  data_stage_4__774_,data_stage_4__773_,data_stage_4__772_,data_stage_4__771_,data_stage_4__770_,
  data_stage_4__769_,data_stage_4__768_,data_stage_4__767_,data_stage_4__766_,
  data_stage_4__765_,data_stage_4__764_,data_stage_4__763_,data_stage_4__762_,
  data_stage_4__761_,data_stage_4__760_,data_stage_4__759_,data_stage_4__758_,
  data_stage_4__757_,data_stage_4__756_,data_stage_4__755_,data_stage_4__754_,
  data_stage_4__753_,data_stage_4__752_,data_stage_4__751_,data_stage_4__750_,data_stage_4__749_,
  data_stage_4__748_,data_stage_4__747_,data_stage_4__746_,data_stage_4__745_,
  data_stage_4__744_,data_stage_4__743_,data_stage_4__742_,data_stage_4__741_,
  data_stage_4__740_,data_stage_4__739_,data_stage_4__738_,data_stage_4__737_,
  data_stage_4__736_,data_stage_4__735_,data_stage_4__734_,data_stage_4__733_,
  data_stage_4__732_,data_stage_4__731_,data_stage_4__730_,data_stage_4__729_,data_stage_4__728_,
  data_stage_4__727_,data_stage_4__726_,data_stage_4__725_,data_stage_4__724_,
  data_stage_4__723_,data_stage_4__722_,data_stage_4__721_,data_stage_4__720_,
  data_stage_4__719_,data_stage_4__718_,data_stage_4__717_,data_stage_4__716_,
  data_stage_4__715_,data_stage_4__714_,data_stage_4__713_,data_stage_4__712_,
  data_stage_4__711_,data_stage_4__710_,data_stage_4__709_,data_stage_4__708_,data_stage_4__707_,
  data_stage_4__706_,data_stage_4__705_,data_stage_4__704_,data_stage_4__703_,
  data_stage_4__702_,data_stage_4__701_,data_stage_4__700_,data_stage_4__699_,
  data_stage_4__698_,data_stage_4__697_,data_stage_4__696_,data_stage_4__695_,
  data_stage_4__694_,data_stage_4__693_,data_stage_4__692_,data_stage_4__691_,data_stage_4__690_,
  data_stage_4__689_,data_stage_4__688_,data_stage_4__687_,data_stage_4__686_,
  data_stage_4__685_,data_stage_4__684_,data_stage_4__683_,data_stage_4__682_,
  data_stage_4__681_,data_stage_4__680_,data_stage_4__679_,data_stage_4__678_,
  data_stage_4__677_,data_stage_4__676_,data_stage_4__675_,data_stage_4__674_,
  data_stage_4__673_,data_stage_4__672_,data_stage_4__671_,data_stage_4__670_,data_stage_4__669_,
  data_stage_4__668_,data_stage_4__667_,data_stage_4__666_,data_stage_4__665_,
  data_stage_4__664_,data_stage_4__663_,data_stage_4__662_,data_stage_4__661_,
  data_stage_4__660_,data_stage_4__659_,data_stage_4__658_,data_stage_4__657_,
  data_stage_4__656_,data_stage_4__655_,data_stage_4__654_,data_stage_4__653_,
  data_stage_4__652_,data_stage_4__651_,data_stage_4__650_,data_stage_4__649_,data_stage_4__648_,
  data_stage_4__647_,data_stage_4__646_,data_stage_4__645_,data_stage_4__644_,
  data_stage_4__643_,data_stage_4__642_,data_stage_4__641_,data_stage_4__640_,
  data_stage_4__639_,data_stage_4__638_,data_stage_4__637_,data_stage_4__636_,
  data_stage_4__635_,data_stage_4__634_,data_stage_4__633_,data_stage_4__632_,
  data_stage_4__631_,data_stage_4__630_,data_stage_4__629_,data_stage_4__628_,data_stage_4__627_,
  data_stage_4__626_,data_stage_4__625_,data_stage_4__624_,data_stage_4__623_,
  data_stage_4__622_,data_stage_4__621_,data_stage_4__620_,data_stage_4__619_,
  data_stage_4__618_,data_stage_4__617_,data_stage_4__616_,data_stage_4__615_,
  data_stage_4__614_,data_stage_4__613_,data_stage_4__612_,data_stage_4__611_,data_stage_4__610_,
  data_stage_4__609_,data_stage_4__608_,data_stage_4__607_,data_stage_4__606_,
  data_stage_4__605_,data_stage_4__604_,data_stage_4__603_,data_stage_4__602_,
  data_stage_4__601_,data_stage_4__600_,data_stage_4__599_,data_stage_4__598_,
  data_stage_4__597_,data_stage_4__596_,data_stage_4__595_,data_stage_4__594_,
  data_stage_4__593_,data_stage_4__592_,data_stage_4__591_,data_stage_4__590_,data_stage_4__589_,
  data_stage_4__588_,data_stage_4__587_,data_stage_4__586_,data_stage_4__585_,
  data_stage_4__584_,data_stage_4__583_,data_stage_4__582_,data_stage_4__581_,
  data_stage_4__580_,data_stage_4__579_,data_stage_4__578_,data_stage_4__577_,
  data_stage_4__576_,data_stage_4__575_,data_stage_4__574_,data_stage_4__573_,
  data_stage_4__572_,data_stage_4__571_,data_stage_4__570_,data_stage_4__569_,data_stage_4__568_,
  data_stage_4__567_,data_stage_4__566_,data_stage_4__565_,data_stage_4__564_,
  data_stage_4__563_,data_stage_4__562_,data_stage_4__561_,data_stage_4__560_,
  data_stage_4__559_,data_stage_4__558_,data_stage_4__557_,data_stage_4__556_,
  data_stage_4__555_,data_stage_4__554_,data_stage_4__553_,data_stage_4__552_,
  data_stage_4__551_,data_stage_4__550_,data_stage_4__549_,data_stage_4__548_,data_stage_4__547_,
  data_stage_4__546_,data_stage_4__545_,data_stage_4__544_,data_stage_4__543_,
  data_stage_4__542_,data_stage_4__541_,data_stage_4__540_,data_stage_4__539_,
  data_stage_4__538_,data_stage_4__537_,data_stage_4__536_,data_stage_4__535_,
  data_stage_4__534_,data_stage_4__533_,data_stage_4__532_,data_stage_4__531_,data_stage_4__530_,
  data_stage_4__529_,data_stage_4__528_,data_stage_4__527_,data_stage_4__526_,
  data_stage_4__525_,data_stage_4__524_,data_stage_4__523_,data_stage_4__522_,
  data_stage_4__521_,data_stage_4__520_,data_stage_4__519_,data_stage_4__518_,
  data_stage_4__517_,data_stage_4__516_,data_stage_4__515_,data_stage_4__514_,
  data_stage_4__513_,data_stage_4__512_,data_stage_4__511_,data_stage_4__510_,data_stage_4__509_,
  data_stage_4__508_,data_stage_4__507_,data_stage_4__506_,data_stage_4__505_,
  data_stage_4__504_,data_stage_4__503_,data_stage_4__502_,data_stage_4__501_,
  data_stage_4__500_,data_stage_4__499_,data_stage_4__498_,data_stage_4__497_,
  data_stage_4__496_,data_stage_4__495_,data_stage_4__494_,data_stage_4__493_,
  data_stage_4__492_,data_stage_4__491_,data_stage_4__490_,data_stage_4__489_,data_stage_4__488_,
  data_stage_4__487_,data_stage_4__486_,data_stage_4__485_,data_stage_4__484_,
  data_stage_4__483_,data_stage_4__482_,data_stage_4__481_,data_stage_4__480_,
  data_stage_4__479_,data_stage_4__478_,data_stage_4__477_,data_stage_4__476_,
  data_stage_4__475_,data_stage_4__474_,data_stage_4__473_,data_stage_4__472_,
  data_stage_4__471_,data_stage_4__470_,data_stage_4__469_,data_stage_4__468_,data_stage_4__467_,
  data_stage_4__466_,data_stage_4__465_,data_stage_4__464_,data_stage_4__463_,
  data_stage_4__462_,data_stage_4__461_,data_stage_4__460_,data_stage_4__459_,
  data_stage_4__458_,data_stage_4__457_,data_stage_4__456_,data_stage_4__455_,
  data_stage_4__454_,data_stage_4__453_,data_stage_4__452_,data_stage_4__451_,data_stage_4__450_,
  data_stage_4__449_,data_stage_4__448_,data_stage_4__447_,data_stage_4__446_,
  data_stage_4__445_,data_stage_4__444_,data_stage_4__443_,data_stage_4__442_,
  data_stage_4__441_,data_stage_4__440_,data_stage_4__439_,data_stage_4__438_,
  data_stage_4__437_,data_stage_4__436_,data_stage_4__435_,data_stage_4__434_,
  data_stage_4__433_,data_stage_4__432_,data_stage_4__431_,data_stage_4__430_,data_stage_4__429_,
  data_stage_4__428_,data_stage_4__427_,data_stage_4__426_,data_stage_4__425_,
  data_stage_4__424_,data_stage_4__423_,data_stage_4__422_,data_stage_4__421_,
  data_stage_4__420_,data_stage_4__419_,data_stage_4__418_,data_stage_4__417_,
  data_stage_4__416_,data_stage_4__415_,data_stage_4__414_,data_stage_4__413_,
  data_stage_4__412_,data_stage_4__411_,data_stage_4__410_,data_stage_4__409_,data_stage_4__408_,
  data_stage_4__407_,data_stage_4__406_,data_stage_4__405_,data_stage_4__404_,
  data_stage_4__403_,data_stage_4__402_,data_stage_4__401_,data_stage_4__400_,
  data_stage_4__399_,data_stage_4__398_,data_stage_4__397_,data_stage_4__396_,
  data_stage_4__395_,data_stage_4__394_,data_stage_4__393_,data_stage_4__392_,
  data_stage_4__391_,data_stage_4__390_,data_stage_4__389_,data_stage_4__388_,data_stage_4__387_,
  data_stage_4__386_,data_stage_4__385_,data_stage_4__384_,data_stage_4__383_,
  data_stage_4__382_,data_stage_4__381_,data_stage_4__380_,data_stage_4__379_,
  data_stage_4__378_,data_stage_4__377_,data_stage_4__376_,data_stage_4__375_,
  data_stage_4__374_,data_stage_4__373_,data_stage_4__372_,data_stage_4__371_,data_stage_4__370_,
  data_stage_4__369_,data_stage_4__368_,data_stage_4__367_,data_stage_4__366_,
  data_stage_4__365_,data_stage_4__364_,data_stage_4__363_,data_stage_4__362_,
  data_stage_4__361_,data_stage_4__360_,data_stage_4__359_,data_stage_4__358_,
  data_stage_4__357_,data_stage_4__356_,data_stage_4__355_,data_stage_4__354_,
  data_stage_4__353_,data_stage_4__352_,data_stage_4__351_,data_stage_4__350_,data_stage_4__349_,
  data_stage_4__348_,data_stage_4__347_,data_stage_4__346_,data_stage_4__345_,
  data_stage_4__344_,data_stage_4__343_,data_stage_4__342_,data_stage_4__341_,
  data_stage_4__340_,data_stage_4__339_,data_stage_4__338_,data_stage_4__337_,
  data_stage_4__336_,data_stage_4__335_,data_stage_4__334_,data_stage_4__333_,
  data_stage_4__332_,data_stage_4__331_,data_stage_4__330_,data_stage_4__329_,data_stage_4__328_,
  data_stage_4__327_,data_stage_4__326_,data_stage_4__325_,data_stage_4__324_,
  data_stage_4__323_,data_stage_4__322_,data_stage_4__321_,data_stage_4__320_,
  data_stage_4__319_,data_stage_4__318_,data_stage_4__317_,data_stage_4__316_,
  data_stage_4__315_,data_stage_4__314_,data_stage_4__313_,data_stage_4__312_,
  data_stage_4__311_,data_stage_4__310_,data_stage_4__309_,data_stage_4__308_,data_stage_4__307_,
  data_stage_4__306_,data_stage_4__305_,data_stage_4__304_,data_stage_4__303_,
  data_stage_4__302_,data_stage_4__301_,data_stage_4__300_,data_stage_4__299_,
  data_stage_4__298_,data_stage_4__297_,data_stage_4__296_,data_stage_4__295_,
  data_stage_4__294_,data_stage_4__293_,data_stage_4__292_,data_stage_4__291_,data_stage_4__290_,
  data_stage_4__289_,data_stage_4__288_,data_stage_4__287_,data_stage_4__286_,
  data_stage_4__285_,data_stage_4__284_,data_stage_4__283_,data_stage_4__282_,
  data_stage_4__281_,data_stage_4__280_,data_stage_4__279_,data_stage_4__278_,
  data_stage_4__277_,data_stage_4__276_,data_stage_4__275_,data_stage_4__274_,
  data_stage_4__273_,data_stage_4__272_,data_stage_4__271_,data_stage_4__270_,data_stage_4__269_,
  data_stage_4__268_,data_stage_4__267_,data_stage_4__266_,data_stage_4__265_,
  data_stage_4__264_,data_stage_4__263_,data_stage_4__262_,data_stage_4__261_,
  data_stage_4__260_,data_stage_4__259_,data_stage_4__258_,data_stage_4__257_,
  data_stage_4__256_,data_stage_4__255_,data_stage_4__254_,data_stage_4__253_,
  data_stage_4__252_,data_stage_4__251_,data_stage_4__250_,data_stage_4__249_,data_stage_4__248_,
  data_stage_4__247_,data_stage_4__246_,data_stage_4__245_,data_stage_4__244_,
  data_stage_4__243_,data_stage_4__242_,data_stage_4__241_,data_stage_4__240_,
  data_stage_4__239_,data_stage_4__238_,data_stage_4__237_,data_stage_4__236_,
  data_stage_4__235_,data_stage_4__234_,data_stage_4__233_,data_stage_4__232_,
  data_stage_4__231_,data_stage_4__230_,data_stage_4__229_,data_stage_4__228_,data_stage_4__227_,
  data_stage_4__226_,data_stage_4__225_,data_stage_4__224_,data_stage_4__223_,
  data_stage_4__222_,data_stage_4__221_,data_stage_4__220_,data_stage_4__219_,
  data_stage_4__218_,data_stage_4__217_,data_stage_4__216_,data_stage_4__215_,
  data_stage_4__214_,data_stage_4__213_,data_stage_4__212_,data_stage_4__211_,data_stage_4__210_,
  data_stage_4__209_,data_stage_4__208_,data_stage_4__207_,data_stage_4__206_,
  data_stage_4__205_,data_stage_4__204_,data_stage_4__203_,data_stage_4__202_,
  data_stage_4__201_,data_stage_4__200_,data_stage_4__199_,data_stage_4__198_,
  data_stage_4__197_,data_stage_4__196_,data_stage_4__195_,data_stage_4__194_,
  data_stage_4__193_,data_stage_4__192_,data_stage_4__191_,data_stage_4__190_,data_stage_4__189_,
  data_stage_4__188_,data_stage_4__187_,data_stage_4__186_,data_stage_4__185_,
  data_stage_4__184_,data_stage_4__183_,data_stage_4__182_,data_stage_4__181_,
  data_stage_4__180_,data_stage_4__179_,data_stage_4__178_,data_stage_4__177_,
  data_stage_4__176_,data_stage_4__175_,data_stage_4__174_,data_stage_4__173_,
  data_stage_4__172_,data_stage_4__171_,data_stage_4__170_,data_stage_4__169_,data_stage_4__168_,
  data_stage_4__167_,data_stage_4__166_,data_stage_4__165_,data_stage_4__164_,
  data_stage_4__163_,data_stage_4__162_,data_stage_4__161_,data_stage_4__160_,
  data_stage_4__159_,data_stage_4__158_,data_stage_4__157_,data_stage_4__156_,
  data_stage_4__155_,data_stage_4__154_,data_stage_4__153_,data_stage_4__152_,
  data_stage_4__151_,data_stage_4__150_,data_stage_4__149_,data_stage_4__148_,data_stage_4__147_,
  data_stage_4__146_,data_stage_4__145_,data_stage_4__144_,data_stage_4__143_,
  data_stage_4__142_,data_stage_4__141_,data_stage_4__140_,data_stage_4__139_,
  data_stage_4__138_,data_stage_4__137_,data_stage_4__136_,data_stage_4__135_,
  data_stage_4__134_,data_stage_4__133_,data_stage_4__132_,data_stage_4__131_,data_stage_4__130_,
  data_stage_4__129_,data_stage_4__128_,data_stage_4__127_,data_stage_4__126_,
  data_stage_4__125_,data_stage_4__124_,data_stage_4__123_,data_stage_4__122_,
  data_stage_4__121_,data_stage_4__120_,data_stage_4__119_,data_stage_4__118_,
  data_stage_4__117_,data_stage_4__116_,data_stage_4__115_,data_stage_4__114_,
  data_stage_4__113_,data_stage_4__112_,data_stage_4__111_,data_stage_4__110_,data_stage_4__109_,
  data_stage_4__108_,data_stage_4__107_,data_stage_4__106_,data_stage_4__105_,
  data_stage_4__104_,data_stage_4__103_,data_stage_4__102_,data_stage_4__101_,
  data_stage_4__100_,data_stage_4__99_,data_stage_4__98_,data_stage_4__97_,
  data_stage_4__96_,data_stage_4__95_,data_stage_4__94_,data_stage_4__93_,data_stage_4__92_,
  data_stage_4__91_,data_stage_4__90_,data_stage_4__89_,data_stage_4__88_,
  data_stage_4__87_,data_stage_4__86_,data_stage_4__85_,data_stage_4__84_,data_stage_4__83_,
  data_stage_4__82_,data_stage_4__81_,data_stage_4__80_,data_stage_4__79_,
  data_stage_4__78_,data_stage_4__77_,data_stage_4__76_,data_stage_4__75_,data_stage_4__74_,
  data_stage_4__73_,data_stage_4__72_,data_stage_4__71_,data_stage_4__70_,
  data_stage_4__69_,data_stage_4__68_,data_stage_4__67_,data_stage_4__66_,data_stage_4__65_,
  data_stage_4__64_,data_stage_4__63_,data_stage_4__62_,data_stage_4__61_,
  data_stage_4__60_,data_stage_4__59_,data_stage_4__58_,data_stage_4__57_,
  data_stage_4__56_,data_stage_4__55_,data_stage_4__54_,data_stage_4__53_,data_stage_4__52_,
  data_stage_4__51_,data_stage_4__50_,data_stage_4__49_,data_stage_4__48_,
  data_stage_4__47_,data_stage_4__46_,data_stage_4__45_,data_stage_4__44_,data_stage_4__43_,
  data_stage_4__42_,data_stage_4__41_,data_stage_4__40_,data_stage_4__39_,
  data_stage_4__38_,data_stage_4__37_,data_stage_4__36_,data_stage_4__35_,data_stage_4__34_,
  data_stage_4__33_,data_stage_4__32_,data_stage_4__31_,data_stage_4__30_,
  data_stage_4__29_,data_stage_4__28_,data_stage_4__27_,data_stage_4__26_,data_stage_4__25_,
  data_stage_4__24_,data_stage_4__23_,data_stage_4__22_,data_stage_4__21_,
  data_stage_4__20_,data_stage_4__19_,data_stage_4__18_,data_stage_4__17_,
  data_stage_4__16_,data_stage_4__15_,data_stage_4__14_,data_stage_4__13_,data_stage_4__12_,
  data_stage_4__11_,data_stage_4__10_,data_stage_4__9_,data_stage_4__8_,
  data_stage_4__7_,data_stage_4__6_,data_stage_4__5_,data_stage_4__4_,data_stage_4__3_,
  data_stage_4__2_,data_stage_4__1_,data_stage_4__0_,data_stage_5__8191_,data_stage_5__8190_,
  data_stage_5__8189_,data_stage_5__8188_,data_stage_5__8187_,data_stage_5__8186_,
  data_stage_5__8185_,data_stage_5__8184_,data_stage_5__8183_,data_stage_5__8182_,
  data_stage_5__8181_,data_stage_5__8180_,data_stage_5__8179_,data_stage_5__8178_,
  data_stage_5__8177_,data_stage_5__8176_,data_stage_5__8175_,data_stage_5__8174_,
  data_stage_5__8173_,data_stage_5__8172_,data_stage_5__8171_,data_stage_5__8170_,
  data_stage_5__8169_,data_stage_5__8168_,data_stage_5__8167_,data_stage_5__8166_,
  data_stage_5__8165_,data_stage_5__8164_,data_stage_5__8163_,data_stage_5__8162_,
  data_stage_5__8161_,data_stage_5__8160_,data_stage_5__8159_,data_stage_5__8158_,
  data_stage_5__8157_,data_stage_5__8156_,data_stage_5__8155_,data_stage_5__8154_,
  data_stage_5__8153_,data_stage_5__8152_,data_stage_5__8151_,data_stage_5__8150_,
  data_stage_5__8149_,data_stage_5__8148_,data_stage_5__8147_,data_stage_5__8146_,
  data_stage_5__8145_,data_stage_5__8144_,data_stage_5__8143_,data_stage_5__8142_,
  data_stage_5__8141_,data_stage_5__8140_,data_stage_5__8139_,data_stage_5__8138_,
  data_stage_5__8137_,data_stage_5__8136_,data_stage_5__8135_,data_stage_5__8134_,
  data_stage_5__8133_,data_stage_5__8132_,data_stage_5__8131_,data_stage_5__8130_,
  data_stage_5__8129_,data_stage_5__8128_,data_stage_5__8127_,data_stage_5__8126_,
  data_stage_5__8125_,data_stage_5__8124_,data_stage_5__8123_,data_stage_5__8122_,
  data_stage_5__8121_,data_stage_5__8120_,data_stage_5__8119_,data_stage_5__8118_,
  data_stage_5__8117_,data_stage_5__8116_,data_stage_5__8115_,data_stage_5__8114_,
  data_stage_5__8113_,data_stage_5__8112_,data_stage_5__8111_,data_stage_5__8110_,
  data_stage_5__8109_,data_stage_5__8108_,data_stage_5__8107_,data_stage_5__8106_,
  data_stage_5__8105_,data_stage_5__8104_,data_stage_5__8103_,data_stage_5__8102_,
  data_stage_5__8101_,data_stage_5__8100_,data_stage_5__8099_,data_stage_5__8098_,
  data_stage_5__8097_,data_stage_5__8096_,data_stage_5__8095_,data_stage_5__8094_,
  data_stage_5__8093_,data_stage_5__8092_,data_stage_5__8091_,data_stage_5__8090_,
  data_stage_5__8089_,data_stage_5__8088_,data_stage_5__8087_,data_stage_5__8086_,
  data_stage_5__8085_,data_stage_5__8084_,data_stage_5__8083_,data_stage_5__8082_,
  data_stage_5__8081_,data_stage_5__8080_,data_stage_5__8079_,data_stage_5__8078_,
  data_stage_5__8077_,data_stage_5__8076_,data_stage_5__8075_,data_stage_5__8074_,
  data_stage_5__8073_,data_stage_5__8072_,data_stage_5__8071_,data_stage_5__8070_,
  data_stage_5__8069_,data_stage_5__8068_,data_stage_5__8067_,data_stage_5__8066_,
  data_stage_5__8065_,data_stage_5__8064_,data_stage_5__8063_,data_stage_5__8062_,
  data_stage_5__8061_,data_stage_5__8060_,data_stage_5__8059_,data_stage_5__8058_,
  data_stage_5__8057_,data_stage_5__8056_,data_stage_5__8055_,data_stage_5__8054_,
  data_stage_5__8053_,data_stage_5__8052_,data_stage_5__8051_,data_stage_5__8050_,
  data_stage_5__8049_,data_stage_5__8048_,data_stage_5__8047_,data_stage_5__8046_,
  data_stage_5__8045_,data_stage_5__8044_,data_stage_5__8043_,data_stage_5__8042_,
  data_stage_5__8041_,data_stage_5__8040_,data_stage_5__8039_,data_stage_5__8038_,
  data_stage_5__8037_,data_stage_5__8036_,data_stage_5__8035_,data_stage_5__8034_,
  data_stage_5__8033_,data_stage_5__8032_,data_stage_5__8031_,data_stage_5__8030_,
  data_stage_5__8029_,data_stage_5__8028_,data_stage_5__8027_,data_stage_5__8026_,
  data_stage_5__8025_,data_stage_5__8024_,data_stage_5__8023_,data_stage_5__8022_,
  data_stage_5__8021_,data_stage_5__8020_,data_stage_5__8019_,data_stage_5__8018_,
  data_stage_5__8017_,data_stage_5__8016_,data_stage_5__8015_,data_stage_5__8014_,
  data_stage_5__8013_,data_stage_5__8012_,data_stage_5__8011_,data_stage_5__8010_,
  data_stage_5__8009_,data_stage_5__8008_,data_stage_5__8007_,data_stage_5__8006_,
  data_stage_5__8005_,data_stage_5__8004_,data_stage_5__8003_,data_stage_5__8002_,
  data_stage_5__8001_,data_stage_5__8000_,data_stage_5__7999_,data_stage_5__7998_,
  data_stage_5__7997_,data_stage_5__7996_,data_stage_5__7995_,data_stage_5__7994_,
  data_stage_5__7993_,data_stage_5__7992_,data_stage_5__7991_,data_stage_5__7990_,
  data_stage_5__7989_,data_stage_5__7988_,data_stage_5__7987_,data_stage_5__7986_,
  data_stage_5__7985_,data_stage_5__7984_,data_stage_5__7983_,data_stage_5__7982_,
  data_stage_5__7981_,data_stage_5__7980_,data_stage_5__7979_,data_stage_5__7978_,
  data_stage_5__7977_,data_stage_5__7976_,data_stage_5__7975_,data_stage_5__7974_,
  data_stage_5__7973_,data_stage_5__7972_,data_stage_5__7971_,data_stage_5__7970_,
  data_stage_5__7969_,data_stage_5__7968_,data_stage_5__7967_,data_stage_5__7966_,
  data_stage_5__7965_,data_stage_5__7964_,data_stage_5__7963_,data_stage_5__7962_,
  data_stage_5__7961_,data_stage_5__7960_,data_stage_5__7959_,data_stage_5__7958_,
  data_stage_5__7957_,data_stage_5__7956_,data_stage_5__7955_,data_stage_5__7954_,
  data_stage_5__7953_,data_stage_5__7952_,data_stage_5__7951_,data_stage_5__7950_,
  data_stage_5__7949_,data_stage_5__7948_,data_stage_5__7947_,data_stage_5__7946_,
  data_stage_5__7945_,data_stage_5__7944_,data_stage_5__7943_,data_stage_5__7942_,
  data_stage_5__7941_,data_stage_5__7940_,data_stage_5__7939_,data_stage_5__7938_,
  data_stage_5__7937_,data_stage_5__7936_,data_stage_5__7935_,data_stage_5__7934_,
  data_stage_5__7933_,data_stage_5__7932_,data_stage_5__7931_,data_stage_5__7930_,
  data_stage_5__7929_,data_stage_5__7928_,data_stage_5__7927_,data_stage_5__7926_,
  data_stage_5__7925_,data_stage_5__7924_,data_stage_5__7923_,data_stage_5__7922_,
  data_stage_5__7921_,data_stage_5__7920_,data_stage_5__7919_,data_stage_5__7918_,
  data_stage_5__7917_,data_stage_5__7916_,data_stage_5__7915_,data_stage_5__7914_,
  data_stage_5__7913_,data_stage_5__7912_,data_stage_5__7911_,data_stage_5__7910_,
  data_stage_5__7909_,data_stage_5__7908_,data_stage_5__7907_,data_stage_5__7906_,
  data_stage_5__7905_,data_stage_5__7904_,data_stage_5__7903_,data_stage_5__7902_,
  data_stage_5__7901_,data_stage_5__7900_,data_stage_5__7899_,data_stage_5__7898_,
  data_stage_5__7897_,data_stage_5__7896_,data_stage_5__7895_,data_stage_5__7894_,
  data_stage_5__7893_,data_stage_5__7892_,data_stage_5__7891_,data_stage_5__7890_,
  data_stage_5__7889_,data_stage_5__7888_,data_stage_5__7887_,data_stage_5__7886_,
  data_stage_5__7885_,data_stage_5__7884_,data_stage_5__7883_,data_stage_5__7882_,
  data_stage_5__7881_,data_stage_5__7880_,data_stage_5__7879_,data_stage_5__7878_,
  data_stage_5__7877_,data_stage_5__7876_,data_stage_5__7875_,data_stage_5__7874_,
  data_stage_5__7873_,data_stage_5__7872_,data_stage_5__7871_,data_stage_5__7870_,
  data_stage_5__7869_,data_stage_5__7868_,data_stage_5__7867_,data_stage_5__7866_,
  data_stage_5__7865_,data_stage_5__7864_,data_stage_5__7863_,data_stage_5__7862_,
  data_stage_5__7861_,data_stage_5__7860_,data_stage_5__7859_,data_stage_5__7858_,
  data_stage_5__7857_,data_stage_5__7856_,data_stage_5__7855_,data_stage_5__7854_,
  data_stage_5__7853_,data_stage_5__7852_,data_stage_5__7851_,data_stage_5__7850_,
  data_stage_5__7849_,data_stage_5__7848_,data_stage_5__7847_,data_stage_5__7846_,
  data_stage_5__7845_,data_stage_5__7844_,data_stage_5__7843_,data_stage_5__7842_,
  data_stage_5__7841_,data_stage_5__7840_,data_stage_5__7839_,data_stage_5__7838_,
  data_stage_5__7837_,data_stage_5__7836_,data_stage_5__7835_,data_stage_5__7834_,
  data_stage_5__7833_,data_stage_5__7832_,data_stage_5__7831_,data_stage_5__7830_,
  data_stage_5__7829_,data_stage_5__7828_,data_stage_5__7827_,data_stage_5__7826_,
  data_stage_5__7825_,data_stage_5__7824_,data_stage_5__7823_,data_stage_5__7822_,
  data_stage_5__7821_,data_stage_5__7820_,data_stage_5__7819_,data_stage_5__7818_,
  data_stage_5__7817_,data_stage_5__7816_,data_stage_5__7815_,data_stage_5__7814_,
  data_stage_5__7813_,data_stage_5__7812_,data_stage_5__7811_,data_stage_5__7810_,
  data_stage_5__7809_,data_stage_5__7808_,data_stage_5__7807_,data_stage_5__7806_,
  data_stage_5__7805_,data_stage_5__7804_,data_stage_5__7803_,data_stage_5__7802_,
  data_stage_5__7801_,data_stage_5__7800_,data_stage_5__7799_,data_stage_5__7798_,
  data_stage_5__7797_,data_stage_5__7796_,data_stage_5__7795_,data_stage_5__7794_,
  data_stage_5__7793_,data_stage_5__7792_,data_stage_5__7791_,data_stage_5__7790_,
  data_stage_5__7789_,data_stage_5__7788_,data_stage_5__7787_,data_stage_5__7786_,
  data_stage_5__7785_,data_stage_5__7784_,data_stage_5__7783_,data_stage_5__7782_,
  data_stage_5__7781_,data_stage_5__7780_,data_stage_5__7779_,data_stage_5__7778_,
  data_stage_5__7777_,data_stage_5__7776_,data_stage_5__7775_,data_stage_5__7774_,
  data_stage_5__7773_,data_stage_5__7772_,data_stage_5__7771_,data_stage_5__7770_,
  data_stage_5__7769_,data_stage_5__7768_,data_stage_5__7767_,data_stage_5__7766_,
  data_stage_5__7765_,data_stage_5__7764_,data_stage_5__7763_,data_stage_5__7762_,
  data_stage_5__7761_,data_stage_5__7760_,data_stage_5__7759_,data_stage_5__7758_,
  data_stage_5__7757_,data_stage_5__7756_,data_stage_5__7755_,data_stage_5__7754_,
  data_stage_5__7753_,data_stage_5__7752_,data_stage_5__7751_,data_stage_5__7750_,
  data_stage_5__7749_,data_stage_5__7748_,data_stage_5__7747_,data_stage_5__7746_,
  data_stage_5__7745_,data_stage_5__7744_,data_stage_5__7743_,data_stage_5__7742_,
  data_stage_5__7741_,data_stage_5__7740_,data_stage_5__7739_,data_stage_5__7738_,
  data_stage_5__7737_,data_stage_5__7736_,data_stage_5__7735_,data_stage_5__7734_,
  data_stage_5__7733_,data_stage_5__7732_,data_stage_5__7731_,data_stage_5__7730_,
  data_stage_5__7729_,data_stage_5__7728_,data_stage_5__7727_,data_stage_5__7726_,
  data_stage_5__7725_,data_stage_5__7724_,data_stage_5__7723_,data_stage_5__7722_,
  data_stage_5__7721_,data_stage_5__7720_,data_stage_5__7719_,data_stage_5__7718_,
  data_stage_5__7717_,data_stage_5__7716_,data_stage_5__7715_,data_stage_5__7714_,
  data_stage_5__7713_,data_stage_5__7712_,data_stage_5__7711_,data_stage_5__7710_,
  data_stage_5__7709_,data_stage_5__7708_,data_stage_5__7707_,data_stage_5__7706_,
  data_stage_5__7705_,data_stage_5__7704_,data_stage_5__7703_,data_stage_5__7702_,
  data_stage_5__7701_,data_stage_5__7700_,data_stage_5__7699_,data_stage_5__7698_,
  data_stage_5__7697_,data_stage_5__7696_,data_stage_5__7695_,data_stage_5__7694_,
  data_stage_5__7693_,data_stage_5__7692_,data_stage_5__7691_,data_stage_5__7690_,
  data_stage_5__7689_,data_stage_5__7688_,data_stage_5__7687_,data_stage_5__7686_,
  data_stage_5__7685_,data_stage_5__7684_,data_stage_5__7683_,data_stage_5__7682_,
  data_stage_5__7681_,data_stage_5__7680_,data_stage_5__7679_,data_stage_5__7678_,
  data_stage_5__7677_,data_stage_5__7676_,data_stage_5__7675_,data_stage_5__7674_,
  data_stage_5__7673_,data_stage_5__7672_,data_stage_5__7671_,data_stage_5__7670_,
  data_stage_5__7669_,data_stage_5__7668_,data_stage_5__7667_,data_stage_5__7666_,
  data_stage_5__7665_,data_stage_5__7664_,data_stage_5__7663_,data_stage_5__7662_,
  data_stage_5__7661_,data_stage_5__7660_,data_stage_5__7659_,data_stage_5__7658_,
  data_stage_5__7657_,data_stage_5__7656_,data_stage_5__7655_,data_stage_5__7654_,
  data_stage_5__7653_,data_stage_5__7652_,data_stage_5__7651_,data_stage_5__7650_,
  data_stage_5__7649_,data_stage_5__7648_,data_stage_5__7647_,data_stage_5__7646_,
  data_stage_5__7645_,data_stage_5__7644_,data_stage_5__7643_,data_stage_5__7642_,
  data_stage_5__7641_,data_stage_5__7640_,data_stage_5__7639_,data_stage_5__7638_,
  data_stage_5__7637_,data_stage_5__7636_,data_stage_5__7635_,data_stage_5__7634_,
  data_stage_5__7633_,data_stage_5__7632_,data_stage_5__7631_,data_stage_5__7630_,
  data_stage_5__7629_,data_stage_5__7628_,data_stage_5__7627_,data_stage_5__7626_,
  data_stage_5__7625_,data_stage_5__7624_,data_stage_5__7623_,data_stage_5__7622_,
  data_stage_5__7621_,data_stage_5__7620_,data_stage_5__7619_,data_stage_5__7618_,
  data_stage_5__7617_,data_stage_5__7616_,data_stage_5__7615_,data_stage_5__7614_,
  data_stage_5__7613_,data_stage_5__7612_,data_stage_5__7611_,data_stage_5__7610_,
  data_stage_5__7609_,data_stage_5__7608_,data_stage_5__7607_,data_stage_5__7606_,
  data_stage_5__7605_,data_stage_5__7604_,data_stage_5__7603_,data_stage_5__7602_,
  data_stage_5__7601_,data_stage_5__7600_,data_stage_5__7599_,data_stage_5__7598_,
  data_stage_5__7597_,data_stage_5__7596_,data_stage_5__7595_,data_stage_5__7594_,
  data_stage_5__7593_,data_stage_5__7592_,data_stage_5__7591_,data_stage_5__7590_,
  data_stage_5__7589_,data_stage_5__7588_,data_stage_5__7587_,data_stage_5__7586_,
  data_stage_5__7585_,data_stage_5__7584_,data_stage_5__7583_,data_stage_5__7582_,
  data_stage_5__7581_,data_stage_5__7580_,data_stage_5__7579_,data_stage_5__7578_,
  data_stage_5__7577_,data_stage_5__7576_,data_stage_5__7575_,data_stage_5__7574_,
  data_stage_5__7573_,data_stage_5__7572_,data_stage_5__7571_,data_stage_5__7570_,
  data_stage_5__7569_,data_stage_5__7568_,data_stage_5__7567_,data_stage_5__7566_,
  data_stage_5__7565_,data_stage_5__7564_,data_stage_5__7563_,data_stage_5__7562_,
  data_stage_5__7561_,data_stage_5__7560_,data_stage_5__7559_,data_stage_5__7558_,
  data_stage_5__7557_,data_stage_5__7556_,data_stage_5__7555_,data_stage_5__7554_,
  data_stage_5__7553_,data_stage_5__7552_,data_stage_5__7551_,data_stage_5__7550_,
  data_stage_5__7549_,data_stage_5__7548_,data_stage_5__7547_,data_stage_5__7546_,
  data_stage_5__7545_,data_stage_5__7544_,data_stage_5__7543_,data_stage_5__7542_,
  data_stage_5__7541_,data_stage_5__7540_,data_stage_5__7539_,data_stage_5__7538_,
  data_stage_5__7537_,data_stage_5__7536_,data_stage_5__7535_,data_stage_5__7534_,
  data_stage_5__7533_,data_stage_5__7532_,data_stage_5__7531_,data_stage_5__7530_,
  data_stage_5__7529_,data_stage_5__7528_,data_stage_5__7527_,data_stage_5__7526_,
  data_stage_5__7525_,data_stage_5__7524_,data_stage_5__7523_,data_stage_5__7522_,
  data_stage_5__7521_,data_stage_5__7520_,data_stage_5__7519_,data_stage_5__7518_,
  data_stage_5__7517_,data_stage_5__7516_,data_stage_5__7515_,data_stage_5__7514_,
  data_stage_5__7513_,data_stage_5__7512_,data_stage_5__7511_,data_stage_5__7510_,
  data_stage_5__7509_,data_stage_5__7508_,data_stage_5__7507_,data_stage_5__7506_,
  data_stage_5__7505_,data_stage_5__7504_,data_stage_5__7503_,data_stage_5__7502_,
  data_stage_5__7501_,data_stage_5__7500_,data_stage_5__7499_,data_stage_5__7498_,
  data_stage_5__7497_,data_stage_5__7496_,data_stage_5__7495_,data_stage_5__7494_,
  data_stage_5__7493_,data_stage_5__7492_,data_stage_5__7491_,data_stage_5__7490_,
  data_stage_5__7489_,data_stage_5__7488_,data_stage_5__7487_,data_stage_5__7486_,
  data_stage_5__7485_,data_stage_5__7484_,data_stage_5__7483_,data_stage_5__7482_,
  data_stage_5__7481_,data_stage_5__7480_,data_stage_5__7479_,data_stage_5__7478_,
  data_stage_5__7477_,data_stage_5__7476_,data_stage_5__7475_,data_stage_5__7474_,
  data_stage_5__7473_,data_stage_5__7472_,data_stage_5__7471_,data_stage_5__7470_,
  data_stage_5__7469_,data_stage_5__7468_,data_stage_5__7467_,data_stage_5__7466_,
  data_stage_5__7465_,data_stage_5__7464_,data_stage_5__7463_,data_stage_5__7462_,
  data_stage_5__7461_,data_stage_5__7460_,data_stage_5__7459_,data_stage_5__7458_,
  data_stage_5__7457_,data_stage_5__7456_,data_stage_5__7455_,data_stage_5__7454_,
  data_stage_5__7453_,data_stage_5__7452_,data_stage_5__7451_,data_stage_5__7450_,
  data_stage_5__7449_,data_stage_5__7448_,data_stage_5__7447_,data_stage_5__7446_,
  data_stage_5__7445_,data_stage_5__7444_,data_stage_5__7443_,data_stage_5__7442_,
  data_stage_5__7441_,data_stage_5__7440_,data_stage_5__7439_,data_stage_5__7438_,
  data_stage_5__7437_,data_stage_5__7436_,data_stage_5__7435_,data_stage_5__7434_,
  data_stage_5__7433_,data_stage_5__7432_,data_stage_5__7431_,data_stage_5__7430_,
  data_stage_5__7429_,data_stage_5__7428_,data_stage_5__7427_,data_stage_5__7426_,
  data_stage_5__7425_,data_stage_5__7424_,data_stage_5__7423_,data_stage_5__7422_,
  data_stage_5__7421_,data_stage_5__7420_,data_stage_5__7419_,data_stage_5__7418_,
  data_stage_5__7417_,data_stage_5__7416_,data_stage_5__7415_,data_stage_5__7414_,
  data_stage_5__7413_,data_stage_5__7412_,data_stage_5__7411_,data_stage_5__7410_,
  data_stage_5__7409_,data_stage_5__7408_,data_stage_5__7407_,data_stage_5__7406_,
  data_stage_5__7405_,data_stage_5__7404_,data_stage_5__7403_,data_stage_5__7402_,
  data_stage_5__7401_,data_stage_5__7400_,data_stage_5__7399_,data_stage_5__7398_,
  data_stage_5__7397_,data_stage_5__7396_,data_stage_5__7395_,data_stage_5__7394_,
  data_stage_5__7393_,data_stage_5__7392_,data_stage_5__7391_,data_stage_5__7390_,
  data_stage_5__7389_,data_stage_5__7388_,data_stage_5__7387_,data_stage_5__7386_,
  data_stage_5__7385_,data_stage_5__7384_,data_stage_5__7383_,data_stage_5__7382_,
  data_stage_5__7381_,data_stage_5__7380_,data_stage_5__7379_,data_stage_5__7378_,
  data_stage_5__7377_,data_stage_5__7376_,data_stage_5__7375_,data_stage_5__7374_,
  data_stage_5__7373_,data_stage_5__7372_,data_stage_5__7371_,data_stage_5__7370_,
  data_stage_5__7369_,data_stage_5__7368_,data_stage_5__7367_,data_stage_5__7366_,
  data_stage_5__7365_,data_stage_5__7364_,data_stage_5__7363_,data_stage_5__7362_,
  data_stage_5__7361_,data_stage_5__7360_,data_stage_5__7359_,data_stage_5__7358_,
  data_stage_5__7357_,data_stage_5__7356_,data_stage_5__7355_,data_stage_5__7354_,
  data_stage_5__7353_,data_stage_5__7352_,data_stage_5__7351_,data_stage_5__7350_,
  data_stage_5__7349_,data_stage_5__7348_,data_stage_5__7347_,data_stage_5__7346_,
  data_stage_5__7345_,data_stage_5__7344_,data_stage_5__7343_,data_stage_5__7342_,
  data_stage_5__7341_,data_stage_5__7340_,data_stage_5__7339_,data_stage_5__7338_,
  data_stage_5__7337_,data_stage_5__7336_,data_stage_5__7335_,data_stage_5__7334_,
  data_stage_5__7333_,data_stage_5__7332_,data_stage_5__7331_,data_stage_5__7330_,
  data_stage_5__7329_,data_stage_5__7328_,data_stage_5__7327_,data_stage_5__7326_,
  data_stage_5__7325_,data_stage_5__7324_,data_stage_5__7323_,data_stage_5__7322_,
  data_stage_5__7321_,data_stage_5__7320_,data_stage_5__7319_,data_stage_5__7318_,
  data_stage_5__7317_,data_stage_5__7316_,data_stage_5__7315_,data_stage_5__7314_,
  data_stage_5__7313_,data_stage_5__7312_,data_stage_5__7311_,data_stage_5__7310_,
  data_stage_5__7309_,data_stage_5__7308_,data_stage_5__7307_,data_stage_5__7306_,
  data_stage_5__7305_,data_stage_5__7304_,data_stage_5__7303_,data_stage_5__7302_,
  data_stage_5__7301_,data_stage_5__7300_,data_stage_5__7299_,data_stage_5__7298_,
  data_stage_5__7297_,data_stage_5__7296_,data_stage_5__7295_,data_stage_5__7294_,
  data_stage_5__7293_,data_stage_5__7292_,data_stage_5__7291_,data_stage_5__7290_,
  data_stage_5__7289_,data_stage_5__7288_,data_stage_5__7287_,data_stage_5__7286_,
  data_stage_5__7285_,data_stage_5__7284_,data_stage_5__7283_,data_stage_5__7282_,
  data_stage_5__7281_,data_stage_5__7280_,data_stage_5__7279_,data_stage_5__7278_,
  data_stage_5__7277_,data_stage_5__7276_,data_stage_5__7275_,data_stage_5__7274_,
  data_stage_5__7273_,data_stage_5__7272_,data_stage_5__7271_,data_stage_5__7270_,
  data_stage_5__7269_,data_stage_5__7268_,data_stage_5__7267_,data_stage_5__7266_,
  data_stage_5__7265_,data_stage_5__7264_,data_stage_5__7263_,data_stage_5__7262_,
  data_stage_5__7261_,data_stage_5__7260_,data_stage_5__7259_,data_stage_5__7258_,
  data_stage_5__7257_,data_stage_5__7256_,data_stage_5__7255_,data_stage_5__7254_,
  data_stage_5__7253_,data_stage_5__7252_,data_stage_5__7251_,data_stage_5__7250_,
  data_stage_5__7249_,data_stage_5__7248_,data_stage_5__7247_,data_stage_5__7246_,
  data_stage_5__7245_,data_stage_5__7244_,data_stage_5__7243_,data_stage_5__7242_,
  data_stage_5__7241_,data_stage_5__7240_,data_stage_5__7239_,data_stage_5__7238_,
  data_stage_5__7237_,data_stage_5__7236_,data_stage_5__7235_,data_stage_5__7234_,
  data_stage_5__7233_,data_stage_5__7232_,data_stage_5__7231_,data_stage_5__7230_,
  data_stage_5__7229_,data_stage_5__7228_,data_stage_5__7227_,data_stage_5__7226_,
  data_stage_5__7225_,data_stage_5__7224_,data_stage_5__7223_,data_stage_5__7222_,
  data_stage_5__7221_,data_stage_5__7220_,data_stage_5__7219_,data_stage_5__7218_,
  data_stage_5__7217_,data_stage_5__7216_,data_stage_5__7215_,data_stage_5__7214_,
  data_stage_5__7213_,data_stage_5__7212_,data_stage_5__7211_,data_stage_5__7210_,
  data_stage_5__7209_,data_stage_5__7208_,data_stage_5__7207_,data_stage_5__7206_,
  data_stage_5__7205_,data_stage_5__7204_,data_stage_5__7203_,data_stage_5__7202_,
  data_stage_5__7201_,data_stage_5__7200_,data_stage_5__7199_,data_stage_5__7198_,
  data_stage_5__7197_,data_stage_5__7196_,data_stage_5__7195_,data_stage_5__7194_,
  data_stage_5__7193_,data_stage_5__7192_,data_stage_5__7191_,data_stage_5__7190_,
  data_stage_5__7189_,data_stage_5__7188_,data_stage_5__7187_,data_stage_5__7186_,
  data_stage_5__7185_,data_stage_5__7184_,data_stage_5__7183_,data_stage_5__7182_,
  data_stage_5__7181_,data_stage_5__7180_,data_stage_5__7179_,data_stage_5__7178_,
  data_stage_5__7177_,data_stage_5__7176_,data_stage_5__7175_,data_stage_5__7174_,
  data_stage_5__7173_,data_stage_5__7172_,data_stage_5__7171_,data_stage_5__7170_,
  data_stage_5__7169_,data_stage_5__7168_,data_stage_5__7167_,data_stage_5__7166_,
  data_stage_5__7165_,data_stage_5__7164_,data_stage_5__7163_,data_stage_5__7162_,
  data_stage_5__7161_,data_stage_5__7160_,data_stage_5__7159_,data_stage_5__7158_,
  data_stage_5__7157_,data_stage_5__7156_,data_stage_5__7155_,data_stage_5__7154_,
  data_stage_5__7153_,data_stage_5__7152_,data_stage_5__7151_,data_stage_5__7150_,
  data_stage_5__7149_,data_stage_5__7148_,data_stage_5__7147_,data_stage_5__7146_,
  data_stage_5__7145_,data_stage_5__7144_,data_stage_5__7143_,data_stage_5__7142_,
  data_stage_5__7141_,data_stage_5__7140_,data_stage_5__7139_,data_stage_5__7138_,
  data_stage_5__7137_,data_stage_5__7136_,data_stage_5__7135_,data_stage_5__7134_,
  data_stage_5__7133_,data_stage_5__7132_,data_stage_5__7131_,data_stage_5__7130_,
  data_stage_5__7129_,data_stage_5__7128_,data_stage_5__7127_,data_stage_5__7126_,
  data_stage_5__7125_,data_stage_5__7124_,data_stage_5__7123_,data_stage_5__7122_,
  data_stage_5__7121_,data_stage_5__7120_,data_stage_5__7119_,data_stage_5__7118_,
  data_stage_5__7117_,data_stage_5__7116_,data_stage_5__7115_,data_stage_5__7114_,
  data_stage_5__7113_,data_stage_5__7112_,data_stage_5__7111_,data_stage_5__7110_,
  data_stage_5__7109_,data_stage_5__7108_,data_stage_5__7107_,data_stage_5__7106_,
  data_stage_5__7105_,data_stage_5__7104_,data_stage_5__7103_,data_stage_5__7102_,
  data_stage_5__7101_,data_stage_5__7100_,data_stage_5__7099_,data_stage_5__7098_,
  data_stage_5__7097_,data_stage_5__7096_,data_stage_5__7095_,data_stage_5__7094_,
  data_stage_5__7093_,data_stage_5__7092_,data_stage_5__7091_,data_stage_5__7090_,
  data_stage_5__7089_,data_stage_5__7088_,data_stage_5__7087_,data_stage_5__7086_,
  data_stage_5__7085_,data_stage_5__7084_,data_stage_5__7083_,data_stage_5__7082_,
  data_stage_5__7081_,data_stage_5__7080_,data_stage_5__7079_,data_stage_5__7078_,
  data_stage_5__7077_,data_stage_5__7076_,data_stage_5__7075_,data_stage_5__7074_,
  data_stage_5__7073_,data_stage_5__7072_,data_stage_5__7071_,data_stage_5__7070_,
  data_stage_5__7069_,data_stage_5__7068_,data_stage_5__7067_,data_stage_5__7066_,
  data_stage_5__7065_,data_stage_5__7064_,data_stage_5__7063_,data_stage_5__7062_,
  data_stage_5__7061_,data_stage_5__7060_,data_stage_5__7059_,data_stage_5__7058_,
  data_stage_5__7057_,data_stage_5__7056_,data_stage_5__7055_,data_stage_5__7054_,
  data_stage_5__7053_,data_stage_5__7052_,data_stage_5__7051_,data_stage_5__7050_,
  data_stage_5__7049_,data_stage_5__7048_,data_stage_5__7047_,data_stage_5__7046_,
  data_stage_5__7045_,data_stage_5__7044_,data_stage_5__7043_,data_stage_5__7042_,
  data_stage_5__7041_,data_stage_5__7040_,data_stage_5__7039_,data_stage_5__7038_,
  data_stage_5__7037_,data_stage_5__7036_,data_stage_5__7035_,data_stage_5__7034_,
  data_stage_5__7033_,data_stage_5__7032_,data_stage_5__7031_,data_stage_5__7030_,
  data_stage_5__7029_,data_stage_5__7028_,data_stage_5__7027_,data_stage_5__7026_,
  data_stage_5__7025_,data_stage_5__7024_,data_stage_5__7023_,data_stage_5__7022_,
  data_stage_5__7021_,data_stage_5__7020_,data_stage_5__7019_,data_stage_5__7018_,
  data_stage_5__7017_,data_stage_5__7016_,data_stage_5__7015_,data_stage_5__7014_,
  data_stage_5__7013_,data_stage_5__7012_,data_stage_5__7011_,data_stage_5__7010_,
  data_stage_5__7009_,data_stage_5__7008_,data_stage_5__7007_,data_stage_5__7006_,
  data_stage_5__7005_,data_stage_5__7004_,data_stage_5__7003_,data_stage_5__7002_,
  data_stage_5__7001_,data_stage_5__7000_,data_stage_5__6999_,data_stage_5__6998_,
  data_stage_5__6997_,data_stage_5__6996_,data_stage_5__6995_,data_stage_5__6994_,
  data_stage_5__6993_,data_stage_5__6992_,data_stage_5__6991_,data_stage_5__6990_,
  data_stage_5__6989_,data_stage_5__6988_,data_stage_5__6987_,data_stage_5__6986_,
  data_stage_5__6985_,data_stage_5__6984_,data_stage_5__6983_,data_stage_5__6982_,
  data_stage_5__6981_,data_stage_5__6980_,data_stage_5__6979_,data_stage_5__6978_,
  data_stage_5__6977_,data_stage_5__6976_,data_stage_5__6975_,data_stage_5__6974_,
  data_stage_5__6973_,data_stage_5__6972_,data_stage_5__6971_,data_stage_5__6970_,
  data_stage_5__6969_,data_stage_5__6968_,data_stage_5__6967_,data_stage_5__6966_,
  data_stage_5__6965_,data_stage_5__6964_,data_stage_5__6963_,data_stage_5__6962_,
  data_stage_5__6961_,data_stage_5__6960_,data_stage_5__6959_,data_stage_5__6958_,
  data_stage_5__6957_,data_stage_5__6956_,data_stage_5__6955_,data_stage_5__6954_,
  data_stage_5__6953_,data_stage_5__6952_,data_stage_5__6951_,data_stage_5__6950_,
  data_stage_5__6949_,data_stage_5__6948_,data_stage_5__6947_,data_stage_5__6946_,
  data_stage_5__6945_,data_stage_5__6944_,data_stage_5__6943_,data_stage_5__6942_,
  data_stage_5__6941_,data_stage_5__6940_,data_stage_5__6939_,data_stage_5__6938_,
  data_stage_5__6937_,data_stage_5__6936_,data_stage_5__6935_,data_stage_5__6934_,
  data_stage_5__6933_,data_stage_5__6932_,data_stage_5__6931_,data_stage_5__6930_,
  data_stage_5__6929_,data_stage_5__6928_,data_stage_5__6927_,data_stage_5__6926_,
  data_stage_5__6925_,data_stage_5__6924_,data_stage_5__6923_,data_stage_5__6922_,
  data_stage_5__6921_,data_stage_5__6920_,data_stage_5__6919_,data_stage_5__6918_,
  data_stage_5__6917_,data_stage_5__6916_,data_stage_5__6915_,data_stage_5__6914_,
  data_stage_5__6913_,data_stage_5__6912_,data_stage_5__6911_,data_stage_5__6910_,
  data_stage_5__6909_,data_stage_5__6908_,data_stage_5__6907_,data_stage_5__6906_,
  data_stage_5__6905_,data_stage_5__6904_,data_stage_5__6903_,data_stage_5__6902_,
  data_stage_5__6901_,data_stage_5__6900_,data_stage_5__6899_,data_stage_5__6898_,
  data_stage_5__6897_,data_stage_5__6896_,data_stage_5__6895_,data_stage_5__6894_,
  data_stage_5__6893_,data_stage_5__6892_,data_stage_5__6891_,data_stage_5__6890_,
  data_stage_5__6889_,data_stage_5__6888_,data_stage_5__6887_,data_stage_5__6886_,
  data_stage_5__6885_,data_stage_5__6884_,data_stage_5__6883_,data_stage_5__6882_,
  data_stage_5__6881_,data_stage_5__6880_,data_stage_5__6879_,data_stage_5__6878_,
  data_stage_5__6877_,data_stage_5__6876_,data_stage_5__6875_,data_stage_5__6874_,
  data_stage_5__6873_,data_stage_5__6872_,data_stage_5__6871_,data_stage_5__6870_,
  data_stage_5__6869_,data_stage_5__6868_,data_stage_5__6867_,data_stage_5__6866_,
  data_stage_5__6865_,data_stage_5__6864_,data_stage_5__6863_,data_stage_5__6862_,
  data_stage_5__6861_,data_stage_5__6860_,data_stage_5__6859_,data_stage_5__6858_,
  data_stage_5__6857_,data_stage_5__6856_,data_stage_5__6855_,data_stage_5__6854_,
  data_stage_5__6853_,data_stage_5__6852_,data_stage_5__6851_,data_stage_5__6850_,
  data_stage_5__6849_,data_stage_5__6848_,data_stage_5__6847_,data_stage_5__6846_,
  data_stage_5__6845_,data_stage_5__6844_,data_stage_5__6843_,data_stage_5__6842_,
  data_stage_5__6841_,data_stage_5__6840_,data_stage_5__6839_,data_stage_5__6838_,
  data_stage_5__6837_,data_stage_5__6836_,data_stage_5__6835_,data_stage_5__6834_,
  data_stage_5__6833_,data_stage_5__6832_,data_stage_5__6831_,data_stage_5__6830_,
  data_stage_5__6829_,data_stage_5__6828_,data_stage_5__6827_,data_stage_5__6826_,
  data_stage_5__6825_,data_stage_5__6824_,data_stage_5__6823_,data_stage_5__6822_,
  data_stage_5__6821_,data_stage_5__6820_,data_stage_5__6819_,data_stage_5__6818_,
  data_stage_5__6817_,data_stage_5__6816_,data_stage_5__6815_,data_stage_5__6814_,
  data_stage_5__6813_,data_stage_5__6812_,data_stage_5__6811_,data_stage_5__6810_,
  data_stage_5__6809_,data_stage_5__6808_,data_stage_5__6807_,data_stage_5__6806_,
  data_stage_5__6805_,data_stage_5__6804_,data_stage_5__6803_,data_stage_5__6802_,
  data_stage_5__6801_,data_stage_5__6800_,data_stage_5__6799_,data_stage_5__6798_,
  data_stage_5__6797_,data_stage_5__6796_,data_stage_5__6795_,data_stage_5__6794_,
  data_stage_5__6793_,data_stage_5__6792_,data_stage_5__6791_,data_stage_5__6790_,
  data_stage_5__6789_,data_stage_5__6788_,data_stage_5__6787_,data_stage_5__6786_,
  data_stage_5__6785_,data_stage_5__6784_,data_stage_5__6783_,data_stage_5__6782_,
  data_stage_5__6781_,data_stage_5__6780_,data_stage_5__6779_,data_stage_5__6778_,
  data_stage_5__6777_,data_stage_5__6776_,data_stage_5__6775_,data_stage_5__6774_,
  data_stage_5__6773_,data_stage_5__6772_,data_stage_5__6771_,data_stage_5__6770_,
  data_stage_5__6769_,data_stage_5__6768_,data_stage_5__6767_,data_stage_5__6766_,
  data_stage_5__6765_,data_stage_5__6764_,data_stage_5__6763_,data_stage_5__6762_,
  data_stage_5__6761_,data_stage_5__6760_,data_stage_5__6759_,data_stage_5__6758_,
  data_stage_5__6757_,data_stage_5__6756_,data_stage_5__6755_,data_stage_5__6754_,
  data_stage_5__6753_,data_stage_5__6752_,data_stage_5__6751_,data_stage_5__6750_,
  data_stage_5__6749_,data_stage_5__6748_,data_stage_5__6747_,data_stage_5__6746_,
  data_stage_5__6745_,data_stage_5__6744_,data_stage_5__6743_,data_stage_5__6742_,
  data_stage_5__6741_,data_stage_5__6740_,data_stage_5__6739_,data_stage_5__6738_,
  data_stage_5__6737_,data_stage_5__6736_,data_stage_5__6735_,data_stage_5__6734_,
  data_stage_5__6733_,data_stage_5__6732_,data_stage_5__6731_,data_stage_5__6730_,
  data_stage_5__6729_,data_stage_5__6728_,data_stage_5__6727_,data_stage_5__6726_,
  data_stage_5__6725_,data_stage_5__6724_,data_stage_5__6723_,data_stage_5__6722_,
  data_stage_5__6721_,data_stage_5__6720_,data_stage_5__6719_,data_stage_5__6718_,
  data_stage_5__6717_,data_stage_5__6716_,data_stage_5__6715_,data_stage_5__6714_,
  data_stage_5__6713_,data_stage_5__6712_,data_stage_5__6711_,data_stage_5__6710_,
  data_stage_5__6709_,data_stage_5__6708_,data_stage_5__6707_,data_stage_5__6706_,
  data_stage_5__6705_,data_stage_5__6704_,data_stage_5__6703_,data_stage_5__6702_,
  data_stage_5__6701_,data_stage_5__6700_,data_stage_5__6699_,data_stage_5__6698_,
  data_stage_5__6697_,data_stage_5__6696_,data_stage_5__6695_,data_stage_5__6694_,
  data_stage_5__6693_,data_stage_5__6692_,data_stage_5__6691_,data_stage_5__6690_,
  data_stage_5__6689_,data_stage_5__6688_,data_stage_5__6687_,data_stage_5__6686_,
  data_stage_5__6685_,data_stage_5__6684_,data_stage_5__6683_,data_stage_5__6682_,
  data_stage_5__6681_,data_stage_5__6680_,data_stage_5__6679_,data_stage_5__6678_,
  data_stage_5__6677_,data_stage_5__6676_,data_stage_5__6675_,data_stage_5__6674_,
  data_stage_5__6673_,data_stage_5__6672_,data_stage_5__6671_,data_stage_5__6670_,
  data_stage_5__6669_,data_stage_5__6668_,data_stage_5__6667_,data_stage_5__6666_,
  data_stage_5__6665_,data_stage_5__6664_,data_stage_5__6663_,data_stage_5__6662_,
  data_stage_5__6661_,data_stage_5__6660_,data_stage_5__6659_,data_stage_5__6658_,
  data_stage_5__6657_,data_stage_5__6656_,data_stage_5__6655_,data_stage_5__6654_,
  data_stage_5__6653_,data_stage_5__6652_,data_stage_5__6651_,data_stage_5__6650_,
  data_stage_5__6649_,data_stage_5__6648_,data_stage_5__6647_,data_stage_5__6646_,
  data_stage_5__6645_,data_stage_5__6644_,data_stage_5__6643_,data_stage_5__6642_,
  data_stage_5__6641_,data_stage_5__6640_,data_stage_5__6639_,data_stage_5__6638_,
  data_stage_5__6637_,data_stage_5__6636_,data_stage_5__6635_,data_stage_5__6634_,
  data_stage_5__6633_,data_stage_5__6632_,data_stage_5__6631_,data_stage_5__6630_,
  data_stage_5__6629_,data_stage_5__6628_,data_stage_5__6627_,data_stage_5__6626_,
  data_stage_5__6625_,data_stage_5__6624_,data_stage_5__6623_,data_stage_5__6622_,
  data_stage_5__6621_,data_stage_5__6620_,data_stage_5__6619_,data_stage_5__6618_,
  data_stage_5__6617_,data_stage_5__6616_,data_stage_5__6615_,data_stage_5__6614_,
  data_stage_5__6613_,data_stage_5__6612_,data_stage_5__6611_,data_stage_5__6610_,
  data_stage_5__6609_,data_stage_5__6608_,data_stage_5__6607_,data_stage_5__6606_,
  data_stage_5__6605_,data_stage_5__6604_,data_stage_5__6603_,data_stage_5__6602_,
  data_stage_5__6601_,data_stage_5__6600_,data_stage_5__6599_,data_stage_5__6598_,
  data_stage_5__6597_,data_stage_5__6596_,data_stage_5__6595_,data_stage_5__6594_,
  data_stage_5__6593_,data_stage_5__6592_,data_stage_5__6591_,data_stage_5__6590_,
  data_stage_5__6589_,data_stage_5__6588_,data_stage_5__6587_,data_stage_5__6586_,
  data_stage_5__6585_,data_stage_5__6584_,data_stage_5__6583_,data_stage_5__6582_,
  data_stage_5__6581_,data_stage_5__6580_,data_stage_5__6579_,data_stage_5__6578_,
  data_stage_5__6577_,data_stage_5__6576_,data_stage_5__6575_,data_stage_5__6574_,
  data_stage_5__6573_,data_stage_5__6572_,data_stage_5__6571_,data_stage_5__6570_,
  data_stage_5__6569_,data_stage_5__6568_,data_stage_5__6567_,data_stage_5__6566_,
  data_stage_5__6565_,data_stage_5__6564_,data_stage_5__6563_,data_stage_5__6562_,
  data_stage_5__6561_,data_stage_5__6560_,data_stage_5__6559_,data_stage_5__6558_,
  data_stage_5__6557_,data_stage_5__6556_,data_stage_5__6555_,data_stage_5__6554_,
  data_stage_5__6553_,data_stage_5__6552_,data_stage_5__6551_,data_stage_5__6550_,
  data_stage_5__6549_,data_stage_5__6548_,data_stage_5__6547_,data_stage_5__6546_,
  data_stage_5__6545_,data_stage_5__6544_,data_stage_5__6543_,data_stage_5__6542_,
  data_stage_5__6541_,data_stage_5__6540_,data_stage_5__6539_,data_stage_5__6538_,
  data_stage_5__6537_,data_stage_5__6536_,data_stage_5__6535_,data_stage_5__6534_,
  data_stage_5__6533_,data_stage_5__6532_,data_stage_5__6531_,data_stage_5__6530_,
  data_stage_5__6529_,data_stage_5__6528_,data_stage_5__6527_,data_stage_5__6526_,
  data_stage_5__6525_,data_stage_5__6524_,data_stage_5__6523_,data_stage_5__6522_,
  data_stage_5__6521_,data_stage_5__6520_,data_stage_5__6519_,data_stage_5__6518_,
  data_stage_5__6517_,data_stage_5__6516_,data_stage_5__6515_,data_stage_5__6514_,
  data_stage_5__6513_,data_stage_5__6512_,data_stage_5__6511_,data_stage_5__6510_,
  data_stage_5__6509_,data_stage_5__6508_,data_stage_5__6507_,data_stage_5__6506_,
  data_stage_5__6505_,data_stage_5__6504_,data_stage_5__6503_,data_stage_5__6502_,
  data_stage_5__6501_,data_stage_5__6500_,data_stage_5__6499_,data_stage_5__6498_,
  data_stage_5__6497_,data_stage_5__6496_,data_stage_5__6495_,data_stage_5__6494_,
  data_stage_5__6493_,data_stage_5__6492_,data_stage_5__6491_,data_stage_5__6490_,
  data_stage_5__6489_,data_stage_5__6488_,data_stage_5__6487_,data_stage_5__6486_,
  data_stage_5__6485_,data_stage_5__6484_,data_stage_5__6483_,data_stage_5__6482_,
  data_stage_5__6481_,data_stage_5__6480_,data_stage_5__6479_,data_stage_5__6478_,
  data_stage_5__6477_,data_stage_5__6476_,data_stage_5__6475_,data_stage_5__6474_,
  data_stage_5__6473_,data_stage_5__6472_,data_stage_5__6471_,data_stage_5__6470_,
  data_stage_5__6469_,data_stage_5__6468_,data_stage_5__6467_,data_stage_5__6466_,
  data_stage_5__6465_,data_stage_5__6464_,data_stage_5__6463_,data_stage_5__6462_,
  data_stage_5__6461_,data_stage_5__6460_,data_stage_5__6459_,data_stage_5__6458_,
  data_stage_5__6457_,data_stage_5__6456_,data_stage_5__6455_,data_stage_5__6454_,
  data_stage_5__6453_,data_stage_5__6452_,data_stage_5__6451_,data_stage_5__6450_,
  data_stage_5__6449_,data_stage_5__6448_,data_stage_5__6447_,data_stage_5__6446_,
  data_stage_5__6445_,data_stage_5__6444_,data_stage_5__6443_,data_stage_5__6442_,
  data_stage_5__6441_,data_stage_5__6440_,data_stage_5__6439_,data_stage_5__6438_,
  data_stage_5__6437_,data_stage_5__6436_,data_stage_5__6435_,data_stage_5__6434_,
  data_stage_5__6433_,data_stage_5__6432_,data_stage_5__6431_,data_stage_5__6430_,
  data_stage_5__6429_,data_stage_5__6428_,data_stage_5__6427_,data_stage_5__6426_,
  data_stage_5__6425_,data_stage_5__6424_,data_stage_5__6423_,data_stage_5__6422_,
  data_stage_5__6421_,data_stage_5__6420_,data_stage_5__6419_,data_stage_5__6418_,
  data_stage_5__6417_,data_stage_5__6416_,data_stage_5__6415_,data_stage_5__6414_,
  data_stage_5__6413_,data_stage_5__6412_,data_stage_5__6411_,data_stage_5__6410_,
  data_stage_5__6409_,data_stage_5__6408_,data_stage_5__6407_,data_stage_5__6406_,
  data_stage_5__6405_,data_stage_5__6404_,data_stage_5__6403_,data_stage_5__6402_,
  data_stage_5__6401_,data_stage_5__6400_,data_stage_5__6399_,data_stage_5__6398_,
  data_stage_5__6397_,data_stage_5__6396_,data_stage_5__6395_,data_stage_5__6394_,
  data_stage_5__6393_,data_stage_5__6392_,data_stage_5__6391_,data_stage_5__6390_,
  data_stage_5__6389_,data_stage_5__6388_,data_stage_5__6387_,data_stage_5__6386_,
  data_stage_5__6385_,data_stage_5__6384_,data_stage_5__6383_,data_stage_5__6382_,
  data_stage_5__6381_,data_stage_5__6380_,data_stage_5__6379_,data_stage_5__6378_,
  data_stage_5__6377_,data_stage_5__6376_,data_stage_5__6375_,data_stage_5__6374_,
  data_stage_5__6373_,data_stage_5__6372_,data_stage_5__6371_,data_stage_5__6370_,
  data_stage_5__6369_,data_stage_5__6368_,data_stage_5__6367_,data_stage_5__6366_,
  data_stage_5__6365_,data_stage_5__6364_,data_stage_5__6363_,data_stage_5__6362_,
  data_stage_5__6361_,data_stage_5__6360_,data_stage_5__6359_,data_stage_5__6358_,
  data_stage_5__6357_,data_stage_5__6356_,data_stage_5__6355_,data_stage_5__6354_,
  data_stage_5__6353_,data_stage_5__6352_,data_stage_5__6351_,data_stage_5__6350_,
  data_stage_5__6349_,data_stage_5__6348_,data_stage_5__6347_,data_stage_5__6346_,
  data_stage_5__6345_,data_stage_5__6344_,data_stage_5__6343_,data_stage_5__6342_,
  data_stage_5__6341_,data_stage_5__6340_,data_stage_5__6339_,data_stage_5__6338_,
  data_stage_5__6337_,data_stage_5__6336_,data_stage_5__6335_,data_stage_5__6334_,
  data_stage_5__6333_,data_stage_5__6332_,data_stage_5__6331_,data_stage_5__6330_,
  data_stage_5__6329_,data_stage_5__6328_,data_stage_5__6327_,data_stage_5__6326_,
  data_stage_5__6325_,data_stage_5__6324_,data_stage_5__6323_,data_stage_5__6322_,
  data_stage_5__6321_,data_stage_5__6320_,data_stage_5__6319_,data_stage_5__6318_,
  data_stage_5__6317_,data_stage_5__6316_,data_stage_5__6315_,data_stage_5__6314_,
  data_stage_5__6313_,data_stage_5__6312_,data_stage_5__6311_,data_stage_5__6310_,
  data_stage_5__6309_,data_stage_5__6308_,data_stage_5__6307_,data_stage_5__6306_,
  data_stage_5__6305_,data_stage_5__6304_,data_stage_5__6303_,data_stage_5__6302_,
  data_stage_5__6301_,data_stage_5__6300_,data_stage_5__6299_,data_stage_5__6298_,
  data_stage_5__6297_,data_stage_5__6296_,data_stage_5__6295_,data_stage_5__6294_,
  data_stage_5__6293_,data_stage_5__6292_,data_stage_5__6291_,data_stage_5__6290_,
  data_stage_5__6289_,data_stage_5__6288_,data_stage_5__6287_,data_stage_5__6286_,
  data_stage_5__6285_,data_stage_5__6284_,data_stage_5__6283_,data_stage_5__6282_,
  data_stage_5__6281_,data_stage_5__6280_,data_stage_5__6279_,data_stage_5__6278_,
  data_stage_5__6277_,data_stage_5__6276_,data_stage_5__6275_,data_stage_5__6274_,
  data_stage_5__6273_,data_stage_5__6272_,data_stage_5__6271_,data_stage_5__6270_,
  data_stage_5__6269_,data_stage_5__6268_,data_stage_5__6267_,data_stage_5__6266_,
  data_stage_5__6265_,data_stage_5__6264_,data_stage_5__6263_,data_stage_5__6262_,
  data_stage_5__6261_,data_stage_5__6260_,data_stage_5__6259_,data_stage_5__6258_,
  data_stage_5__6257_,data_stage_5__6256_,data_stage_5__6255_,data_stage_5__6254_,
  data_stage_5__6253_,data_stage_5__6252_,data_stage_5__6251_,data_stage_5__6250_,
  data_stage_5__6249_,data_stage_5__6248_,data_stage_5__6247_,data_stage_5__6246_,
  data_stage_5__6245_,data_stage_5__6244_,data_stage_5__6243_,data_stage_5__6242_,
  data_stage_5__6241_,data_stage_5__6240_,data_stage_5__6239_,data_stage_5__6238_,
  data_stage_5__6237_,data_stage_5__6236_,data_stage_5__6235_,data_stage_5__6234_,
  data_stage_5__6233_,data_stage_5__6232_,data_stage_5__6231_,data_stage_5__6230_,
  data_stage_5__6229_,data_stage_5__6228_,data_stage_5__6227_,data_stage_5__6226_,
  data_stage_5__6225_,data_stage_5__6224_,data_stage_5__6223_,data_stage_5__6222_,
  data_stage_5__6221_,data_stage_5__6220_,data_stage_5__6219_,data_stage_5__6218_,
  data_stage_5__6217_,data_stage_5__6216_,data_stage_5__6215_,data_stage_5__6214_,
  data_stage_5__6213_,data_stage_5__6212_,data_stage_5__6211_,data_stage_5__6210_,
  data_stage_5__6209_,data_stage_5__6208_,data_stage_5__6207_,data_stage_5__6206_,
  data_stage_5__6205_,data_stage_5__6204_,data_stage_5__6203_,data_stage_5__6202_,
  data_stage_5__6201_,data_stage_5__6200_,data_stage_5__6199_,data_stage_5__6198_,
  data_stage_5__6197_,data_stage_5__6196_,data_stage_5__6195_,data_stage_5__6194_,
  data_stage_5__6193_,data_stage_5__6192_,data_stage_5__6191_,data_stage_5__6190_,
  data_stage_5__6189_,data_stage_5__6188_,data_stage_5__6187_,data_stage_5__6186_,
  data_stage_5__6185_,data_stage_5__6184_,data_stage_5__6183_,data_stage_5__6182_,
  data_stage_5__6181_,data_stage_5__6180_,data_stage_5__6179_,data_stage_5__6178_,
  data_stage_5__6177_,data_stage_5__6176_,data_stage_5__6175_,data_stage_5__6174_,
  data_stage_5__6173_,data_stage_5__6172_,data_stage_5__6171_,data_stage_5__6170_,
  data_stage_5__6169_,data_stage_5__6168_,data_stage_5__6167_,data_stage_5__6166_,
  data_stage_5__6165_,data_stage_5__6164_,data_stage_5__6163_,data_stage_5__6162_,
  data_stage_5__6161_,data_stage_5__6160_,data_stage_5__6159_,data_stage_5__6158_,
  data_stage_5__6157_,data_stage_5__6156_,data_stage_5__6155_,data_stage_5__6154_,
  data_stage_5__6153_,data_stage_5__6152_,data_stage_5__6151_,data_stage_5__6150_,
  data_stage_5__6149_,data_stage_5__6148_,data_stage_5__6147_,data_stage_5__6146_,
  data_stage_5__6145_,data_stage_5__6144_,data_stage_5__6143_,data_stage_5__6142_,
  data_stage_5__6141_,data_stage_5__6140_,data_stage_5__6139_,data_stage_5__6138_,
  data_stage_5__6137_,data_stage_5__6136_,data_stage_5__6135_,data_stage_5__6134_,
  data_stage_5__6133_,data_stage_5__6132_,data_stage_5__6131_,data_stage_5__6130_,
  data_stage_5__6129_,data_stage_5__6128_,data_stage_5__6127_,data_stage_5__6126_,
  data_stage_5__6125_,data_stage_5__6124_,data_stage_5__6123_,data_stage_5__6122_,
  data_stage_5__6121_,data_stage_5__6120_,data_stage_5__6119_,data_stage_5__6118_,
  data_stage_5__6117_,data_stage_5__6116_,data_stage_5__6115_,data_stage_5__6114_,
  data_stage_5__6113_,data_stage_5__6112_,data_stage_5__6111_,data_stage_5__6110_,
  data_stage_5__6109_,data_stage_5__6108_,data_stage_5__6107_,data_stage_5__6106_,
  data_stage_5__6105_,data_stage_5__6104_,data_stage_5__6103_,data_stage_5__6102_,
  data_stage_5__6101_,data_stage_5__6100_,data_stage_5__6099_,data_stage_5__6098_,
  data_stage_5__6097_,data_stage_5__6096_,data_stage_5__6095_,data_stage_5__6094_,
  data_stage_5__6093_,data_stage_5__6092_,data_stage_5__6091_,data_stage_5__6090_,
  data_stage_5__6089_,data_stage_5__6088_,data_stage_5__6087_,data_stage_5__6086_,
  data_stage_5__6085_,data_stage_5__6084_,data_stage_5__6083_,data_stage_5__6082_,
  data_stage_5__6081_,data_stage_5__6080_,data_stage_5__6079_,data_stage_5__6078_,
  data_stage_5__6077_,data_stage_5__6076_,data_stage_5__6075_,data_stage_5__6074_,
  data_stage_5__6073_,data_stage_5__6072_,data_stage_5__6071_,data_stage_5__6070_,
  data_stage_5__6069_,data_stage_5__6068_,data_stage_5__6067_,data_stage_5__6066_,
  data_stage_5__6065_,data_stage_5__6064_,data_stage_5__6063_,data_stage_5__6062_,
  data_stage_5__6061_,data_stage_5__6060_,data_stage_5__6059_,data_stage_5__6058_,
  data_stage_5__6057_,data_stage_5__6056_,data_stage_5__6055_,data_stage_5__6054_,
  data_stage_5__6053_,data_stage_5__6052_,data_stage_5__6051_,data_stage_5__6050_,
  data_stage_5__6049_,data_stage_5__6048_,data_stage_5__6047_,data_stage_5__6046_,
  data_stage_5__6045_,data_stage_5__6044_,data_stage_5__6043_,data_stage_5__6042_,
  data_stage_5__6041_,data_stage_5__6040_,data_stage_5__6039_,data_stage_5__6038_,
  data_stage_5__6037_,data_stage_5__6036_,data_stage_5__6035_,data_stage_5__6034_,
  data_stage_5__6033_,data_stage_5__6032_,data_stage_5__6031_,data_stage_5__6030_,
  data_stage_5__6029_,data_stage_5__6028_,data_stage_5__6027_,data_stage_5__6026_,
  data_stage_5__6025_,data_stage_5__6024_,data_stage_5__6023_,data_stage_5__6022_,
  data_stage_5__6021_,data_stage_5__6020_,data_stage_5__6019_,data_stage_5__6018_,
  data_stage_5__6017_,data_stage_5__6016_,data_stage_5__6015_,data_stage_5__6014_,
  data_stage_5__6013_,data_stage_5__6012_,data_stage_5__6011_,data_stage_5__6010_,
  data_stage_5__6009_,data_stage_5__6008_,data_stage_5__6007_,data_stage_5__6006_,
  data_stage_5__6005_,data_stage_5__6004_,data_stage_5__6003_,data_stage_5__6002_,
  data_stage_5__6001_,data_stage_5__6000_,data_stage_5__5999_,data_stage_5__5998_,
  data_stage_5__5997_,data_stage_5__5996_,data_stage_5__5995_,data_stage_5__5994_,
  data_stage_5__5993_,data_stage_5__5992_,data_stage_5__5991_,data_stage_5__5990_,
  data_stage_5__5989_,data_stage_5__5988_,data_stage_5__5987_,data_stage_5__5986_,
  data_stage_5__5985_,data_stage_5__5984_,data_stage_5__5983_,data_stage_5__5982_,
  data_stage_5__5981_,data_stage_5__5980_,data_stage_5__5979_,data_stage_5__5978_,
  data_stage_5__5977_,data_stage_5__5976_,data_stage_5__5975_,data_stage_5__5974_,
  data_stage_5__5973_,data_stage_5__5972_,data_stage_5__5971_,data_stage_5__5970_,
  data_stage_5__5969_,data_stage_5__5968_,data_stage_5__5967_,data_stage_5__5966_,
  data_stage_5__5965_,data_stage_5__5964_,data_stage_5__5963_,data_stage_5__5962_,
  data_stage_5__5961_,data_stage_5__5960_,data_stage_5__5959_,data_stage_5__5958_,
  data_stage_5__5957_,data_stage_5__5956_,data_stage_5__5955_,data_stage_5__5954_,
  data_stage_5__5953_,data_stage_5__5952_,data_stage_5__5951_,data_stage_5__5950_,
  data_stage_5__5949_,data_stage_5__5948_,data_stage_5__5947_,data_stage_5__5946_,
  data_stage_5__5945_,data_stage_5__5944_,data_stage_5__5943_,data_stage_5__5942_,
  data_stage_5__5941_,data_stage_5__5940_,data_stage_5__5939_,data_stage_5__5938_,
  data_stage_5__5937_,data_stage_5__5936_,data_stage_5__5935_,data_stage_5__5934_,
  data_stage_5__5933_,data_stage_5__5932_,data_stage_5__5931_,data_stage_5__5930_,
  data_stage_5__5929_,data_stage_5__5928_,data_stage_5__5927_,data_stage_5__5926_,
  data_stage_5__5925_,data_stage_5__5924_,data_stage_5__5923_,data_stage_5__5922_,
  data_stage_5__5921_,data_stage_5__5920_,data_stage_5__5919_,data_stage_5__5918_,
  data_stage_5__5917_,data_stage_5__5916_,data_stage_5__5915_,data_stage_5__5914_,
  data_stage_5__5913_,data_stage_5__5912_,data_stage_5__5911_,data_stage_5__5910_,
  data_stage_5__5909_,data_stage_5__5908_,data_stage_5__5907_,data_stage_5__5906_,
  data_stage_5__5905_,data_stage_5__5904_,data_stage_5__5903_,data_stage_5__5902_,
  data_stage_5__5901_,data_stage_5__5900_,data_stage_5__5899_,data_stage_5__5898_,
  data_stage_5__5897_,data_stage_5__5896_,data_stage_5__5895_,data_stage_5__5894_,
  data_stage_5__5893_,data_stage_5__5892_,data_stage_5__5891_,data_stage_5__5890_,
  data_stage_5__5889_,data_stage_5__5888_,data_stage_5__5887_,data_stage_5__5886_,
  data_stage_5__5885_,data_stage_5__5884_,data_stage_5__5883_,data_stage_5__5882_,
  data_stage_5__5881_,data_stage_5__5880_,data_stage_5__5879_,data_stage_5__5878_,
  data_stage_5__5877_,data_stage_5__5876_,data_stage_5__5875_,data_stage_5__5874_,
  data_stage_5__5873_,data_stage_5__5872_,data_stage_5__5871_,data_stage_5__5870_,
  data_stage_5__5869_,data_stage_5__5868_,data_stage_5__5867_,data_stage_5__5866_,
  data_stage_5__5865_,data_stage_5__5864_,data_stage_5__5863_,data_stage_5__5862_,
  data_stage_5__5861_,data_stage_5__5860_,data_stage_5__5859_,data_stage_5__5858_,
  data_stage_5__5857_,data_stage_5__5856_,data_stage_5__5855_,data_stage_5__5854_,
  data_stage_5__5853_,data_stage_5__5852_,data_stage_5__5851_,data_stage_5__5850_,
  data_stage_5__5849_,data_stage_5__5848_,data_stage_5__5847_,data_stage_5__5846_,
  data_stage_5__5845_,data_stage_5__5844_,data_stage_5__5843_,data_stage_5__5842_,
  data_stage_5__5841_,data_stage_5__5840_,data_stage_5__5839_,data_stage_5__5838_,
  data_stage_5__5837_,data_stage_5__5836_,data_stage_5__5835_,data_stage_5__5834_,
  data_stage_5__5833_,data_stage_5__5832_,data_stage_5__5831_,data_stage_5__5830_,
  data_stage_5__5829_,data_stage_5__5828_,data_stage_5__5827_,data_stage_5__5826_,
  data_stage_5__5825_,data_stage_5__5824_,data_stage_5__5823_,data_stage_5__5822_,
  data_stage_5__5821_,data_stage_5__5820_,data_stage_5__5819_,data_stage_5__5818_,
  data_stage_5__5817_,data_stage_5__5816_,data_stage_5__5815_,data_stage_5__5814_,
  data_stage_5__5813_,data_stage_5__5812_,data_stage_5__5811_,data_stage_5__5810_,
  data_stage_5__5809_,data_stage_5__5808_,data_stage_5__5807_,data_stage_5__5806_,
  data_stage_5__5805_,data_stage_5__5804_,data_stage_5__5803_,data_stage_5__5802_,
  data_stage_5__5801_,data_stage_5__5800_,data_stage_5__5799_,data_stage_5__5798_,
  data_stage_5__5797_,data_stage_5__5796_,data_stage_5__5795_,data_stage_5__5794_,
  data_stage_5__5793_,data_stage_5__5792_,data_stage_5__5791_,data_stage_5__5790_,
  data_stage_5__5789_,data_stage_5__5788_,data_stage_5__5787_,data_stage_5__5786_,
  data_stage_5__5785_,data_stage_5__5784_,data_stage_5__5783_,data_stage_5__5782_,
  data_stage_5__5781_,data_stage_5__5780_,data_stage_5__5779_,data_stage_5__5778_,
  data_stage_5__5777_,data_stage_5__5776_,data_stage_5__5775_,data_stage_5__5774_,
  data_stage_5__5773_,data_stage_5__5772_,data_stage_5__5771_,data_stage_5__5770_,
  data_stage_5__5769_,data_stage_5__5768_,data_stage_5__5767_,data_stage_5__5766_,
  data_stage_5__5765_,data_stage_5__5764_,data_stage_5__5763_,data_stage_5__5762_,
  data_stage_5__5761_,data_stage_5__5760_,data_stage_5__5759_,data_stage_5__5758_,
  data_stage_5__5757_,data_stage_5__5756_,data_stage_5__5755_,data_stage_5__5754_,
  data_stage_5__5753_,data_stage_5__5752_,data_stage_5__5751_,data_stage_5__5750_,
  data_stage_5__5749_,data_stage_5__5748_,data_stage_5__5747_,data_stage_5__5746_,
  data_stage_5__5745_,data_stage_5__5744_,data_stage_5__5743_,data_stage_5__5742_,
  data_stage_5__5741_,data_stage_5__5740_,data_stage_5__5739_,data_stage_5__5738_,
  data_stage_5__5737_,data_stage_5__5736_,data_stage_5__5735_,data_stage_5__5734_,
  data_stage_5__5733_,data_stage_5__5732_,data_stage_5__5731_,data_stage_5__5730_,
  data_stage_5__5729_,data_stage_5__5728_,data_stage_5__5727_,data_stage_5__5726_,
  data_stage_5__5725_,data_stage_5__5724_,data_stage_5__5723_,data_stage_5__5722_,
  data_stage_5__5721_,data_stage_5__5720_,data_stage_5__5719_,data_stage_5__5718_,
  data_stage_5__5717_,data_stage_5__5716_,data_stage_5__5715_,data_stage_5__5714_,
  data_stage_5__5713_,data_stage_5__5712_,data_stage_5__5711_,data_stage_5__5710_,
  data_stage_5__5709_,data_stage_5__5708_,data_stage_5__5707_,data_stage_5__5706_,
  data_stage_5__5705_,data_stage_5__5704_,data_stage_5__5703_,data_stage_5__5702_,
  data_stage_5__5701_,data_stage_5__5700_,data_stage_5__5699_,data_stage_5__5698_,
  data_stage_5__5697_,data_stage_5__5696_,data_stage_5__5695_,data_stage_5__5694_,
  data_stage_5__5693_,data_stage_5__5692_,data_stage_5__5691_,data_stage_5__5690_,
  data_stage_5__5689_,data_stage_5__5688_,data_stage_5__5687_,data_stage_5__5686_,
  data_stage_5__5685_,data_stage_5__5684_,data_stage_5__5683_,data_stage_5__5682_,
  data_stage_5__5681_,data_stage_5__5680_,data_stage_5__5679_,data_stage_5__5678_,
  data_stage_5__5677_,data_stage_5__5676_,data_stage_5__5675_,data_stage_5__5674_,
  data_stage_5__5673_,data_stage_5__5672_,data_stage_5__5671_,data_stage_5__5670_,
  data_stage_5__5669_,data_stage_5__5668_,data_stage_5__5667_,data_stage_5__5666_,
  data_stage_5__5665_,data_stage_5__5664_,data_stage_5__5663_,data_stage_5__5662_,
  data_stage_5__5661_,data_stage_5__5660_,data_stage_5__5659_,data_stage_5__5658_,
  data_stage_5__5657_,data_stage_5__5656_,data_stage_5__5655_,data_stage_5__5654_,
  data_stage_5__5653_,data_stage_5__5652_,data_stage_5__5651_,data_stage_5__5650_,
  data_stage_5__5649_,data_stage_5__5648_,data_stage_5__5647_,data_stage_5__5646_,
  data_stage_5__5645_,data_stage_5__5644_,data_stage_5__5643_,data_stage_5__5642_,
  data_stage_5__5641_,data_stage_5__5640_,data_stage_5__5639_,data_stage_5__5638_,
  data_stage_5__5637_,data_stage_5__5636_,data_stage_5__5635_,data_stage_5__5634_,
  data_stage_5__5633_,data_stage_5__5632_,data_stage_5__5631_,data_stage_5__5630_,
  data_stage_5__5629_,data_stage_5__5628_,data_stage_5__5627_,data_stage_5__5626_,
  data_stage_5__5625_,data_stage_5__5624_,data_stage_5__5623_,data_stage_5__5622_,
  data_stage_5__5621_,data_stage_5__5620_,data_stage_5__5619_,data_stage_5__5618_,
  data_stage_5__5617_,data_stage_5__5616_,data_stage_5__5615_,data_stage_5__5614_,
  data_stage_5__5613_,data_stage_5__5612_,data_stage_5__5611_,data_stage_5__5610_,
  data_stage_5__5609_,data_stage_5__5608_,data_stage_5__5607_,data_stage_5__5606_,
  data_stage_5__5605_,data_stage_5__5604_,data_stage_5__5603_,data_stage_5__5602_,
  data_stage_5__5601_,data_stage_5__5600_,data_stage_5__5599_,data_stage_5__5598_,
  data_stage_5__5597_,data_stage_5__5596_,data_stage_5__5595_,data_stage_5__5594_,
  data_stage_5__5593_,data_stage_5__5592_,data_stage_5__5591_,data_stage_5__5590_,
  data_stage_5__5589_,data_stage_5__5588_,data_stage_5__5587_,data_stage_5__5586_,
  data_stage_5__5585_,data_stage_5__5584_,data_stage_5__5583_,data_stage_5__5582_,
  data_stage_5__5581_,data_stage_5__5580_,data_stage_5__5579_,data_stage_5__5578_,
  data_stage_5__5577_,data_stage_5__5576_,data_stage_5__5575_,data_stage_5__5574_,
  data_stage_5__5573_,data_stage_5__5572_,data_stage_5__5571_,data_stage_5__5570_,
  data_stage_5__5569_,data_stage_5__5568_,data_stage_5__5567_,data_stage_5__5566_,
  data_stage_5__5565_,data_stage_5__5564_,data_stage_5__5563_,data_stage_5__5562_,
  data_stage_5__5561_,data_stage_5__5560_,data_stage_5__5559_,data_stage_5__5558_,
  data_stage_5__5557_,data_stage_5__5556_,data_stage_5__5555_,data_stage_5__5554_,
  data_stage_5__5553_,data_stage_5__5552_,data_stage_5__5551_,data_stage_5__5550_,
  data_stage_5__5549_,data_stage_5__5548_,data_stage_5__5547_,data_stage_5__5546_,
  data_stage_5__5545_,data_stage_5__5544_,data_stage_5__5543_,data_stage_5__5542_,
  data_stage_5__5541_,data_stage_5__5540_,data_stage_5__5539_,data_stage_5__5538_,
  data_stage_5__5537_,data_stage_5__5536_,data_stage_5__5535_,data_stage_5__5534_,
  data_stage_5__5533_,data_stage_5__5532_,data_stage_5__5531_,data_stage_5__5530_,
  data_stage_5__5529_,data_stage_5__5528_,data_stage_5__5527_,data_stage_5__5526_,
  data_stage_5__5525_,data_stage_5__5524_,data_stage_5__5523_,data_stage_5__5522_,
  data_stage_5__5521_,data_stage_5__5520_,data_stage_5__5519_,data_stage_5__5518_,
  data_stage_5__5517_,data_stage_5__5516_,data_stage_5__5515_,data_stage_5__5514_,
  data_stage_5__5513_,data_stage_5__5512_,data_stage_5__5511_,data_stage_5__5510_,
  data_stage_5__5509_,data_stage_5__5508_,data_stage_5__5507_,data_stage_5__5506_,
  data_stage_5__5505_,data_stage_5__5504_,data_stage_5__5503_,data_stage_5__5502_,
  data_stage_5__5501_,data_stage_5__5500_,data_stage_5__5499_,data_stage_5__5498_,
  data_stage_5__5497_,data_stage_5__5496_,data_stage_5__5495_,data_stage_5__5494_,
  data_stage_5__5493_,data_stage_5__5492_,data_stage_5__5491_,data_stage_5__5490_,
  data_stage_5__5489_,data_stage_5__5488_,data_stage_5__5487_,data_stage_5__5486_,
  data_stage_5__5485_,data_stage_5__5484_,data_stage_5__5483_,data_stage_5__5482_,
  data_stage_5__5481_,data_stage_5__5480_,data_stage_5__5479_,data_stage_5__5478_,
  data_stage_5__5477_,data_stage_5__5476_,data_stage_5__5475_,data_stage_5__5474_,
  data_stage_5__5473_,data_stage_5__5472_,data_stage_5__5471_,data_stage_5__5470_,
  data_stage_5__5469_,data_stage_5__5468_,data_stage_5__5467_,data_stage_5__5466_,
  data_stage_5__5465_,data_stage_5__5464_,data_stage_5__5463_,data_stage_5__5462_,
  data_stage_5__5461_,data_stage_5__5460_,data_stage_5__5459_,data_stage_5__5458_,
  data_stage_5__5457_,data_stage_5__5456_,data_stage_5__5455_,data_stage_5__5454_,
  data_stage_5__5453_,data_stage_5__5452_,data_stage_5__5451_,data_stage_5__5450_,
  data_stage_5__5449_,data_stage_5__5448_,data_stage_5__5447_,data_stage_5__5446_,
  data_stage_5__5445_,data_stage_5__5444_,data_stage_5__5443_,data_stage_5__5442_,
  data_stage_5__5441_,data_stage_5__5440_,data_stage_5__5439_,data_stage_5__5438_,
  data_stage_5__5437_,data_stage_5__5436_,data_stage_5__5435_,data_stage_5__5434_,
  data_stage_5__5433_,data_stage_5__5432_,data_stage_5__5431_,data_stage_5__5430_,
  data_stage_5__5429_,data_stage_5__5428_,data_stage_5__5427_,data_stage_5__5426_,
  data_stage_5__5425_,data_stage_5__5424_,data_stage_5__5423_,data_stage_5__5422_,
  data_stage_5__5421_,data_stage_5__5420_,data_stage_5__5419_,data_stage_5__5418_,
  data_stage_5__5417_,data_stage_5__5416_,data_stage_5__5415_,data_stage_5__5414_,
  data_stage_5__5413_,data_stage_5__5412_,data_stage_5__5411_,data_stage_5__5410_,
  data_stage_5__5409_,data_stage_5__5408_,data_stage_5__5407_,data_stage_5__5406_,
  data_stage_5__5405_,data_stage_5__5404_,data_stage_5__5403_,data_stage_5__5402_,
  data_stage_5__5401_,data_stage_5__5400_,data_stage_5__5399_,data_stage_5__5398_,
  data_stage_5__5397_,data_stage_5__5396_,data_stage_5__5395_,data_stage_5__5394_,
  data_stage_5__5393_,data_stage_5__5392_,data_stage_5__5391_,data_stage_5__5390_,
  data_stage_5__5389_,data_stage_5__5388_,data_stage_5__5387_,data_stage_5__5386_,
  data_stage_5__5385_,data_stage_5__5384_,data_stage_5__5383_,data_stage_5__5382_,
  data_stage_5__5381_,data_stage_5__5380_,data_stage_5__5379_,data_stage_5__5378_,
  data_stage_5__5377_,data_stage_5__5376_,data_stage_5__5375_,data_stage_5__5374_,
  data_stage_5__5373_,data_stage_5__5372_,data_stage_5__5371_,data_stage_5__5370_,
  data_stage_5__5369_,data_stage_5__5368_,data_stage_5__5367_,data_stage_5__5366_,
  data_stage_5__5365_,data_stage_5__5364_,data_stage_5__5363_,data_stage_5__5362_,
  data_stage_5__5361_,data_stage_5__5360_,data_stage_5__5359_,data_stage_5__5358_,
  data_stage_5__5357_,data_stage_5__5356_,data_stage_5__5355_,data_stage_5__5354_,
  data_stage_5__5353_,data_stage_5__5352_,data_stage_5__5351_,data_stage_5__5350_,
  data_stage_5__5349_,data_stage_5__5348_,data_stage_5__5347_,data_stage_5__5346_,
  data_stage_5__5345_,data_stage_5__5344_,data_stage_5__5343_,data_stage_5__5342_,
  data_stage_5__5341_,data_stage_5__5340_,data_stage_5__5339_,data_stage_5__5338_,
  data_stage_5__5337_,data_stage_5__5336_,data_stage_5__5335_,data_stage_5__5334_,
  data_stage_5__5333_,data_stage_5__5332_,data_stage_5__5331_,data_stage_5__5330_,
  data_stage_5__5329_,data_stage_5__5328_,data_stage_5__5327_,data_stage_5__5326_,
  data_stage_5__5325_,data_stage_5__5324_,data_stage_5__5323_,data_stage_5__5322_,
  data_stage_5__5321_,data_stage_5__5320_,data_stage_5__5319_,data_stage_5__5318_,
  data_stage_5__5317_,data_stage_5__5316_,data_stage_5__5315_,data_stage_5__5314_,
  data_stage_5__5313_,data_stage_5__5312_,data_stage_5__5311_,data_stage_5__5310_,
  data_stage_5__5309_,data_stage_5__5308_,data_stage_5__5307_,data_stage_5__5306_,
  data_stage_5__5305_,data_stage_5__5304_,data_stage_5__5303_,data_stage_5__5302_,
  data_stage_5__5301_,data_stage_5__5300_,data_stage_5__5299_,data_stage_5__5298_,
  data_stage_5__5297_,data_stage_5__5296_,data_stage_5__5295_,data_stage_5__5294_,
  data_stage_5__5293_,data_stage_5__5292_,data_stage_5__5291_,data_stage_5__5290_,
  data_stage_5__5289_,data_stage_5__5288_,data_stage_5__5287_,data_stage_5__5286_,
  data_stage_5__5285_,data_stage_5__5284_,data_stage_5__5283_,data_stage_5__5282_,
  data_stage_5__5281_,data_stage_5__5280_,data_stage_5__5279_,data_stage_5__5278_,
  data_stage_5__5277_,data_stage_5__5276_,data_stage_5__5275_,data_stage_5__5274_,
  data_stage_5__5273_,data_stage_5__5272_,data_stage_5__5271_,data_stage_5__5270_,
  data_stage_5__5269_,data_stage_5__5268_,data_stage_5__5267_,data_stage_5__5266_,
  data_stage_5__5265_,data_stage_5__5264_,data_stage_5__5263_,data_stage_5__5262_,
  data_stage_5__5261_,data_stage_5__5260_,data_stage_5__5259_,data_stage_5__5258_,
  data_stage_5__5257_,data_stage_5__5256_,data_stage_5__5255_,data_stage_5__5254_,
  data_stage_5__5253_,data_stage_5__5252_,data_stage_5__5251_,data_stage_5__5250_,
  data_stage_5__5249_,data_stage_5__5248_,data_stage_5__5247_,data_stage_5__5246_,
  data_stage_5__5245_,data_stage_5__5244_,data_stage_5__5243_,data_stage_5__5242_,
  data_stage_5__5241_,data_stage_5__5240_,data_stage_5__5239_,data_stage_5__5238_,
  data_stage_5__5237_,data_stage_5__5236_,data_stage_5__5235_,data_stage_5__5234_,
  data_stage_5__5233_,data_stage_5__5232_,data_stage_5__5231_,data_stage_5__5230_,
  data_stage_5__5229_,data_stage_5__5228_,data_stage_5__5227_,data_stage_5__5226_,
  data_stage_5__5225_,data_stage_5__5224_,data_stage_5__5223_,data_stage_5__5222_,
  data_stage_5__5221_,data_stage_5__5220_,data_stage_5__5219_,data_stage_5__5218_,
  data_stage_5__5217_,data_stage_5__5216_,data_stage_5__5215_,data_stage_5__5214_,
  data_stage_5__5213_,data_stage_5__5212_,data_stage_5__5211_,data_stage_5__5210_,
  data_stage_5__5209_,data_stage_5__5208_,data_stage_5__5207_,data_stage_5__5206_,
  data_stage_5__5205_,data_stage_5__5204_,data_stage_5__5203_,data_stage_5__5202_,
  data_stage_5__5201_,data_stage_5__5200_,data_stage_5__5199_,data_stage_5__5198_,
  data_stage_5__5197_,data_stage_5__5196_,data_stage_5__5195_,data_stage_5__5194_,
  data_stage_5__5193_,data_stage_5__5192_,data_stage_5__5191_,data_stage_5__5190_,
  data_stage_5__5189_,data_stage_5__5188_,data_stage_5__5187_,data_stage_5__5186_,
  data_stage_5__5185_,data_stage_5__5184_,data_stage_5__5183_,data_stage_5__5182_,
  data_stage_5__5181_,data_stage_5__5180_,data_stage_5__5179_,data_stage_5__5178_,
  data_stage_5__5177_,data_stage_5__5176_,data_stage_5__5175_,data_stage_5__5174_,
  data_stage_5__5173_,data_stage_5__5172_,data_stage_5__5171_,data_stage_5__5170_,
  data_stage_5__5169_,data_stage_5__5168_,data_stage_5__5167_,data_stage_5__5166_,
  data_stage_5__5165_,data_stage_5__5164_,data_stage_5__5163_,data_stage_5__5162_,
  data_stage_5__5161_,data_stage_5__5160_,data_stage_5__5159_,data_stage_5__5158_,
  data_stage_5__5157_,data_stage_5__5156_,data_stage_5__5155_,data_stage_5__5154_,
  data_stage_5__5153_,data_stage_5__5152_,data_stage_5__5151_,data_stage_5__5150_,
  data_stage_5__5149_,data_stage_5__5148_,data_stage_5__5147_,data_stage_5__5146_,
  data_stage_5__5145_,data_stage_5__5144_,data_stage_5__5143_,data_stage_5__5142_,
  data_stage_5__5141_,data_stage_5__5140_,data_stage_5__5139_,data_stage_5__5138_,
  data_stage_5__5137_,data_stage_5__5136_,data_stage_5__5135_,data_stage_5__5134_,
  data_stage_5__5133_,data_stage_5__5132_,data_stage_5__5131_,data_stage_5__5130_,
  data_stage_5__5129_,data_stage_5__5128_,data_stage_5__5127_,data_stage_5__5126_,
  data_stage_5__5125_,data_stage_5__5124_,data_stage_5__5123_,data_stage_5__5122_,
  data_stage_5__5121_,data_stage_5__5120_,data_stage_5__5119_,data_stage_5__5118_,
  data_stage_5__5117_,data_stage_5__5116_,data_stage_5__5115_,data_stage_5__5114_,
  data_stage_5__5113_,data_stage_5__5112_,data_stage_5__5111_,data_stage_5__5110_,
  data_stage_5__5109_,data_stage_5__5108_,data_stage_5__5107_,data_stage_5__5106_,
  data_stage_5__5105_,data_stage_5__5104_,data_stage_5__5103_,data_stage_5__5102_,
  data_stage_5__5101_,data_stage_5__5100_,data_stage_5__5099_,data_stage_5__5098_,
  data_stage_5__5097_,data_stage_5__5096_,data_stage_5__5095_,data_stage_5__5094_,
  data_stage_5__5093_,data_stage_5__5092_,data_stage_5__5091_,data_stage_5__5090_,
  data_stage_5__5089_,data_stage_5__5088_,data_stage_5__5087_,data_stage_5__5086_,
  data_stage_5__5085_,data_stage_5__5084_,data_stage_5__5083_,data_stage_5__5082_,
  data_stage_5__5081_,data_stage_5__5080_,data_stage_5__5079_,data_stage_5__5078_,
  data_stage_5__5077_,data_stage_5__5076_,data_stage_5__5075_,data_stage_5__5074_,
  data_stage_5__5073_,data_stage_5__5072_,data_stage_5__5071_,data_stage_5__5070_,
  data_stage_5__5069_,data_stage_5__5068_,data_stage_5__5067_,data_stage_5__5066_,
  data_stage_5__5065_,data_stage_5__5064_,data_stage_5__5063_,data_stage_5__5062_,
  data_stage_5__5061_,data_stage_5__5060_,data_stage_5__5059_,data_stage_5__5058_,
  data_stage_5__5057_,data_stage_5__5056_,data_stage_5__5055_,data_stage_5__5054_,
  data_stage_5__5053_,data_stage_5__5052_,data_stage_5__5051_,data_stage_5__5050_,
  data_stage_5__5049_,data_stage_5__5048_,data_stage_5__5047_,data_stage_5__5046_,
  data_stage_5__5045_,data_stage_5__5044_,data_stage_5__5043_,data_stage_5__5042_,
  data_stage_5__5041_,data_stage_5__5040_,data_stage_5__5039_,data_stage_5__5038_,
  data_stage_5__5037_,data_stage_5__5036_,data_stage_5__5035_,data_stage_5__5034_,
  data_stage_5__5033_,data_stage_5__5032_,data_stage_5__5031_,data_stage_5__5030_,
  data_stage_5__5029_,data_stage_5__5028_,data_stage_5__5027_,data_stage_5__5026_,
  data_stage_5__5025_,data_stage_5__5024_,data_stage_5__5023_,data_stage_5__5022_,
  data_stage_5__5021_,data_stage_5__5020_,data_stage_5__5019_,data_stage_5__5018_,
  data_stage_5__5017_,data_stage_5__5016_,data_stage_5__5015_,data_stage_5__5014_,
  data_stage_5__5013_,data_stage_5__5012_,data_stage_5__5011_,data_stage_5__5010_,
  data_stage_5__5009_,data_stage_5__5008_,data_stage_5__5007_,data_stage_5__5006_,
  data_stage_5__5005_,data_stage_5__5004_,data_stage_5__5003_,data_stage_5__5002_,
  data_stage_5__5001_,data_stage_5__5000_,data_stage_5__4999_,data_stage_5__4998_,
  data_stage_5__4997_,data_stage_5__4996_,data_stage_5__4995_,data_stage_5__4994_,
  data_stage_5__4993_,data_stage_5__4992_,data_stage_5__4991_,data_stage_5__4990_,
  data_stage_5__4989_,data_stage_5__4988_,data_stage_5__4987_,data_stage_5__4986_,
  data_stage_5__4985_,data_stage_5__4984_,data_stage_5__4983_,data_stage_5__4982_,
  data_stage_5__4981_,data_stage_5__4980_,data_stage_5__4979_,data_stage_5__4978_,
  data_stage_5__4977_,data_stage_5__4976_,data_stage_5__4975_,data_stage_5__4974_,
  data_stage_5__4973_,data_stage_5__4972_,data_stage_5__4971_,data_stage_5__4970_,
  data_stage_5__4969_,data_stage_5__4968_,data_stage_5__4967_,data_stage_5__4966_,
  data_stage_5__4965_,data_stage_5__4964_,data_stage_5__4963_,data_stage_5__4962_,
  data_stage_5__4961_,data_stage_5__4960_,data_stage_5__4959_,data_stage_5__4958_,
  data_stage_5__4957_,data_stage_5__4956_,data_stage_5__4955_,data_stage_5__4954_,
  data_stage_5__4953_,data_stage_5__4952_,data_stage_5__4951_,data_stage_5__4950_,
  data_stage_5__4949_,data_stage_5__4948_,data_stage_5__4947_,data_stage_5__4946_,
  data_stage_5__4945_,data_stage_5__4944_,data_stage_5__4943_,data_stage_5__4942_,
  data_stage_5__4941_,data_stage_5__4940_,data_stage_5__4939_,data_stage_5__4938_,
  data_stage_5__4937_,data_stage_5__4936_,data_stage_5__4935_,data_stage_5__4934_,
  data_stage_5__4933_,data_stage_5__4932_,data_stage_5__4931_,data_stage_5__4930_,
  data_stage_5__4929_,data_stage_5__4928_,data_stage_5__4927_,data_stage_5__4926_,
  data_stage_5__4925_,data_stage_5__4924_,data_stage_5__4923_,data_stage_5__4922_,
  data_stage_5__4921_,data_stage_5__4920_,data_stage_5__4919_,data_stage_5__4918_,
  data_stage_5__4917_,data_stage_5__4916_,data_stage_5__4915_,data_stage_5__4914_,
  data_stage_5__4913_,data_stage_5__4912_,data_stage_5__4911_,data_stage_5__4910_,
  data_stage_5__4909_,data_stage_5__4908_,data_stage_5__4907_,data_stage_5__4906_,
  data_stage_5__4905_,data_stage_5__4904_,data_stage_5__4903_,data_stage_5__4902_,
  data_stage_5__4901_,data_stage_5__4900_,data_stage_5__4899_,data_stage_5__4898_,
  data_stage_5__4897_,data_stage_5__4896_,data_stage_5__4895_,data_stage_5__4894_,
  data_stage_5__4893_,data_stage_5__4892_,data_stage_5__4891_,data_stage_5__4890_,
  data_stage_5__4889_,data_stage_5__4888_,data_stage_5__4887_,data_stage_5__4886_,
  data_stage_5__4885_,data_stage_5__4884_,data_stage_5__4883_,data_stage_5__4882_,
  data_stage_5__4881_,data_stage_5__4880_,data_stage_5__4879_,data_stage_5__4878_,
  data_stage_5__4877_,data_stage_5__4876_,data_stage_5__4875_,data_stage_5__4874_,
  data_stage_5__4873_,data_stage_5__4872_,data_stage_5__4871_,data_stage_5__4870_,
  data_stage_5__4869_,data_stage_5__4868_,data_stage_5__4867_,data_stage_5__4866_,
  data_stage_5__4865_,data_stage_5__4864_,data_stage_5__4863_,data_stage_5__4862_,
  data_stage_5__4861_,data_stage_5__4860_,data_stage_5__4859_,data_stage_5__4858_,
  data_stage_5__4857_,data_stage_5__4856_,data_stage_5__4855_,data_stage_5__4854_,
  data_stage_5__4853_,data_stage_5__4852_,data_stage_5__4851_,data_stage_5__4850_,
  data_stage_5__4849_,data_stage_5__4848_,data_stage_5__4847_,data_stage_5__4846_,
  data_stage_5__4845_,data_stage_5__4844_,data_stage_5__4843_,data_stage_5__4842_,
  data_stage_5__4841_,data_stage_5__4840_,data_stage_5__4839_,data_stage_5__4838_,
  data_stage_5__4837_,data_stage_5__4836_,data_stage_5__4835_,data_stage_5__4834_,
  data_stage_5__4833_,data_stage_5__4832_,data_stage_5__4831_,data_stage_5__4830_,
  data_stage_5__4829_,data_stage_5__4828_,data_stage_5__4827_,data_stage_5__4826_,
  data_stage_5__4825_,data_stage_5__4824_,data_stage_5__4823_,data_stage_5__4822_,
  data_stage_5__4821_,data_stage_5__4820_,data_stage_5__4819_,data_stage_5__4818_,
  data_stage_5__4817_,data_stage_5__4816_,data_stage_5__4815_,data_stage_5__4814_,
  data_stage_5__4813_,data_stage_5__4812_,data_stage_5__4811_,data_stage_5__4810_,
  data_stage_5__4809_,data_stage_5__4808_,data_stage_5__4807_,data_stage_5__4806_,
  data_stage_5__4805_,data_stage_5__4804_,data_stage_5__4803_,data_stage_5__4802_,
  data_stage_5__4801_,data_stage_5__4800_,data_stage_5__4799_,data_stage_5__4798_,
  data_stage_5__4797_,data_stage_5__4796_,data_stage_5__4795_,data_stage_5__4794_,
  data_stage_5__4793_,data_stage_5__4792_,data_stage_5__4791_,data_stage_5__4790_,
  data_stage_5__4789_,data_stage_5__4788_,data_stage_5__4787_,data_stage_5__4786_,
  data_stage_5__4785_,data_stage_5__4784_,data_stage_5__4783_,data_stage_5__4782_,
  data_stage_5__4781_,data_stage_5__4780_,data_stage_5__4779_,data_stage_5__4778_,
  data_stage_5__4777_,data_stage_5__4776_,data_stage_5__4775_,data_stage_5__4774_,
  data_stage_5__4773_,data_stage_5__4772_,data_stage_5__4771_,data_stage_5__4770_,
  data_stage_5__4769_,data_stage_5__4768_,data_stage_5__4767_,data_stage_5__4766_,
  data_stage_5__4765_,data_stage_5__4764_,data_stage_5__4763_,data_stage_5__4762_,
  data_stage_5__4761_,data_stage_5__4760_,data_stage_5__4759_,data_stage_5__4758_,
  data_stage_5__4757_,data_stage_5__4756_,data_stage_5__4755_,data_stage_5__4754_,
  data_stage_5__4753_,data_stage_5__4752_,data_stage_5__4751_,data_stage_5__4750_,
  data_stage_5__4749_,data_stage_5__4748_,data_stage_5__4747_,data_stage_5__4746_,
  data_stage_5__4745_,data_stage_5__4744_,data_stage_5__4743_,data_stage_5__4742_,
  data_stage_5__4741_,data_stage_5__4740_,data_stage_5__4739_,data_stage_5__4738_,
  data_stage_5__4737_,data_stage_5__4736_,data_stage_5__4735_,data_stage_5__4734_,
  data_stage_5__4733_,data_stage_5__4732_,data_stage_5__4731_,data_stage_5__4730_,
  data_stage_5__4729_,data_stage_5__4728_,data_stage_5__4727_,data_stage_5__4726_,
  data_stage_5__4725_,data_stage_5__4724_,data_stage_5__4723_,data_stage_5__4722_,
  data_stage_5__4721_,data_stage_5__4720_,data_stage_5__4719_,data_stage_5__4718_,
  data_stage_5__4717_,data_stage_5__4716_,data_stage_5__4715_,data_stage_5__4714_,
  data_stage_5__4713_,data_stage_5__4712_,data_stage_5__4711_,data_stage_5__4710_,
  data_stage_5__4709_,data_stage_5__4708_,data_stage_5__4707_,data_stage_5__4706_,
  data_stage_5__4705_,data_stage_5__4704_,data_stage_5__4703_,data_stage_5__4702_,
  data_stage_5__4701_,data_stage_5__4700_,data_stage_5__4699_,data_stage_5__4698_,
  data_stage_5__4697_,data_stage_5__4696_,data_stage_5__4695_,data_stage_5__4694_,
  data_stage_5__4693_,data_stage_5__4692_,data_stage_5__4691_,data_stage_5__4690_,
  data_stage_5__4689_,data_stage_5__4688_,data_stage_5__4687_,data_stage_5__4686_,
  data_stage_5__4685_,data_stage_5__4684_,data_stage_5__4683_,data_stage_5__4682_,
  data_stage_5__4681_,data_stage_5__4680_,data_stage_5__4679_,data_stage_5__4678_,
  data_stage_5__4677_,data_stage_5__4676_,data_stage_5__4675_,data_stage_5__4674_,
  data_stage_5__4673_,data_stage_5__4672_,data_stage_5__4671_,data_stage_5__4670_,
  data_stage_5__4669_,data_stage_5__4668_,data_stage_5__4667_,data_stage_5__4666_,
  data_stage_5__4665_,data_stage_5__4664_,data_stage_5__4663_,data_stage_5__4662_,
  data_stage_5__4661_,data_stage_5__4660_,data_stage_5__4659_,data_stage_5__4658_,
  data_stage_5__4657_,data_stage_5__4656_,data_stage_5__4655_,data_stage_5__4654_,
  data_stage_5__4653_,data_stage_5__4652_,data_stage_5__4651_,data_stage_5__4650_,
  data_stage_5__4649_,data_stage_5__4648_,data_stage_5__4647_,data_stage_5__4646_,
  data_stage_5__4645_,data_stage_5__4644_,data_stage_5__4643_,data_stage_5__4642_,
  data_stage_5__4641_,data_stage_5__4640_,data_stage_5__4639_,data_stage_5__4638_,
  data_stage_5__4637_,data_stage_5__4636_,data_stage_5__4635_,data_stage_5__4634_,
  data_stage_5__4633_,data_stage_5__4632_,data_stage_5__4631_,data_stage_5__4630_,
  data_stage_5__4629_,data_stage_5__4628_,data_stage_5__4627_,data_stage_5__4626_,
  data_stage_5__4625_,data_stage_5__4624_,data_stage_5__4623_,data_stage_5__4622_,
  data_stage_5__4621_,data_stage_5__4620_,data_stage_5__4619_,data_stage_5__4618_,
  data_stage_5__4617_,data_stage_5__4616_,data_stage_5__4615_,data_stage_5__4614_,
  data_stage_5__4613_,data_stage_5__4612_,data_stage_5__4611_,data_stage_5__4610_,
  data_stage_5__4609_,data_stage_5__4608_,data_stage_5__4607_,data_stage_5__4606_,
  data_stage_5__4605_,data_stage_5__4604_,data_stage_5__4603_,data_stage_5__4602_,
  data_stage_5__4601_,data_stage_5__4600_,data_stage_5__4599_,data_stage_5__4598_,
  data_stage_5__4597_,data_stage_5__4596_,data_stage_5__4595_,data_stage_5__4594_,
  data_stage_5__4593_,data_stage_5__4592_,data_stage_5__4591_,data_stage_5__4590_,
  data_stage_5__4589_,data_stage_5__4588_,data_stage_5__4587_,data_stage_5__4586_,
  data_stage_5__4585_,data_stage_5__4584_,data_stage_5__4583_,data_stage_5__4582_,
  data_stage_5__4581_,data_stage_5__4580_,data_stage_5__4579_,data_stage_5__4578_,
  data_stage_5__4577_,data_stage_5__4576_,data_stage_5__4575_,data_stage_5__4574_,
  data_stage_5__4573_,data_stage_5__4572_,data_stage_5__4571_,data_stage_5__4570_,
  data_stage_5__4569_,data_stage_5__4568_,data_stage_5__4567_,data_stage_5__4566_,
  data_stage_5__4565_,data_stage_5__4564_,data_stage_5__4563_,data_stage_5__4562_,
  data_stage_5__4561_,data_stage_5__4560_,data_stage_5__4559_,data_stage_5__4558_,
  data_stage_5__4557_,data_stage_5__4556_,data_stage_5__4555_,data_stage_5__4554_,
  data_stage_5__4553_,data_stage_5__4552_,data_stage_5__4551_,data_stage_5__4550_,
  data_stage_5__4549_,data_stage_5__4548_,data_stage_5__4547_,data_stage_5__4546_,
  data_stage_5__4545_,data_stage_5__4544_,data_stage_5__4543_,data_stage_5__4542_,
  data_stage_5__4541_,data_stage_5__4540_,data_stage_5__4539_,data_stage_5__4538_,
  data_stage_5__4537_,data_stage_5__4536_,data_stage_5__4535_,data_stage_5__4534_,
  data_stage_5__4533_,data_stage_5__4532_,data_stage_5__4531_,data_stage_5__4530_,
  data_stage_5__4529_,data_stage_5__4528_,data_stage_5__4527_,data_stage_5__4526_,
  data_stage_5__4525_,data_stage_5__4524_,data_stage_5__4523_,data_stage_5__4522_,
  data_stage_5__4521_,data_stage_5__4520_,data_stage_5__4519_,data_stage_5__4518_,
  data_stage_5__4517_,data_stage_5__4516_,data_stage_5__4515_,data_stage_5__4514_,
  data_stage_5__4513_,data_stage_5__4512_,data_stage_5__4511_,data_stage_5__4510_,
  data_stage_5__4509_,data_stage_5__4508_,data_stage_5__4507_,data_stage_5__4506_,
  data_stage_5__4505_,data_stage_5__4504_,data_stage_5__4503_,data_stage_5__4502_,
  data_stage_5__4501_,data_stage_5__4500_,data_stage_5__4499_,data_stage_5__4498_,
  data_stage_5__4497_,data_stage_5__4496_,data_stage_5__4495_,data_stage_5__4494_,
  data_stage_5__4493_,data_stage_5__4492_,data_stage_5__4491_,data_stage_5__4490_,
  data_stage_5__4489_,data_stage_5__4488_,data_stage_5__4487_,data_stage_5__4486_,
  data_stage_5__4485_,data_stage_5__4484_,data_stage_5__4483_,data_stage_5__4482_,
  data_stage_5__4481_,data_stage_5__4480_,data_stage_5__4479_,data_stage_5__4478_,
  data_stage_5__4477_,data_stage_5__4476_,data_stage_5__4475_,data_stage_5__4474_,
  data_stage_5__4473_,data_stage_5__4472_,data_stage_5__4471_,data_stage_5__4470_,
  data_stage_5__4469_,data_stage_5__4468_,data_stage_5__4467_,data_stage_5__4466_,
  data_stage_5__4465_,data_stage_5__4464_,data_stage_5__4463_,data_stage_5__4462_,
  data_stage_5__4461_,data_stage_5__4460_,data_stage_5__4459_,data_stage_5__4458_,
  data_stage_5__4457_,data_stage_5__4456_,data_stage_5__4455_,data_stage_5__4454_,
  data_stage_5__4453_,data_stage_5__4452_,data_stage_5__4451_,data_stage_5__4450_,
  data_stage_5__4449_,data_stage_5__4448_,data_stage_5__4447_,data_stage_5__4446_,
  data_stage_5__4445_,data_stage_5__4444_,data_stage_5__4443_,data_stage_5__4442_,
  data_stage_5__4441_,data_stage_5__4440_,data_stage_5__4439_,data_stage_5__4438_,
  data_stage_5__4437_,data_stage_5__4436_,data_stage_5__4435_,data_stage_5__4434_,
  data_stage_5__4433_,data_stage_5__4432_,data_stage_5__4431_,data_stage_5__4430_,
  data_stage_5__4429_,data_stage_5__4428_,data_stage_5__4427_,data_stage_5__4426_,
  data_stage_5__4425_,data_stage_5__4424_,data_stage_5__4423_,data_stage_5__4422_,
  data_stage_5__4421_,data_stage_5__4420_,data_stage_5__4419_,data_stage_5__4418_,
  data_stage_5__4417_,data_stage_5__4416_,data_stage_5__4415_,data_stage_5__4414_,
  data_stage_5__4413_,data_stage_5__4412_,data_stage_5__4411_,data_stage_5__4410_,
  data_stage_5__4409_,data_stage_5__4408_,data_stage_5__4407_,data_stage_5__4406_,
  data_stage_5__4405_,data_stage_5__4404_,data_stage_5__4403_,data_stage_5__4402_,
  data_stage_5__4401_,data_stage_5__4400_,data_stage_5__4399_,data_stage_5__4398_,
  data_stage_5__4397_,data_stage_5__4396_,data_stage_5__4395_,data_stage_5__4394_,
  data_stage_5__4393_,data_stage_5__4392_,data_stage_5__4391_,data_stage_5__4390_,
  data_stage_5__4389_,data_stage_5__4388_,data_stage_5__4387_,data_stage_5__4386_,
  data_stage_5__4385_,data_stage_5__4384_,data_stage_5__4383_,data_stage_5__4382_,
  data_stage_5__4381_,data_stage_5__4380_,data_stage_5__4379_,data_stage_5__4378_,
  data_stage_5__4377_,data_stage_5__4376_,data_stage_5__4375_,data_stage_5__4374_,
  data_stage_5__4373_,data_stage_5__4372_,data_stage_5__4371_,data_stage_5__4370_,
  data_stage_5__4369_,data_stage_5__4368_,data_stage_5__4367_,data_stage_5__4366_,
  data_stage_5__4365_,data_stage_5__4364_,data_stage_5__4363_,data_stage_5__4362_,
  data_stage_5__4361_,data_stage_5__4360_,data_stage_5__4359_,data_stage_5__4358_,
  data_stage_5__4357_,data_stage_5__4356_,data_stage_5__4355_,data_stage_5__4354_,
  data_stage_5__4353_,data_stage_5__4352_,data_stage_5__4351_,data_stage_5__4350_,
  data_stage_5__4349_,data_stage_5__4348_,data_stage_5__4347_,data_stage_5__4346_,
  data_stage_5__4345_,data_stage_5__4344_,data_stage_5__4343_,data_stage_5__4342_,
  data_stage_5__4341_,data_stage_5__4340_,data_stage_5__4339_,data_stage_5__4338_,
  data_stage_5__4337_,data_stage_5__4336_,data_stage_5__4335_,data_stage_5__4334_,
  data_stage_5__4333_,data_stage_5__4332_,data_stage_5__4331_,data_stage_5__4330_,
  data_stage_5__4329_,data_stage_5__4328_,data_stage_5__4327_,data_stage_5__4326_,
  data_stage_5__4325_,data_stage_5__4324_,data_stage_5__4323_,data_stage_5__4322_,
  data_stage_5__4321_,data_stage_5__4320_,data_stage_5__4319_,data_stage_5__4318_,
  data_stage_5__4317_,data_stage_5__4316_,data_stage_5__4315_,data_stage_5__4314_,
  data_stage_5__4313_,data_stage_5__4312_,data_stage_5__4311_,data_stage_5__4310_,
  data_stage_5__4309_,data_stage_5__4308_,data_stage_5__4307_,data_stage_5__4306_,
  data_stage_5__4305_,data_stage_5__4304_,data_stage_5__4303_,data_stage_5__4302_,
  data_stage_5__4301_,data_stage_5__4300_,data_stage_5__4299_,data_stage_5__4298_,
  data_stage_5__4297_,data_stage_5__4296_,data_stage_5__4295_,data_stage_5__4294_,
  data_stage_5__4293_,data_stage_5__4292_,data_stage_5__4291_,data_stage_5__4290_,
  data_stage_5__4289_,data_stage_5__4288_,data_stage_5__4287_,data_stage_5__4286_,
  data_stage_5__4285_,data_stage_5__4284_,data_stage_5__4283_,data_stage_5__4282_,
  data_stage_5__4281_,data_stage_5__4280_,data_stage_5__4279_,data_stage_5__4278_,
  data_stage_5__4277_,data_stage_5__4276_,data_stage_5__4275_,data_stage_5__4274_,
  data_stage_5__4273_,data_stage_5__4272_,data_stage_5__4271_,data_stage_5__4270_,
  data_stage_5__4269_,data_stage_5__4268_,data_stage_5__4267_,data_stage_5__4266_,
  data_stage_5__4265_,data_stage_5__4264_,data_stage_5__4263_,data_stage_5__4262_,
  data_stage_5__4261_,data_stage_5__4260_,data_stage_5__4259_,data_stage_5__4258_,
  data_stage_5__4257_,data_stage_5__4256_,data_stage_5__4255_,data_stage_5__4254_,
  data_stage_5__4253_,data_stage_5__4252_,data_stage_5__4251_,data_stage_5__4250_,
  data_stage_5__4249_,data_stage_5__4248_,data_stage_5__4247_,data_stage_5__4246_,
  data_stage_5__4245_,data_stage_5__4244_,data_stage_5__4243_,data_stage_5__4242_,
  data_stage_5__4241_,data_stage_5__4240_,data_stage_5__4239_,data_stage_5__4238_,
  data_stage_5__4237_,data_stage_5__4236_,data_stage_5__4235_,data_stage_5__4234_,
  data_stage_5__4233_,data_stage_5__4232_,data_stage_5__4231_,data_stage_5__4230_,
  data_stage_5__4229_,data_stage_5__4228_,data_stage_5__4227_,data_stage_5__4226_,
  data_stage_5__4225_,data_stage_5__4224_,data_stage_5__4223_,data_stage_5__4222_,
  data_stage_5__4221_,data_stage_5__4220_,data_stage_5__4219_,data_stage_5__4218_,
  data_stage_5__4217_,data_stage_5__4216_,data_stage_5__4215_,data_stage_5__4214_,
  data_stage_5__4213_,data_stage_5__4212_,data_stage_5__4211_,data_stage_5__4210_,
  data_stage_5__4209_,data_stage_5__4208_,data_stage_5__4207_,data_stage_5__4206_,
  data_stage_5__4205_,data_stage_5__4204_,data_stage_5__4203_,data_stage_5__4202_,
  data_stage_5__4201_,data_stage_5__4200_,data_stage_5__4199_,data_stage_5__4198_,
  data_stage_5__4197_,data_stage_5__4196_,data_stage_5__4195_,data_stage_5__4194_,
  data_stage_5__4193_,data_stage_5__4192_,data_stage_5__4191_,data_stage_5__4190_,
  data_stage_5__4189_,data_stage_5__4188_,data_stage_5__4187_,data_stage_5__4186_,
  data_stage_5__4185_,data_stage_5__4184_,data_stage_5__4183_,data_stage_5__4182_,
  data_stage_5__4181_,data_stage_5__4180_,data_stage_5__4179_,data_stage_5__4178_,
  data_stage_5__4177_,data_stage_5__4176_,data_stage_5__4175_,data_stage_5__4174_,
  data_stage_5__4173_,data_stage_5__4172_,data_stage_5__4171_,data_stage_5__4170_,
  data_stage_5__4169_,data_stage_5__4168_,data_stage_5__4167_,data_stage_5__4166_,
  data_stage_5__4165_,data_stage_5__4164_,data_stage_5__4163_,data_stage_5__4162_,
  data_stage_5__4161_,data_stage_5__4160_,data_stage_5__4159_,data_stage_5__4158_,
  data_stage_5__4157_,data_stage_5__4156_,data_stage_5__4155_,data_stage_5__4154_,
  data_stage_5__4153_,data_stage_5__4152_,data_stage_5__4151_,data_stage_5__4150_,
  data_stage_5__4149_,data_stage_5__4148_,data_stage_5__4147_,data_stage_5__4146_,
  data_stage_5__4145_,data_stage_5__4144_,data_stage_5__4143_,data_stage_5__4142_,
  data_stage_5__4141_,data_stage_5__4140_,data_stage_5__4139_,data_stage_5__4138_,
  data_stage_5__4137_,data_stage_5__4136_,data_stage_5__4135_,data_stage_5__4134_,
  data_stage_5__4133_,data_stage_5__4132_,data_stage_5__4131_,data_stage_5__4130_,
  data_stage_5__4129_,data_stage_5__4128_,data_stage_5__4127_,data_stage_5__4126_,
  data_stage_5__4125_,data_stage_5__4124_,data_stage_5__4123_,data_stage_5__4122_,
  data_stage_5__4121_,data_stage_5__4120_,data_stage_5__4119_,data_stage_5__4118_,
  data_stage_5__4117_,data_stage_5__4116_,data_stage_5__4115_,data_stage_5__4114_,
  data_stage_5__4113_,data_stage_5__4112_,data_stage_5__4111_,data_stage_5__4110_,
  data_stage_5__4109_,data_stage_5__4108_,data_stage_5__4107_,data_stage_5__4106_,
  data_stage_5__4105_,data_stage_5__4104_,data_stage_5__4103_,data_stage_5__4102_,
  data_stage_5__4101_,data_stage_5__4100_,data_stage_5__4099_,data_stage_5__4098_,
  data_stage_5__4097_,data_stage_5__4096_,data_stage_5__4095_,data_stage_5__4094_,
  data_stage_5__4093_,data_stage_5__4092_,data_stage_5__4091_,data_stage_5__4090_,
  data_stage_5__4089_,data_stage_5__4088_,data_stage_5__4087_,data_stage_5__4086_,
  data_stage_5__4085_,data_stage_5__4084_,data_stage_5__4083_,data_stage_5__4082_,
  data_stage_5__4081_,data_stage_5__4080_,data_stage_5__4079_,data_stage_5__4078_,
  data_stage_5__4077_,data_stage_5__4076_,data_stage_5__4075_,data_stage_5__4074_,
  data_stage_5__4073_,data_stage_5__4072_,data_stage_5__4071_,data_stage_5__4070_,
  data_stage_5__4069_,data_stage_5__4068_,data_stage_5__4067_,data_stage_5__4066_,
  data_stage_5__4065_,data_stage_5__4064_,data_stage_5__4063_,data_stage_5__4062_,
  data_stage_5__4061_,data_stage_5__4060_,data_stage_5__4059_,data_stage_5__4058_,
  data_stage_5__4057_,data_stage_5__4056_,data_stage_5__4055_,data_stage_5__4054_,
  data_stage_5__4053_,data_stage_5__4052_,data_stage_5__4051_,data_stage_5__4050_,
  data_stage_5__4049_,data_stage_5__4048_,data_stage_5__4047_,data_stage_5__4046_,
  data_stage_5__4045_,data_stage_5__4044_,data_stage_5__4043_,data_stage_5__4042_,
  data_stage_5__4041_,data_stage_5__4040_,data_stage_5__4039_,data_stage_5__4038_,
  data_stage_5__4037_,data_stage_5__4036_,data_stage_5__4035_,data_stage_5__4034_,
  data_stage_5__4033_,data_stage_5__4032_,data_stage_5__4031_,data_stage_5__4030_,
  data_stage_5__4029_,data_stage_5__4028_,data_stage_5__4027_,data_stage_5__4026_,
  data_stage_5__4025_,data_stage_5__4024_,data_stage_5__4023_,data_stage_5__4022_,
  data_stage_5__4021_,data_stage_5__4020_,data_stage_5__4019_,data_stage_5__4018_,
  data_stage_5__4017_,data_stage_5__4016_,data_stage_5__4015_,data_stage_5__4014_,
  data_stage_5__4013_,data_stage_5__4012_,data_stage_5__4011_,data_stage_5__4010_,
  data_stage_5__4009_,data_stage_5__4008_,data_stage_5__4007_,data_stage_5__4006_,
  data_stage_5__4005_,data_stage_5__4004_,data_stage_5__4003_,data_stage_5__4002_,
  data_stage_5__4001_,data_stage_5__4000_,data_stage_5__3999_,data_stage_5__3998_,
  data_stage_5__3997_,data_stage_5__3996_,data_stage_5__3995_,data_stage_5__3994_,
  data_stage_5__3993_,data_stage_5__3992_,data_stage_5__3991_,data_stage_5__3990_,
  data_stage_5__3989_,data_stage_5__3988_,data_stage_5__3987_,data_stage_5__3986_,
  data_stage_5__3985_,data_stage_5__3984_,data_stage_5__3983_,data_stage_5__3982_,
  data_stage_5__3981_,data_stage_5__3980_,data_stage_5__3979_,data_stage_5__3978_,
  data_stage_5__3977_,data_stage_5__3976_,data_stage_5__3975_,data_stage_5__3974_,
  data_stage_5__3973_,data_stage_5__3972_,data_stage_5__3971_,data_stage_5__3970_,
  data_stage_5__3969_,data_stage_5__3968_,data_stage_5__3967_,data_stage_5__3966_,
  data_stage_5__3965_,data_stage_5__3964_,data_stage_5__3963_,data_stage_5__3962_,
  data_stage_5__3961_,data_stage_5__3960_,data_stage_5__3959_,data_stage_5__3958_,
  data_stage_5__3957_,data_stage_5__3956_,data_stage_5__3955_,data_stage_5__3954_,
  data_stage_5__3953_,data_stage_5__3952_,data_stage_5__3951_,data_stage_5__3950_,
  data_stage_5__3949_,data_stage_5__3948_,data_stage_5__3947_,data_stage_5__3946_,
  data_stage_5__3945_,data_stage_5__3944_,data_stage_5__3943_,data_stage_5__3942_,
  data_stage_5__3941_,data_stage_5__3940_,data_stage_5__3939_,data_stage_5__3938_,
  data_stage_5__3937_,data_stage_5__3936_,data_stage_5__3935_,data_stage_5__3934_,
  data_stage_5__3933_,data_stage_5__3932_,data_stage_5__3931_,data_stage_5__3930_,
  data_stage_5__3929_,data_stage_5__3928_,data_stage_5__3927_,data_stage_5__3926_,
  data_stage_5__3925_,data_stage_5__3924_,data_stage_5__3923_,data_stage_5__3922_,
  data_stage_5__3921_,data_stage_5__3920_,data_stage_5__3919_,data_stage_5__3918_,
  data_stage_5__3917_,data_stage_5__3916_,data_stage_5__3915_,data_stage_5__3914_,
  data_stage_5__3913_,data_stage_5__3912_,data_stage_5__3911_,data_stage_5__3910_,
  data_stage_5__3909_,data_stage_5__3908_,data_stage_5__3907_,data_stage_5__3906_,
  data_stage_5__3905_,data_stage_5__3904_,data_stage_5__3903_,data_stage_5__3902_,
  data_stage_5__3901_,data_stage_5__3900_,data_stage_5__3899_,data_stage_5__3898_,
  data_stage_5__3897_,data_stage_5__3896_,data_stage_5__3895_,data_stage_5__3894_,
  data_stage_5__3893_,data_stage_5__3892_,data_stage_5__3891_,data_stage_5__3890_,
  data_stage_5__3889_,data_stage_5__3888_,data_stage_5__3887_,data_stage_5__3886_,
  data_stage_5__3885_,data_stage_5__3884_,data_stage_5__3883_,data_stage_5__3882_,
  data_stage_5__3881_,data_stage_5__3880_,data_stage_5__3879_,data_stage_5__3878_,
  data_stage_5__3877_,data_stage_5__3876_,data_stage_5__3875_,data_stage_5__3874_,
  data_stage_5__3873_,data_stage_5__3872_,data_stage_5__3871_,data_stage_5__3870_,
  data_stage_5__3869_,data_stage_5__3868_,data_stage_5__3867_,data_stage_5__3866_,
  data_stage_5__3865_,data_stage_5__3864_,data_stage_5__3863_,data_stage_5__3862_,
  data_stage_5__3861_,data_stage_5__3860_,data_stage_5__3859_,data_stage_5__3858_,
  data_stage_5__3857_,data_stage_5__3856_,data_stage_5__3855_,data_stage_5__3854_,
  data_stage_5__3853_,data_stage_5__3852_,data_stage_5__3851_,data_stage_5__3850_,
  data_stage_5__3849_,data_stage_5__3848_,data_stage_5__3847_,data_stage_5__3846_,
  data_stage_5__3845_,data_stage_5__3844_,data_stage_5__3843_,data_stage_5__3842_,
  data_stage_5__3841_,data_stage_5__3840_,data_stage_5__3839_,data_stage_5__3838_,
  data_stage_5__3837_,data_stage_5__3836_,data_stage_5__3835_,data_stage_5__3834_,
  data_stage_5__3833_,data_stage_5__3832_,data_stage_5__3831_,data_stage_5__3830_,
  data_stage_5__3829_,data_stage_5__3828_,data_stage_5__3827_,data_stage_5__3826_,
  data_stage_5__3825_,data_stage_5__3824_,data_stage_5__3823_,data_stage_5__3822_,
  data_stage_5__3821_,data_stage_5__3820_,data_stage_5__3819_,data_stage_5__3818_,
  data_stage_5__3817_,data_stage_5__3816_,data_stage_5__3815_,data_stage_5__3814_,
  data_stage_5__3813_,data_stage_5__3812_,data_stage_5__3811_,data_stage_5__3810_,
  data_stage_5__3809_,data_stage_5__3808_,data_stage_5__3807_,data_stage_5__3806_,
  data_stage_5__3805_,data_stage_5__3804_,data_stage_5__3803_,data_stage_5__3802_,
  data_stage_5__3801_,data_stage_5__3800_,data_stage_5__3799_,data_stage_5__3798_,
  data_stage_5__3797_,data_stage_5__3796_,data_stage_5__3795_,data_stage_5__3794_,
  data_stage_5__3793_,data_stage_5__3792_,data_stage_5__3791_,data_stage_5__3790_,
  data_stage_5__3789_,data_stage_5__3788_,data_stage_5__3787_,data_stage_5__3786_,
  data_stage_5__3785_,data_stage_5__3784_,data_stage_5__3783_,data_stage_5__3782_,
  data_stage_5__3781_,data_stage_5__3780_,data_stage_5__3779_,data_stage_5__3778_,
  data_stage_5__3777_,data_stage_5__3776_,data_stage_5__3775_,data_stage_5__3774_,
  data_stage_5__3773_,data_stage_5__3772_,data_stage_5__3771_,data_stage_5__3770_,
  data_stage_5__3769_,data_stage_5__3768_,data_stage_5__3767_,data_stage_5__3766_,
  data_stage_5__3765_,data_stage_5__3764_,data_stage_5__3763_,data_stage_5__3762_,
  data_stage_5__3761_,data_stage_5__3760_,data_stage_5__3759_,data_stage_5__3758_,
  data_stage_5__3757_,data_stage_5__3756_,data_stage_5__3755_,data_stage_5__3754_,
  data_stage_5__3753_,data_stage_5__3752_,data_stage_5__3751_,data_stage_5__3750_,
  data_stage_5__3749_,data_stage_5__3748_,data_stage_5__3747_,data_stage_5__3746_,
  data_stage_5__3745_,data_stage_5__3744_,data_stage_5__3743_,data_stage_5__3742_,
  data_stage_5__3741_,data_stage_5__3740_,data_stage_5__3739_,data_stage_5__3738_,
  data_stage_5__3737_,data_stage_5__3736_,data_stage_5__3735_,data_stage_5__3734_,
  data_stage_5__3733_,data_stage_5__3732_,data_stage_5__3731_,data_stage_5__3730_,
  data_stage_5__3729_,data_stage_5__3728_,data_stage_5__3727_,data_stage_5__3726_,
  data_stage_5__3725_,data_stage_5__3724_,data_stage_5__3723_,data_stage_5__3722_,
  data_stage_5__3721_,data_stage_5__3720_,data_stage_5__3719_,data_stage_5__3718_,
  data_stage_5__3717_,data_stage_5__3716_,data_stage_5__3715_,data_stage_5__3714_,
  data_stage_5__3713_,data_stage_5__3712_,data_stage_5__3711_,data_stage_5__3710_,
  data_stage_5__3709_,data_stage_5__3708_,data_stage_5__3707_,data_stage_5__3706_,
  data_stage_5__3705_,data_stage_5__3704_,data_stage_5__3703_,data_stage_5__3702_,
  data_stage_5__3701_,data_stage_5__3700_,data_stage_5__3699_,data_stage_5__3698_,
  data_stage_5__3697_,data_stage_5__3696_,data_stage_5__3695_,data_stage_5__3694_,
  data_stage_5__3693_,data_stage_5__3692_,data_stage_5__3691_,data_stage_5__3690_,
  data_stage_5__3689_,data_stage_5__3688_,data_stage_5__3687_,data_stage_5__3686_,
  data_stage_5__3685_,data_stage_5__3684_,data_stage_5__3683_,data_stage_5__3682_,
  data_stage_5__3681_,data_stage_5__3680_,data_stage_5__3679_,data_stage_5__3678_,
  data_stage_5__3677_,data_stage_5__3676_,data_stage_5__3675_,data_stage_5__3674_,
  data_stage_5__3673_,data_stage_5__3672_,data_stage_5__3671_,data_stage_5__3670_,
  data_stage_5__3669_,data_stage_5__3668_,data_stage_5__3667_,data_stage_5__3666_,
  data_stage_5__3665_,data_stage_5__3664_,data_stage_5__3663_,data_stage_5__3662_,
  data_stage_5__3661_,data_stage_5__3660_,data_stage_5__3659_,data_stage_5__3658_,
  data_stage_5__3657_,data_stage_5__3656_,data_stage_5__3655_,data_stage_5__3654_,
  data_stage_5__3653_,data_stage_5__3652_,data_stage_5__3651_,data_stage_5__3650_,
  data_stage_5__3649_,data_stage_5__3648_,data_stage_5__3647_,data_stage_5__3646_,
  data_stage_5__3645_,data_stage_5__3644_,data_stage_5__3643_,data_stage_5__3642_,
  data_stage_5__3641_,data_stage_5__3640_,data_stage_5__3639_,data_stage_5__3638_,
  data_stage_5__3637_,data_stage_5__3636_,data_stage_5__3635_,data_stage_5__3634_,
  data_stage_5__3633_,data_stage_5__3632_,data_stage_5__3631_,data_stage_5__3630_,
  data_stage_5__3629_,data_stage_5__3628_,data_stage_5__3627_,data_stage_5__3626_,
  data_stage_5__3625_,data_stage_5__3624_,data_stage_5__3623_,data_stage_5__3622_,
  data_stage_5__3621_,data_stage_5__3620_,data_stage_5__3619_,data_stage_5__3618_,
  data_stage_5__3617_,data_stage_5__3616_,data_stage_5__3615_,data_stage_5__3614_,
  data_stage_5__3613_,data_stage_5__3612_,data_stage_5__3611_,data_stage_5__3610_,
  data_stage_5__3609_,data_stage_5__3608_,data_stage_5__3607_,data_stage_5__3606_,
  data_stage_5__3605_,data_stage_5__3604_,data_stage_5__3603_,data_stage_5__3602_,
  data_stage_5__3601_,data_stage_5__3600_,data_stage_5__3599_,data_stage_5__3598_,
  data_stage_5__3597_,data_stage_5__3596_,data_stage_5__3595_,data_stage_5__3594_,
  data_stage_5__3593_,data_stage_5__3592_,data_stage_5__3591_,data_stage_5__3590_,
  data_stage_5__3589_,data_stage_5__3588_,data_stage_5__3587_,data_stage_5__3586_,
  data_stage_5__3585_,data_stage_5__3584_,data_stage_5__3583_,data_stage_5__3582_,
  data_stage_5__3581_,data_stage_5__3580_,data_stage_5__3579_,data_stage_5__3578_,
  data_stage_5__3577_,data_stage_5__3576_,data_stage_5__3575_,data_stage_5__3574_,
  data_stage_5__3573_,data_stage_5__3572_,data_stage_5__3571_,data_stage_5__3570_,
  data_stage_5__3569_,data_stage_5__3568_,data_stage_5__3567_,data_stage_5__3566_,
  data_stage_5__3565_,data_stage_5__3564_,data_stage_5__3563_,data_stage_5__3562_,
  data_stage_5__3561_,data_stage_5__3560_,data_stage_5__3559_,data_stage_5__3558_,
  data_stage_5__3557_,data_stage_5__3556_,data_stage_5__3555_,data_stage_5__3554_,
  data_stage_5__3553_,data_stage_5__3552_,data_stage_5__3551_,data_stage_5__3550_,
  data_stage_5__3549_,data_stage_5__3548_,data_stage_5__3547_,data_stage_5__3546_,
  data_stage_5__3545_,data_stage_5__3544_,data_stage_5__3543_,data_stage_5__3542_,
  data_stage_5__3541_,data_stage_5__3540_,data_stage_5__3539_,data_stage_5__3538_,
  data_stage_5__3537_,data_stage_5__3536_,data_stage_5__3535_,data_stage_5__3534_,
  data_stage_5__3533_,data_stage_5__3532_,data_stage_5__3531_,data_stage_5__3530_,
  data_stage_5__3529_,data_stage_5__3528_,data_stage_5__3527_,data_stage_5__3526_,
  data_stage_5__3525_,data_stage_5__3524_,data_stage_5__3523_,data_stage_5__3522_,
  data_stage_5__3521_,data_stage_5__3520_,data_stage_5__3519_,data_stage_5__3518_,
  data_stage_5__3517_,data_stage_5__3516_,data_stage_5__3515_,data_stage_5__3514_,
  data_stage_5__3513_,data_stage_5__3512_,data_stage_5__3511_,data_stage_5__3510_,
  data_stage_5__3509_,data_stage_5__3508_,data_stage_5__3507_,data_stage_5__3506_,
  data_stage_5__3505_,data_stage_5__3504_,data_stage_5__3503_,data_stage_5__3502_,
  data_stage_5__3501_,data_stage_5__3500_,data_stage_5__3499_,data_stage_5__3498_,
  data_stage_5__3497_,data_stage_5__3496_,data_stage_5__3495_,data_stage_5__3494_,
  data_stage_5__3493_,data_stage_5__3492_,data_stage_5__3491_,data_stage_5__3490_,
  data_stage_5__3489_,data_stage_5__3488_,data_stage_5__3487_,data_stage_5__3486_,
  data_stage_5__3485_,data_stage_5__3484_,data_stage_5__3483_,data_stage_5__3482_,
  data_stage_5__3481_,data_stage_5__3480_,data_stage_5__3479_,data_stage_5__3478_,
  data_stage_5__3477_,data_stage_5__3476_,data_stage_5__3475_,data_stage_5__3474_,
  data_stage_5__3473_,data_stage_5__3472_,data_stage_5__3471_,data_stage_5__3470_,
  data_stage_5__3469_,data_stage_5__3468_,data_stage_5__3467_,data_stage_5__3466_,
  data_stage_5__3465_,data_stage_5__3464_,data_stage_5__3463_,data_stage_5__3462_,
  data_stage_5__3461_,data_stage_5__3460_,data_stage_5__3459_,data_stage_5__3458_,
  data_stage_5__3457_,data_stage_5__3456_,data_stage_5__3455_,data_stage_5__3454_,
  data_stage_5__3453_,data_stage_5__3452_,data_stage_5__3451_,data_stage_5__3450_,
  data_stage_5__3449_,data_stage_5__3448_,data_stage_5__3447_,data_stage_5__3446_,
  data_stage_5__3445_,data_stage_5__3444_,data_stage_5__3443_,data_stage_5__3442_,
  data_stage_5__3441_,data_stage_5__3440_,data_stage_5__3439_,data_stage_5__3438_,
  data_stage_5__3437_,data_stage_5__3436_,data_stage_5__3435_,data_stage_5__3434_,
  data_stage_5__3433_,data_stage_5__3432_,data_stage_5__3431_,data_stage_5__3430_,
  data_stage_5__3429_,data_stage_5__3428_,data_stage_5__3427_,data_stage_5__3426_,
  data_stage_5__3425_,data_stage_5__3424_,data_stage_5__3423_,data_stage_5__3422_,
  data_stage_5__3421_,data_stage_5__3420_,data_stage_5__3419_,data_stage_5__3418_,
  data_stage_5__3417_,data_stage_5__3416_,data_stage_5__3415_,data_stage_5__3414_,
  data_stage_5__3413_,data_stage_5__3412_,data_stage_5__3411_,data_stage_5__3410_,
  data_stage_5__3409_,data_stage_5__3408_,data_stage_5__3407_,data_stage_5__3406_,
  data_stage_5__3405_,data_stage_5__3404_,data_stage_5__3403_,data_stage_5__3402_,
  data_stage_5__3401_,data_stage_5__3400_,data_stage_5__3399_,data_stage_5__3398_,
  data_stage_5__3397_,data_stage_5__3396_,data_stage_5__3395_,data_stage_5__3394_,
  data_stage_5__3393_,data_stage_5__3392_,data_stage_5__3391_,data_stage_5__3390_,
  data_stage_5__3389_,data_stage_5__3388_,data_stage_5__3387_,data_stage_5__3386_,
  data_stage_5__3385_,data_stage_5__3384_,data_stage_5__3383_,data_stage_5__3382_,
  data_stage_5__3381_,data_stage_5__3380_,data_stage_5__3379_,data_stage_5__3378_,
  data_stage_5__3377_,data_stage_5__3376_,data_stage_5__3375_,data_stage_5__3374_,
  data_stage_5__3373_,data_stage_5__3372_,data_stage_5__3371_,data_stage_5__3370_,
  data_stage_5__3369_,data_stage_5__3368_,data_stage_5__3367_,data_stage_5__3366_,
  data_stage_5__3365_,data_stage_5__3364_,data_stage_5__3363_,data_stage_5__3362_,
  data_stage_5__3361_,data_stage_5__3360_,data_stage_5__3359_,data_stage_5__3358_,
  data_stage_5__3357_,data_stage_5__3356_,data_stage_5__3355_,data_stage_5__3354_,
  data_stage_5__3353_,data_stage_5__3352_,data_stage_5__3351_,data_stage_5__3350_,
  data_stage_5__3349_,data_stage_5__3348_,data_stage_5__3347_,data_stage_5__3346_,
  data_stage_5__3345_,data_stage_5__3344_,data_stage_5__3343_,data_stage_5__3342_,
  data_stage_5__3341_,data_stage_5__3340_,data_stage_5__3339_,data_stage_5__3338_,
  data_stage_5__3337_,data_stage_5__3336_,data_stage_5__3335_,data_stage_5__3334_,
  data_stage_5__3333_,data_stage_5__3332_,data_stage_5__3331_,data_stage_5__3330_,
  data_stage_5__3329_,data_stage_5__3328_,data_stage_5__3327_,data_stage_5__3326_,
  data_stage_5__3325_,data_stage_5__3324_,data_stage_5__3323_,data_stage_5__3322_,
  data_stage_5__3321_,data_stage_5__3320_,data_stage_5__3319_,data_stage_5__3318_,
  data_stage_5__3317_,data_stage_5__3316_,data_stage_5__3315_,data_stage_5__3314_,
  data_stage_5__3313_,data_stage_5__3312_,data_stage_5__3311_,data_stage_5__3310_,
  data_stage_5__3309_,data_stage_5__3308_,data_stage_5__3307_,data_stage_5__3306_,
  data_stage_5__3305_,data_stage_5__3304_,data_stage_5__3303_,data_stage_5__3302_,
  data_stage_5__3301_,data_stage_5__3300_,data_stage_5__3299_,data_stage_5__3298_,
  data_stage_5__3297_,data_stage_5__3296_,data_stage_5__3295_,data_stage_5__3294_,
  data_stage_5__3293_,data_stage_5__3292_,data_stage_5__3291_,data_stage_5__3290_,
  data_stage_5__3289_,data_stage_5__3288_,data_stage_5__3287_,data_stage_5__3286_,
  data_stage_5__3285_,data_stage_5__3284_,data_stage_5__3283_,data_stage_5__3282_,
  data_stage_5__3281_,data_stage_5__3280_,data_stage_5__3279_,data_stage_5__3278_,
  data_stage_5__3277_,data_stage_5__3276_,data_stage_5__3275_,data_stage_5__3274_,
  data_stage_5__3273_,data_stage_5__3272_,data_stage_5__3271_,data_stage_5__3270_,
  data_stage_5__3269_,data_stage_5__3268_,data_stage_5__3267_,data_stage_5__3266_,
  data_stage_5__3265_,data_stage_5__3264_,data_stage_5__3263_,data_stage_5__3262_,
  data_stage_5__3261_,data_stage_5__3260_,data_stage_5__3259_,data_stage_5__3258_,
  data_stage_5__3257_,data_stage_5__3256_,data_stage_5__3255_,data_stage_5__3254_,
  data_stage_5__3253_,data_stage_5__3252_,data_stage_5__3251_,data_stage_5__3250_,
  data_stage_5__3249_,data_stage_5__3248_,data_stage_5__3247_,data_stage_5__3246_,
  data_stage_5__3245_,data_stage_5__3244_,data_stage_5__3243_,data_stage_5__3242_,
  data_stage_5__3241_,data_stage_5__3240_,data_stage_5__3239_,data_stage_5__3238_,
  data_stage_5__3237_,data_stage_5__3236_,data_stage_5__3235_,data_stage_5__3234_,
  data_stage_5__3233_,data_stage_5__3232_,data_stage_5__3231_,data_stage_5__3230_,
  data_stage_5__3229_,data_stage_5__3228_,data_stage_5__3227_,data_stage_5__3226_,
  data_stage_5__3225_,data_stage_5__3224_,data_stage_5__3223_,data_stage_5__3222_,
  data_stage_5__3221_,data_stage_5__3220_,data_stage_5__3219_,data_stage_5__3218_,
  data_stage_5__3217_,data_stage_5__3216_,data_stage_5__3215_,data_stage_5__3214_,
  data_stage_5__3213_,data_stage_5__3212_,data_stage_5__3211_,data_stage_5__3210_,
  data_stage_5__3209_,data_stage_5__3208_,data_stage_5__3207_,data_stage_5__3206_,
  data_stage_5__3205_,data_stage_5__3204_,data_stage_5__3203_,data_stage_5__3202_,
  data_stage_5__3201_,data_stage_5__3200_,data_stage_5__3199_,data_stage_5__3198_,
  data_stage_5__3197_,data_stage_5__3196_,data_stage_5__3195_,data_stage_5__3194_,
  data_stage_5__3193_,data_stage_5__3192_,data_stage_5__3191_,data_stage_5__3190_,
  data_stage_5__3189_,data_stage_5__3188_,data_stage_5__3187_,data_stage_5__3186_,
  data_stage_5__3185_,data_stage_5__3184_,data_stage_5__3183_,data_stage_5__3182_,
  data_stage_5__3181_,data_stage_5__3180_,data_stage_5__3179_,data_stage_5__3178_,
  data_stage_5__3177_,data_stage_5__3176_,data_stage_5__3175_,data_stage_5__3174_,
  data_stage_5__3173_,data_stage_5__3172_,data_stage_5__3171_,data_stage_5__3170_,
  data_stage_5__3169_,data_stage_5__3168_,data_stage_5__3167_,data_stage_5__3166_,
  data_stage_5__3165_,data_stage_5__3164_,data_stage_5__3163_,data_stage_5__3162_,
  data_stage_5__3161_,data_stage_5__3160_,data_stage_5__3159_,data_stage_5__3158_,
  data_stage_5__3157_,data_stage_5__3156_,data_stage_5__3155_,data_stage_5__3154_,
  data_stage_5__3153_,data_stage_5__3152_,data_stage_5__3151_,data_stage_5__3150_,
  data_stage_5__3149_,data_stage_5__3148_,data_stage_5__3147_,data_stage_5__3146_,
  data_stage_5__3145_,data_stage_5__3144_,data_stage_5__3143_,data_stage_5__3142_,
  data_stage_5__3141_,data_stage_5__3140_,data_stage_5__3139_,data_stage_5__3138_,
  data_stage_5__3137_,data_stage_5__3136_,data_stage_5__3135_,data_stage_5__3134_,
  data_stage_5__3133_,data_stage_5__3132_,data_stage_5__3131_,data_stage_5__3130_,
  data_stage_5__3129_,data_stage_5__3128_,data_stage_5__3127_,data_stage_5__3126_,
  data_stage_5__3125_,data_stage_5__3124_,data_stage_5__3123_,data_stage_5__3122_,
  data_stage_5__3121_,data_stage_5__3120_,data_stage_5__3119_,data_stage_5__3118_,
  data_stage_5__3117_,data_stage_5__3116_,data_stage_5__3115_,data_stage_5__3114_,
  data_stage_5__3113_,data_stage_5__3112_,data_stage_5__3111_,data_stage_5__3110_,
  data_stage_5__3109_,data_stage_5__3108_,data_stage_5__3107_,data_stage_5__3106_,
  data_stage_5__3105_,data_stage_5__3104_,data_stage_5__3103_,data_stage_5__3102_,
  data_stage_5__3101_,data_stage_5__3100_,data_stage_5__3099_,data_stage_5__3098_,
  data_stage_5__3097_,data_stage_5__3096_,data_stage_5__3095_,data_stage_5__3094_,
  data_stage_5__3093_,data_stage_5__3092_,data_stage_5__3091_,data_stage_5__3090_,
  data_stage_5__3089_,data_stage_5__3088_,data_stage_5__3087_,data_stage_5__3086_,
  data_stage_5__3085_,data_stage_5__3084_,data_stage_5__3083_,data_stage_5__3082_,
  data_stage_5__3081_,data_stage_5__3080_,data_stage_5__3079_,data_stage_5__3078_,
  data_stage_5__3077_,data_stage_5__3076_,data_stage_5__3075_,data_stage_5__3074_,
  data_stage_5__3073_,data_stage_5__3072_,data_stage_5__3071_,data_stage_5__3070_,
  data_stage_5__3069_,data_stage_5__3068_,data_stage_5__3067_,data_stage_5__3066_,
  data_stage_5__3065_,data_stage_5__3064_,data_stage_5__3063_,data_stage_5__3062_,
  data_stage_5__3061_,data_stage_5__3060_,data_stage_5__3059_,data_stage_5__3058_,
  data_stage_5__3057_,data_stage_5__3056_,data_stage_5__3055_,data_stage_5__3054_,
  data_stage_5__3053_,data_stage_5__3052_,data_stage_5__3051_,data_stage_5__3050_,
  data_stage_5__3049_,data_stage_5__3048_,data_stage_5__3047_,data_stage_5__3046_,
  data_stage_5__3045_,data_stage_5__3044_,data_stage_5__3043_,data_stage_5__3042_,
  data_stage_5__3041_,data_stage_5__3040_,data_stage_5__3039_,data_stage_5__3038_,
  data_stage_5__3037_,data_stage_5__3036_,data_stage_5__3035_,data_stage_5__3034_,
  data_stage_5__3033_,data_stage_5__3032_,data_stage_5__3031_,data_stage_5__3030_,
  data_stage_5__3029_,data_stage_5__3028_,data_stage_5__3027_,data_stage_5__3026_,
  data_stage_5__3025_,data_stage_5__3024_,data_stage_5__3023_,data_stage_5__3022_,
  data_stage_5__3021_,data_stage_5__3020_,data_stage_5__3019_,data_stage_5__3018_,
  data_stage_5__3017_,data_stage_5__3016_,data_stage_5__3015_,data_stage_5__3014_,
  data_stage_5__3013_,data_stage_5__3012_,data_stage_5__3011_,data_stage_5__3010_,
  data_stage_5__3009_,data_stage_5__3008_,data_stage_5__3007_,data_stage_5__3006_,
  data_stage_5__3005_,data_stage_5__3004_,data_stage_5__3003_,data_stage_5__3002_,
  data_stage_5__3001_,data_stage_5__3000_,data_stage_5__2999_,data_stage_5__2998_,
  data_stage_5__2997_,data_stage_5__2996_,data_stage_5__2995_,data_stage_5__2994_,
  data_stage_5__2993_,data_stage_5__2992_,data_stage_5__2991_,data_stage_5__2990_,
  data_stage_5__2989_,data_stage_5__2988_,data_stage_5__2987_,data_stage_5__2986_,
  data_stage_5__2985_,data_stage_5__2984_,data_stage_5__2983_,data_stage_5__2982_,
  data_stage_5__2981_,data_stage_5__2980_,data_stage_5__2979_,data_stage_5__2978_,
  data_stage_5__2977_,data_stage_5__2976_,data_stage_5__2975_,data_stage_5__2974_,
  data_stage_5__2973_,data_stage_5__2972_,data_stage_5__2971_,data_stage_5__2970_,
  data_stage_5__2969_,data_stage_5__2968_,data_stage_5__2967_,data_stage_5__2966_,
  data_stage_5__2965_,data_stage_5__2964_,data_stage_5__2963_,data_stage_5__2962_,
  data_stage_5__2961_,data_stage_5__2960_,data_stage_5__2959_,data_stage_5__2958_,
  data_stage_5__2957_,data_stage_5__2956_,data_stage_5__2955_,data_stage_5__2954_,
  data_stage_5__2953_,data_stage_5__2952_,data_stage_5__2951_,data_stage_5__2950_,
  data_stage_5__2949_,data_stage_5__2948_,data_stage_5__2947_,data_stage_5__2946_,
  data_stage_5__2945_,data_stage_5__2944_,data_stage_5__2943_,data_stage_5__2942_,
  data_stage_5__2941_,data_stage_5__2940_,data_stage_5__2939_,data_stage_5__2938_,
  data_stage_5__2937_,data_stage_5__2936_,data_stage_5__2935_,data_stage_5__2934_,
  data_stage_5__2933_,data_stage_5__2932_,data_stage_5__2931_,data_stage_5__2930_,
  data_stage_5__2929_,data_stage_5__2928_,data_stage_5__2927_,data_stage_5__2926_,
  data_stage_5__2925_,data_stage_5__2924_,data_stage_5__2923_,data_stage_5__2922_,
  data_stage_5__2921_,data_stage_5__2920_,data_stage_5__2919_,data_stage_5__2918_,
  data_stage_5__2917_,data_stage_5__2916_,data_stage_5__2915_,data_stage_5__2914_,
  data_stage_5__2913_,data_stage_5__2912_,data_stage_5__2911_,data_stage_5__2910_,
  data_stage_5__2909_,data_stage_5__2908_,data_stage_5__2907_,data_stage_5__2906_,
  data_stage_5__2905_,data_stage_5__2904_,data_stage_5__2903_,data_stage_5__2902_,
  data_stage_5__2901_,data_stage_5__2900_,data_stage_5__2899_,data_stage_5__2898_,
  data_stage_5__2897_,data_stage_5__2896_,data_stage_5__2895_,data_stage_5__2894_,
  data_stage_5__2893_,data_stage_5__2892_,data_stage_5__2891_,data_stage_5__2890_,
  data_stage_5__2889_,data_stage_5__2888_,data_stage_5__2887_,data_stage_5__2886_,
  data_stage_5__2885_,data_stage_5__2884_,data_stage_5__2883_,data_stage_5__2882_,
  data_stage_5__2881_,data_stage_5__2880_,data_stage_5__2879_,data_stage_5__2878_,
  data_stage_5__2877_,data_stage_5__2876_,data_stage_5__2875_,data_stage_5__2874_,
  data_stage_5__2873_,data_stage_5__2872_,data_stage_5__2871_,data_stage_5__2870_,
  data_stage_5__2869_,data_stage_5__2868_,data_stage_5__2867_,data_stage_5__2866_,
  data_stage_5__2865_,data_stage_5__2864_,data_stage_5__2863_,data_stage_5__2862_,
  data_stage_5__2861_,data_stage_5__2860_,data_stage_5__2859_,data_stage_5__2858_,
  data_stage_5__2857_,data_stage_5__2856_,data_stage_5__2855_,data_stage_5__2854_,
  data_stage_5__2853_,data_stage_5__2852_,data_stage_5__2851_,data_stage_5__2850_,
  data_stage_5__2849_,data_stage_5__2848_,data_stage_5__2847_,data_stage_5__2846_,
  data_stage_5__2845_,data_stage_5__2844_,data_stage_5__2843_,data_stage_5__2842_,
  data_stage_5__2841_,data_stage_5__2840_,data_stage_5__2839_,data_stage_5__2838_,
  data_stage_5__2837_,data_stage_5__2836_,data_stage_5__2835_,data_stage_5__2834_,
  data_stage_5__2833_,data_stage_5__2832_,data_stage_5__2831_,data_stage_5__2830_,
  data_stage_5__2829_,data_stage_5__2828_,data_stage_5__2827_,data_stage_5__2826_,
  data_stage_5__2825_,data_stage_5__2824_,data_stage_5__2823_,data_stage_5__2822_,
  data_stage_5__2821_,data_stage_5__2820_,data_stage_5__2819_,data_stage_5__2818_,
  data_stage_5__2817_,data_stage_5__2816_,data_stage_5__2815_,data_stage_5__2814_,
  data_stage_5__2813_,data_stage_5__2812_,data_stage_5__2811_,data_stage_5__2810_,
  data_stage_5__2809_,data_stage_5__2808_,data_stage_5__2807_,data_stage_5__2806_,
  data_stage_5__2805_,data_stage_5__2804_,data_stage_5__2803_,data_stage_5__2802_,
  data_stage_5__2801_,data_stage_5__2800_,data_stage_5__2799_,data_stage_5__2798_,
  data_stage_5__2797_,data_stage_5__2796_,data_stage_5__2795_,data_stage_5__2794_,
  data_stage_5__2793_,data_stage_5__2792_,data_stage_5__2791_,data_stage_5__2790_,
  data_stage_5__2789_,data_stage_5__2788_,data_stage_5__2787_,data_stage_5__2786_,
  data_stage_5__2785_,data_stage_5__2784_,data_stage_5__2783_,data_stage_5__2782_,
  data_stage_5__2781_,data_stage_5__2780_,data_stage_5__2779_,data_stage_5__2778_,
  data_stage_5__2777_,data_stage_5__2776_,data_stage_5__2775_,data_stage_5__2774_,
  data_stage_5__2773_,data_stage_5__2772_,data_stage_5__2771_,data_stage_5__2770_,
  data_stage_5__2769_,data_stage_5__2768_,data_stage_5__2767_,data_stage_5__2766_,
  data_stage_5__2765_,data_stage_5__2764_,data_stage_5__2763_,data_stage_5__2762_,
  data_stage_5__2761_,data_stage_5__2760_,data_stage_5__2759_,data_stage_5__2758_,
  data_stage_5__2757_,data_stage_5__2756_,data_stage_5__2755_,data_stage_5__2754_,
  data_stage_5__2753_,data_stage_5__2752_,data_stage_5__2751_,data_stage_5__2750_,
  data_stage_5__2749_,data_stage_5__2748_,data_stage_5__2747_,data_stage_5__2746_,
  data_stage_5__2745_,data_stage_5__2744_,data_stage_5__2743_,data_stage_5__2742_,
  data_stage_5__2741_,data_stage_5__2740_,data_stage_5__2739_,data_stage_5__2738_,
  data_stage_5__2737_,data_stage_5__2736_,data_stage_5__2735_,data_stage_5__2734_,
  data_stage_5__2733_,data_stage_5__2732_,data_stage_5__2731_,data_stage_5__2730_,
  data_stage_5__2729_,data_stage_5__2728_,data_stage_5__2727_,data_stage_5__2726_,
  data_stage_5__2725_,data_stage_5__2724_,data_stage_5__2723_,data_stage_5__2722_,
  data_stage_5__2721_,data_stage_5__2720_,data_stage_5__2719_,data_stage_5__2718_,
  data_stage_5__2717_,data_stage_5__2716_,data_stage_5__2715_,data_stage_5__2714_,
  data_stage_5__2713_,data_stage_5__2712_,data_stage_5__2711_,data_stage_5__2710_,
  data_stage_5__2709_,data_stage_5__2708_,data_stage_5__2707_,data_stage_5__2706_,
  data_stage_5__2705_,data_stage_5__2704_,data_stage_5__2703_,data_stage_5__2702_,
  data_stage_5__2701_,data_stage_5__2700_,data_stage_5__2699_,data_stage_5__2698_,
  data_stage_5__2697_,data_stage_5__2696_,data_stage_5__2695_,data_stage_5__2694_,
  data_stage_5__2693_,data_stage_5__2692_,data_stage_5__2691_,data_stage_5__2690_,
  data_stage_5__2689_,data_stage_5__2688_,data_stage_5__2687_,data_stage_5__2686_,
  data_stage_5__2685_,data_stage_5__2684_,data_stage_5__2683_,data_stage_5__2682_,
  data_stage_5__2681_,data_stage_5__2680_,data_stage_5__2679_,data_stage_5__2678_,
  data_stage_5__2677_,data_stage_5__2676_,data_stage_5__2675_,data_stage_5__2674_,
  data_stage_5__2673_,data_stage_5__2672_,data_stage_5__2671_,data_stage_5__2670_,
  data_stage_5__2669_,data_stage_5__2668_,data_stage_5__2667_,data_stage_5__2666_,
  data_stage_5__2665_,data_stage_5__2664_,data_stage_5__2663_,data_stage_5__2662_,
  data_stage_5__2661_,data_stage_5__2660_,data_stage_5__2659_,data_stage_5__2658_,
  data_stage_5__2657_,data_stage_5__2656_,data_stage_5__2655_,data_stage_5__2654_,
  data_stage_5__2653_,data_stage_5__2652_,data_stage_5__2651_,data_stage_5__2650_,
  data_stage_5__2649_,data_stage_5__2648_,data_stage_5__2647_,data_stage_5__2646_,
  data_stage_5__2645_,data_stage_5__2644_,data_stage_5__2643_,data_stage_5__2642_,
  data_stage_5__2641_,data_stage_5__2640_,data_stage_5__2639_,data_stage_5__2638_,
  data_stage_5__2637_,data_stage_5__2636_,data_stage_5__2635_,data_stage_5__2634_,
  data_stage_5__2633_,data_stage_5__2632_,data_stage_5__2631_,data_stage_5__2630_,
  data_stage_5__2629_,data_stage_5__2628_,data_stage_5__2627_,data_stage_5__2626_,
  data_stage_5__2625_,data_stage_5__2624_,data_stage_5__2623_,data_stage_5__2622_,
  data_stage_5__2621_,data_stage_5__2620_,data_stage_5__2619_,data_stage_5__2618_,
  data_stage_5__2617_,data_stage_5__2616_,data_stage_5__2615_,data_stage_5__2614_,
  data_stage_5__2613_,data_stage_5__2612_,data_stage_5__2611_,data_stage_5__2610_,
  data_stage_5__2609_,data_stage_5__2608_,data_stage_5__2607_,data_stage_5__2606_,
  data_stage_5__2605_,data_stage_5__2604_,data_stage_5__2603_,data_stage_5__2602_,
  data_stage_5__2601_,data_stage_5__2600_,data_stage_5__2599_,data_stage_5__2598_,
  data_stage_5__2597_,data_stage_5__2596_,data_stage_5__2595_,data_stage_5__2594_,
  data_stage_5__2593_,data_stage_5__2592_,data_stage_5__2591_,data_stage_5__2590_,
  data_stage_5__2589_,data_stage_5__2588_,data_stage_5__2587_,data_stage_5__2586_,
  data_stage_5__2585_,data_stage_5__2584_,data_stage_5__2583_,data_stage_5__2582_,
  data_stage_5__2581_,data_stage_5__2580_,data_stage_5__2579_,data_stage_5__2578_,
  data_stage_5__2577_,data_stage_5__2576_,data_stage_5__2575_,data_stage_5__2574_,
  data_stage_5__2573_,data_stage_5__2572_,data_stage_5__2571_,data_stage_5__2570_,
  data_stage_5__2569_,data_stage_5__2568_,data_stage_5__2567_,data_stage_5__2566_,
  data_stage_5__2565_,data_stage_5__2564_,data_stage_5__2563_,data_stage_5__2562_,
  data_stage_5__2561_,data_stage_5__2560_,data_stage_5__2559_,data_stage_5__2558_,
  data_stage_5__2557_,data_stage_5__2556_,data_stage_5__2555_,data_stage_5__2554_,
  data_stage_5__2553_,data_stage_5__2552_,data_stage_5__2551_,data_stage_5__2550_,
  data_stage_5__2549_,data_stage_5__2548_,data_stage_5__2547_,data_stage_5__2546_,
  data_stage_5__2545_,data_stage_5__2544_,data_stage_5__2543_,data_stage_5__2542_,
  data_stage_5__2541_,data_stage_5__2540_,data_stage_5__2539_,data_stage_5__2538_,
  data_stage_5__2537_,data_stage_5__2536_,data_stage_5__2535_,data_stage_5__2534_,
  data_stage_5__2533_,data_stage_5__2532_,data_stage_5__2531_,data_stage_5__2530_,
  data_stage_5__2529_,data_stage_5__2528_,data_stage_5__2527_,data_stage_5__2526_,
  data_stage_5__2525_,data_stage_5__2524_,data_stage_5__2523_,data_stage_5__2522_,
  data_stage_5__2521_,data_stage_5__2520_,data_stage_5__2519_,data_stage_5__2518_,
  data_stage_5__2517_,data_stage_5__2516_,data_stage_5__2515_,data_stage_5__2514_,
  data_stage_5__2513_,data_stage_5__2512_,data_stage_5__2511_,data_stage_5__2510_,
  data_stage_5__2509_,data_stage_5__2508_,data_stage_5__2507_,data_stage_5__2506_,
  data_stage_5__2505_,data_stage_5__2504_,data_stage_5__2503_,data_stage_5__2502_,
  data_stage_5__2501_,data_stage_5__2500_,data_stage_5__2499_,data_stage_5__2498_,
  data_stage_5__2497_,data_stage_5__2496_,data_stage_5__2495_,data_stage_5__2494_,
  data_stage_5__2493_,data_stage_5__2492_,data_stage_5__2491_,data_stage_5__2490_,
  data_stage_5__2489_,data_stage_5__2488_,data_stage_5__2487_,data_stage_5__2486_,
  data_stage_5__2485_,data_stage_5__2484_,data_stage_5__2483_,data_stage_5__2482_,
  data_stage_5__2481_,data_stage_5__2480_,data_stage_5__2479_,data_stage_5__2478_,
  data_stage_5__2477_,data_stage_5__2476_,data_stage_5__2475_,data_stage_5__2474_,
  data_stage_5__2473_,data_stage_5__2472_,data_stage_5__2471_,data_stage_5__2470_,
  data_stage_5__2469_,data_stage_5__2468_,data_stage_5__2467_,data_stage_5__2466_,
  data_stage_5__2465_,data_stage_5__2464_,data_stage_5__2463_,data_stage_5__2462_,
  data_stage_5__2461_,data_stage_5__2460_,data_stage_5__2459_,data_stage_5__2458_,
  data_stage_5__2457_,data_stage_5__2456_,data_stage_5__2455_,data_stage_5__2454_,
  data_stage_5__2453_,data_stage_5__2452_,data_stage_5__2451_,data_stage_5__2450_,
  data_stage_5__2449_,data_stage_5__2448_,data_stage_5__2447_,data_stage_5__2446_,
  data_stage_5__2445_,data_stage_5__2444_,data_stage_5__2443_,data_stage_5__2442_,
  data_stage_5__2441_,data_stage_5__2440_,data_stage_5__2439_,data_stage_5__2438_,
  data_stage_5__2437_,data_stage_5__2436_,data_stage_5__2435_,data_stage_5__2434_,
  data_stage_5__2433_,data_stage_5__2432_,data_stage_5__2431_,data_stage_5__2430_,
  data_stage_5__2429_,data_stage_5__2428_,data_stage_5__2427_,data_stage_5__2426_,
  data_stage_5__2425_,data_stage_5__2424_,data_stage_5__2423_,data_stage_5__2422_,
  data_stage_5__2421_,data_stage_5__2420_,data_stage_5__2419_,data_stage_5__2418_,
  data_stage_5__2417_,data_stage_5__2416_,data_stage_5__2415_,data_stage_5__2414_,
  data_stage_5__2413_,data_stage_5__2412_,data_stage_5__2411_,data_stage_5__2410_,
  data_stage_5__2409_,data_stage_5__2408_,data_stage_5__2407_,data_stage_5__2406_,
  data_stage_5__2405_,data_stage_5__2404_,data_stage_5__2403_,data_stage_5__2402_,
  data_stage_5__2401_,data_stage_5__2400_,data_stage_5__2399_,data_stage_5__2398_,
  data_stage_5__2397_,data_stage_5__2396_,data_stage_5__2395_,data_stage_5__2394_,
  data_stage_5__2393_,data_stage_5__2392_,data_stage_5__2391_,data_stage_5__2390_,
  data_stage_5__2389_,data_stage_5__2388_,data_stage_5__2387_,data_stage_5__2386_,
  data_stage_5__2385_,data_stage_5__2384_,data_stage_5__2383_,data_stage_5__2382_,
  data_stage_5__2381_,data_stage_5__2380_,data_stage_5__2379_,data_stage_5__2378_,
  data_stage_5__2377_,data_stage_5__2376_,data_stage_5__2375_,data_stage_5__2374_,
  data_stage_5__2373_,data_stage_5__2372_,data_stage_5__2371_,data_stage_5__2370_,
  data_stage_5__2369_,data_stage_5__2368_,data_stage_5__2367_,data_stage_5__2366_,
  data_stage_5__2365_,data_stage_5__2364_,data_stage_5__2363_,data_stage_5__2362_,
  data_stage_5__2361_,data_stage_5__2360_,data_stage_5__2359_,data_stage_5__2358_,
  data_stage_5__2357_,data_stage_5__2356_,data_stage_5__2355_,data_stage_5__2354_,
  data_stage_5__2353_,data_stage_5__2352_,data_stage_5__2351_,data_stage_5__2350_,
  data_stage_5__2349_,data_stage_5__2348_,data_stage_5__2347_,data_stage_5__2346_,
  data_stage_5__2345_,data_stage_5__2344_,data_stage_5__2343_,data_stage_5__2342_,
  data_stage_5__2341_,data_stage_5__2340_,data_stage_5__2339_,data_stage_5__2338_,
  data_stage_5__2337_,data_stage_5__2336_,data_stage_5__2335_,data_stage_5__2334_,
  data_stage_5__2333_,data_stage_5__2332_,data_stage_5__2331_,data_stage_5__2330_,
  data_stage_5__2329_,data_stage_5__2328_,data_stage_5__2327_,data_stage_5__2326_,
  data_stage_5__2325_,data_stage_5__2324_,data_stage_5__2323_,data_stage_5__2322_,
  data_stage_5__2321_,data_stage_5__2320_,data_stage_5__2319_,data_stage_5__2318_,
  data_stage_5__2317_,data_stage_5__2316_,data_stage_5__2315_,data_stage_5__2314_,
  data_stage_5__2313_,data_stage_5__2312_,data_stage_5__2311_,data_stage_5__2310_,
  data_stage_5__2309_,data_stage_5__2308_,data_stage_5__2307_,data_stage_5__2306_,
  data_stage_5__2305_,data_stage_5__2304_,data_stage_5__2303_,data_stage_5__2302_,
  data_stage_5__2301_,data_stage_5__2300_,data_stage_5__2299_,data_stage_5__2298_,
  data_stage_5__2297_,data_stage_5__2296_,data_stage_5__2295_,data_stage_5__2294_,
  data_stage_5__2293_,data_stage_5__2292_,data_stage_5__2291_,data_stage_5__2290_,
  data_stage_5__2289_,data_stage_5__2288_,data_stage_5__2287_,data_stage_5__2286_,
  data_stage_5__2285_,data_stage_5__2284_,data_stage_5__2283_,data_stage_5__2282_,
  data_stage_5__2281_,data_stage_5__2280_,data_stage_5__2279_,data_stage_5__2278_,
  data_stage_5__2277_,data_stage_5__2276_,data_stage_5__2275_,data_stage_5__2274_,
  data_stage_5__2273_,data_stage_5__2272_,data_stage_5__2271_,data_stage_5__2270_,
  data_stage_5__2269_,data_stage_5__2268_,data_stage_5__2267_,data_stage_5__2266_,
  data_stage_5__2265_,data_stage_5__2264_,data_stage_5__2263_,data_stage_5__2262_,
  data_stage_5__2261_,data_stage_5__2260_,data_stage_5__2259_,data_stage_5__2258_,
  data_stage_5__2257_,data_stage_5__2256_,data_stage_5__2255_,data_stage_5__2254_,
  data_stage_5__2253_,data_stage_5__2252_,data_stage_5__2251_,data_stage_5__2250_,
  data_stage_5__2249_,data_stage_5__2248_,data_stage_5__2247_,data_stage_5__2246_,
  data_stage_5__2245_,data_stage_5__2244_,data_stage_5__2243_,data_stage_5__2242_,
  data_stage_5__2241_,data_stage_5__2240_,data_stage_5__2239_,data_stage_5__2238_,
  data_stage_5__2237_,data_stage_5__2236_,data_stage_5__2235_,data_stage_5__2234_,
  data_stage_5__2233_,data_stage_5__2232_,data_stage_5__2231_,data_stage_5__2230_,
  data_stage_5__2229_,data_stage_5__2228_,data_stage_5__2227_,data_stage_5__2226_,
  data_stage_5__2225_,data_stage_5__2224_,data_stage_5__2223_,data_stage_5__2222_,
  data_stage_5__2221_,data_stage_5__2220_,data_stage_5__2219_,data_stage_5__2218_,
  data_stage_5__2217_,data_stage_5__2216_,data_stage_5__2215_,data_stage_5__2214_,
  data_stage_5__2213_,data_stage_5__2212_,data_stage_5__2211_,data_stage_5__2210_,
  data_stage_5__2209_,data_stage_5__2208_,data_stage_5__2207_,data_stage_5__2206_,
  data_stage_5__2205_,data_stage_5__2204_,data_stage_5__2203_,data_stage_5__2202_,
  data_stage_5__2201_,data_stage_5__2200_,data_stage_5__2199_,data_stage_5__2198_,
  data_stage_5__2197_,data_stage_5__2196_,data_stage_5__2195_,data_stage_5__2194_,
  data_stage_5__2193_,data_stage_5__2192_,data_stage_5__2191_,data_stage_5__2190_,
  data_stage_5__2189_,data_stage_5__2188_,data_stage_5__2187_,data_stage_5__2186_,
  data_stage_5__2185_,data_stage_5__2184_,data_stage_5__2183_,data_stage_5__2182_,
  data_stage_5__2181_,data_stage_5__2180_,data_stage_5__2179_,data_stage_5__2178_,
  data_stage_5__2177_,data_stage_5__2176_,data_stage_5__2175_,data_stage_5__2174_,
  data_stage_5__2173_,data_stage_5__2172_,data_stage_5__2171_,data_stage_5__2170_,
  data_stage_5__2169_,data_stage_5__2168_,data_stage_5__2167_,data_stage_5__2166_,
  data_stage_5__2165_,data_stage_5__2164_,data_stage_5__2163_,data_stage_5__2162_,
  data_stage_5__2161_,data_stage_5__2160_,data_stage_5__2159_,data_stage_5__2158_,
  data_stage_5__2157_,data_stage_5__2156_,data_stage_5__2155_,data_stage_5__2154_,
  data_stage_5__2153_,data_stage_5__2152_,data_stage_5__2151_,data_stage_5__2150_,
  data_stage_5__2149_,data_stage_5__2148_,data_stage_5__2147_,data_stage_5__2146_,
  data_stage_5__2145_,data_stage_5__2144_,data_stage_5__2143_,data_stage_5__2142_,
  data_stage_5__2141_,data_stage_5__2140_,data_stage_5__2139_,data_stage_5__2138_,
  data_stage_5__2137_,data_stage_5__2136_,data_stage_5__2135_,data_stage_5__2134_,
  data_stage_5__2133_,data_stage_5__2132_,data_stage_5__2131_,data_stage_5__2130_,
  data_stage_5__2129_,data_stage_5__2128_,data_stage_5__2127_,data_stage_5__2126_,
  data_stage_5__2125_,data_stage_5__2124_,data_stage_5__2123_,data_stage_5__2122_,
  data_stage_5__2121_,data_stage_5__2120_,data_stage_5__2119_,data_stage_5__2118_,
  data_stage_5__2117_,data_stage_5__2116_,data_stage_5__2115_,data_stage_5__2114_,
  data_stage_5__2113_,data_stage_5__2112_,data_stage_5__2111_,data_stage_5__2110_,
  data_stage_5__2109_,data_stage_5__2108_,data_stage_5__2107_,data_stage_5__2106_,
  data_stage_5__2105_,data_stage_5__2104_,data_stage_5__2103_,data_stage_5__2102_,
  data_stage_5__2101_,data_stage_5__2100_,data_stage_5__2099_,data_stage_5__2098_,
  data_stage_5__2097_,data_stage_5__2096_,data_stage_5__2095_,data_stage_5__2094_,
  data_stage_5__2093_,data_stage_5__2092_,data_stage_5__2091_,data_stage_5__2090_,
  data_stage_5__2089_,data_stage_5__2088_,data_stage_5__2087_,data_stage_5__2086_,
  data_stage_5__2085_,data_stage_5__2084_,data_stage_5__2083_,data_stage_5__2082_,
  data_stage_5__2081_,data_stage_5__2080_,data_stage_5__2079_,data_stage_5__2078_,
  data_stage_5__2077_,data_stage_5__2076_,data_stage_5__2075_,data_stage_5__2074_,
  data_stage_5__2073_,data_stage_5__2072_,data_stage_5__2071_,data_stage_5__2070_,
  data_stage_5__2069_,data_stage_5__2068_,data_stage_5__2067_,data_stage_5__2066_,
  data_stage_5__2065_,data_stage_5__2064_,data_stage_5__2063_,data_stage_5__2062_,
  data_stage_5__2061_,data_stage_5__2060_,data_stage_5__2059_,data_stage_5__2058_,
  data_stage_5__2057_,data_stage_5__2056_,data_stage_5__2055_,data_stage_5__2054_,
  data_stage_5__2053_,data_stage_5__2052_,data_stage_5__2051_,data_stage_5__2050_,
  data_stage_5__2049_,data_stage_5__2048_,data_stage_5__2047_,data_stage_5__2046_,
  data_stage_5__2045_,data_stage_5__2044_,data_stage_5__2043_,data_stage_5__2042_,
  data_stage_5__2041_,data_stage_5__2040_,data_stage_5__2039_,data_stage_5__2038_,
  data_stage_5__2037_,data_stage_5__2036_,data_stage_5__2035_,data_stage_5__2034_,
  data_stage_5__2033_,data_stage_5__2032_,data_stage_5__2031_,data_stage_5__2030_,
  data_stage_5__2029_,data_stage_5__2028_,data_stage_5__2027_,data_stage_5__2026_,
  data_stage_5__2025_,data_stage_5__2024_,data_stage_5__2023_,data_stage_5__2022_,
  data_stage_5__2021_,data_stage_5__2020_,data_stage_5__2019_,data_stage_5__2018_,
  data_stage_5__2017_,data_stage_5__2016_,data_stage_5__2015_,data_stage_5__2014_,
  data_stage_5__2013_,data_stage_5__2012_,data_stage_5__2011_,data_stage_5__2010_,
  data_stage_5__2009_,data_stage_5__2008_,data_stage_5__2007_,data_stage_5__2006_,
  data_stage_5__2005_,data_stage_5__2004_,data_stage_5__2003_,data_stage_5__2002_,
  data_stage_5__2001_,data_stage_5__2000_,data_stage_5__1999_,data_stage_5__1998_,
  data_stage_5__1997_,data_stage_5__1996_,data_stage_5__1995_,data_stage_5__1994_,
  data_stage_5__1993_,data_stage_5__1992_,data_stage_5__1991_,data_stage_5__1990_,
  data_stage_5__1989_,data_stage_5__1988_,data_stage_5__1987_,data_stage_5__1986_,
  data_stage_5__1985_,data_stage_5__1984_,data_stage_5__1983_,data_stage_5__1982_,
  data_stage_5__1981_,data_stage_5__1980_,data_stage_5__1979_,data_stage_5__1978_,
  data_stage_5__1977_,data_stage_5__1976_,data_stage_5__1975_,data_stage_5__1974_,
  data_stage_5__1973_,data_stage_5__1972_,data_stage_5__1971_,data_stage_5__1970_,
  data_stage_5__1969_,data_stage_5__1968_,data_stage_5__1967_,data_stage_5__1966_,
  data_stage_5__1965_,data_stage_5__1964_,data_stage_5__1963_,data_stage_5__1962_,
  data_stage_5__1961_,data_stage_5__1960_,data_stage_5__1959_,data_stage_5__1958_,
  data_stage_5__1957_,data_stage_5__1956_,data_stage_5__1955_,data_stage_5__1954_,
  data_stage_5__1953_,data_stage_5__1952_,data_stage_5__1951_,data_stage_5__1950_,
  data_stage_5__1949_,data_stage_5__1948_,data_stage_5__1947_,data_stage_5__1946_,
  data_stage_5__1945_,data_stage_5__1944_,data_stage_5__1943_,data_stage_5__1942_,
  data_stage_5__1941_,data_stage_5__1940_,data_stage_5__1939_,data_stage_5__1938_,
  data_stage_5__1937_,data_stage_5__1936_,data_stage_5__1935_,data_stage_5__1934_,
  data_stage_5__1933_,data_stage_5__1932_,data_stage_5__1931_,data_stage_5__1930_,
  data_stage_5__1929_,data_stage_5__1928_,data_stage_5__1927_,data_stage_5__1926_,
  data_stage_5__1925_,data_stage_5__1924_,data_stage_5__1923_,data_stage_5__1922_,
  data_stage_5__1921_,data_stage_5__1920_,data_stage_5__1919_,data_stage_5__1918_,
  data_stage_5__1917_,data_stage_5__1916_,data_stage_5__1915_,data_stage_5__1914_,
  data_stage_5__1913_,data_stage_5__1912_,data_stage_5__1911_,data_stage_5__1910_,
  data_stage_5__1909_,data_stage_5__1908_,data_stage_5__1907_,data_stage_5__1906_,
  data_stage_5__1905_,data_stage_5__1904_,data_stage_5__1903_,data_stage_5__1902_,
  data_stage_5__1901_,data_stage_5__1900_,data_stage_5__1899_,data_stage_5__1898_,
  data_stage_5__1897_,data_stage_5__1896_,data_stage_5__1895_,data_stage_5__1894_,
  data_stage_5__1893_,data_stage_5__1892_,data_stage_5__1891_,data_stage_5__1890_,
  data_stage_5__1889_,data_stage_5__1888_,data_stage_5__1887_,data_stage_5__1886_,
  data_stage_5__1885_,data_stage_5__1884_,data_stage_5__1883_,data_stage_5__1882_,
  data_stage_5__1881_,data_stage_5__1880_,data_stage_5__1879_,data_stage_5__1878_,
  data_stage_5__1877_,data_stage_5__1876_,data_stage_5__1875_,data_stage_5__1874_,
  data_stage_5__1873_,data_stage_5__1872_,data_stage_5__1871_,data_stage_5__1870_,
  data_stage_5__1869_,data_stage_5__1868_,data_stage_5__1867_,data_stage_5__1866_,
  data_stage_5__1865_,data_stage_5__1864_,data_stage_5__1863_,data_stage_5__1862_,
  data_stage_5__1861_,data_stage_5__1860_,data_stage_5__1859_,data_stage_5__1858_,
  data_stage_5__1857_,data_stage_5__1856_,data_stage_5__1855_,data_stage_5__1854_,
  data_stage_5__1853_,data_stage_5__1852_,data_stage_5__1851_,data_stage_5__1850_,
  data_stage_5__1849_,data_stage_5__1848_,data_stage_5__1847_,data_stage_5__1846_,
  data_stage_5__1845_,data_stage_5__1844_,data_stage_5__1843_,data_stage_5__1842_,
  data_stage_5__1841_,data_stage_5__1840_,data_stage_5__1839_,data_stage_5__1838_,
  data_stage_5__1837_,data_stage_5__1836_,data_stage_5__1835_,data_stage_5__1834_,
  data_stage_5__1833_,data_stage_5__1832_,data_stage_5__1831_,data_stage_5__1830_,
  data_stage_5__1829_,data_stage_5__1828_,data_stage_5__1827_,data_stage_5__1826_,
  data_stage_5__1825_,data_stage_5__1824_,data_stage_5__1823_,data_stage_5__1822_,
  data_stage_5__1821_,data_stage_5__1820_,data_stage_5__1819_,data_stage_5__1818_,
  data_stage_5__1817_,data_stage_5__1816_,data_stage_5__1815_,data_stage_5__1814_,
  data_stage_5__1813_,data_stage_5__1812_,data_stage_5__1811_,data_stage_5__1810_,
  data_stage_5__1809_,data_stage_5__1808_,data_stage_5__1807_,data_stage_5__1806_,
  data_stage_5__1805_,data_stage_5__1804_,data_stage_5__1803_,data_stage_5__1802_,
  data_stage_5__1801_,data_stage_5__1800_,data_stage_5__1799_,data_stage_5__1798_,
  data_stage_5__1797_,data_stage_5__1796_,data_stage_5__1795_,data_stage_5__1794_,
  data_stage_5__1793_,data_stage_5__1792_,data_stage_5__1791_,data_stage_5__1790_,
  data_stage_5__1789_,data_stage_5__1788_,data_stage_5__1787_,data_stage_5__1786_,
  data_stage_5__1785_,data_stage_5__1784_,data_stage_5__1783_,data_stage_5__1782_,
  data_stage_5__1781_,data_stage_5__1780_,data_stage_5__1779_,data_stage_5__1778_,
  data_stage_5__1777_,data_stage_5__1776_,data_stage_5__1775_,data_stage_5__1774_,
  data_stage_5__1773_,data_stage_5__1772_,data_stage_5__1771_,data_stage_5__1770_,
  data_stage_5__1769_,data_stage_5__1768_,data_stage_5__1767_,data_stage_5__1766_,
  data_stage_5__1765_,data_stage_5__1764_,data_stage_5__1763_,data_stage_5__1762_,
  data_stage_5__1761_,data_stage_5__1760_,data_stage_5__1759_,data_stage_5__1758_,
  data_stage_5__1757_,data_stage_5__1756_,data_stage_5__1755_,data_stage_5__1754_,
  data_stage_5__1753_,data_stage_5__1752_,data_stage_5__1751_,data_stage_5__1750_,
  data_stage_5__1749_,data_stage_5__1748_,data_stage_5__1747_,data_stage_5__1746_,
  data_stage_5__1745_,data_stage_5__1744_,data_stage_5__1743_,data_stage_5__1742_,
  data_stage_5__1741_,data_stage_5__1740_,data_stage_5__1739_,data_stage_5__1738_,
  data_stage_5__1737_,data_stage_5__1736_,data_stage_5__1735_,data_stage_5__1734_,
  data_stage_5__1733_,data_stage_5__1732_,data_stage_5__1731_,data_stage_5__1730_,
  data_stage_5__1729_,data_stage_5__1728_,data_stage_5__1727_,data_stage_5__1726_,
  data_stage_5__1725_,data_stage_5__1724_,data_stage_5__1723_,data_stage_5__1722_,
  data_stage_5__1721_,data_stage_5__1720_,data_stage_5__1719_,data_stage_5__1718_,
  data_stage_5__1717_,data_stage_5__1716_,data_stage_5__1715_,data_stage_5__1714_,
  data_stage_5__1713_,data_stage_5__1712_,data_stage_5__1711_,data_stage_5__1710_,
  data_stage_5__1709_,data_stage_5__1708_,data_stage_5__1707_,data_stage_5__1706_,
  data_stage_5__1705_,data_stage_5__1704_,data_stage_5__1703_,data_stage_5__1702_,
  data_stage_5__1701_,data_stage_5__1700_,data_stage_5__1699_,data_stage_5__1698_,
  data_stage_5__1697_,data_stage_5__1696_,data_stage_5__1695_,data_stage_5__1694_,
  data_stage_5__1693_,data_stage_5__1692_,data_stage_5__1691_,data_stage_5__1690_,
  data_stage_5__1689_,data_stage_5__1688_,data_stage_5__1687_,data_stage_5__1686_,
  data_stage_5__1685_,data_stage_5__1684_,data_stage_5__1683_,data_stage_5__1682_,
  data_stage_5__1681_,data_stage_5__1680_,data_stage_5__1679_,data_stage_5__1678_,
  data_stage_5__1677_,data_stage_5__1676_,data_stage_5__1675_,data_stage_5__1674_,
  data_stage_5__1673_,data_stage_5__1672_,data_stage_5__1671_,data_stage_5__1670_,
  data_stage_5__1669_,data_stage_5__1668_,data_stage_5__1667_,data_stage_5__1666_,
  data_stage_5__1665_,data_stage_5__1664_,data_stage_5__1663_,data_stage_5__1662_,
  data_stage_5__1661_,data_stage_5__1660_,data_stage_5__1659_,data_stage_5__1658_,
  data_stage_5__1657_,data_stage_5__1656_,data_stage_5__1655_,data_stage_5__1654_,
  data_stage_5__1653_,data_stage_5__1652_,data_stage_5__1651_,data_stage_5__1650_,
  data_stage_5__1649_,data_stage_5__1648_,data_stage_5__1647_,data_stage_5__1646_,
  data_stage_5__1645_,data_stage_5__1644_,data_stage_5__1643_,data_stage_5__1642_,
  data_stage_5__1641_,data_stage_5__1640_,data_stage_5__1639_,data_stage_5__1638_,
  data_stage_5__1637_,data_stage_5__1636_,data_stage_5__1635_,data_stage_5__1634_,
  data_stage_5__1633_,data_stage_5__1632_,data_stage_5__1631_,data_stage_5__1630_,
  data_stage_5__1629_,data_stage_5__1628_,data_stage_5__1627_,data_stage_5__1626_,
  data_stage_5__1625_,data_stage_5__1624_,data_stage_5__1623_,data_stage_5__1622_,
  data_stage_5__1621_,data_stage_5__1620_,data_stage_5__1619_,data_stage_5__1618_,
  data_stage_5__1617_,data_stage_5__1616_,data_stage_5__1615_,data_stage_5__1614_,
  data_stage_5__1613_,data_stage_5__1612_,data_stage_5__1611_,data_stage_5__1610_,
  data_stage_5__1609_,data_stage_5__1608_,data_stage_5__1607_,data_stage_5__1606_,
  data_stage_5__1605_,data_stage_5__1604_,data_stage_5__1603_,data_stage_5__1602_,
  data_stage_5__1601_,data_stage_5__1600_,data_stage_5__1599_,data_stage_5__1598_,
  data_stage_5__1597_,data_stage_5__1596_,data_stage_5__1595_,data_stage_5__1594_,
  data_stage_5__1593_,data_stage_5__1592_,data_stage_5__1591_,data_stage_5__1590_,
  data_stage_5__1589_,data_stage_5__1588_,data_stage_5__1587_,data_stage_5__1586_,
  data_stage_5__1585_,data_stage_5__1584_,data_stage_5__1583_,data_stage_5__1582_,
  data_stage_5__1581_,data_stage_5__1580_,data_stage_5__1579_,data_stage_5__1578_,
  data_stage_5__1577_,data_stage_5__1576_,data_stage_5__1575_,data_stage_5__1574_,
  data_stage_5__1573_,data_stage_5__1572_,data_stage_5__1571_,data_stage_5__1570_,
  data_stage_5__1569_,data_stage_5__1568_,data_stage_5__1567_,data_stage_5__1566_,
  data_stage_5__1565_,data_stage_5__1564_,data_stage_5__1563_,data_stage_5__1562_,
  data_stage_5__1561_,data_stage_5__1560_,data_stage_5__1559_,data_stage_5__1558_,
  data_stage_5__1557_,data_stage_5__1556_,data_stage_5__1555_,data_stage_5__1554_,
  data_stage_5__1553_,data_stage_5__1552_,data_stage_5__1551_,data_stage_5__1550_,
  data_stage_5__1549_,data_stage_5__1548_,data_stage_5__1547_,data_stage_5__1546_,
  data_stage_5__1545_,data_stage_5__1544_,data_stage_5__1543_,data_stage_5__1542_,
  data_stage_5__1541_,data_stage_5__1540_,data_stage_5__1539_,data_stage_5__1538_,
  data_stage_5__1537_,data_stage_5__1536_,data_stage_5__1535_,data_stage_5__1534_,
  data_stage_5__1533_,data_stage_5__1532_,data_stage_5__1531_,data_stage_5__1530_,
  data_stage_5__1529_,data_stage_5__1528_,data_stage_5__1527_,data_stage_5__1526_,
  data_stage_5__1525_,data_stage_5__1524_,data_stage_5__1523_,data_stage_5__1522_,
  data_stage_5__1521_,data_stage_5__1520_,data_stage_5__1519_,data_stage_5__1518_,
  data_stage_5__1517_,data_stage_5__1516_,data_stage_5__1515_,data_stage_5__1514_,
  data_stage_5__1513_,data_stage_5__1512_,data_stage_5__1511_,data_stage_5__1510_,
  data_stage_5__1509_,data_stage_5__1508_,data_stage_5__1507_,data_stage_5__1506_,
  data_stage_5__1505_,data_stage_5__1504_,data_stage_5__1503_,data_stage_5__1502_,
  data_stage_5__1501_,data_stage_5__1500_,data_stage_5__1499_,data_stage_5__1498_,
  data_stage_5__1497_,data_stage_5__1496_,data_stage_5__1495_,data_stage_5__1494_,
  data_stage_5__1493_,data_stage_5__1492_,data_stage_5__1491_,data_stage_5__1490_,
  data_stage_5__1489_,data_stage_5__1488_,data_stage_5__1487_,data_stage_5__1486_,
  data_stage_5__1485_,data_stage_5__1484_,data_stage_5__1483_,data_stage_5__1482_,
  data_stage_5__1481_,data_stage_5__1480_,data_stage_5__1479_,data_stage_5__1478_,
  data_stage_5__1477_,data_stage_5__1476_,data_stage_5__1475_,data_stage_5__1474_,
  data_stage_5__1473_,data_stage_5__1472_,data_stage_5__1471_,data_stage_5__1470_,
  data_stage_5__1469_,data_stage_5__1468_,data_stage_5__1467_,data_stage_5__1466_,
  data_stage_5__1465_,data_stage_5__1464_,data_stage_5__1463_,data_stage_5__1462_,
  data_stage_5__1461_,data_stage_5__1460_,data_stage_5__1459_,data_stage_5__1458_,
  data_stage_5__1457_,data_stage_5__1456_,data_stage_5__1455_,data_stage_5__1454_,
  data_stage_5__1453_,data_stage_5__1452_,data_stage_5__1451_,data_stage_5__1450_,
  data_stage_5__1449_,data_stage_5__1448_,data_stage_5__1447_,data_stage_5__1446_,
  data_stage_5__1445_,data_stage_5__1444_,data_stage_5__1443_,data_stage_5__1442_,
  data_stage_5__1441_,data_stage_5__1440_,data_stage_5__1439_,data_stage_5__1438_,
  data_stage_5__1437_,data_stage_5__1436_,data_stage_5__1435_,data_stage_5__1434_,
  data_stage_5__1433_,data_stage_5__1432_,data_stage_5__1431_,data_stage_5__1430_,
  data_stage_5__1429_,data_stage_5__1428_,data_stage_5__1427_,data_stage_5__1426_,
  data_stage_5__1425_,data_stage_5__1424_,data_stage_5__1423_,data_stage_5__1422_,
  data_stage_5__1421_,data_stage_5__1420_,data_stage_5__1419_,data_stage_5__1418_,
  data_stage_5__1417_,data_stage_5__1416_,data_stage_5__1415_,data_stage_5__1414_,
  data_stage_5__1413_,data_stage_5__1412_,data_stage_5__1411_,data_stage_5__1410_,
  data_stage_5__1409_,data_stage_5__1408_,data_stage_5__1407_,data_stage_5__1406_,
  data_stage_5__1405_,data_stage_5__1404_,data_stage_5__1403_,data_stage_5__1402_,
  data_stage_5__1401_,data_stage_5__1400_,data_stage_5__1399_,data_stage_5__1398_,
  data_stage_5__1397_,data_stage_5__1396_,data_stage_5__1395_,data_stage_5__1394_,
  data_stage_5__1393_,data_stage_5__1392_,data_stage_5__1391_,data_stage_5__1390_,
  data_stage_5__1389_,data_stage_5__1388_,data_stage_5__1387_,data_stage_5__1386_,
  data_stage_5__1385_,data_stage_5__1384_,data_stage_5__1383_,data_stage_5__1382_,
  data_stage_5__1381_,data_stage_5__1380_,data_stage_5__1379_,data_stage_5__1378_,
  data_stage_5__1377_,data_stage_5__1376_,data_stage_5__1375_,data_stage_5__1374_,
  data_stage_5__1373_,data_stage_5__1372_,data_stage_5__1371_,data_stage_5__1370_,
  data_stage_5__1369_,data_stage_5__1368_,data_stage_5__1367_,data_stage_5__1366_,
  data_stage_5__1365_,data_stage_5__1364_,data_stage_5__1363_,data_stage_5__1362_,
  data_stage_5__1361_,data_stage_5__1360_,data_stage_5__1359_,data_stage_5__1358_,
  data_stage_5__1357_,data_stage_5__1356_,data_stage_5__1355_,data_stage_5__1354_,
  data_stage_5__1353_,data_stage_5__1352_,data_stage_5__1351_,data_stage_5__1350_,
  data_stage_5__1349_,data_stage_5__1348_,data_stage_5__1347_,data_stage_5__1346_,
  data_stage_5__1345_,data_stage_5__1344_,data_stage_5__1343_,data_stage_5__1342_,
  data_stage_5__1341_,data_stage_5__1340_,data_stage_5__1339_,data_stage_5__1338_,
  data_stage_5__1337_,data_stage_5__1336_,data_stage_5__1335_,data_stage_5__1334_,
  data_stage_5__1333_,data_stage_5__1332_,data_stage_5__1331_,data_stage_5__1330_,
  data_stage_5__1329_,data_stage_5__1328_,data_stage_5__1327_,data_stage_5__1326_,
  data_stage_5__1325_,data_stage_5__1324_,data_stage_5__1323_,data_stage_5__1322_,
  data_stage_5__1321_,data_stage_5__1320_,data_stage_5__1319_,data_stage_5__1318_,
  data_stage_5__1317_,data_stage_5__1316_,data_stage_5__1315_,data_stage_5__1314_,
  data_stage_5__1313_,data_stage_5__1312_,data_stage_5__1311_,data_stage_5__1310_,
  data_stage_5__1309_,data_stage_5__1308_,data_stage_5__1307_,data_stage_5__1306_,
  data_stage_5__1305_,data_stage_5__1304_,data_stage_5__1303_,data_stage_5__1302_,
  data_stage_5__1301_,data_stage_5__1300_,data_stage_5__1299_,data_stage_5__1298_,
  data_stage_5__1297_,data_stage_5__1296_,data_stage_5__1295_,data_stage_5__1294_,
  data_stage_5__1293_,data_stage_5__1292_,data_stage_5__1291_,data_stage_5__1290_,
  data_stage_5__1289_,data_stage_5__1288_,data_stage_5__1287_,data_stage_5__1286_,
  data_stage_5__1285_,data_stage_5__1284_,data_stage_5__1283_,data_stage_5__1282_,
  data_stage_5__1281_,data_stage_5__1280_,data_stage_5__1279_,data_stage_5__1278_,
  data_stage_5__1277_,data_stage_5__1276_,data_stage_5__1275_,data_stage_5__1274_,
  data_stage_5__1273_,data_stage_5__1272_,data_stage_5__1271_,data_stage_5__1270_,
  data_stage_5__1269_,data_stage_5__1268_,data_stage_5__1267_,data_stage_5__1266_,
  data_stage_5__1265_,data_stage_5__1264_,data_stage_5__1263_,data_stage_5__1262_,
  data_stage_5__1261_,data_stage_5__1260_,data_stage_5__1259_,data_stage_5__1258_,
  data_stage_5__1257_,data_stage_5__1256_,data_stage_5__1255_,data_stage_5__1254_,
  data_stage_5__1253_,data_stage_5__1252_,data_stage_5__1251_,data_stage_5__1250_,
  data_stage_5__1249_,data_stage_5__1248_,data_stage_5__1247_,data_stage_5__1246_,
  data_stage_5__1245_,data_stage_5__1244_,data_stage_5__1243_,data_stage_5__1242_,
  data_stage_5__1241_,data_stage_5__1240_,data_stage_5__1239_,data_stage_5__1238_,
  data_stage_5__1237_,data_stage_5__1236_,data_stage_5__1235_,data_stage_5__1234_,
  data_stage_5__1233_,data_stage_5__1232_,data_stage_5__1231_,data_stage_5__1230_,
  data_stage_5__1229_,data_stage_5__1228_,data_stage_5__1227_,data_stage_5__1226_,
  data_stage_5__1225_,data_stage_5__1224_,data_stage_5__1223_,data_stage_5__1222_,
  data_stage_5__1221_,data_stage_5__1220_,data_stage_5__1219_,data_stage_5__1218_,
  data_stage_5__1217_,data_stage_5__1216_,data_stage_5__1215_,data_stage_5__1214_,
  data_stage_5__1213_,data_stage_5__1212_,data_stage_5__1211_,data_stage_5__1210_,
  data_stage_5__1209_,data_stage_5__1208_,data_stage_5__1207_,data_stage_5__1206_,
  data_stage_5__1205_,data_stage_5__1204_,data_stage_5__1203_,data_stage_5__1202_,
  data_stage_5__1201_,data_stage_5__1200_,data_stage_5__1199_,data_stage_5__1198_,
  data_stage_5__1197_,data_stage_5__1196_,data_stage_5__1195_,data_stage_5__1194_,
  data_stage_5__1193_,data_stage_5__1192_,data_stage_5__1191_,data_stage_5__1190_,
  data_stage_5__1189_,data_stage_5__1188_,data_stage_5__1187_,data_stage_5__1186_,
  data_stage_5__1185_,data_stage_5__1184_,data_stage_5__1183_,data_stage_5__1182_,
  data_stage_5__1181_,data_stage_5__1180_,data_stage_5__1179_,data_stage_5__1178_,
  data_stage_5__1177_,data_stage_5__1176_,data_stage_5__1175_,data_stage_5__1174_,
  data_stage_5__1173_,data_stage_5__1172_,data_stage_5__1171_,data_stage_5__1170_,
  data_stage_5__1169_,data_stage_5__1168_,data_stage_5__1167_,data_stage_5__1166_,
  data_stage_5__1165_,data_stage_5__1164_,data_stage_5__1163_,data_stage_5__1162_,
  data_stage_5__1161_,data_stage_5__1160_,data_stage_5__1159_,data_stage_5__1158_,
  data_stage_5__1157_,data_stage_5__1156_,data_stage_5__1155_,data_stage_5__1154_,
  data_stage_5__1153_,data_stage_5__1152_,data_stage_5__1151_,data_stage_5__1150_,
  data_stage_5__1149_,data_stage_5__1148_,data_stage_5__1147_,data_stage_5__1146_,
  data_stage_5__1145_,data_stage_5__1144_,data_stage_5__1143_,data_stage_5__1142_,
  data_stage_5__1141_,data_stage_5__1140_,data_stage_5__1139_,data_stage_5__1138_,
  data_stage_5__1137_,data_stage_5__1136_,data_stage_5__1135_,data_stage_5__1134_,
  data_stage_5__1133_,data_stage_5__1132_,data_stage_5__1131_,data_stage_5__1130_,
  data_stage_5__1129_,data_stage_5__1128_,data_stage_5__1127_,data_stage_5__1126_,
  data_stage_5__1125_,data_stage_5__1124_,data_stage_5__1123_,data_stage_5__1122_,
  data_stage_5__1121_,data_stage_5__1120_,data_stage_5__1119_,data_stage_5__1118_,
  data_stage_5__1117_,data_stage_5__1116_,data_stage_5__1115_,data_stage_5__1114_,
  data_stage_5__1113_,data_stage_5__1112_,data_stage_5__1111_,data_stage_5__1110_,
  data_stage_5__1109_,data_stage_5__1108_,data_stage_5__1107_,data_stage_5__1106_,
  data_stage_5__1105_,data_stage_5__1104_,data_stage_5__1103_,data_stage_5__1102_,
  data_stage_5__1101_,data_stage_5__1100_,data_stage_5__1099_,data_stage_5__1098_,
  data_stage_5__1097_,data_stage_5__1096_,data_stage_5__1095_,data_stage_5__1094_,
  data_stage_5__1093_,data_stage_5__1092_,data_stage_5__1091_,data_stage_5__1090_,
  data_stage_5__1089_,data_stage_5__1088_,data_stage_5__1087_,data_stage_5__1086_,
  data_stage_5__1085_,data_stage_5__1084_,data_stage_5__1083_,data_stage_5__1082_,
  data_stage_5__1081_,data_stage_5__1080_,data_stage_5__1079_,data_stage_5__1078_,
  data_stage_5__1077_,data_stage_5__1076_,data_stage_5__1075_,data_stage_5__1074_,
  data_stage_5__1073_,data_stage_5__1072_,data_stage_5__1071_,data_stage_5__1070_,
  data_stage_5__1069_,data_stage_5__1068_,data_stage_5__1067_,data_stage_5__1066_,
  data_stage_5__1065_,data_stage_5__1064_,data_stage_5__1063_,data_stage_5__1062_,
  data_stage_5__1061_,data_stage_5__1060_,data_stage_5__1059_,data_stage_5__1058_,
  data_stage_5__1057_,data_stage_5__1056_,data_stage_5__1055_,data_stage_5__1054_,
  data_stage_5__1053_,data_stage_5__1052_,data_stage_5__1051_,data_stage_5__1050_,
  data_stage_5__1049_,data_stage_5__1048_,data_stage_5__1047_,data_stage_5__1046_,
  data_stage_5__1045_,data_stage_5__1044_,data_stage_5__1043_,data_stage_5__1042_,
  data_stage_5__1041_,data_stage_5__1040_,data_stage_5__1039_,data_stage_5__1038_,
  data_stage_5__1037_,data_stage_5__1036_,data_stage_5__1035_,data_stage_5__1034_,
  data_stage_5__1033_,data_stage_5__1032_,data_stage_5__1031_,data_stage_5__1030_,
  data_stage_5__1029_,data_stage_5__1028_,data_stage_5__1027_,data_stage_5__1026_,
  data_stage_5__1025_,data_stage_5__1024_,data_stage_5__1023_,data_stage_5__1022_,
  data_stage_5__1021_,data_stage_5__1020_,data_stage_5__1019_,data_stage_5__1018_,
  data_stage_5__1017_,data_stage_5__1016_,data_stage_5__1015_,data_stage_5__1014_,
  data_stage_5__1013_,data_stage_5__1012_,data_stage_5__1011_,data_stage_5__1010_,
  data_stage_5__1009_,data_stage_5__1008_,data_stage_5__1007_,data_stage_5__1006_,
  data_stage_5__1005_,data_stage_5__1004_,data_stage_5__1003_,data_stage_5__1002_,
  data_stage_5__1001_,data_stage_5__1000_,data_stage_5__999_,data_stage_5__998_,
  data_stage_5__997_,data_stage_5__996_,data_stage_5__995_,data_stage_5__994_,
  data_stage_5__993_,data_stage_5__992_,data_stage_5__991_,data_stage_5__990_,
  data_stage_5__989_,data_stage_5__988_,data_stage_5__987_,data_stage_5__986_,
  data_stage_5__985_,data_stage_5__984_,data_stage_5__983_,data_stage_5__982_,
  data_stage_5__981_,data_stage_5__980_,data_stage_5__979_,data_stage_5__978_,data_stage_5__977_,
  data_stage_5__976_,data_stage_5__975_,data_stage_5__974_,data_stage_5__973_,
  data_stage_5__972_,data_stage_5__971_,data_stage_5__970_,data_stage_5__969_,
  data_stage_5__968_,data_stage_5__967_,data_stage_5__966_,data_stage_5__965_,
  data_stage_5__964_,data_stage_5__963_,data_stage_5__962_,data_stage_5__961_,data_stage_5__960_,
  data_stage_5__959_,data_stage_5__958_,data_stage_5__957_,data_stage_5__956_,
  data_stage_5__955_,data_stage_5__954_,data_stage_5__953_,data_stage_5__952_,
  data_stage_5__951_,data_stage_5__950_,data_stage_5__949_,data_stage_5__948_,
  data_stage_5__947_,data_stage_5__946_,data_stage_5__945_,data_stage_5__944_,
  data_stage_5__943_,data_stage_5__942_,data_stage_5__941_,data_stage_5__940_,data_stage_5__939_,
  data_stage_5__938_,data_stage_5__937_,data_stage_5__936_,data_stage_5__935_,
  data_stage_5__934_,data_stage_5__933_,data_stage_5__932_,data_stage_5__931_,
  data_stage_5__930_,data_stage_5__929_,data_stage_5__928_,data_stage_5__927_,
  data_stage_5__926_,data_stage_5__925_,data_stage_5__924_,data_stage_5__923_,
  data_stage_5__922_,data_stage_5__921_,data_stage_5__920_,data_stage_5__919_,data_stage_5__918_,
  data_stage_5__917_,data_stage_5__916_,data_stage_5__915_,data_stage_5__914_,
  data_stage_5__913_,data_stage_5__912_,data_stage_5__911_,data_stage_5__910_,
  data_stage_5__909_,data_stage_5__908_,data_stage_5__907_,data_stage_5__906_,
  data_stage_5__905_,data_stage_5__904_,data_stage_5__903_,data_stage_5__902_,
  data_stage_5__901_,data_stage_5__900_,data_stage_5__899_,data_stage_5__898_,data_stage_5__897_,
  data_stage_5__896_,data_stage_5__895_,data_stage_5__894_,data_stage_5__893_,
  data_stage_5__892_,data_stage_5__891_,data_stage_5__890_,data_stage_5__889_,
  data_stage_5__888_,data_stage_5__887_,data_stage_5__886_,data_stage_5__885_,
  data_stage_5__884_,data_stage_5__883_,data_stage_5__882_,data_stage_5__881_,data_stage_5__880_,
  data_stage_5__879_,data_stage_5__878_,data_stage_5__877_,data_stage_5__876_,
  data_stage_5__875_,data_stage_5__874_,data_stage_5__873_,data_stage_5__872_,
  data_stage_5__871_,data_stage_5__870_,data_stage_5__869_,data_stage_5__868_,
  data_stage_5__867_,data_stage_5__866_,data_stage_5__865_,data_stage_5__864_,
  data_stage_5__863_,data_stage_5__862_,data_stage_5__861_,data_stage_5__860_,data_stage_5__859_,
  data_stage_5__858_,data_stage_5__857_,data_stage_5__856_,data_stage_5__855_,
  data_stage_5__854_,data_stage_5__853_,data_stage_5__852_,data_stage_5__851_,
  data_stage_5__850_,data_stage_5__849_,data_stage_5__848_,data_stage_5__847_,
  data_stage_5__846_,data_stage_5__845_,data_stage_5__844_,data_stage_5__843_,
  data_stage_5__842_,data_stage_5__841_,data_stage_5__840_,data_stage_5__839_,data_stage_5__838_,
  data_stage_5__837_,data_stage_5__836_,data_stage_5__835_,data_stage_5__834_,
  data_stage_5__833_,data_stage_5__832_,data_stage_5__831_,data_stage_5__830_,
  data_stage_5__829_,data_stage_5__828_,data_stage_5__827_,data_stage_5__826_,
  data_stage_5__825_,data_stage_5__824_,data_stage_5__823_,data_stage_5__822_,
  data_stage_5__821_,data_stage_5__820_,data_stage_5__819_,data_stage_5__818_,data_stage_5__817_,
  data_stage_5__816_,data_stage_5__815_,data_stage_5__814_,data_stage_5__813_,
  data_stage_5__812_,data_stage_5__811_,data_stage_5__810_,data_stage_5__809_,
  data_stage_5__808_,data_stage_5__807_,data_stage_5__806_,data_stage_5__805_,
  data_stage_5__804_,data_stage_5__803_,data_stage_5__802_,data_stage_5__801_,data_stage_5__800_,
  data_stage_5__799_,data_stage_5__798_,data_stage_5__797_,data_stage_5__796_,
  data_stage_5__795_,data_stage_5__794_,data_stage_5__793_,data_stage_5__792_,
  data_stage_5__791_,data_stage_5__790_,data_stage_5__789_,data_stage_5__788_,
  data_stage_5__787_,data_stage_5__786_,data_stage_5__785_,data_stage_5__784_,
  data_stage_5__783_,data_stage_5__782_,data_stage_5__781_,data_stage_5__780_,data_stage_5__779_,
  data_stage_5__778_,data_stage_5__777_,data_stage_5__776_,data_stage_5__775_,
  data_stage_5__774_,data_stage_5__773_,data_stage_5__772_,data_stage_5__771_,
  data_stage_5__770_,data_stage_5__769_,data_stage_5__768_,data_stage_5__767_,
  data_stage_5__766_,data_stage_5__765_,data_stage_5__764_,data_stage_5__763_,
  data_stage_5__762_,data_stage_5__761_,data_stage_5__760_,data_stage_5__759_,data_stage_5__758_,
  data_stage_5__757_,data_stage_5__756_,data_stage_5__755_,data_stage_5__754_,
  data_stage_5__753_,data_stage_5__752_,data_stage_5__751_,data_stage_5__750_,
  data_stage_5__749_,data_stage_5__748_,data_stage_5__747_,data_stage_5__746_,
  data_stage_5__745_,data_stage_5__744_,data_stage_5__743_,data_stage_5__742_,
  data_stage_5__741_,data_stage_5__740_,data_stage_5__739_,data_stage_5__738_,data_stage_5__737_,
  data_stage_5__736_,data_stage_5__735_,data_stage_5__734_,data_stage_5__733_,
  data_stage_5__732_,data_stage_5__731_,data_stage_5__730_,data_stage_5__729_,
  data_stage_5__728_,data_stage_5__727_,data_stage_5__726_,data_stage_5__725_,
  data_stage_5__724_,data_stage_5__723_,data_stage_5__722_,data_stage_5__721_,data_stage_5__720_,
  data_stage_5__719_,data_stage_5__718_,data_stage_5__717_,data_stage_5__716_,
  data_stage_5__715_,data_stage_5__714_,data_stage_5__713_,data_stage_5__712_,
  data_stage_5__711_,data_stage_5__710_,data_stage_5__709_,data_stage_5__708_,
  data_stage_5__707_,data_stage_5__706_,data_stage_5__705_,data_stage_5__704_,
  data_stage_5__703_,data_stage_5__702_,data_stage_5__701_,data_stage_5__700_,data_stage_5__699_,
  data_stage_5__698_,data_stage_5__697_,data_stage_5__696_,data_stage_5__695_,
  data_stage_5__694_,data_stage_5__693_,data_stage_5__692_,data_stage_5__691_,
  data_stage_5__690_,data_stage_5__689_,data_stage_5__688_,data_stage_5__687_,
  data_stage_5__686_,data_stage_5__685_,data_stage_5__684_,data_stage_5__683_,
  data_stage_5__682_,data_stage_5__681_,data_stage_5__680_,data_stage_5__679_,data_stage_5__678_,
  data_stage_5__677_,data_stage_5__676_,data_stage_5__675_,data_stage_5__674_,
  data_stage_5__673_,data_stage_5__672_,data_stage_5__671_,data_stage_5__670_,
  data_stage_5__669_,data_stage_5__668_,data_stage_5__667_,data_stage_5__666_,
  data_stage_5__665_,data_stage_5__664_,data_stage_5__663_,data_stage_5__662_,
  data_stage_5__661_,data_stage_5__660_,data_stage_5__659_,data_stage_5__658_,data_stage_5__657_,
  data_stage_5__656_,data_stage_5__655_,data_stage_5__654_,data_stage_5__653_,
  data_stage_5__652_,data_stage_5__651_,data_stage_5__650_,data_stage_5__649_,
  data_stage_5__648_,data_stage_5__647_,data_stage_5__646_,data_stage_5__645_,
  data_stage_5__644_,data_stage_5__643_,data_stage_5__642_,data_stage_5__641_,data_stage_5__640_,
  data_stage_5__639_,data_stage_5__638_,data_stage_5__637_,data_stage_5__636_,
  data_stage_5__635_,data_stage_5__634_,data_stage_5__633_,data_stage_5__632_,
  data_stage_5__631_,data_stage_5__630_,data_stage_5__629_,data_stage_5__628_,
  data_stage_5__627_,data_stage_5__626_,data_stage_5__625_,data_stage_5__624_,
  data_stage_5__623_,data_stage_5__622_,data_stage_5__621_,data_stage_5__620_,data_stage_5__619_,
  data_stage_5__618_,data_stage_5__617_,data_stage_5__616_,data_stage_5__615_,
  data_stage_5__614_,data_stage_5__613_,data_stage_5__612_,data_stage_5__611_,
  data_stage_5__610_,data_stage_5__609_,data_stage_5__608_,data_stage_5__607_,
  data_stage_5__606_,data_stage_5__605_,data_stage_5__604_,data_stage_5__603_,
  data_stage_5__602_,data_stage_5__601_,data_stage_5__600_,data_stage_5__599_,data_stage_5__598_,
  data_stage_5__597_,data_stage_5__596_,data_stage_5__595_,data_stage_5__594_,
  data_stage_5__593_,data_stage_5__592_,data_stage_5__591_,data_stage_5__590_,
  data_stage_5__589_,data_stage_5__588_,data_stage_5__587_,data_stage_5__586_,
  data_stage_5__585_,data_stage_5__584_,data_stage_5__583_,data_stage_5__582_,
  data_stage_5__581_,data_stage_5__580_,data_stage_5__579_,data_stage_5__578_,data_stage_5__577_,
  data_stage_5__576_,data_stage_5__575_,data_stage_5__574_,data_stage_5__573_,
  data_stage_5__572_,data_stage_5__571_,data_stage_5__570_,data_stage_5__569_,
  data_stage_5__568_,data_stage_5__567_,data_stage_5__566_,data_stage_5__565_,
  data_stage_5__564_,data_stage_5__563_,data_stage_5__562_,data_stage_5__561_,data_stage_5__560_,
  data_stage_5__559_,data_stage_5__558_,data_stage_5__557_,data_stage_5__556_,
  data_stage_5__555_,data_stage_5__554_,data_stage_5__553_,data_stage_5__552_,
  data_stage_5__551_,data_stage_5__550_,data_stage_5__549_,data_stage_5__548_,
  data_stage_5__547_,data_stage_5__546_,data_stage_5__545_,data_stage_5__544_,
  data_stage_5__543_,data_stage_5__542_,data_stage_5__541_,data_stage_5__540_,data_stage_5__539_,
  data_stage_5__538_,data_stage_5__537_,data_stage_5__536_,data_stage_5__535_,
  data_stage_5__534_,data_stage_5__533_,data_stage_5__532_,data_stage_5__531_,
  data_stage_5__530_,data_stage_5__529_,data_stage_5__528_,data_stage_5__527_,
  data_stage_5__526_,data_stage_5__525_,data_stage_5__524_,data_stage_5__523_,
  data_stage_5__522_,data_stage_5__521_,data_stage_5__520_,data_stage_5__519_,data_stage_5__518_,
  data_stage_5__517_,data_stage_5__516_,data_stage_5__515_,data_stage_5__514_,
  data_stage_5__513_,data_stage_5__512_,data_stage_5__511_,data_stage_5__510_,
  data_stage_5__509_,data_stage_5__508_,data_stage_5__507_,data_stage_5__506_,
  data_stage_5__505_,data_stage_5__504_,data_stage_5__503_,data_stage_5__502_,
  data_stage_5__501_,data_stage_5__500_,data_stage_5__499_,data_stage_5__498_,data_stage_5__497_,
  data_stage_5__496_,data_stage_5__495_,data_stage_5__494_,data_stage_5__493_,
  data_stage_5__492_,data_stage_5__491_,data_stage_5__490_,data_stage_5__489_,
  data_stage_5__488_,data_stage_5__487_,data_stage_5__486_,data_stage_5__485_,
  data_stage_5__484_,data_stage_5__483_,data_stage_5__482_,data_stage_5__481_,data_stage_5__480_,
  data_stage_5__479_,data_stage_5__478_,data_stage_5__477_,data_stage_5__476_,
  data_stage_5__475_,data_stage_5__474_,data_stage_5__473_,data_stage_5__472_,
  data_stage_5__471_,data_stage_5__470_,data_stage_5__469_,data_stage_5__468_,
  data_stage_5__467_,data_stage_5__466_,data_stage_5__465_,data_stage_5__464_,
  data_stage_5__463_,data_stage_5__462_,data_stage_5__461_,data_stage_5__460_,data_stage_5__459_,
  data_stage_5__458_,data_stage_5__457_,data_stage_5__456_,data_stage_5__455_,
  data_stage_5__454_,data_stage_5__453_,data_stage_5__452_,data_stage_5__451_,
  data_stage_5__450_,data_stage_5__449_,data_stage_5__448_,data_stage_5__447_,
  data_stage_5__446_,data_stage_5__445_,data_stage_5__444_,data_stage_5__443_,
  data_stage_5__442_,data_stage_5__441_,data_stage_5__440_,data_stage_5__439_,data_stage_5__438_,
  data_stage_5__437_,data_stage_5__436_,data_stage_5__435_,data_stage_5__434_,
  data_stage_5__433_,data_stage_5__432_,data_stage_5__431_,data_stage_5__430_,
  data_stage_5__429_,data_stage_5__428_,data_stage_5__427_,data_stage_5__426_,
  data_stage_5__425_,data_stage_5__424_,data_stage_5__423_,data_stage_5__422_,
  data_stage_5__421_,data_stage_5__420_,data_stage_5__419_,data_stage_5__418_,data_stage_5__417_,
  data_stage_5__416_,data_stage_5__415_,data_stage_5__414_,data_stage_5__413_,
  data_stage_5__412_,data_stage_5__411_,data_stage_5__410_,data_stage_5__409_,
  data_stage_5__408_,data_stage_5__407_,data_stage_5__406_,data_stage_5__405_,
  data_stage_5__404_,data_stage_5__403_,data_stage_5__402_,data_stage_5__401_,data_stage_5__400_,
  data_stage_5__399_,data_stage_5__398_,data_stage_5__397_,data_stage_5__396_,
  data_stage_5__395_,data_stage_5__394_,data_stage_5__393_,data_stage_5__392_,
  data_stage_5__391_,data_stage_5__390_,data_stage_5__389_,data_stage_5__388_,
  data_stage_5__387_,data_stage_5__386_,data_stage_5__385_,data_stage_5__384_,
  data_stage_5__383_,data_stage_5__382_,data_stage_5__381_,data_stage_5__380_,data_stage_5__379_,
  data_stage_5__378_,data_stage_5__377_,data_stage_5__376_,data_stage_5__375_,
  data_stage_5__374_,data_stage_5__373_,data_stage_5__372_,data_stage_5__371_,
  data_stage_5__370_,data_stage_5__369_,data_stage_5__368_,data_stage_5__367_,
  data_stage_5__366_,data_stage_5__365_,data_stage_5__364_,data_stage_5__363_,
  data_stage_5__362_,data_stage_5__361_,data_stage_5__360_,data_stage_5__359_,data_stage_5__358_,
  data_stage_5__357_,data_stage_5__356_,data_stage_5__355_,data_stage_5__354_,
  data_stage_5__353_,data_stage_5__352_,data_stage_5__351_,data_stage_5__350_,
  data_stage_5__349_,data_stage_5__348_,data_stage_5__347_,data_stage_5__346_,
  data_stage_5__345_,data_stage_5__344_,data_stage_5__343_,data_stage_5__342_,
  data_stage_5__341_,data_stage_5__340_,data_stage_5__339_,data_stage_5__338_,data_stage_5__337_,
  data_stage_5__336_,data_stage_5__335_,data_stage_5__334_,data_stage_5__333_,
  data_stage_5__332_,data_stage_5__331_,data_stage_5__330_,data_stage_5__329_,
  data_stage_5__328_,data_stage_5__327_,data_stage_5__326_,data_stage_5__325_,
  data_stage_5__324_,data_stage_5__323_,data_stage_5__322_,data_stage_5__321_,data_stage_5__320_,
  data_stage_5__319_,data_stage_5__318_,data_stage_5__317_,data_stage_5__316_,
  data_stage_5__315_,data_stage_5__314_,data_stage_5__313_,data_stage_5__312_,
  data_stage_5__311_,data_stage_5__310_,data_stage_5__309_,data_stage_5__308_,
  data_stage_5__307_,data_stage_5__306_,data_stage_5__305_,data_stage_5__304_,
  data_stage_5__303_,data_stage_5__302_,data_stage_5__301_,data_stage_5__300_,data_stage_5__299_,
  data_stage_5__298_,data_stage_5__297_,data_stage_5__296_,data_stage_5__295_,
  data_stage_5__294_,data_stage_5__293_,data_stage_5__292_,data_stage_5__291_,
  data_stage_5__290_,data_stage_5__289_,data_stage_5__288_,data_stage_5__287_,
  data_stage_5__286_,data_stage_5__285_,data_stage_5__284_,data_stage_5__283_,
  data_stage_5__282_,data_stage_5__281_,data_stage_5__280_,data_stage_5__279_,data_stage_5__278_,
  data_stage_5__277_,data_stage_5__276_,data_stage_5__275_,data_stage_5__274_,
  data_stage_5__273_,data_stage_5__272_,data_stage_5__271_,data_stage_5__270_,
  data_stage_5__269_,data_stage_5__268_,data_stage_5__267_,data_stage_5__266_,
  data_stage_5__265_,data_stage_5__264_,data_stage_5__263_,data_stage_5__262_,
  data_stage_5__261_,data_stage_5__260_,data_stage_5__259_,data_stage_5__258_,data_stage_5__257_,
  data_stage_5__256_,data_stage_5__255_,data_stage_5__254_,data_stage_5__253_,
  data_stage_5__252_,data_stage_5__251_,data_stage_5__250_,data_stage_5__249_,
  data_stage_5__248_,data_stage_5__247_,data_stage_5__246_,data_stage_5__245_,
  data_stage_5__244_,data_stage_5__243_,data_stage_5__242_,data_stage_5__241_,data_stage_5__240_,
  data_stage_5__239_,data_stage_5__238_,data_stage_5__237_,data_stage_5__236_,
  data_stage_5__235_,data_stage_5__234_,data_stage_5__233_,data_stage_5__232_,
  data_stage_5__231_,data_stage_5__230_,data_stage_5__229_,data_stage_5__228_,
  data_stage_5__227_,data_stage_5__226_,data_stage_5__225_,data_stage_5__224_,
  data_stage_5__223_,data_stage_5__222_,data_stage_5__221_,data_stage_5__220_,data_stage_5__219_,
  data_stage_5__218_,data_stage_5__217_,data_stage_5__216_,data_stage_5__215_,
  data_stage_5__214_,data_stage_5__213_,data_stage_5__212_,data_stage_5__211_,
  data_stage_5__210_,data_stage_5__209_,data_stage_5__208_,data_stage_5__207_,
  data_stage_5__206_,data_stage_5__205_,data_stage_5__204_,data_stage_5__203_,
  data_stage_5__202_,data_stage_5__201_,data_stage_5__200_,data_stage_5__199_,data_stage_5__198_,
  data_stage_5__197_,data_stage_5__196_,data_stage_5__195_,data_stage_5__194_,
  data_stage_5__193_,data_stage_5__192_,data_stage_5__191_,data_stage_5__190_,
  data_stage_5__189_,data_stage_5__188_,data_stage_5__187_,data_stage_5__186_,
  data_stage_5__185_,data_stage_5__184_,data_stage_5__183_,data_stage_5__182_,
  data_stage_5__181_,data_stage_5__180_,data_stage_5__179_,data_stage_5__178_,data_stage_5__177_,
  data_stage_5__176_,data_stage_5__175_,data_stage_5__174_,data_stage_5__173_,
  data_stage_5__172_,data_stage_5__171_,data_stage_5__170_,data_stage_5__169_,
  data_stage_5__168_,data_stage_5__167_,data_stage_5__166_,data_stage_5__165_,
  data_stage_5__164_,data_stage_5__163_,data_stage_5__162_,data_stage_5__161_,data_stage_5__160_,
  data_stage_5__159_,data_stage_5__158_,data_stage_5__157_,data_stage_5__156_,
  data_stage_5__155_,data_stage_5__154_,data_stage_5__153_,data_stage_5__152_,
  data_stage_5__151_,data_stage_5__150_,data_stage_5__149_,data_stage_5__148_,
  data_stage_5__147_,data_stage_5__146_,data_stage_5__145_,data_stage_5__144_,
  data_stage_5__143_,data_stage_5__142_,data_stage_5__141_,data_stage_5__140_,data_stage_5__139_,
  data_stage_5__138_,data_stage_5__137_,data_stage_5__136_,data_stage_5__135_,
  data_stage_5__134_,data_stage_5__133_,data_stage_5__132_,data_stage_5__131_,
  data_stage_5__130_,data_stage_5__129_,data_stage_5__128_,data_stage_5__127_,
  data_stage_5__126_,data_stage_5__125_,data_stage_5__124_,data_stage_5__123_,
  data_stage_5__122_,data_stage_5__121_,data_stage_5__120_,data_stage_5__119_,data_stage_5__118_,
  data_stage_5__117_,data_stage_5__116_,data_stage_5__115_,data_stage_5__114_,
  data_stage_5__113_,data_stage_5__112_,data_stage_5__111_,data_stage_5__110_,
  data_stage_5__109_,data_stage_5__108_,data_stage_5__107_,data_stage_5__106_,
  data_stage_5__105_,data_stage_5__104_,data_stage_5__103_,data_stage_5__102_,
  data_stage_5__101_,data_stage_5__100_,data_stage_5__99_,data_stage_5__98_,data_stage_5__97_,
  data_stage_5__96_,data_stage_5__95_,data_stage_5__94_,data_stage_5__93_,
  data_stage_5__92_,data_stage_5__91_,data_stage_5__90_,data_stage_5__89_,data_stage_5__88_,
  data_stage_5__87_,data_stage_5__86_,data_stage_5__85_,data_stage_5__84_,
  data_stage_5__83_,data_stage_5__82_,data_stage_5__81_,data_stage_5__80_,data_stage_5__79_,
  data_stage_5__78_,data_stage_5__77_,data_stage_5__76_,data_stage_5__75_,
  data_stage_5__74_,data_stage_5__73_,data_stage_5__72_,data_stage_5__71_,data_stage_5__70_,
  data_stage_5__69_,data_stage_5__68_,data_stage_5__67_,data_stage_5__66_,
  data_stage_5__65_,data_stage_5__64_,data_stage_5__63_,data_stage_5__62_,
  data_stage_5__61_,data_stage_5__60_,data_stage_5__59_,data_stage_5__58_,data_stage_5__57_,
  data_stage_5__56_,data_stage_5__55_,data_stage_5__54_,data_stage_5__53_,
  data_stage_5__52_,data_stage_5__51_,data_stage_5__50_,data_stage_5__49_,data_stage_5__48_,
  data_stage_5__47_,data_stage_5__46_,data_stage_5__45_,data_stage_5__44_,
  data_stage_5__43_,data_stage_5__42_,data_stage_5__41_,data_stage_5__40_,data_stage_5__39_,
  data_stage_5__38_,data_stage_5__37_,data_stage_5__36_,data_stage_5__35_,
  data_stage_5__34_,data_stage_5__33_,data_stage_5__32_,data_stage_5__31_,data_stage_5__30_,
  data_stage_5__29_,data_stage_5__28_,data_stage_5__27_,data_stage_5__26_,
  data_stage_5__25_,data_stage_5__24_,data_stage_5__23_,data_stage_5__22_,
  data_stage_5__21_,data_stage_5__20_,data_stage_5__19_,data_stage_5__18_,data_stage_5__17_,
  data_stage_5__16_,data_stage_5__15_,data_stage_5__14_,data_stage_5__13_,
  data_stage_5__12_,data_stage_5__11_,data_stage_5__10_,data_stage_5__9_,data_stage_5__8_,
  data_stage_5__7_,data_stage_5__6_,data_stage_5__5_,data_stage_5__4_,data_stage_5__3_,
  data_stage_5__2_,data_stage_5__1_,data_stage_5__0_;

  bsg_swap_width_p128
  mux_stage_0__mux_swap_0__swap_inst
  (
    .data_i(data_i[255:0]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_, data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_, data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_, data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_1__swap_inst
  (
    .data_i(data_i[511:256]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_, data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_, data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_, data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_2__swap_inst
  (
    .data_i(data_i[767:512]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__767_, data_stage_1__766_, data_stage_1__765_, data_stage_1__764_, data_stage_1__763_, data_stage_1__762_, data_stage_1__761_, data_stage_1__760_, data_stage_1__759_, data_stage_1__758_, data_stage_1__757_, data_stage_1__756_, data_stage_1__755_, data_stage_1__754_, data_stage_1__753_, data_stage_1__752_, data_stage_1__751_, data_stage_1__750_, data_stage_1__749_, data_stage_1__748_, data_stage_1__747_, data_stage_1__746_, data_stage_1__745_, data_stage_1__744_, data_stage_1__743_, data_stage_1__742_, data_stage_1__741_, data_stage_1__740_, data_stage_1__739_, data_stage_1__738_, data_stage_1__737_, data_stage_1__736_, data_stage_1__735_, data_stage_1__734_, data_stage_1__733_, data_stage_1__732_, data_stage_1__731_, data_stage_1__730_, data_stage_1__729_, data_stage_1__728_, data_stage_1__727_, data_stage_1__726_, data_stage_1__725_, data_stage_1__724_, data_stage_1__723_, data_stage_1__722_, data_stage_1__721_, data_stage_1__720_, data_stage_1__719_, data_stage_1__718_, data_stage_1__717_, data_stage_1__716_, data_stage_1__715_, data_stage_1__714_, data_stage_1__713_, data_stage_1__712_, data_stage_1__711_, data_stage_1__710_, data_stage_1__709_, data_stage_1__708_, data_stage_1__707_, data_stage_1__706_, data_stage_1__705_, data_stage_1__704_, data_stage_1__703_, data_stage_1__702_, data_stage_1__701_, data_stage_1__700_, data_stage_1__699_, data_stage_1__698_, data_stage_1__697_, data_stage_1__696_, data_stage_1__695_, data_stage_1__694_, data_stage_1__693_, data_stage_1__692_, data_stage_1__691_, data_stage_1__690_, data_stage_1__689_, data_stage_1__688_, data_stage_1__687_, data_stage_1__686_, data_stage_1__685_, data_stage_1__684_, data_stage_1__683_, data_stage_1__682_, data_stage_1__681_, data_stage_1__680_, data_stage_1__679_, data_stage_1__678_, data_stage_1__677_, data_stage_1__676_, data_stage_1__675_, data_stage_1__674_, data_stage_1__673_, data_stage_1__672_, data_stage_1__671_, data_stage_1__670_, data_stage_1__669_, data_stage_1__668_, data_stage_1__667_, data_stage_1__666_, data_stage_1__665_, data_stage_1__664_, data_stage_1__663_, data_stage_1__662_, data_stage_1__661_, data_stage_1__660_, data_stage_1__659_, data_stage_1__658_, data_stage_1__657_, data_stage_1__656_, data_stage_1__655_, data_stage_1__654_, data_stage_1__653_, data_stage_1__652_, data_stage_1__651_, data_stage_1__650_, data_stage_1__649_, data_stage_1__648_, data_stage_1__647_, data_stage_1__646_, data_stage_1__645_, data_stage_1__644_, data_stage_1__643_, data_stage_1__642_, data_stage_1__641_, data_stage_1__640_, data_stage_1__639_, data_stage_1__638_, data_stage_1__637_, data_stage_1__636_, data_stage_1__635_, data_stage_1__634_, data_stage_1__633_, data_stage_1__632_, data_stage_1__631_, data_stage_1__630_, data_stage_1__629_, data_stage_1__628_, data_stage_1__627_, data_stage_1__626_, data_stage_1__625_, data_stage_1__624_, data_stage_1__623_, data_stage_1__622_, data_stage_1__621_, data_stage_1__620_, data_stage_1__619_, data_stage_1__618_, data_stage_1__617_, data_stage_1__616_, data_stage_1__615_, data_stage_1__614_, data_stage_1__613_, data_stage_1__612_, data_stage_1__611_, data_stage_1__610_, data_stage_1__609_, data_stage_1__608_, data_stage_1__607_, data_stage_1__606_, data_stage_1__605_, data_stage_1__604_, data_stage_1__603_, data_stage_1__602_, data_stage_1__601_, data_stage_1__600_, data_stage_1__599_, data_stage_1__598_, data_stage_1__597_, data_stage_1__596_, data_stage_1__595_, data_stage_1__594_, data_stage_1__593_, data_stage_1__592_, data_stage_1__591_, data_stage_1__590_, data_stage_1__589_, data_stage_1__588_, data_stage_1__587_, data_stage_1__586_, data_stage_1__585_, data_stage_1__584_, data_stage_1__583_, data_stage_1__582_, data_stage_1__581_, data_stage_1__580_, data_stage_1__579_, data_stage_1__578_, data_stage_1__577_, data_stage_1__576_, data_stage_1__575_, data_stage_1__574_, data_stage_1__573_, data_stage_1__572_, data_stage_1__571_, data_stage_1__570_, data_stage_1__569_, data_stage_1__568_, data_stage_1__567_, data_stage_1__566_, data_stage_1__565_, data_stage_1__564_, data_stage_1__563_, data_stage_1__562_, data_stage_1__561_, data_stage_1__560_, data_stage_1__559_, data_stage_1__558_, data_stage_1__557_, data_stage_1__556_, data_stage_1__555_, data_stage_1__554_, data_stage_1__553_, data_stage_1__552_, data_stage_1__551_, data_stage_1__550_, data_stage_1__549_, data_stage_1__548_, data_stage_1__547_, data_stage_1__546_, data_stage_1__545_, data_stage_1__544_, data_stage_1__543_, data_stage_1__542_, data_stage_1__541_, data_stage_1__540_, data_stage_1__539_, data_stage_1__538_, data_stage_1__537_, data_stage_1__536_, data_stage_1__535_, data_stage_1__534_, data_stage_1__533_, data_stage_1__532_, data_stage_1__531_, data_stage_1__530_, data_stage_1__529_, data_stage_1__528_, data_stage_1__527_, data_stage_1__526_, data_stage_1__525_, data_stage_1__524_, data_stage_1__523_, data_stage_1__522_, data_stage_1__521_, data_stage_1__520_, data_stage_1__519_, data_stage_1__518_, data_stage_1__517_, data_stage_1__516_, data_stage_1__515_, data_stage_1__514_, data_stage_1__513_, data_stage_1__512_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_3__swap_inst
  (
    .data_i(data_i[1023:768]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1023_, data_stage_1__1022_, data_stage_1__1021_, data_stage_1__1020_, data_stage_1__1019_, data_stage_1__1018_, data_stage_1__1017_, data_stage_1__1016_, data_stage_1__1015_, data_stage_1__1014_, data_stage_1__1013_, data_stage_1__1012_, data_stage_1__1011_, data_stage_1__1010_, data_stage_1__1009_, data_stage_1__1008_, data_stage_1__1007_, data_stage_1__1006_, data_stage_1__1005_, data_stage_1__1004_, data_stage_1__1003_, data_stage_1__1002_, data_stage_1__1001_, data_stage_1__1000_, data_stage_1__999_, data_stage_1__998_, data_stage_1__997_, data_stage_1__996_, data_stage_1__995_, data_stage_1__994_, data_stage_1__993_, data_stage_1__992_, data_stage_1__991_, data_stage_1__990_, data_stage_1__989_, data_stage_1__988_, data_stage_1__987_, data_stage_1__986_, data_stage_1__985_, data_stage_1__984_, data_stage_1__983_, data_stage_1__982_, data_stage_1__981_, data_stage_1__980_, data_stage_1__979_, data_stage_1__978_, data_stage_1__977_, data_stage_1__976_, data_stage_1__975_, data_stage_1__974_, data_stage_1__973_, data_stage_1__972_, data_stage_1__971_, data_stage_1__970_, data_stage_1__969_, data_stage_1__968_, data_stage_1__967_, data_stage_1__966_, data_stage_1__965_, data_stage_1__964_, data_stage_1__963_, data_stage_1__962_, data_stage_1__961_, data_stage_1__960_, data_stage_1__959_, data_stage_1__958_, data_stage_1__957_, data_stage_1__956_, data_stage_1__955_, data_stage_1__954_, data_stage_1__953_, data_stage_1__952_, data_stage_1__951_, data_stage_1__950_, data_stage_1__949_, data_stage_1__948_, data_stage_1__947_, data_stage_1__946_, data_stage_1__945_, data_stage_1__944_, data_stage_1__943_, data_stage_1__942_, data_stage_1__941_, data_stage_1__940_, data_stage_1__939_, data_stage_1__938_, data_stage_1__937_, data_stage_1__936_, data_stage_1__935_, data_stage_1__934_, data_stage_1__933_, data_stage_1__932_, data_stage_1__931_, data_stage_1__930_, data_stage_1__929_, data_stage_1__928_, data_stage_1__927_, data_stage_1__926_, data_stage_1__925_, data_stage_1__924_, data_stage_1__923_, data_stage_1__922_, data_stage_1__921_, data_stage_1__920_, data_stage_1__919_, data_stage_1__918_, data_stage_1__917_, data_stage_1__916_, data_stage_1__915_, data_stage_1__914_, data_stage_1__913_, data_stage_1__912_, data_stage_1__911_, data_stage_1__910_, data_stage_1__909_, data_stage_1__908_, data_stage_1__907_, data_stage_1__906_, data_stage_1__905_, data_stage_1__904_, data_stage_1__903_, data_stage_1__902_, data_stage_1__901_, data_stage_1__900_, data_stage_1__899_, data_stage_1__898_, data_stage_1__897_, data_stage_1__896_, data_stage_1__895_, data_stage_1__894_, data_stage_1__893_, data_stage_1__892_, data_stage_1__891_, data_stage_1__890_, data_stage_1__889_, data_stage_1__888_, data_stage_1__887_, data_stage_1__886_, data_stage_1__885_, data_stage_1__884_, data_stage_1__883_, data_stage_1__882_, data_stage_1__881_, data_stage_1__880_, data_stage_1__879_, data_stage_1__878_, data_stage_1__877_, data_stage_1__876_, data_stage_1__875_, data_stage_1__874_, data_stage_1__873_, data_stage_1__872_, data_stage_1__871_, data_stage_1__870_, data_stage_1__869_, data_stage_1__868_, data_stage_1__867_, data_stage_1__866_, data_stage_1__865_, data_stage_1__864_, data_stage_1__863_, data_stage_1__862_, data_stage_1__861_, data_stage_1__860_, data_stage_1__859_, data_stage_1__858_, data_stage_1__857_, data_stage_1__856_, data_stage_1__855_, data_stage_1__854_, data_stage_1__853_, data_stage_1__852_, data_stage_1__851_, data_stage_1__850_, data_stage_1__849_, data_stage_1__848_, data_stage_1__847_, data_stage_1__846_, data_stage_1__845_, data_stage_1__844_, data_stage_1__843_, data_stage_1__842_, data_stage_1__841_, data_stage_1__840_, data_stage_1__839_, data_stage_1__838_, data_stage_1__837_, data_stage_1__836_, data_stage_1__835_, data_stage_1__834_, data_stage_1__833_, data_stage_1__832_, data_stage_1__831_, data_stage_1__830_, data_stage_1__829_, data_stage_1__828_, data_stage_1__827_, data_stage_1__826_, data_stage_1__825_, data_stage_1__824_, data_stage_1__823_, data_stage_1__822_, data_stage_1__821_, data_stage_1__820_, data_stage_1__819_, data_stage_1__818_, data_stage_1__817_, data_stage_1__816_, data_stage_1__815_, data_stage_1__814_, data_stage_1__813_, data_stage_1__812_, data_stage_1__811_, data_stage_1__810_, data_stage_1__809_, data_stage_1__808_, data_stage_1__807_, data_stage_1__806_, data_stage_1__805_, data_stage_1__804_, data_stage_1__803_, data_stage_1__802_, data_stage_1__801_, data_stage_1__800_, data_stage_1__799_, data_stage_1__798_, data_stage_1__797_, data_stage_1__796_, data_stage_1__795_, data_stage_1__794_, data_stage_1__793_, data_stage_1__792_, data_stage_1__791_, data_stage_1__790_, data_stage_1__789_, data_stage_1__788_, data_stage_1__787_, data_stage_1__786_, data_stage_1__785_, data_stage_1__784_, data_stage_1__783_, data_stage_1__782_, data_stage_1__781_, data_stage_1__780_, data_stage_1__779_, data_stage_1__778_, data_stage_1__777_, data_stage_1__776_, data_stage_1__775_, data_stage_1__774_, data_stage_1__773_, data_stage_1__772_, data_stage_1__771_, data_stage_1__770_, data_stage_1__769_, data_stage_1__768_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_4__swap_inst
  (
    .data_i(data_i[1279:1024]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1279_, data_stage_1__1278_, data_stage_1__1277_, data_stage_1__1276_, data_stage_1__1275_, data_stage_1__1274_, data_stage_1__1273_, data_stage_1__1272_, data_stage_1__1271_, data_stage_1__1270_, data_stage_1__1269_, data_stage_1__1268_, data_stage_1__1267_, data_stage_1__1266_, data_stage_1__1265_, data_stage_1__1264_, data_stage_1__1263_, data_stage_1__1262_, data_stage_1__1261_, data_stage_1__1260_, data_stage_1__1259_, data_stage_1__1258_, data_stage_1__1257_, data_stage_1__1256_, data_stage_1__1255_, data_stage_1__1254_, data_stage_1__1253_, data_stage_1__1252_, data_stage_1__1251_, data_stage_1__1250_, data_stage_1__1249_, data_stage_1__1248_, data_stage_1__1247_, data_stage_1__1246_, data_stage_1__1245_, data_stage_1__1244_, data_stage_1__1243_, data_stage_1__1242_, data_stage_1__1241_, data_stage_1__1240_, data_stage_1__1239_, data_stage_1__1238_, data_stage_1__1237_, data_stage_1__1236_, data_stage_1__1235_, data_stage_1__1234_, data_stage_1__1233_, data_stage_1__1232_, data_stage_1__1231_, data_stage_1__1230_, data_stage_1__1229_, data_stage_1__1228_, data_stage_1__1227_, data_stage_1__1226_, data_stage_1__1225_, data_stage_1__1224_, data_stage_1__1223_, data_stage_1__1222_, data_stage_1__1221_, data_stage_1__1220_, data_stage_1__1219_, data_stage_1__1218_, data_stage_1__1217_, data_stage_1__1216_, data_stage_1__1215_, data_stage_1__1214_, data_stage_1__1213_, data_stage_1__1212_, data_stage_1__1211_, data_stage_1__1210_, data_stage_1__1209_, data_stage_1__1208_, data_stage_1__1207_, data_stage_1__1206_, data_stage_1__1205_, data_stage_1__1204_, data_stage_1__1203_, data_stage_1__1202_, data_stage_1__1201_, data_stage_1__1200_, data_stage_1__1199_, data_stage_1__1198_, data_stage_1__1197_, data_stage_1__1196_, data_stage_1__1195_, data_stage_1__1194_, data_stage_1__1193_, data_stage_1__1192_, data_stage_1__1191_, data_stage_1__1190_, data_stage_1__1189_, data_stage_1__1188_, data_stage_1__1187_, data_stage_1__1186_, data_stage_1__1185_, data_stage_1__1184_, data_stage_1__1183_, data_stage_1__1182_, data_stage_1__1181_, data_stage_1__1180_, data_stage_1__1179_, data_stage_1__1178_, data_stage_1__1177_, data_stage_1__1176_, data_stage_1__1175_, data_stage_1__1174_, data_stage_1__1173_, data_stage_1__1172_, data_stage_1__1171_, data_stage_1__1170_, data_stage_1__1169_, data_stage_1__1168_, data_stage_1__1167_, data_stage_1__1166_, data_stage_1__1165_, data_stage_1__1164_, data_stage_1__1163_, data_stage_1__1162_, data_stage_1__1161_, data_stage_1__1160_, data_stage_1__1159_, data_stage_1__1158_, data_stage_1__1157_, data_stage_1__1156_, data_stage_1__1155_, data_stage_1__1154_, data_stage_1__1153_, data_stage_1__1152_, data_stage_1__1151_, data_stage_1__1150_, data_stage_1__1149_, data_stage_1__1148_, data_stage_1__1147_, data_stage_1__1146_, data_stage_1__1145_, data_stage_1__1144_, data_stage_1__1143_, data_stage_1__1142_, data_stage_1__1141_, data_stage_1__1140_, data_stage_1__1139_, data_stage_1__1138_, data_stage_1__1137_, data_stage_1__1136_, data_stage_1__1135_, data_stage_1__1134_, data_stage_1__1133_, data_stage_1__1132_, data_stage_1__1131_, data_stage_1__1130_, data_stage_1__1129_, data_stage_1__1128_, data_stage_1__1127_, data_stage_1__1126_, data_stage_1__1125_, data_stage_1__1124_, data_stage_1__1123_, data_stage_1__1122_, data_stage_1__1121_, data_stage_1__1120_, data_stage_1__1119_, data_stage_1__1118_, data_stage_1__1117_, data_stage_1__1116_, data_stage_1__1115_, data_stage_1__1114_, data_stage_1__1113_, data_stage_1__1112_, data_stage_1__1111_, data_stage_1__1110_, data_stage_1__1109_, data_stage_1__1108_, data_stage_1__1107_, data_stage_1__1106_, data_stage_1__1105_, data_stage_1__1104_, data_stage_1__1103_, data_stage_1__1102_, data_stage_1__1101_, data_stage_1__1100_, data_stage_1__1099_, data_stage_1__1098_, data_stage_1__1097_, data_stage_1__1096_, data_stage_1__1095_, data_stage_1__1094_, data_stage_1__1093_, data_stage_1__1092_, data_stage_1__1091_, data_stage_1__1090_, data_stage_1__1089_, data_stage_1__1088_, data_stage_1__1087_, data_stage_1__1086_, data_stage_1__1085_, data_stage_1__1084_, data_stage_1__1083_, data_stage_1__1082_, data_stage_1__1081_, data_stage_1__1080_, data_stage_1__1079_, data_stage_1__1078_, data_stage_1__1077_, data_stage_1__1076_, data_stage_1__1075_, data_stage_1__1074_, data_stage_1__1073_, data_stage_1__1072_, data_stage_1__1071_, data_stage_1__1070_, data_stage_1__1069_, data_stage_1__1068_, data_stage_1__1067_, data_stage_1__1066_, data_stage_1__1065_, data_stage_1__1064_, data_stage_1__1063_, data_stage_1__1062_, data_stage_1__1061_, data_stage_1__1060_, data_stage_1__1059_, data_stage_1__1058_, data_stage_1__1057_, data_stage_1__1056_, data_stage_1__1055_, data_stage_1__1054_, data_stage_1__1053_, data_stage_1__1052_, data_stage_1__1051_, data_stage_1__1050_, data_stage_1__1049_, data_stage_1__1048_, data_stage_1__1047_, data_stage_1__1046_, data_stage_1__1045_, data_stage_1__1044_, data_stage_1__1043_, data_stage_1__1042_, data_stage_1__1041_, data_stage_1__1040_, data_stage_1__1039_, data_stage_1__1038_, data_stage_1__1037_, data_stage_1__1036_, data_stage_1__1035_, data_stage_1__1034_, data_stage_1__1033_, data_stage_1__1032_, data_stage_1__1031_, data_stage_1__1030_, data_stage_1__1029_, data_stage_1__1028_, data_stage_1__1027_, data_stage_1__1026_, data_stage_1__1025_, data_stage_1__1024_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_5__swap_inst
  (
    .data_i(data_i[1535:1280]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1535_, data_stage_1__1534_, data_stage_1__1533_, data_stage_1__1532_, data_stage_1__1531_, data_stage_1__1530_, data_stage_1__1529_, data_stage_1__1528_, data_stage_1__1527_, data_stage_1__1526_, data_stage_1__1525_, data_stage_1__1524_, data_stage_1__1523_, data_stage_1__1522_, data_stage_1__1521_, data_stage_1__1520_, data_stage_1__1519_, data_stage_1__1518_, data_stage_1__1517_, data_stage_1__1516_, data_stage_1__1515_, data_stage_1__1514_, data_stage_1__1513_, data_stage_1__1512_, data_stage_1__1511_, data_stage_1__1510_, data_stage_1__1509_, data_stage_1__1508_, data_stage_1__1507_, data_stage_1__1506_, data_stage_1__1505_, data_stage_1__1504_, data_stage_1__1503_, data_stage_1__1502_, data_stage_1__1501_, data_stage_1__1500_, data_stage_1__1499_, data_stage_1__1498_, data_stage_1__1497_, data_stage_1__1496_, data_stage_1__1495_, data_stage_1__1494_, data_stage_1__1493_, data_stage_1__1492_, data_stage_1__1491_, data_stage_1__1490_, data_stage_1__1489_, data_stage_1__1488_, data_stage_1__1487_, data_stage_1__1486_, data_stage_1__1485_, data_stage_1__1484_, data_stage_1__1483_, data_stage_1__1482_, data_stage_1__1481_, data_stage_1__1480_, data_stage_1__1479_, data_stage_1__1478_, data_stage_1__1477_, data_stage_1__1476_, data_stage_1__1475_, data_stage_1__1474_, data_stage_1__1473_, data_stage_1__1472_, data_stage_1__1471_, data_stage_1__1470_, data_stage_1__1469_, data_stage_1__1468_, data_stage_1__1467_, data_stage_1__1466_, data_stage_1__1465_, data_stage_1__1464_, data_stage_1__1463_, data_stage_1__1462_, data_stage_1__1461_, data_stage_1__1460_, data_stage_1__1459_, data_stage_1__1458_, data_stage_1__1457_, data_stage_1__1456_, data_stage_1__1455_, data_stage_1__1454_, data_stage_1__1453_, data_stage_1__1452_, data_stage_1__1451_, data_stage_1__1450_, data_stage_1__1449_, data_stage_1__1448_, data_stage_1__1447_, data_stage_1__1446_, data_stage_1__1445_, data_stage_1__1444_, data_stage_1__1443_, data_stage_1__1442_, data_stage_1__1441_, data_stage_1__1440_, data_stage_1__1439_, data_stage_1__1438_, data_stage_1__1437_, data_stage_1__1436_, data_stage_1__1435_, data_stage_1__1434_, data_stage_1__1433_, data_stage_1__1432_, data_stage_1__1431_, data_stage_1__1430_, data_stage_1__1429_, data_stage_1__1428_, data_stage_1__1427_, data_stage_1__1426_, data_stage_1__1425_, data_stage_1__1424_, data_stage_1__1423_, data_stage_1__1422_, data_stage_1__1421_, data_stage_1__1420_, data_stage_1__1419_, data_stage_1__1418_, data_stage_1__1417_, data_stage_1__1416_, data_stage_1__1415_, data_stage_1__1414_, data_stage_1__1413_, data_stage_1__1412_, data_stage_1__1411_, data_stage_1__1410_, data_stage_1__1409_, data_stage_1__1408_, data_stage_1__1407_, data_stage_1__1406_, data_stage_1__1405_, data_stage_1__1404_, data_stage_1__1403_, data_stage_1__1402_, data_stage_1__1401_, data_stage_1__1400_, data_stage_1__1399_, data_stage_1__1398_, data_stage_1__1397_, data_stage_1__1396_, data_stage_1__1395_, data_stage_1__1394_, data_stage_1__1393_, data_stage_1__1392_, data_stage_1__1391_, data_stage_1__1390_, data_stage_1__1389_, data_stage_1__1388_, data_stage_1__1387_, data_stage_1__1386_, data_stage_1__1385_, data_stage_1__1384_, data_stage_1__1383_, data_stage_1__1382_, data_stage_1__1381_, data_stage_1__1380_, data_stage_1__1379_, data_stage_1__1378_, data_stage_1__1377_, data_stage_1__1376_, data_stage_1__1375_, data_stage_1__1374_, data_stage_1__1373_, data_stage_1__1372_, data_stage_1__1371_, data_stage_1__1370_, data_stage_1__1369_, data_stage_1__1368_, data_stage_1__1367_, data_stage_1__1366_, data_stage_1__1365_, data_stage_1__1364_, data_stage_1__1363_, data_stage_1__1362_, data_stage_1__1361_, data_stage_1__1360_, data_stage_1__1359_, data_stage_1__1358_, data_stage_1__1357_, data_stage_1__1356_, data_stage_1__1355_, data_stage_1__1354_, data_stage_1__1353_, data_stage_1__1352_, data_stage_1__1351_, data_stage_1__1350_, data_stage_1__1349_, data_stage_1__1348_, data_stage_1__1347_, data_stage_1__1346_, data_stage_1__1345_, data_stage_1__1344_, data_stage_1__1343_, data_stage_1__1342_, data_stage_1__1341_, data_stage_1__1340_, data_stage_1__1339_, data_stage_1__1338_, data_stage_1__1337_, data_stage_1__1336_, data_stage_1__1335_, data_stage_1__1334_, data_stage_1__1333_, data_stage_1__1332_, data_stage_1__1331_, data_stage_1__1330_, data_stage_1__1329_, data_stage_1__1328_, data_stage_1__1327_, data_stage_1__1326_, data_stage_1__1325_, data_stage_1__1324_, data_stage_1__1323_, data_stage_1__1322_, data_stage_1__1321_, data_stage_1__1320_, data_stage_1__1319_, data_stage_1__1318_, data_stage_1__1317_, data_stage_1__1316_, data_stage_1__1315_, data_stage_1__1314_, data_stage_1__1313_, data_stage_1__1312_, data_stage_1__1311_, data_stage_1__1310_, data_stage_1__1309_, data_stage_1__1308_, data_stage_1__1307_, data_stage_1__1306_, data_stage_1__1305_, data_stage_1__1304_, data_stage_1__1303_, data_stage_1__1302_, data_stage_1__1301_, data_stage_1__1300_, data_stage_1__1299_, data_stage_1__1298_, data_stage_1__1297_, data_stage_1__1296_, data_stage_1__1295_, data_stage_1__1294_, data_stage_1__1293_, data_stage_1__1292_, data_stage_1__1291_, data_stage_1__1290_, data_stage_1__1289_, data_stage_1__1288_, data_stage_1__1287_, data_stage_1__1286_, data_stage_1__1285_, data_stage_1__1284_, data_stage_1__1283_, data_stage_1__1282_, data_stage_1__1281_, data_stage_1__1280_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_6__swap_inst
  (
    .data_i(data_i[1791:1536]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1791_, data_stage_1__1790_, data_stage_1__1789_, data_stage_1__1788_, data_stage_1__1787_, data_stage_1__1786_, data_stage_1__1785_, data_stage_1__1784_, data_stage_1__1783_, data_stage_1__1782_, data_stage_1__1781_, data_stage_1__1780_, data_stage_1__1779_, data_stage_1__1778_, data_stage_1__1777_, data_stage_1__1776_, data_stage_1__1775_, data_stage_1__1774_, data_stage_1__1773_, data_stage_1__1772_, data_stage_1__1771_, data_stage_1__1770_, data_stage_1__1769_, data_stage_1__1768_, data_stage_1__1767_, data_stage_1__1766_, data_stage_1__1765_, data_stage_1__1764_, data_stage_1__1763_, data_stage_1__1762_, data_stage_1__1761_, data_stage_1__1760_, data_stage_1__1759_, data_stage_1__1758_, data_stage_1__1757_, data_stage_1__1756_, data_stage_1__1755_, data_stage_1__1754_, data_stage_1__1753_, data_stage_1__1752_, data_stage_1__1751_, data_stage_1__1750_, data_stage_1__1749_, data_stage_1__1748_, data_stage_1__1747_, data_stage_1__1746_, data_stage_1__1745_, data_stage_1__1744_, data_stage_1__1743_, data_stage_1__1742_, data_stage_1__1741_, data_stage_1__1740_, data_stage_1__1739_, data_stage_1__1738_, data_stage_1__1737_, data_stage_1__1736_, data_stage_1__1735_, data_stage_1__1734_, data_stage_1__1733_, data_stage_1__1732_, data_stage_1__1731_, data_stage_1__1730_, data_stage_1__1729_, data_stage_1__1728_, data_stage_1__1727_, data_stage_1__1726_, data_stage_1__1725_, data_stage_1__1724_, data_stage_1__1723_, data_stage_1__1722_, data_stage_1__1721_, data_stage_1__1720_, data_stage_1__1719_, data_stage_1__1718_, data_stage_1__1717_, data_stage_1__1716_, data_stage_1__1715_, data_stage_1__1714_, data_stage_1__1713_, data_stage_1__1712_, data_stage_1__1711_, data_stage_1__1710_, data_stage_1__1709_, data_stage_1__1708_, data_stage_1__1707_, data_stage_1__1706_, data_stage_1__1705_, data_stage_1__1704_, data_stage_1__1703_, data_stage_1__1702_, data_stage_1__1701_, data_stage_1__1700_, data_stage_1__1699_, data_stage_1__1698_, data_stage_1__1697_, data_stage_1__1696_, data_stage_1__1695_, data_stage_1__1694_, data_stage_1__1693_, data_stage_1__1692_, data_stage_1__1691_, data_stage_1__1690_, data_stage_1__1689_, data_stage_1__1688_, data_stage_1__1687_, data_stage_1__1686_, data_stage_1__1685_, data_stage_1__1684_, data_stage_1__1683_, data_stage_1__1682_, data_stage_1__1681_, data_stage_1__1680_, data_stage_1__1679_, data_stage_1__1678_, data_stage_1__1677_, data_stage_1__1676_, data_stage_1__1675_, data_stage_1__1674_, data_stage_1__1673_, data_stage_1__1672_, data_stage_1__1671_, data_stage_1__1670_, data_stage_1__1669_, data_stage_1__1668_, data_stage_1__1667_, data_stage_1__1666_, data_stage_1__1665_, data_stage_1__1664_, data_stage_1__1663_, data_stage_1__1662_, data_stage_1__1661_, data_stage_1__1660_, data_stage_1__1659_, data_stage_1__1658_, data_stage_1__1657_, data_stage_1__1656_, data_stage_1__1655_, data_stage_1__1654_, data_stage_1__1653_, data_stage_1__1652_, data_stage_1__1651_, data_stage_1__1650_, data_stage_1__1649_, data_stage_1__1648_, data_stage_1__1647_, data_stage_1__1646_, data_stage_1__1645_, data_stage_1__1644_, data_stage_1__1643_, data_stage_1__1642_, data_stage_1__1641_, data_stage_1__1640_, data_stage_1__1639_, data_stage_1__1638_, data_stage_1__1637_, data_stage_1__1636_, data_stage_1__1635_, data_stage_1__1634_, data_stage_1__1633_, data_stage_1__1632_, data_stage_1__1631_, data_stage_1__1630_, data_stage_1__1629_, data_stage_1__1628_, data_stage_1__1627_, data_stage_1__1626_, data_stage_1__1625_, data_stage_1__1624_, data_stage_1__1623_, data_stage_1__1622_, data_stage_1__1621_, data_stage_1__1620_, data_stage_1__1619_, data_stage_1__1618_, data_stage_1__1617_, data_stage_1__1616_, data_stage_1__1615_, data_stage_1__1614_, data_stage_1__1613_, data_stage_1__1612_, data_stage_1__1611_, data_stage_1__1610_, data_stage_1__1609_, data_stage_1__1608_, data_stage_1__1607_, data_stage_1__1606_, data_stage_1__1605_, data_stage_1__1604_, data_stage_1__1603_, data_stage_1__1602_, data_stage_1__1601_, data_stage_1__1600_, data_stage_1__1599_, data_stage_1__1598_, data_stage_1__1597_, data_stage_1__1596_, data_stage_1__1595_, data_stage_1__1594_, data_stage_1__1593_, data_stage_1__1592_, data_stage_1__1591_, data_stage_1__1590_, data_stage_1__1589_, data_stage_1__1588_, data_stage_1__1587_, data_stage_1__1586_, data_stage_1__1585_, data_stage_1__1584_, data_stage_1__1583_, data_stage_1__1582_, data_stage_1__1581_, data_stage_1__1580_, data_stage_1__1579_, data_stage_1__1578_, data_stage_1__1577_, data_stage_1__1576_, data_stage_1__1575_, data_stage_1__1574_, data_stage_1__1573_, data_stage_1__1572_, data_stage_1__1571_, data_stage_1__1570_, data_stage_1__1569_, data_stage_1__1568_, data_stage_1__1567_, data_stage_1__1566_, data_stage_1__1565_, data_stage_1__1564_, data_stage_1__1563_, data_stage_1__1562_, data_stage_1__1561_, data_stage_1__1560_, data_stage_1__1559_, data_stage_1__1558_, data_stage_1__1557_, data_stage_1__1556_, data_stage_1__1555_, data_stage_1__1554_, data_stage_1__1553_, data_stage_1__1552_, data_stage_1__1551_, data_stage_1__1550_, data_stage_1__1549_, data_stage_1__1548_, data_stage_1__1547_, data_stage_1__1546_, data_stage_1__1545_, data_stage_1__1544_, data_stage_1__1543_, data_stage_1__1542_, data_stage_1__1541_, data_stage_1__1540_, data_stage_1__1539_, data_stage_1__1538_, data_stage_1__1537_, data_stage_1__1536_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_7__swap_inst
  (
    .data_i(data_i[2047:1792]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2047_, data_stage_1__2046_, data_stage_1__2045_, data_stage_1__2044_, data_stage_1__2043_, data_stage_1__2042_, data_stage_1__2041_, data_stage_1__2040_, data_stage_1__2039_, data_stage_1__2038_, data_stage_1__2037_, data_stage_1__2036_, data_stage_1__2035_, data_stage_1__2034_, data_stage_1__2033_, data_stage_1__2032_, data_stage_1__2031_, data_stage_1__2030_, data_stage_1__2029_, data_stage_1__2028_, data_stage_1__2027_, data_stage_1__2026_, data_stage_1__2025_, data_stage_1__2024_, data_stage_1__2023_, data_stage_1__2022_, data_stage_1__2021_, data_stage_1__2020_, data_stage_1__2019_, data_stage_1__2018_, data_stage_1__2017_, data_stage_1__2016_, data_stage_1__2015_, data_stage_1__2014_, data_stage_1__2013_, data_stage_1__2012_, data_stage_1__2011_, data_stage_1__2010_, data_stage_1__2009_, data_stage_1__2008_, data_stage_1__2007_, data_stage_1__2006_, data_stage_1__2005_, data_stage_1__2004_, data_stage_1__2003_, data_stage_1__2002_, data_stage_1__2001_, data_stage_1__2000_, data_stage_1__1999_, data_stage_1__1998_, data_stage_1__1997_, data_stage_1__1996_, data_stage_1__1995_, data_stage_1__1994_, data_stage_1__1993_, data_stage_1__1992_, data_stage_1__1991_, data_stage_1__1990_, data_stage_1__1989_, data_stage_1__1988_, data_stage_1__1987_, data_stage_1__1986_, data_stage_1__1985_, data_stage_1__1984_, data_stage_1__1983_, data_stage_1__1982_, data_stage_1__1981_, data_stage_1__1980_, data_stage_1__1979_, data_stage_1__1978_, data_stage_1__1977_, data_stage_1__1976_, data_stage_1__1975_, data_stage_1__1974_, data_stage_1__1973_, data_stage_1__1972_, data_stage_1__1971_, data_stage_1__1970_, data_stage_1__1969_, data_stage_1__1968_, data_stage_1__1967_, data_stage_1__1966_, data_stage_1__1965_, data_stage_1__1964_, data_stage_1__1963_, data_stage_1__1962_, data_stage_1__1961_, data_stage_1__1960_, data_stage_1__1959_, data_stage_1__1958_, data_stage_1__1957_, data_stage_1__1956_, data_stage_1__1955_, data_stage_1__1954_, data_stage_1__1953_, data_stage_1__1952_, data_stage_1__1951_, data_stage_1__1950_, data_stage_1__1949_, data_stage_1__1948_, data_stage_1__1947_, data_stage_1__1946_, data_stage_1__1945_, data_stage_1__1944_, data_stage_1__1943_, data_stage_1__1942_, data_stage_1__1941_, data_stage_1__1940_, data_stage_1__1939_, data_stage_1__1938_, data_stage_1__1937_, data_stage_1__1936_, data_stage_1__1935_, data_stage_1__1934_, data_stage_1__1933_, data_stage_1__1932_, data_stage_1__1931_, data_stage_1__1930_, data_stage_1__1929_, data_stage_1__1928_, data_stage_1__1927_, data_stage_1__1926_, data_stage_1__1925_, data_stage_1__1924_, data_stage_1__1923_, data_stage_1__1922_, data_stage_1__1921_, data_stage_1__1920_, data_stage_1__1919_, data_stage_1__1918_, data_stage_1__1917_, data_stage_1__1916_, data_stage_1__1915_, data_stage_1__1914_, data_stage_1__1913_, data_stage_1__1912_, data_stage_1__1911_, data_stage_1__1910_, data_stage_1__1909_, data_stage_1__1908_, data_stage_1__1907_, data_stage_1__1906_, data_stage_1__1905_, data_stage_1__1904_, data_stage_1__1903_, data_stage_1__1902_, data_stage_1__1901_, data_stage_1__1900_, data_stage_1__1899_, data_stage_1__1898_, data_stage_1__1897_, data_stage_1__1896_, data_stage_1__1895_, data_stage_1__1894_, data_stage_1__1893_, data_stage_1__1892_, data_stage_1__1891_, data_stage_1__1890_, data_stage_1__1889_, data_stage_1__1888_, data_stage_1__1887_, data_stage_1__1886_, data_stage_1__1885_, data_stage_1__1884_, data_stage_1__1883_, data_stage_1__1882_, data_stage_1__1881_, data_stage_1__1880_, data_stage_1__1879_, data_stage_1__1878_, data_stage_1__1877_, data_stage_1__1876_, data_stage_1__1875_, data_stage_1__1874_, data_stage_1__1873_, data_stage_1__1872_, data_stage_1__1871_, data_stage_1__1870_, data_stage_1__1869_, data_stage_1__1868_, data_stage_1__1867_, data_stage_1__1866_, data_stage_1__1865_, data_stage_1__1864_, data_stage_1__1863_, data_stage_1__1862_, data_stage_1__1861_, data_stage_1__1860_, data_stage_1__1859_, data_stage_1__1858_, data_stage_1__1857_, data_stage_1__1856_, data_stage_1__1855_, data_stage_1__1854_, data_stage_1__1853_, data_stage_1__1852_, data_stage_1__1851_, data_stage_1__1850_, data_stage_1__1849_, data_stage_1__1848_, data_stage_1__1847_, data_stage_1__1846_, data_stage_1__1845_, data_stage_1__1844_, data_stage_1__1843_, data_stage_1__1842_, data_stage_1__1841_, data_stage_1__1840_, data_stage_1__1839_, data_stage_1__1838_, data_stage_1__1837_, data_stage_1__1836_, data_stage_1__1835_, data_stage_1__1834_, data_stage_1__1833_, data_stage_1__1832_, data_stage_1__1831_, data_stage_1__1830_, data_stage_1__1829_, data_stage_1__1828_, data_stage_1__1827_, data_stage_1__1826_, data_stage_1__1825_, data_stage_1__1824_, data_stage_1__1823_, data_stage_1__1822_, data_stage_1__1821_, data_stage_1__1820_, data_stage_1__1819_, data_stage_1__1818_, data_stage_1__1817_, data_stage_1__1816_, data_stage_1__1815_, data_stage_1__1814_, data_stage_1__1813_, data_stage_1__1812_, data_stage_1__1811_, data_stage_1__1810_, data_stage_1__1809_, data_stage_1__1808_, data_stage_1__1807_, data_stage_1__1806_, data_stage_1__1805_, data_stage_1__1804_, data_stage_1__1803_, data_stage_1__1802_, data_stage_1__1801_, data_stage_1__1800_, data_stage_1__1799_, data_stage_1__1798_, data_stage_1__1797_, data_stage_1__1796_, data_stage_1__1795_, data_stage_1__1794_, data_stage_1__1793_, data_stage_1__1792_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_8__swap_inst
  (
    .data_i(data_i[2303:2048]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2303_, data_stage_1__2302_, data_stage_1__2301_, data_stage_1__2300_, data_stage_1__2299_, data_stage_1__2298_, data_stage_1__2297_, data_stage_1__2296_, data_stage_1__2295_, data_stage_1__2294_, data_stage_1__2293_, data_stage_1__2292_, data_stage_1__2291_, data_stage_1__2290_, data_stage_1__2289_, data_stage_1__2288_, data_stage_1__2287_, data_stage_1__2286_, data_stage_1__2285_, data_stage_1__2284_, data_stage_1__2283_, data_stage_1__2282_, data_stage_1__2281_, data_stage_1__2280_, data_stage_1__2279_, data_stage_1__2278_, data_stage_1__2277_, data_stage_1__2276_, data_stage_1__2275_, data_stage_1__2274_, data_stage_1__2273_, data_stage_1__2272_, data_stage_1__2271_, data_stage_1__2270_, data_stage_1__2269_, data_stage_1__2268_, data_stage_1__2267_, data_stage_1__2266_, data_stage_1__2265_, data_stage_1__2264_, data_stage_1__2263_, data_stage_1__2262_, data_stage_1__2261_, data_stage_1__2260_, data_stage_1__2259_, data_stage_1__2258_, data_stage_1__2257_, data_stage_1__2256_, data_stage_1__2255_, data_stage_1__2254_, data_stage_1__2253_, data_stage_1__2252_, data_stage_1__2251_, data_stage_1__2250_, data_stage_1__2249_, data_stage_1__2248_, data_stage_1__2247_, data_stage_1__2246_, data_stage_1__2245_, data_stage_1__2244_, data_stage_1__2243_, data_stage_1__2242_, data_stage_1__2241_, data_stage_1__2240_, data_stage_1__2239_, data_stage_1__2238_, data_stage_1__2237_, data_stage_1__2236_, data_stage_1__2235_, data_stage_1__2234_, data_stage_1__2233_, data_stage_1__2232_, data_stage_1__2231_, data_stage_1__2230_, data_stage_1__2229_, data_stage_1__2228_, data_stage_1__2227_, data_stage_1__2226_, data_stage_1__2225_, data_stage_1__2224_, data_stage_1__2223_, data_stage_1__2222_, data_stage_1__2221_, data_stage_1__2220_, data_stage_1__2219_, data_stage_1__2218_, data_stage_1__2217_, data_stage_1__2216_, data_stage_1__2215_, data_stage_1__2214_, data_stage_1__2213_, data_stage_1__2212_, data_stage_1__2211_, data_stage_1__2210_, data_stage_1__2209_, data_stage_1__2208_, data_stage_1__2207_, data_stage_1__2206_, data_stage_1__2205_, data_stage_1__2204_, data_stage_1__2203_, data_stage_1__2202_, data_stage_1__2201_, data_stage_1__2200_, data_stage_1__2199_, data_stage_1__2198_, data_stage_1__2197_, data_stage_1__2196_, data_stage_1__2195_, data_stage_1__2194_, data_stage_1__2193_, data_stage_1__2192_, data_stage_1__2191_, data_stage_1__2190_, data_stage_1__2189_, data_stage_1__2188_, data_stage_1__2187_, data_stage_1__2186_, data_stage_1__2185_, data_stage_1__2184_, data_stage_1__2183_, data_stage_1__2182_, data_stage_1__2181_, data_stage_1__2180_, data_stage_1__2179_, data_stage_1__2178_, data_stage_1__2177_, data_stage_1__2176_, data_stage_1__2175_, data_stage_1__2174_, data_stage_1__2173_, data_stage_1__2172_, data_stage_1__2171_, data_stage_1__2170_, data_stage_1__2169_, data_stage_1__2168_, data_stage_1__2167_, data_stage_1__2166_, data_stage_1__2165_, data_stage_1__2164_, data_stage_1__2163_, data_stage_1__2162_, data_stage_1__2161_, data_stage_1__2160_, data_stage_1__2159_, data_stage_1__2158_, data_stage_1__2157_, data_stage_1__2156_, data_stage_1__2155_, data_stage_1__2154_, data_stage_1__2153_, data_stage_1__2152_, data_stage_1__2151_, data_stage_1__2150_, data_stage_1__2149_, data_stage_1__2148_, data_stage_1__2147_, data_stage_1__2146_, data_stage_1__2145_, data_stage_1__2144_, data_stage_1__2143_, data_stage_1__2142_, data_stage_1__2141_, data_stage_1__2140_, data_stage_1__2139_, data_stage_1__2138_, data_stage_1__2137_, data_stage_1__2136_, data_stage_1__2135_, data_stage_1__2134_, data_stage_1__2133_, data_stage_1__2132_, data_stage_1__2131_, data_stage_1__2130_, data_stage_1__2129_, data_stage_1__2128_, data_stage_1__2127_, data_stage_1__2126_, data_stage_1__2125_, data_stage_1__2124_, data_stage_1__2123_, data_stage_1__2122_, data_stage_1__2121_, data_stage_1__2120_, data_stage_1__2119_, data_stage_1__2118_, data_stage_1__2117_, data_stage_1__2116_, data_stage_1__2115_, data_stage_1__2114_, data_stage_1__2113_, data_stage_1__2112_, data_stage_1__2111_, data_stage_1__2110_, data_stage_1__2109_, data_stage_1__2108_, data_stage_1__2107_, data_stage_1__2106_, data_stage_1__2105_, data_stage_1__2104_, data_stage_1__2103_, data_stage_1__2102_, data_stage_1__2101_, data_stage_1__2100_, data_stage_1__2099_, data_stage_1__2098_, data_stage_1__2097_, data_stage_1__2096_, data_stage_1__2095_, data_stage_1__2094_, data_stage_1__2093_, data_stage_1__2092_, data_stage_1__2091_, data_stage_1__2090_, data_stage_1__2089_, data_stage_1__2088_, data_stage_1__2087_, data_stage_1__2086_, data_stage_1__2085_, data_stage_1__2084_, data_stage_1__2083_, data_stage_1__2082_, data_stage_1__2081_, data_stage_1__2080_, data_stage_1__2079_, data_stage_1__2078_, data_stage_1__2077_, data_stage_1__2076_, data_stage_1__2075_, data_stage_1__2074_, data_stage_1__2073_, data_stage_1__2072_, data_stage_1__2071_, data_stage_1__2070_, data_stage_1__2069_, data_stage_1__2068_, data_stage_1__2067_, data_stage_1__2066_, data_stage_1__2065_, data_stage_1__2064_, data_stage_1__2063_, data_stage_1__2062_, data_stage_1__2061_, data_stage_1__2060_, data_stage_1__2059_, data_stage_1__2058_, data_stage_1__2057_, data_stage_1__2056_, data_stage_1__2055_, data_stage_1__2054_, data_stage_1__2053_, data_stage_1__2052_, data_stage_1__2051_, data_stage_1__2050_, data_stage_1__2049_, data_stage_1__2048_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_9__swap_inst
  (
    .data_i(data_i[2559:2304]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2559_, data_stage_1__2558_, data_stage_1__2557_, data_stage_1__2556_, data_stage_1__2555_, data_stage_1__2554_, data_stage_1__2553_, data_stage_1__2552_, data_stage_1__2551_, data_stage_1__2550_, data_stage_1__2549_, data_stage_1__2548_, data_stage_1__2547_, data_stage_1__2546_, data_stage_1__2545_, data_stage_1__2544_, data_stage_1__2543_, data_stage_1__2542_, data_stage_1__2541_, data_stage_1__2540_, data_stage_1__2539_, data_stage_1__2538_, data_stage_1__2537_, data_stage_1__2536_, data_stage_1__2535_, data_stage_1__2534_, data_stage_1__2533_, data_stage_1__2532_, data_stage_1__2531_, data_stage_1__2530_, data_stage_1__2529_, data_stage_1__2528_, data_stage_1__2527_, data_stage_1__2526_, data_stage_1__2525_, data_stage_1__2524_, data_stage_1__2523_, data_stage_1__2522_, data_stage_1__2521_, data_stage_1__2520_, data_stage_1__2519_, data_stage_1__2518_, data_stage_1__2517_, data_stage_1__2516_, data_stage_1__2515_, data_stage_1__2514_, data_stage_1__2513_, data_stage_1__2512_, data_stage_1__2511_, data_stage_1__2510_, data_stage_1__2509_, data_stage_1__2508_, data_stage_1__2507_, data_stage_1__2506_, data_stage_1__2505_, data_stage_1__2504_, data_stage_1__2503_, data_stage_1__2502_, data_stage_1__2501_, data_stage_1__2500_, data_stage_1__2499_, data_stage_1__2498_, data_stage_1__2497_, data_stage_1__2496_, data_stage_1__2495_, data_stage_1__2494_, data_stage_1__2493_, data_stage_1__2492_, data_stage_1__2491_, data_stage_1__2490_, data_stage_1__2489_, data_stage_1__2488_, data_stage_1__2487_, data_stage_1__2486_, data_stage_1__2485_, data_stage_1__2484_, data_stage_1__2483_, data_stage_1__2482_, data_stage_1__2481_, data_stage_1__2480_, data_stage_1__2479_, data_stage_1__2478_, data_stage_1__2477_, data_stage_1__2476_, data_stage_1__2475_, data_stage_1__2474_, data_stage_1__2473_, data_stage_1__2472_, data_stage_1__2471_, data_stage_1__2470_, data_stage_1__2469_, data_stage_1__2468_, data_stage_1__2467_, data_stage_1__2466_, data_stage_1__2465_, data_stage_1__2464_, data_stage_1__2463_, data_stage_1__2462_, data_stage_1__2461_, data_stage_1__2460_, data_stage_1__2459_, data_stage_1__2458_, data_stage_1__2457_, data_stage_1__2456_, data_stage_1__2455_, data_stage_1__2454_, data_stage_1__2453_, data_stage_1__2452_, data_stage_1__2451_, data_stage_1__2450_, data_stage_1__2449_, data_stage_1__2448_, data_stage_1__2447_, data_stage_1__2446_, data_stage_1__2445_, data_stage_1__2444_, data_stage_1__2443_, data_stage_1__2442_, data_stage_1__2441_, data_stage_1__2440_, data_stage_1__2439_, data_stage_1__2438_, data_stage_1__2437_, data_stage_1__2436_, data_stage_1__2435_, data_stage_1__2434_, data_stage_1__2433_, data_stage_1__2432_, data_stage_1__2431_, data_stage_1__2430_, data_stage_1__2429_, data_stage_1__2428_, data_stage_1__2427_, data_stage_1__2426_, data_stage_1__2425_, data_stage_1__2424_, data_stage_1__2423_, data_stage_1__2422_, data_stage_1__2421_, data_stage_1__2420_, data_stage_1__2419_, data_stage_1__2418_, data_stage_1__2417_, data_stage_1__2416_, data_stage_1__2415_, data_stage_1__2414_, data_stage_1__2413_, data_stage_1__2412_, data_stage_1__2411_, data_stage_1__2410_, data_stage_1__2409_, data_stage_1__2408_, data_stage_1__2407_, data_stage_1__2406_, data_stage_1__2405_, data_stage_1__2404_, data_stage_1__2403_, data_stage_1__2402_, data_stage_1__2401_, data_stage_1__2400_, data_stage_1__2399_, data_stage_1__2398_, data_stage_1__2397_, data_stage_1__2396_, data_stage_1__2395_, data_stage_1__2394_, data_stage_1__2393_, data_stage_1__2392_, data_stage_1__2391_, data_stage_1__2390_, data_stage_1__2389_, data_stage_1__2388_, data_stage_1__2387_, data_stage_1__2386_, data_stage_1__2385_, data_stage_1__2384_, data_stage_1__2383_, data_stage_1__2382_, data_stage_1__2381_, data_stage_1__2380_, data_stage_1__2379_, data_stage_1__2378_, data_stage_1__2377_, data_stage_1__2376_, data_stage_1__2375_, data_stage_1__2374_, data_stage_1__2373_, data_stage_1__2372_, data_stage_1__2371_, data_stage_1__2370_, data_stage_1__2369_, data_stage_1__2368_, data_stage_1__2367_, data_stage_1__2366_, data_stage_1__2365_, data_stage_1__2364_, data_stage_1__2363_, data_stage_1__2362_, data_stage_1__2361_, data_stage_1__2360_, data_stage_1__2359_, data_stage_1__2358_, data_stage_1__2357_, data_stage_1__2356_, data_stage_1__2355_, data_stage_1__2354_, data_stage_1__2353_, data_stage_1__2352_, data_stage_1__2351_, data_stage_1__2350_, data_stage_1__2349_, data_stage_1__2348_, data_stage_1__2347_, data_stage_1__2346_, data_stage_1__2345_, data_stage_1__2344_, data_stage_1__2343_, data_stage_1__2342_, data_stage_1__2341_, data_stage_1__2340_, data_stage_1__2339_, data_stage_1__2338_, data_stage_1__2337_, data_stage_1__2336_, data_stage_1__2335_, data_stage_1__2334_, data_stage_1__2333_, data_stage_1__2332_, data_stage_1__2331_, data_stage_1__2330_, data_stage_1__2329_, data_stage_1__2328_, data_stage_1__2327_, data_stage_1__2326_, data_stage_1__2325_, data_stage_1__2324_, data_stage_1__2323_, data_stage_1__2322_, data_stage_1__2321_, data_stage_1__2320_, data_stage_1__2319_, data_stage_1__2318_, data_stage_1__2317_, data_stage_1__2316_, data_stage_1__2315_, data_stage_1__2314_, data_stage_1__2313_, data_stage_1__2312_, data_stage_1__2311_, data_stage_1__2310_, data_stage_1__2309_, data_stage_1__2308_, data_stage_1__2307_, data_stage_1__2306_, data_stage_1__2305_, data_stage_1__2304_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_10__swap_inst
  (
    .data_i(data_i[2815:2560]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__2815_, data_stage_1__2814_, data_stage_1__2813_, data_stage_1__2812_, data_stage_1__2811_, data_stage_1__2810_, data_stage_1__2809_, data_stage_1__2808_, data_stage_1__2807_, data_stage_1__2806_, data_stage_1__2805_, data_stage_1__2804_, data_stage_1__2803_, data_stage_1__2802_, data_stage_1__2801_, data_stage_1__2800_, data_stage_1__2799_, data_stage_1__2798_, data_stage_1__2797_, data_stage_1__2796_, data_stage_1__2795_, data_stage_1__2794_, data_stage_1__2793_, data_stage_1__2792_, data_stage_1__2791_, data_stage_1__2790_, data_stage_1__2789_, data_stage_1__2788_, data_stage_1__2787_, data_stage_1__2786_, data_stage_1__2785_, data_stage_1__2784_, data_stage_1__2783_, data_stage_1__2782_, data_stage_1__2781_, data_stage_1__2780_, data_stage_1__2779_, data_stage_1__2778_, data_stage_1__2777_, data_stage_1__2776_, data_stage_1__2775_, data_stage_1__2774_, data_stage_1__2773_, data_stage_1__2772_, data_stage_1__2771_, data_stage_1__2770_, data_stage_1__2769_, data_stage_1__2768_, data_stage_1__2767_, data_stage_1__2766_, data_stage_1__2765_, data_stage_1__2764_, data_stage_1__2763_, data_stage_1__2762_, data_stage_1__2761_, data_stage_1__2760_, data_stage_1__2759_, data_stage_1__2758_, data_stage_1__2757_, data_stage_1__2756_, data_stage_1__2755_, data_stage_1__2754_, data_stage_1__2753_, data_stage_1__2752_, data_stage_1__2751_, data_stage_1__2750_, data_stage_1__2749_, data_stage_1__2748_, data_stage_1__2747_, data_stage_1__2746_, data_stage_1__2745_, data_stage_1__2744_, data_stage_1__2743_, data_stage_1__2742_, data_stage_1__2741_, data_stage_1__2740_, data_stage_1__2739_, data_stage_1__2738_, data_stage_1__2737_, data_stage_1__2736_, data_stage_1__2735_, data_stage_1__2734_, data_stage_1__2733_, data_stage_1__2732_, data_stage_1__2731_, data_stage_1__2730_, data_stage_1__2729_, data_stage_1__2728_, data_stage_1__2727_, data_stage_1__2726_, data_stage_1__2725_, data_stage_1__2724_, data_stage_1__2723_, data_stage_1__2722_, data_stage_1__2721_, data_stage_1__2720_, data_stage_1__2719_, data_stage_1__2718_, data_stage_1__2717_, data_stage_1__2716_, data_stage_1__2715_, data_stage_1__2714_, data_stage_1__2713_, data_stage_1__2712_, data_stage_1__2711_, data_stage_1__2710_, data_stage_1__2709_, data_stage_1__2708_, data_stage_1__2707_, data_stage_1__2706_, data_stage_1__2705_, data_stage_1__2704_, data_stage_1__2703_, data_stage_1__2702_, data_stage_1__2701_, data_stage_1__2700_, data_stage_1__2699_, data_stage_1__2698_, data_stage_1__2697_, data_stage_1__2696_, data_stage_1__2695_, data_stage_1__2694_, data_stage_1__2693_, data_stage_1__2692_, data_stage_1__2691_, data_stage_1__2690_, data_stage_1__2689_, data_stage_1__2688_, data_stage_1__2687_, data_stage_1__2686_, data_stage_1__2685_, data_stage_1__2684_, data_stage_1__2683_, data_stage_1__2682_, data_stage_1__2681_, data_stage_1__2680_, data_stage_1__2679_, data_stage_1__2678_, data_stage_1__2677_, data_stage_1__2676_, data_stage_1__2675_, data_stage_1__2674_, data_stage_1__2673_, data_stage_1__2672_, data_stage_1__2671_, data_stage_1__2670_, data_stage_1__2669_, data_stage_1__2668_, data_stage_1__2667_, data_stage_1__2666_, data_stage_1__2665_, data_stage_1__2664_, data_stage_1__2663_, data_stage_1__2662_, data_stage_1__2661_, data_stage_1__2660_, data_stage_1__2659_, data_stage_1__2658_, data_stage_1__2657_, data_stage_1__2656_, data_stage_1__2655_, data_stage_1__2654_, data_stage_1__2653_, data_stage_1__2652_, data_stage_1__2651_, data_stage_1__2650_, data_stage_1__2649_, data_stage_1__2648_, data_stage_1__2647_, data_stage_1__2646_, data_stage_1__2645_, data_stage_1__2644_, data_stage_1__2643_, data_stage_1__2642_, data_stage_1__2641_, data_stage_1__2640_, data_stage_1__2639_, data_stage_1__2638_, data_stage_1__2637_, data_stage_1__2636_, data_stage_1__2635_, data_stage_1__2634_, data_stage_1__2633_, data_stage_1__2632_, data_stage_1__2631_, data_stage_1__2630_, data_stage_1__2629_, data_stage_1__2628_, data_stage_1__2627_, data_stage_1__2626_, data_stage_1__2625_, data_stage_1__2624_, data_stage_1__2623_, data_stage_1__2622_, data_stage_1__2621_, data_stage_1__2620_, data_stage_1__2619_, data_stage_1__2618_, data_stage_1__2617_, data_stage_1__2616_, data_stage_1__2615_, data_stage_1__2614_, data_stage_1__2613_, data_stage_1__2612_, data_stage_1__2611_, data_stage_1__2610_, data_stage_1__2609_, data_stage_1__2608_, data_stage_1__2607_, data_stage_1__2606_, data_stage_1__2605_, data_stage_1__2604_, data_stage_1__2603_, data_stage_1__2602_, data_stage_1__2601_, data_stage_1__2600_, data_stage_1__2599_, data_stage_1__2598_, data_stage_1__2597_, data_stage_1__2596_, data_stage_1__2595_, data_stage_1__2594_, data_stage_1__2593_, data_stage_1__2592_, data_stage_1__2591_, data_stage_1__2590_, data_stage_1__2589_, data_stage_1__2588_, data_stage_1__2587_, data_stage_1__2586_, data_stage_1__2585_, data_stage_1__2584_, data_stage_1__2583_, data_stage_1__2582_, data_stage_1__2581_, data_stage_1__2580_, data_stage_1__2579_, data_stage_1__2578_, data_stage_1__2577_, data_stage_1__2576_, data_stage_1__2575_, data_stage_1__2574_, data_stage_1__2573_, data_stage_1__2572_, data_stage_1__2571_, data_stage_1__2570_, data_stage_1__2569_, data_stage_1__2568_, data_stage_1__2567_, data_stage_1__2566_, data_stage_1__2565_, data_stage_1__2564_, data_stage_1__2563_, data_stage_1__2562_, data_stage_1__2561_, data_stage_1__2560_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_11__swap_inst
  (
    .data_i(data_i[3071:2816]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3071_, data_stage_1__3070_, data_stage_1__3069_, data_stage_1__3068_, data_stage_1__3067_, data_stage_1__3066_, data_stage_1__3065_, data_stage_1__3064_, data_stage_1__3063_, data_stage_1__3062_, data_stage_1__3061_, data_stage_1__3060_, data_stage_1__3059_, data_stage_1__3058_, data_stage_1__3057_, data_stage_1__3056_, data_stage_1__3055_, data_stage_1__3054_, data_stage_1__3053_, data_stage_1__3052_, data_stage_1__3051_, data_stage_1__3050_, data_stage_1__3049_, data_stage_1__3048_, data_stage_1__3047_, data_stage_1__3046_, data_stage_1__3045_, data_stage_1__3044_, data_stage_1__3043_, data_stage_1__3042_, data_stage_1__3041_, data_stage_1__3040_, data_stage_1__3039_, data_stage_1__3038_, data_stage_1__3037_, data_stage_1__3036_, data_stage_1__3035_, data_stage_1__3034_, data_stage_1__3033_, data_stage_1__3032_, data_stage_1__3031_, data_stage_1__3030_, data_stage_1__3029_, data_stage_1__3028_, data_stage_1__3027_, data_stage_1__3026_, data_stage_1__3025_, data_stage_1__3024_, data_stage_1__3023_, data_stage_1__3022_, data_stage_1__3021_, data_stage_1__3020_, data_stage_1__3019_, data_stage_1__3018_, data_stage_1__3017_, data_stage_1__3016_, data_stage_1__3015_, data_stage_1__3014_, data_stage_1__3013_, data_stage_1__3012_, data_stage_1__3011_, data_stage_1__3010_, data_stage_1__3009_, data_stage_1__3008_, data_stage_1__3007_, data_stage_1__3006_, data_stage_1__3005_, data_stage_1__3004_, data_stage_1__3003_, data_stage_1__3002_, data_stage_1__3001_, data_stage_1__3000_, data_stage_1__2999_, data_stage_1__2998_, data_stage_1__2997_, data_stage_1__2996_, data_stage_1__2995_, data_stage_1__2994_, data_stage_1__2993_, data_stage_1__2992_, data_stage_1__2991_, data_stage_1__2990_, data_stage_1__2989_, data_stage_1__2988_, data_stage_1__2987_, data_stage_1__2986_, data_stage_1__2985_, data_stage_1__2984_, data_stage_1__2983_, data_stage_1__2982_, data_stage_1__2981_, data_stage_1__2980_, data_stage_1__2979_, data_stage_1__2978_, data_stage_1__2977_, data_stage_1__2976_, data_stage_1__2975_, data_stage_1__2974_, data_stage_1__2973_, data_stage_1__2972_, data_stage_1__2971_, data_stage_1__2970_, data_stage_1__2969_, data_stage_1__2968_, data_stage_1__2967_, data_stage_1__2966_, data_stage_1__2965_, data_stage_1__2964_, data_stage_1__2963_, data_stage_1__2962_, data_stage_1__2961_, data_stage_1__2960_, data_stage_1__2959_, data_stage_1__2958_, data_stage_1__2957_, data_stage_1__2956_, data_stage_1__2955_, data_stage_1__2954_, data_stage_1__2953_, data_stage_1__2952_, data_stage_1__2951_, data_stage_1__2950_, data_stage_1__2949_, data_stage_1__2948_, data_stage_1__2947_, data_stage_1__2946_, data_stage_1__2945_, data_stage_1__2944_, data_stage_1__2943_, data_stage_1__2942_, data_stage_1__2941_, data_stage_1__2940_, data_stage_1__2939_, data_stage_1__2938_, data_stage_1__2937_, data_stage_1__2936_, data_stage_1__2935_, data_stage_1__2934_, data_stage_1__2933_, data_stage_1__2932_, data_stage_1__2931_, data_stage_1__2930_, data_stage_1__2929_, data_stage_1__2928_, data_stage_1__2927_, data_stage_1__2926_, data_stage_1__2925_, data_stage_1__2924_, data_stage_1__2923_, data_stage_1__2922_, data_stage_1__2921_, data_stage_1__2920_, data_stage_1__2919_, data_stage_1__2918_, data_stage_1__2917_, data_stage_1__2916_, data_stage_1__2915_, data_stage_1__2914_, data_stage_1__2913_, data_stage_1__2912_, data_stage_1__2911_, data_stage_1__2910_, data_stage_1__2909_, data_stage_1__2908_, data_stage_1__2907_, data_stage_1__2906_, data_stage_1__2905_, data_stage_1__2904_, data_stage_1__2903_, data_stage_1__2902_, data_stage_1__2901_, data_stage_1__2900_, data_stage_1__2899_, data_stage_1__2898_, data_stage_1__2897_, data_stage_1__2896_, data_stage_1__2895_, data_stage_1__2894_, data_stage_1__2893_, data_stage_1__2892_, data_stage_1__2891_, data_stage_1__2890_, data_stage_1__2889_, data_stage_1__2888_, data_stage_1__2887_, data_stage_1__2886_, data_stage_1__2885_, data_stage_1__2884_, data_stage_1__2883_, data_stage_1__2882_, data_stage_1__2881_, data_stage_1__2880_, data_stage_1__2879_, data_stage_1__2878_, data_stage_1__2877_, data_stage_1__2876_, data_stage_1__2875_, data_stage_1__2874_, data_stage_1__2873_, data_stage_1__2872_, data_stage_1__2871_, data_stage_1__2870_, data_stage_1__2869_, data_stage_1__2868_, data_stage_1__2867_, data_stage_1__2866_, data_stage_1__2865_, data_stage_1__2864_, data_stage_1__2863_, data_stage_1__2862_, data_stage_1__2861_, data_stage_1__2860_, data_stage_1__2859_, data_stage_1__2858_, data_stage_1__2857_, data_stage_1__2856_, data_stage_1__2855_, data_stage_1__2854_, data_stage_1__2853_, data_stage_1__2852_, data_stage_1__2851_, data_stage_1__2850_, data_stage_1__2849_, data_stage_1__2848_, data_stage_1__2847_, data_stage_1__2846_, data_stage_1__2845_, data_stage_1__2844_, data_stage_1__2843_, data_stage_1__2842_, data_stage_1__2841_, data_stage_1__2840_, data_stage_1__2839_, data_stage_1__2838_, data_stage_1__2837_, data_stage_1__2836_, data_stage_1__2835_, data_stage_1__2834_, data_stage_1__2833_, data_stage_1__2832_, data_stage_1__2831_, data_stage_1__2830_, data_stage_1__2829_, data_stage_1__2828_, data_stage_1__2827_, data_stage_1__2826_, data_stage_1__2825_, data_stage_1__2824_, data_stage_1__2823_, data_stage_1__2822_, data_stage_1__2821_, data_stage_1__2820_, data_stage_1__2819_, data_stage_1__2818_, data_stage_1__2817_, data_stage_1__2816_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_12__swap_inst
  (
    .data_i(data_i[3327:3072]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3327_, data_stage_1__3326_, data_stage_1__3325_, data_stage_1__3324_, data_stage_1__3323_, data_stage_1__3322_, data_stage_1__3321_, data_stage_1__3320_, data_stage_1__3319_, data_stage_1__3318_, data_stage_1__3317_, data_stage_1__3316_, data_stage_1__3315_, data_stage_1__3314_, data_stage_1__3313_, data_stage_1__3312_, data_stage_1__3311_, data_stage_1__3310_, data_stage_1__3309_, data_stage_1__3308_, data_stage_1__3307_, data_stage_1__3306_, data_stage_1__3305_, data_stage_1__3304_, data_stage_1__3303_, data_stage_1__3302_, data_stage_1__3301_, data_stage_1__3300_, data_stage_1__3299_, data_stage_1__3298_, data_stage_1__3297_, data_stage_1__3296_, data_stage_1__3295_, data_stage_1__3294_, data_stage_1__3293_, data_stage_1__3292_, data_stage_1__3291_, data_stage_1__3290_, data_stage_1__3289_, data_stage_1__3288_, data_stage_1__3287_, data_stage_1__3286_, data_stage_1__3285_, data_stage_1__3284_, data_stage_1__3283_, data_stage_1__3282_, data_stage_1__3281_, data_stage_1__3280_, data_stage_1__3279_, data_stage_1__3278_, data_stage_1__3277_, data_stage_1__3276_, data_stage_1__3275_, data_stage_1__3274_, data_stage_1__3273_, data_stage_1__3272_, data_stage_1__3271_, data_stage_1__3270_, data_stage_1__3269_, data_stage_1__3268_, data_stage_1__3267_, data_stage_1__3266_, data_stage_1__3265_, data_stage_1__3264_, data_stage_1__3263_, data_stage_1__3262_, data_stage_1__3261_, data_stage_1__3260_, data_stage_1__3259_, data_stage_1__3258_, data_stage_1__3257_, data_stage_1__3256_, data_stage_1__3255_, data_stage_1__3254_, data_stage_1__3253_, data_stage_1__3252_, data_stage_1__3251_, data_stage_1__3250_, data_stage_1__3249_, data_stage_1__3248_, data_stage_1__3247_, data_stage_1__3246_, data_stage_1__3245_, data_stage_1__3244_, data_stage_1__3243_, data_stage_1__3242_, data_stage_1__3241_, data_stage_1__3240_, data_stage_1__3239_, data_stage_1__3238_, data_stage_1__3237_, data_stage_1__3236_, data_stage_1__3235_, data_stage_1__3234_, data_stage_1__3233_, data_stage_1__3232_, data_stage_1__3231_, data_stage_1__3230_, data_stage_1__3229_, data_stage_1__3228_, data_stage_1__3227_, data_stage_1__3226_, data_stage_1__3225_, data_stage_1__3224_, data_stage_1__3223_, data_stage_1__3222_, data_stage_1__3221_, data_stage_1__3220_, data_stage_1__3219_, data_stage_1__3218_, data_stage_1__3217_, data_stage_1__3216_, data_stage_1__3215_, data_stage_1__3214_, data_stage_1__3213_, data_stage_1__3212_, data_stage_1__3211_, data_stage_1__3210_, data_stage_1__3209_, data_stage_1__3208_, data_stage_1__3207_, data_stage_1__3206_, data_stage_1__3205_, data_stage_1__3204_, data_stage_1__3203_, data_stage_1__3202_, data_stage_1__3201_, data_stage_1__3200_, data_stage_1__3199_, data_stage_1__3198_, data_stage_1__3197_, data_stage_1__3196_, data_stage_1__3195_, data_stage_1__3194_, data_stage_1__3193_, data_stage_1__3192_, data_stage_1__3191_, data_stage_1__3190_, data_stage_1__3189_, data_stage_1__3188_, data_stage_1__3187_, data_stage_1__3186_, data_stage_1__3185_, data_stage_1__3184_, data_stage_1__3183_, data_stage_1__3182_, data_stage_1__3181_, data_stage_1__3180_, data_stage_1__3179_, data_stage_1__3178_, data_stage_1__3177_, data_stage_1__3176_, data_stage_1__3175_, data_stage_1__3174_, data_stage_1__3173_, data_stage_1__3172_, data_stage_1__3171_, data_stage_1__3170_, data_stage_1__3169_, data_stage_1__3168_, data_stage_1__3167_, data_stage_1__3166_, data_stage_1__3165_, data_stage_1__3164_, data_stage_1__3163_, data_stage_1__3162_, data_stage_1__3161_, data_stage_1__3160_, data_stage_1__3159_, data_stage_1__3158_, data_stage_1__3157_, data_stage_1__3156_, data_stage_1__3155_, data_stage_1__3154_, data_stage_1__3153_, data_stage_1__3152_, data_stage_1__3151_, data_stage_1__3150_, data_stage_1__3149_, data_stage_1__3148_, data_stage_1__3147_, data_stage_1__3146_, data_stage_1__3145_, data_stage_1__3144_, data_stage_1__3143_, data_stage_1__3142_, data_stage_1__3141_, data_stage_1__3140_, data_stage_1__3139_, data_stage_1__3138_, data_stage_1__3137_, data_stage_1__3136_, data_stage_1__3135_, data_stage_1__3134_, data_stage_1__3133_, data_stage_1__3132_, data_stage_1__3131_, data_stage_1__3130_, data_stage_1__3129_, data_stage_1__3128_, data_stage_1__3127_, data_stage_1__3126_, data_stage_1__3125_, data_stage_1__3124_, data_stage_1__3123_, data_stage_1__3122_, data_stage_1__3121_, data_stage_1__3120_, data_stage_1__3119_, data_stage_1__3118_, data_stage_1__3117_, data_stage_1__3116_, data_stage_1__3115_, data_stage_1__3114_, data_stage_1__3113_, data_stage_1__3112_, data_stage_1__3111_, data_stage_1__3110_, data_stage_1__3109_, data_stage_1__3108_, data_stage_1__3107_, data_stage_1__3106_, data_stage_1__3105_, data_stage_1__3104_, data_stage_1__3103_, data_stage_1__3102_, data_stage_1__3101_, data_stage_1__3100_, data_stage_1__3099_, data_stage_1__3098_, data_stage_1__3097_, data_stage_1__3096_, data_stage_1__3095_, data_stage_1__3094_, data_stage_1__3093_, data_stage_1__3092_, data_stage_1__3091_, data_stage_1__3090_, data_stage_1__3089_, data_stage_1__3088_, data_stage_1__3087_, data_stage_1__3086_, data_stage_1__3085_, data_stage_1__3084_, data_stage_1__3083_, data_stage_1__3082_, data_stage_1__3081_, data_stage_1__3080_, data_stage_1__3079_, data_stage_1__3078_, data_stage_1__3077_, data_stage_1__3076_, data_stage_1__3075_, data_stage_1__3074_, data_stage_1__3073_, data_stage_1__3072_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_13__swap_inst
  (
    .data_i(data_i[3583:3328]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3583_, data_stage_1__3582_, data_stage_1__3581_, data_stage_1__3580_, data_stage_1__3579_, data_stage_1__3578_, data_stage_1__3577_, data_stage_1__3576_, data_stage_1__3575_, data_stage_1__3574_, data_stage_1__3573_, data_stage_1__3572_, data_stage_1__3571_, data_stage_1__3570_, data_stage_1__3569_, data_stage_1__3568_, data_stage_1__3567_, data_stage_1__3566_, data_stage_1__3565_, data_stage_1__3564_, data_stage_1__3563_, data_stage_1__3562_, data_stage_1__3561_, data_stage_1__3560_, data_stage_1__3559_, data_stage_1__3558_, data_stage_1__3557_, data_stage_1__3556_, data_stage_1__3555_, data_stage_1__3554_, data_stage_1__3553_, data_stage_1__3552_, data_stage_1__3551_, data_stage_1__3550_, data_stage_1__3549_, data_stage_1__3548_, data_stage_1__3547_, data_stage_1__3546_, data_stage_1__3545_, data_stage_1__3544_, data_stage_1__3543_, data_stage_1__3542_, data_stage_1__3541_, data_stage_1__3540_, data_stage_1__3539_, data_stage_1__3538_, data_stage_1__3537_, data_stage_1__3536_, data_stage_1__3535_, data_stage_1__3534_, data_stage_1__3533_, data_stage_1__3532_, data_stage_1__3531_, data_stage_1__3530_, data_stage_1__3529_, data_stage_1__3528_, data_stage_1__3527_, data_stage_1__3526_, data_stage_1__3525_, data_stage_1__3524_, data_stage_1__3523_, data_stage_1__3522_, data_stage_1__3521_, data_stage_1__3520_, data_stage_1__3519_, data_stage_1__3518_, data_stage_1__3517_, data_stage_1__3516_, data_stage_1__3515_, data_stage_1__3514_, data_stage_1__3513_, data_stage_1__3512_, data_stage_1__3511_, data_stage_1__3510_, data_stage_1__3509_, data_stage_1__3508_, data_stage_1__3507_, data_stage_1__3506_, data_stage_1__3505_, data_stage_1__3504_, data_stage_1__3503_, data_stage_1__3502_, data_stage_1__3501_, data_stage_1__3500_, data_stage_1__3499_, data_stage_1__3498_, data_stage_1__3497_, data_stage_1__3496_, data_stage_1__3495_, data_stage_1__3494_, data_stage_1__3493_, data_stage_1__3492_, data_stage_1__3491_, data_stage_1__3490_, data_stage_1__3489_, data_stage_1__3488_, data_stage_1__3487_, data_stage_1__3486_, data_stage_1__3485_, data_stage_1__3484_, data_stage_1__3483_, data_stage_1__3482_, data_stage_1__3481_, data_stage_1__3480_, data_stage_1__3479_, data_stage_1__3478_, data_stage_1__3477_, data_stage_1__3476_, data_stage_1__3475_, data_stage_1__3474_, data_stage_1__3473_, data_stage_1__3472_, data_stage_1__3471_, data_stage_1__3470_, data_stage_1__3469_, data_stage_1__3468_, data_stage_1__3467_, data_stage_1__3466_, data_stage_1__3465_, data_stage_1__3464_, data_stage_1__3463_, data_stage_1__3462_, data_stage_1__3461_, data_stage_1__3460_, data_stage_1__3459_, data_stage_1__3458_, data_stage_1__3457_, data_stage_1__3456_, data_stage_1__3455_, data_stage_1__3454_, data_stage_1__3453_, data_stage_1__3452_, data_stage_1__3451_, data_stage_1__3450_, data_stage_1__3449_, data_stage_1__3448_, data_stage_1__3447_, data_stage_1__3446_, data_stage_1__3445_, data_stage_1__3444_, data_stage_1__3443_, data_stage_1__3442_, data_stage_1__3441_, data_stage_1__3440_, data_stage_1__3439_, data_stage_1__3438_, data_stage_1__3437_, data_stage_1__3436_, data_stage_1__3435_, data_stage_1__3434_, data_stage_1__3433_, data_stage_1__3432_, data_stage_1__3431_, data_stage_1__3430_, data_stage_1__3429_, data_stage_1__3428_, data_stage_1__3427_, data_stage_1__3426_, data_stage_1__3425_, data_stage_1__3424_, data_stage_1__3423_, data_stage_1__3422_, data_stage_1__3421_, data_stage_1__3420_, data_stage_1__3419_, data_stage_1__3418_, data_stage_1__3417_, data_stage_1__3416_, data_stage_1__3415_, data_stage_1__3414_, data_stage_1__3413_, data_stage_1__3412_, data_stage_1__3411_, data_stage_1__3410_, data_stage_1__3409_, data_stage_1__3408_, data_stage_1__3407_, data_stage_1__3406_, data_stage_1__3405_, data_stage_1__3404_, data_stage_1__3403_, data_stage_1__3402_, data_stage_1__3401_, data_stage_1__3400_, data_stage_1__3399_, data_stage_1__3398_, data_stage_1__3397_, data_stage_1__3396_, data_stage_1__3395_, data_stage_1__3394_, data_stage_1__3393_, data_stage_1__3392_, data_stage_1__3391_, data_stage_1__3390_, data_stage_1__3389_, data_stage_1__3388_, data_stage_1__3387_, data_stage_1__3386_, data_stage_1__3385_, data_stage_1__3384_, data_stage_1__3383_, data_stage_1__3382_, data_stage_1__3381_, data_stage_1__3380_, data_stage_1__3379_, data_stage_1__3378_, data_stage_1__3377_, data_stage_1__3376_, data_stage_1__3375_, data_stage_1__3374_, data_stage_1__3373_, data_stage_1__3372_, data_stage_1__3371_, data_stage_1__3370_, data_stage_1__3369_, data_stage_1__3368_, data_stage_1__3367_, data_stage_1__3366_, data_stage_1__3365_, data_stage_1__3364_, data_stage_1__3363_, data_stage_1__3362_, data_stage_1__3361_, data_stage_1__3360_, data_stage_1__3359_, data_stage_1__3358_, data_stage_1__3357_, data_stage_1__3356_, data_stage_1__3355_, data_stage_1__3354_, data_stage_1__3353_, data_stage_1__3352_, data_stage_1__3351_, data_stage_1__3350_, data_stage_1__3349_, data_stage_1__3348_, data_stage_1__3347_, data_stage_1__3346_, data_stage_1__3345_, data_stage_1__3344_, data_stage_1__3343_, data_stage_1__3342_, data_stage_1__3341_, data_stage_1__3340_, data_stage_1__3339_, data_stage_1__3338_, data_stage_1__3337_, data_stage_1__3336_, data_stage_1__3335_, data_stage_1__3334_, data_stage_1__3333_, data_stage_1__3332_, data_stage_1__3331_, data_stage_1__3330_, data_stage_1__3329_, data_stage_1__3328_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_14__swap_inst
  (
    .data_i(data_i[3839:3584]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__3839_, data_stage_1__3838_, data_stage_1__3837_, data_stage_1__3836_, data_stage_1__3835_, data_stage_1__3834_, data_stage_1__3833_, data_stage_1__3832_, data_stage_1__3831_, data_stage_1__3830_, data_stage_1__3829_, data_stage_1__3828_, data_stage_1__3827_, data_stage_1__3826_, data_stage_1__3825_, data_stage_1__3824_, data_stage_1__3823_, data_stage_1__3822_, data_stage_1__3821_, data_stage_1__3820_, data_stage_1__3819_, data_stage_1__3818_, data_stage_1__3817_, data_stage_1__3816_, data_stage_1__3815_, data_stage_1__3814_, data_stage_1__3813_, data_stage_1__3812_, data_stage_1__3811_, data_stage_1__3810_, data_stage_1__3809_, data_stage_1__3808_, data_stage_1__3807_, data_stage_1__3806_, data_stage_1__3805_, data_stage_1__3804_, data_stage_1__3803_, data_stage_1__3802_, data_stage_1__3801_, data_stage_1__3800_, data_stage_1__3799_, data_stage_1__3798_, data_stage_1__3797_, data_stage_1__3796_, data_stage_1__3795_, data_stage_1__3794_, data_stage_1__3793_, data_stage_1__3792_, data_stage_1__3791_, data_stage_1__3790_, data_stage_1__3789_, data_stage_1__3788_, data_stage_1__3787_, data_stage_1__3786_, data_stage_1__3785_, data_stage_1__3784_, data_stage_1__3783_, data_stage_1__3782_, data_stage_1__3781_, data_stage_1__3780_, data_stage_1__3779_, data_stage_1__3778_, data_stage_1__3777_, data_stage_1__3776_, data_stage_1__3775_, data_stage_1__3774_, data_stage_1__3773_, data_stage_1__3772_, data_stage_1__3771_, data_stage_1__3770_, data_stage_1__3769_, data_stage_1__3768_, data_stage_1__3767_, data_stage_1__3766_, data_stage_1__3765_, data_stage_1__3764_, data_stage_1__3763_, data_stage_1__3762_, data_stage_1__3761_, data_stage_1__3760_, data_stage_1__3759_, data_stage_1__3758_, data_stage_1__3757_, data_stage_1__3756_, data_stage_1__3755_, data_stage_1__3754_, data_stage_1__3753_, data_stage_1__3752_, data_stage_1__3751_, data_stage_1__3750_, data_stage_1__3749_, data_stage_1__3748_, data_stage_1__3747_, data_stage_1__3746_, data_stage_1__3745_, data_stage_1__3744_, data_stage_1__3743_, data_stage_1__3742_, data_stage_1__3741_, data_stage_1__3740_, data_stage_1__3739_, data_stage_1__3738_, data_stage_1__3737_, data_stage_1__3736_, data_stage_1__3735_, data_stage_1__3734_, data_stage_1__3733_, data_stage_1__3732_, data_stage_1__3731_, data_stage_1__3730_, data_stage_1__3729_, data_stage_1__3728_, data_stage_1__3727_, data_stage_1__3726_, data_stage_1__3725_, data_stage_1__3724_, data_stage_1__3723_, data_stage_1__3722_, data_stage_1__3721_, data_stage_1__3720_, data_stage_1__3719_, data_stage_1__3718_, data_stage_1__3717_, data_stage_1__3716_, data_stage_1__3715_, data_stage_1__3714_, data_stage_1__3713_, data_stage_1__3712_, data_stage_1__3711_, data_stage_1__3710_, data_stage_1__3709_, data_stage_1__3708_, data_stage_1__3707_, data_stage_1__3706_, data_stage_1__3705_, data_stage_1__3704_, data_stage_1__3703_, data_stage_1__3702_, data_stage_1__3701_, data_stage_1__3700_, data_stage_1__3699_, data_stage_1__3698_, data_stage_1__3697_, data_stage_1__3696_, data_stage_1__3695_, data_stage_1__3694_, data_stage_1__3693_, data_stage_1__3692_, data_stage_1__3691_, data_stage_1__3690_, data_stage_1__3689_, data_stage_1__3688_, data_stage_1__3687_, data_stage_1__3686_, data_stage_1__3685_, data_stage_1__3684_, data_stage_1__3683_, data_stage_1__3682_, data_stage_1__3681_, data_stage_1__3680_, data_stage_1__3679_, data_stage_1__3678_, data_stage_1__3677_, data_stage_1__3676_, data_stage_1__3675_, data_stage_1__3674_, data_stage_1__3673_, data_stage_1__3672_, data_stage_1__3671_, data_stage_1__3670_, data_stage_1__3669_, data_stage_1__3668_, data_stage_1__3667_, data_stage_1__3666_, data_stage_1__3665_, data_stage_1__3664_, data_stage_1__3663_, data_stage_1__3662_, data_stage_1__3661_, data_stage_1__3660_, data_stage_1__3659_, data_stage_1__3658_, data_stage_1__3657_, data_stage_1__3656_, data_stage_1__3655_, data_stage_1__3654_, data_stage_1__3653_, data_stage_1__3652_, data_stage_1__3651_, data_stage_1__3650_, data_stage_1__3649_, data_stage_1__3648_, data_stage_1__3647_, data_stage_1__3646_, data_stage_1__3645_, data_stage_1__3644_, data_stage_1__3643_, data_stage_1__3642_, data_stage_1__3641_, data_stage_1__3640_, data_stage_1__3639_, data_stage_1__3638_, data_stage_1__3637_, data_stage_1__3636_, data_stage_1__3635_, data_stage_1__3634_, data_stage_1__3633_, data_stage_1__3632_, data_stage_1__3631_, data_stage_1__3630_, data_stage_1__3629_, data_stage_1__3628_, data_stage_1__3627_, data_stage_1__3626_, data_stage_1__3625_, data_stage_1__3624_, data_stage_1__3623_, data_stage_1__3622_, data_stage_1__3621_, data_stage_1__3620_, data_stage_1__3619_, data_stage_1__3618_, data_stage_1__3617_, data_stage_1__3616_, data_stage_1__3615_, data_stage_1__3614_, data_stage_1__3613_, data_stage_1__3612_, data_stage_1__3611_, data_stage_1__3610_, data_stage_1__3609_, data_stage_1__3608_, data_stage_1__3607_, data_stage_1__3606_, data_stage_1__3605_, data_stage_1__3604_, data_stage_1__3603_, data_stage_1__3602_, data_stage_1__3601_, data_stage_1__3600_, data_stage_1__3599_, data_stage_1__3598_, data_stage_1__3597_, data_stage_1__3596_, data_stage_1__3595_, data_stage_1__3594_, data_stage_1__3593_, data_stage_1__3592_, data_stage_1__3591_, data_stage_1__3590_, data_stage_1__3589_, data_stage_1__3588_, data_stage_1__3587_, data_stage_1__3586_, data_stage_1__3585_, data_stage_1__3584_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_15__swap_inst
  (
    .data_i(data_i[4095:3840]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__4095_, data_stage_1__4094_, data_stage_1__4093_, data_stage_1__4092_, data_stage_1__4091_, data_stage_1__4090_, data_stage_1__4089_, data_stage_1__4088_, data_stage_1__4087_, data_stage_1__4086_, data_stage_1__4085_, data_stage_1__4084_, data_stage_1__4083_, data_stage_1__4082_, data_stage_1__4081_, data_stage_1__4080_, data_stage_1__4079_, data_stage_1__4078_, data_stage_1__4077_, data_stage_1__4076_, data_stage_1__4075_, data_stage_1__4074_, data_stage_1__4073_, data_stage_1__4072_, data_stage_1__4071_, data_stage_1__4070_, data_stage_1__4069_, data_stage_1__4068_, data_stage_1__4067_, data_stage_1__4066_, data_stage_1__4065_, data_stage_1__4064_, data_stage_1__4063_, data_stage_1__4062_, data_stage_1__4061_, data_stage_1__4060_, data_stage_1__4059_, data_stage_1__4058_, data_stage_1__4057_, data_stage_1__4056_, data_stage_1__4055_, data_stage_1__4054_, data_stage_1__4053_, data_stage_1__4052_, data_stage_1__4051_, data_stage_1__4050_, data_stage_1__4049_, data_stage_1__4048_, data_stage_1__4047_, data_stage_1__4046_, data_stage_1__4045_, data_stage_1__4044_, data_stage_1__4043_, data_stage_1__4042_, data_stage_1__4041_, data_stage_1__4040_, data_stage_1__4039_, data_stage_1__4038_, data_stage_1__4037_, data_stage_1__4036_, data_stage_1__4035_, data_stage_1__4034_, data_stage_1__4033_, data_stage_1__4032_, data_stage_1__4031_, data_stage_1__4030_, data_stage_1__4029_, data_stage_1__4028_, data_stage_1__4027_, data_stage_1__4026_, data_stage_1__4025_, data_stage_1__4024_, data_stage_1__4023_, data_stage_1__4022_, data_stage_1__4021_, data_stage_1__4020_, data_stage_1__4019_, data_stage_1__4018_, data_stage_1__4017_, data_stage_1__4016_, data_stage_1__4015_, data_stage_1__4014_, data_stage_1__4013_, data_stage_1__4012_, data_stage_1__4011_, data_stage_1__4010_, data_stage_1__4009_, data_stage_1__4008_, data_stage_1__4007_, data_stage_1__4006_, data_stage_1__4005_, data_stage_1__4004_, data_stage_1__4003_, data_stage_1__4002_, data_stage_1__4001_, data_stage_1__4000_, data_stage_1__3999_, data_stage_1__3998_, data_stage_1__3997_, data_stage_1__3996_, data_stage_1__3995_, data_stage_1__3994_, data_stage_1__3993_, data_stage_1__3992_, data_stage_1__3991_, data_stage_1__3990_, data_stage_1__3989_, data_stage_1__3988_, data_stage_1__3987_, data_stage_1__3986_, data_stage_1__3985_, data_stage_1__3984_, data_stage_1__3983_, data_stage_1__3982_, data_stage_1__3981_, data_stage_1__3980_, data_stage_1__3979_, data_stage_1__3978_, data_stage_1__3977_, data_stage_1__3976_, data_stage_1__3975_, data_stage_1__3974_, data_stage_1__3973_, data_stage_1__3972_, data_stage_1__3971_, data_stage_1__3970_, data_stage_1__3969_, data_stage_1__3968_, data_stage_1__3967_, data_stage_1__3966_, data_stage_1__3965_, data_stage_1__3964_, data_stage_1__3963_, data_stage_1__3962_, data_stage_1__3961_, data_stage_1__3960_, data_stage_1__3959_, data_stage_1__3958_, data_stage_1__3957_, data_stage_1__3956_, data_stage_1__3955_, data_stage_1__3954_, data_stage_1__3953_, data_stage_1__3952_, data_stage_1__3951_, data_stage_1__3950_, data_stage_1__3949_, data_stage_1__3948_, data_stage_1__3947_, data_stage_1__3946_, data_stage_1__3945_, data_stage_1__3944_, data_stage_1__3943_, data_stage_1__3942_, data_stage_1__3941_, data_stage_1__3940_, data_stage_1__3939_, data_stage_1__3938_, data_stage_1__3937_, data_stage_1__3936_, data_stage_1__3935_, data_stage_1__3934_, data_stage_1__3933_, data_stage_1__3932_, data_stage_1__3931_, data_stage_1__3930_, data_stage_1__3929_, data_stage_1__3928_, data_stage_1__3927_, data_stage_1__3926_, data_stage_1__3925_, data_stage_1__3924_, data_stage_1__3923_, data_stage_1__3922_, data_stage_1__3921_, data_stage_1__3920_, data_stage_1__3919_, data_stage_1__3918_, data_stage_1__3917_, data_stage_1__3916_, data_stage_1__3915_, data_stage_1__3914_, data_stage_1__3913_, data_stage_1__3912_, data_stage_1__3911_, data_stage_1__3910_, data_stage_1__3909_, data_stage_1__3908_, data_stage_1__3907_, data_stage_1__3906_, data_stage_1__3905_, data_stage_1__3904_, data_stage_1__3903_, data_stage_1__3902_, data_stage_1__3901_, data_stage_1__3900_, data_stage_1__3899_, data_stage_1__3898_, data_stage_1__3897_, data_stage_1__3896_, data_stage_1__3895_, data_stage_1__3894_, data_stage_1__3893_, data_stage_1__3892_, data_stage_1__3891_, data_stage_1__3890_, data_stage_1__3889_, data_stage_1__3888_, data_stage_1__3887_, data_stage_1__3886_, data_stage_1__3885_, data_stage_1__3884_, data_stage_1__3883_, data_stage_1__3882_, data_stage_1__3881_, data_stage_1__3880_, data_stage_1__3879_, data_stage_1__3878_, data_stage_1__3877_, data_stage_1__3876_, data_stage_1__3875_, data_stage_1__3874_, data_stage_1__3873_, data_stage_1__3872_, data_stage_1__3871_, data_stage_1__3870_, data_stage_1__3869_, data_stage_1__3868_, data_stage_1__3867_, data_stage_1__3866_, data_stage_1__3865_, data_stage_1__3864_, data_stage_1__3863_, data_stage_1__3862_, data_stage_1__3861_, data_stage_1__3860_, data_stage_1__3859_, data_stage_1__3858_, data_stage_1__3857_, data_stage_1__3856_, data_stage_1__3855_, data_stage_1__3854_, data_stage_1__3853_, data_stage_1__3852_, data_stage_1__3851_, data_stage_1__3850_, data_stage_1__3849_, data_stage_1__3848_, data_stage_1__3847_, data_stage_1__3846_, data_stage_1__3845_, data_stage_1__3844_, data_stage_1__3843_, data_stage_1__3842_, data_stage_1__3841_, data_stage_1__3840_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_16__swap_inst
  (
    .data_i(data_i[4351:4096]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__4351_, data_stage_1__4350_, data_stage_1__4349_, data_stage_1__4348_, data_stage_1__4347_, data_stage_1__4346_, data_stage_1__4345_, data_stage_1__4344_, data_stage_1__4343_, data_stage_1__4342_, data_stage_1__4341_, data_stage_1__4340_, data_stage_1__4339_, data_stage_1__4338_, data_stage_1__4337_, data_stage_1__4336_, data_stage_1__4335_, data_stage_1__4334_, data_stage_1__4333_, data_stage_1__4332_, data_stage_1__4331_, data_stage_1__4330_, data_stage_1__4329_, data_stage_1__4328_, data_stage_1__4327_, data_stage_1__4326_, data_stage_1__4325_, data_stage_1__4324_, data_stage_1__4323_, data_stage_1__4322_, data_stage_1__4321_, data_stage_1__4320_, data_stage_1__4319_, data_stage_1__4318_, data_stage_1__4317_, data_stage_1__4316_, data_stage_1__4315_, data_stage_1__4314_, data_stage_1__4313_, data_stage_1__4312_, data_stage_1__4311_, data_stage_1__4310_, data_stage_1__4309_, data_stage_1__4308_, data_stage_1__4307_, data_stage_1__4306_, data_stage_1__4305_, data_stage_1__4304_, data_stage_1__4303_, data_stage_1__4302_, data_stage_1__4301_, data_stage_1__4300_, data_stage_1__4299_, data_stage_1__4298_, data_stage_1__4297_, data_stage_1__4296_, data_stage_1__4295_, data_stage_1__4294_, data_stage_1__4293_, data_stage_1__4292_, data_stage_1__4291_, data_stage_1__4290_, data_stage_1__4289_, data_stage_1__4288_, data_stage_1__4287_, data_stage_1__4286_, data_stage_1__4285_, data_stage_1__4284_, data_stage_1__4283_, data_stage_1__4282_, data_stage_1__4281_, data_stage_1__4280_, data_stage_1__4279_, data_stage_1__4278_, data_stage_1__4277_, data_stage_1__4276_, data_stage_1__4275_, data_stage_1__4274_, data_stage_1__4273_, data_stage_1__4272_, data_stage_1__4271_, data_stage_1__4270_, data_stage_1__4269_, data_stage_1__4268_, data_stage_1__4267_, data_stage_1__4266_, data_stage_1__4265_, data_stage_1__4264_, data_stage_1__4263_, data_stage_1__4262_, data_stage_1__4261_, data_stage_1__4260_, data_stage_1__4259_, data_stage_1__4258_, data_stage_1__4257_, data_stage_1__4256_, data_stage_1__4255_, data_stage_1__4254_, data_stage_1__4253_, data_stage_1__4252_, data_stage_1__4251_, data_stage_1__4250_, data_stage_1__4249_, data_stage_1__4248_, data_stage_1__4247_, data_stage_1__4246_, data_stage_1__4245_, data_stage_1__4244_, data_stage_1__4243_, data_stage_1__4242_, data_stage_1__4241_, data_stage_1__4240_, data_stage_1__4239_, data_stage_1__4238_, data_stage_1__4237_, data_stage_1__4236_, data_stage_1__4235_, data_stage_1__4234_, data_stage_1__4233_, data_stage_1__4232_, data_stage_1__4231_, data_stage_1__4230_, data_stage_1__4229_, data_stage_1__4228_, data_stage_1__4227_, data_stage_1__4226_, data_stage_1__4225_, data_stage_1__4224_, data_stage_1__4223_, data_stage_1__4222_, data_stage_1__4221_, data_stage_1__4220_, data_stage_1__4219_, data_stage_1__4218_, data_stage_1__4217_, data_stage_1__4216_, data_stage_1__4215_, data_stage_1__4214_, data_stage_1__4213_, data_stage_1__4212_, data_stage_1__4211_, data_stage_1__4210_, data_stage_1__4209_, data_stage_1__4208_, data_stage_1__4207_, data_stage_1__4206_, data_stage_1__4205_, data_stage_1__4204_, data_stage_1__4203_, data_stage_1__4202_, data_stage_1__4201_, data_stage_1__4200_, data_stage_1__4199_, data_stage_1__4198_, data_stage_1__4197_, data_stage_1__4196_, data_stage_1__4195_, data_stage_1__4194_, data_stage_1__4193_, data_stage_1__4192_, data_stage_1__4191_, data_stage_1__4190_, data_stage_1__4189_, data_stage_1__4188_, data_stage_1__4187_, data_stage_1__4186_, data_stage_1__4185_, data_stage_1__4184_, data_stage_1__4183_, data_stage_1__4182_, data_stage_1__4181_, data_stage_1__4180_, data_stage_1__4179_, data_stage_1__4178_, data_stage_1__4177_, data_stage_1__4176_, data_stage_1__4175_, data_stage_1__4174_, data_stage_1__4173_, data_stage_1__4172_, data_stage_1__4171_, data_stage_1__4170_, data_stage_1__4169_, data_stage_1__4168_, data_stage_1__4167_, data_stage_1__4166_, data_stage_1__4165_, data_stage_1__4164_, data_stage_1__4163_, data_stage_1__4162_, data_stage_1__4161_, data_stage_1__4160_, data_stage_1__4159_, data_stage_1__4158_, data_stage_1__4157_, data_stage_1__4156_, data_stage_1__4155_, data_stage_1__4154_, data_stage_1__4153_, data_stage_1__4152_, data_stage_1__4151_, data_stage_1__4150_, data_stage_1__4149_, data_stage_1__4148_, data_stage_1__4147_, data_stage_1__4146_, data_stage_1__4145_, data_stage_1__4144_, data_stage_1__4143_, data_stage_1__4142_, data_stage_1__4141_, data_stage_1__4140_, data_stage_1__4139_, data_stage_1__4138_, data_stage_1__4137_, data_stage_1__4136_, data_stage_1__4135_, data_stage_1__4134_, data_stage_1__4133_, data_stage_1__4132_, data_stage_1__4131_, data_stage_1__4130_, data_stage_1__4129_, data_stage_1__4128_, data_stage_1__4127_, data_stage_1__4126_, data_stage_1__4125_, data_stage_1__4124_, data_stage_1__4123_, data_stage_1__4122_, data_stage_1__4121_, data_stage_1__4120_, data_stage_1__4119_, data_stage_1__4118_, data_stage_1__4117_, data_stage_1__4116_, data_stage_1__4115_, data_stage_1__4114_, data_stage_1__4113_, data_stage_1__4112_, data_stage_1__4111_, data_stage_1__4110_, data_stage_1__4109_, data_stage_1__4108_, data_stage_1__4107_, data_stage_1__4106_, data_stage_1__4105_, data_stage_1__4104_, data_stage_1__4103_, data_stage_1__4102_, data_stage_1__4101_, data_stage_1__4100_, data_stage_1__4099_, data_stage_1__4098_, data_stage_1__4097_, data_stage_1__4096_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_17__swap_inst
  (
    .data_i(data_i[4607:4352]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__4607_, data_stage_1__4606_, data_stage_1__4605_, data_stage_1__4604_, data_stage_1__4603_, data_stage_1__4602_, data_stage_1__4601_, data_stage_1__4600_, data_stage_1__4599_, data_stage_1__4598_, data_stage_1__4597_, data_stage_1__4596_, data_stage_1__4595_, data_stage_1__4594_, data_stage_1__4593_, data_stage_1__4592_, data_stage_1__4591_, data_stage_1__4590_, data_stage_1__4589_, data_stage_1__4588_, data_stage_1__4587_, data_stage_1__4586_, data_stage_1__4585_, data_stage_1__4584_, data_stage_1__4583_, data_stage_1__4582_, data_stage_1__4581_, data_stage_1__4580_, data_stage_1__4579_, data_stage_1__4578_, data_stage_1__4577_, data_stage_1__4576_, data_stage_1__4575_, data_stage_1__4574_, data_stage_1__4573_, data_stage_1__4572_, data_stage_1__4571_, data_stage_1__4570_, data_stage_1__4569_, data_stage_1__4568_, data_stage_1__4567_, data_stage_1__4566_, data_stage_1__4565_, data_stage_1__4564_, data_stage_1__4563_, data_stage_1__4562_, data_stage_1__4561_, data_stage_1__4560_, data_stage_1__4559_, data_stage_1__4558_, data_stage_1__4557_, data_stage_1__4556_, data_stage_1__4555_, data_stage_1__4554_, data_stage_1__4553_, data_stage_1__4552_, data_stage_1__4551_, data_stage_1__4550_, data_stage_1__4549_, data_stage_1__4548_, data_stage_1__4547_, data_stage_1__4546_, data_stage_1__4545_, data_stage_1__4544_, data_stage_1__4543_, data_stage_1__4542_, data_stage_1__4541_, data_stage_1__4540_, data_stage_1__4539_, data_stage_1__4538_, data_stage_1__4537_, data_stage_1__4536_, data_stage_1__4535_, data_stage_1__4534_, data_stage_1__4533_, data_stage_1__4532_, data_stage_1__4531_, data_stage_1__4530_, data_stage_1__4529_, data_stage_1__4528_, data_stage_1__4527_, data_stage_1__4526_, data_stage_1__4525_, data_stage_1__4524_, data_stage_1__4523_, data_stage_1__4522_, data_stage_1__4521_, data_stage_1__4520_, data_stage_1__4519_, data_stage_1__4518_, data_stage_1__4517_, data_stage_1__4516_, data_stage_1__4515_, data_stage_1__4514_, data_stage_1__4513_, data_stage_1__4512_, data_stage_1__4511_, data_stage_1__4510_, data_stage_1__4509_, data_stage_1__4508_, data_stage_1__4507_, data_stage_1__4506_, data_stage_1__4505_, data_stage_1__4504_, data_stage_1__4503_, data_stage_1__4502_, data_stage_1__4501_, data_stage_1__4500_, data_stage_1__4499_, data_stage_1__4498_, data_stage_1__4497_, data_stage_1__4496_, data_stage_1__4495_, data_stage_1__4494_, data_stage_1__4493_, data_stage_1__4492_, data_stage_1__4491_, data_stage_1__4490_, data_stage_1__4489_, data_stage_1__4488_, data_stage_1__4487_, data_stage_1__4486_, data_stage_1__4485_, data_stage_1__4484_, data_stage_1__4483_, data_stage_1__4482_, data_stage_1__4481_, data_stage_1__4480_, data_stage_1__4479_, data_stage_1__4478_, data_stage_1__4477_, data_stage_1__4476_, data_stage_1__4475_, data_stage_1__4474_, data_stage_1__4473_, data_stage_1__4472_, data_stage_1__4471_, data_stage_1__4470_, data_stage_1__4469_, data_stage_1__4468_, data_stage_1__4467_, data_stage_1__4466_, data_stage_1__4465_, data_stage_1__4464_, data_stage_1__4463_, data_stage_1__4462_, data_stage_1__4461_, data_stage_1__4460_, data_stage_1__4459_, data_stage_1__4458_, data_stage_1__4457_, data_stage_1__4456_, data_stage_1__4455_, data_stage_1__4454_, data_stage_1__4453_, data_stage_1__4452_, data_stage_1__4451_, data_stage_1__4450_, data_stage_1__4449_, data_stage_1__4448_, data_stage_1__4447_, data_stage_1__4446_, data_stage_1__4445_, data_stage_1__4444_, data_stage_1__4443_, data_stage_1__4442_, data_stage_1__4441_, data_stage_1__4440_, data_stage_1__4439_, data_stage_1__4438_, data_stage_1__4437_, data_stage_1__4436_, data_stage_1__4435_, data_stage_1__4434_, data_stage_1__4433_, data_stage_1__4432_, data_stage_1__4431_, data_stage_1__4430_, data_stage_1__4429_, data_stage_1__4428_, data_stage_1__4427_, data_stage_1__4426_, data_stage_1__4425_, data_stage_1__4424_, data_stage_1__4423_, data_stage_1__4422_, data_stage_1__4421_, data_stage_1__4420_, data_stage_1__4419_, data_stage_1__4418_, data_stage_1__4417_, data_stage_1__4416_, data_stage_1__4415_, data_stage_1__4414_, data_stage_1__4413_, data_stage_1__4412_, data_stage_1__4411_, data_stage_1__4410_, data_stage_1__4409_, data_stage_1__4408_, data_stage_1__4407_, data_stage_1__4406_, data_stage_1__4405_, data_stage_1__4404_, data_stage_1__4403_, data_stage_1__4402_, data_stage_1__4401_, data_stage_1__4400_, data_stage_1__4399_, data_stage_1__4398_, data_stage_1__4397_, data_stage_1__4396_, data_stage_1__4395_, data_stage_1__4394_, data_stage_1__4393_, data_stage_1__4392_, data_stage_1__4391_, data_stage_1__4390_, data_stage_1__4389_, data_stage_1__4388_, data_stage_1__4387_, data_stage_1__4386_, data_stage_1__4385_, data_stage_1__4384_, data_stage_1__4383_, data_stage_1__4382_, data_stage_1__4381_, data_stage_1__4380_, data_stage_1__4379_, data_stage_1__4378_, data_stage_1__4377_, data_stage_1__4376_, data_stage_1__4375_, data_stage_1__4374_, data_stage_1__4373_, data_stage_1__4372_, data_stage_1__4371_, data_stage_1__4370_, data_stage_1__4369_, data_stage_1__4368_, data_stage_1__4367_, data_stage_1__4366_, data_stage_1__4365_, data_stage_1__4364_, data_stage_1__4363_, data_stage_1__4362_, data_stage_1__4361_, data_stage_1__4360_, data_stage_1__4359_, data_stage_1__4358_, data_stage_1__4357_, data_stage_1__4356_, data_stage_1__4355_, data_stage_1__4354_, data_stage_1__4353_, data_stage_1__4352_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_18__swap_inst
  (
    .data_i(data_i[4863:4608]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__4863_, data_stage_1__4862_, data_stage_1__4861_, data_stage_1__4860_, data_stage_1__4859_, data_stage_1__4858_, data_stage_1__4857_, data_stage_1__4856_, data_stage_1__4855_, data_stage_1__4854_, data_stage_1__4853_, data_stage_1__4852_, data_stage_1__4851_, data_stage_1__4850_, data_stage_1__4849_, data_stage_1__4848_, data_stage_1__4847_, data_stage_1__4846_, data_stage_1__4845_, data_stage_1__4844_, data_stage_1__4843_, data_stage_1__4842_, data_stage_1__4841_, data_stage_1__4840_, data_stage_1__4839_, data_stage_1__4838_, data_stage_1__4837_, data_stage_1__4836_, data_stage_1__4835_, data_stage_1__4834_, data_stage_1__4833_, data_stage_1__4832_, data_stage_1__4831_, data_stage_1__4830_, data_stage_1__4829_, data_stage_1__4828_, data_stage_1__4827_, data_stage_1__4826_, data_stage_1__4825_, data_stage_1__4824_, data_stage_1__4823_, data_stage_1__4822_, data_stage_1__4821_, data_stage_1__4820_, data_stage_1__4819_, data_stage_1__4818_, data_stage_1__4817_, data_stage_1__4816_, data_stage_1__4815_, data_stage_1__4814_, data_stage_1__4813_, data_stage_1__4812_, data_stage_1__4811_, data_stage_1__4810_, data_stage_1__4809_, data_stage_1__4808_, data_stage_1__4807_, data_stage_1__4806_, data_stage_1__4805_, data_stage_1__4804_, data_stage_1__4803_, data_stage_1__4802_, data_stage_1__4801_, data_stage_1__4800_, data_stage_1__4799_, data_stage_1__4798_, data_stage_1__4797_, data_stage_1__4796_, data_stage_1__4795_, data_stage_1__4794_, data_stage_1__4793_, data_stage_1__4792_, data_stage_1__4791_, data_stage_1__4790_, data_stage_1__4789_, data_stage_1__4788_, data_stage_1__4787_, data_stage_1__4786_, data_stage_1__4785_, data_stage_1__4784_, data_stage_1__4783_, data_stage_1__4782_, data_stage_1__4781_, data_stage_1__4780_, data_stage_1__4779_, data_stage_1__4778_, data_stage_1__4777_, data_stage_1__4776_, data_stage_1__4775_, data_stage_1__4774_, data_stage_1__4773_, data_stage_1__4772_, data_stage_1__4771_, data_stage_1__4770_, data_stage_1__4769_, data_stage_1__4768_, data_stage_1__4767_, data_stage_1__4766_, data_stage_1__4765_, data_stage_1__4764_, data_stage_1__4763_, data_stage_1__4762_, data_stage_1__4761_, data_stage_1__4760_, data_stage_1__4759_, data_stage_1__4758_, data_stage_1__4757_, data_stage_1__4756_, data_stage_1__4755_, data_stage_1__4754_, data_stage_1__4753_, data_stage_1__4752_, data_stage_1__4751_, data_stage_1__4750_, data_stage_1__4749_, data_stage_1__4748_, data_stage_1__4747_, data_stage_1__4746_, data_stage_1__4745_, data_stage_1__4744_, data_stage_1__4743_, data_stage_1__4742_, data_stage_1__4741_, data_stage_1__4740_, data_stage_1__4739_, data_stage_1__4738_, data_stage_1__4737_, data_stage_1__4736_, data_stage_1__4735_, data_stage_1__4734_, data_stage_1__4733_, data_stage_1__4732_, data_stage_1__4731_, data_stage_1__4730_, data_stage_1__4729_, data_stage_1__4728_, data_stage_1__4727_, data_stage_1__4726_, data_stage_1__4725_, data_stage_1__4724_, data_stage_1__4723_, data_stage_1__4722_, data_stage_1__4721_, data_stage_1__4720_, data_stage_1__4719_, data_stage_1__4718_, data_stage_1__4717_, data_stage_1__4716_, data_stage_1__4715_, data_stage_1__4714_, data_stage_1__4713_, data_stage_1__4712_, data_stage_1__4711_, data_stage_1__4710_, data_stage_1__4709_, data_stage_1__4708_, data_stage_1__4707_, data_stage_1__4706_, data_stage_1__4705_, data_stage_1__4704_, data_stage_1__4703_, data_stage_1__4702_, data_stage_1__4701_, data_stage_1__4700_, data_stage_1__4699_, data_stage_1__4698_, data_stage_1__4697_, data_stage_1__4696_, data_stage_1__4695_, data_stage_1__4694_, data_stage_1__4693_, data_stage_1__4692_, data_stage_1__4691_, data_stage_1__4690_, data_stage_1__4689_, data_stage_1__4688_, data_stage_1__4687_, data_stage_1__4686_, data_stage_1__4685_, data_stage_1__4684_, data_stage_1__4683_, data_stage_1__4682_, data_stage_1__4681_, data_stage_1__4680_, data_stage_1__4679_, data_stage_1__4678_, data_stage_1__4677_, data_stage_1__4676_, data_stage_1__4675_, data_stage_1__4674_, data_stage_1__4673_, data_stage_1__4672_, data_stage_1__4671_, data_stage_1__4670_, data_stage_1__4669_, data_stage_1__4668_, data_stage_1__4667_, data_stage_1__4666_, data_stage_1__4665_, data_stage_1__4664_, data_stage_1__4663_, data_stage_1__4662_, data_stage_1__4661_, data_stage_1__4660_, data_stage_1__4659_, data_stage_1__4658_, data_stage_1__4657_, data_stage_1__4656_, data_stage_1__4655_, data_stage_1__4654_, data_stage_1__4653_, data_stage_1__4652_, data_stage_1__4651_, data_stage_1__4650_, data_stage_1__4649_, data_stage_1__4648_, data_stage_1__4647_, data_stage_1__4646_, data_stage_1__4645_, data_stage_1__4644_, data_stage_1__4643_, data_stage_1__4642_, data_stage_1__4641_, data_stage_1__4640_, data_stage_1__4639_, data_stage_1__4638_, data_stage_1__4637_, data_stage_1__4636_, data_stage_1__4635_, data_stage_1__4634_, data_stage_1__4633_, data_stage_1__4632_, data_stage_1__4631_, data_stage_1__4630_, data_stage_1__4629_, data_stage_1__4628_, data_stage_1__4627_, data_stage_1__4626_, data_stage_1__4625_, data_stage_1__4624_, data_stage_1__4623_, data_stage_1__4622_, data_stage_1__4621_, data_stage_1__4620_, data_stage_1__4619_, data_stage_1__4618_, data_stage_1__4617_, data_stage_1__4616_, data_stage_1__4615_, data_stage_1__4614_, data_stage_1__4613_, data_stage_1__4612_, data_stage_1__4611_, data_stage_1__4610_, data_stage_1__4609_, data_stage_1__4608_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_19__swap_inst
  (
    .data_i(data_i[5119:4864]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__5119_, data_stage_1__5118_, data_stage_1__5117_, data_stage_1__5116_, data_stage_1__5115_, data_stage_1__5114_, data_stage_1__5113_, data_stage_1__5112_, data_stage_1__5111_, data_stage_1__5110_, data_stage_1__5109_, data_stage_1__5108_, data_stage_1__5107_, data_stage_1__5106_, data_stage_1__5105_, data_stage_1__5104_, data_stage_1__5103_, data_stage_1__5102_, data_stage_1__5101_, data_stage_1__5100_, data_stage_1__5099_, data_stage_1__5098_, data_stage_1__5097_, data_stage_1__5096_, data_stage_1__5095_, data_stage_1__5094_, data_stage_1__5093_, data_stage_1__5092_, data_stage_1__5091_, data_stage_1__5090_, data_stage_1__5089_, data_stage_1__5088_, data_stage_1__5087_, data_stage_1__5086_, data_stage_1__5085_, data_stage_1__5084_, data_stage_1__5083_, data_stage_1__5082_, data_stage_1__5081_, data_stage_1__5080_, data_stage_1__5079_, data_stage_1__5078_, data_stage_1__5077_, data_stage_1__5076_, data_stage_1__5075_, data_stage_1__5074_, data_stage_1__5073_, data_stage_1__5072_, data_stage_1__5071_, data_stage_1__5070_, data_stage_1__5069_, data_stage_1__5068_, data_stage_1__5067_, data_stage_1__5066_, data_stage_1__5065_, data_stage_1__5064_, data_stage_1__5063_, data_stage_1__5062_, data_stage_1__5061_, data_stage_1__5060_, data_stage_1__5059_, data_stage_1__5058_, data_stage_1__5057_, data_stage_1__5056_, data_stage_1__5055_, data_stage_1__5054_, data_stage_1__5053_, data_stage_1__5052_, data_stage_1__5051_, data_stage_1__5050_, data_stage_1__5049_, data_stage_1__5048_, data_stage_1__5047_, data_stage_1__5046_, data_stage_1__5045_, data_stage_1__5044_, data_stage_1__5043_, data_stage_1__5042_, data_stage_1__5041_, data_stage_1__5040_, data_stage_1__5039_, data_stage_1__5038_, data_stage_1__5037_, data_stage_1__5036_, data_stage_1__5035_, data_stage_1__5034_, data_stage_1__5033_, data_stage_1__5032_, data_stage_1__5031_, data_stage_1__5030_, data_stage_1__5029_, data_stage_1__5028_, data_stage_1__5027_, data_stage_1__5026_, data_stage_1__5025_, data_stage_1__5024_, data_stage_1__5023_, data_stage_1__5022_, data_stage_1__5021_, data_stage_1__5020_, data_stage_1__5019_, data_stage_1__5018_, data_stage_1__5017_, data_stage_1__5016_, data_stage_1__5015_, data_stage_1__5014_, data_stage_1__5013_, data_stage_1__5012_, data_stage_1__5011_, data_stage_1__5010_, data_stage_1__5009_, data_stage_1__5008_, data_stage_1__5007_, data_stage_1__5006_, data_stage_1__5005_, data_stage_1__5004_, data_stage_1__5003_, data_stage_1__5002_, data_stage_1__5001_, data_stage_1__5000_, data_stage_1__4999_, data_stage_1__4998_, data_stage_1__4997_, data_stage_1__4996_, data_stage_1__4995_, data_stage_1__4994_, data_stage_1__4993_, data_stage_1__4992_, data_stage_1__4991_, data_stage_1__4990_, data_stage_1__4989_, data_stage_1__4988_, data_stage_1__4987_, data_stage_1__4986_, data_stage_1__4985_, data_stage_1__4984_, data_stage_1__4983_, data_stage_1__4982_, data_stage_1__4981_, data_stage_1__4980_, data_stage_1__4979_, data_stage_1__4978_, data_stage_1__4977_, data_stage_1__4976_, data_stage_1__4975_, data_stage_1__4974_, data_stage_1__4973_, data_stage_1__4972_, data_stage_1__4971_, data_stage_1__4970_, data_stage_1__4969_, data_stage_1__4968_, data_stage_1__4967_, data_stage_1__4966_, data_stage_1__4965_, data_stage_1__4964_, data_stage_1__4963_, data_stage_1__4962_, data_stage_1__4961_, data_stage_1__4960_, data_stage_1__4959_, data_stage_1__4958_, data_stage_1__4957_, data_stage_1__4956_, data_stage_1__4955_, data_stage_1__4954_, data_stage_1__4953_, data_stage_1__4952_, data_stage_1__4951_, data_stage_1__4950_, data_stage_1__4949_, data_stage_1__4948_, data_stage_1__4947_, data_stage_1__4946_, data_stage_1__4945_, data_stage_1__4944_, data_stage_1__4943_, data_stage_1__4942_, data_stage_1__4941_, data_stage_1__4940_, data_stage_1__4939_, data_stage_1__4938_, data_stage_1__4937_, data_stage_1__4936_, data_stage_1__4935_, data_stage_1__4934_, data_stage_1__4933_, data_stage_1__4932_, data_stage_1__4931_, data_stage_1__4930_, data_stage_1__4929_, data_stage_1__4928_, data_stage_1__4927_, data_stage_1__4926_, data_stage_1__4925_, data_stage_1__4924_, data_stage_1__4923_, data_stage_1__4922_, data_stage_1__4921_, data_stage_1__4920_, data_stage_1__4919_, data_stage_1__4918_, data_stage_1__4917_, data_stage_1__4916_, data_stage_1__4915_, data_stage_1__4914_, data_stage_1__4913_, data_stage_1__4912_, data_stage_1__4911_, data_stage_1__4910_, data_stage_1__4909_, data_stage_1__4908_, data_stage_1__4907_, data_stage_1__4906_, data_stage_1__4905_, data_stage_1__4904_, data_stage_1__4903_, data_stage_1__4902_, data_stage_1__4901_, data_stage_1__4900_, data_stage_1__4899_, data_stage_1__4898_, data_stage_1__4897_, data_stage_1__4896_, data_stage_1__4895_, data_stage_1__4894_, data_stage_1__4893_, data_stage_1__4892_, data_stage_1__4891_, data_stage_1__4890_, data_stage_1__4889_, data_stage_1__4888_, data_stage_1__4887_, data_stage_1__4886_, data_stage_1__4885_, data_stage_1__4884_, data_stage_1__4883_, data_stage_1__4882_, data_stage_1__4881_, data_stage_1__4880_, data_stage_1__4879_, data_stage_1__4878_, data_stage_1__4877_, data_stage_1__4876_, data_stage_1__4875_, data_stage_1__4874_, data_stage_1__4873_, data_stage_1__4872_, data_stage_1__4871_, data_stage_1__4870_, data_stage_1__4869_, data_stage_1__4868_, data_stage_1__4867_, data_stage_1__4866_, data_stage_1__4865_, data_stage_1__4864_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_20__swap_inst
  (
    .data_i(data_i[5375:5120]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__5375_, data_stage_1__5374_, data_stage_1__5373_, data_stage_1__5372_, data_stage_1__5371_, data_stage_1__5370_, data_stage_1__5369_, data_stage_1__5368_, data_stage_1__5367_, data_stage_1__5366_, data_stage_1__5365_, data_stage_1__5364_, data_stage_1__5363_, data_stage_1__5362_, data_stage_1__5361_, data_stage_1__5360_, data_stage_1__5359_, data_stage_1__5358_, data_stage_1__5357_, data_stage_1__5356_, data_stage_1__5355_, data_stage_1__5354_, data_stage_1__5353_, data_stage_1__5352_, data_stage_1__5351_, data_stage_1__5350_, data_stage_1__5349_, data_stage_1__5348_, data_stage_1__5347_, data_stage_1__5346_, data_stage_1__5345_, data_stage_1__5344_, data_stage_1__5343_, data_stage_1__5342_, data_stage_1__5341_, data_stage_1__5340_, data_stage_1__5339_, data_stage_1__5338_, data_stage_1__5337_, data_stage_1__5336_, data_stage_1__5335_, data_stage_1__5334_, data_stage_1__5333_, data_stage_1__5332_, data_stage_1__5331_, data_stage_1__5330_, data_stage_1__5329_, data_stage_1__5328_, data_stage_1__5327_, data_stage_1__5326_, data_stage_1__5325_, data_stage_1__5324_, data_stage_1__5323_, data_stage_1__5322_, data_stage_1__5321_, data_stage_1__5320_, data_stage_1__5319_, data_stage_1__5318_, data_stage_1__5317_, data_stage_1__5316_, data_stage_1__5315_, data_stage_1__5314_, data_stage_1__5313_, data_stage_1__5312_, data_stage_1__5311_, data_stage_1__5310_, data_stage_1__5309_, data_stage_1__5308_, data_stage_1__5307_, data_stage_1__5306_, data_stage_1__5305_, data_stage_1__5304_, data_stage_1__5303_, data_stage_1__5302_, data_stage_1__5301_, data_stage_1__5300_, data_stage_1__5299_, data_stage_1__5298_, data_stage_1__5297_, data_stage_1__5296_, data_stage_1__5295_, data_stage_1__5294_, data_stage_1__5293_, data_stage_1__5292_, data_stage_1__5291_, data_stage_1__5290_, data_stage_1__5289_, data_stage_1__5288_, data_stage_1__5287_, data_stage_1__5286_, data_stage_1__5285_, data_stage_1__5284_, data_stage_1__5283_, data_stage_1__5282_, data_stage_1__5281_, data_stage_1__5280_, data_stage_1__5279_, data_stage_1__5278_, data_stage_1__5277_, data_stage_1__5276_, data_stage_1__5275_, data_stage_1__5274_, data_stage_1__5273_, data_stage_1__5272_, data_stage_1__5271_, data_stage_1__5270_, data_stage_1__5269_, data_stage_1__5268_, data_stage_1__5267_, data_stage_1__5266_, data_stage_1__5265_, data_stage_1__5264_, data_stage_1__5263_, data_stage_1__5262_, data_stage_1__5261_, data_stage_1__5260_, data_stage_1__5259_, data_stage_1__5258_, data_stage_1__5257_, data_stage_1__5256_, data_stage_1__5255_, data_stage_1__5254_, data_stage_1__5253_, data_stage_1__5252_, data_stage_1__5251_, data_stage_1__5250_, data_stage_1__5249_, data_stage_1__5248_, data_stage_1__5247_, data_stage_1__5246_, data_stage_1__5245_, data_stage_1__5244_, data_stage_1__5243_, data_stage_1__5242_, data_stage_1__5241_, data_stage_1__5240_, data_stage_1__5239_, data_stage_1__5238_, data_stage_1__5237_, data_stage_1__5236_, data_stage_1__5235_, data_stage_1__5234_, data_stage_1__5233_, data_stage_1__5232_, data_stage_1__5231_, data_stage_1__5230_, data_stage_1__5229_, data_stage_1__5228_, data_stage_1__5227_, data_stage_1__5226_, data_stage_1__5225_, data_stage_1__5224_, data_stage_1__5223_, data_stage_1__5222_, data_stage_1__5221_, data_stage_1__5220_, data_stage_1__5219_, data_stage_1__5218_, data_stage_1__5217_, data_stage_1__5216_, data_stage_1__5215_, data_stage_1__5214_, data_stage_1__5213_, data_stage_1__5212_, data_stage_1__5211_, data_stage_1__5210_, data_stage_1__5209_, data_stage_1__5208_, data_stage_1__5207_, data_stage_1__5206_, data_stage_1__5205_, data_stage_1__5204_, data_stage_1__5203_, data_stage_1__5202_, data_stage_1__5201_, data_stage_1__5200_, data_stage_1__5199_, data_stage_1__5198_, data_stage_1__5197_, data_stage_1__5196_, data_stage_1__5195_, data_stage_1__5194_, data_stage_1__5193_, data_stage_1__5192_, data_stage_1__5191_, data_stage_1__5190_, data_stage_1__5189_, data_stage_1__5188_, data_stage_1__5187_, data_stage_1__5186_, data_stage_1__5185_, data_stage_1__5184_, data_stage_1__5183_, data_stage_1__5182_, data_stage_1__5181_, data_stage_1__5180_, data_stage_1__5179_, data_stage_1__5178_, data_stage_1__5177_, data_stage_1__5176_, data_stage_1__5175_, data_stage_1__5174_, data_stage_1__5173_, data_stage_1__5172_, data_stage_1__5171_, data_stage_1__5170_, data_stage_1__5169_, data_stage_1__5168_, data_stage_1__5167_, data_stage_1__5166_, data_stage_1__5165_, data_stage_1__5164_, data_stage_1__5163_, data_stage_1__5162_, data_stage_1__5161_, data_stage_1__5160_, data_stage_1__5159_, data_stage_1__5158_, data_stage_1__5157_, data_stage_1__5156_, data_stage_1__5155_, data_stage_1__5154_, data_stage_1__5153_, data_stage_1__5152_, data_stage_1__5151_, data_stage_1__5150_, data_stage_1__5149_, data_stage_1__5148_, data_stage_1__5147_, data_stage_1__5146_, data_stage_1__5145_, data_stage_1__5144_, data_stage_1__5143_, data_stage_1__5142_, data_stage_1__5141_, data_stage_1__5140_, data_stage_1__5139_, data_stage_1__5138_, data_stage_1__5137_, data_stage_1__5136_, data_stage_1__5135_, data_stage_1__5134_, data_stage_1__5133_, data_stage_1__5132_, data_stage_1__5131_, data_stage_1__5130_, data_stage_1__5129_, data_stage_1__5128_, data_stage_1__5127_, data_stage_1__5126_, data_stage_1__5125_, data_stage_1__5124_, data_stage_1__5123_, data_stage_1__5122_, data_stage_1__5121_, data_stage_1__5120_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_21__swap_inst
  (
    .data_i(data_i[5631:5376]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__5631_, data_stage_1__5630_, data_stage_1__5629_, data_stage_1__5628_, data_stage_1__5627_, data_stage_1__5626_, data_stage_1__5625_, data_stage_1__5624_, data_stage_1__5623_, data_stage_1__5622_, data_stage_1__5621_, data_stage_1__5620_, data_stage_1__5619_, data_stage_1__5618_, data_stage_1__5617_, data_stage_1__5616_, data_stage_1__5615_, data_stage_1__5614_, data_stage_1__5613_, data_stage_1__5612_, data_stage_1__5611_, data_stage_1__5610_, data_stage_1__5609_, data_stage_1__5608_, data_stage_1__5607_, data_stage_1__5606_, data_stage_1__5605_, data_stage_1__5604_, data_stage_1__5603_, data_stage_1__5602_, data_stage_1__5601_, data_stage_1__5600_, data_stage_1__5599_, data_stage_1__5598_, data_stage_1__5597_, data_stage_1__5596_, data_stage_1__5595_, data_stage_1__5594_, data_stage_1__5593_, data_stage_1__5592_, data_stage_1__5591_, data_stage_1__5590_, data_stage_1__5589_, data_stage_1__5588_, data_stage_1__5587_, data_stage_1__5586_, data_stage_1__5585_, data_stage_1__5584_, data_stage_1__5583_, data_stage_1__5582_, data_stage_1__5581_, data_stage_1__5580_, data_stage_1__5579_, data_stage_1__5578_, data_stage_1__5577_, data_stage_1__5576_, data_stage_1__5575_, data_stage_1__5574_, data_stage_1__5573_, data_stage_1__5572_, data_stage_1__5571_, data_stage_1__5570_, data_stage_1__5569_, data_stage_1__5568_, data_stage_1__5567_, data_stage_1__5566_, data_stage_1__5565_, data_stage_1__5564_, data_stage_1__5563_, data_stage_1__5562_, data_stage_1__5561_, data_stage_1__5560_, data_stage_1__5559_, data_stage_1__5558_, data_stage_1__5557_, data_stage_1__5556_, data_stage_1__5555_, data_stage_1__5554_, data_stage_1__5553_, data_stage_1__5552_, data_stage_1__5551_, data_stage_1__5550_, data_stage_1__5549_, data_stage_1__5548_, data_stage_1__5547_, data_stage_1__5546_, data_stage_1__5545_, data_stage_1__5544_, data_stage_1__5543_, data_stage_1__5542_, data_stage_1__5541_, data_stage_1__5540_, data_stage_1__5539_, data_stage_1__5538_, data_stage_1__5537_, data_stage_1__5536_, data_stage_1__5535_, data_stage_1__5534_, data_stage_1__5533_, data_stage_1__5532_, data_stage_1__5531_, data_stage_1__5530_, data_stage_1__5529_, data_stage_1__5528_, data_stage_1__5527_, data_stage_1__5526_, data_stage_1__5525_, data_stage_1__5524_, data_stage_1__5523_, data_stage_1__5522_, data_stage_1__5521_, data_stage_1__5520_, data_stage_1__5519_, data_stage_1__5518_, data_stage_1__5517_, data_stage_1__5516_, data_stage_1__5515_, data_stage_1__5514_, data_stage_1__5513_, data_stage_1__5512_, data_stage_1__5511_, data_stage_1__5510_, data_stage_1__5509_, data_stage_1__5508_, data_stage_1__5507_, data_stage_1__5506_, data_stage_1__5505_, data_stage_1__5504_, data_stage_1__5503_, data_stage_1__5502_, data_stage_1__5501_, data_stage_1__5500_, data_stage_1__5499_, data_stage_1__5498_, data_stage_1__5497_, data_stage_1__5496_, data_stage_1__5495_, data_stage_1__5494_, data_stage_1__5493_, data_stage_1__5492_, data_stage_1__5491_, data_stage_1__5490_, data_stage_1__5489_, data_stage_1__5488_, data_stage_1__5487_, data_stage_1__5486_, data_stage_1__5485_, data_stage_1__5484_, data_stage_1__5483_, data_stage_1__5482_, data_stage_1__5481_, data_stage_1__5480_, data_stage_1__5479_, data_stage_1__5478_, data_stage_1__5477_, data_stage_1__5476_, data_stage_1__5475_, data_stage_1__5474_, data_stage_1__5473_, data_stage_1__5472_, data_stage_1__5471_, data_stage_1__5470_, data_stage_1__5469_, data_stage_1__5468_, data_stage_1__5467_, data_stage_1__5466_, data_stage_1__5465_, data_stage_1__5464_, data_stage_1__5463_, data_stage_1__5462_, data_stage_1__5461_, data_stage_1__5460_, data_stage_1__5459_, data_stage_1__5458_, data_stage_1__5457_, data_stage_1__5456_, data_stage_1__5455_, data_stage_1__5454_, data_stage_1__5453_, data_stage_1__5452_, data_stage_1__5451_, data_stage_1__5450_, data_stage_1__5449_, data_stage_1__5448_, data_stage_1__5447_, data_stage_1__5446_, data_stage_1__5445_, data_stage_1__5444_, data_stage_1__5443_, data_stage_1__5442_, data_stage_1__5441_, data_stage_1__5440_, data_stage_1__5439_, data_stage_1__5438_, data_stage_1__5437_, data_stage_1__5436_, data_stage_1__5435_, data_stage_1__5434_, data_stage_1__5433_, data_stage_1__5432_, data_stage_1__5431_, data_stage_1__5430_, data_stage_1__5429_, data_stage_1__5428_, data_stage_1__5427_, data_stage_1__5426_, data_stage_1__5425_, data_stage_1__5424_, data_stage_1__5423_, data_stage_1__5422_, data_stage_1__5421_, data_stage_1__5420_, data_stage_1__5419_, data_stage_1__5418_, data_stage_1__5417_, data_stage_1__5416_, data_stage_1__5415_, data_stage_1__5414_, data_stage_1__5413_, data_stage_1__5412_, data_stage_1__5411_, data_stage_1__5410_, data_stage_1__5409_, data_stage_1__5408_, data_stage_1__5407_, data_stage_1__5406_, data_stage_1__5405_, data_stage_1__5404_, data_stage_1__5403_, data_stage_1__5402_, data_stage_1__5401_, data_stage_1__5400_, data_stage_1__5399_, data_stage_1__5398_, data_stage_1__5397_, data_stage_1__5396_, data_stage_1__5395_, data_stage_1__5394_, data_stage_1__5393_, data_stage_1__5392_, data_stage_1__5391_, data_stage_1__5390_, data_stage_1__5389_, data_stage_1__5388_, data_stage_1__5387_, data_stage_1__5386_, data_stage_1__5385_, data_stage_1__5384_, data_stage_1__5383_, data_stage_1__5382_, data_stage_1__5381_, data_stage_1__5380_, data_stage_1__5379_, data_stage_1__5378_, data_stage_1__5377_, data_stage_1__5376_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_22__swap_inst
  (
    .data_i(data_i[5887:5632]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__5887_, data_stage_1__5886_, data_stage_1__5885_, data_stage_1__5884_, data_stage_1__5883_, data_stage_1__5882_, data_stage_1__5881_, data_stage_1__5880_, data_stage_1__5879_, data_stage_1__5878_, data_stage_1__5877_, data_stage_1__5876_, data_stage_1__5875_, data_stage_1__5874_, data_stage_1__5873_, data_stage_1__5872_, data_stage_1__5871_, data_stage_1__5870_, data_stage_1__5869_, data_stage_1__5868_, data_stage_1__5867_, data_stage_1__5866_, data_stage_1__5865_, data_stage_1__5864_, data_stage_1__5863_, data_stage_1__5862_, data_stage_1__5861_, data_stage_1__5860_, data_stage_1__5859_, data_stage_1__5858_, data_stage_1__5857_, data_stage_1__5856_, data_stage_1__5855_, data_stage_1__5854_, data_stage_1__5853_, data_stage_1__5852_, data_stage_1__5851_, data_stage_1__5850_, data_stage_1__5849_, data_stage_1__5848_, data_stage_1__5847_, data_stage_1__5846_, data_stage_1__5845_, data_stage_1__5844_, data_stage_1__5843_, data_stage_1__5842_, data_stage_1__5841_, data_stage_1__5840_, data_stage_1__5839_, data_stage_1__5838_, data_stage_1__5837_, data_stage_1__5836_, data_stage_1__5835_, data_stage_1__5834_, data_stage_1__5833_, data_stage_1__5832_, data_stage_1__5831_, data_stage_1__5830_, data_stage_1__5829_, data_stage_1__5828_, data_stage_1__5827_, data_stage_1__5826_, data_stage_1__5825_, data_stage_1__5824_, data_stage_1__5823_, data_stage_1__5822_, data_stage_1__5821_, data_stage_1__5820_, data_stage_1__5819_, data_stage_1__5818_, data_stage_1__5817_, data_stage_1__5816_, data_stage_1__5815_, data_stage_1__5814_, data_stage_1__5813_, data_stage_1__5812_, data_stage_1__5811_, data_stage_1__5810_, data_stage_1__5809_, data_stage_1__5808_, data_stage_1__5807_, data_stage_1__5806_, data_stage_1__5805_, data_stage_1__5804_, data_stage_1__5803_, data_stage_1__5802_, data_stage_1__5801_, data_stage_1__5800_, data_stage_1__5799_, data_stage_1__5798_, data_stage_1__5797_, data_stage_1__5796_, data_stage_1__5795_, data_stage_1__5794_, data_stage_1__5793_, data_stage_1__5792_, data_stage_1__5791_, data_stage_1__5790_, data_stage_1__5789_, data_stage_1__5788_, data_stage_1__5787_, data_stage_1__5786_, data_stage_1__5785_, data_stage_1__5784_, data_stage_1__5783_, data_stage_1__5782_, data_stage_1__5781_, data_stage_1__5780_, data_stage_1__5779_, data_stage_1__5778_, data_stage_1__5777_, data_stage_1__5776_, data_stage_1__5775_, data_stage_1__5774_, data_stage_1__5773_, data_stage_1__5772_, data_stage_1__5771_, data_stage_1__5770_, data_stage_1__5769_, data_stage_1__5768_, data_stage_1__5767_, data_stage_1__5766_, data_stage_1__5765_, data_stage_1__5764_, data_stage_1__5763_, data_stage_1__5762_, data_stage_1__5761_, data_stage_1__5760_, data_stage_1__5759_, data_stage_1__5758_, data_stage_1__5757_, data_stage_1__5756_, data_stage_1__5755_, data_stage_1__5754_, data_stage_1__5753_, data_stage_1__5752_, data_stage_1__5751_, data_stage_1__5750_, data_stage_1__5749_, data_stage_1__5748_, data_stage_1__5747_, data_stage_1__5746_, data_stage_1__5745_, data_stage_1__5744_, data_stage_1__5743_, data_stage_1__5742_, data_stage_1__5741_, data_stage_1__5740_, data_stage_1__5739_, data_stage_1__5738_, data_stage_1__5737_, data_stage_1__5736_, data_stage_1__5735_, data_stage_1__5734_, data_stage_1__5733_, data_stage_1__5732_, data_stage_1__5731_, data_stage_1__5730_, data_stage_1__5729_, data_stage_1__5728_, data_stage_1__5727_, data_stage_1__5726_, data_stage_1__5725_, data_stage_1__5724_, data_stage_1__5723_, data_stage_1__5722_, data_stage_1__5721_, data_stage_1__5720_, data_stage_1__5719_, data_stage_1__5718_, data_stage_1__5717_, data_stage_1__5716_, data_stage_1__5715_, data_stage_1__5714_, data_stage_1__5713_, data_stage_1__5712_, data_stage_1__5711_, data_stage_1__5710_, data_stage_1__5709_, data_stage_1__5708_, data_stage_1__5707_, data_stage_1__5706_, data_stage_1__5705_, data_stage_1__5704_, data_stage_1__5703_, data_stage_1__5702_, data_stage_1__5701_, data_stage_1__5700_, data_stage_1__5699_, data_stage_1__5698_, data_stage_1__5697_, data_stage_1__5696_, data_stage_1__5695_, data_stage_1__5694_, data_stage_1__5693_, data_stage_1__5692_, data_stage_1__5691_, data_stage_1__5690_, data_stage_1__5689_, data_stage_1__5688_, data_stage_1__5687_, data_stage_1__5686_, data_stage_1__5685_, data_stage_1__5684_, data_stage_1__5683_, data_stage_1__5682_, data_stage_1__5681_, data_stage_1__5680_, data_stage_1__5679_, data_stage_1__5678_, data_stage_1__5677_, data_stage_1__5676_, data_stage_1__5675_, data_stage_1__5674_, data_stage_1__5673_, data_stage_1__5672_, data_stage_1__5671_, data_stage_1__5670_, data_stage_1__5669_, data_stage_1__5668_, data_stage_1__5667_, data_stage_1__5666_, data_stage_1__5665_, data_stage_1__5664_, data_stage_1__5663_, data_stage_1__5662_, data_stage_1__5661_, data_stage_1__5660_, data_stage_1__5659_, data_stage_1__5658_, data_stage_1__5657_, data_stage_1__5656_, data_stage_1__5655_, data_stage_1__5654_, data_stage_1__5653_, data_stage_1__5652_, data_stage_1__5651_, data_stage_1__5650_, data_stage_1__5649_, data_stage_1__5648_, data_stage_1__5647_, data_stage_1__5646_, data_stage_1__5645_, data_stage_1__5644_, data_stage_1__5643_, data_stage_1__5642_, data_stage_1__5641_, data_stage_1__5640_, data_stage_1__5639_, data_stage_1__5638_, data_stage_1__5637_, data_stage_1__5636_, data_stage_1__5635_, data_stage_1__5634_, data_stage_1__5633_, data_stage_1__5632_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_23__swap_inst
  (
    .data_i(data_i[6143:5888]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__6143_, data_stage_1__6142_, data_stage_1__6141_, data_stage_1__6140_, data_stage_1__6139_, data_stage_1__6138_, data_stage_1__6137_, data_stage_1__6136_, data_stage_1__6135_, data_stage_1__6134_, data_stage_1__6133_, data_stage_1__6132_, data_stage_1__6131_, data_stage_1__6130_, data_stage_1__6129_, data_stage_1__6128_, data_stage_1__6127_, data_stage_1__6126_, data_stage_1__6125_, data_stage_1__6124_, data_stage_1__6123_, data_stage_1__6122_, data_stage_1__6121_, data_stage_1__6120_, data_stage_1__6119_, data_stage_1__6118_, data_stage_1__6117_, data_stage_1__6116_, data_stage_1__6115_, data_stage_1__6114_, data_stage_1__6113_, data_stage_1__6112_, data_stage_1__6111_, data_stage_1__6110_, data_stage_1__6109_, data_stage_1__6108_, data_stage_1__6107_, data_stage_1__6106_, data_stage_1__6105_, data_stage_1__6104_, data_stage_1__6103_, data_stage_1__6102_, data_stage_1__6101_, data_stage_1__6100_, data_stage_1__6099_, data_stage_1__6098_, data_stage_1__6097_, data_stage_1__6096_, data_stage_1__6095_, data_stage_1__6094_, data_stage_1__6093_, data_stage_1__6092_, data_stage_1__6091_, data_stage_1__6090_, data_stage_1__6089_, data_stage_1__6088_, data_stage_1__6087_, data_stage_1__6086_, data_stage_1__6085_, data_stage_1__6084_, data_stage_1__6083_, data_stage_1__6082_, data_stage_1__6081_, data_stage_1__6080_, data_stage_1__6079_, data_stage_1__6078_, data_stage_1__6077_, data_stage_1__6076_, data_stage_1__6075_, data_stage_1__6074_, data_stage_1__6073_, data_stage_1__6072_, data_stage_1__6071_, data_stage_1__6070_, data_stage_1__6069_, data_stage_1__6068_, data_stage_1__6067_, data_stage_1__6066_, data_stage_1__6065_, data_stage_1__6064_, data_stage_1__6063_, data_stage_1__6062_, data_stage_1__6061_, data_stage_1__6060_, data_stage_1__6059_, data_stage_1__6058_, data_stage_1__6057_, data_stage_1__6056_, data_stage_1__6055_, data_stage_1__6054_, data_stage_1__6053_, data_stage_1__6052_, data_stage_1__6051_, data_stage_1__6050_, data_stage_1__6049_, data_stage_1__6048_, data_stage_1__6047_, data_stage_1__6046_, data_stage_1__6045_, data_stage_1__6044_, data_stage_1__6043_, data_stage_1__6042_, data_stage_1__6041_, data_stage_1__6040_, data_stage_1__6039_, data_stage_1__6038_, data_stage_1__6037_, data_stage_1__6036_, data_stage_1__6035_, data_stage_1__6034_, data_stage_1__6033_, data_stage_1__6032_, data_stage_1__6031_, data_stage_1__6030_, data_stage_1__6029_, data_stage_1__6028_, data_stage_1__6027_, data_stage_1__6026_, data_stage_1__6025_, data_stage_1__6024_, data_stage_1__6023_, data_stage_1__6022_, data_stage_1__6021_, data_stage_1__6020_, data_stage_1__6019_, data_stage_1__6018_, data_stage_1__6017_, data_stage_1__6016_, data_stage_1__6015_, data_stage_1__6014_, data_stage_1__6013_, data_stage_1__6012_, data_stage_1__6011_, data_stage_1__6010_, data_stage_1__6009_, data_stage_1__6008_, data_stage_1__6007_, data_stage_1__6006_, data_stage_1__6005_, data_stage_1__6004_, data_stage_1__6003_, data_stage_1__6002_, data_stage_1__6001_, data_stage_1__6000_, data_stage_1__5999_, data_stage_1__5998_, data_stage_1__5997_, data_stage_1__5996_, data_stage_1__5995_, data_stage_1__5994_, data_stage_1__5993_, data_stage_1__5992_, data_stage_1__5991_, data_stage_1__5990_, data_stage_1__5989_, data_stage_1__5988_, data_stage_1__5987_, data_stage_1__5986_, data_stage_1__5985_, data_stage_1__5984_, data_stage_1__5983_, data_stage_1__5982_, data_stage_1__5981_, data_stage_1__5980_, data_stage_1__5979_, data_stage_1__5978_, data_stage_1__5977_, data_stage_1__5976_, data_stage_1__5975_, data_stage_1__5974_, data_stage_1__5973_, data_stage_1__5972_, data_stage_1__5971_, data_stage_1__5970_, data_stage_1__5969_, data_stage_1__5968_, data_stage_1__5967_, data_stage_1__5966_, data_stage_1__5965_, data_stage_1__5964_, data_stage_1__5963_, data_stage_1__5962_, data_stage_1__5961_, data_stage_1__5960_, data_stage_1__5959_, data_stage_1__5958_, data_stage_1__5957_, data_stage_1__5956_, data_stage_1__5955_, data_stage_1__5954_, data_stage_1__5953_, data_stage_1__5952_, data_stage_1__5951_, data_stage_1__5950_, data_stage_1__5949_, data_stage_1__5948_, data_stage_1__5947_, data_stage_1__5946_, data_stage_1__5945_, data_stage_1__5944_, data_stage_1__5943_, data_stage_1__5942_, data_stage_1__5941_, data_stage_1__5940_, data_stage_1__5939_, data_stage_1__5938_, data_stage_1__5937_, data_stage_1__5936_, data_stage_1__5935_, data_stage_1__5934_, data_stage_1__5933_, data_stage_1__5932_, data_stage_1__5931_, data_stage_1__5930_, data_stage_1__5929_, data_stage_1__5928_, data_stage_1__5927_, data_stage_1__5926_, data_stage_1__5925_, data_stage_1__5924_, data_stage_1__5923_, data_stage_1__5922_, data_stage_1__5921_, data_stage_1__5920_, data_stage_1__5919_, data_stage_1__5918_, data_stage_1__5917_, data_stage_1__5916_, data_stage_1__5915_, data_stage_1__5914_, data_stage_1__5913_, data_stage_1__5912_, data_stage_1__5911_, data_stage_1__5910_, data_stage_1__5909_, data_stage_1__5908_, data_stage_1__5907_, data_stage_1__5906_, data_stage_1__5905_, data_stage_1__5904_, data_stage_1__5903_, data_stage_1__5902_, data_stage_1__5901_, data_stage_1__5900_, data_stage_1__5899_, data_stage_1__5898_, data_stage_1__5897_, data_stage_1__5896_, data_stage_1__5895_, data_stage_1__5894_, data_stage_1__5893_, data_stage_1__5892_, data_stage_1__5891_, data_stage_1__5890_, data_stage_1__5889_, data_stage_1__5888_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_24__swap_inst
  (
    .data_i(data_i[6399:6144]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__6399_, data_stage_1__6398_, data_stage_1__6397_, data_stage_1__6396_, data_stage_1__6395_, data_stage_1__6394_, data_stage_1__6393_, data_stage_1__6392_, data_stage_1__6391_, data_stage_1__6390_, data_stage_1__6389_, data_stage_1__6388_, data_stage_1__6387_, data_stage_1__6386_, data_stage_1__6385_, data_stage_1__6384_, data_stage_1__6383_, data_stage_1__6382_, data_stage_1__6381_, data_stage_1__6380_, data_stage_1__6379_, data_stage_1__6378_, data_stage_1__6377_, data_stage_1__6376_, data_stage_1__6375_, data_stage_1__6374_, data_stage_1__6373_, data_stage_1__6372_, data_stage_1__6371_, data_stage_1__6370_, data_stage_1__6369_, data_stage_1__6368_, data_stage_1__6367_, data_stage_1__6366_, data_stage_1__6365_, data_stage_1__6364_, data_stage_1__6363_, data_stage_1__6362_, data_stage_1__6361_, data_stage_1__6360_, data_stage_1__6359_, data_stage_1__6358_, data_stage_1__6357_, data_stage_1__6356_, data_stage_1__6355_, data_stage_1__6354_, data_stage_1__6353_, data_stage_1__6352_, data_stage_1__6351_, data_stage_1__6350_, data_stage_1__6349_, data_stage_1__6348_, data_stage_1__6347_, data_stage_1__6346_, data_stage_1__6345_, data_stage_1__6344_, data_stage_1__6343_, data_stage_1__6342_, data_stage_1__6341_, data_stage_1__6340_, data_stage_1__6339_, data_stage_1__6338_, data_stage_1__6337_, data_stage_1__6336_, data_stage_1__6335_, data_stage_1__6334_, data_stage_1__6333_, data_stage_1__6332_, data_stage_1__6331_, data_stage_1__6330_, data_stage_1__6329_, data_stage_1__6328_, data_stage_1__6327_, data_stage_1__6326_, data_stage_1__6325_, data_stage_1__6324_, data_stage_1__6323_, data_stage_1__6322_, data_stage_1__6321_, data_stage_1__6320_, data_stage_1__6319_, data_stage_1__6318_, data_stage_1__6317_, data_stage_1__6316_, data_stage_1__6315_, data_stage_1__6314_, data_stage_1__6313_, data_stage_1__6312_, data_stage_1__6311_, data_stage_1__6310_, data_stage_1__6309_, data_stage_1__6308_, data_stage_1__6307_, data_stage_1__6306_, data_stage_1__6305_, data_stage_1__6304_, data_stage_1__6303_, data_stage_1__6302_, data_stage_1__6301_, data_stage_1__6300_, data_stage_1__6299_, data_stage_1__6298_, data_stage_1__6297_, data_stage_1__6296_, data_stage_1__6295_, data_stage_1__6294_, data_stage_1__6293_, data_stage_1__6292_, data_stage_1__6291_, data_stage_1__6290_, data_stage_1__6289_, data_stage_1__6288_, data_stage_1__6287_, data_stage_1__6286_, data_stage_1__6285_, data_stage_1__6284_, data_stage_1__6283_, data_stage_1__6282_, data_stage_1__6281_, data_stage_1__6280_, data_stage_1__6279_, data_stage_1__6278_, data_stage_1__6277_, data_stage_1__6276_, data_stage_1__6275_, data_stage_1__6274_, data_stage_1__6273_, data_stage_1__6272_, data_stage_1__6271_, data_stage_1__6270_, data_stage_1__6269_, data_stage_1__6268_, data_stage_1__6267_, data_stage_1__6266_, data_stage_1__6265_, data_stage_1__6264_, data_stage_1__6263_, data_stage_1__6262_, data_stage_1__6261_, data_stage_1__6260_, data_stage_1__6259_, data_stage_1__6258_, data_stage_1__6257_, data_stage_1__6256_, data_stage_1__6255_, data_stage_1__6254_, data_stage_1__6253_, data_stage_1__6252_, data_stage_1__6251_, data_stage_1__6250_, data_stage_1__6249_, data_stage_1__6248_, data_stage_1__6247_, data_stage_1__6246_, data_stage_1__6245_, data_stage_1__6244_, data_stage_1__6243_, data_stage_1__6242_, data_stage_1__6241_, data_stage_1__6240_, data_stage_1__6239_, data_stage_1__6238_, data_stage_1__6237_, data_stage_1__6236_, data_stage_1__6235_, data_stage_1__6234_, data_stage_1__6233_, data_stage_1__6232_, data_stage_1__6231_, data_stage_1__6230_, data_stage_1__6229_, data_stage_1__6228_, data_stage_1__6227_, data_stage_1__6226_, data_stage_1__6225_, data_stage_1__6224_, data_stage_1__6223_, data_stage_1__6222_, data_stage_1__6221_, data_stage_1__6220_, data_stage_1__6219_, data_stage_1__6218_, data_stage_1__6217_, data_stage_1__6216_, data_stage_1__6215_, data_stage_1__6214_, data_stage_1__6213_, data_stage_1__6212_, data_stage_1__6211_, data_stage_1__6210_, data_stage_1__6209_, data_stage_1__6208_, data_stage_1__6207_, data_stage_1__6206_, data_stage_1__6205_, data_stage_1__6204_, data_stage_1__6203_, data_stage_1__6202_, data_stage_1__6201_, data_stage_1__6200_, data_stage_1__6199_, data_stage_1__6198_, data_stage_1__6197_, data_stage_1__6196_, data_stage_1__6195_, data_stage_1__6194_, data_stage_1__6193_, data_stage_1__6192_, data_stage_1__6191_, data_stage_1__6190_, data_stage_1__6189_, data_stage_1__6188_, data_stage_1__6187_, data_stage_1__6186_, data_stage_1__6185_, data_stage_1__6184_, data_stage_1__6183_, data_stage_1__6182_, data_stage_1__6181_, data_stage_1__6180_, data_stage_1__6179_, data_stage_1__6178_, data_stage_1__6177_, data_stage_1__6176_, data_stage_1__6175_, data_stage_1__6174_, data_stage_1__6173_, data_stage_1__6172_, data_stage_1__6171_, data_stage_1__6170_, data_stage_1__6169_, data_stage_1__6168_, data_stage_1__6167_, data_stage_1__6166_, data_stage_1__6165_, data_stage_1__6164_, data_stage_1__6163_, data_stage_1__6162_, data_stage_1__6161_, data_stage_1__6160_, data_stage_1__6159_, data_stage_1__6158_, data_stage_1__6157_, data_stage_1__6156_, data_stage_1__6155_, data_stage_1__6154_, data_stage_1__6153_, data_stage_1__6152_, data_stage_1__6151_, data_stage_1__6150_, data_stage_1__6149_, data_stage_1__6148_, data_stage_1__6147_, data_stage_1__6146_, data_stage_1__6145_, data_stage_1__6144_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_25__swap_inst
  (
    .data_i(data_i[6655:6400]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__6655_, data_stage_1__6654_, data_stage_1__6653_, data_stage_1__6652_, data_stage_1__6651_, data_stage_1__6650_, data_stage_1__6649_, data_stage_1__6648_, data_stage_1__6647_, data_stage_1__6646_, data_stage_1__6645_, data_stage_1__6644_, data_stage_1__6643_, data_stage_1__6642_, data_stage_1__6641_, data_stage_1__6640_, data_stage_1__6639_, data_stage_1__6638_, data_stage_1__6637_, data_stage_1__6636_, data_stage_1__6635_, data_stage_1__6634_, data_stage_1__6633_, data_stage_1__6632_, data_stage_1__6631_, data_stage_1__6630_, data_stage_1__6629_, data_stage_1__6628_, data_stage_1__6627_, data_stage_1__6626_, data_stage_1__6625_, data_stage_1__6624_, data_stage_1__6623_, data_stage_1__6622_, data_stage_1__6621_, data_stage_1__6620_, data_stage_1__6619_, data_stage_1__6618_, data_stage_1__6617_, data_stage_1__6616_, data_stage_1__6615_, data_stage_1__6614_, data_stage_1__6613_, data_stage_1__6612_, data_stage_1__6611_, data_stage_1__6610_, data_stage_1__6609_, data_stage_1__6608_, data_stage_1__6607_, data_stage_1__6606_, data_stage_1__6605_, data_stage_1__6604_, data_stage_1__6603_, data_stage_1__6602_, data_stage_1__6601_, data_stage_1__6600_, data_stage_1__6599_, data_stage_1__6598_, data_stage_1__6597_, data_stage_1__6596_, data_stage_1__6595_, data_stage_1__6594_, data_stage_1__6593_, data_stage_1__6592_, data_stage_1__6591_, data_stage_1__6590_, data_stage_1__6589_, data_stage_1__6588_, data_stage_1__6587_, data_stage_1__6586_, data_stage_1__6585_, data_stage_1__6584_, data_stage_1__6583_, data_stage_1__6582_, data_stage_1__6581_, data_stage_1__6580_, data_stage_1__6579_, data_stage_1__6578_, data_stage_1__6577_, data_stage_1__6576_, data_stage_1__6575_, data_stage_1__6574_, data_stage_1__6573_, data_stage_1__6572_, data_stage_1__6571_, data_stage_1__6570_, data_stage_1__6569_, data_stage_1__6568_, data_stage_1__6567_, data_stage_1__6566_, data_stage_1__6565_, data_stage_1__6564_, data_stage_1__6563_, data_stage_1__6562_, data_stage_1__6561_, data_stage_1__6560_, data_stage_1__6559_, data_stage_1__6558_, data_stage_1__6557_, data_stage_1__6556_, data_stage_1__6555_, data_stage_1__6554_, data_stage_1__6553_, data_stage_1__6552_, data_stage_1__6551_, data_stage_1__6550_, data_stage_1__6549_, data_stage_1__6548_, data_stage_1__6547_, data_stage_1__6546_, data_stage_1__6545_, data_stage_1__6544_, data_stage_1__6543_, data_stage_1__6542_, data_stage_1__6541_, data_stage_1__6540_, data_stage_1__6539_, data_stage_1__6538_, data_stage_1__6537_, data_stage_1__6536_, data_stage_1__6535_, data_stage_1__6534_, data_stage_1__6533_, data_stage_1__6532_, data_stage_1__6531_, data_stage_1__6530_, data_stage_1__6529_, data_stage_1__6528_, data_stage_1__6527_, data_stage_1__6526_, data_stage_1__6525_, data_stage_1__6524_, data_stage_1__6523_, data_stage_1__6522_, data_stage_1__6521_, data_stage_1__6520_, data_stage_1__6519_, data_stage_1__6518_, data_stage_1__6517_, data_stage_1__6516_, data_stage_1__6515_, data_stage_1__6514_, data_stage_1__6513_, data_stage_1__6512_, data_stage_1__6511_, data_stage_1__6510_, data_stage_1__6509_, data_stage_1__6508_, data_stage_1__6507_, data_stage_1__6506_, data_stage_1__6505_, data_stage_1__6504_, data_stage_1__6503_, data_stage_1__6502_, data_stage_1__6501_, data_stage_1__6500_, data_stage_1__6499_, data_stage_1__6498_, data_stage_1__6497_, data_stage_1__6496_, data_stage_1__6495_, data_stage_1__6494_, data_stage_1__6493_, data_stage_1__6492_, data_stage_1__6491_, data_stage_1__6490_, data_stage_1__6489_, data_stage_1__6488_, data_stage_1__6487_, data_stage_1__6486_, data_stage_1__6485_, data_stage_1__6484_, data_stage_1__6483_, data_stage_1__6482_, data_stage_1__6481_, data_stage_1__6480_, data_stage_1__6479_, data_stage_1__6478_, data_stage_1__6477_, data_stage_1__6476_, data_stage_1__6475_, data_stage_1__6474_, data_stage_1__6473_, data_stage_1__6472_, data_stage_1__6471_, data_stage_1__6470_, data_stage_1__6469_, data_stage_1__6468_, data_stage_1__6467_, data_stage_1__6466_, data_stage_1__6465_, data_stage_1__6464_, data_stage_1__6463_, data_stage_1__6462_, data_stage_1__6461_, data_stage_1__6460_, data_stage_1__6459_, data_stage_1__6458_, data_stage_1__6457_, data_stage_1__6456_, data_stage_1__6455_, data_stage_1__6454_, data_stage_1__6453_, data_stage_1__6452_, data_stage_1__6451_, data_stage_1__6450_, data_stage_1__6449_, data_stage_1__6448_, data_stage_1__6447_, data_stage_1__6446_, data_stage_1__6445_, data_stage_1__6444_, data_stage_1__6443_, data_stage_1__6442_, data_stage_1__6441_, data_stage_1__6440_, data_stage_1__6439_, data_stage_1__6438_, data_stage_1__6437_, data_stage_1__6436_, data_stage_1__6435_, data_stage_1__6434_, data_stage_1__6433_, data_stage_1__6432_, data_stage_1__6431_, data_stage_1__6430_, data_stage_1__6429_, data_stage_1__6428_, data_stage_1__6427_, data_stage_1__6426_, data_stage_1__6425_, data_stage_1__6424_, data_stage_1__6423_, data_stage_1__6422_, data_stage_1__6421_, data_stage_1__6420_, data_stage_1__6419_, data_stage_1__6418_, data_stage_1__6417_, data_stage_1__6416_, data_stage_1__6415_, data_stage_1__6414_, data_stage_1__6413_, data_stage_1__6412_, data_stage_1__6411_, data_stage_1__6410_, data_stage_1__6409_, data_stage_1__6408_, data_stage_1__6407_, data_stage_1__6406_, data_stage_1__6405_, data_stage_1__6404_, data_stage_1__6403_, data_stage_1__6402_, data_stage_1__6401_, data_stage_1__6400_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_26__swap_inst
  (
    .data_i(data_i[6911:6656]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__6911_, data_stage_1__6910_, data_stage_1__6909_, data_stage_1__6908_, data_stage_1__6907_, data_stage_1__6906_, data_stage_1__6905_, data_stage_1__6904_, data_stage_1__6903_, data_stage_1__6902_, data_stage_1__6901_, data_stage_1__6900_, data_stage_1__6899_, data_stage_1__6898_, data_stage_1__6897_, data_stage_1__6896_, data_stage_1__6895_, data_stage_1__6894_, data_stage_1__6893_, data_stage_1__6892_, data_stage_1__6891_, data_stage_1__6890_, data_stage_1__6889_, data_stage_1__6888_, data_stage_1__6887_, data_stage_1__6886_, data_stage_1__6885_, data_stage_1__6884_, data_stage_1__6883_, data_stage_1__6882_, data_stage_1__6881_, data_stage_1__6880_, data_stage_1__6879_, data_stage_1__6878_, data_stage_1__6877_, data_stage_1__6876_, data_stage_1__6875_, data_stage_1__6874_, data_stage_1__6873_, data_stage_1__6872_, data_stage_1__6871_, data_stage_1__6870_, data_stage_1__6869_, data_stage_1__6868_, data_stage_1__6867_, data_stage_1__6866_, data_stage_1__6865_, data_stage_1__6864_, data_stage_1__6863_, data_stage_1__6862_, data_stage_1__6861_, data_stage_1__6860_, data_stage_1__6859_, data_stage_1__6858_, data_stage_1__6857_, data_stage_1__6856_, data_stage_1__6855_, data_stage_1__6854_, data_stage_1__6853_, data_stage_1__6852_, data_stage_1__6851_, data_stage_1__6850_, data_stage_1__6849_, data_stage_1__6848_, data_stage_1__6847_, data_stage_1__6846_, data_stage_1__6845_, data_stage_1__6844_, data_stage_1__6843_, data_stage_1__6842_, data_stage_1__6841_, data_stage_1__6840_, data_stage_1__6839_, data_stage_1__6838_, data_stage_1__6837_, data_stage_1__6836_, data_stage_1__6835_, data_stage_1__6834_, data_stage_1__6833_, data_stage_1__6832_, data_stage_1__6831_, data_stage_1__6830_, data_stage_1__6829_, data_stage_1__6828_, data_stage_1__6827_, data_stage_1__6826_, data_stage_1__6825_, data_stage_1__6824_, data_stage_1__6823_, data_stage_1__6822_, data_stage_1__6821_, data_stage_1__6820_, data_stage_1__6819_, data_stage_1__6818_, data_stage_1__6817_, data_stage_1__6816_, data_stage_1__6815_, data_stage_1__6814_, data_stage_1__6813_, data_stage_1__6812_, data_stage_1__6811_, data_stage_1__6810_, data_stage_1__6809_, data_stage_1__6808_, data_stage_1__6807_, data_stage_1__6806_, data_stage_1__6805_, data_stage_1__6804_, data_stage_1__6803_, data_stage_1__6802_, data_stage_1__6801_, data_stage_1__6800_, data_stage_1__6799_, data_stage_1__6798_, data_stage_1__6797_, data_stage_1__6796_, data_stage_1__6795_, data_stage_1__6794_, data_stage_1__6793_, data_stage_1__6792_, data_stage_1__6791_, data_stage_1__6790_, data_stage_1__6789_, data_stage_1__6788_, data_stage_1__6787_, data_stage_1__6786_, data_stage_1__6785_, data_stage_1__6784_, data_stage_1__6783_, data_stage_1__6782_, data_stage_1__6781_, data_stage_1__6780_, data_stage_1__6779_, data_stage_1__6778_, data_stage_1__6777_, data_stage_1__6776_, data_stage_1__6775_, data_stage_1__6774_, data_stage_1__6773_, data_stage_1__6772_, data_stage_1__6771_, data_stage_1__6770_, data_stage_1__6769_, data_stage_1__6768_, data_stage_1__6767_, data_stage_1__6766_, data_stage_1__6765_, data_stage_1__6764_, data_stage_1__6763_, data_stage_1__6762_, data_stage_1__6761_, data_stage_1__6760_, data_stage_1__6759_, data_stage_1__6758_, data_stage_1__6757_, data_stage_1__6756_, data_stage_1__6755_, data_stage_1__6754_, data_stage_1__6753_, data_stage_1__6752_, data_stage_1__6751_, data_stage_1__6750_, data_stage_1__6749_, data_stage_1__6748_, data_stage_1__6747_, data_stage_1__6746_, data_stage_1__6745_, data_stage_1__6744_, data_stage_1__6743_, data_stage_1__6742_, data_stage_1__6741_, data_stage_1__6740_, data_stage_1__6739_, data_stage_1__6738_, data_stage_1__6737_, data_stage_1__6736_, data_stage_1__6735_, data_stage_1__6734_, data_stage_1__6733_, data_stage_1__6732_, data_stage_1__6731_, data_stage_1__6730_, data_stage_1__6729_, data_stage_1__6728_, data_stage_1__6727_, data_stage_1__6726_, data_stage_1__6725_, data_stage_1__6724_, data_stage_1__6723_, data_stage_1__6722_, data_stage_1__6721_, data_stage_1__6720_, data_stage_1__6719_, data_stage_1__6718_, data_stage_1__6717_, data_stage_1__6716_, data_stage_1__6715_, data_stage_1__6714_, data_stage_1__6713_, data_stage_1__6712_, data_stage_1__6711_, data_stage_1__6710_, data_stage_1__6709_, data_stage_1__6708_, data_stage_1__6707_, data_stage_1__6706_, data_stage_1__6705_, data_stage_1__6704_, data_stage_1__6703_, data_stage_1__6702_, data_stage_1__6701_, data_stage_1__6700_, data_stage_1__6699_, data_stage_1__6698_, data_stage_1__6697_, data_stage_1__6696_, data_stage_1__6695_, data_stage_1__6694_, data_stage_1__6693_, data_stage_1__6692_, data_stage_1__6691_, data_stage_1__6690_, data_stage_1__6689_, data_stage_1__6688_, data_stage_1__6687_, data_stage_1__6686_, data_stage_1__6685_, data_stage_1__6684_, data_stage_1__6683_, data_stage_1__6682_, data_stage_1__6681_, data_stage_1__6680_, data_stage_1__6679_, data_stage_1__6678_, data_stage_1__6677_, data_stage_1__6676_, data_stage_1__6675_, data_stage_1__6674_, data_stage_1__6673_, data_stage_1__6672_, data_stage_1__6671_, data_stage_1__6670_, data_stage_1__6669_, data_stage_1__6668_, data_stage_1__6667_, data_stage_1__6666_, data_stage_1__6665_, data_stage_1__6664_, data_stage_1__6663_, data_stage_1__6662_, data_stage_1__6661_, data_stage_1__6660_, data_stage_1__6659_, data_stage_1__6658_, data_stage_1__6657_, data_stage_1__6656_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_27__swap_inst
  (
    .data_i(data_i[7167:6912]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__7167_, data_stage_1__7166_, data_stage_1__7165_, data_stage_1__7164_, data_stage_1__7163_, data_stage_1__7162_, data_stage_1__7161_, data_stage_1__7160_, data_stage_1__7159_, data_stage_1__7158_, data_stage_1__7157_, data_stage_1__7156_, data_stage_1__7155_, data_stage_1__7154_, data_stage_1__7153_, data_stage_1__7152_, data_stage_1__7151_, data_stage_1__7150_, data_stage_1__7149_, data_stage_1__7148_, data_stage_1__7147_, data_stage_1__7146_, data_stage_1__7145_, data_stage_1__7144_, data_stage_1__7143_, data_stage_1__7142_, data_stage_1__7141_, data_stage_1__7140_, data_stage_1__7139_, data_stage_1__7138_, data_stage_1__7137_, data_stage_1__7136_, data_stage_1__7135_, data_stage_1__7134_, data_stage_1__7133_, data_stage_1__7132_, data_stage_1__7131_, data_stage_1__7130_, data_stage_1__7129_, data_stage_1__7128_, data_stage_1__7127_, data_stage_1__7126_, data_stage_1__7125_, data_stage_1__7124_, data_stage_1__7123_, data_stage_1__7122_, data_stage_1__7121_, data_stage_1__7120_, data_stage_1__7119_, data_stage_1__7118_, data_stage_1__7117_, data_stage_1__7116_, data_stage_1__7115_, data_stage_1__7114_, data_stage_1__7113_, data_stage_1__7112_, data_stage_1__7111_, data_stage_1__7110_, data_stage_1__7109_, data_stage_1__7108_, data_stage_1__7107_, data_stage_1__7106_, data_stage_1__7105_, data_stage_1__7104_, data_stage_1__7103_, data_stage_1__7102_, data_stage_1__7101_, data_stage_1__7100_, data_stage_1__7099_, data_stage_1__7098_, data_stage_1__7097_, data_stage_1__7096_, data_stage_1__7095_, data_stage_1__7094_, data_stage_1__7093_, data_stage_1__7092_, data_stage_1__7091_, data_stage_1__7090_, data_stage_1__7089_, data_stage_1__7088_, data_stage_1__7087_, data_stage_1__7086_, data_stage_1__7085_, data_stage_1__7084_, data_stage_1__7083_, data_stage_1__7082_, data_stage_1__7081_, data_stage_1__7080_, data_stage_1__7079_, data_stage_1__7078_, data_stage_1__7077_, data_stage_1__7076_, data_stage_1__7075_, data_stage_1__7074_, data_stage_1__7073_, data_stage_1__7072_, data_stage_1__7071_, data_stage_1__7070_, data_stage_1__7069_, data_stage_1__7068_, data_stage_1__7067_, data_stage_1__7066_, data_stage_1__7065_, data_stage_1__7064_, data_stage_1__7063_, data_stage_1__7062_, data_stage_1__7061_, data_stage_1__7060_, data_stage_1__7059_, data_stage_1__7058_, data_stage_1__7057_, data_stage_1__7056_, data_stage_1__7055_, data_stage_1__7054_, data_stage_1__7053_, data_stage_1__7052_, data_stage_1__7051_, data_stage_1__7050_, data_stage_1__7049_, data_stage_1__7048_, data_stage_1__7047_, data_stage_1__7046_, data_stage_1__7045_, data_stage_1__7044_, data_stage_1__7043_, data_stage_1__7042_, data_stage_1__7041_, data_stage_1__7040_, data_stage_1__7039_, data_stage_1__7038_, data_stage_1__7037_, data_stage_1__7036_, data_stage_1__7035_, data_stage_1__7034_, data_stage_1__7033_, data_stage_1__7032_, data_stage_1__7031_, data_stage_1__7030_, data_stage_1__7029_, data_stage_1__7028_, data_stage_1__7027_, data_stage_1__7026_, data_stage_1__7025_, data_stage_1__7024_, data_stage_1__7023_, data_stage_1__7022_, data_stage_1__7021_, data_stage_1__7020_, data_stage_1__7019_, data_stage_1__7018_, data_stage_1__7017_, data_stage_1__7016_, data_stage_1__7015_, data_stage_1__7014_, data_stage_1__7013_, data_stage_1__7012_, data_stage_1__7011_, data_stage_1__7010_, data_stage_1__7009_, data_stage_1__7008_, data_stage_1__7007_, data_stage_1__7006_, data_stage_1__7005_, data_stage_1__7004_, data_stage_1__7003_, data_stage_1__7002_, data_stage_1__7001_, data_stage_1__7000_, data_stage_1__6999_, data_stage_1__6998_, data_stage_1__6997_, data_stage_1__6996_, data_stage_1__6995_, data_stage_1__6994_, data_stage_1__6993_, data_stage_1__6992_, data_stage_1__6991_, data_stage_1__6990_, data_stage_1__6989_, data_stage_1__6988_, data_stage_1__6987_, data_stage_1__6986_, data_stage_1__6985_, data_stage_1__6984_, data_stage_1__6983_, data_stage_1__6982_, data_stage_1__6981_, data_stage_1__6980_, data_stage_1__6979_, data_stage_1__6978_, data_stage_1__6977_, data_stage_1__6976_, data_stage_1__6975_, data_stage_1__6974_, data_stage_1__6973_, data_stage_1__6972_, data_stage_1__6971_, data_stage_1__6970_, data_stage_1__6969_, data_stage_1__6968_, data_stage_1__6967_, data_stage_1__6966_, data_stage_1__6965_, data_stage_1__6964_, data_stage_1__6963_, data_stage_1__6962_, data_stage_1__6961_, data_stage_1__6960_, data_stage_1__6959_, data_stage_1__6958_, data_stage_1__6957_, data_stage_1__6956_, data_stage_1__6955_, data_stage_1__6954_, data_stage_1__6953_, data_stage_1__6952_, data_stage_1__6951_, data_stage_1__6950_, data_stage_1__6949_, data_stage_1__6948_, data_stage_1__6947_, data_stage_1__6946_, data_stage_1__6945_, data_stage_1__6944_, data_stage_1__6943_, data_stage_1__6942_, data_stage_1__6941_, data_stage_1__6940_, data_stage_1__6939_, data_stage_1__6938_, data_stage_1__6937_, data_stage_1__6936_, data_stage_1__6935_, data_stage_1__6934_, data_stage_1__6933_, data_stage_1__6932_, data_stage_1__6931_, data_stage_1__6930_, data_stage_1__6929_, data_stage_1__6928_, data_stage_1__6927_, data_stage_1__6926_, data_stage_1__6925_, data_stage_1__6924_, data_stage_1__6923_, data_stage_1__6922_, data_stage_1__6921_, data_stage_1__6920_, data_stage_1__6919_, data_stage_1__6918_, data_stage_1__6917_, data_stage_1__6916_, data_stage_1__6915_, data_stage_1__6914_, data_stage_1__6913_, data_stage_1__6912_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_28__swap_inst
  (
    .data_i(data_i[7423:7168]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__7423_, data_stage_1__7422_, data_stage_1__7421_, data_stage_1__7420_, data_stage_1__7419_, data_stage_1__7418_, data_stage_1__7417_, data_stage_1__7416_, data_stage_1__7415_, data_stage_1__7414_, data_stage_1__7413_, data_stage_1__7412_, data_stage_1__7411_, data_stage_1__7410_, data_stage_1__7409_, data_stage_1__7408_, data_stage_1__7407_, data_stage_1__7406_, data_stage_1__7405_, data_stage_1__7404_, data_stage_1__7403_, data_stage_1__7402_, data_stage_1__7401_, data_stage_1__7400_, data_stage_1__7399_, data_stage_1__7398_, data_stage_1__7397_, data_stage_1__7396_, data_stage_1__7395_, data_stage_1__7394_, data_stage_1__7393_, data_stage_1__7392_, data_stage_1__7391_, data_stage_1__7390_, data_stage_1__7389_, data_stage_1__7388_, data_stage_1__7387_, data_stage_1__7386_, data_stage_1__7385_, data_stage_1__7384_, data_stage_1__7383_, data_stage_1__7382_, data_stage_1__7381_, data_stage_1__7380_, data_stage_1__7379_, data_stage_1__7378_, data_stage_1__7377_, data_stage_1__7376_, data_stage_1__7375_, data_stage_1__7374_, data_stage_1__7373_, data_stage_1__7372_, data_stage_1__7371_, data_stage_1__7370_, data_stage_1__7369_, data_stage_1__7368_, data_stage_1__7367_, data_stage_1__7366_, data_stage_1__7365_, data_stage_1__7364_, data_stage_1__7363_, data_stage_1__7362_, data_stage_1__7361_, data_stage_1__7360_, data_stage_1__7359_, data_stage_1__7358_, data_stage_1__7357_, data_stage_1__7356_, data_stage_1__7355_, data_stage_1__7354_, data_stage_1__7353_, data_stage_1__7352_, data_stage_1__7351_, data_stage_1__7350_, data_stage_1__7349_, data_stage_1__7348_, data_stage_1__7347_, data_stage_1__7346_, data_stage_1__7345_, data_stage_1__7344_, data_stage_1__7343_, data_stage_1__7342_, data_stage_1__7341_, data_stage_1__7340_, data_stage_1__7339_, data_stage_1__7338_, data_stage_1__7337_, data_stage_1__7336_, data_stage_1__7335_, data_stage_1__7334_, data_stage_1__7333_, data_stage_1__7332_, data_stage_1__7331_, data_stage_1__7330_, data_stage_1__7329_, data_stage_1__7328_, data_stage_1__7327_, data_stage_1__7326_, data_stage_1__7325_, data_stage_1__7324_, data_stage_1__7323_, data_stage_1__7322_, data_stage_1__7321_, data_stage_1__7320_, data_stage_1__7319_, data_stage_1__7318_, data_stage_1__7317_, data_stage_1__7316_, data_stage_1__7315_, data_stage_1__7314_, data_stage_1__7313_, data_stage_1__7312_, data_stage_1__7311_, data_stage_1__7310_, data_stage_1__7309_, data_stage_1__7308_, data_stage_1__7307_, data_stage_1__7306_, data_stage_1__7305_, data_stage_1__7304_, data_stage_1__7303_, data_stage_1__7302_, data_stage_1__7301_, data_stage_1__7300_, data_stage_1__7299_, data_stage_1__7298_, data_stage_1__7297_, data_stage_1__7296_, data_stage_1__7295_, data_stage_1__7294_, data_stage_1__7293_, data_stage_1__7292_, data_stage_1__7291_, data_stage_1__7290_, data_stage_1__7289_, data_stage_1__7288_, data_stage_1__7287_, data_stage_1__7286_, data_stage_1__7285_, data_stage_1__7284_, data_stage_1__7283_, data_stage_1__7282_, data_stage_1__7281_, data_stage_1__7280_, data_stage_1__7279_, data_stage_1__7278_, data_stage_1__7277_, data_stage_1__7276_, data_stage_1__7275_, data_stage_1__7274_, data_stage_1__7273_, data_stage_1__7272_, data_stage_1__7271_, data_stage_1__7270_, data_stage_1__7269_, data_stage_1__7268_, data_stage_1__7267_, data_stage_1__7266_, data_stage_1__7265_, data_stage_1__7264_, data_stage_1__7263_, data_stage_1__7262_, data_stage_1__7261_, data_stage_1__7260_, data_stage_1__7259_, data_stage_1__7258_, data_stage_1__7257_, data_stage_1__7256_, data_stage_1__7255_, data_stage_1__7254_, data_stage_1__7253_, data_stage_1__7252_, data_stage_1__7251_, data_stage_1__7250_, data_stage_1__7249_, data_stage_1__7248_, data_stage_1__7247_, data_stage_1__7246_, data_stage_1__7245_, data_stage_1__7244_, data_stage_1__7243_, data_stage_1__7242_, data_stage_1__7241_, data_stage_1__7240_, data_stage_1__7239_, data_stage_1__7238_, data_stage_1__7237_, data_stage_1__7236_, data_stage_1__7235_, data_stage_1__7234_, data_stage_1__7233_, data_stage_1__7232_, data_stage_1__7231_, data_stage_1__7230_, data_stage_1__7229_, data_stage_1__7228_, data_stage_1__7227_, data_stage_1__7226_, data_stage_1__7225_, data_stage_1__7224_, data_stage_1__7223_, data_stage_1__7222_, data_stage_1__7221_, data_stage_1__7220_, data_stage_1__7219_, data_stage_1__7218_, data_stage_1__7217_, data_stage_1__7216_, data_stage_1__7215_, data_stage_1__7214_, data_stage_1__7213_, data_stage_1__7212_, data_stage_1__7211_, data_stage_1__7210_, data_stage_1__7209_, data_stage_1__7208_, data_stage_1__7207_, data_stage_1__7206_, data_stage_1__7205_, data_stage_1__7204_, data_stage_1__7203_, data_stage_1__7202_, data_stage_1__7201_, data_stage_1__7200_, data_stage_1__7199_, data_stage_1__7198_, data_stage_1__7197_, data_stage_1__7196_, data_stage_1__7195_, data_stage_1__7194_, data_stage_1__7193_, data_stage_1__7192_, data_stage_1__7191_, data_stage_1__7190_, data_stage_1__7189_, data_stage_1__7188_, data_stage_1__7187_, data_stage_1__7186_, data_stage_1__7185_, data_stage_1__7184_, data_stage_1__7183_, data_stage_1__7182_, data_stage_1__7181_, data_stage_1__7180_, data_stage_1__7179_, data_stage_1__7178_, data_stage_1__7177_, data_stage_1__7176_, data_stage_1__7175_, data_stage_1__7174_, data_stage_1__7173_, data_stage_1__7172_, data_stage_1__7171_, data_stage_1__7170_, data_stage_1__7169_, data_stage_1__7168_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_29__swap_inst
  (
    .data_i(data_i[7679:7424]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__7679_, data_stage_1__7678_, data_stage_1__7677_, data_stage_1__7676_, data_stage_1__7675_, data_stage_1__7674_, data_stage_1__7673_, data_stage_1__7672_, data_stage_1__7671_, data_stage_1__7670_, data_stage_1__7669_, data_stage_1__7668_, data_stage_1__7667_, data_stage_1__7666_, data_stage_1__7665_, data_stage_1__7664_, data_stage_1__7663_, data_stage_1__7662_, data_stage_1__7661_, data_stage_1__7660_, data_stage_1__7659_, data_stage_1__7658_, data_stage_1__7657_, data_stage_1__7656_, data_stage_1__7655_, data_stage_1__7654_, data_stage_1__7653_, data_stage_1__7652_, data_stage_1__7651_, data_stage_1__7650_, data_stage_1__7649_, data_stage_1__7648_, data_stage_1__7647_, data_stage_1__7646_, data_stage_1__7645_, data_stage_1__7644_, data_stage_1__7643_, data_stage_1__7642_, data_stage_1__7641_, data_stage_1__7640_, data_stage_1__7639_, data_stage_1__7638_, data_stage_1__7637_, data_stage_1__7636_, data_stage_1__7635_, data_stage_1__7634_, data_stage_1__7633_, data_stage_1__7632_, data_stage_1__7631_, data_stage_1__7630_, data_stage_1__7629_, data_stage_1__7628_, data_stage_1__7627_, data_stage_1__7626_, data_stage_1__7625_, data_stage_1__7624_, data_stage_1__7623_, data_stage_1__7622_, data_stage_1__7621_, data_stage_1__7620_, data_stage_1__7619_, data_stage_1__7618_, data_stage_1__7617_, data_stage_1__7616_, data_stage_1__7615_, data_stage_1__7614_, data_stage_1__7613_, data_stage_1__7612_, data_stage_1__7611_, data_stage_1__7610_, data_stage_1__7609_, data_stage_1__7608_, data_stage_1__7607_, data_stage_1__7606_, data_stage_1__7605_, data_stage_1__7604_, data_stage_1__7603_, data_stage_1__7602_, data_stage_1__7601_, data_stage_1__7600_, data_stage_1__7599_, data_stage_1__7598_, data_stage_1__7597_, data_stage_1__7596_, data_stage_1__7595_, data_stage_1__7594_, data_stage_1__7593_, data_stage_1__7592_, data_stage_1__7591_, data_stage_1__7590_, data_stage_1__7589_, data_stage_1__7588_, data_stage_1__7587_, data_stage_1__7586_, data_stage_1__7585_, data_stage_1__7584_, data_stage_1__7583_, data_stage_1__7582_, data_stage_1__7581_, data_stage_1__7580_, data_stage_1__7579_, data_stage_1__7578_, data_stage_1__7577_, data_stage_1__7576_, data_stage_1__7575_, data_stage_1__7574_, data_stage_1__7573_, data_stage_1__7572_, data_stage_1__7571_, data_stage_1__7570_, data_stage_1__7569_, data_stage_1__7568_, data_stage_1__7567_, data_stage_1__7566_, data_stage_1__7565_, data_stage_1__7564_, data_stage_1__7563_, data_stage_1__7562_, data_stage_1__7561_, data_stage_1__7560_, data_stage_1__7559_, data_stage_1__7558_, data_stage_1__7557_, data_stage_1__7556_, data_stage_1__7555_, data_stage_1__7554_, data_stage_1__7553_, data_stage_1__7552_, data_stage_1__7551_, data_stage_1__7550_, data_stage_1__7549_, data_stage_1__7548_, data_stage_1__7547_, data_stage_1__7546_, data_stage_1__7545_, data_stage_1__7544_, data_stage_1__7543_, data_stage_1__7542_, data_stage_1__7541_, data_stage_1__7540_, data_stage_1__7539_, data_stage_1__7538_, data_stage_1__7537_, data_stage_1__7536_, data_stage_1__7535_, data_stage_1__7534_, data_stage_1__7533_, data_stage_1__7532_, data_stage_1__7531_, data_stage_1__7530_, data_stage_1__7529_, data_stage_1__7528_, data_stage_1__7527_, data_stage_1__7526_, data_stage_1__7525_, data_stage_1__7524_, data_stage_1__7523_, data_stage_1__7522_, data_stage_1__7521_, data_stage_1__7520_, data_stage_1__7519_, data_stage_1__7518_, data_stage_1__7517_, data_stage_1__7516_, data_stage_1__7515_, data_stage_1__7514_, data_stage_1__7513_, data_stage_1__7512_, data_stage_1__7511_, data_stage_1__7510_, data_stage_1__7509_, data_stage_1__7508_, data_stage_1__7507_, data_stage_1__7506_, data_stage_1__7505_, data_stage_1__7504_, data_stage_1__7503_, data_stage_1__7502_, data_stage_1__7501_, data_stage_1__7500_, data_stage_1__7499_, data_stage_1__7498_, data_stage_1__7497_, data_stage_1__7496_, data_stage_1__7495_, data_stage_1__7494_, data_stage_1__7493_, data_stage_1__7492_, data_stage_1__7491_, data_stage_1__7490_, data_stage_1__7489_, data_stage_1__7488_, data_stage_1__7487_, data_stage_1__7486_, data_stage_1__7485_, data_stage_1__7484_, data_stage_1__7483_, data_stage_1__7482_, data_stage_1__7481_, data_stage_1__7480_, data_stage_1__7479_, data_stage_1__7478_, data_stage_1__7477_, data_stage_1__7476_, data_stage_1__7475_, data_stage_1__7474_, data_stage_1__7473_, data_stage_1__7472_, data_stage_1__7471_, data_stage_1__7470_, data_stage_1__7469_, data_stage_1__7468_, data_stage_1__7467_, data_stage_1__7466_, data_stage_1__7465_, data_stage_1__7464_, data_stage_1__7463_, data_stage_1__7462_, data_stage_1__7461_, data_stage_1__7460_, data_stage_1__7459_, data_stage_1__7458_, data_stage_1__7457_, data_stage_1__7456_, data_stage_1__7455_, data_stage_1__7454_, data_stage_1__7453_, data_stage_1__7452_, data_stage_1__7451_, data_stage_1__7450_, data_stage_1__7449_, data_stage_1__7448_, data_stage_1__7447_, data_stage_1__7446_, data_stage_1__7445_, data_stage_1__7444_, data_stage_1__7443_, data_stage_1__7442_, data_stage_1__7441_, data_stage_1__7440_, data_stage_1__7439_, data_stage_1__7438_, data_stage_1__7437_, data_stage_1__7436_, data_stage_1__7435_, data_stage_1__7434_, data_stage_1__7433_, data_stage_1__7432_, data_stage_1__7431_, data_stage_1__7430_, data_stage_1__7429_, data_stage_1__7428_, data_stage_1__7427_, data_stage_1__7426_, data_stage_1__7425_, data_stage_1__7424_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_30__swap_inst
  (
    .data_i(data_i[7935:7680]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__7935_, data_stage_1__7934_, data_stage_1__7933_, data_stage_1__7932_, data_stage_1__7931_, data_stage_1__7930_, data_stage_1__7929_, data_stage_1__7928_, data_stage_1__7927_, data_stage_1__7926_, data_stage_1__7925_, data_stage_1__7924_, data_stage_1__7923_, data_stage_1__7922_, data_stage_1__7921_, data_stage_1__7920_, data_stage_1__7919_, data_stage_1__7918_, data_stage_1__7917_, data_stage_1__7916_, data_stage_1__7915_, data_stage_1__7914_, data_stage_1__7913_, data_stage_1__7912_, data_stage_1__7911_, data_stage_1__7910_, data_stage_1__7909_, data_stage_1__7908_, data_stage_1__7907_, data_stage_1__7906_, data_stage_1__7905_, data_stage_1__7904_, data_stage_1__7903_, data_stage_1__7902_, data_stage_1__7901_, data_stage_1__7900_, data_stage_1__7899_, data_stage_1__7898_, data_stage_1__7897_, data_stage_1__7896_, data_stage_1__7895_, data_stage_1__7894_, data_stage_1__7893_, data_stage_1__7892_, data_stage_1__7891_, data_stage_1__7890_, data_stage_1__7889_, data_stage_1__7888_, data_stage_1__7887_, data_stage_1__7886_, data_stage_1__7885_, data_stage_1__7884_, data_stage_1__7883_, data_stage_1__7882_, data_stage_1__7881_, data_stage_1__7880_, data_stage_1__7879_, data_stage_1__7878_, data_stage_1__7877_, data_stage_1__7876_, data_stage_1__7875_, data_stage_1__7874_, data_stage_1__7873_, data_stage_1__7872_, data_stage_1__7871_, data_stage_1__7870_, data_stage_1__7869_, data_stage_1__7868_, data_stage_1__7867_, data_stage_1__7866_, data_stage_1__7865_, data_stage_1__7864_, data_stage_1__7863_, data_stage_1__7862_, data_stage_1__7861_, data_stage_1__7860_, data_stage_1__7859_, data_stage_1__7858_, data_stage_1__7857_, data_stage_1__7856_, data_stage_1__7855_, data_stage_1__7854_, data_stage_1__7853_, data_stage_1__7852_, data_stage_1__7851_, data_stage_1__7850_, data_stage_1__7849_, data_stage_1__7848_, data_stage_1__7847_, data_stage_1__7846_, data_stage_1__7845_, data_stage_1__7844_, data_stage_1__7843_, data_stage_1__7842_, data_stage_1__7841_, data_stage_1__7840_, data_stage_1__7839_, data_stage_1__7838_, data_stage_1__7837_, data_stage_1__7836_, data_stage_1__7835_, data_stage_1__7834_, data_stage_1__7833_, data_stage_1__7832_, data_stage_1__7831_, data_stage_1__7830_, data_stage_1__7829_, data_stage_1__7828_, data_stage_1__7827_, data_stage_1__7826_, data_stage_1__7825_, data_stage_1__7824_, data_stage_1__7823_, data_stage_1__7822_, data_stage_1__7821_, data_stage_1__7820_, data_stage_1__7819_, data_stage_1__7818_, data_stage_1__7817_, data_stage_1__7816_, data_stage_1__7815_, data_stage_1__7814_, data_stage_1__7813_, data_stage_1__7812_, data_stage_1__7811_, data_stage_1__7810_, data_stage_1__7809_, data_stage_1__7808_, data_stage_1__7807_, data_stage_1__7806_, data_stage_1__7805_, data_stage_1__7804_, data_stage_1__7803_, data_stage_1__7802_, data_stage_1__7801_, data_stage_1__7800_, data_stage_1__7799_, data_stage_1__7798_, data_stage_1__7797_, data_stage_1__7796_, data_stage_1__7795_, data_stage_1__7794_, data_stage_1__7793_, data_stage_1__7792_, data_stage_1__7791_, data_stage_1__7790_, data_stage_1__7789_, data_stage_1__7788_, data_stage_1__7787_, data_stage_1__7786_, data_stage_1__7785_, data_stage_1__7784_, data_stage_1__7783_, data_stage_1__7782_, data_stage_1__7781_, data_stage_1__7780_, data_stage_1__7779_, data_stage_1__7778_, data_stage_1__7777_, data_stage_1__7776_, data_stage_1__7775_, data_stage_1__7774_, data_stage_1__7773_, data_stage_1__7772_, data_stage_1__7771_, data_stage_1__7770_, data_stage_1__7769_, data_stage_1__7768_, data_stage_1__7767_, data_stage_1__7766_, data_stage_1__7765_, data_stage_1__7764_, data_stage_1__7763_, data_stage_1__7762_, data_stage_1__7761_, data_stage_1__7760_, data_stage_1__7759_, data_stage_1__7758_, data_stage_1__7757_, data_stage_1__7756_, data_stage_1__7755_, data_stage_1__7754_, data_stage_1__7753_, data_stage_1__7752_, data_stage_1__7751_, data_stage_1__7750_, data_stage_1__7749_, data_stage_1__7748_, data_stage_1__7747_, data_stage_1__7746_, data_stage_1__7745_, data_stage_1__7744_, data_stage_1__7743_, data_stage_1__7742_, data_stage_1__7741_, data_stage_1__7740_, data_stage_1__7739_, data_stage_1__7738_, data_stage_1__7737_, data_stage_1__7736_, data_stage_1__7735_, data_stage_1__7734_, data_stage_1__7733_, data_stage_1__7732_, data_stage_1__7731_, data_stage_1__7730_, data_stage_1__7729_, data_stage_1__7728_, data_stage_1__7727_, data_stage_1__7726_, data_stage_1__7725_, data_stage_1__7724_, data_stage_1__7723_, data_stage_1__7722_, data_stage_1__7721_, data_stage_1__7720_, data_stage_1__7719_, data_stage_1__7718_, data_stage_1__7717_, data_stage_1__7716_, data_stage_1__7715_, data_stage_1__7714_, data_stage_1__7713_, data_stage_1__7712_, data_stage_1__7711_, data_stage_1__7710_, data_stage_1__7709_, data_stage_1__7708_, data_stage_1__7707_, data_stage_1__7706_, data_stage_1__7705_, data_stage_1__7704_, data_stage_1__7703_, data_stage_1__7702_, data_stage_1__7701_, data_stage_1__7700_, data_stage_1__7699_, data_stage_1__7698_, data_stage_1__7697_, data_stage_1__7696_, data_stage_1__7695_, data_stage_1__7694_, data_stage_1__7693_, data_stage_1__7692_, data_stage_1__7691_, data_stage_1__7690_, data_stage_1__7689_, data_stage_1__7688_, data_stage_1__7687_, data_stage_1__7686_, data_stage_1__7685_, data_stage_1__7684_, data_stage_1__7683_, data_stage_1__7682_, data_stage_1__7681_, data_stage_1__7680_ })
  );


  bsg_swap_width_p128
  mux_stage_0__mux_swap_31__swap_inst
  (
    .data_i(data_i[8191:7936]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__8191_, data_stage_1__8190_, data_stage_1__8189_, data_stage_1__8188_, data_stage_1__8187_, data_stage_1__8186_, data_stage_1__8185_, data_stage_1__8184_, data_stage_1__8183_, data_stage_1__8182_, data_stage_1__8181_, data_stage_1__8180_, data_stage_1__8179_, data_stage_1__8178_, data_stage_1__8177_, data_stage_1__8176_, data_stage_1__8175_, data_stage_1__8174_, data_stage_1__8173_, data_stage_1__8172_, data_stage_1__8171_, data_stage_1__8170_, data_stage_1__8169_, data_stage_1__8168_, data_stage_1__8167_, data_stage_1__8166_, data_stage_1__8165_, data_stage_1__8164_, data_stage_1__8163_, data_stage_1__8162_, data_stage_1__8161_, data_stage_1__8160_, data_stage_1__8159_, data_stage_1__8158_, data_stage_1__8157_, data_stage_1__8156_, data_stage_1__8155_, data_stage_1__8154_, data_stage_1__8153_, data_stage_1__8152_, data_stage_1__8151_, data_stage_1__8150_, data_stage_1__8149_, data_stage_1__8148_, data_stage_1__8147_, data_stage_1__8146_, data_stage_1__8145_, data_stage_1__8144_, data_stage_1__8143_, data_stage_1__8142_, data_stage_1__8141_, data_stage_1__8140_, data_stage_1__8139_, data_stage_1__8138_, data_stage_1__8137_, data_stage_1__8136_, data_stage_1__8135_, data_stage_1__8134_, data_stage_1__8133_, data_stage_1__8132_, data_stage_1__8131_, data_stage_1__8130_, data_stage_1__8129_, data_stage_1__8128_, data_stage_1__8127_, data_stage_1__8126_, data_stage_1__8125_, data_stage_1__8124_, data_stage_1__8123_, data_stage_1__8122_, data_stage_1__8121_, data_stage_1__8120_, data_stage_1__8119_, data_stage_1__8118_, data_stage_1__8117_, data_stage_1__8116_, data_stage_1__8115_, data_stage_1__8114_, data_stage_1__8113_, data_stage_1__8112_, data_stage_1__8111_, data_stage_1__8110_, data_stage_1__8109_, data_stage_1__8108_, data_stage_1__8107_, data_stage_1__8106_, data_stage_1__8105_, data_stage_1__8104_, data_stage_1__8103_, data_stage_1__8102_, data_stage_1__8101_, data_stage_1__8100_, data_stage_1__8099_, data_stage_1__8098_, data_stage_1__8097_, data_stage_1__8096_, data_stage_1__8095_, data_stage_1__8094_, data_stage_1__8093_, data_stage_1__8092_, data_stage_1__8091_, data_stage_1__8090_, data_stage_1__8089_, data_stage_1__8088_, data_stage_1__8087_, data_stage_1__8086_, data_stage_1__8085_, data_stage_1__8084_, data_stage_1__8083_, data_stage_1__8082_, data_stage_1__8081_, data_stage_1__8080_, data_stage_1__8079_, data_stage_1__8078_, data_stage_1__8077_, data_stage_1__8076_, data_stage_1__8075_, data_stage_1__8074_, data_stage_1__8073_, data_stage_1__8072_, data_stage_1__8071_, data_stage_1__8070_, data_stage_1__8069_, data_stage_1__8068_, data_stage_1__8067_, data_stage_1__8066_, data_stage_1__8065_, data_stage_1__8064_, data_stage_1__8063_, data_stage_1__8062_, data_stage_1__8061_, data_stage_1__8060_, data_stage_1__8059_, data_stage_1__8058_, data_stage_1__8057_, data_stage_1__8056_, data_stage_1__8055_, data_stage_1__8054_, data_stage_1__8053_, data_stage_1__8052_, data_stage_1__8051_, data_stage_1__8050_, data_stage_1__8049_, data_stage_1__8048_, data_stage_1__8047_, data_stage_1__8046_, data_stage_1__8045_, data_stage_1__8044_, data_stage_1__8043_, data_stage_1__8042_, data_stage_1__8041_, data_stage_1__8040_, data_stage_1__8039_, data_stage_1__8038_, data_stage_1__8037_, data_stage_1__8036_, data_stage_1__8035_, data_stage_1__8034_, data_stage_1__8033_, data_stage_1__8032_, data_stage_1__8031_, data_stage_1__8030_, data_stage_1__8029_, data_stage_1__8028_, data_stage_1__8027_, data_stage_1__8026_, data_stage_1__8025_, data_stage_1__8024_, data_stage_1__8023_, data_stage_1__8022_, data_stage_1__8021_, data_stage_1__8020_, data_stage_1__8019_, data_stage_1__8018_, data_stage_1__8017_, data_stage_1__8016_, data_stage_1__8015_, data_stage_1__8014_, data_stage_1__8013_, data_stage_1__8012_, data_stage_1__8011_, data_stage_1__8010_, data_stage_1__8009_, data_stage_1__8008_, data_stage_1__8007_, data_stage_1__8006_, data_stage_1__8005_, data_stage_1__8004_, data_stage_1__8003_, data_stage_1__8002_, data_stage_1__8001_, data_stage_1__8000_, data_stage_1__7999_, data_stage_1__7998_, data_stage_1__7997_, data_stage_1__7996_, data_stage_1__7995_, data_stage_1__7994_, data_stage_1__7993_, data_stage_1__7992_, data_stage_1__7991_, data_stage_1__7990_, data_stage_1__7989_, data_stage_1__7988_, data_stage_1__7987_, data_stage_1__7986_, data_stage_1__7985_, data_stage_1__7984_, data_stage_1__7983_, data_stage_1__7982_, data_stage_1__7981_, data_stage_1__7980_, data_stage_1__7979_, data_stage_1__7978_, data_stage_1__7977_, data_stage_1__7976_, data_stage_1__7975_, data_stage_1__7974_, data_stage_1__7973_, data_stage_1__7972_, data_stage_1__7971_, data_stage_1__7970_, data_stage_1__7969_, data_stage_1__7968_, data_stage_1__7967_, data_stage_1__7966_, data_stage_1__7965_, data_stage_1__7964_, data_stage_1__7963_, data_stage_1__7962_, data_stage_1__7961_, data_stage_1__7960_, data_stage_1__7959_, data_stage_1__7958_, data_stage_1__7957_, data_stage_1__7956_, data_stage_1__7955_, data_stage_1__7954_, data_stage_1__7953_, data_stage_1__7952_, data_stage_1__7951_, data_stage_1__7950_, data_stage_1__7949_, data_stage_1__7948_, data_stage_1__7947_, data_stage_1__7946_, data_stage_1__7945_, data_stage_1__7944_, data_stage_1__7943_, data_stage_1__7942_, data_stage_1__7941_, data_stage_1__7940_, data_stage_1__7939_, data_stage_1__7938_, data_stage_1__7937_, data_stage_1__7936_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_, data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_, data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_, data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_, data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_, data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_, data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_, data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_, data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_, data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_, data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_1__1023_, data_stage_1__1022_, data_stage_1__1021_, data_stage_1__1020_, data_stage_1__1019_, data_stage_1__1018_, data_stage_1__1017_, data_stage_1__1016_, data_stage_1__1015_, data_stage_1__1014_, data_stage_1__1013_, data_stage_1__1012_, data_stage_1__1011_, data_stage_1__1010_, data_stage_1__1009_, data_stage_1__1008_, data_stage_1__1007_, data_stage_1__1006_, data_stage_1__1005_, data_stage_1__1004_, data_stage_1__1003_, data_stage_1__1002_, data_stage_1__1001_, data_stage_1__1000_, data_stage_1__999_, data_stage_1__998_, data_stage_1__997_, data_stage_1__996_, data_stage_1__995_, data_stage_1__994_, data_stage_1__993_, data_stage_1__992_, data_stage_1__991_, data_stage_1__990_, data_stage_1__989_, data_stage_1__988_, data_stage_1__987_, data_stage_1__986_, data_stage_1__985_, data_stage_1__984_, data_stage_1__983_, data_stage_1__982_, data_stage_1__981_, data_stage_1__980_, data_stage_1__979_, data_stage_1__978_, data_stage_1__977_, data_stage_1__976_, data_stage_1__975_, data_stage_1__974_, data_stage_1__973_, data_stage_1__972_, data_stage_1__971_, data_stage_1__970_, data_stage_1__969_, data_stage_1__968_, data_stage_1__967_, data_stage_1__966_, data_stage_1__965_, data_stage_1__964_, data_stage_1__963_, data_stage_1__962_, data_stage_1__961_, data_stage_1__960_, data_stage_1__959_, data_stage_1__958_, data_stage_1__957_, data_stage_1__956_, data_stage_1__955_, data_stage_1__954_, data_stage_1__953_, data_stage_1__952_, data_stage_1__951_, data_stage_1__950_, data_stage_1__949_, data_stage_1__948_, data_stage_1__947_, data_stage_1__946_, data_stage_1__945_, data_stage_1__944_, data_stage_1__943_, data_stage_1__942_, data_stage_1__941_, data_stage_1__940_, data_stage_1__939_, data_stage_1__938_, data_stage_1__937_, data_stage_1__936_, data_stage_1__935_, data_stage_1__934_, data_stage_1__933_, data_stage_1__932_, data_stage_1__931_, data_stage_1__930_, data_stage_1__929_, data_stage_1__928_, data_stage_1__927_, data_stage_1__926_, data_stage_1__925_, data_stage_1__924_, data_stage_1__923_, data_stage_1__922_, data_stage_1__921_, data_stage_1__920_, data_stage_1__919_, data_stage_1__918_, data_stage_1__917_, data_stage_1__916_, data_stage_1__915_, data_stage_1__914_, data_stage_1__913_, data_stage_1__912_, data_stage_1__911_, data_stage_1__910_, data_stage_1__909_, data_stage_1__908_, data_stage_1__907_, data_stage_1__906_, data_stage_1__905_, data_stage_1__904_, data_stage_1__903_, data_stage_1__902_, data_stage_1__901_, data_stage_1__900_, data_stage_1__899_, data_stage_1__898_, data_stage_1__897_, data_stage_1__896_, data_stage_1__895_, data_stage_1__894_, data_stage_1__893_, data_stage_1__892_, data_stage_1__891_, data_stage_1__890_, data_stage_1__889_, data_stage_1__888_, data_stage_1__887_, data_stage_1__886_, data_stage_1__885_, data_stage_1__884_, data_stage_1__883_, data_stage_1__882_, data_stage_1__881_, data_stage_1__880_, data_stage_1__879_, data_stage_1__878_, data_stage_1__877_, data_stage_1__876_, data_stage_1__875_, data_stage_1__874_, data_stage_1__873_, data_stage_1__872_, data_stage_1__871_, data_stage_1__870_, data_stage_1__869_, data_stage_1__868_, data_stage_1__867_, data_stage_1__866_, data_stage_1__865_, data_stage_1__864_, data_stage_1__863_, data_stage_1__862_, data_stage_1__861_, data_stage_1__860_, data_stage_1__859_, data_stage_1__858_, data_stage_1__857_, data_stage_1__856_, data_stage_1__855_, data_stage_1__854_, data_stage_1__853_, data_stage_1__852_, data_stage_1__851_, data_stage_1__850_, data_stage_1__849_, data_stage_1__848_, data_stage_1__847_, data_stage_1__846_, data_stage_1__845_, data_stage_1__844_, data_stage_1__843_, data_stage_1__842_, data_stage_1__841_, data_stage_1__840_, data_stage_1__839_, data_stage_1__838_, data_stage_1__837_, data_stage_1__836_, data_stage_1__835_, data_stage_1__834_, data_stage_1__833_, data_stage_1__832_, data_stage_1__831_, data_stage_1__830_, data_stage_1__829_, data_stage_1__828_, data_stage_1__827_, data_stage_1__826_, data_stage_1__825_, data_stage_1__824_, data_stage_1__823_, data_stage_1__822_, data_stage_1__821_, data_stage_1__820_, data_stage_1__819_, data_stage_1__818_, data_stage_1__817_, data_stage_1__816_, data_stage_1__815_, data_stage_1__814_, data_stage_1__813_, data_stage_1__812_, data_stage_1__811_, data_stage_1__810_, data_stage_1__809_, data_stage_1__808_, data_stage_1__807_, data_stage_1__806_, data_stage_1__805_, data_stage_1__804_, data_stage_1__803_, data_stage_1__802_, data_stage_1__801_, data_stage_1__800_, data_stage_1__799_, data_stage_1__798_, data_stage_1__797_, data_stage_1__796_, data_stage_1__795_, data_stage_1__794_, data_stage_1__793_, data_stage_1__792_, data_stage_1__791_, data_stage_1__790_, data_stage_1__789_, data_stage_1__788_, data_stage_1__787_, data_stage_1__786_, data_stage_1__785_, data_stage_1__784_, data_stage_1__783_, data_stage_1__782_, data_stage_1__781_, data_stage_1__780_, data_stage_1__779_, data_stage_1__778_, data_stage_1__777_, data_stage_1__776_, data_stage_1__775_, data_stage_1__774_, data_stage_1__773_, data_stage_1__772_, data_stage_1__771_, data_stage_1__770_, data_stage_1__769_, data_stage_1__768_, data_stage_1__767_, data_stage_1__766_, data_stage_1__765_, data_stage_1__764_, data_stage_1__763_, data_stage_1__762_, data_stage_1__761_, data_stage_1__760_, data_stage_1__759_, data_stage_1__758_, data_stage_1__757_, data_stage_1__756_, data_stage_1__755_, data_stage_1__754_, data_stage_1__753_, data_stage_1__752_, data_stage_1__751_, data_stage_1__750_, data_stage_1__749_, data_stage_1__748_, data_stage_1__747_, data_stage_1__746_, data_stage_1__745_, data_stage_1__744_, data_stage_1__743_, data_stage_1__742_, data_stage_1__741_, data_stage_1__740_, data_stage_1__739_, data_stage_1__738_, data_stage_1__737_, data_stage_1__736_, data_stage_1__735_, data_stage_1__734_, data_stage_1__733_, data_stage_1__732_, data_stage_1__731_, data_stage_1__730_, data_stage_1__729_, data_stage_1__728_, data_stage_1__727_, data_stage_1__726_, data_stage_1__725_, data_stage_1__724_, data_stage_1__723_, data_stage_1__722_, data_stage_1__721_, data_stage_1__720_, data_stage_1__719_, data_stage_1__718_, data_stage_1__717_, data_stage_1__716_, data_stage_1__715_, data_stage_1__714_, data_stage_1__713_, data_stage_1__712_, data_stage_1__711_, data_stage_1__710_, data_stage_1__709_, data_stage_1__708_, data_stage_1__707_, data_stage_1__706_, data_stage_1__705_, data_stage_1__704_, data_stage_1__703_, data_stage_1__702_, data_stage_1__701_, data_stage_1__700_, data_stage_1__699_, data_stage_1__698_, data_stage_1__697_, data_stage_1__696_, data_stage_1__695_, data_stage_1__694_, data_stage_1__693_, data_stage_1__692_, data_stage_1__691_, data_stage_1__690_, data_stage_1__689_, data_stage_1__688_, data_stage_1__687_, data_stage_1__686_, data_stage_1__685_, data_stage_1__684_, data_stage_1__683_, data_stage_1__682_, data_stage_1__681_, data_stage_1__680_, data_stage_1__679_, data_stage_1__678_, data_stage_1__677_, data_stage_1__676_, data_stage_1__675_, data_stage_1__674_, data_stage_1__673_, data_stage_1__672_, data_stage_1__671_, data_stage_1__670_, data_stage_1__669_, data_stage_1__668_, data_stage_1__667_, data_stage_1__666_, data_stage_1__665_, data_stage_1__664_, data_stage_1__663_, data_stage_1__662_, data_stage_1__661_, data_stage_1__660_, data_stage_1__659_, data_stage_1__658_, data_stage_1__657_, data_stage_1__656_, data_stage_1__655_, data_stage_1__654_, data_stage_1__653_, data_stage_1__652_, data_stage_1__651_, data_stage_1__650_, data_stage_1__649_, data_stage_1__648_, data_stage_1__647_, data_stage_1__646_, data_stage_1__645_, data_stage_1__644_, data_stage_1__643_, data_stage_1__642_, data_stage_1__641_, data_stage_1__640_, data_stage_1__639_, data_stage_1__638_, data_stage_1__637_, data_stage_1__636_, data_stage_1__635_, data_stage_1__634_, data_stage_1__633_, data_stage_1__632_, data_stage_1__631_, data_stage_1__630_, data_stage_1__629_, data_stage_1__628_, data_stage_1__627_, data_stage_1__626_, data_stage_1__625_, data_stage_1__624_, data_stage_1__623_, data_stage_1__622_, data_stage_1__621_, data_stage_1__620_, data_stage_1__619_, data_stage_1__618_, data_stage_1__617_, data_stage_1__616_, data_stage_1__615_, data_stage_1__614_, data_stage_1__613_, data_stage_1__612_, data_stage_1__611_, data_stage_1__610_, data_stage_1__609_, data_stage_1__608_, data_stage_1__607_, data_stage_1__606_, data_stage_1__605_, data_stage_1__604_, data_stage_1__603_, data_stage_1__602_, data_stage_1__601_, data_stage_1__600_, data_stage_1__599_, data_stage_1__598_, data_stage_1__597_, data_stage_1__596_, data_stage_1__595_, data_stage_1__594_, data_stage_1__593_, data_stage_1__592_, data_stage_1__591_, data_stage_1__590_, data_stage_1__589_, data_stage_1__588_, data_stage_1__587_, data_stage_1__586_, data_stage_1__585_, data_stage_1__584_, data_stage_1__583_, data_stage_1__582_, data_stage_1__581_, data_stage_1__580_, data_stage_1__579_, data_stage_1__578_, data_stage_1__577_, data_stage_1__576_, data_stage_1__575_, data_stage_1__574_, data_stage_1__573_, data_stage_1__572_, data_stage_1__571_, data_stage_1__570_, data_stage_1__569_, data_stage_1__568_, data_stage_1__567_, data_stage_1__566_, data_stage_1__565_, data_stage_1__564_, data_stage_1__563_, data_stage_1__562_, data_stage_1__561_, data_stage_1__560_, data_stage_1__559_, data_stage_1__558_, data_stage_1__557_, data_stage_1__556_, data_stage_1__555_, data_stage_1__554_, data_stage_1__553_, data_stage_1__552_, data_stage_1__551_, data_stage_1__550_, data_stage_1__549_, data_stage_1__548_, data_stage_1__547_, data_stage_1__546_, data_stage_1__545_, data_stage_1__544_, data_stage_1__543_, data_stage_1__542_, data_stage_1__541_, data_stage_1__540_, data_stage_1__539_, data_stage_1__538_, data_stage_1__537_, data_stage_1__536_, data_stage_1__535_, data_stage_1__534_, data_stage_1__533_, data_stage_1__532_, data_stage_1__531_, data_stage_1__530_, data_stage_1__529_, data_stage_1__528_, data_stage_1__527_, data_stage_1__526_, data_stage_1__525_, data_stage_1__524_, data_stage_1__523_, data_stage_1__522_, data_stage_1__521_, data_stage_1__520_, data_stage_1__519_, data_stage_1__518_, data_stage_1__517_, data_stage_1__516_, data_stage_1__515_, data_stage_1__514_, data_stage_1__513_, data_stage_1__512_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__1023_, data_stage_2__1022_, data_stage_2__1021_, data_stage_2__1020_, data_stage_2__1019_, data_stage_2__1018_, data_stage_2__1017_, data_stage_2__1016_, data_stage_2__1015_, data_stage_2__1014_, data_stage_2__1013_, data_stage_2__1012_, data_stage_2__1011_, data_stage_2__1010_, data_stage_2__1009_, data_stage_2__1008_, data_stage_2__1007_, data_stage_2__1006_, data_stage_2__1005_, data_stage_2__1004_, data_stage_2__1003_, data_stage_2__1002_, data_stage_2__1001_, data_stage_2__1000_, data_stage_2__999_, data_stage_2__998_, data_stage_2__997_, data_stage_2__996_, data_stage_2__995_, data_stage_2__994_, data_stage_2__993_, data_stage_2__992_, data_stage_2__991_, data_stage_2__990_, data_stage_2__989_, data_stage_2__988_, data_stage_2__987_, data_stage_2__986_, data_stage_2__985_, data_stage_2__984_, data_stage_2__983_, data_stage_2__982_, data_stage_2__981_, data_stage_2__980_, data_stage_2__979_, data_stage_2__978_, data_stage_2__977_, data_stage_2__976_, data_stage_2__975_, data_stage_2__974_, data_stage_2__973_, data_stage_2__972_, data_stage_2__971_, data_stage_2__970_, data_stage_2__969_, data_stage_2__968_, data_stage_2__967_, data_stage_2__966_, data_stage_2__965_, data_stage_2__964_, data_stage_2__963_, data_stage_2__962_, data_stage_2__961_, data_stage_2__960_, data_stage_2__959_, data_stage_2__958_, data_stage_2__957_, data_stage_2__956_, data_stage_2__955_, data_stage_2__954_, data_stage_2__953_, data_stage_2__952_, data_stage_2__951_, data_stage_2__950_, data_stage_2__949_, data_stage_2__948_, data_stage_2__947_, data_stage_2__946_, data_stage_2__945_, data_stage_2__944_, data_stage_2__943_, data_stage_2__942_, data_stage_2__941_, data_stage_2__940_, data_stage_2__939_, data_stage_2__938_, data_stage_2__937_, data_stage_2__936_, data_stage_2__935_, data_stage_2__934_, data_stage_2__933_, data_stage_2__932_, data_stage_2__931_, data_stage_2__930_, data_stage_2__929_, data_stage_2__928_, data_stage_2__927_, data_stage_2__926_, data_stage_2__925_, data_stage_2__924_, data_stage_2__923_, data_stage_2__922_, data_stage_2__921_, data_stage_2__920_, data_stage_2__919_, data_stage_2__918_, data_stage_2__917_, data_stage_2__916_, data_stage_2__915_, data_stage_2__914_, data_stage_2__913_, data_stage_2__912_, data_stage_2__911_, data_stage_2__910_, data_stage_2__909_, data_stage_2__908_, data_stage_2__907_, data_stage_2__906_, data_stage_2__905_, data_stage_2__904_, data_stage_2__903_, data_stage_2__902_, data_stage_2__901_, data_stage_2__900_, data_stage_2__899_, data_stage_2__898_, data_stage_2__897_, data_stage_2__896_, data_stage_2__895_, data_stage_2__894_, data_stage_2__893_, data_stage_2__892_, data_stage_2__891_, data_stage_2__890_, data_stage_2__889_, data_stage_2__888_, data_stage_2__887_, data_stage_2__886_, data_stage_2__885_, data_stage_2__884_, data_stage_2__883_, data_stage_2__882_, data_stage_2__881_, data_stage_2__880_, data_stage_2__879_, data_stage_2__878_, data_stage_2__877_, data_stage_2__876_, data_stage_2__875_, data_stage_2__874_, data_stage_2__873_, data_stage_2__872_, data_stage_2__871_, data_stage_2__870_, data_stage_2__869_, data_stage_2__868_, data_stage_2__867_, data_stage_2__866_, data_stage_2__865_, data_stage_2__864_, data_stage_2__863_, data_stage_2__862_, data_stage_2__861_, data_stage_2__860_, data_stage_2__859_, data_stage_2__858_, data_stage_2__857_, data_stage_2__856_, data_stage_2__855_, data_stage_2__854_, data_stage_2__853_, data_stage_2__852_, data_stage_2__851_, data_stage_2__850_, data_stage_2__849_, data_stage_2__848_, data_stage_2__847_, data_stage_2__846_, data_stage_2__845_, data_stage_2__844_, data_stage_2__843_, data_stage_2__842_, data_stage_2__841_, data_stage_2__840_, data_stage_2__839_, data_stage_2__838_, data_stage_2__837_, data_stage_2__836_, data_stage_2__835_, data_stage_2__834_, data_stage_2__833_, data_stage_2__832_, data_stage_2__831_, data_stage_2__830_, data_stage_2__829_, data_stage_2__828_, data_stage_2__827_, data_stage_2__826_, data_stage_2__825_, data_stage_2__824_, data_stage_2__823_, data_stage_2__822_, data_stage_2__821_, data_stage_2__820_, data_stage_2__819_, data_stage_2__818_, data_stage_2__817_, data_stage_2__816_, data_stage_2__815_, data_stage_2__814_, data_stage_2__813_, data_stage_2__812_, data_stage_2__811_, data_stage_2__810_, data_stage_2__809_, data_stage_2__808_, data_stage_2__807_, data_stage_2__806_, data_stage_2__805_, data_stage_2__804_, data_stage_2__803_, data_stage_2__802_, data_stage_2__801_, data_stage_2__800_, data_stage_2__799_, data_stage_2__798_, data_stage_2__797_, data_stage_2__796_, data_stage_2__795_, data_stage_2__794_, data_stage_2__793_, data_stage_2__792_, data_stage_2__791_, data_stage_2__790_, data_stage_2__789_, data_stage_2__788_, data_stage_2__787_, data_stage_2__786_, data_stage_2__785_, data_stage_2__784_, data_stage_2__783_, data_stage_2__782_, data_stage_2__781_, data_stage_2__780_, data_stage_2__779_, data_stage_2__778_, data_stage_2__777_, data_stage_2__776_, data_stage_2__775_, data_stage_2__774_, data_stage_2__773_, data_stage_2__772_, data_stage_2__771_, data_stage_2__770_, data_stage_2__769_, data_stage_2__768_, data_stage_2__767_, data_stage_2__766_, data_stage_2__765_, data_stage_2__764_, data_stage_2__763_, data_stage_2__762_, data_stage_2__761_, data_stage_2__760_, data_stage_2__759_, data_stage_2__758_, data_stage_2__757_, data_stage_2__756_, data_stage_2__755_, data_stage_2__754_, data_stage_2__753_, data_stage_2__752_, data_stage_2__751_, data_stage_2__750_, data_stage_2__749_, data_stage_2__748_, data_stage_2__747_, data_stage_2__746_, data_stage_2__745_, data_stage_2__744_, data_stage_2__743_, data_stage_2__742_, data_stage_2__741_, data_stage_2__740_, data_stage_2__739_, data_stage_2__738_, data_stage_2__737_, data_stage_2__736_, data_stage_2__735_, data_stage_2__734_, data_stage_2__733_, data_stage_2__732_, data_stage_2__731_, data_stage_2__730_, data_stage_2__729_, data_stage_2__728_, data_stage_2__727_, data_stage_2__726_, data_stage_2__725_, data_stage_2__724_, data_stage_2__723_, data_stage_2__722_, data_stage_2__721_, data_stage_2__720_, data_stage_2__719_, data_stage_2__718_, data_stage_2__717_, data_stage_2__716_, data_stage_2__715_, data_stage_2__714_, data_stage_2__713_, data_stage_2__712_, data_stage_2__711_, data_stage_2__710_, data_stage_2__709_, data_stage_2__708_, data_stage_2__707_, data_stage_2__706_, data_stage_2__705_, data_stage_2__704_, data_stage_2__703_, data_stage_2__702_, data_stage_2__701_, data_stage_2__700_, data_stage_2__699_, data_stage_2__698_, data_stage_2__697_, data_stage_2__696_, data_stage_2__695_, data_stage_2__694_, data_stage_2__693_, data_stage_2__692_, data_stage_2__691_, data_stage_2__690_, data_stage_2__689_, data_stage_2__688_, data_stage_2__687_, data_stage_2__686_, data_stage_2__685_, data_stage_2__684_, data_stage_2__683_, data_stage_2__682_, data_stage_2__681_, data_stage_2__680_, data_stage_2__679_, data_stage_2__678_, data_stage_2__677_, data_stage_2__676_, data_stage_2__675_, data_stage_2__674_, data_stage_2__673_, data_stage_2__672_, data_stage_2__671_, data_stage_2__670_, data_stage_2__669_, data_stage_2__668_, data_stage_2__667_, data_stage_2__666_, data_stage_2__665_, data_stage_2__664_, data_stage_2__663_, data_stage_2__662_, data_stage_2__661_, data_stage_2__660_, data_stage_2__659_, data_stage_2__658_, data_stage_2__657_, data_stage_2__656_, data_stage_2__655_, data_stage_2__654_, data_stage_2__653_, data_stage_2__652_, data_stage_2__651_, data_stage_2__650_, data_stage_2__649_, data_stage_2__648_, data_stage_2__647_, data_stage_2__646_, data_stage_2__645_, data_stage_2__644_, data_stage_2__643_, data_stage_2__642_, data_stage_2__641_, data_stage_2__640_, data_stage_2__639_, data_stage_2__638_, data_stage_2__637_, data_stage_2__636_, data_stage_2__635_, data_stage_2__634_, data_stage_2__633_, data_stage_2__632_, data_stage_2__631_, data_stage_2__630_, data_stage_2__629_, data_stage_2__628_, data_stage_2__627_, data_stage_2__626_, data_stage_2__625_, data_stage_2__624_, data_stage_2__623_, data_stage_2__622_, data_stage_2__621_, data_stage_2__620_, data_stage_2__619_, data_stage_2__618_, data_stage_2__617_, data_stage_2__616_, data_stage_2__615_, data_stage_2__614_, data_stage_2__613_, data_stage_2__612_, data_stage_2__611_, data_stage_2__610_, data_stage_2__609_, data_stage_2__608_, data_stage_2__607_, data_stage_2__606_, data_stage_2__605_, data_stage_2__604_, data_stage_2__603_, data_stage_2__602_, data_stage_2__601_, data_stage_2__600_, data_stage_2__599_, data_stage_2__598_, data_stage_2__597_, data_stage_2__596_, data_stage_2__595_, data_stage_2__594_, data_stage_2__593_, data_stage_2__592_, data_stage_2__591_, data_stage_2__590_, data_stage_2__589_, data_stage_2__588_, data_stage_2__587_, data_stage_2__586_, data_stage_2__585_, data_stage_2__584_, data_stage_2__583_, data_stage_2__582_, data_stage_2__581_, data_stage_2__580_, data_stage_2__579_, data_stage_2__578_, data_stage_2__577_, data_stage_2__576_, data_stage_2__575_, data_stage_2__574_, data_stage_2__573_, data_stage_2__572_, data_stage_2__571_, data_stage_2__570_, data_stage_2__569_, data_stage_2__568_, data_stage_2__567_, data_stage_2__566_, data_stage_2__565_, data_stage_2__564_, data_stage_2__563_, data_stage_2__562_, data_stage_2__561_, data_stage_2__560_, data_stage_2__559_, data_stage_2__558_, data_stage_2__557_, data_stage_2__556_, data_stage_2__555_, data_stage_2__554_, data_stage_2__553_, data_stage_2__552_, data_stage_2__551_, data_stage_2__550_, data_stage_2__549_, data_stage_2__548_, data_stage_2__547_, data_stage_2__546_, data_stage_2__545_, data_stage_2__544_, data_stage_2__543_, data_stage_2__542_, data_stage_2__541_, data_stage_2__540_, data_stage_2__539_, data_stage_2__538_, data_stage_2__537_, data_stage_2__536_, data_stage_2__535_, data_stage_2__534_, data_stage_2__533_, data_stage_2__532_, data_stage_2__531_, data_stage_2__530_, data_stage_2__529_, data_stage_2__528_, data_stage_2__527_, data_stage_2__526_, data_stage_2__525_, data_stage_2__524_, data_stage_2__523_, data_stage_2__522_, data_stage_2__521_, data_stage_2__520_, data_stage_2__519_, data_stage_2__518_, data_stage_2__517_, data_stage_2__516_, data_stage_2__515_, data_stage_2__514_, data_stage_2__513_, data_stage_2__512_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_2__swap_inst
  (
    .data_i({ data_stage_1__1535_, data_stage_1__1534_, data_stage_1__1533_, data_stage_1__1532_, data_stage_1__1531_, data_stage_1__1530_, data_stage_1__1529_, data_stage_1__1528_, data_stage_1__1527_, data_stage_1__1526_, data_stage_1__1525_, data_stage_1__1524_, data_stage_1__1523_, data_stage_1__1522_, data_stage_1__1521_, data_stage_1__1520_, data_stage_1__1519_, data_stage_1__1518_, data_stage_1__1517_, data_stage_1__1516_, data_stage_1__1515_, data_stage_1__1514_, data_stage_1__1513_, data_stage_1__1512_, data_stage_1__1511_, data_stage_1__1510_, data_stage_1__1509_, data_stage_1__1508_, data_stage_1__1507_, data_stage_1__1506_, data_stage_1__1505_, data_stage_1__1504_, data_stage_1__1503_, data_stage_1__1502_, data_stage_1__1501_, data_stage_1__1500_, data_stage_1__1499_, data_stage_1__1498_, data_stage_1__1497_, data_stage_1__1496_, data_stage_1__1495_, data_stage_1__1494_, data_stage_1__1493_, data_stage_1__1492_, data_stage_1__1491_, data_stage_1__1490_, data_stage_1__1489_, data_stage_1__1488_, data_stage_1__1487_, data_stage_1__1486_, data_stage_1__1485_, data_stage_1__1484_, data_stage_1__1483_, data_stage_1__1482_, data_stage_1__1481_, data_stage_1__1480_, data_stage_1__1479_, data_stage_1__1478_, data_stage_1__1477_, data_stage_1__1476_, data_stage_1__1475_, data_stage_1__1474_, data_stage_1__1473_, data_stage_1__1472_, data_stage_1__1471_, data_stage_1__1470_, data_stage_1__1469_, data_stage_1__1468_, data_stage_1__1467_, data_stage_1__1466_, data_stage_1__1465_, data_stage_1__1464_, data_stage_1__1463_, data_stage_1__1462_, data_stage_1__1461_, data_stage_1__1460_, data_stage_1__1459_, data_stage_1__1458_, data_stage_1__1457_, data_stage_1__1456_, data_stage_1__1455_, data_stage_1__1454_, data_stage_1__1453_, data_stage_1__1452_, data_stage_1__1451_, data_stage_1__1450_, data_stage_1__1449_, data_stage_1__1448_, data_stage_1__1447_, data_stage_1__1446_, data_stage_1__1445_, data_stage_1__1444_, data_stage_1__1443_, data_stage_1__1442_, data_stage_1__1441_, data_stage_1__1440_, data_stage_1__1439_, data_stage_1__1438_, data_stage_1__1437_, data_stage_1__1436_, data_stage_1__1435_, data_stage_1__1434_, data_stage_1__1433_, data_stage_1__1432_, data_stage_1__1431_, data_stage_1__1430_, data_stage_1__1429_, data_stage_1__1428_, data_stage_1__1427_, data_stage_1__1426_, data_stage_1__1425_, data_stage_1__1424_, data_stage_1__1423_, data_stage_1__1422_, data_stage_1__1421_, data_stage_1__1420_, data_stage_1__1419_, data_stage_1__1418_, data_stage_1__1417_, data_stage_1__1416_, data_stage_1__1415_, data_stage_1__1414_, data_stage_1__1413_, data_stage_1__1412_, data_stage_1__1411_, data_stage_1__1410_, data_stage_1__1409_, data_stage_1__1408_, data_stage_1__1407_, data_stage_1__1406_, data_stage_1__1405_, data_stage_1__1404_, data_stage_1__1403_, data_stage_1__1402_, data_stage_1__1401_, data_stage_1__1400_, data_stage_1__1399_, data_stage_1__1398_, data_stage_1__1397_, data_stage_1__1396_, data_stage_1__1395_, data_stage_1__1394_, data_stage_1__1393_, data_stage_1__1392_, data_stage_1__1391_, data_stage_1__1390_, data_stage_1__1389_, data_stage_1__1388_, data_stage_1__1387_, data_stage_1__1386_, data_stage_1__1385_, data_stage_1__1384_, data_stage_1__1383_, data_stage_1__1382_, data_stage_1__1381_, data_stage_1__1380_, data_stage_1__1379_, data_stage_1__1378_, data_stage_1__1377_, data_stage_1__1376_, data_stage_1__1375_, data_stage_1__1374_, data_stage_1__1373_, data_stage_1__1372_, data_stage_1__1371_, data_stage_1__1370_, data_stage_1__1369_, data_stage_1__1368_, data_stage_1__1367_, data_stage_1__1366_, data_stage_1__1365_, data_stage_1__1364_, data_stage_1__1363_, data_stage_1__1362_, data_stage_1__1361_, data_stage_1__1360_, data_stage_1__1359_, data_stage_1__1358_, data_stage_1__1357_, data_stage_1__1356_, data_stage_1__1355_, data_stage_1__1354_, data_stage_1__1353_, data_stage_1__1352_, data_stage_1__1351_, data_stage_1__1350_, data_stage_1__1349_, data_stage_1__1348_, data_stage_1__1347_, data_stage_1__1346_, data_stage_1__1345_, data_stage_1__1344_, data_stage_1__1343_, data_stage_1__1342_, data_stage_1__1341_, data_stage_1__1340_, data_stage_1__1339_, data_stage_1__1338_, data_stage_1__1337_, data_stage_1__1336_, data_stage_1__1335_, data_stage_1__1334_, data_stage_1__1333_, data_stage_1__1332_, data_stage_1__1331_, data_stage_1__1330_, data_stage_1__1329_, data_stage_1__1328_, data_stage_1__1327_, data_stage_1__1326_, data_stage_1__1325_, data_stage_1__1324_, data_stage_1__1323_, data_stage_1__1322_, data_stage_1__1321_, data_stage_1__1320_, data_stage_1__1319_, data_stage_1__1318_, data_stage_1__1317_, data_stage_1__1316_, data_stage_1__1315_, data_stage_1__1314_, data_stage_1__1313_, data_stage_1__1312_, data_stage_1__1311_, data_stage_1__1310_, data_stage_1__1309_, data_stage_1__1308_, data_stage_1__1307_, data_stage_1__1306_, data_stage_1__1305_, data_stage_1__1304_, data_stage_1__1303_, data_stage_1__1302_, data_stage_1__1301_, data_stage_1__1300_, data_stage_1__1299_, data_stage_1__1298_, data_stage_1__1297_, data_stage_1__1296_, data_stage_1__1295_, data_stage_1__1294_, data_stage_1__1293_, data_stage_1__1292_, data_stage_1__1291_, data_stage_1__1290_, data_stage_1__1289_, data_stage_1__1288_, data_stage_1__1287_, data_stage_1__1286_, data_stage_1__1285_, data_stage_1__1284_, data_stage_1__1283_, data_stage_1__1282_, data_stage_1__1281_, data_stage_1__1280_, data_stage_1__1279_, data_stage_1__1278_, data_stage_1__1277_, data_stage_1__1276_, data_stage_1__1275_, data_stage_1__1274_, data_stage_1__1273_, data_stage_1__1272_, data_stage_1__1271_, data_stage_1__1270_, data_stage_1__1269_, data_stage_1__1268_, data_stage_1__1267_, data_stage_1__1266_, data_stage_1__1265_, data_stage_1__1264_, data_stage_1__1263_, data_stage_1__1262_, data_stage_1__1261_, data_stage_1__1260_, data_stage_1__1259_, data_stage_1__1258_, data_stage_1__1257_, data_stage_1__1256_, data_stage_1__1255_, data_stage_1__1254_, data_stage_1__1253_, data_stage_1__1252_, data_stage_1__1251_, data_stage_1__1250_, data_stage_1__1249_, data_stage_1__1248_, data_stage_1__1247_, data_stage_1__1246_, data_stage_1__1245_, data_stage_1__1244_, data_stage_1__1243_, data_stage_1__1242_, data_stage_1__1241_, data_stage_1__1240_, data_stage_1__1239_, data_stage_1__1238_, data_stage_1__1237_, data_stage_1__1236_, data_stage_1__1235_, data_stage_1__1234_, data_stage_1__1233_, data_stage_1__1232_, data_stage_1__1231_, data_stage_1__1230_, data_stage_1__1229_, data_stage_1__1228_, data_stage_1__1227_, data_stage_1__1226_, data_stage_1__1225_, data_stage_1__1224_, data_stage_1__1223_, data_stage_1__1222_, data_stage_1__1221_, data_stage_1__1220_, data_stage_1__1219_, data_stage_1__1218_, data_stage_1__1217_, data_stage_1__1216_, data_stage_1__1215_, data_stage_1__1214_, data_stage_1__1213_, data_stage_1__1212_, data_stage_1__1211_, data_stage_1__1210_, data_stage_1__1209_, data_stage_1__1208_, data_stage_1__1207_, data_stage_1__1206_, data_stage_1__1205_, data_stage_1__1204_, data_stage_1__1203_, data_stage_1__1202_, data_stage_1__1201_, data_stage_1__1200_, data_stage_1__1199_, data_stage_1__1198_, data_stage_1__1197_, data_stage_1__1196_, data_stage_1__1195_, data_stage_1__1194_, data_stage_1__1193_, data_stage_1__1192_, data_stage_1__1191_, data_stage_1__1190_, data_stage_1__1189_, data_stage_1__1188_, data_stage_1__1187_, data_stage_1__1186_, data_stage_1__1185_, data_stage_1__1184_, data_stage_1__1183_, data_stage_1__1182_, data_stage_1__1181_, data_stage_1__1180_, data_stage_1__1179_, data_stage_1__1178_, data_stage_1__1177_, data_stage_1__1176_, data_stage_1__1175_, data_stage_1__1174_, data_stage_1__1173_, data_stage_1__1172_, data_stage_1__1171_, data_stage_1__1170_, data_stage_1__1169_, data_stage_1__1168_, data_stage_1__1167_, data_stage_1__1166_, data_stage_1__1165_, data_stage_1__1164_, data_stage_1__1163_, data_stage_1__1162_, data_stage_1__1161_, data_stage_1__1160_, data_stage_1__1159_, data_stage_1__1158_, data_stage_1__1157_, data_stage_1__1156_, data_stage_1__1155_, data_stage_1__1154_, data_stage_1__1153_, data_stage_1__1152_, data_stage_1__1151_, data_stage_1__1150_, data_stage_1__1149_, data_stage_1__1148_, data_stage_1__1147_, data_stage_1__1146_, data_stage_1__1145_, data_stage_1__1144_, data_stage_1__1143_, data_stage_1__1142_, data_stage_1__1141_, data_stage_1__1140_, data_stage_1__1139_, data_stage_1__1138_, data_stage_1__1137_, data_stage_1__1136_, data_stage_1__1135_, data_stage_1__1134_, data_stage_1__1133_, data_stage_1__1132_, data_stage_1__1131_, data_stage_1__1130_, data_stage_1__1129_, data_stage_1__1128_, data_stage_1__1127_, data_stage_1__1126_, data_stage_1__1125_, data_stage_1__1124_, data_stage_1__1123_, data_stage_1__1122_, data_stage_1__1121_, data_stage_1__1120_, data_stage_1__1119_, data_stage_1__1118_, data_stage_1__1117_, data_stage_1__1116_, data_stage_1__1115_, data_stage_1__1114_, data_stage_1__1113_, data_stage_1__1112_, data_stage_1__1111_, data_stage_1__1110_, data_stage_1__1109_, data_stage_1__1108_, data_stage_1__1107_, data_stage_1__1106_, data_stage_1__1105_, data_stage_1__1104_, data_stage_1__1103_, data_stage_1__1102_, data_stage_1__1101_, data_stage_1__1100_, data_stage_1__1099_, data_stage_1__1098_, data_stage_1__1097_, data_stage_1__1096_, data_stage_1__1095_, data_stage_1__1094_, data_stage_1__1093_, data_stage_1__1092_, data_stage_1__1091_, data_stage_1__1090_, data_stage_1__1089_, data_stage_1__1088_, data_stage_1__1087_, data_stage_1__1086_, data_stage_1__1085_, data_stage_1__1084_, data_stage_1__1083_, data_stage_1__1082_, data_stage_1__1081_, data_stage_1__1080_, data_stage_1__1079_, data_stage_1__1078_, data_stage_1__1077_, data_stage_1__1076_, data_stage_1__1075_, data_stage_1__1074_, data_stage_1__1073_, data_stage_1__1072_, data_stage_1__1071_, data_stage_1__1070_, data_stage_1__1069_, data_stage_1__1068_, data_stage_1__1067_, data_stage_1__1066_, data_stage_1__1065_, data_stage_1__1064_, data_stage_1__1063_, data_stage_1__1062_, data_stage_1__1061_, data_stage_1__1060_, data_stage_1__1059_, data_stage_1__1058_, data_stage_1__1057_, data_stage_1__1056_, data_stage_1__1055_, data_stage_1__1054_, data_stage_1__1053_, data_stage_1__1052_, data_stage_1__1051_, data_stage_1__1050_, data_stage_1__1049_, data_stage_1__1048_, data_stage_1__1047_, data_stage_1__1046_, data_stage_1__1045_, data_stage_1__1044_, data_stage_1__1043_, data_stage_1__1042_, data_stage_1__1041_, data_stage_1__1040_, data_stage_1__1039_, data_stage_1__1038_, data_stage_1__1037_, data_stage_1__1036_, data_stage_1__1035_, data_stage_1__1034_, data_stage_1__1033_, data_stage_1__1032_, data_stage_1__1031_, data_stage_1__1030_, data_stage_1__1029_, data_stage_1__1028_, data_stage_1__1027_, data_stage_1__1026_, data_stage_1__1025_, data_stage_1__1024_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__1535_, data_stage_2__1534_, data_stage_2__1533_, data_stage_2__1532_, data_stage_2__1531_, data_stage_2__1530_, data_stage_2__1529_, data_stage_2__1528_, data_stage_2__1527_, data_stage_2__1526_, data_stage_2__1525_, data_stage_2__1524_, data_stage_2__1523_, data_stage_2__1522_, data_stage_2__1521_, data_stage_2__1520_, data_stage_2__1519_, data_stage_2__1518_, data_stage_2__1517_, data_stage_2__1516_, data_stage_2__1515_, data_stage_2__1514_, data_stage_2__1513_, data_stage_2__1512_, data_stage_2__1511_, data_stage_2__1510_, data_stage_2__1509_, data_stage_2__1508_, data_stage_2__1507_, data_stage_2__1506_, data_stage_2__1505_, data_stage_2__1504_, data_stage_2__1503_, data_stage_2__1502_, data_stage_2__1501_, data_stage_2__1500_, data_stage_2__1499_, data_stage_2__1498_, data_stage_2__1497_, data_stage_2__1496_, data_stage_2__1495_, data_stage_2__1494_, data_stage_2__1493_, data_stage_2__1492_, data_stage_2__1491_, data_stage_2__1490_, data_stage_2__1489_, data_stage_2__1488_, data_stage_2__1487_, data_stage_2__1486_, data_stage_2__1485_, data_stage_2__1484_, data_stage_2__1483_, data_stage_2__1482_, data_stage_2__1481_, data_stage_2__1480_, data_stage_2__1479_, data_stage_2__1478_, data_stage_2__1477_, data_stage_2__1476_, data_stage_2__1475_, data_stage_2__1474_, data_stage_2__1473_, data_stage_2__1472_, data_stage_2__1471_, data_stage_2__1470_, data_stage_2__1469_, data_stage_2__1468_, data_stage_2__1467_, data_stage_2__1466_, data_stage_2__1465_, data_stage_2__1464_, data_stage_2__1463_, data_stage_2__1462_, data_stage_2__1461_, data_stage_2__1460_, data_stage_2__1459_, data_stage_2__1458_, data_stage_2__1457_, data_stage_2__1456_, data_stage_2__1455_, data_stage_2__1454_, data_stage_2__1453_, data_stage_2__1452_, data_stage_2__1451_, data_stage_2__1450_, data_stage_2__1449_, data_stage_2__1448_, data_stage_2__1447_, data_stage_2__1446_, data_stage_2__1445_, data_stage_2__1444_, data_stage_2__1443_, data_stage_2__1442_, data_stage_2__1441_, data_stage_2__1440_, data_stage_2__1439_, data_stage_2__1438_, data_stage_2__1437_, data_stage_2__1436_, data_stage_2__1435_, data_stage_2__1434_, data_stage_2__1433_, data_stage_2__1432_, data_stage_2__1431_, data_stage_2__1430_, data_stage_2__1429_, data_stage_2__1428_, data_stage_2__1427_, data_stage_2__1426_, data_stage_2__1425_, data_stage_2__1424_, data_stage_2__1423_, data_stage_2__1422_, data_stage_2__1421_, data_stage_2__1420_, data_stage_2__1419_, data_stage_2__1418_, data_stage_2__1417_, data_stage_2__1416_, data_stage_2__1415_, data_stage_2__1414_, data_stage_2__1413_, data_stage_2__1412_, data_stage_2__1411_, data_stage_2__1410_, data_stage_2__1409_, data_stage_2__1408_, data_stage_2__1407_, data_stage_2__1406_, data_stage_2__1405_, data_stage_2__1404_, data_stage_2__1403_, data_stage_2__1402_, data_stage_2__1401_, data_stage_2__1400_, data_stage_2__1399_, data_stage_2__1398_, data_stage_2__1397_, data_stage_2__1396_, data_stage_2__1395_, data_stage_2__1394_, data_stage_2__1393_, data_stage_2__1392_, data_stage_2__1391_, data_stage_2__1390_, data_stage_2__1389_, data_stage_2__1388_, data_stage_2__1387_, data_stage_2__1386_, data_stage_2__1385_, data_stage_2__1384_, data_stage_2__1383_, data_stage_2__1382_, data_stage_2__1381_, data_stage_2__1380_, data_stage_2__1379_, data_stage_2__1378_, data_stage_2__1377_, data_stage_2__1376_, data_stage_2__1375_, data_stage_2__1374_, data_stage_2__1373_, data_stage_2__1372_, data_stage_2__1371_, data_stage_2__1370_, data_stage_2__1369_, data_stage_2__1368_, data_stage_2__1367_, data_stage_2__1366_, data_stage_2__1365_, data_stage_2__1364_, data_stage_2__1363_, data_stage_2__1362_, data_stage_2__1361_, data_stage_2__1360_, data_stage_2__1359_, data_stage_2__1358_, data_stage_2__1357_, data_stage_2__1356_, data_stage_2__1355_, data_stage_2__1354_, data_stage_2__1353_, data_stage_2__1352_, data_stage_2__1351_, data_stage_2__1350_, data_stage_2__1349_, data_stage_2__1348_, data_stage_2__1347_, data_stage_2__1346_, data_stage_2__1345_, data_stage_2__1344_, data_stage_2__1343_, data_stage_2__1342_, data_stage_2__1341_, data_stage_2__1340_, data_stage_2__1339_, data_stage_2__1338_, data_stage_2__1337_, data_stage_2__1336_, data_stage_2__1335_, data_stage_2__1334_, data_stage_2__1333_, data_stage_2__1332_, data_stage_2__1331_, data_stage_2__1330_, data_stage_2__1329_, data_stage_2__1328_, data_stage_2__1327_, data_stage_2__1326_, data_stage_2__1325_, data_stage_2__1324_, data_stage_2__1323_, data_stage_2__1322_, data_stage_2__1321_, data_stage_2__1320_, data_stage_2__1319_, data_stage_2__1318_, data_stage_2__1317_, data_stage_2__1316_, data_stage_2__1315_, data_stage_2__1314_, data_stage_2__1313_, data_stage_2__1312_, data_stage_2__1311_, data_stage_2__1310_, data_stage_2__1309_, data_stage_2__1308_, data_stage_2__1307_, data_stage_2__1306_, data_stage_2__1305_, data_stage_2__1304_, data_stage_2__1303_, data_stage_2__1302_, data_stage_2__1301_, data_stage_2__1300_, data_stage_2__1299_, data_stage_2__1298_, data_stage_2__1297_, data_stage_2__1296_, data_stage_2__1295_, data_stage_2__1294_, data_stage_2__1293_, data_stage_2__1292_, data_stage_2__1291_, data_stage_2__1290_, data_stage_2__1289_, data_stage_2__1288_, data_stage_2__1287_, data_stage_2__1286_, data_stage_2__1285_, data_stage_2__1284_, data_stage_2__1283_, data_stage_2__1282_, data_stage_2__1281_, data_stage_2__1280_, data_stage_2__1279_, data_stage_2__1278_, data_stage_2__1277_, data_stage_2__1276_, data_stage_2__1275_, data_stage_2__1274_, data_stage_2__1273_, data_stage_2__1272_, data_stage_2__1271_, data_stage_2__1270_, data_stage_2__1269_, data_stage_2__1268_, data_stage_2__1267_, data_stage_2__1266_, data_stage_2__1265_, data_stage_2__1264_, data_stage_2__1263_, data_stage_2__1262_, data_stage_2__1261_, data_stage_2__1260_, data_stage_2__1259_, data_stage_2__1258_, data_stage_2__1257_, data_stage_2__1256_, data_stage_2__1255_, data_stage_2__1254_, data_stage_2__1253_, data_stage_2__1252_, data_stage_2__1251_, data_stage_2__1250_, data_stage_2__1249_, data_stage_2__1248_, data_stage_2__1247_, data_stage_2__1246_, data_stage_2__1245_, data_stage_2__1244_, data_stage_2__1243_, data_stage_2__1242_, data_stage_2__1241_, data_stage_2__1240_, data_stage_2__1239_, data_stage_2__1238_, data_stage_2__1237_, data_stage_2__1236_, data_stage_2__1235_, data_stage_2__1234_, data_stage_2__1233_, data_stage_2__1232_, data_stage_2__1231_, data_stage_2__1230_, data_stage_2__1229_, data_stage_2__1228_, data_stage_2__1227_, data_stage_2__1226_, data_stage_2__1225_, data_stage_2__1224_, data_stage_2__1223_, data_stage_2__1222_, data_stage_2__1221_, data_stage_2__1220_, data_stage_2__1219_, data_stage_2__1218_, data_stage_2__1217_, data_stage_2__1216_, data_stage_2__1215_, data_stage_2__1214_, data_stage_2__1213_, data_stage_2__1212_, data_stage_2__1211_, data_stage_2__1210_, data_stage_2__1209_, data_stage_2__1208_, data_stage_2__1207_, data_stage_2__1206_, data_stage_2__1205_, data_stage_2__1204_, data_stage_2__1203_, data_stage_2__1202_, data_stage_2__1201_, data_stage_2__1200_, data_stage_2__1199_, data_stage_2__1198_, data_stage_2__1197_, data_stage_2__1196_, data_stage_2__1195_, data_stage_2__1194_, data_stage_2__1193_, data_stage_2__1192_, data_stage_2__1191_, data_stage_2__1190_, data_stage_2__1189_, data_stage_2__1188_, data_stage_2__1187_, data_stage_2__1186_, data_stage_2__1185_, data_stage_2__1184_, data_stage_2__1183_, data_stage_2__1182_, data_stage_2__1181_, data_stage_2__1180_, data_stage_2__1179_, data_stage_2__1178_, data_stage_2__1177_, data_stage_2__1176_, data_stage_2__1175_, data_stage_2__1174_, data_stage_2__1173_, data_stage_2__1172_, data_stage_2__1171_, data_stage_2__1170_, data_stage_2__1169_, data_stage_2__1168_, data_stage_2__1167_, data_stage_2__1166_, data_stage_2__1165_, data_stage_2__1164_, data_stage_2__1163_, data_stage_2__1162_, data_stage_2__1161_, data_stage_2__1160_, data_stage_2__1159_, data_stage_2__1158_, data_stage_2__1157_, data_stage_2__1156_, data_stage_2__1155_, data_stage_2__1154_, data_stage_2__1153_, data_stage_2__1152_, data_stage_2__1151_, data_stage_2__1150_, data_stage_2__1149_, data_stage_2__1148_, data_stage_2__1147_, data_stage_2__1146_, data_stage_2__1145_, data_stage_2__1144_, data_stage_2__1143_, data_stage_2__1142_, data_stage_2__1141_, data_stage_2__1140_, data_stage_2__1139_, data_stage_2__1138_, data_stage_2__1137_, data_stage_2__1136_, data_stage_2__1135_, data_stage_2__1134_, data_stage_2__1133_, data_stage_2__1132_, data_stage_2__1131_, data_stage_2__1130_, data_stage_2__1129_, data_stage_2__1128_, data_stage_2__1127_, data_stage_2__1126_, data_stage_2__1125_, data_stage_2__1124_, data_stage_2__1123_, data_stage_2__1122_, data_stage_2__1121_, data_stage_2__1120_, data_stage_2__1119_, data_stage_2__1118_, data_stage_2__1117_, data_stage_2__1116_, data_stage_2__1115_, data_stage_2__1114_, data_stage_2__1113_, data_stage_2__1112_, data_stage_2__1111_, data_stage_2__1110_, data_stage_2__1109_, data_stage_2__1108_, data_stage_2__1107_, data_stage_2__1106_, data_stage_2__1105_, data_stage_2__1104_, data_stage_2__1103_, data_stage_2__1102_, data_stage_2__1101_, data_stage_2__1100_, data_stage_2__1099_, data_stage_2__1098_, data_stage_2__1097_, data_stage_2__1096_, data_stage_2__1095_, data_stage_2__1094_, data_stage_2__1093_, data_stage_2__1092_, data_stage_2__1091_, data_stage_2__1090_, data_stage_2__1089_, data_stage_2__1088_, data_stage_2__1087_, data_stage_2__1086_, data_stage_2__1085_, data_stage_2__1084_, data_stage_2__1083_, data_stage_2__1082_, data_stage_2__1081_, data_stage_2__1080_, data_stage_2__1079_, data_stage_2__1078_, data_stage_2__1077_, data_stage_2__1076_, data_stage_2__1075_, data_stage_2__1074_, data_stage_2__1073_, data_stage_2__1072_, data_stage_2__1071_, data_stage_2__1070_, data_stage_2__1069_, data_stage_2__1068_, data_stage_2__1067_, data_stage_2__1066_, data_stage_2__1065_, data_stage_2__1064_, data_stage_2__1063_, data_stage_2__1062_, data_stage_2__1061_, data_stage_2__1060_, data_stage_2__1059_, data_stage_2__1058_, data_stage_2__1057_, data_stage_2__1056_, data_stage_2__1055_, data_stage_2__1054_, data_stage_2__1053_, data_stage_2__1052_, data_stage_2__1051_, data_stage_2__1050_, data_stage_2__1049_, data_stage_2__1048_, data_stage_2__1047_, data_stage_2__1046_, data_stage_2__1045_, data_stage_2__1044_, data_stage_2__1043_, data_stage_2__1042_, data_stage_2__1041_, data_stage_2__1040_, data_stage_2__1039_, data_stage_2__1038_, data_stage_2__1037_, data_stage_2__1036_, data_stage_2__1035_, data_stage_2__1034_, data_stage_2__1033_, data_stage_2__1032_, data_stage_2__1031_, data_stage_2__1030_, data_stage_2__1029_, data_stage_2__1028_, data_stage_2__1027_, data_stage_2__1026_, data_stage_2__1025_, data_stage_2__1024_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_3__swap_inst
  (
    .data_i({ data_stage_1__2047_, data_stage_1__2046_, data_stage_1__2045_, data_stage_1__2044_, data_stage_1__2043_, data_stage_1__2042_, data_stage_1__2041_, data_stage_1__2040_, data_stage_1__2039_, data_stage_1__2038_, data_stage_1__2037_, data_stage_1__2036_, data_stage_1__2035_, data_stage_1__2034_, data_stage_1__2033_, data_stage_1__2032_, data_stage_1__2031_, data_stage_1__2030_, data_stage_1__2029_, data_stage_1__2028_, data_stage_1__2027_, data_stage_1__2026_, data_stage_1__2025_, data_stage_1__2024_, data_stage_1__2023_, data_stage_1__2022_, data_stage_1__2021_, data_stage_1__2020_, data_stage_1__2019_, data_stage_1__2018_, data_stage_1__2017_, data_stage_1__2016_, data_stage_1__2015_, data_stage_1__2014_, data_stage_1__2013_, data_stage_1__2012_, data_stage_1__2011_, data_stage_1__2010_, data_stage_1__2009_, data_stage_1__2008_, data_stage_1__2007_, data_stage_1__2006_, data_stage_1__2005_, data_stage_1__2004_, data_stage_1__2003_, data_stage_1__2002_, data_stage_1__2001_, data_stage_1__2000_, data_stage_1__1999_, data_stage_1__1998_, data_stage_1__1997_, data_stage_1__1996_, data_stage_1__1995_, data_stage_1__1994_, data_stage_1__1993_, data_stage_1__1992_, data_stage_1__1991_, data_stage_1__1990_, data_stage_1__1989_, data_stage_1__1988_, data_stage_1__1987_, data_stage_1__1986_, data_stage_1__1985_, data_stage_1__1984_, data_stage_1__1983_, data_stage_1__1982_, data_stage_1__1981_, data_stage_1__1980_, data_stage_1__1979_, data_stage_1__1978_, data_stage_1__1977_, data_stage_1__1976_, data_stage_1__1975_, data_stage_1__1974_, data_stage_1__1973_, data_stage_1__1972_, data_stage_1__1971_, data_stage_1__1970_, data_stage_1__1969_, data_stage_1__1968_, data_stage_1__1967_, data_stage_1__1966_, data_stage_1__1965_, data_stage_1__1964_, data_stage_1__1963_, data_stage_1__1962_, data_stage_1__1961_, data_stage_1__1960_, data_stage_1__1959_, data_stage_1__1958_, data_stage_1__1957_, data_stage_1__1956_, data_stage_1__1955_, data_stage_1__1954_, data_stage_1__1953_, data_stage_1__1952_, data_stage_1__1951_, data_stage_1__1950_, data_stage_1__1949_, data_stage_1__1948_, data_stage_1__1947_, data_stage_1__1946_, data_stage_1__1945_, data_stage_1__1944_, data_stage_1__1943_, data_stage_1__1942_, data_stage_1__1941_, data_stage_1__1940_, data_stage_1__1939_, data_stage_1__1938_, data_stage_1__1937_, data_stage_1__1936_, data_stage_1__1935_, data_stage_1__1934_, data_stage_1__1933_, data_stage_1__1932_, data_stage_1__1931_, data_stage_1__1930_, data_stage_1__1929_, data_stage_1__1928_, data_stage_1__1927_, data_stage_1__1926_, data_stage_1__1925_, data_stage_1__1924_, data_stage_1__1923_, data_stage_1__1922_, data_stage_1__1921_, data_stage_1__1920_, data_stage_1__1919_, data_stage_1__1918_, data_stage_1__1917_, data_stage_1__1916_, data_stage_1__1915_, data_stage_1__1914_, data_stage_1__1913_, data_stage_1__1912_, data_stage_1__1911_, data_stage_1__1910_, data_stage_1__1909_, data_stage_1__1908_, data_stage_1__1907_, data_stage_1__1906_, data_stage_1__1905_, data_stage_1__1904_, data_stage_1__1903_, data_stage_1__1902_, data_stage_1__1901_, data_stage_1__1900_, data_stage_1__1899_, data_stage_1__1898_, data_stage_1__1897_, data_stage_1__1896_, data_stage_1__1895_, data_stage_1__1894_, data_stage_1__1893_, data_stage_1__1892_, data_stage_1__1891_, data_stage_1__1890_, data_stage_1__1889_, data_stage_1__1888_, data_stage_1__1887_, data_stage_1__1886_, data_stage_1__1885_, data_stage_1__1884_, data_stage_1__1883_, data_stage_1__1882_, data_stage_1__1881_, data_stage_1__1880_, data_stage_1__1879_, data_stage_1__1878_, data_stage_1__1877_, data_stage_1__1876_, data_stage_1__1875_, data_stage_1__1874_, data_stage_1__1873_, data_stage_1__1872_, data_stage_1__1871_, data_stage_1__1870_, data_stage_1__1869_, data_stage_1__1868_, data_stage_1__1867_, data_stage_1__1866_, data_stage_1__1865_, data_stage_1__1864_, data_stage_1__1863_, data_stage_1__1862_, data_stage_1__1861_, data_stage_1__1860_, data_stage_1__1859_, data_stage_1__1858_, data_stage_1__1857_, data_stage_1__1856_, data_stage_1__1855_, data_stage_1__1854_, data_stage_1__1853_, data_stage_1__1852_, data_stage_1__1851_, data_stage_1__1850_, data_stage_1__1849_, data_stage_1__1848_, data_stage_1__1847_, data_stage_1__1846_, data_stage_1__1845_, data_stage_1__1844_, data_stage_1__1843_, data_stage_1__1842_, data_stage_1__1841_, data_stage_1__1840_, data_stage_1__1839_, data_stage_1__1838_, data_stage_1__1837_, data_stage_1__1836_, data_stage_1__1835_, data_stage_1__1834_, data_stage_1__1833_, data_stage_1__1832_, data_stage_1__1831_, data_stage_1__1830_, data_stage_1__1829_, data_stage_1__1828_, data_stage_1__1827_, data_stage_1__1826_, data_stage_1__1825_, data_stage_1__1824_, data_stage_1__1823_, data_stage_1__1822_, data_stage_1__1821_, data_stage_1__1820_, data_stage_1__1819_, data_stage_1__1818_, data_stage_1__1817_, data_stage_1__1816_, data_stage_1__1815_, data_stage_1__1814_, data_stage_1__1813_, data_stage_1__1812_, data_stage_1__1811_, data_stage_1__1810_, data_stage_1__1809_, data_stage_1__1808_, data_stage_1__1807_, data_stage_1__1806_, data_stage_1__1805_, data_stage_1__1804_, data_stage_1__1803_, data_stage_1__1802_, data_stage_1__1801_, data_stage_1__1800_, data_stage_1__1799_, data_stage_1__1798_, data_stage_1__1797_, data_stage_1__1796_, data_stage_1__1795_, data_stage_1__1794_, data_stage_1__1793_, data_stage_1__1792_, data_stage_1__1791_, data_stage_1__1790_, data_stage_1__1789_, data_stage_1__1788_, data_stage_1__1787_, data_stage_1__1786_, data_stage_1__1785_, data_stage_1__1784_, data_stage_1__1783_, data_stage_1__1782_, data_stage_1__1781_, data_stage_1__1780_, data_stage_1__1779_, data_stage_1__1778_, data_stage_1__1777_, data_stage_1__1776_, data_stage_1__1775_, data_stage_1__1774_, data_stage_1__1773_, data_stage_1__1772_, data_stage_1__1771_, data_stage_1__1770_, data_stage_1__1769_, data_stage_1__1768_, data_stage_1__1767_, data_stage_1__1766_, data_stage_1__1765_, data_stage_1__1764_, data_stage_1__1763_, data_stage_1__1762_, data_stage_1__1761_, data_stage_1__1760_, data_stage_1__1759_, data_stage_1__1758_, data_stage_1__1757_, data_stage_1__1756_, data_stage_1__1755_, data_stage_1__1754_, data_stage_1__1753_, data_stage_1__1752_, data_stage_1__1751_, data_stage_1__1750_, data_stage_1__1749_, data_stage_1__1748_, data_stage_1__1747_, data_stage_1__1746_, data_stage_1__1745_, data_stage_1__1744_, data_stage_1__1743_, data_stage_1__1742_, data_stage_1__1741_, data_stage_1__1740_, data_stage_1__1739_, data_stage_1__1738_, data_stage_1__1737_, data_stage_1__1736_, data_stage_1__1735_, data_stage_1__1734_, data_stage_1__1733_, data_stage_1__1732_, data_stage_1__1731_, data_stage_1__1730_, data_stage_1__1729_, data_stage_1__1728_, data_stage_1__1727_, data_stage_1__1726_, data_stage_1__1725_, data_stage_1__1724_, data_stage_1__1723_, data_stage_1__1722_, data_stage_1__1721_, data_stage_1__1720_, data_stage_1__1719_, data_stage_1__1718_, data_stage_1__1717_, data_stage_1__1716_, data_stage_1__1715_, data_stage_1__1714_, data_stage_1__1713_, data_stage_1__1712_, data_stage_1__1711_, data_stage_1__1710_, data_stage_1__1709_, data_stage_1__1708_, data_stage_1__1707_, data_stage_1__1706_, data_stage_1__1705_, data_stage_1__1704_, data_stage_1__1703_, data_stage_1__1702_, data_stage_1__1701_, data_stage_1__1700_, data_stage_1__1699_, data_stage_1__1698_, data_stage_1__1697_, data_stage_1__1696_, data_stage_1__1695_, data_stage_1__1694_, data_stage_1__1693_, data_stage_1__1692_, data_stage_1__1691_, data_stage_1__1690_, data_stage_1__1689_, data_stage_1__1688_, data_stage_1__1687_, data_stage_1__1686_, data_stage_1__1685_, data_stage_1__1684_, data_stage_1__1683_, data_stage_1__1682_, data_stage_1__1681_, data_stage_1__1680_, data_stage_1__1679_, data_stage_1__1678_, data_stage_1__1677_, data_stage_1__1676_, data_stage_1__1675_, data_stage_1__1674_, data_stage_1__1673_, data_stage_1__1672_, data_stage_1__1671_, data_stage_1__1670_, data_stage_1__1669_, data_stage_1__1668_, data_stage_1__1667_, data_stage_1__1666_, data_stage_1__1665_, data_stage_1__1664_, data_stage_1__1663_, data_stage_1__1662_, data_stage_1__1661_, data_stage_1__1660_, data_stage_1__1659_, data_stage_1__1658_, data_stage_1__1657_, data_stage_1__1656_, data_stage_1__1655_, data_stage_1__1654_, data_stage_1__1653_, data_stage_1__1652_, data_stage_1__1651_, data_stage_1__1650_, data_stage_1__1649_, data_stage_1__1648_, data_stage_1__1647_, data_stage_1__1646_, data_stage_1__1645_, data_stage_1__1644_, data_stage_1__1643_, data_stage_1__1642_, data_stage_1__1641_, data_stage_1__1640_, data_stage_1__1639_, data_stage_1__1638_, data_stage_1__1637_, data_stage_1__1636_, data_stage_1__1635_, data_stage_1__1634_, data_stage_1__1633_, data_stage_1__1632_, data_stage_1__1631_, data_stage_1__1630_, data_stage_1__1629_, data_stage_1__1628_, data_stage_1__1627_, data_stage_1__1626_, data_stage_1__1625_, data_stage_1__1624_, data_stage_1__1623_, data_stage_1__1622_, data_stage_1__1621_, data_stage_1__1620_, data_stage_1__1619_, data_stage_1__1618_, data_stage_1__1617_, data_stage_1__1616_, data_stage_1__1615_, data_stage_1__1614_, data_stage_1__1613_, data_stage_1__1612_, data_stage_1__1611_, data_stage_1__1610_, data_stage_1__1609_, data_stage_1__1608_, data_stage_1__1607_, data_stage_1__1606_, data_stage_1__1605_, data_stage_1__1604_, data_stage_1__1603_, data_stage_1__1602_, data_stage_1__1601_, data_stage_1__1600_, data_stage_1__1599_, data_stage_1__1598_, data_stage_1__1597_, data_stage_1__1596_, data_stage_1__1595_, data_stage_1__1594_, data_stage_1__1593_, data_stage_1__1592_, data_stage_1__1591_, data_stage_1__1590_, data_stage_1__1589_, data_stage_1__1588_, data_stage_1__1587_, data_stage_1__1586_, data_stage_1__1585_, data_stage_1__1584_, data_stage_1__1583_, data_stage_1__1582_, data_stage_1__1581_, data_stage_1__1580_, data_stage_1__1579_, data_stage_1__1578_, data_stage_1__1577_, data_stage_1__1576_, data_stage_1__1575_, data_stage_1__1574_, data_stage_1__1573_, data_stage_1__1572_, data_stage_1__1571_, data_stage_1__1570_, data_stage_1__1569_, data_stage_1__1568_, data_stage_1__1567_, data_stage_1__1566_, data_stage_1__1565_, data_stage_1__1564_, data_stage_1__1563_, data_stage_1__1562_, data_stage_1__1561_, data_stage_1__1560_, data_stage_1__1559_, data_stage_1__1558_, data_stage_1__1557_, data_stage_1__1556_, data_stage_1__1555_, data_stage_1__1554_, data_stage_1__1553_, data_stage_1__1552_, data_stage_1__1551_, data_stage_1__1550_, data_stage_1__1549_, data_stage_1__1548_, data_stage_1__1547_, data_stage_1__1546_, data_stage_1__1545_, data_stage_1__1544_, data_stage_1__1543_, data_stage_1__1542_, data_stage_1__1541_, data_stage_1__1540_, data_stage_1__1539_, data_stage_1__1538_, data_stage_1__1537_, data_stage_1__1536_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__2047_, data_stage_2__2046_, data_stage_2__2045_, data_stage_2__2044_, data_stage_2__2043_, data_stage_2__2042_, data_stage_2__2041_, data_stage_2__2040_, data_stage_2__2039_, data_stage_2__2038_, data_stage_2__2037_, data_stage_2__2036_, data_stage_2__2035_, data_stage_2__2034_, data_stage_2__2033_, data_stage_2__2032_, data_stage_2__2031_, data_stage_2__2030_, data_stage_2__2029_, data_stage_2__2028_, data_stage_2__2027_, data_stage_2__2026_, data_stage_2__2025_, data_stage_2__2024_, data_stage_2__2023_, data_stage_2__2022_, data_stage_2__2021_, data_stage_2__2020_, data_stage_2__2019_, data_stage_2__2018_, data_stage_2__2017_, data_stage_2__2016_, data_stage_2__2015_, data_stage_2__2014_, data_stage_2__2013_, data_stage_2__2012_, data_stage_2__2011_, data_stage_2__2010_, data_stage_2__2009_, data_stage_2__2008_, data_stage_2__2007_, data_stage_2__2006_, data_stage_2__2005_, data_stage_2__2004_, data_stage_2__2003_, data_stage_2__2002_, data_stage_2__2001_, data_stage_2__2000_, data_stage_2__1999_, data_stage_2__1998_, data_stage_2__1997_, data_stage_2__1996_, data_stage_2__1995_, data_stage_2__1994_, data_stage_2__1993_, data_stage_2__1992_, data_stage_2__1991_, data_stage_2__1990_, data_stage_2__1989_, data_stage_2__1988_, data_stage_2__1987_, data_stage_2__1986_, data_stage_2__1985_, data_stage_2__1984_, data_stage_2__1983_, data_stage_2__1982_, data_stage_2__1981_, data_stage_2__1980_, data_stage_2__1979_, data_stage_2__1978_, data_stage_2__1977_, data_stage_2__1976_, data_stage_2__1975_, data_stage_2__1974_, data_stage_2__1973_, data_stage_2__1972_, data_stage_2__1971_, data_stage_2__1970_, data_stage_2__1969_, data_stage_2__1968_, data_stage_2__1967_, data_stage_2__1966_, data_stage_2__1965_, data_stage_2__1964_, data_stage_2__1963_, data_stage_2__1962_, data_stage_2__1961_, data_stage_2__1960_, data_stage_2__1959_, data_stage_2__1958_, data_stage_2__1957_, data_stage_2__1956_, data_stage_2__1955_, data_stage_2__1954_, data_stage_2__1953_, data_stage_2__1952_, data_stage_2__1951_, data_stage_2__1950_, data_stage_2__1949_, data_stage_2__1948_, data_stage_2__1947_, data_stage_2__1946_, data_stage_2__1945_, data_stage_2__1944_, data_stage_2__1943_, data_stage_2__1942_, data_stage_2__1941_, data_stage_2__1940_, data_stage_2__1939_, data_stage_2__1938_, data_stage_2__1937_, data_stage_2__1936_, data_stage_2__1935_, data_stage_2__1934_, data_stage_2__1933_, data_stage_2__1932_, data_stage_2__1931_, data_stage_2__1930_, data_stage_2__1929_, data_stage_2__1928_, data_stage_2__1927_, data_stage_2__1926_, data_stage_2__1925_, data_stage_2__1924_, data_stage_2__1923_, data_stage_2__1922_, data_stage_2__1921_, data_stage_2__1920_, data_stage_2__1919_, data_stage_2__1918_, data_stage_2__1917_, data_stage_2__1916_, data_stage_2__1915_, data_stage_2__1914_, data_stage_2__1913_, data_stage_2__1912_, data_stage_2__1911_, data_stage_2__1910_, data_stage_2__1909_, data_stage_2__1908_, data_stage_2__1907_, data_stage_2__1906_, data_stage_2__1905_, data_stage_2__1904_, data_stage_2__1903_, data_stage_2__1902_, data_stage_2__1901_, data_stage_2__1900_, data_stage_2__1899_, data_stage_2__1898_, data_stage_2__1897_, data_stage_2__1896_, data_stage_2__1895_, data_stage_2__1894_, data_stage_2__1893_, data_stage_2__1892_, data_stage_2__1891_, data_stage_2__1890_, data_stage_2__1889_, data_stage_2__1888_, data_stage_2__1887_, data_stage_2__1886_, data_stage_2__1885_, data_stage_2__1884_, data_stage_2__1883_, data_stage_2__1882_, data_stage_2__1881_, data_stage_2__1880_, data_stage_2__1879_, data_stage_2__1878_, data_stage_2__1877_, data_stage_2__1876_, data_stage_2__1875_, data_stage_2__1874_, data_stage_2__1873_, data_stage_2__1872_, data_stage_2__1871_, data_stage_2__1870_, data_stage_2__1869_, data_stage_2__1868_, data_stage_2__1867_, data_stage_2__1866_, data_stage_2__1865_, data_stage_2__1864_, data_stage_2__1863_, data_stage_2__1862_, data_stage_2__1861_, data_stage_2__1860_, data_stage_2__1859_, data_stage_2__1858_, data_stage_2__1857_, data_stage_2__1856_, data_stage_2__1855_, data_stage_2__1854_, data_stage_2__1853_, data_stage_2__1852_, data_stage_2__1851_, data_stage_2__1850_, data_stage_2__1849_, data_stage_2__1848_, data_stage_2__1847_, data_stage_2__1846_, data_stage_2__1845_, data_stage_2__1844_, data_stage_2__1843_, data_stage_2__1842_, data_stage_2__1841_, data_stage_2__1840_, data_stage_2__1839_, data_stage_2__1838_, data_stage_2__1837_, data_stage_2__1836_, data_stage_2__1835_, data_stage_2__1834_, data_stage_2__1833_, data_stage_2__1832_, data_stage_2__1831_, data_stage_2__1830_, data_stage_2__1829_, data_stage_2__1828_, data_stage_2__1827_, data_stage_2__1826_, data_stage_2__1825_, data_stage_2__1824_, data_stage_2__1823_, data_stage_2__1822_, data_stage_2__1821_, data_stage_2__1820_, data_stage_2__1819_, data_stage_2__1818_, data_stage_2__1817_, data_stage_2__1816_, data_stage_2__1815_, data_stage_2__1814_, data_stage_2__1813_, data_stage_2__1812_, data_stage_2__1811_, data_stage_2__1810_, data_stage_2__1809_, data_stage_2__1808_, data_stage_2__1807_, data_stage_2__1806_, data_stage_2__1805_, data_stage_2__1804_, data_stage_2__1803_, data_stage_2__1802_, data_stage_2__1801_, data_stage_2__1800_, data_stage_2__1799_, data_stage_2__1798_, data_stage_2__1797_, data_stage_2__1796_, data_stage_2__1795_, data_stage_2__1794_, data_stage_2__1793_, data_stage_2__1792_, data_stage_2__1791_, data_stage_2__1790_, data_stage_2__1789_, data_stage_2__1788_, data_stage_2__1787_, data_stage_2__1786_, data_stage_2__1785_, data_stage_2__1784_, data_stage_2__1783_, data_stage_2__1782_, data_stage_2__1781_, data_stage_2__1780_, data_stage_2__1779_, data_stage_2__1778_, data_stage_2__1777_, data_stage_2__1776_, data_stage_2__1775_, data_stage_2__1774_, data_stage_2__1773_, data_stage_2__1772_, data_stage_2__1771_, data_stage_2__1770_, data_stage_2__1769_, data_stage_2__1768_, data_stage_2__1767_, data_stage_2__1766_, data_stage_2__1765_, data_stage_2__1764_, data_stage_2__1763_, data_stage_2__1762_, data_stage_2__1761_, data_stage_2__1760_, data_stage_2__1759_, data_stage_2__1758_, data_stage_2__1757_, data_stage_2__1756_, data_stage_2__1755_, data_stage_2__1754_, data_stage_2__1753_, data_stage_2__1752_, data_stage_2__1751_, data_stage_2__1750_, data_stage_2__1749_, data_stage_2__1748_, data_stage_2__1747_, data_stage_2__1746_, data_stage_2__1745_, data_stage_2__1744_, data_stage_2__1743_, data_stage_2__1742_, data_stage_2__1741_, data_stage_2__1740_, data_stage_2__1739_, data_stage_2__1738_, data_stage_2__1737_, data_stage_2__1736_, data_stage_2__1735_, data_stage_2__1734_, data_stage_2__1733_, data_stage_2__1732_, data_stage_2__1731_, data_stage_2__1730_, data_stage_2__1729_, data_stage_2__1728_, data_stage_2__1727_, data_stage_2__1726_, data_stage_2__1725_, data_stage_2__1724_, data_stage_2__1723_, data_stage_2__1722_, data_stage_2__1721_, data_stage_2__1720_, data_stage_2__1719_, data_stage_2__1718_, data_stage_2__1717_, data_stage_2__1716_, data_stage_2__1715_, data_stage_2__1714_, data_stage_2__1713_, data_stage_2__1712_, data_stage_2__1711_, data_stage_2__1710_, data_stage_2__1709_, data_stage_2__1708_, data_stage_2__1707_, data_stage_2__1706_, data_stage_2__1705_, data_stage_2__1704_, data_stage_2__1703_, data_stage_2__1702_, data_stage_2__1701_, data_stage_2__1700_, data_stage_2__1699_, data_stage_2__1698_, data_stage_2__1697_, data_stage_2__1696_, data_stage_2__1695_, data_stage_2__1694_, data_stage_2__1693_, data_stage_2__1692_, data_stage_2__1691_, data_stage_2__1690_, data_stage_2__1689_, data_stage_2__1688_, data_stage_2__1687_, data_stage_2__1686_, data_stage_2__1685_, data_stage_2__1684_, data_stage_2__1683_, data_stage_2__1682_, data_stage_2__1681_, data_stage_2__1680_, data_stage_2__1679_, data_stage_2__1678_, data_stage_2__1677_, data_stage_2__1676_, data_stage_2__1675_, data_stage_2__1674_, data_stage_2__1673_, data_stage_2__1672_, data_stage_2__1671_, data_stage_2__1670_, data_stage_2__1669_, data_stage_2__1668_, data_stage_2__1667_, data_stage_2__1666_, data_stage_2__1665_, data_stage_2__1664_, data_stage_2__1663_, data_stage_2__1662_, data_stage_2__1661_, data_stage_2__1660_, data_stage_2__1659_, data_stage_2__1658_, data_stage_2__1657_, data_stage_2__1656_, data_stage_2__1655_, data_stage_2__1654_, data_stage_2__1653_, data_stage_2__1652_, data_stage_2__1651_, data_stage_2__1650_, data_stage_2__1649_, data_stage_2__1648_, data_stage_2__1647_, data_stage_2__1646_, data_stage_2__1645_, data_stage_2__1644_, data_stage_2__1643_, data_stage_2__1642_, data_stage_2__1641_, data_stage_2__1640_, data_stage_2__1639_, data_stage_2__1638_, data_stage_2__1637_, data_stage_2__1636_, data_stage_2__1635_, data_stage_2__1634_, data_stage_2__1633_, data_stage_2__1632_, data_stage_2__1631_, data_stage_2__1630_, data_stage_2__1629_, data_stage_2__1628_, data_stage_2__1627_, data_stage_2__1626_, data_stage_2__1625_, data_stage_2__1624_, data_stage_2__1623_, data_stage_2__1622_, data_stage_2__1621_, data_stage_2__1620_, data_stage_2__1619_, data_stage_2__1618_, data_stage_2__1617_, data_stage_2__1616_, data_stage_2__1615_, data_stage_2__1614_, data_stage_2__1613_, data_stage_2__1612_, data_stage_2__1611_, data_stage_2__1610_, data_stage_2__1609_, data_stage_2__1608_, data_stage_2__1607_, data_stage_2__1606_, data_stage_2__1605_, data_stage_2__1604_, data_stage_2__1603_, data_stage_2__1602_, data_stage_2__1601_, data_stage_2__1600_, data_stage_2__1599_, data_stage_2__1598_, data_stage_2__1597_, data_stage_2__1596_, data_stage_2__1595_, data_stage_2__1594_, data_stage_2__1593_, data_stage_2__1592_, data_stage_2__1591_, data_stage_2__1590_, data_stage_2__1589_, data_stage_2__1588_, data_stage_2__1587_, data_stage_2__1586_, data_stage_2__1585_, data_stage_2__1584_, data_stage_2__1583_, data_stage_2__1582_, data_stage_2__1581_, data_stage_2__1580_, data_stage_2__1579_, data_stage_2__1578_, data_stage_2__1577_, data_stage_2__1576_, data_stage_2__1575_, data_stage_2__1574_, data_stage_2__1573_, data_stage_2__1572_, data_stage_2__1571_, data_stage_2__1570_, data_stage_2__1569_, data_stage_2__1568_, data_stage_2__1567_, data_stage_2__1566_, data_stage_2__1565_, data_stage_2__1564_, data_stage_2__1563_, data_stage_2__1562_, data_stage_2__1561_, data_stage_2__1560_, data_stage_2__1559_, data_stage_2__1558_, data_stage_2__1557_, data_stage_2__1556_, data_stage_2__1555_, data_stage_2__1554_, data_stage_2__1553_, data_stage_2__1552_, data_stage_2__1551_, data_stage_2__1550_, data_stage_2__1549_, data_stage_2__1548_, data_stage_2__1547_, data_stage_2__1546_, data_stage_2__1545_, data_stage_2__1544_, data_stage_2__1543_, data_stage_2__1542_, data_stage_2__1541_, data_stage_2__1540_, data_stage_2__1539_, data_stage_2__1538_, data_stage_2__1537_, data_stage_2__1536_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_4__swap_inst
  (
    .data_i({ data_stage_1__2559_, data_stage_1__2558_, data_stage_1__2557_, data_stage_1__2556_, data_stage_1__2555_, data_stage_1__2554_, data_stage_1__2553_, data_stage_1__2552_, data_stage_1__2551_, data_stage_1__2550_, data_stage_1__2549_, data_stage_1__2548_, data_stage_1__2547_, data_stage_1__2546_, data_stage_1__2545_, data_stage_1__2544_, data_stage_1__2543_, data_stage_1__2542_, data_stage_1__2541_, data_stage_1__2540_, data_stage_1__2539_, data_stage_1__2538_, data_stage_1__2537_, data_stage_1__2536_, data_stage_1__2535_, data_stage_1__2534_, data_stage_1__2533_, data_stage_1__2532_, data_stage_1__2531_, data_stage_1__2530_, data_stage_1__2529_, data_stage_1__2528_, data_stage_1__2527_, data_stage_1__2526_, data_stage_1__2525_, data_stage_1__2524_, data_stage_1__2523_, data_stage_1__2522_, data_stage_1__2521_, data_stage_1__2520_, data_stage_1__2519_, data_stage_1__2518_, data_stage_1__2517_, data_stage_1__2516_, data_stage_1__2515_, data_stage_1__2514_, data_stage_1__2513_, data_stage_1__2512_, data_stage_1__2511_, data_stage_1__2510_, data_stage_1__2509_, data_stage_1__2508_, data_stage_1__2507_, data_stage_1__2506_, data_stage_1__2505_, data_stage_1__2504_, data_stage_1__2503_, data_stage_1__2502_, data_stage_1__2501_, data_stage_1__2500_, data_stage_1__2499_, data_stage_1__2498_, data_stage_1__2497_, data_stage_1__2496_, data_stage_1__2495_, data_stage_1__2494_, data_stage_1__2493_, data_stage_1__2492_, data_stage_1__2491_, data_stage_1__2490_, data_stage_1__2489_, data_stage_1__2488_, data_stage_1__2487_, data_stage_1__2486_, data_stage_1__2485_, data_stage_1__2484_, data_stage_1__2483_, data_stage_1__2482_, data_stage_1__2481_, data_stage_1__2480_, data_stage_1__2479_, data_stage_1__2478_, data_stage_1__2477_, data_stage_1__2476_, data_stage_1__2475_, data_stage_1__2474_, data_stage_1__2473_, data_stage_1__2472_, data_stage_1__2471_, data_stage_1__2470_, data_stage_1__2469_, data_stage_1__2468_, data_stage_1__2467_, data_stage_1__2466_, data_stage_1__2465_, data_stage_1__2464_, data_stage_1__2463_, data_stage_1__2462_, data_stage_1__2461_, data_stage_1__2460_, data_stage_1__2459_, data_stage_1__2458_, data_stage_1__2457_, data_stage_1__2456_, data_stage_1__2455_, data_stage_1__2454_, data_stage_1__2453_, data_stage_1__2452_, data_stage_1__2451_, data_stage_1__2450_, data_stage_1__2449_, data_stage_1__2448_, data_stage_1__2447_, data_stage_1__2446_, data_stage_1__2445_, data_stage_1__2444_, data_stage_1__2443_, data_stage_1__2442_, data_stage_1__2441_, data_stage_1__2440_, data_stage_1__2439_, data_stage_1__2438_, data_stage_1__2437_, data_stage_1__2436_, data_stage_1__2435_, data_stage_1__2434_, data_stage_1__2433_, data_stage_1__2432_, data_stage_1__2431_, data_stage_1__2430_, data_stage_1__2429_, data_stage_1__2428_, data_stage_1__2427_, data_stage_1__2426_, data_stage_1__2425_, data_stage_1__2424_, data_stage_1__2423_, data_stage_1__2422_, data_stage_1__2421_, data_stage_1__2420_, data_stage_1__2419_, data_stage_1__2418_, data_stage_1__2417_, data_stage_1__2416_, data_stage_1__2415_, data_stage_1__2414_, data_stage_1__2413_, data_stage_1__2412_, data_stage_1__2411_, data_stage_1__2410_, data_stage_1__2409_, data_stage_1__2408_, data_stage_1__2407_, data_stage_1__2406_, data_stage_1__2405_, data_stage_1__2404_, data_stage_1__2403_, data_stage_1__2402_, data_stage_1__2401_, data_stage_1__2400_, data_stage_1__2399_, data_stage_1__2398_, data_stage_1__2397_, data_stage_1__2396_, data_stage_1__2395_, data_stage_1__2394_, data_stage_1__2393_, data_stage_1__2392_, data_stage_1__2391_, data_stage_1__2390_, data_stage_1__2389_, data_stage_1__2388_, data_stage_1__2387_, data_stage_1__2386_, data_stage_1__2385_, data_stage_1__2384_, data_stage_1__2383_, data_stage_1__2382_, data_stage_1__2381_, data_stage_1__2380_, data_stage_1__2379_, data_stage_1__2378_, data_stage_1__2377_, data_stage_1__2376_, data_stage_1__2375_, data_stage_1__2374_, data_stage_1__2373_, data_stage_1__2372_, data_stage_1__2371_, data_stage_1__2370_, data_stage_1__2369_, data_stage_1__2368_, data_stage_1__2367_, data_stage_1__2366_, data_stage_1__2365_, data_stage_1__2364_, data_stage_1__2363_, data_stage_1__2362_, data_stage_1__2361_, data_stage_1__2360_, data_stage_1__2359_, data_stage_1__2358_, data_stage_1__2357_, data_stage_1__2356_, data_stage_1__2355_, data_stage_1__2354_, data_stage_1__2353_, data_stage_1__2352_, data_stage_1__2351_, data_stage_1__2350_, data_stage_1__2349_, data_stage_1__2348_, data_stage_1__2347_, data_stage_1__2346_, data_stage_1__2345_, data_stage_1__2344_, data_stage_1__2343_, data_stage_1__2342_, data_stage_1__2341_, data_stage_1__2340_, data_stage_1__2339_, data_stage_1__2338_, data_stage_1__2337_, data_stage_1__2336_, data_stage_1__2335_, data_stage_1__2334_, data_stage_1__2333_, data_stage_1__2332_, data_stage_1__2331_, data_stage_1__2330_, data_stage_1__2329_, data_stage_1__2328_, data_stage_1__2327_, data_stage_1__2326_, data_stage_1__2325_, data_stage_1__2324_, data_stage_1__2323_, data_stage_1__2322_, data_stage_1__2321_, data_stage_1__2320_, data_stage_1__2319_, data_stage_1__2318_, data_stage_1__2317_, data_stage_1__2316_, data_stage_1__2315_, data_stage_1__2314_, data_stage_1__2313_, data_stage_1__2312_, data_stage_1__2311_, data_stage_1__2310_, data_stage_1__2309_, data_stage_1__2308_, data_stage_1__2307_, data_stage_1__2306_, data_stage_1__2305_, data_stage_1__2304_, data_stage_1__2303_, data_stage_1__2302_, data_stage_1__2301_, data_stage_1__2300_, data_stage_1__2299_, data_stage_1__2298_, data_stage_1__2297_, data_stage_1__2296_, data_stage_1__2295_, data_stage_1__2294_, data_stage_1__2293_, data_stage_1__2292_, data_stage_1__2291_, data_stage_1__2290_, data_stage_1__2289_, data_stage_1__2288_, data_stage_1__2287_, data_stage_1__2286_, data_stage_1__2285_, data_stage_1__2284_, data_stage_1__2283_, data_stage_1__2282_, data_stage_1__2281_, data_stage_1__2280_, data_stage_1__2279_, data_stage_1__2278_, data_stage_1__2277_, data_stage_1__2276_, data_stage_1__2275_, data_stage_1__2274_, data_stage_1__2273_, data_stage_1__2272_, data_stage_1__2271_, data_stage_1__2270_, data_stage_1__2269_, data_stage_1__2268_, data_stage_1__2267_, data_stage_1__2266_, data_stage_1__2265_, data_stage_1__2264_, data_stage_1__2263_, data_stage_1__2262_, data_stage_1__2261_, data_stage_1__2260_, data_stage_1__2259_, data_stage_1__2258_, data_stage_1__2257_, data_stage_1__2256_, data_stage_1__2255_, data_stage_1__2254_, data_stage_1__2253_, data_stage_1__2252_, data_stage_1__2251_, data_stage_1__2250_, data_stage_1__2249_, data_stage_1__2248_, data_stage_1__2247_, data_stage_1__2246_, data_stage_1__2245_, data_stage_1__2244_, data_stage_1__2243_, data_stage_1__2242_, data_stage_1__2241_, data_stage_1__2240_, data_stage_1__2239_, data_stage_1__2238_, data_stage_1__2237_, data_stage_1__2236_, data_stage_1__2235_, data_stage_1__2234_, data_stage_1__2233_, data_stage_1__2232_, data_stage_1__2231_, data_stage_1__2230_, data_stage_1__2229_, data_stage_1__2228_, data_stage_1__2227_, data_stage_1__2226_, data_stage_1__2225_, data_stage_1__2224_, data_stage_1__2223_, data_stage_1__2222_, data_stage_1__2221_, data_stage_1__2220_, data_stage_1__2219_, data_stage_1__2218_, data_stage_1__2217_, data_stage_1__2216_, data_stage_1__2215_, data_stage_1__2214_, data_stage_1__2213_, data_stage_1__2212_, data_stage_1__2211_, data_stage_1__2210_, data_stage_1__2209_, data_stage_1__2208_, data_stage_1__2207_, data_stage_1__2206_, data_stage_1__2205_, data_stage_1__2204_, data_stage_1__2203_, data_stage_1__2202_, data_stage_1__2201_, data_stage_1__2200_, data_stage_1__2199_, data_stage_1__2198_, data_stage_1__2197_, data_stage_1__2196_, data_stage_1__2195_, data_stage_1__2194_, data_stage_1__2193_, data_stage_1__2192_, data_stage_1__2191_, data_stage_1__2190_, data_stage_1__2189_, data_stage_1__2188_, data_stage_1__2187_, data_stage_1__2186_, data_stage_1__2185_, data_stage_1__2184_, data_stage_1__2183_, data_stage_1__2182_, data_stage_1__2181_, data_stage_1__2180_, data_stage_1__2179_, data_stage_1__2178_, data_stage_1__2177_, data_stage_1__2176_, data_stage_1__2175_, data_stage_1__2174_, data_stage_1__2173_, data_stage_1__2172_, data_stage_1__2171_, data_stage_1__2170_, data_stage_1__2169_, data_stage_1__2168_, data_stage_1__2167_, data_stage_1__2166_, data_stage_1__2165_, data_stage_1__2164_, data_stage_1__2163_, data_stage_1__2162_, data_stage_1__2161_, data_stage_1__2160_, data_stage_1__2159_, data_stage_1__2158_, data_stage_1__2157_, data_stage_1__2156_, data_stage_1__2155_, data_stage_1__2154_, data_stage_1__2153_, data_stage_1__2152_, data_stage_1__2151_, data_stage_1__2150_, data_stage_1__2149_, data_stage_1__2148_, data_stage_1__2147_, data_stage_1__2146_, data_stage_1__2145_, data_stage_1__2144_, data_stage_1__2143_, data_stage_1__2142_, data_stage_1__2141_, data_stage_1__2140_, data_stage_1__2139_, data_stage_1__2138_, data_stage_1__2137_, data_stage_1__2136_, data_stage_1__2135_, data_stage_1__2134_, data_stage_1__2133_, data_stage_1__2132_, data_stage_1__2131_, data_stage_1__2130_, data_stage_1__2129_, data_stage_1__2128_, data_stage_1__2127_, data_stage_1__2126_, data_stage_1__2125_, data_stage_1__2124_, data_stage_1__2123_, data_stage_1__2122_, data_stage_1__2121_, data_stage_1__2120_, data_stage_1__2119_, data_stage_1__2118_, data_stage_1__2117_, data_stage_1__2116_, data_stage_1__2115_, data_stage_1__2114_, data_stage_1__2113_, data_stage_1__2112_, data_stage_1__2111_, data_stage_1__2110_, data_stage_1__2109_, data_stage_1__2108_, data_stage_1__2107_, data_stage_1__2106_, data_stage_1__2105_, data_stage_1__2104_, data_stage_1__2103_, data_stage_1__2102_, data_stage_1__2101_, data_stage_1__2100_, data_stage_1__2099_, data_stage_1__2098_, data_stage_1__2097_, data_stage_1__2096_, data_stage_1__2095_, data_stage_1__2094_, data_stage_1__2093_, data_stage_1__2092_, data_stage_1__2091_, data_stage_1__2090_, data_stage_1__2089_, data_stage_1__2088_, data_stage_1__2087_, data_stage_1__2086_, data_stage_1__2085_, data_stage_1__2084_, data_stage_1__2083_, data_stage_1__2082_, data_stage_1__2081_, data_stage_1__2080_, data_stage_1__2079_, data_stage_1__2078_, data_stage_1__2077_, data_stage_1__2076_, data_stage_1__2075_, data_stage_1__2074_, data_stage_1__2073_, data_stage_1__2072_, data_stage_1__2071_, data_stage_1__2070_, data_stage_1__2069_, data_stage_1__2068_, data_stage_1__2067_, data_stage_1__2066_, data_stage_1__2065_, data_stage_1__2064_, data_stage_1__2063_, data_stage_1__2062_, data_stage_1__2061_, data_stage_1__2060_, data_stage_1__2059_, data_stage_1__2058_, data_stage_1__2057_, data_stage_1__2056_, data_stage_1__2055_, data_stage_1__2054_, data_stage_1__2053_, data_stage_1__2052_, data_stage_1__2051_, data_stage_1__2050_, data_stage_1__2049_, data_stage_1__2048_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__2559_, data_stage_2__2558_, data_stage_2__2557_, data_stage_2__2556_, data_stage_2__2555_, data_stage_2__2554_, data_stage_2__2553_, data_stage_2__2552_, data_stage_2__2551_, data_stage_2__2550_, data_stage_2__2549_, data_stage_2__2548_, data_stage_2__2547_, data_stage_2__2546_, data_stage_2__2545_, data_stage_2__2544_, data_stage_2__2543_, data_stage_2__2542_, data_stage_2__2541_, data_stage_2__2540_, data_stage_2__2539_, data_stage_2__2538_, data_stage_2__2537_, data_stage_2__2536_, data_stage_2__2535_, data_stage_2__2534_, data_stage_2__2533_, data_stage_2__2532_, data_stage_2__2531_, data_stage_2__2530_, data_stage_2__2529_, data_stage_2__2528_, data_stage_2__2527_, data_stage_2__2526_, data_stage_2__2525_, data_stage_2__2524_, data_stage_2__2523_, data_stage_2__2522_, data_stage_2__2521_, data_stage_2__2520_, data_stage_2__2519_, data_stage_2__2518_, data_stage_2__2517_, data_stage_2__2516_, data_stage_2__2515_, data_stage_2__2514_, data_stage_2__2513_, data_stage_2__2512_, data_stage_2__2511_, data_stage_2__2510_, data_stage_2__2509_, data_stage_2__2508_, data_stage_2__2507_, data_stage_2__2506_, data_stage_2__2505_, data_stage_2__2504_, data_stage_2__2503_, data_stage_2__2502_, data_stage_2__2501_, data_stage_2__2500_, data_stage_2__2499_, data_stage_2__2498_, data_stage_2__2497_, data_stage_2__2496_, data_stage_2__2495_, data_stage_2__2494_, data_stage_2__2493_, data_stage_2__2492_, data_stage_2__2491_, data_stage_2__2490_, data_stage_2__2489_, data_stage_2__2488_, data_stage_2__2487_, data_stage_2__2486_, data_stage_2__2485_, data_stage_2__2484_, data_stage_2__2483_, data_stage_2__2482_, data_stage_2__2481_, data_stage_2__2480_, data_stage_2__2479_, data_stage_2__2478_, data_stage_2__2477_, data_stage_2__2476_, data_stage_2__2475_, data_stage_2__2474_, data_stage_2__2473_, data_stage_2__2472_, data_stage_2__2471_, data_stage_2__2470_, data_stage_2__2469_, data_stage_2__2468_, data_stage_2__2467_, data_stage_2__2466_, data_stage_2__2465_, data_stage_2__2464_, data_stage_2__2463_, data_stage_2__2462_, data_stage_2__2461_, data_stage_2__2460_, data_stage_2__2459_, data_stage_2__2458_, data_stage_2__2457_, data_stage_2__2456_, data_stage_2__2455_, data_stage_2__2454_, data_stage_2__2453_, data_stage_2__2452_, data_stage_2__2451_, data_stage_2__2450_, data_stage_2__2449_, data_stage_2__2448_, data_stage_2__2447_, data_stage_2__2446_, data_stage_2__2445_, data_stage_2__2444_, data_stage_2__2443_, data_stage_2__2442_, data_stage_2__2441_, data_stage_2__2440_, data_stage_2__2439_, data_stage_2__2438_, data_stage_2__2437_, data_stage_2__2436_, data_stage_2__2435_, data_stage_2__2434_, data_stage_2__2433_, data_stage_2__2432_, data_stage_2__2431_, data_stage_2__2430_, data_stage_2__2429_, data_stage_2__2428_, data_stage_2__2427_, data_stage_2__2426_, data_stage_2__2425_, data_stage_2__2424_, data_stage_2__2423_, data_stage_2__2422_, data_stage_2__2421_, data_stage_2__2420_, data_stage_2__2419_, data_stage_2__2418_, data_stage_2__2417_, data_stage_2__2416_, data_stage_2__2415_, data_stage_2__2414_, data_stage_2__2413_, data_stage_2__2412_, data_stage_2__2411_, data_stage_2__2410_, data_stage_2__2409_, data_stage_2__2408_, data_stage_2__2407_, data_stage_2__2406_, data_stage_2__2405_, data_stage_2__2404_, data_stage_2__2403_, data_stage_2__2402_, data_stage_2__2401_, data_stage_2__2400_, data_stage_2__2399_, data_stage_2__2398_, data_stage_2__2397_, data_stage_2__2396_, data_stage_2__2395_, data_stage_2__2394_, data_stage_2__2393_, data_stage_2__2392_, data_stage_2__2391_, data_stage_2__2390_, data_stage_2__2389_, data_stage_2__2388_, data_stage_2__2387_, data_stage_2__2386_, data_stage_2__2385_, data_stage_2__2384_, data_stage_2__2383_, data_stage_2__2382_, data_stage_2__2381_, data_stage_2__2380_, data_stage_2__2379_, data_stage_2__2378_, data_stage_2__2377_, data_stage_2__2376_, data_stage_2__2375_, data_stage_2__2374_, data_stage_2__2373_, data_stage_2__2372_, data_stage_2__2371_, data_stage_2__2370_, data_stage_2__2369_, data_stage_2__2368_, data_stage_2__2367_, data_stage_2__2366_, data_stage_2__2365_, data_stage_2__2364_, data_stage_2__2363_, data_stage_2__2362_, data_stage_2__2361_, data_stage_2__2360_, data_stage_2__2359_, data_stage_2__2358_, data_stage_2__2357_, data_stage_2__2356_, data_stage_2__2355_, data_stage_2__2354_, data_stage_2__2353_, data_stage_2__2352_, data_stage_2__2351_, data_stage_2__2350_, data_stage_2__2349_, data_stage_2__2348_, data_stage_2__2347_, data_stage_2__2346_, data_stage_2__2345_, data_stage_2__2344_, data_stage_2__2343_, data_stage_2__2342_, data_stage_2__2341_, data_stage_2__2340_, data_stage_2__2339_, data_stage_2__2338_, data_stage_2__2337_, data_stage_2__2336_, data_stage_2__2335_, data_stage_2__2334_, data_stage_2__2333_, data_stage_2__2332_, data_stage_2__2331_, data_stage_2__2330_, data_stage_2__2329_, data_stage_2__2328_, data_stage_2__2327_, data_stage_2__2326_, data_stage_2__2325_, data_stage_2__2324_, data_stage_2__2323_, data_stage_2__2322_, data_stage_2__2321_, data_stage_2__2320_, data_stage_2__2319_, data_stage_2__2318_, data_stage_2__2317_, data_stage_2__2316_, data_stage_2__2315_, data_stage_2__2314_, data_stage_2__2313_, data_stage_2__2312_, data_stage_2__2311_, data_stage_2__2310_, data_stage_2__2309_, data_stage_2__2308_, data_stage_2__2307_, data_stage_2__2306_, data_stage_2__2305_, data_stage_2__2304_, data_stage_2__2303_, data_stage_2__2302_, data_stage_2__2301_, data_stage_2__2300_, data_stage_2__2299_, data_stage_2__2298_, data_stage_2__2297_, data_stage_2__2296_, data_stage_2__2295_, data_stage_2__2294_, data_stage_2__2293_, data_stage_2__2292_, data_stage_2__2291_, data_stage_2__2290_, data_stage_2__2289_, data_stage_2__2288_, data_stage_2__2287_, data_stage_2__2286_, data_stage_2__2285_, data_stage_2__2284_, data_stage_2__2283_, data_stage_2__2282_, data_stage_2__2281_, data_stage_2__2280_, data_stage_2__2279_, data_stage_2__2278_, data_stage_2__2277_, data_stage_2__2276_, data_stage_2__2275_, data_stage_2__2274_, data_stage_2__2273_, data_stage_2__2272_, data_stage_2__2271_, data_stage_2__2270_, data_stage_2__2269_, data_stage_2__2268_, data_stage_2__2267_, data_stage_2__2266_, data_stage_2__2265_, data_stage_2__2264_, data_stage_2__2263_, data_stage_2__2262_, data_stage_2__2261_, data_stage_2__2260_, data_stage_2__2259_, data_stage_2__2258_, data_stage_2__2257_, data_stage_2__2256_, data_stage_2__2255_, data_stage_2__2254_, data_stage_2__2253_, data_stage_2__2252_, data_stage_2__2251_, data_stage_2__2250_, data_stage_2__2249_, data_stage_2__2248_, data_stage_2__2247_, data_stage_2__2246_, data_stage_2__2245_, data_stage_2__2244_, data_stage_2__2243_, data_stage_2__2242_, data_stage_2__2241_, data_stage_2__2240_, data_stage_2__2239_, data_stage_2__2238_, data_stage_2__2237_, data_stage_2__2236_, data_stage_2__2235_, data_stage_2__2234_, data_stage_2__2233_, data_stage_2__2232_, data_stage_2__2231_, data_stage_2__2230_, data_stage_2__2229_, data_stage_2__2228_, data_stage_2__2227_, data_stage_2__2226_, data_stage_2__2225_, data_stage_2__2224_, data_stage_2__2223_, data_stage_2__2222_, data_stage_2__2221_, data_stage_2__2220_, data_stage_2__2219_, data_stage_2__2218_, data_stage_2__2217_, data_stage_2__2216_, data_stage_2__2215_, data_stage_2__2214_, data_stage_2__2213_, data_stage_2__2212_, data_stage_2__2211_, data_stage_2__2210_, data_stage_2__2209_, data_stage_2__2208_, data_stage_2__2207_, data_stage_2__2206_, data_stage_2__2205_, data_stage_2__2204_, data_stage_2__2203_, data_stage_2__2202_, data_stage_2__2201_, data_stage_2__2200_, data_stage_2__2199_, data_stage_2__2198_, data_stage_2__2197_, data_stage_2__2196_, data_stage_2__2195_, data_stage_2__2194_, data_stage_2__2193_, data_stage_2__2192_, data_stage_2__2191_, data_stage_2__2190_, data_stage_2__2189_, data_stage_2__2188_, data_stage_2__2187_, data_stage_2__2186_, data_stage_2__2185_, data_stage_2__2184_, data_stage_2__2183_, data_stage_2__2182_, data_stage_2__2181_, data_stage_2__2180_, data_stage_2__2179_, data_stage_2__2178_, data_stage_2__2177_, data_stage_2__2176_, data_stage_2__2175_, data_stage_2__2174_, data_stage_2__2173_, data_stage_2__2172_, data_stage_2__2171_, data_stage_2__2170_, data_stage_2__2169_, data_stage_2__2168_, data_stage_2__2167_, data_stage_2__2166_, data_stage_2__2165_, data_stage_2__2164_, data_stage_2__2163_, data_stage_2__2162_, data_stage_2__2161_, data_stage_2__2160_, data_stage_2__2159_, data_stage_2__2158_, data_stage_2__2157_, data_stage_2__2156_, data_stage_2__2155_, data_stage_2__2154_, data_stage_2__2153_, data_stage_2__2152_, data_stage_2__2151_, data_stage_2__2150_, data_stage_2__2149_, data_stage_2__2148_, data_stage_2__2147_, data_stage_2__2146_, data_stage_2__2145_, data_stage_2__2144_, data_stage_2__2143_, data_stage_2__2142_, data_stage_2__2141_, data_stage_2__2140_, data_stage_2__2139_, data_stage_2__2138_, data_stage_2__2137_, data_stage_2__2136_, data_stage_2__2135_, data_stage_2__2134_, data_stage_2__2133_, data_stage_2__2132_, data_stage_2__2131_, data_stage_2__2130_, data_stage_2__2129_, data_stage_2__2128_, data_stage_2__2127_, data_stage_2__2126_, data_stage_2__2125_, data_stage_2__2124_, data_stage_2__2123_, data_stage_2__2122_, data_stage_2__2121_, data_stage_2__2120_, data_stage_2__2119_, data_stage_2__2118_, data_stage_2__2117_, data_stage_2__2116_, data_stage_2__2115_, data_stage_2__2114_, data_stage_2__2113_, data_stage_2__2112_, data_stage_2__2111_, data_stage_2__2110_, data_stage_2__2109_, data_stage_2__2108_, data_stage_2__2107_, data_stage_2__2106_, data_stage_2__2105_, data_stage_2__2104_, data_stage_2__2103_, data_stage_2__2102_, data_stage_2__2101_, data_stage_2__2100_, data_stage_2__2099_, data_stage_2__2098_, data_stage_2__2097_, data_stage_2__2096_, data_stage_2__2095_, data_stage_2__2094_, data_stage_2__2093_, data_stage_2__2092_, data_stage_2__2091_, data_stage_2__2090_, data_stage_2__2089_, data_stage_2__2088_, data_stage_2__2087_, data_stage_2__2086_, data_stage_2__2085_, data_stage_2__2084_, data_stage_2__2083_, data_stage_2__2082_, data_stage_2__2081_, data_stage_2__2080_, data_stage_2__2079_, data_stage_2__2078_, data_stage_2__2077_, data_stage_2__2076_, data_stage_2__2075_, data_stage_2__2074_, data_stage_2__2073_, data_stage_2__2072_, data_stage_2__2071_, data_stage_2__2070_, data_stage_2__2069_, data_stage_2__2068_, data_stage_2__2067_, data_stage_2__2066_, data_stage_2__2065_, data_stage_2__2064_, data_stage_2__2063_, data_stage_2__2062_, data_stage_2__2061_, data_stage_2__2060_, data_stage_2__2059_, data_stage_2__2058_, data_stage_2__2057_, data_stage_2__2056_, data_stage_2__2055_, data_stage_2__2054_, data_stage_2__2053_, data_stage_2__2052_, data_stage_2__2051_, data_stage_2__2050_, data_stage_2__2049_, data_stage_2__2048_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_5__swap_inst
  (
    .data_i({ data_stage_1__3071_, data_stage_1__3070_, data_stage_1__3069_, data_stage_1__3068_, data_stage_1__3067_, data_stage_1__3066_, data_stage_1__3065_, data_stage_1__3064_, data_stage_1__3063_, data_stage_1__3062_, data_stage_1__3061_, data_stage_1__3060_, data_stage_1__3059_, data_stage_1__3058_, data_stage_1__3057_, data_stage_1__3056_, data_stage_1__3055_, data_stage_1__3054_, data_stage_1__3053_, data_stage_1__3052_, data_stage_1__3051_, data_stage_1__3050_, data_stage_1__3049_, data_stage_1__3048_, data_stage_1__3047_, data_stage_1__3046_, data_stage_1__3045_, data_stage_1__3044_, data_stage_1__3043_, data_stage_1__3042_, data_stage_1__3041_, data_stage_1__3040_, data_stage_1__3039_, data_stage_1__3038_, data_stage_1__3037_, data_stage_1__3036_, data_stage_1__3035_, data_stage_1__3034_, data_stage_1__3033_, data_stage_1__3032_, data_stage_1__3031_, data_stage_1__3030_, data_stage_1__3029_, data_stage_1__3028_, data_stage_1__3027_, data_stage_1__3026_, data_stage_1__3025_, data_stage_1__3024_, data_stage_1__3023_, data_stage_1__3022_, data_stage_1__3021_, data_stage_1__3020_, data_stage_1__3019_, data_stage_1__3018_, data_stage_1__3017_, data_stage_1__3016_, data_stage_1__3015_, data_stage_1__3014_, data_stage_1__3013_, data_stage_1__3012_, data_stage_1__3011_, data_stage_1__3010_, data_stage_1__3009_, data_stage_1__3008_, data_stage_1__3007_, data_stage_1__3006_, data_stage_1__3005_, data_stage_1__3004_, data_stage_1__3003_, data_stage_1__3002_, data_stage_1__3001_, data_stage_1__3000_, data_stage_1__2999_, data_stage_1__2998_, data_stage_1__2997_, data_stage_1__2996_, data_stage_1__2995_, data_stage_1__2994_, data_stage_1__2993_, data_stage_1__2992_, data_stage_1__2991_, data_stage_1__2990_, data_stage_1__2989_, data_stage_1__2988_, data_stage_1__2987_, data_stage_1__2986_, data_stage_1__2985_, data_stage_1__2984_, data_stage_1__2983_, data_stage_1__2982_, data_stage_1__2981_, data_stage_1__2980_, data_stage_1__2979_, data_stage_1__2978_, data_stage_1__2977_, data_stage_1__2976_, data_stage_1__2975_, data_stage_1__2974_, data_stage_1__2973_, data_stage_1__2972_, data_stage_1__2971_, data_stage_1__2970_, data_stage_1__2969_, data_stage_1__2968_, data_stage_1__2967_, data_stage_1__2966_, data_stage_1__2965_, data_stage_1__2964_, data_stage_1__2963_, data_stage_1__2962_, data_stage_1__2961_, data_stage_1__2960_, data_stage_1__2959_, data_stage_1__2958_, data_stage_1__2957_, data_stage_1__2956_, data_stage_1__2955_, data_stage_1__2954_, data_stage_1__2953_, data_stage_1__2952_, data_stage_1__2951_, data_stage_1__2950_, data_stage_1__2949_, data_stage_1__2948_, data_stage_1__2947_, data_stage_1__2946_, data_stage_1__2945_, data_stage_1__2944_, data_stage_1__2943_, data_stage_1__2942_, data_stage_1__2941_, data_stage_1__2940_, data_stage_1__2939_, data_stage_1__2938_, data_stage_1__2937_, data_stage_1__2936_, data_stage_1__2935_, data_stage_1__2934_, data_stage_1__2933_, data_stage_1__2932_, data_stage_1__2931_, data_stage_1__2930_, data_stage_1__2929_, data_stage_1__2928_, data_stage_1__2927_, data_stage_1__2926_, data_stage_1__2925_, data_stage_1__2924_, data_stage_1__2923_, data_stage_1__2922_, data_stage_1__2921_, data_stage_1__2920_, data_stage_1__2919_, data_stage_1__2918_, data_stage_1__2917_, data_stage_1__2916_, data_stage_1__2915_, data_stage_1__2914_, data_stage_1__2913_, data_stage_1__2912_, data_stage_1__2911_, data_stage_1__2910_, data_stage_1__2909_, data_stage_1__2908_, data_stage_1__2907_, data_stage_1__2906_, data_stage_1__2905_, data_stage_1__2904_, data_stage_1__2903_, data_stage_1__2902_, data_stage_1__2901_, data_stage_1__2900_, data_stage_1__2899_, data_stage_1__2898_, data_stage_1__2897_, data_stage_1__2896_, data_stage_1__2895_, data_stage_1__2894_, data_stage_1__2893_, data_stage_1__2892_, data_stage_1__2891_, data_stage_1__2890_, data_stage_1__2889_, data_stage_1__2888_, data_stage_1__2887_, data_stage_1__2886_, data_stage_1__2885_, data_stage_1__2884_, data_stage_1__2883_, data_stage_1__2882_, data_stage_1__2881_, data_stage_1__2880_, data_stage_1__2879_, data_stage_1__2878_, data_stage_1__2877_, data_stage_1__2876_, data_stage_1__2875_, data_stage_1__2874_, data_stage_1__2873_, data_stage_1__2872_, data_stage_1__2871_, data_stage_1__2870_, data_stage_1__2869_, data_stage_1__2868_, data_stage_1__2867_, data_stage_1__2866_, data_stage_1__2865_, data_stage_1__2864_, data_stage_1__2863_, data_stage_1__2862_, data_stage_1__2861_, data_stage_1__2860_, data_stage_1__2859_, data_stage_1__2858_, data_stage_1__2857_, data_stage_1__2856_, data_stage_1__2855_, data_stage_1__2854_, data_stage_1__2853_, data_stage_1__2852_, data_stage_1__2851_, data_stage_1__2850_, data_stage_1__2849_, data_stage_1__2848_, data_stage_1__2847_, data_stage_1__2846_, data_stage_1__2845_, data_stage_1__2844_, data_stage_1__2843_, data_stage_1__2842_, data_stage_1__2841_, data_stage_1__2840_, data_stage_1__2839_, data_stage_1__2838_, data_stage_1__2837_, data_stage_1__2836_, data_stage_1__2835_, data_stage_1__2834_, data_stage_1__2833_, data_stage_1__2832_, data_stage_1__2831_, data_stage_1__2830_, data_stage_1__2829_, data_stage_1__2828_, data_stage_1__2827_, data_stage_1__2826_, data_stage_1__2825_, data_stage_1__2824_, data_stage_1__2823_, data_stage_1__2822_, data_stage_1__2821_, data_stage_1__2820_, data_stage_1__2819_, data_stage_1__2818_, data_stage_1__2817_, data_stage_1__2816_, data_stage_1__2815_, data_stage_1__2814_, data_stage_1__2813_, data_stage_1__2812_, data_stage_1__2811_, data_stage_1__2810_, data_stage_1__2809_, data_stage_1__2808_, data_stage_1__2807_, data_stage_1__2806_, data_stage_1__2805_, data_stage_1__2804_, data_stage_1__2803_, data_stage_1__2802_, data_stage_1__2801_, data_stage_1__2800_, data_stage_1__2799_, data_stage_1__2798_, data_stage_1__2797_, data_stage_1__2796_, data_stage_1__2795_, data_stage_1__2794_, data_stage_1__2793_, data_stage_1__2792_, data_stage_1__2791_, data_stage_1__2790_, data_stage_1__2789_, data_stage_1__2788_, data_stage_1__2787_, data_stage_1__2786_, data_stage_1__2785_, data_stage_1__2784_, data_stage_1__2783_, data_stage_1__2782_, data_stage_1__2781_, data_stage_1__2780_, data_stage_1__2779_, data_stage_1__2778_, data_stage_1__2777_, data_stage_1__2776_, data_stage_1__2775_, data_stage_1__2774_, data_stage_1__2773_, data_stage_1__2772_, data_stage_1__2771_, data_stage_1__2770_, data_stage_1__2769_, data_stage_1__2768_, data_stage_1__2767_, data_stage_1__2766_, data_stage_1__2765_, data_stage_1__2764_, data_stage_1__2763_, data_stage_1__2762_, data_stage_1__2761_, data_stage_1__2760_, data_stage_1__2759_, data_stage_1__2758_, data_stage_1__2757_, data_stage_1__2756_, data_stage_1__2755_, data_stage_1__2754_, data_stage_1__2753_, data_stage_1__2752_, data_stage_1__2751_, data_stage_1__2750_, data_stage_1__2749_, data_stage_1__2748_, data_stage_1__2747_, data_stage_1__2746_, data_stage_1__2745_, data_stage_1__2744_, data_stage_1__2743_, data_stage_1__2742_, data_stage_1__2741_, data_stage_1__2740_, data_stage_1__2739_, data_stage_1__2738_, data_stage_1__2737_, data_stage_1__2736_, data_stage_1__2735_, data_stage_1__2734_, data_stage_1__2733_, data_stage_1__2732_, data_stage_1__2731_, data_stage_1__2730_, data_stage_1__2729_, data_stage_1__2728_, data_stage_1__2727_, data_stage_1__2726_, data_stage_1__2725_, data_stage_1__2724_, data_stage_1__2723_, data_stage_1__2722_, data_stage_1__2721_, data_stage_1__2720_, data_stage_1__2719_, data_stage_1__2718_, data_stage_1__2717_, data_stage_1__2716_, data_stage_1__2715_, data_stage_1__2714_, data_stage_1__2713_, data_stage_1__2712_, data_stage_1__2711_, data_stage_1__2710_, data_stage_1__2709_, data_stage_1__2708_, data_stage_1__2707_, data_stage_1__2706_, data_stage_1__2705_, data_stage_1__2704_, data_stage_1__2703_, data_stage_1__2702_, data_stage_1__2701_, data_stage_1__2700_, data_stage_1__2699_, data_stage_1__2698_, data_stage_1__2697_, data_stage_1__2696_, data_stage_1__2695_, data_stage_1__2694_, data_stage_1__2693_, data_stage_1__2692_, data_stage_1__2691_, data_stage_1__2690_, data_stage_1__2689_, data_stage_1__2688_, data_stage_1__2687_, data_stage_1__2686_, data_stage_1__2685_, data_stage_1__2684_, data_stage_1__2683_, data_stage_1__2682_, data_stage_1__2681_, data_stage_1__2680_, data_stage_1__2679_, data_stage_1__2678_, data_stage_1__2677_, data_stage_1__2676_, data_stage_1__2675_, data_stage_1__2674_, data_stage_1__2673_, data_stage_1__2672_, data_stage_1__2671_, data_stage_1__2670_, data_stage_1__2669_, data_stage_1__2668_, data_stage_1__2667_, data_stage_1__2666_, data_stage_1__2665_, data_stage_1__2664_, data_stage_1__2663_, data_stage_1__2662_, data_stage_1__2661_, data_stage_1__2660_, data_stage_1__2659_, data_stage_1__2658_, data_stage_1__2657_, data_stage_1__2656_, data_stage_1__2655_, data_stage_1__2654_, data_stage_1__2653_, data_stage_1__2652_, data_stage_1__2651_, data_stage_1__2650_, data_stage_1__2649_, data_stage_1__2648_, data_stage_1__2647_, data_stage_1__2646_, data_stage_1__2645_, data_stage_1__2644_, data_stage_1__2643_, data_stage_1__2642_, data_stage_1__2641_, data_stage_1__2640_, data_stage_1__2639_, data_stage_1__2638_, data_stage_1__2637_, data_stage_1__2636_, data_stage_1__2635_, data_stage_1__2634_, data_stage_1__2633_, data_stage_1__2632_, data_stage_1__2631_, data_stage_1__2630_, data_stage_1__2629_, data_stage_1__2628_, data_stage_1__2627_, data_stage_1__2626_, data_stage_1__2625_, data_stage_1__2624_, data_stage_1__2623_, data_stage_1__2622_, data_stage_1__2621_, data_stage_1__2620_, data_stage_1__2619_, data_stage_1__2618_, data_stage_1__2617_, data_stage_1__2616_, data_stage_1__2615_, data_stage_1__2614_, data_stage_1__2613_, data_stage_1__2612_, data_stage_1__2611_, data_stage_1__2610_, data_stage_1__2609_, data_stage_1__2608_, data_stage_1__2607_, data_stage_1__2606_, data_stage_1__2605_, data_stage_1__2604_, data_stage_1__2603_, data_stage_1__2602_, data_stage_1__2601_, data_stage_1__2600_, data_stage_1__2599_, data_stage_1__2598_, data_stage_1__2597_, data_stage_1__2596_, data_stage_1__2595_, data_stage_1__2594_, data_stage_1__2593_, data_stage_1__2592_, data_stage_1__2591_, data_stage_1__2590_, data_stage_1__2589_, data_stage_1__2588_, data_stage_1__2587_, data_stage_1__2586_, data_stage_1__2585_, data_stage_1__2584_, data_stage_1__2583_, data_stage_1__2582_, data_stage_1__2581_, data_stage_1__2580_, data_stage_1__2579_, data_stage_1__2578_, data_stage_1__2577_, data_stage_1__2576_, data_stage_1__2575_, data_stage_1__2574_, data_stage_1__2573_, data_stage_1__2572_, data_stage_1__2571_, data_stage_1__2570_, data_stage_1__2569_, data_stage_1__2568_, data_stage_1__2567_, data_stage_1__2566_, data_stage_1__2565_, data_stage_1__2564_, data_stage_1__2563_, data_stage_1__2562_, data_stage_1__2561_, data_stage_1__2560_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__3071_, data_stage_2__3070_, data_stage_2__3069_, data_stage_2__3068_, data_stage_2__3067_, data_stage_2__3066_, data_stage_2__3065_, data_stage_2__3064_, data_stage_2__3063_, data_stage_2__3062_, data_stage_2__3061_, data_stage_2__3060_, data_stage_2__3059_, data_stage_2__3058_, data_stage_2__3057_, data_stage_2__3056_, data_stage_2__3055_, data_stage_2__3054_, data_stage_2__3053_, data_stage_2__3052_, data_stage_2__3051_, data_stage_2__3050_, data_stage_2__3049_, data_stage_2__3048_, data_stage_2__3047_, data_stage_2__3046_, data_stage_2__3045_, data_stage_2__3044_, data_stage_2__3043_, data_stage_2__3042_, data_stage_2__3041_, data_stage_2__3040_, data_stage_2__3039_, data_stage_2__3038_, data_stage_2__3037_, data_stage_2__3036_, data_stage_2__3035_, data_stage_2__3034_, data_stage_2__3033_, data_stage_2__3032_, data_stage_2__3031_, data_stage_2__3030_, data_stage_2__3029_, data_stage_2__3028_, data_stage_2__3027_, data_stage_2__3026_, data_stage_2__3025_, data_stage_2__3024_, data_stage_2__3023_, data_stage_2__3022_, data_stage_2__3021_, data_stage_2__3020_, data_stage_2__3019_, data_stage_2__3018_, data_stage_2__3017_, data_stage_2__3016_, data_stage_2__3015_, data_stage_2__3014_, data_stage_2__3013_, data_stage_2__3012_, data_stage_2__3011_, data_stage_2__3010_, data_stage_2__3009_, data_stage_2__3008_, data_stage_2__3007_, data_stage_2__3006_, data_stage_2__3005_, data_stage_2__3004_, data_stage_2__3003_, data_stage_2__3002_, data_stage_2__3001_, data_stage_2__3000_, data_stage_2__2999_, data_stage_2__2998_, data_stage_2__2997_, data_stage_2__2996_, data_stage_2__2995_, data_stage_2__2994_, data_stage_2__2993_, data_stage_2__2992_, data_stage_2__2991_, data_stage_2__2990_, data_stage_2__2989_, data_stage_2__2988_, data_stage_2__2987_, data_stage_2__2986_, data_stage_2__2985_, data_stage_2__2984_, data_stage_2__2983_, data_stage_2__2982_, data_stage_2__2981_, data_stage_2__2980_, data_stage_2__2979_, data_stage_2__2978_, data_stage_2__2977_, data_stage_2__2976_, data_stage_2__2975_, data_stage_2__2974_, data_stage_2__2973_, data_stage_2__2972_, data_stage_2__2971_, data_stage_2__2970_, data_stage_2__2969_, data_stage_2__2968_, data_stage_2__2967_, data_stage_2__2966_, data_stage_2__2965_, data_stage_2__2964_, data_stage_2__2963_, data_stage_2__2962_, data_stage_2__2961_, data_stage_2__2960_, data_stage_2__2959_, data_stage_2__2958_, data_stage_2__2957_, data_stage_2__2956_, data_stage_2__2955_, data_stage_2__2954_, data_stage_2__2953_, data_stage_2__2952_, data_stage_2__2951_, data_stage_2__2950_, data_stage_2__2949_, data_stage_2__2948_, data_stage_2__2947_, data_stage_2__2946_, data_stage_2__2945_, data_stage_2__2944_, data_stage_2__2943_, data_stage_2__2942_, data_stage_2__2941_, data_stage_2__2940_, data_stage_2__2939_, data_stage_2__2938_, data_stage_2__2937_, data_stage_2__2936_, data_stage_2__2935_, data_stage_2__2934_, data_stage_2__2933_, data_stage_2__2932_, data_stage_2__2931_, data_stage_2__2930_, data_stage_2__2929_, data_stage_2__2928_, data_stage_2__2927_, data_stage_2__2926_, data_stage_2__2925_, data_stage_2__2924_, data_stage_2__2923_, data_stage_2__2922_, data_stage_2__2921_, data_stage_2__2920_, data_stage_2__2919_, data_stage_2__2918_, data_stage_2__2917_, data_stage_2__2916_, data_stage_2__2915_, data_stage_2__2914_, data_stage_2__2913_, data_stage_2__2912_, data_stage_2__2911_, data_stage_2__2910_, data_stage_2__2909_, data_stage_2__2908_, data_stage_2__2907_, data_stage_2__2906_, data_stage_2__2905_, data_stage_2__2904_, data_stage_2__2903_, data_stage_2__2902_, data_stage_2__2901_, data_stage_2__2900_, data_stage_2__2899_, data_stage_2__2898_, data_stage_2__2897_, data_stage_2__2896_, data_stage_2__2895_, data_stage_2__2894_, data_stage_2__2893_, data_stage_2__2892_, data_stage_2__2891_, data_stage_2__2890_, data_stage_2__2889_, data_stage_2__2888_, data_stage_2__2887_, data_stage_2__2886_, data_stage_2__2885_, data_stage_2__2884_, data_stage_2__2883_, data_stage_2__2882_, data_stage_2__2881_, data_stage_2__2880_, data_stage_2__2879_, data_stage_2__2878_, data_stage_2__2877_, data_stage_2__2876_, data_stage_2__2875_, data_stage_2__2874_, data_stage_2__2873_, data_stage_2__2872_, data_stage_2__2871_, data_stage_2__2870_, data_stage_2__2869_, data_stage_2__2868_, data_stage_2__2867_, data_stage_2__2866_, data_stage_2__2865_, data_stage_2__2864_, data_stage_2__2863_, data_stage_2__2862_, data_stage_2__2861_, data_stage_2__2860_, data_stage_2__2859_, data_stage_2__2858_, data_stage_2__2857_, data_stage_2__2856_, data_stage_2__2855_, data_stage_2__2854_, data_stage_2__2853_, data_stage_2__2852_, data_stage_2__2851_, data_stage_2__2850_, data_stage_2__2849_, data_stage_2__2848_, data_stage_2__2847_, data_stage_2__2846_, data_stage_2__2845_, data_stage_2__2844_, data_stage_2__2843_, data_stage_2__2842_, data_stage_2__2841_, data_stage_2__2840_, data_stage_2__2839_, data_stage_2__2838_, data_stage_2__2837_, data_stage_2__2836_, data_stage_2__2835_, data_stage_2__2834_, data_stage_2__2833_, data_stage_2__2832_, data_stage_2__2831_, data_stage_2__2830_, data_stage_2__2829_, data_stage_2__2828_, data_stage_2__2827_, data_stage_2__2826_, data_stage_2__2825_, data_stage_2__2824_, data_stage_2__2823_, data_stage_2__2822_, data_stage_2__2821_, data_stage_2__2820_, data_stage_2__2819_, data_stage_2__2818_, data_stage_2__2817_, data_stage_2__2816_, data_stage_2__2815_, data_stage_2__2814_, data_stage_2__2813_, data_stage_2__2812_, data_stage_2__2811_, data_stage_2__2810_, data_stage_2__2809_, data_stage_2__2808_, data_stage_2__2807_, data_stage_2__2806_, data_stage_2__2805_, data_stage_2__2804_, data_stage_2__2803_, data_stage_2__2802_, data_stage_2__2801_, data_stage_2__2800_, data_stage_2__2799_, data_stage_2__2798_, data_stage_2__2797_, data_stage_2__2796_, data_stage_2__2795_, data_stage_2__2794_, data_stage_2__2793_, data_stage_2__2792_, data_stage_2__2791_, data_stage_2__2790_, data_stage_2__2789_, data_stage_2__2788_, data_stage_2__2787_, data_stage_2__2786_, data_stage_2__2785_, data_stage_2__2784_, data_stage_2__2783_, data_stage_2__2782_, data_stage_2__2781_, data_stage_2__2780_, data_stage_2__2779_, data_stage_2__2778_, data_stage_2__2777_, data_stage_2__2776_, data_stage_2__2775_, data_stage_2__2774_, data_stage_2__2773_, data_stage_2__2772_, data_stage_2__2771_, data_stage_2__2770_, data_stage_2__2769_, data_stage_2__2768_, data_stage_2__2767_, data_stage_2__2766_, data_stage_2__2765_, data_stage_2__2764_, data_stage_2__2763_, data_stage_2__2762_, data_stage_2__2761_, data_stage_2__2760_, data_stage_2__2759_, data_stage_2__2758_, data_stage_2__2757_, data_stage_2__2756_, data_stage_2__2755_, data_stage_2__2754_, data_stage_2__2753_, data_stage_2__2752_, data_stage_2__2751_, data_stage_2__2750_, data_stage_2__2749_, data_stage_2__2748_, data_stage_2__2747_, data_stage_2__2746_, data_stage_2__2745_, data_stage_2__2744_, data_stage_2__2743_, data_stage_2__2742_, data_stage_2__2741_, data_stage_2__2740_, data_stage_2__2739_, data_stage_2__2738_, data_stage_2__2737_, data_stage_2__2736_, data_stage_2__2735_, data_stage_2__2734_, data_stage_2__2733_, data_stage_2__2732_, data_stage_2__2731_, data_stage_2__2730_, data_stage_2__2729_, data_stage_2__2728_, data_stage_2__2727_, data_stage_2__2726_, data_stage_2__2725_, data_stage_2__2724_, data_stage_2__2723_, data_stage_2__2722_, data_stage_2__2721_, data_stage_2__2720_, data_stage_2__2719_, data_stage_2__2718_, data_stage_2__2717_, data_stage_2__2716_, data_stage_2__2715_, data_stage_2__2714_, data_stage_2__2713_, data_stage_2__2712_, data_stage_2__2711_, data_stage_2__2710_, data_stage_2__2709_, data_stage_2__2708_, data_stage_2__2707_, data_stage_2__2706_, data_stage_2__2705_, data_stage_2__2704_, data_stage_2__2703_, data_stage_2__2702_, data_stage_2__2701_, data_stage_2__2700_, data_stage_2__2699_, data_stage_2__2698_, data_stage_2__2697_, data_stage_2__2696_, data_stage_2__2695_, data_stage_2__2694_, data_stage_2__2693_, data_stage_2__2692_, data_stage_2__2691_, data_stage_2__2690_, data_stage_2__2689_, data_stage_2__2688_, data_stage_2__2687_, data_stage_2__2686_, data_stage_2__2685_, data_stage_2__2684_, data_stage_2__2683_, data_stage_2__2682_, data_stage_2__2681_, data_stage_2__2680_, data_stage_2__2679_, data_stage_2__2678_, data_stage_2__2677_, data_stage_2__2676_, data_stage_2__2675_, data_stage_2__2674_, data_stage_2__2673_, data_stage_2__2672_, data_stage_2__2671_, data_stage_2__2670_, data_stage_2__2669_, data_stage_2__2668_, data_stage_2__2667_, data_stage_2__2666_, data_stage_2__2665_, data_stage_2__2664_, data_stage_2__2663_, data_stage_2__2662_, data_stage_2__2661_, data_stage_2__2660_, data_stage_2__2659_, data_stage_2__2658_, data_stage_2__2657_, data_stage_2__2656_, data_stage_2__2655_, data_stage_2__2654_, data_stage_2__2653_, data_stage_2__2652_, data_stage_2__2651_, data_stage_2__2650_, data_stage_2__2649_, data_stage_2__2648_, data_stage_2__2647_, data_stage_2__2646_, data_stage_2__2645_, data_stage_2__2644_, data_stage_2__2643_, data_stage_2__2642_, data_stage_2__2641_, data_stage_2__2640_, data_stage_2__2639_, data_stage_2__2638_, data_stage_2__2637_, data_stage_2__2636_, data_stage_2__2635_, data_stage_2__2634_, data_stage_2__2633_, data_stage_2__2632_, data_stage_2__2631_, data_stage_2__2630_, data_stage_2__2629_, data_stage_2__2628_, data_stage_2__2627_, data_stage_2__2626_, data_stage_2__2625_, data_stage_2__2624_, data_stage_2__2623_, data_stage_2__2622_, data_stage_2__2621_, data_stage_2__2620_, data_stage_2__2619_, data_stage_2__2618_, data_stage_2__2617_, data_stage_2__2616_, data_stage_2__2615_, data_stage_2__2614_, data_stage_2__2613_, data_stage_2__2612_, data_stage_2__2611_, data_stage_2__2610_, data_stage_2__2609_, data_stage_2__2608_, data_stage_2__2607_, data_stage_2__2606_, data_stage_2__2605_, data_stage_2__2604_, data_stage_2__2603_, data_stage_2__2602_, data_stage_2__2601_, data_stage_2__2600_, data_stage_2__2599_, data_stage_2__2598_, data_stage_2__2597_, data_stage_2__2596_, data_stage_2__2595_, data_stage_2__2594_, data_stage_2__2593_, data_stage_2__2592_, data_stage_2__2591_, data_stage_2__2590_, data_stage_2__2589_, data_stage_2__2588_, data_stage_2__2587_, data_stage_2__2586_, data_stage_2__2585_, data_stage_2__2584_, data_stage_2__2583_, data_stage_2__2582_, data_stage_2__2581_, data_stage_2__2580_, data_stage_2__2579_, data_stage_2__2578_, data_stage_2__2577_, data_stage_2__2576_, data_stage_2__2575_, data_stage_2__2574_, data_stage_2__2573_, data_stage_2__2572_, data_stage_2__2571_, data_stage_2__2570_, data_stage_2__2569_, data_stage_2__2568_, data_stage_2__2567_, data_stage_2__2566_, data_stage_2__2565_, data_stage_2__2564_, data_stage_2__2563_, data_stage_2__2562_, data_stage_2__2561_, data_stage_2__2560_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_6__swap_inst
  (
    .data_i({ data_stage_1__3583_, data_stage_1__3582_, data_stage_1__3581_, data_stage_1__3580_, data_stage_1__3579_, data_stage_1__3578_, data_stage_1__3577_, data_stage_1__3576_, data_stage_1__3575_, data_stage_1__3574_, data_stage_1__3573_, data_stage_1__3572_, data_stage_1__3571_, data_stage_1__3570_, data_stage_1__3569_, data_stage_1__3568_, data_stage_1__3567_, data_stage_1__3566_, data_stage_1__3565_, data_stage_1__3564_, data_stage_1__3563_, data_stage_1__3562_, data_stage_1__3561_, data_stage_1__3560_, data_stage_1__3559_, data_stage_1__3558_, data_stage_1__3557_, data_stage_1__3556_, data_stage_1__3555_, data_stage_1__3554_, data_stage_1__3553_, data_stage_1__3552_, data_stage_1__3551_, data_stage_1__3550_, data_stage_1__3549_, data_stage_1__3548_, data_stage_1__3547_, data_stage_1__3546_, data_stage_1__3545_, data_stage_1__3544_, data_stage_1__3543_, data_stage_1__3542_, data_stage_1__3541_, data_stage_1__3540_, data_stage_1__3539_, data_stage_1__3538_, data_stage_1__3537_, data_stage_1__3536_, data_stage_1__3535_, data_stage_1__3534_, data_stage_1__3533_, data_stage_1__3532_, data_stage_1__3531_, data_stage_1__3530_, data_stage_1__3529_, data_stage_1__3528_, data_stage_1__3527_, data_stage_1__3526_, data_stage_1__3525_, data_stage_1__3524_, data_stage_1__3523_, data_stage_1__3522_, data_stage_1__3521_, data_stage_1__3520_, data_stage_1__3519_, data_stage_1__3518_, data_stage_1__3517_, data_stage_1__3516_, data_stage_1__3515_, data_stage_1__3514_, data_stage_1__3513_, data_stage_1__3512_, data_stage_1__3511_, data_stage_1__3510_, data_stage_1__3509_, data_stage_1__3508_, data_stage_1__3507_, data_stage_1__3506_, data_stage_1__3505_, data_stage_1__3504_, data_stage_1__3503_, data_stage_1__3502_, data_stage_1__3501_, data_stage_1__3500_, data_stage_1__3499_, data_stage_1__3498_, data_stage_1__3497_, data_stage_1__3496_, data_stage_1__3495_, data_stage_1__3494_, data_stage_1__3493_, data_stage_1__3492_, data_stage_1__3491_, data_stage_1__3490_, data_stage_1__3489_, data_stage_1__3488_, data_stage_1__3487_, data_stage_1__3486_, data_stage_1__3485_, data_stage_1__3484_, data_stage_1__3483_, data_stage_1__3482_, data_stage_1__3481_, data_stage_1__3480_, data_stage_1__3479_, data_stage_1__3478_, data_stage_1__3477_, data_stage_1__3476_, data_stage_1__3475_, data_stage_1__3474_, data_stage_1__3473_, data_stage_1__3472_, data_stage_1__3471_, data_stage_1__3470_, data_stage_1__3469_, data_stage_1__3468_, data_stage_1__3467_, data_stage_1__3466_, data_stage_1__3465_, data_stage_1__3464_, data_stage_1__3463_, data_stage_1__3462_, data_stage_1__3461_, data_stage_1__3460_, data_stage_1__3459_, data_stage_1__3458_, data_stage_1__3457_, data_stage_1__3456_, data_stage_1__3455_, data_stage_1__3454_, data_stage_1__3453_, data_stage_1__3452_, data_stage_1__3451_, data_stage_1__3450_, data_stage_1__3449_, data_stage_1__3448_, data_stage_1__3447_, data_stage_1__3446_, data_stage_1__3445_, data_stage_1__3444_, data_stage_1__3443_, data_stage_1__3442_, data_stage_1__3441_, data_stage_1__3440_, data_stage_1__3439_, data_stage_1__3438_, data_stage_1__3437_, data_stage_1__3436_, data_stage_1__3435_, data_stage_1__3434_, data_stage_1__3433_, data_stage_1__3432_, data_stage_1__3431_, data_stage_1__3430_, data_stage_1__3429_, data_stage_1__3428_, data_stage_1__3427_, data_stage_1__3426_, data_stage_1__3425_, data_stage_1__3424_, data_stage_1__3423_, data_stage_1__3422_, data_stage_1__3421_, data_stage_1__3420_, data_stage_1__3419_, data_stage_1__3418_, data_stage_1__3417_, data_stage_1__3416_, data_stage_1__3415_, data_stage_1__3414_, data_stage_1__3413_, data_stage_1__3412_, data_stage_1__3411_, data_stage_1__3410_, data_stage_1__3409_, data_stage_1__3408_, data_stage_1__3407_, data_stage_1__3406_, data_stage_1__3405_, data_stage_1__3404_, data_stage_1__3403_, data_stage_1__3402_, data_stage_1__3401_, data_stage_1__3400_, data_stage_1__3399_, data_stage_1__3398_, data_stage_1__3397_, data_stage_1__3396_, data_stage_1__3395_, data_stage_1__3394_, data_stage_1__3393_, data_stage_1__3392_, data_stage_1__3391_, data_stage_1__3390_, data_stage_1__3389_, data_stage_1__3388_, data_stage_1__3387_, data_stage_1__3386_, data_stage_1__3385_, data_stage_1__3384_, data_stage_1__3383_, data_stage_1__3382_, data_stage_1__3381_, data_stage_1__3380_, data_stage_1__3379_, data_stage_1__3378_, data_stage_1__3377_, data_stage_1__3376_, data_stage_1__3375_, data_stage_1__3374_, data_stage_1__3373_, data_stage_1__3372_, data_stage_1__3371_, data_stage_1__3370_, data_stage_1__3369_, data_stage_1__3368_, data_stage_1__3367_, data_stage_1__3366_, data_stage_1__3365_, data_stage_1__3364_, data_stage_1__3363_, data_stage_1__3362_, data_stage_1__3361_, data_stage_1__3360_, data_stage_1__3359_, data_stage_1__3358_, data_stage_1__3357_, data_stage_1__3356_, data_stage_1__3355_, data_stage_1__3354_, data_stage_1__3353_, data_stage_1__3352_, data_stage_1__3351_, data_stage_1__3350_, data_stage_1__3349_, data_stage_1__3348_, data_stage_1__3347_, data_stage_1__3346_, data_stage_1__3345_, data_stage_1__3344_, data_stage_1__3343_, data_stage_1__3342_, data_stage_1__3341_, data_stage_1__3340_, data_stage_1__3339_, data_stage_1__3338_, data_stage_1__3337_, data_stage_1__3336_, data_stage_1__3335_, data_stage_1__3334_, data_stage_1__3333_, data_stage_1__3332_, data_stage_1__3331_, data_stage_1__3330_, data_stage_1__3329_, data_stage_1__3328_, data_stage_1__3327_, data_stage_1__3326_, data_stage_1__3325_, data_stage_1__3324_, data_stage_1__3323_, data_stage_1__3322_, data_stage_1__3321_, data_stage_1__3320_, data_stage_1__3319_, data_stage_1__3318_, data_stage_1__3317_, data_stage_1__3316_, data_stage_1__3315_, data_stage_1__3314_, data_stage_1__3313_, data_stage_1__3312_, data_stage_1__3311_, data_stage_1__3310_, data_stage_1__3309_, data_stage_1__3308_, data_stage_1__3307_, data_stage_1__3306_, data_stage_1__3305_, data_stage_1__3304_, data_stage_1__3303_, data_stage_1__3302_, data_stage_1__3301_, data_stage_1__3300_, data_stage_1__3299_, data_stage_1__3298_, data_stage_1__3297_, data_stage_1__3296_, data_stage_1__3295_, data_stage_1__3294_, data_stage_1__3293_, data_stage_1__3292_, data_stage_1__3291_, data_stage_1__3290_, data_stage_1__3289_, data_stage_1__3288_, data_stage_1__3287_, data_stage_1__3286_, data_stage_1__3285_, data_stage_1__3284_, data_stage_1__3283_, data_stage_1__3282_, data_stage_1__3281_, data_stage_1__3280_, data_stage_1__3279_, data_stage_1__3278_, data_stage_1__3277_, data_stage_1__3276_, data_stage_1__3275_, data_stage_1__3274_, data_stage_1__3273_, data_stage_1__3272_, data_stage_1__3271_, data_stage_1__3270_, data_stage_1__3269_, data_stage_1__3268_, data_stage_1__3267_, data_stage_1__3266_, data_stage_1__3265_, data_stage_1__3264_, data_stage_1__3263_, data_stage_1__3262_, data_stage_1__3261_, data_stage_1__3260_, data_stage_1__3259_, data_stage_1__3258_, data_stage_1__3257_, data_stage_1__3256_, data_stage_1__3255_, data_stage_1__3254_, data_stage_1__3253_, data_stage_1__3252_, data_stage_1__3251_, data_stage_1__3250_, data_stage_1__3249_, data_stage_1__3248_, data_stage_1__3247_, data_stage_1__3246_, data_stage_1__3245_, data_stage_1__3244_, data_stage_1__3243_, data_stage_1__3242_, data_stage_1__3241_, data_stage_1__3240_, data_stage_1__3239_, data_stage_1__3238_, data_stage_1__3237_, data_stage_1__3236_, data_stage_1__3235_, data_stage_1__3234_, data_stage_1__3233_, data_stage_1__3232_, data_stage_1__3231_, data_stage_1__3230_, data_stage_1__3229_, data_stage_1__3228_, data_stage_1__3227_, data_stage_1__3226_, data_stage_1__3225_, data_stage_1__3224_, data_stage_1__3223_, data_stage_1__3222_, data_stage_1__3221_, data_stage_1__3220_, data_stage_1__3219_, data_stage_1__3218_, data_stage_1__3217_, data_stage_1__3216_, data_stage_1__3215_, data_stage_1__3214_, data_stage_1__3213_, data_stage_1__3212_, data_stage_1__3211_, data_stage_1__3210_, data_stage_1__3209_, data_stage_1__3208_, data_stage_1__3207_, data_stage_1__3206_, data_stage_1__3205_, data_stage_1__3204_, data_stage_1__3203_, data_stage_1__3202_, data_stage_1__3201_, data_stage_1__3200_, data_stage_1__3199_, data_stage_1__3198_, data_stage_1__3197_, data_stage_1__3196_, data_stage_1__3195_, data_stage_1__3194_, data_stage_1__3193_, data_stage_1__3192_, data_stage_1__3191_, data_stage_1__3190_, data_stage_1__3189_, data_stage_1__3188_, data_stage_1__3187_, data_stage_1__3186_, data_stage_1__3185_, data_stage_1__3184_, data_stage_1__3183_, data_stage_1__3182_, data_stage_1__3181_, data_stage_1__3180_, data_stage_1__3179_, data_stage_1__3178_, data_stage_1__3177_, data_stage_1__3176_, data_stage_1__3175_, data_stage_1__3174_, data_stage_1__3173_, data_stage_1__3172_, data_stage_1__3171_, data_stage_1__3170_, data_stage_1__3169_, data_stage_1__3168_, data_stage_1__3167_, data_stage_1__3166_, data_stage_1__3165_, data_stage_1__3164_, data_stage_1__3163_, data_stage_1__3162_, data_stage_1__3161_, data_stage_1__3160_, data_stage_1__3159_, data_stage_1__3158_, data_stage_1__3157_, data_stage_1__3156_, data_stage_1__3155_, data_stage_1__3154_, data_stage_1__3153_, data_stage_1__3152_, data_stage_1__3151_, data_stage_1__3150_, data_stage_1__3149_, data_stage_1__3148_, data_stage_1__3147_, data_stage_1__3146_, data_stage_1__3145_, data_stage_1__3144_, data_stage_1__3143_, data_stage_1__3142_, data_stage_1__3141_, data_stage_1__3140_, data_stage_1__3139_, data_stage_1__3138_, data_stage_1__3137_, data_stage_1__3136_, data_stage_1__3135_, data_stage_1__3134_, data_stage_1__3133_, data_stage_1__3132_, data_stage_1__3131_, data_stage_1__3130_, data_stage_1__3129_, data_stage_1__3128_, data_stage_1__3127_, data_stage_1__3126_, data_stage_1__3125_, data_stage_1__3124_, data_stage_1__3123_, data_stage_1__3122_, data_stage_1__3121_, data_stage_1__3120_, data_stage_1__3119_, data_stage_1__3118_, data_stage_1__3117_, data_stage_1__3116_, data_stage_1__3115_, data_stage_1__3114_, data_stage_1__3113_, data_stage_1__3112_, data_stage_1__3111_, data_stage_1__3110_, data_stage_1__3109_, data_stage_1__3108_, data_stage_1__3107_, data_stage_1__3106_, data_stage_1__3105_, data_stage_1__3104_, data_stage_1__3103_, data_stage_1__3102_, data_stage_1__3101_, data_stage_1__3100_, data_stage_1__3099_, data_stage_1__3098_, data_stage_1__3097_, data_stage_1__3096_, data_stage_1__3095_, data_stage_1__3094_, data_stage_1__3093_, data_stage_1__3092_, data_stage_1__3091_, data_stage_1__3090_, data_stage_1__3089_, data_stage_1__3088_, data_stage_1__3087_, data_stage_1__3086_, data_stage_1__3085_, data_stage_1__3084_, data_stage_1__3083_, data_stage_1__3082_, data_stage_1__3081_, data_stage_1__3080_, data_stage_1__3079_, data_stage_1__3078_, data_stage_1__3077_, data_stage_1__3076_, data_stage_1__3075_, data_stage_1__3074_, data_stage_1__3073_, data_stage_1__3072_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__3583_, data_stage_2__3582_, data_stage_2__3581_, data_stage_2__3580_, data_stage_2__3579_, data_stage_2__3578_, data_stage_2__3577_, data_stage_2__3576_, data_stage_2__3575_, data_stage_2__3574_, data_stage_2__3573_, data_stage_2__3572_, data_stage_2__3571_, data_stage_2__3570_, data_stage_2__3569_, data_stage_2__3568_, data_stage_2__3567_, data_stage_2__3566_, data_stage_2__3565_, data_stage_2__3564_, data_stage_2__3563_, data_stage_2__3562_, data_stage_2__3561_, data_stage_2__3560_, data_stage_2__3559_, data_stage_2__3558_, data_stage_2__3557_, data_stage_2__3556_, data_stage_2__3555_, data_stage_2__3554_, data_stage_2__3553_, data_stage_2__3552_, data_stage_2__3551_, data_stage_2__3550_, data_stage_2__3549_, data_stage_2__3548_, data_stage_2__3547_, data_stage_2__3546_, data_stage_2__3545_, data_stage_2__3544_, data_stage_2__3543_, data_stage_2__3542_, data_stage_2__3541_, data_stage_2__3540_, data_stage_2__3539_, data_stage_2__3538_, data_stage_2__3537_, data_stage_2__3536_, data_stage_2__3535_, data_stage_2__3534_, data_stage_2__3533_, data_stage_2__3532_, data_stage_2__3531_, data_stage_2__3530_, data_stage_2__3529_, data_stage_2__3528_, data_stage_2__3527_, data_stage_2__3526_, data_stage_2__3525_, data_stage_2__3524_, data_stage_2__3523_, data_stage_2__3522_, data_stage_2__3521_, data_stage_2__3520_, data_stage_2__3519_, data_stage_2__3518_, data_stage_2__3517_, data_stage_2__3516_, data_stage_2__3515_, data_stage_2__3514_, data_stage_2__3513_, data_stage_2__3512_, data_stage_2__3511_, data_stage_2__3510_, data_stage_2__3509_, data_stage_2__3508_, data_stage_2__3507_, data_stage_2__3506_, data_stage_2__3505_, data_stage_2__3504_, data_stage_2__3503_, data_stage_2__3502_, data_stage_2__3501_, data_stage_2__3500_, data_stage_2__3499_, data_stage_2__3498_, data_stage_2__3497_, data_stage_2__3496_, data_stage_2__3495_, data_stage_2__3494_, data_stage_2__3493_, data_stage_2__3492_, data_stage_2__3491_, data_stage_2__3490_, data_stage_2__3489_, data_stage_2__3488_, data_stage_2__3487_, data_stage_2__3486_, data_stage_2__3485_, data_stage_2__3484_, data_stage_2__3483_, data_stage_2__3482_, data_stage_2__3481_, data_stage_2__3480_, data_stage_2__3479_, data_stage_2__3478_, data_stage_2__3477_, data_stage_2__3476_, data_stage_2__3475_, data_stage_2__3474_, data_stage_2__3473_, data_stage_2__3472_, data_stage_2__3471_, data_stage_2__3470_, data_stage_2__3469_, data_stage_2__3468_, data_stage_2__3467_, data_stage_2__3466_, data_stage_2__3465_, data_stage_2__3464_, data_stage_2__3463_, data_stage_2__3462_, data_stage_2__3461_, data_stage_2__3460_, data_stage_2__3459_, data_stage_2__3458_, data_stage_2__3457_, data_stage_2__3456_, data_stage_2__3455_, data_stage_2__3454_, data_stage_2__3453_, data_stage_2__3452_, data_stage_2__3451_, data_stage_2__3450_, data_stage_2__3449_, data_stage_2__3448_, data_stage_2__3447_, data_stage_2__3446_, data_stage_2__3445_, data_stage_2__3444_, data_stage_2__3443_, data_stage_2__3442_, data_stage_2__3441_, data_stage_2__3440_, data_stage_2__3439_, data_stage_2__3438_, data_stage_2__3437_, data_stage_2__3436_, data_stage_2__3435_, data_stage_2__3434_, data_stage_2__3433_, data_stage_2__3432_, data_stage_2__3431_, data_stage_2__3430_, data_stage_2__3429_, data_stage_2__3428_, data_stage_2__3427_, data_stage_2__3426_, data_stage_2__3425_, data_stage_2__3424_, data_stage_2__3423_, data_stage_2__3422_, data_stage_2__3421_, data_stage_2__3420_, data_stage_2__3419_, data_stage_2__3418_, data_stage_2__3417_, data_stage_2__3416_, data_stage_2__3415_, data_stage_2__3414_, data_stage_2__3413_, data_stage_2__3412_, data_stage_2__3411_, data_stage_2__3410_, data_stage_2__3409_, data_stage_2__3408_, data_stage_2__3407_, data_stage_2__3406_, data_stage_2__3405_, data_stage_2__3404_, data_stage_2__3403_, data_stage_2__3402_, data_stage_2__3401_, data_stage_2__3400_, data_stage_2__3399_, data_stage_2__3398_, data_stage_2__3397_, data_stage_2__3396_, data_stage_2__3395_, data_stage_2__3394_, data_stage_2__3393_, data_stage_2__3392_, data_stage_2__3391_, data_stage_2__3390_, data_stage_2__3389_, data_stage_2__3388_, data_stage_2__3387_, data_stage_2__3386_, data_stage_2__3385_, data_stage_2__3384_, data_stage_2__3383_, data_stage_2__3382_, data_stage_2__3381_, data_stage_2__3380_, data_stage_2__3379_, data_stage_2__3378_, data_stage_2__3377_, data_stage_2__3376_, data_stage_2__3375_, data_stage_2__3374_, data_stage_2__3373_, data_stage_2__3372_, data_stage_2__3371_, data_stage_2__3370_, data_stage_2__3369_, data_stage_2__3368_, data_stage_2__3367_, data_stage_2__3366_, data_stage_2__3365_, data_stage_2__3364_, data_stage_2__3363_, data_stage_2__3362_, data_stage_2__3361_, data_stage_2__3360_, data_stage_2__3359_, data_stage_2__3358_, data_stage_2__3357_, data_stage_2__3356_, data_stage_2__3355_, data_stage_2__3354_, data_stage_2__3353_, data_stage_2__3352_, data_stage_2__3351_, data_stage_2__3350_, data_stage_2__3349_, data_stage_2__3348_, data_stage_2__3347_, data_stage_2__3346_, data_stage_2__3345_, data_stage_2__3344_, data_stage_2__3343_, data_stage_2__3342_, data_stage_2__3341_, data_stage_2__3340_, data_stage_2__3339_, data_stage_2__3338_, data_stage_2__3337_, data_stage_2__3336_, data_stage_2__3335_, data_stage_2__3334_, data_stage_2__3333_, data_stage_2__3332_, data_stage_2__3331_, data_stage_2__3330_, data_stage_2__3329_, data_stage_2__3328_, data_stage_2__3327_, data_stage_2__3326_, data_stage_2__3325_, data_stage_2__3324_, data_stage_2__3323_, data_stage_2__3322_, data_stage_2__3321_, data_stage_2__3320_, data_stage_2__3319_, data_stage_2__3318_, data_stage_2__3317_, data_stage_2__3316_, data_stage_2__3315_, data_stage_2__3314_, data_stage_2__3313_, data_stage_2__3312_, data_stage_2__3311_, data_stage_2__3310_, data_stage_2__3309_, data_stage_2__3308_, data_stage_2__3307_, data_stage_2__3306_, data_stage_2__3305_, data_stage_2__3304_, data_stage_2__3303_, data_stage_2__3302_, data_stage_2__3301_, data_stage_2__3300_, data_stage_2__3299_, data_stage_2__3298_, data_stage_2__3297_, data_stage_2__3296_, data_stage_2__3295_, data_stage_2__3294_, data_stage_2__3293_, data_stage_2__3292_, data_stage_2__3291_, data_stage_2__3290_, data_stage_2__3289_, data_stage_2__3288_, data_stage_2__3287_, data_stage_2__3286_, data_stage_2__3285_, data_stage_2__3284_, data_stage_2__3283_, data_stage_2__3282_, data_stage_2__3281_, data_stage_2__3280_, data_stage_2__3279_, data_stage_2__3278_, data_stage_2__3277_, data_stage_2__3276_, data_stage_2__3275_, data_stage_2__3274_, data_stage_2__3273_, data_stage_2__3272_, data_stage_2__3271_, data_stage_2__3270_, data_stage_2__3269_, data_stage_2__3268_, data_stage_2__3267_, data_stage_2__3266_, data_stage_2__3265_, data_stage_2__3264_, data_stage_2__3263_, data_stage_2__3262_, data_stage_2__3261_, data_stage_2__3260_, data_stage_2__3259_, data_stage_2__3258_, data_stage_2__3257_, data_stage_2__3256_, data_stage_2__3255_, data_stage_2__3254_, data_stage_2__3253_, data_stage_2__3252_, data_stage_2__3251_, data_stage_2__3250_, data_stage_2__3249_, data_stage_2__3248_, data_stage_2__3247_, data_stage_2__3246_, data_stage_2__3245_, data_stage_2__3244_, data_stage_2__3243_, data_stage_2__3242_, data_stage_2__3241_, data_stage_2__3240_, data_stage_2__3239_, data_stage_2__3238_, data_stage_2__3237_, data_stage_2__3236_, data_stage_2__3235_, data_stage_2__3234_, data_stage_2__3233_, data_stage_2__3232_, data_stage_2__3231_, data_stage_2__3230_, data_stage_2__3229_, data_stage_2__3228_, data_stage_2__3227_, data_stage_2__3226_, data_stage_2__3225_, data_stage_2__3224_, data_stage_2__3223_, data_stage_2__3222_, data_stage_2__3221_, data_stage_2__3220_, data_stage_2__3219_, data_stage_2__3218_, data_stage_2__3217_, data_stage_2__3216_, data_stage_2__3215_, data_stage_2__3214_, data_stage_2__3213_, data_stage_2__3212_, data_stage_2__3211_, data_stage_2__3210_, data_stage_2__3209_, data_stage_2__3208_, data_stage_2__3207_, data_stage_2__3206_, data_stage_2__3205_, data_stage_2__3204_, data_stage_2__3203_, data_stage_2__3202_, data_stage_2__3201_, data_stage_2__3200_, data_stage_2__3199_, data_stage_2__3198_, data_stage_2__3197_, data_stage_2__3196_, data_stage_2__3195_, data_stage_2__3194_, data_stage_2__3193_, data_stage_2__3192_, data_stage_2__3191_, data_stage_2__3190_, data_stage_2__3189_, data_stage_2__3188_, data_stage_2__3187_, data_stage_2__3186_, data_stage_2__3185_, data_stage_2__3184_, data_stage_2__3183_, data_stage_2__3182_, data_stage_2__3181_, data_stage_2__3180_, data_stage_2__3179_, data_stage_2__3178_, data_stage_2__3177_, data_stage_2__3176_, data_stage_2__3175_, data_stage_2__3174_, data_stage_2__3173_, data_stage_2__3172_, data_stage_2__3171_, data_stage_2__3170_, data_stage_2__3169_, data_stage_2__3168_, data_stage_2__3167_, data_stage_2__3166_, data_stage_2__3165_, data_stage_2__3164_, data_stage_2__3163_, data_stage_2__3162_, data_stage_2__3161_, data_stage_2__3160_, data_stage_2__3159_, data_stage_2__3158_, data_stage_2__3157_, data_stage_2__3156_, data_stage_2__3155_, data_stage_2__3154_, data_stage_2__3153_, data_stage_2__3152_, data_stage_2__3151_, data_stage_2__3150_, data_stage_2__3149_, data_stage_2__3148_, data_stage_2__3147_, data_stage_2__3146_, data_stage_2__3145_, data_stage_2__3144_, data_stage_2__3143_, data_stage_2__3142_, data_stage_2__3141_, data_stage_2__3140_, data_stage_2__3139_, data_stage_2__3138_, data_stage_2__3137_, data_stage_2__3136_, data_stage_2__3135_, data_stage_2__3134_, data_stage_2__3133_, data_stage_2__3132_, data_stage_2__3131_, data_stage_2__3130_, data_stage_2__3129_, data_stage_2__3128_, data_stage_2__3127_, data_stage_2__3126_, data_stage_2__3125_, data_stage_2__3124_, data_stage_2__3123_, data_stage_2__3122_, data_stage_2__3121_, data_stage_2__3120_, data_stage_2__3119_, data_stage_2__3118_, data_stage_2__3117_, data_stage_2__3116_, data_stage_2__3115_, data_stage_2__3114_, data_stage_2__3113_, data_stage_2__3112_, data_stage_2__3111_, data_stage_2__3110_, data_stage_2__3109_, data_stage_2__3108_, data_stage_2__3107_, data_stage_2__3106_, data_stage_2__3105_, data_stage_2__3104_, data_stage_2__3103_, data_stage_2__3102_, data_stage_2__3101_, data_stage_2__3100_, data_stage_2__3099_, data_stage_2__3098_, data_stage_2__3097_, data_stage_2__3096_, data_stage_2__3095_, data_stage_2__3094_, data_stage_2__3093_, data_stage_2__3092_, data_stage_2__3091_, data_stage_2__3090_, data_stage_2__3089_, data_stage_2__3088_, data_stage_2__3087_, data_stage_2__3086_, data_stage_2__3085_, data_stage_2__3084_, data_stage_2__3083_, data_stage_2__3082_, data_stage_2__3081_, data_stage_2__3080_, data_stage_2__3079_, data_stage_2__3078_, data_stage_2__3077_, data_stage_2__3076_, data_stage_2__3075_, data_stage_2__3074_, data_stage_2__3073_, data_stage_2__3072_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_7__swap_inst
  (
    .data_i({ data_stage_1__4095_, data_stage_1__4094_, data_stage_1__4093_, data_stage_1__4092_, data_stage_1__4091_, data_stage_1__4090_, data_stage_1__4089_, data_stage_1__4088_, data_stage_1__4087_, data_stage_1__4086_, data_stage_1__4085_, data_stage_1__4084_, data_stage_1__4083_, data_stage_1__4082_, data_stage_1__4081_, data_stage_1__4080_, data_stage_1__4079_, data_stage_1__4078_, data_stage_1__4077_, data_stage_1__4076_, data_stage_1__4075_, data_stage_1__4074_, data_stage_1__4073_, data_stage_1__4072_, data_stage_1__4071_, data_stage_1__4070_, data_stage_1__4069_, data_stage_1__4068_, data_stage_1__4067_, data_stage_1__4066_, data_stage_1__4065_, data_stage_1__4064_, data_stage_1__4063_, data_stage_1__4062_, data_stage_1__4061_, data_stage_1__4060_, data_stage_1__4059_, data_stage_1__4058_, data_stage_1__4057_, data_stage_1__4056_, data_stage_1__4055_, data_stage_1__4054_, data_stage_1__4053_, data_stage_1__4052_, data_stage_1__4051_, data_stage_1__4050_, data_stage_1__4049_, data_stage_1__4048_, data_stage_1__4047_, data_stage_1__4046_, data_stage_1__4045_, data_stage_1__4044_, data_stage_1__4043_, data_stage_1__4042_, data_stage_1__4041_, data_stage_1__4040_, data_stage_1__4039_, data_stage_1__4038_, data_stage_1__4037_, data_stage_1__4036_, data_stage_1__4035_, data_stage_1__4034_, data_stage_1__4033_, data_stage_1__4032_, data_stage_1__4031_, data_stage_1__4030_, data_stage_1__4029_, data_stage_1__4028_, data_stage_1__4027_, data_stage_1__4026_, data_stage_1__4025_, data_stage_1__4024_, data_stage_1__4023_, data_stage_1__4022_, data_stage_1__4021_, data_stage_1__4020_, data_stage_1__4019_, data_stage_1__4018_, data_stage_1__4017_, data_stage_1__4016_, data_stage_1__4015_, data_stage_1__4014_, data_stage_1__4013_, data_stage_1__4012_, data_stage_1__4011_, data_stage_1__4010_, data_stage_1__4009_, data_stage_1__4008_, data_stage_1__4007_, data_stage_1__4006_, data_stage_1__4005_, data_stage_1__4004_, data_stage_1__4003_, data_stage_1__4002_, data_stage_1__4001_, data_stage_1__4000_, data_stage_1__3999_, data_stage_1__3998_, data_stage_1__3997_, data_stage_1__3996_, data_stage_1__3995_, data_stage_1__3994_, data_stage_1__3993_, data_stage_1__3992_, data_stage_1__3991_, data_stage_1__3990_, data_stage_1__3989_, data_stage_1__3988_, data_stage_1__3987_, data_stage_1__3986_, data_stage_1__3985_, data_stage_1__3984_, data_stage_1__3983_, data_stage_1__3982_, data_stage_1__3981_, data_stage_1__3980_, data_stage_1__3979_, data_stage_1__3978_, data_stage_1__3977_, data_stage_1__3976_, data_stage_1__3975_, data_stage_1__3974_, data_stage_1__3973_, data_stage_1__3972_, data_stage_1__3971_, data_stage_1__3970_, data_stage_1__3969_, data_stage_1__3968_, data_stage_1__3967_, data_stage_1__3966_, data_stage_1__3965_, data_stage_1__3964_, data_stage_1__3963_, data_stage_1__3962_, data_stage_1__3961_, data_stage_1__3960_, data_stage_1__3959_, data_stage_1__3958_, data_stage_1__3957_, data_stage_1__3956_, data_stage_1__3955_, data_stage_1__3954_, data_stage_1__3953_, data_stage_1__3952_, data_stage_1__3951_, data_stage_1__3950_, data_stage_1__3949_, data_stage_1__3948_, data_stage_1__3947_, data_stage_1__3946_, data_stage_1__3945_, data_stage_1__3944_, data_stage_1__3943_, data_stage_1__3942_, data_stage_1__3941_, data_stage_1__3940_, data_stage_1__3939_, data_stage_1__3938_, data_stage_1__3937_, data_stage_1__3936_, data_stage_1__3935_, data_stage_1__3934_, data_stage_1__3933_, data_stage_1__3932_, data_stage_1__3931_, data_stage_1__3930_, data_stage_1__3929_, data_stage_1__3928_, data_stage_1__3927_, data_stage_1__3926_, data_stage_1__3925_, data_stage_1__3924_, data_stage_1__3923_, data_stage_1__3922_, data_stage_1__3921_, data_stage_1__3920_, data_stage_1__3919_, data_stage_1__3918_, data_stage_1__3917_, data_stage_1__3916_, data_stage_1__3915_, data_stage_1__3914_, data_stage_1__3913_, data_stage_1__3912_, data_stage_1__3911_, data_stage_1__3910_, data_stage_1__3909_, data_stage_1__3908_, data_stage_1__3907_, data_stage_1__3906_, data_stage_1__3905_, data_stage_1__3904_, data_stage_1__3903_, data_stage_1__3902_, data_stage_1__3901_, data_stage_1__3900_, data_stage_1__3899_, data_stage_1__3898_, data_stage_1__3897_, data_stage_1__3896_, data_stage_1__3895_, data_stage_1__3894_, data_stage_1__3893_, data_stage_1__3892_, data_stage_1__3891_, data_stage_1__3890_, data_stage_1__3889_, data_stage_1__3888_, data_stage_1__3887_, data_stage_1__3886_, data_stage_1__3885_, data_stage_1__3884_, data_stage_1__3883_, data_stage_1__3882_, data_stage_1__3881_, data_stage_1__3880_, data_stage_1__3879_, data_stage_1__3878_, data_stage_1__3877_, data_stage_1__3876_, data_stage_1__3875_, data_stage_1__3874_, data_stage_1__3873_, data_stage_1__3872_, data_stage_1__3871_, data_stage_1__3870_, data_stage_1__3869_, data_stage_1__3868_, data_stage_1__3867_, data_stage_1__3866_, data_stage_1__3865_, data_stage_1__3864_, data_stage_1__3863_, data_stage_1__3862_, data_stage_1__3861_, data_stage_1__3860_, data_stage_1__3859_, data_stage_1__3858_, data_stage_1__3857_, data_stage_1__3856_, data_stage_1__3855_, data_stage_1__3854_, data_stage_1__3853_, data_stage_1__3852_, data_stage_1__3851_, data_stage_1__3850_, data_stage_1__3849_, data_stage_1__3848_, data_stage_1__3847_, data_stage_1__3846_, data_stage_1__3845_, data_stage_1__3844_, data_stage_1__3843_, data_stage_1__3842_, data_stage_1__3841_, data_stage_1__3840_, data_stage_1__3839_, data_stage_1__3838_, data_stage_1__3837_, data_stage_1__3836_, data_stage_1__3835_, data_stage_1__3834_, data_stage_1__3833_, data_stage_1__3832_, data_stage_1__3831_, data_stage_1__3830_, data_stage_1__3829_, data_stage_1__3828_, data_stage_1__3827_, data_stage_1__3826_, data_stage_1__3825_, data_stage_1__3824_, data_stage_1__3823_, data_stage_1__3822_, data_stage_1__3821_, data_stage_1__3820_, data_stage_1__3819_, data_stage_1__3818_, data_stage_1__3817_, data_stage_1__3816_, data_stage_1__3815_, data_stage_1__3814_, data_stage_1__3813_, data_stage_1__3812_, data_stage_1__3811_, data_stage_1__3810_, data_stage_1__3809_, data_stage_1__3808_, data_stage_1__3807_, data_stage_1__3806_, data_stage_1__3805_, data_stage_1__3804_, data_stage_1__3803_, data_stage_1__3802_, data_stage_1__3801_, data_stage_1__3800_, data_stage_1__3799_, data_stage_1__3798_, data_stage_1__3797_, data_stage_1__3796_, data_stage_1__3795_, data_stage_1__3794_, data_stage_1__3793_, data_stage_1__3792_, data_stage_1__3791_, data_stage_1__3790_, data_stage_1__3789_, data_stage_1__3788_, data_stage_1__3787_, data_stage_1__3786_, data_stage_1__3785_, data_stage_1__3784_, data_stage_1__3783_, data_stage_1__3782_, data_stage_1__3781_, data_stage_1__3780_, data_stage_1__3779_, data_stage_1__3778_, data_stage_1__3777_, data_stage_1__3776_, data_stage_1__3775_, data_stage_1__3774_, data_stage_1__3773_, data_stage_1__3772_, data_stage_1__3771_, data_stage_1__3770_, data_stage_1__3769_, data_stage_1__3768_, data_stage_1__3767_, data_stage_1__3766_, data_stage_1__3765_, data_stage_1__3764_, data_stage_1__3763_, data_stage_1__3762_, data_stage_1__3761_, data_stage_1__3760_, data_stage_1__3759_, data_stage_1__3758_, data_stage_1__3757_, data_stage_1__3756_, data_stage_1__3755_, data_stage_1__3754_, data_stage_1__3753_, data_stage_1__3752_, data_stage_1__3751_, data_stage_1__3750_, data_stage_1__3749_, data_stage_1__3748_, data_stage_1__3747_, data_stage_1__3746_, data_stage_1__3745_, data_stage_1__3744_, data_stage_1__3743_, data_stage_1__3742_, data_stage_1__3741_, data_stage_1__3740_, data_stage_1__3739_, data_stage_1__3738_, data_stage_1__3737_, data_stage_1__3736_, data_stage_1__3735_, data_stage_1__3734_, data_stage_1__3733_, data_stage_1__3732_, data_stage_1__3731_, data_stage_1__3730_, data_stage_1__3729_, data_stage_1__3728_, data_stage_1__3727_, data_stage_1__3726_, data_stage_1__3725_, data_stage_1__3724_, data_stage_1__3723_, data_stage_1__3722_, data_stage_1__3721_, data_stage_1__3720_, data_stage_1__3719_, data_stage_1__3718_, data_stage_1__3717_, data_stage_1__3716_, data_stage_1__3715_, data_stage_1__3714_, data_stage_1__3713_, data_stage_1__3712_, data_stage_1__3711_, data_stage_1__3710_, data_stage_1__3709_, data_stage_1__3708_, data_stage_1__3707_, data_stage_1__3706_, data_stage_1__3705_, data_stage_1__3704_, data_stage_1__3703_, data_stage_1__3702_, data_stage_1__3701_, data_stage_1__3700_, data_stage_1__3699_, data_stage_1__3698_, data_stage_1__3697_, data_stage_1__3696_, data_stage_1__3695_, data_stage_1__3694_, data_stage_1__3693_, data_stage_1__3692_, data_stage_1__3691_, data_stage_1__3690_, data_stage_1__3689_, data_stage_1__3688_, data_stage_1__3687_, data_stage_1__3686_, data_stage_1__3685_, data_stage_1__3684_, data_stage_1__3683_, data_stage_1__3682_, data_stage_1__3681_, data_stage_1__3680_, data_stage_1__3679_, data_stage_1__3678_, data_stage_1__3677_, data_stage_1__3676_, data_stage_1__3675_, data_stage_1__3674_, data_stage_1__3673_, data_stage_1__3672_, data_stage_1__3671_, data_stage_1__3670_, data_stage_1__3669_, data_stage_1__3668_, data_stage_1__3667_, data_stage_1__3666_, data_stage_1__3665_, data_stage_1__3664_, data_stage_1__3663_, data_stage_1__3662_, data_stage_1__3661_, data_stage_1__3660_, data_stage_1__3659_, data_stage_1__3658_, data_stage_1__3657_, data_stage_1__3656_, data_stage_1__3655_, data_stage_1__3654_, data_stage_1__3653_, data_stage_1__3652_, data_stage_1__3651_, data_stage_1__3650_, data_stage_1__3649_, data_stage_1__3648_, data_stage_1__3647_, data_stage_1__3646_, data_stage_1__3645_, data_stage_1__3644_, data_stage_1__3643_, data_stage_1__3642_, data_stage_1__3641_, data_stage_1__3640_, data_stage_1__3639_, data_stage_1__3638_, data_stage_1__3637_, data_stage_1__3636_, data_stage_1__3635_, data_stage_1__3634_, data_stage_1__3633_, data_stage_1__3632_, data_stage_1__3631_, data_stage_1__3630_, data_stage_1__3629_, data_stage_1__3628_, data_stage_1__3627_, data_stage_1__3626_, data_stage_1__3625_, data_stage_1__3624_, data_stage_1__3623_, data_stage_1__3622_, data_stage_1__3621_, data_stage_1__3620_, data_stage_1__3619_, data_stage_1__3618_, data_stage_1__3617_, data_stage_1__3616_, data_stage_1__3615_, data_stage_1__3614_, data_stage_1__3613_, data_stage_1__3612_, data_stage_1__3611_, data_stage_1__3610_, data_stage_1__3609_, data_stage_1__3608_, data_stage_1__3607_, data_stage_1__3606_, data_stage_1__3605_, data_stage_1__3604_, data_stage_1__3603_, data_stage_1__3602_, data_stage_1__3601_, data_stage_1__3600_, data_stage_1__3599_, data_stage_1__3598_, data_stage_1__3597_, data_stage_1__3596_, data_stage_1__3595_, data_stage_1__3594_, data_stage_1__3593_, data_stage_1__3592_, data_stage_1__3591_, data_stage_1__3590_, data_stage_1__3589_, data_stage_1__3588_, data_stage_1__3587_, data_stage_1__3586_, data_stage_1__3585_, data_stage_1__3584_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__4095_, data_stage_2__4094_, data_stage_2__4093_, data_stage_2__4092_, data_stage_2__4091_, data_stage_2__4090_, data_stage_2__4089_, data_stage_2__4088_, data_stage_2__4087_, data_stage_2__4086_, data_stage_2__4085_, data_stage_2__4084_, data_stage_2__4083_, data_stage_2__4082_, data_stage_2__4081_, data_stage_2__4080_, data_stage_2__4079_, data_stage_2__4078_, data_stage_2__4077_, data_stage_2__4076_, data_stage_2__4075_, data_stage_2__4074_, data_stage_2__4073_, data_stage_2__4072_, data_stage_2__4071_, data_stage_2__4070_, data_stage_2__4069_, data_stage_2__4068_, data_stage_2__4067_, data_stage_2__4066_, data_stage_2__4065_, data_stage_2__4064_, data_stage_2__4063_, data_stage_2__4062_, data_stage_2__4061_, data_stage_2__4060_, data_stage_2__4059_, data_stage_2__4058_, data_stage_2__4057_, data_stage_2__4056_, data_stage_2__4055_, data_stage_2__4054_, data_stage_2__4053_, data_stage_2__4052_, data_stage_2__4051_, data_stage_2__4050_, data_stage_2__4049_, data_stage_2__4048_, data_stage_2__4047_, data_stage_2__4046_, data_stage_2__4045_, data_stage_2__4044_, data_stage_2__4043_, data_stage_2__4042_, data_stage_2__4041_, data_stage_2__4040_, data_stage_2__4039_, data_stage_2__4038_, data_stage_2__4037_, data_stage_2__4036_, data_stage_2__4035_, data_stage_2__4034_, data_stage_2__4033_, data_stage_2__4032_, data_stage_2__4031_, data_stage_2__4030_, data_stage_2__4029_, data_stage_2__4028_, data_stage_2__4027_, data_stage_2__4026_, data_stage_2__4025_, data_stage_2__4024_, data_stage_2__4023_, data_stage_2__4022_, data_stage_2__4021_, data_stage_2__4020_, data_stage_2__4019_, data_stage_2__4018_, data_stage_2__4017_, data_stage_2__4016_, data_stage_2__4015_, data_stage_2__4014_, data_stage_2__4013_, data_stage_2__4012_, data_stage_2__4011_, data_stage_2__4010_, data_stage_2__4009_, data_stage_2__4008_, data_stage_2__4007_, data_stage_2__4006_, data_stage_2__4005_, data_stage_2__4004_, data_stage_2__4003_, data_stage_2__4002_, data_stage_2__4001_, data_stage_2__4000_, data_stage_2__3999_, data_stage_2__3998_, data_stage_2__3997_, data_stage_2__3996_, data_stage_2__3995_, data_stage_2__3994_, data_stage_2__3993_, data_stage_2__3992_, data_stage_2__3991_, data_stage_2__3990_, data_stage_2__3989_, data_stage_2__3988_, data_stage_2__3987_, data_stage_2__3986_, data_stage_2__3985_, data_stage_2__3984_, data_stage_2__3983_, data_stage_2__3982_, data_stage_2__3981_, data_stage_2__3980_, data_stage_2__3979_, data_stage_2__3978_, data_stage_2__3977_, data_stage_2__3976_, data_stage_2__3975_, data_stage_2__3974_, data_stage_2__3973_, data_stage_2__3972_, data_stage_2__3971_, data_stage_2__3970_, data_stage_2__3969_, data_stage_2__3968_, data_stage_2__3967_, data_stage_2__3966_, data_stage_2__3965_, data_stage_2__3964_, data_stage_2__3963_, data_stage_2__3962_, data_stage_2__3961_, data_stage_2__3960_, data_stage_2__3959_, data_stage_2__3958_, data_stage_2__3957_, data_stage_2__3956_, data_stage_2__3955_, data_stage_2__3954_, data_stage_2__3953_, data_stage_2__3952_, data_stage_2__3951_, data_stage_2__3950_, data_stage_2__3949_, data_stage_2__3948_, data_stage_2__3947_, data_stage_2__3946_, data_stage_2__3945_, data_stage_2__3944_, data_stage_2__3943_, data_stage_2__3942_, data_stage_2__3941_, data_stage_2__3940_, data_stage_2__3939_, data_stage_2__3938_, data_stage_2__3937_, data_stage_2__3936_, data_stage_2__3935_, data_stage_2__3934_, data_stage_2__3933_, data_stage_2__3932_, data_stage_2__3931_, data_stage_2__3930_, data_stage_2__3929_, data_stage_2__3928_, data_stage_2__3927_, data_stage_2__3926_, data_stage_2__3925_, data_stage_2__3924_, data_stage_2__3923_, data_stage_2__3922_, data_stage_2__3921_, data_stage_2__3920_, data_stage_2__3919_, data_stage_2__3918_, data_stage_2__3917_, data_stage_2__3916_, data_stage_2__3915_, data_stage_2__3914_, data_stage_2__3913_, data_stage_2__3912_, data_stage_2__3911_, data_stage_2__3910_, data_stage_2__3909_, data_stage_2__3908_, data_stage_2__3907_, data_stage_2__3906_, data_stage_2__3905_, data_stage_2__3904_, data_stage_2__3903_, data_stage_2__3902_, data_stage_2__3901_, data_stage_2__3900_, data_stage_2__3899_, data_stage_2__3898_, data_stage_2__3897_, data_stage_2__3896_, data_stage_2__3895_, data_stage_2__3894_, data_stage_2__3893_, data_stage_2__3892_, data_stage_2__3891_, data_stage_2__3890_, data_stage_2__3889_, data_stage_2__3888_, data_stage_2__3887_, data_stage_2__3886_, data_stage_2__3885_, data_stage_2__3884_, data_stage_2__3883_, data_stage_2__3882_, data_stage_2__3881_, data_stage_2__3880_, data_stage_2__3879_, data_stage_2__3878_, data_stage_2__3877_, data_stage_2__3876_, data_stage_2__3875_, data_stage_2__3874_, data_stage_2__3873_, data_stage_2__3872_, data_stage_2__3871_, data_stage_2__3870_, data_stage_2__3869_, data_stage_2__3868_, data_stage_2__3867_, data_stage_2__3866_, data_stage_2__3865_, data_stage_2__3864_, data_stage_2__3863_, data_stage_2__3862_, data_stage_2__3861_, data_stage_2__3860_, data_stage_2__3859_, data_stage_2__3858_, data_stage_2__3857_, data_stage_2__3856_, data_stage_2__3855_, data_stage_2__3854_, data_stage_2__3853_, data_stage_2__3852_, data_stage_2__3851_, data_stage_2__3850_, data_stage_2__3849_, data_stage_2__3848_, data_stage_2__3847_, data_stage_2__3846_, data_stage_2__3845_, data_stage_2__3844_, data_stage_2__3843_, data_stage_2__3842_, data_stage_2__3841_, data_stage_2__3840_, data_stage_2__3839_, data_stage_2__3838_, data_stage_2__3837_, data_stage_2__3836_, data_stage_2__3835_, data_stage_2__3834_, data_stage_2__3833_, data_stage_2__3832_, data_stage_2__3831_, data_stage_2__3830_, data_stage_2__3829_, data_stage_2__3828_, data_stage_2__3827_, data_stage_2__3826_, data_stage_2__3825_, data_stage_2__3824_, data_stage_2__3823_, data_stage_2__3822_, data_stage_2__3821_, data_stage_2__3820_, data_stage_2__3819_, data_stage_2__3818_, data_stage_2__3817_, data_stage_2__3816_, data_stage_2__3815_, data_stage_2__3814_, data_stage_2__3813_, data_stage_2__3812_, data_stage_2__3811_, data_stage_2__3810_, data_stage_2__3809_, data_stage_2__3808_, data_stage_2__3807_, data_stage_2__3806_, data_stage_2__3805_, data_stage_2__3804_, data_stage_2__3803_, data_stage_2__3802_, data_stage_2__3801_, data_stage_2__3800_, data_stage_2__3799_, data_stage_2__3798_, data_stage_2__3797_, data_stage_2__3796_, data_stage_2__3795_, data_stage_2__3794_, data_stage_2__3793_, data_stage_2__3792_, data_stage_2__3791_, data_stage_2__3790_, data_stage_2__3789_, data_stage_2__3788_, data_stage_2__3787_, data_stage_2__3786_, data_stage_2__3785_, data_stage_2__3784_, data_stage_2__3783_, data_stage_2__3782_, data_stage_2__3781_, data_stage_2__3780_, data_stage_2__3779_, data_stage_2__3778_, data_stage_2__3777_, data_stage_2__3776_, data_stage_2__3775_, data_stage_2__3774_, data_stage_2__3773_, data_stage_2__3772_, data_stage_2__3771_, data_stage_2__3770_, data_stage_2__3769_, data_stage_2__3768_, data_stage_2__3767_, data_stage_2__3766_, data_stage_2__3765_, data_stage_2__3764_, data_stage_2__3763_, data_stage_2__3762_, data_stage_2__3761_, data_stage_2__3760_, data_stage_2__3759_, data_stage_2__3758_, data_stage_2__3757_, data_stage_2__3756_, data_stage_2__3755_, data_stage_2__3754_, data_stage_2__3753_, data_stage_2__3752_, data_stage_2__3751_, data_stage_2__3750_, data_stage_2__3749_, data_stage_2__3748_, data_stage_2__3747_, data_stage_2__3746_, data_stage_2__3745_, data_stage_2__3744_, data_stage_2__3743_, data_stage_2__3742_, data_stage_2__3741_, data_stage_2__3740_, data_stage_2__3739_, data_stage_2__3738_, data_stage_2__3737_, data_stage_2__3736_, data_stage_2__3735_, data_stage_2__3734_, data_stage_2__3733_, data_stage_2__3732_, data_stage_2__3731_, data_stage_2__3730_, data_stage_2__3729_, data_stage_2__3728_, data_stage_2__3727_, data_stage_2__3726_, data_stage_2__3725_, data_stage_2__3724_, data_stage_2__3723_, data_stage_2__3722_, data_stage_2__3721_, data_stage_2__3720_, data_stage_2__3719_, data_stage_2__3718_, data_stage_2__3717_, data_stage_2__3716_, data_stage_2__3715_, data_stage_2__3714_, data_stage_2__3713_, data_stage_2__3712_, data_stage_2__3711_, data_stage_2__3710_, data_stage_2__3709_, data_stage_2__3708_, data_stage_2__3707_, data_stage_2__3706_, data_stage_2__3705_, data_stage_2__3704_, data_stage_2__3703_, data_stage_2__3702_, data_stage_2__3701_, data_stage_2__3700_, data_stage_2__3699_, data_stage_2__3698_, data_stage_2__3697_, data_stage_2__3696_, data_stage_2__3695_, data_stage_2__3694_, data_stage_2__3693_, data_stage_2__3692_, data_stage_2__3691_, data_stage_2__3690_, data_stage_2__3689_, data_stage_2__3688_, data_stage_2__3687_, data_stage_2__3686_, data_stage_2__3685_, data_stage_2__3684_, data_stage_2__3683_, data_stage_2__3682_, data_stage_2__3681_, data_stage_2__3680_, data_stage_2__3679_, data_stage_2__3678_, data_stage_2__3677_, data_stage_2__3676_, data_stage_2__3675_, data_stage_2__3674_, data_stage_2__3673_, data_stage_2__3672_, data_stage_2__3671_, data_stage_2__3670_, data_stage_2__3669_, data_stage_2__3668_, data_stage_2__3667_, data_stage_2__3666_, data_stage_2__3665_, data_stage_2__3664_, data_stage_2__3663_, data_stage_2__3662_, data_stage_2__3661_, data_stage_2__3660_, data_stage_2__3659_, data_stage_2__3658_, data_stage_2__3657_, data_stage_2__3656_, data_stage_2__3655_, data_stage_2__3654_, data_stage_2__3653_, data_stage_2__3652_, data_stage_2__3651_, data_stage_2__3650_, data_stage_2__3649_, data_stage_2__3648_, data_stage_2__3647_, data_stage_2__3646_, data_stage_2__3645_, data_stage_2__3644_, data_stage_2__3643_, data_stage_2__3642_, data_stage_2__3641_, data_stage_2__3640_, data_stage_2__3639_, data_stage_2__3638_, data_stage_2__3637_, data_stage_2__3636_, data_stage_2__3635_, data_stage_2__3634_, data_stage_2__3633_, data_stage_2__3632_, data_stage_2__3631_, data_stage_2__3630_, data_stage_2__3629_, data_stage_2__3628_, data_stage_2__3627_, data_stage_2__3626_, data_stage_2__3625_, data_stage_2__3624_, data_stage_2__3623_, data_stage_2__3622_, data_stage_2__3621_, data_stage_2__3620_, data_stage_2__3619_, data_stage_2__3618_, data_stage_2__3617_, data_stage_2__3616_, data_stage_2__3615_, data_stage_2__3614_, data_stage_2__3613_, data_stage_2__3612_, data_stage_2__3611_, data_stage_2__3610_, data_stage_2__3609_, data_stage_2__3608_, data_stage_2__3607_, data_stage_2__3606_, data_stage_2__3605_, data_stage_2__3604_, data_stage_2__3603_, data_stage_2__3602_, data_stage_2__3601_, data_stage_2__3600_, data_stage_2__3599_, data_stage_2__3598_, data_stage_2__3597_, data_stage_2__3596_, data_stage_2__3595_, data_stage_2__3594_, data_stage_2__3593_, data_stage_2__3592_, data_stage_2__3591_, data_stage_2__3590_, data_stage_2__3589_, data_stage_2__3588_, data_stage_2__3587_, data_stage_2__3586_, data_stage_2__3585_, data_stage_2__3584_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_8__swap_inst
  (
    .data_i({ data_stage_1__4607_, data_stage_1__4606_, data_stage_1__4605_, data_stage_1__4604_, data_stage_1__4603_, data_stage_1__4602_, data_stage_1__4601_, data_stage_1__4600_, data_stage_1__4599_, data_stage_1__4598_, data_stage_1__4597_, data_stage_1__4596_, data_stage_1__4595_, data_stage_1__4594_, data_stage_1__4593_, data_stage_1__4592_, data_stage_1__4591_, data_stage_1__4590_, data_stage_1__4589_, data_stage_1__4588_, data_stage_1__4587_, data_stage_1__4586_, data_stage_1__4585_, data_stage_1__4584_, data_stage_1__4583_, data_stage_1__4582_, data_stage_1__4581_, data_stage_1__4580_, data_stage_1__4579_, data_stage_1__4578_, data_stage_1__4577_, data_stage_1__4576_, data_stage_1__4575_, data_stage_1__4574_, data_stage_1__4573_, data_stage_1__4572_, data_stage_1__4571_, data_stage_1__4570_, data_stage_1__4569_, data_stage_1__4568_, data_stage_1__4567_, data_stage_1__4566_, data_stage_1__4565_, data_stage_1__4564_, data_stage_1__4563_, data_stage_1__4562_, data_stage_1__4561_, data_stage_1__4560_, data_stage_1__4559_, data_stage_1__4558_, data_stage_1__4557_, data_stage_1__4556_, data_stage_1__4555_, data_stage_1__4554_, data_stage_1__4553_, data_stage_1__4552_, data_stage_1__4551_, data_stage_1__4550_, data_stage_1__4549_, data_stage_1__4548_, data_stage_1__4547_, data_stage_1__4546_, data_stage_1__4545_, data_stage_1__4544_, data_stage_1__4543_, data_stage_1__4542_, data_stage_1__4541_, data_stage_1__4540_, data_stage_1__4539_, data_stage_1__4538_, data_stage_1__4537_, data_stage_1__4536_, data_stage_1__4535_, data_stage_1__4534_, data_stage_1__4533_, data_stage_1__4532_, data_stage_1__4531_, data_stage_1__4530_, data_stage_1__4529_, data_stage_1__4528_, data_stage_1__4527_, data_stage_1__4526_, data_stage_1__4525_, data_stage_1__4524_, data_stage_1__4523_, data_stage_1__4522_, data_stage_1__4521_, data_stage_1__4520_, data_stage_1__4519_, data_stage_1__4518_, data_stage_1__4517_, data_stage_1__4516_, data_stage_1__4515_, data_stage_1__4514_, data_stage_1__4513_, data_stage_1__4512_, data_stage_1__4511_, data_stage_1__4510_, data_stage_1__4509_, data_stage_1__4508_, data_stage_1__4507_, data_stage_1__4506_, data_stage_1__4505_, data_stage_1__4504_, data_stage_1__4503_, data_stage_1__4502_, data_stage_1__4501_, data_stage_1__4500_, data_stage_1__4499_, data_stage_1__4498_, data_stage_1__4497_, data_stage_1__4496_, data_stage_1__4495_, data_stage_1__4494_, data_stage_1__4493_, data_stage_1__4492_, data_stage_1__4491_, data_stage_1__4490_, data_stage_1__4489_, data_stage_1__4488_, data_stage_1__4487_, data_stage_1__4486_, data_stage_1__4485_, data_stage_1__4484_, data_stage_1__4483_, data_stage_1__4482_, data_stage_1__4481_, data_stage_1__4480_, data_stage_1__4479_, data_stage_1__4478_, data_stage_1__4477_, data_stage_1__4476_, data_stage_1__4475_, data_stage_1__4474_, data_stage_1__4473_, data_stage_1__4472_, data_stage_1__4471_, data_stage_1__4470_, data_stage_1__4469_, data_stage_1__4468_, data_stage_1__4467_, data_stage_1__4466_, data_stage_1__4465_, data_stage_1__4464_, data_stage_1__4463_, data_stage_1__4462_, data_stage_1__4461_, data_stage_1__4460_, data_stage_1__4459_, data_stage_1__4458_, data_stage_1__4457_, data_stage_1__4456_, data_stage_1__4455_, data_stage_1__4454_, data_stage_1__4453_, data_stage_1__4452_, data_stage_1__4451_, data_stage_1__4450_, data_stage_1__4449_, data_stage_1__4448_, data_stage_1__4447_, data_stage_1__4446_, data_stage_1__4445_, data_stage_1__4444_, data_stage_1__4443_, data_stage_1__4442_, data_stage_1__4441_, data_stage_1__4440_, data_stage_1__4439_, data_stage_1__4438_, data_stage_1__4437_, data_stage_1__4436_, data_stage_1__4435_, data_stage_1__4434_, data_stage_1__4433_, data_stage_1__4432_, data_stage_1__4431_, data_stage_1__4430_, data_stage_1__4429_, data_stage_1__4428_, data_stage_1__4427_, data_stage_1__4426_, data_stage_1__4425_, data_stage_1__4424_, data_stage_1__4423_, data_stage_1__4422_, data_stage_1__4421_, data_stage_1__4420_, data_stage_1__4419_, data_stage_1__4418_, data_stage_1__4417_, data_stage_1__4416_, data_stage_1__4415_, data_stage_1__4414_, data_stage_1__4413_, data_stage_1__4412_, data_stage_1__4411_, data_stage_1__4410_, data_stage_1__4409_, data_stage_1__4408_, data_stage_1__4407_, data_stage_1__4406_, data_stage_1__4405_, data_stage_1__4404_, data_stage_1__4403_, data_stage_1__4402_, data_stage_1__4401_, data_stage_1__4400_, data_stage_1__4399_, data_stage_1__4398_, data_stage_1__4397_, data_stage_1__4396_, data_stage_1__4395_, data_stage_1__4394_, data_stage_1__4393_, data_stage_1__4392_, data_stage_1__4391_, data_stage_1__4390_, data_stage_1__4389_, data_stage_1__4388_, data_stage_1__4387_, data_stage_1__4386_, data_stage_1__4385_, data_stage_1__4384_, data_stage_1__4383_, data_stage_1__4382_, data_stage_1__4381_, data_stage_1__4380_, data_stage_1__4379_, data_stage_1__4378_, data_stage_1__4377_, data_stage_1__4376_, data_stage_1__4375_, data_stage_1__4374_, data_stage_1__4373_, data_stage_1__4372_, data_stage_1__4371_, data_stage_1__4370_, data_stage_1__4369_, data_stage_1__4368_, data_stage_1__4367_, data_stage_1__4366_, data_stage_1__4365_, data_stage_1__4364_, data_stage_1__4363_, data_stage_1__4362_, data_stage_1__4361_, data_stage_1__4360_, data_stage_1__4359_, data_stage_1__4358_, data_stage_1__4357_, data_stage_1__4356_, data_stage_1__4355_, data_stage_1__4354_, data_stage_1__4353_, data_stage_1__4352_, data_stage_1__4351_, data_stage_1__4350_, data_stage_1__4349_, data_stage_1__4348_, data_stage_1__4347_, data_stage_1__4346_, data_stage_1__4345_, data_stage_1__4344_, data_stage_1__4343_, data_stage_1__4342_, data_stage_1__4341_, data_stage_1__4340_, data_stage_1__4339_, data_stage_1__4338_, data_stage_1__4337_, data_stage_1__4336_, data_stage_1__4335_, data_stage_1__4334_, data_stage_1__4333_, data_stage_1__4332_, data_stage_1__4331_, data_stage_1__4330_, data_stage_1__4329_, data_stage_1__4328_, data_stage_1__4327_, data_stage_1__4326_, data_stage_1__4325_, data_stage_1__4324_, data_stage_1__4323_, data_stage_1__4322_, data_stage_1__4321_, data_stage_1__4320_, data_stage_1__4319_, data_stage_1__4318_, data_stage_1__4317_, data_stage_1__4316_, data_stage_1__4315_, data_stage_1__4314_, data_stage_1__4313_, data_stage_1__4312_, data_stage_1__4311_, data_stage_1__4310_, data_stage_1__4309_, data_stage_1__4308_, data_stage_1__4307_, data_stage_1__4306_, data_stage_1__4305_, data_stage_1__4304_, data_stage_1__4303_, data_stage_1__4302_, data_stage_1__4301_, data_stage_1__4300_, data_stage_1__4299_, data_stage_1__4298_, data_stage_1__4297_, data_stage_1__4296_, data_stage_1__4295_, data_stage_1__4294_, data_stage_1__4293_, data_stage_1__4292_, data_stage_1__4291_, data_stage_1__4290_, data_stage_1__4289_, data_stage_1__4288_, data_stage_1__4287_, data_stage_1__4286_, data_stage_1__4285_, data_stage_1__4284_, data_stage_1__4283_, data_stage_1__4282_, data_stage_1__4281_, data_stage_1__4280_, data_stage_1__4279_, data_stage_1__4278_, data_stage_1__4277_, data_stage_1__4276_, data_stage_1__4275_, data_stage_1__4274_, data_stage_1__4273_, data_stage_1__4272_, data_stage_1__4271_, data_stage_1__4270_, data_stage_1__4269_, data_stage_1__4268_, data_stage_1__4267_, data_stage_1__4266_, data_stage_1__4265_, data_stage_1__4264_, data_stage_1__4263_, data_stage_1__4262_, data_stage_1__4261_, data_stage_1__4260_, data_stage_1__4259_, data_stage_1__4258_, data_stage_1__4257_, data_stage_1__4256_, data_stage_1__4255_, data_stage_1__4254_, data_stage_1__4253_, data_stage_1__4252_, data_stage_1__4251_, data_stage_1__4250_, data_stage_1__4249_, data_stage_1__4248_, data_stage_1__4247_, data_stage_1__4246_, data_stage_1__4245_, data_stage_1__4244_, data_stage_1__4243_, data_stage_1__4242_, data_stage_1__4241_, data_stage_1__4240_, data_stage_1__4239_, data_stage_1__4238_, data_stage_1__4237_, data_stage_1__4236_, data_stage_1__4235_, data_stage_1__4234_, data_stage_1__4233_, data_stage_1__4232_, data_stage_1__4231_, data_stage_1__4230_, data_stage_1__4229_, data_stage_1__4228_, data_stage_1__4227_, data_stage_1__4226_, data_stage_1__4225_, data_stage_1__4224_, data_stage_1__4223_, data_stage_1__4222_, data_stage_1__4221_, data_stage_1__4220_, data_stage_1__4219_, data_stage_1__4218_, data_stage_1__4217_, data_stage_1__4216_, data_stage_1__4215_, data_stage_1__4214_, data_stage_1__4213_, data_stage_1__4212_, data_stage_1__4211_, data_stage_1__4210_, data_stage_1__4209_, data_stage_1__4208_, data_stage_1__4207_, data_stage_1__4206_, data_stage_1__4205_, data_stage_1__4204_, data_stage_1__4203_, data_stage_1__4202_, data_stage_1__4201_, data_stage_1__4200_, data_stage_1__4199_, data_stage_1__4198_, data_stage_1__4197_, data_stage_1__4196_, data_stage_1__4195_, data_stage_1__4194_, data_stage_1__4193_, data_stage_1__4192_, data_stage_1__4191_, data_stage_1__4190_, data_stage_1__4189_, data_stage_1__4188_, data_stage_1__4187_, data_stage_1__4186_, data_stage_1__4185_, data_stage_1__4184_, data_stage_1__4183_, data_stage_1__4182_, data_stage_1__4181_, data_stage_1__4180_, data_stage_1__4179_, data_stage_1__4178_, data_stage_1__4177_, data_stage_1__4176_, data_stage_1__4175_, data_stage_1__4174_, data_stage_1__4173_, data_stage_1__4172_, data_stage_1__4171_, data_stage_1__4170_, data_stage_1__4169_, data_stage_1__4168_, data_stage_1__4167_, data_stage_1__4166_, data_stage_1__4165_, data_stage_1__4164_, data_stage_1__4163_, data_stage_1__4162_, data_stage_1__4161_, data_stage_1__4160_, data_stage_1__4159_, data_stage_1__4158_, data_stage_1__4157_, data_stage_1__4156_, data_stage_1__4155_, data_stage_1__4154_, data_stage_1__4153_, data_stage_1__4152_, data_stage_1__4151_, data_stage_1__4150_, data_stage_1__4149_, data_stage_1__4148_, data_stage_1__4147_, data_stage_1__4146_, data_stage_1__4145_, data_stage_1__4144_, data_stage_1__4143_, data_stage_1__4142_, data_stage_1__4141_, data_stage_1__4140_, data_stage_1__4139_, data_stage_1__4138_, data_stage_1__4137_, data_stage_1__4136_, data_stage_1__4135_, data_stage_1__4134_, data_stage_1__4133_, data_stage_1__4132_, data_stage_1__4131_, data_stage_1__4130_, data_stage_1__4129_, data_stage_1__4128_, data_stage_1__4127_, data_stage_1__4126_, data_stage_1__4125_, data_stage_1__4124_, data_stage_1__4123_, data_stage_1__4122_, data_stage_1__4121_, data_stage_1__4120_, data_stage_1__4119_, data_stage_1__4118_, data_stage_1__4117_, data_stage_1__4116_, data_stage_1__4115_, data_stage_1__4114_, data_stage_1__4113_, data_stage_1__4112_, data_stage_1__4111_, data_stage_1__4110_, data_stage_1__4109_, data_stage_1__4108_, data_stage_1__4107_, data_stage_1__4106_, data_stage_1__4105_, data_stage_1__4104_, data_stage_1__4103_, data_stage_1__4102_, data_stage_1__4101_, data_stage_1__4100_, data_stage_1__4099_, data_stage_1__4098_, data_stage_1__4097_, data_stage_1__4096_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__4607_, data_stage_2__4606_, data_stage_2__4605_, data_stage_2__4604_, data_stage_2__4603_, data_stage_2__4602_, data_stage_2__4601_, data_stage_2__4600_, data_stage_2__4599_, data_stage_2__4598_, data_stage_2__4597_, data_stage_2__4596_, data_stage_2__4595_, data_stage_2__4594_, data_stage_2__4593_, data_stage_2__4592_, data_stage_2__4591_, data_stage_2__4590_, data_stage_2__4589_, data_stage_2__4588_, data_stage_2__4587_, data_stage_2__4586_, data_stage_2__4585_, data_stage_2__4584_, data_stage_2__4583_, data_stage_2__4582_, data_stage_2__4581_, data_stage_2__4580_, data_stage_2__4579_, data_stage_2__4578_, data_stage_2__4577_, data_stage_2__4576_, data_stage_2__4575_, data_stage_2__4574_, data_stage_2__4573_, data_stage_2__4572_, data_stage_2__4571_, data_stage_2__4570_, data_stage_2__4569_, data_stage_2__4568_, data_stage_2__4567_, data_stage_2__4566_, data_stage_2__4565_, data_stage_2__4564_, data_stage_2__4563_, data_stage_2__4562_, data_stage_2__4561_, data_stage_2__4560_, data_stage_2__4559_, data_stage_2__4558_, data_stage_2__4557_, data_stage_2__4556_, data_stage_2__4555_, data_stage_2__4554_, data_stage_2__4553_, data_stage_2__4552_, data_stage_2__4551_, data_stage_2__4550_, data_stage_2__4549_, data_stage_2__4548_, data_stage_2__4547_, data_stage_2__4546_, data_stage_2__4545_, data_stage_2__4544_, data_stage_2__4543_, data_stage_2__4542_, data_stage_2__4541_, data_stage_2__4540_, data_stage_2__4539_, data_stage_2__4538_, data_stage_2__4537_, data_stage_2__4536_, data_stage_2__4535_, data_stage_2__4534_, data_stage_2__4533_, data_stage_2__4532_, data_stage_2__4531_, data_stage_2__4530_, data_stage_2__4529_, data_stage_2__4528_, data_stage_2__4527_, data_stage_2__4526_, data_stage_2__4525_, data_stage_2__4524_, data_stage_2__4523_, data_stage_2__4522_, data_stage_2__4521_, data_stage_2__4520_, data_stage_2__4519_, data_stage_2__4518_, data_stage_2__4517_, data_stage_2__4516_, data_stage_2__4515_, data_stage_2__4514_, data_stage_2__4513_, data_stage_2__4512_, data_stage_2__4511_, data_stage_2__4510_, data_stage_2__4509_, data_stage_2__4508_, data_stage_2__4507_, data_stage_2__4506_, data_stage_2__4505_, data_stage_2__4504_, data_stage_2__4503_, data_stage_2__4502_, data_stage_2__4501_, data_stage_2__4500_, data_stage_2__4499_, data_stage_2__4498_, data_stage_2__4497_, data_stage_2__4496_, data_stage_2__4495_, data_stage_2__4494_, data_stage_2__4493_, data_stage_2__4492_, data_stage_2__4491_, data_stage_2__4490_, data_stage_2__4489_, data_stage_2__4488_, data_stage_2__4487_, data_stage_2__4486_, data_stage_2__4485_, data_stage_2__4484_, data_stage_2__4483_, data_stage_2__4482_, data_stage_2__4481_, data_stage_2__4480_, data_stage_2__4479_, data_stage_2__4478_, data_stage_2__4477_, data_stage_2__4476_, data_stage_2__4475_, data_stage_2__4474_, data_stage_2__4473_, data_stage_2__4472_, data_stage_2__4471_, data_stage_2__4470_, data_stage_2__4469_, data_stage_2__4468_, data_stage_2__4467_, data_stage_2__4466_, data_stage_2__4465_, data_stage_2__4464_, data_stage_2__4463_, data_stage_2__4462_, data_stage_2__4461_, data_stage_2__4460_, data_stage_2__4459_, data_stage_2__4458_, data_stage_2__4457_, data_stage_2__4456_, data_stage_2__4455_, data_stage_2__4454_, data_stage_2__4453_, data_stage_2__4452_, data_stage_2__4451_, data_stage_2__4450_, data_stage_2__4449_, data_stage_2__4448_, data_stage_2__4447_, data_stage_2__4446_, data_stage_2__4445_, data_stage_2__4444_, data_stage_2__4443_, data_stage_2__4442_, data_stage_2__4441_, data_stage_2__4440_, data_stage_2__4439_, data_stage_2__4438_, data_stage_2__4437_, data_stage_2__4436_, data_stage_2__4435_, data_stage_2__4434_, data_stage_2__4433_, data_stage_2__4432_, data_stage_2__4431_, data_stage_2__4430_, data_stage_2__4429_, data_stage_2__4428_, data_stage_2__4427_, data_stage_2__4426_, data_stage_2__4425_, data_stage_2__4424_, data_stage_2__4423_, data_stage_2__4422_, data_stage_2__4421_, data_stage_2__4420_, data_stage_2__4419_, data_stage_2__4418_, data_stage_2__4417_, data_stage_2__4416_, data_stage_2__4415_, data_stage_2__4414_, data_stage_2__4413_, data_stage_2__4412_, data_stage_2__4411_, data_stage_2__4410_, data_stage_2__4409_, data_stage_2__4408_, data_stage_2__4407_, data_stage_2__4406_, data_stage_2__4405_, data_stage_2__4404_, data_stage_2__4403_, data_stage_2__4402_, data_stage_2__4401_, data_stage_2__4400_, data_stage_2__4399_, data_stage_2__4398_, data_stage_2__4397_, data_stage_2__4396_, data_stage_2__4395_, data_stage_2__4394_, data_stage_2__4393_, data_stage_2__4392_, data_stage_2__4391_, data_stage_2__4390_, data_stage_2__4389_, data_stage_2__4388_, data_stage_2__4387_, data_stage_2__4386_, data_stage_2__4385_, data_stage_2__4384_, data_stage_2__4383_, data_stage_2__4382_, data_stage_2__4381_, data_stage_2__4380_, data_stage_2__4379_, data_stage_2__4378_, data_stage_2__4377_, data_stage_2__4376_, data_stage_2__4375_, data_stage_2__4374_, data_stage_2__4373_, data_stage_2__4372_, data_stage_2__4371_, data_stage_2__4370_, data_stage_2__4369_, data_stage_2__4368_, data_stage_2__4367_, data_stage_2__4366_, data_stage_2__4365_, data_stage_2__4364_, data_stage_2__4363_, data_stage_2__4362_, data_stage_2__4361_, data_stage_2__4360_, data_stage_2__4359_, data_stage_2__4358_, data_stage_2__4357_, data_stage_2__4356_, data_stage_2__4355_, data_stage_2__4354_, data_stage_2__4353_, data_stage_2__4352_, data_stage_2__4351_, data_stage_2__4350_, data_stage_2__4349_, data_stage_2__4348_, data_stage_2__4347_, data_stage_2__4346_, data_stage_2__4345_, data_stage_2__4344_, data_stage_2__4343_, data_stage_2__4342_, data_stage_2__4341_, data_stage_2__4340_, data_stage_2__4339_, data_stage_2__4338_, data_stage_2__4337_, data_stage_2__4336_, data_stage_2__4335_, data_stage_2__4334_, data_stage_2__4333_, data_stage_2__4332_, data_stage_2__4331_, data_stage_2__4330_, data_stage_2__4329_, data_stage_2__4328_, data_stage_2__4327_, data_stage_2__4326_, data_stage_2__4325_, data_stage_2__4324_, data_stage_2__4323_, data_stage_2__4322_, data_stage_2__4321_, data_stage_2__4320_, data_stage_2__4319_, data_stage_2__4318_, data_stage_2__4317_, data_stage_2__4316_, data_stage_2__4315_, data_stage_2__4314_, data_stage_2__4313_, data_stage_2__4312_, data_stage_2__4311_, data_stage_2__4310_, data_stage_2__4309_, data_stage_2__4308_, data_stage_2__4307_, data_stage_2__4306_, data_stage_2__4305_, data_stage_2__4304_, data_stage_2__4303_, data_stage_2__4302_, data_stage_2__4301_, data_stage_2__4300_, data_stage_2__4299_, data_stage_2__4298_, data_stage_2__4297_, data_stage_2__4296_, data_stage_2__4295_, data_stage_2__4294_, data_stage_2__4293_, data_stage_2__4292_, data_stage_2__4291_, data_stage_2__4290_, data_stage_2__4289_, data_stage_2__4288_, data_stage_2__4287_, data_stage_2__4286_, data_stage_2__4285_, data_stage_2__4284_, data_stage_2__4283_, data_stage_2__4282_, data_stage_2__4281_, data_stage_2__4280_, data_stage_2__4279_, data_stage_2__4278_, data_stage_2__4277_, data_stage_2__4276_, data_stage_2__4275_, data_stage_2__4274_, data_stage_2__4273_, data_stage_2__4272_, data_stage_2__4271_, data_stage_2__4270_, data_stage_2__4269_, data_stage_2__4268_, data_stage_2__4267_, data_stage_2__4266_, data_stage_2__4265_, data_stage_2__4264_, data_stage_2__4263_, data_stage_2__4262_, data_stage_2__4261_, data_stage_2__4260_, data_stage_2__4259_, data_stage_2__4258_, data_stage_2__4257_, data_stage_2__4256_, data_stage_2__4255_, data_stage_2__4254_, data_stage_2__4253_, data_stage_2__4252_, data_stage_2__4251_, data_stage_2__4250_, data_stage_2__4249_, data_stage_2__4248_, data_stage_2__4247_, data_stage_2__4246_, data_stage_2__4245_, data_stage_2__4244_, data_stage_2__4243_, data_stage_2__4242_, data_stage_2__4241_, data_stage_2__4240_, data_stage_2__4239_, data_stage_2__4238_, data_stage_2__4237_, data_stage_2__4236_, data_stage_2__4235_, data_stage_2__4234_, data_stage_2__4233_, data_stage_2__4232_, data_stage_2__4231_, data_stage_2__4230_, data_stage_2__4229_, data_stage_2__4228_, data_stage_2__4227_, data_stage_2__4226_, data_stage_2__4225_, data_stage_2__4224_, data_stage_2__4223_, data_stage_2__4222_, data_stage_2__4221_, data_stage_2__4220_, data_stage_2__4219_, data_stage_2__4218_, data_stage_2__4217_, data_stage_2__4216_, data_stage_2__4215_, data_stage_2__4214_, data_stage_2__4213_, data_stage_2__4212_, data_stage_2__4211_, data_stage_2__4210_, data_stage_2__4209_, data_stage_2__4208_, data_stage_2__4207_, data_stage_2__4206_, data_stage_2__4205_, data_stage_2__4204_, data_stage_2__4203_, data_stage_2__4202_, data_stage_2__4201_, data_stage_2__4200_, data_stage_2__4199_, data_stage_2__4198_, data_stage_2__4197_, data_stage_2__4196_, data_stage_2__4195_, data_stage_2__4194_, data_stage_2__4193_, data_stage_2__4192_, data_stage_2__4191_, data_stage_2__4190_, data_stage_2__4189_, data_stage_2__4188_, data_stage_2__4187_, data_stage_2__4186_, data_stage_2__4185_, data_stage_2__4184_, data_stage_2__4183_, data_stage_2__4182_, data_stage_2__4181_, data_stage_2__4180_, data_stage_2__4179_, data_stage_2__4178_, data_stage_2__4177_, data_stage_2__4176_, data_stage_2__4175_, data_stage_2__4174_, data_stage_2__4173_, data_stage_2__4172_, data_stage_2__4171_, data_stage_2__4170_, data_stage_2__4169_, data_stage_2__4168_, data_stage_2__4167_, data_stage_2__4166_, data_stage_2__4165_, data_stage_2__4164_, data_stage_2__4163_, data_stage_2__4162_, data_stage_2__4161_, data_stage_2__4160_, data_stage_2__4159_, data_stage_2__4158_, data_stage_2__4157_, data_stage_2__4156_, data_stage_2__4155_, data_stage_2__4154_, data_stage_2__4153_, data_stage_2__4152_, data_stage_2__4151_, data_stage_2__4150_, data_stage_2__4149_, data_stage_2__4148_, data_stage_2__4147_, data_stage_2__4146_, data_stage_2__4145_, data_stage_2__4144_, data_stage_2__4143_, data_stage_2__4142_, data_stage_2__4141_, data_stage_2__4140_, data_stage_2__4139_, data_stage_2__4138_, data_stage_2__4137_, data_stage_2__4136_, data_stage_2__4135_, data_stage_2__4134_, data_stage_2__4133_, data_stage_2__4132_, data_stage_2__4131_, data_stage_2__4130_, data_stage_2__4129_, data_stage_2__4128_, data_stage_2__4127_, data_stage_2__4126_, data_stage_2__4125_, data_stage_2__4124_, data_stage_2__4123_, data_stage_2__4122_, data_stage_2__4121_, data_stage_2__4120_, data_stage_2__4119_, data_stage_2__4118_, data_stage_2__4117_, data_stage_2__4116_, data_stage_2__4115_, data_stage_2__4114_, data_stage_2__4113_, data_stage_2__4112_, data_stage_2__4111_, data_stage_2__4110_, data_stage_2__4109_, data_stage_2__4108_, data_stage_2__4107_, data_stage_2__4106_, data_stage_2__4105_, data_stage_2__4104_, data_stage_2__4103_, data_stage_2__4102_, data_stage_2__4101_, data_stage_2__4100_, data_stage_2__4099_, data_stage_2__4098_, data_stage_2__4097_, data_stage_2__4096_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_9__swap_inst
  (
    .data_i({ data_stage_1__5119_, data_stage_1__5118_, data_stage_1__5117_, data_stage_1__5116_, data_stage_1__5115_, data_stage_1__5114_, data_stage_1__5113_, data_stage_1__5112_, data_stage_1__5111_, data_stage_1__5110_, data_stage_1__5109_, data_stage_1__5108_, data_stage_1__5107_, data_stage_1__5106_, data_stage_1__5105_, data_stage_1__5104_, data_stage_1__5103_, data_stage_1__5102_, data_stage_1__5101_, data_stage_1__5100_, data_stage_1__5099_, data_stage_1__5098_, data_stage_1__5097_, data_stage_1__5096_, data_stage_1__5095_, data_stage_1__5094_, data_stage_1__5093_, data_stage_1__5092_, data_stage_1__5091_, data_stage_1__5090_, data_stage_1__5089_, data_stage_1__5088_, data_stage_1__5087_, data_stage_1__5086_, data_stage_1__5085_, data_stage_1__5084_, data_stage_1__5083_, data_stage_1__5082_, data_stage_1__5081_, data_stage_1__5080_, data_stage_1__5079_, data_stage_1__5078_, data_stage_1__5077_, data_stage_1__5076_, data_stage_1__5075_, data_stage_1__5074_, data_stage_1__5073_, data_stage_1__5072_, data_stage_1__5071_, data_stage_1__5070_, data_stage_1__5069_, data_stage_1__5068_, data_stage_1__5067_, data_stage_1__5066_, data_stage_1__5065_, data_stage_1__5064_, data_stage_1__5063_, data_stage_1__5062_, data_stage_1__5061_, data_stage_1__5060_, data_stage_1__5059_, data_stage_1__5058_, data_stage_1__5057_, data_stage_1__5056_, data_stage_1__5055_, data_stage_1__5054_, data_stage_1__5053_, data_stage_1__5052_, data_stage_1__5051_, data_stage_1__5050_, data_stage_1__5049_, data_stage_1__5048_, data_stage_1__5047_, data_stage_1__5046_, data_stage_1__5045_, data_stage_1__5044_, data_stage_1__5043_, data_stage_1__5042_, data_stage_1__5041_, data_stage_1__5040_, data_stage_1__5039_, data_stage_1__5038_, data_stage_1__5037_, data_stage_1__5036_, data_stage_1__5035_, data_stage_1__5034_, data_stage_1__5033_, data_stage_1__5032_, data_stage_1__5031_, data_stage_1__5030_, data_stage_1__5029_, data_stage_1__5028_, data_stage_1__5027_, data_stage_1__5026_, data_stage_1__5025_, data_stage_1__5024_, data_stage_1__5023_, data_stage_1__5022_, data_stage_1__5021_, data_stage_1__5020_, data_stage_1__5019_, data_stage_1__5018_, data_stage_1__5017_, data_stage_1__5016_, data_stage_1__5015_, data_stage_1__5014_, data_stage_1__5013_, data_stage_1__5012_, data_stage_1__5011_, data_stage_1__5010_, data_stage_1__5009_, data_stage_1__5008_, data_stage_1__5007_, data_stage_1__5006_, data_stage_1__5005_, data_stage_1__5004_, data_stage_1__5003_, data_stage_1__5002_, data_stage_1__5001_, data_stage_1__5000_, data_stage_1__4999_, data_stage_1__4998_, data_stage_1__4997_, data_stage_1__4996_, data_stage_1__4995_, data_stage_1__4994_, data_stage_1__4993_, data_stage_1__4992_, data_stage_1__4991_, data_stage_1__4990_, data_stage_1__4989_, data_stage_1__4988_, data_stage_1__4987_, data_stage_1__4986_, data_stage_1__4985_, data_stage_1__4984_, data_stage_1__4983_, data_stage_1__4982_, data_stage_1__4981_, data_stage_1__4980_, data_stage_1__4979_, data_stage_1__4978_, data_stage_1__4977_, data_stage_1__4976_, data_stage_1__4975_, data_stage_1__4974_, data_stage_1__4973_, data_stage_1__4972_, data_stage_1__4971_, data_stage_1__4970_, data_stage_1__4969_, data_stage_1__4968_, data_stage_1__4967_, data_stage_1__4966_, data_stage_1__4965_, data_stage_1__4964_, data_stage_1__4963_, data_stage_1__4962_, data_stage_1__4961_, data_stage_1__4960_, data_stage_1__4959_, data_stage_1__4958_, data_stage_1__4957_, data_stage_1__4956_, data_stage_1__4955_, data_stage_1__4954_, data_stage_1__4953_, data_stage_1__4952_, data_stage_1__4951_, data_stage_1__4950_, data_stage_1__4949_, data_stage_1__4948_, data_stage_1__4947_, data_stage_1__4946_, data_stage_1__4945_, data_stage_1__4944_, data_stage_1__4943_, data_stage_1__4942_, data_stage_1__4941_, data_stage_1__4940_, data_stage_1__4939_, data_stage_1__4938_, data_stage_1__4937_, data_stage_1__4936_, data_stage_1__4935_, data_stage_1__4934_, data_stage_1__4933_, data_stage_1__4932_, data_stage_1__4931_, data_stage_1__4930_, data_stage_1__4929_, data_stage_1__4928_, data_stage_1__4927_, data_stage_1__4926_, data_stage_1__4925_, data_stage_1__4924_, data_stage_1__4923_, data_stage_1__4922_, data_stage_1__4921_, data_stage_1__4920_, data_stage_1__4919_, data_stage_1__4918_, data_stage_1__4917_, data_stage_1__4916_, data_stage_1__4915_, data_stage_1__4914_, data_stage_1__4913_, data_stage_1__4912_, data_stage_1__4911_, data_stage_1__4910_, data_stage_1__4909_, data_stage_1__4908_, data_stage_1__4907_, data_stage_1__4906_, data_stage_1__4905_, data_stage_1__4904_, data_stage_1__4903_, data_stage_1__4902_, data_stage_1__4901_, data_stage_1__4900_, data_stage_1__4899_, data_stage_1__4898_, data_stage_1__4897_, data_stage_1__4896_, data_stage_1__4895_, data_stage_1__4894_, data_stage_1__4893_, data_stage_1__4892_, data_stage_1__4891_, data_stage_1__4890_, data_stage_1__4889_, data_stage_1__4888_, data_stage_1__4887_, data_stage_1__4886_, data_stage_1__4885_, data_stage_1__4884_, data_stage_1__4883_, data_stage_1__4882_, data_stage_1__4881_, data_stage_1__4880_, data_stage_1__4879_, data_stage_1__4878_, data_stage_1__4877_, data_stage_1__4876_, data_stage_1__4875_, data_stage_1__4874_, data_stage_1__4873_, data_stage_1__4872_, data_stage_1__4871_, data_stage_1__4870_, data_stage_1__4869_, data_stage_1__4868_, data_stage_1__4867_, data_stage_1__4866_, data_stage_1__4865_, data_stage_1__4864_, data_stage_1__4863_, data_stage_1__4862_, data_stage_1__4861_, data_stage_1__4860_, data_stage_1__4859_, data_stage_1__4858_, data_stage_1__4857_, data_stage_1__4856_, data_stage_1__4855_, data_stage_1__4854_, data_stage_1__4853_, data_stage_1__4852_, data_stage_1__4851_, data_stage_1__4850_, data_stage_1__4849_, data_stage_1__4848_, data_stage_1__4847_, data_stage_1__4846_, data_stage_1__4845_, data_stage_1__4844_, data_stage_1__4843_, data_stage_1__4842_, data_stage_1__4841_, data_stage_1__4840_, data_stage_1__4839_, data_stage_1__4838_, data_stage_1__4837_, data_stage_1__4836_, data_stage_1__4835_, data_stage_1__4834_, data_stage_1__4833_, data_stage_1__4832_, data_stage_1__4831_, data_stage_1__4830_, data_stage_1__4829_, data_stage_1__4828_, data_stage_1__4827_, data_stage_1__4826_, data_stage_1__4825_, data_stage_1__4824_, data_stage_1__4823_, data_stage_1__4822_, data_stage_1__4821_, data_stage_1__4820_, data_stage_1__4819_, data_stage_1__4818_, data_stage_1__4817_, data_stage_1__4816_, data_stage_1__4815_, data_stage_1__4814_, data_stage_1__4813_, data_stage_1__4812_, data_stage_1__4811_, data_stage_1__4810_, data_stage_1__4809_, data_stage_1__4808_, data_stage_1__4807_, data_stage_1__4806_, data_stage_1__4805_, data_stage_1__4804_, data_stage_1__4803_, data_stage_1__4802_, data_stage_1__4801_, data_stage_1__4800_, data_stage_1__4799_, data_stage_1__4798_, data_stage_1__4797_, data_stage_1__4796_, data_stage_1__4795_, data_stage_1__4794_, data_stage_1__4793_, data_stage_1__4792_, data_stage_1__4791_, data_stage_1__4790_, data_stage_1__4789_, data_stage_1__4788_, data_stage_1__4787_, data_stage_1__4786_, data_stage_1__4785_, data_stage_1__4784_, data_stage_1__4783_, data_stage_1__4782_, data_stage_1__4781_, data_stage_1__4780_, data_stage_1__4779_, data_stage_1__4778_, data_stage_1__4777_, data_stage_1__4776_, data_stage_1__4775_, data_stage_1__4774_, data_stage_1__4773_, data_stage_1__4772_, data_stage_1__4771_, data_stage_1__4770_, data_stage_1__4769_, data_stage_1__4768_, data_stage_1__4767_, data_stage_1__4766_, data_stage_1__4765_, data_stage_1__4764_, data_stage_1__4763_, data_stage_1__4762_, data_stage_1__4761_, data_stage_1__4760_, data_stage_1__4759_, data_stage_1__4758_, data_stage_1__4757_, data_stage_1__4756_, data_stage_1__4755_, data_stage_1__4754_, data_stage_1__4753_, data_stage_1__4752_, data_stage_1__4751_, data_stage_1__4750_, data_stage_1__4749_, data_stage_1__4748_, data_stage_1__4747_, data_stage_1__4746_, data_stage_1__4745_, data_stage_1__4744_, data_stage_1__4743_, data_stage_1__4742_, data_stage_1__4741_, data_stage_1__4740_, data_stage_1__4739_, data_stage_1__4738_, data_stage_1__4737_, data_stage_1__4736_, data_stage_1__4735_, data_stage_1__4734_, data_stage_1__4733_, data_stage_1__4732_, data_stage_1__4731_, data_stage_1__4730_, data_stage_1__4729_, data_stage_1__4728_, data_stage_1__4727_, data_stage_1__4726_, data_stage_1__4725_, data_stage_1__4724_, data_stage_1__4723_, data_stage_1__4722_, data_stage_1__4721_, data_stage_1__4720_, data_stage_1__4719_, data_stage_1__4718_, data_stage_1__4717_, data_stage_1__4716_, data_stage_1__4715_, data_stage_1__4714_, data_stage_1__4713_, data_stage_1__4712_, data_stage_1__4711_, data_stage_1__4710_, data_stage_1__4709_, data_stage_1__4708_, data_stage_1__4707_, data_stage_1__4706_, data_stage_1__4705_, data_stage_1__4704_, data_stage_1__4703_, data_stage_1__4702_, data_stage_1__4701_, data_stage_1__4700_, data_stage_1__4699_, data_stage_1__4698_, data_stage_1__4697_, data_stage_1__4696_, data_stage_1__4695_, data_stage_1__4694_, data_stage_1__4693_, data_stage_1__4692_, data_stage_1__4691_, data_stage_1__4690_, data_stage_1__4689_, data_stage_1__4688_, data_stage_1__4687_, data_stage_1__4686_, data_stage_1__4685_, data_stage_1__4684_, data_stage_1__4683_, data_stage_1__4682_, data_stage_1__4681_, data_stage_1__4680_, data_stage_1__4679_, data_stage_1__4678_, data_stage_1__4677_, data_stage_1__4676_, data_stage_1__4675_, data_stage_1__4674_, data_stage_1__4673_, data_stage_1__4672_, data_stage_1__4671_, data_stage_1__4670_, data_stage_1__4669_, data_stage_1__4668_, data_stage_1__4667_, data_stage_1__4666_, data_stage_1__4665_, data_stage_1__4664_, data_stage_1__4663_, data_stage_1__4662_, data_stage_1__4661_, data_stage_1__4660_, data_stage_1__4659_, data_stage_1__4658_, data_stage_1__4657_, data_stage_1__4656_, data_stage_1__4655_, data_stage_1__4654_, data_stage_1__4653_, data_stage_1__4652_, data_stage_1__4651_, data_stage_1__4650_, data_stage_1__4649_, data_stage_1__4648_, data_stage_1__4647_, data_stage_1__4646_, data_stage_1__4645_, data_stage_1__4644_, data_stage_1__4643_, data_stage_1__4642_, data_stage_1__4641_, data_stage_1__4640_, data_stage_1__4639_, data_stage_1__4638_, data_stage_1__4637_, data_stage_1__4636_, data_stage_1__4635_, data_stage_1__4634_, data_stage_1__4633_, data_stage_1__4632_, data_stage_1__4631_, data_stage_1__4630_, data_stage_1__4629_, data_stage_1__4628_, data_stage_1__4627_, data_stage_1__4626_, data_stage_1__4625_, data_stage_1__4624_, data_stage_1__4623_, data_stage_1__4622_, data_stage_1__4621_, data_stage_1__4620_, data_stage_1__4619_, data_stage_1__4618_, data_stage_1__4617_, data_stage_1__4616_, data_stage_1__4615_, data_stage_1__4614_, data_stage_1__4613_, data_stage_1__4612_, data_stage_1__4611_, data_stage_1__4610_, data_stage_1__4609_, data_stage_1__4608_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__5119_, data_stage_2__5118_, data_stage_2__5117_, data_stage_2__5116_, data_stage_2__5115_, data_stage_2__5114_, data_stage_2__5113_, data_stage_2__5112_, data_stage_2__5111_, data_stage_2__5110_, data_stage_2__5109_, data_stage_2__5108_, data_stage_2__5107_, data_stage_2__5106_, data_stage_2__5105_, data_stage_2__5104_, data_stage_2__5103_, data_stage_2__5102_, data_stage_2__5101_, data_stage_2__5100_, data_stage_2__5099_, data_stage_2__5098_, data_stage_2__5097_, data_stage_2__5096_, data_stage_2__5095_, data_stage_2__5094_, data_stage_2__5093_, data_stage_2__5092_, data_stage_2__5091_, data_stage_2__5090_, data_stage_2__5089_, data_stage_2__5088_, data_stage_2__5087_, data_stage_2__5086_, data_stage_2__5085_, data_stage_2__5084_, data_stage_2__5083_, data_stage_2__5082_, data_stage_2__5081_, data_stage_2__5080_, data_stage_2__5079_, data_stage_2__5078_, data_stage_2__5077_, data_stage_2__5076_, data_stage_2__5075_, data_stage_2__5074_, data_stage_2__5073_, data_stage_2__5072_, data_stage_2__5071_, data_stage_2__5070_, data_stage_2__5069_, data_stage_2__5068_, data_stage_2__5067_, data_stage_2__5066_, data_stage_2__5065_, data_stage_2__5064_, data_stage_2__5063_, data_stage_2__5062_, data_stage_2__5061_, data_stage_2__5060_, data_stage_2__5059_, data_stage_2__5058_, data_stage_2__5057_, data_stage_2__5056_, data_stage_2__5055_, data_stage_2__5054_, data_stage_2__5053_, data_stage_2__5052_, data_stage_2__5051_, data_stage_2__5050_, data_stage_2__5049_, data_stage_2__5048_, data_stage_2__5047_, data_stage_2__5046_, data_stage_2__5045_, data_stage_2__5044_, data_stage_2__5043_, data_stage_2__5042_, data_stage_2__5041_, data_stage_2__5040_, data_stage_2__5039_, data_stage_2__5038_, data_stage_2__5037_, data_stage_2__5036_, data_stage_2__5035_, data_stage_2__5034_, data_stage_2__5033_, data_stage_2__5032_, data_stage_2__5031_, data_stage_2__5030_, data_stage_2__5029_, data_stage_2__5028_, data_stage_2__5027_, data_stage_2__5026_, data_stage_2__5025_, data_stage_2__5024_, data_stage_2__5023_, data_stage_2__5022_, data_stage_2__5021_, data_stage_2__5020_, data_stage_2__5019_, data_stage_2__5018_, data_stage_2__5017_, data_stage_2__5016_, data_stage_2__5015_, data_stage_2__5014_, data_stage_2__5013_, data_stage_2__5012_, data_stage_2__5011_, data_stage_2__5010_, data_stage_2__5009_, data_stage_2__5008_, data_stage_2__5007_, data_stage_2__5006_, data_stage_2__5005_, data_stage_2__5004_, data_stage_2__5003_, data_stage_2__5002_, data_stage_2__5001_, data_stage_2__5000_, data_stage_2__4999_, data_stage_2__4998_, data_stage_2__4997_, data_stage_2__4996_, data_stage_2__4995_, data_stage_2__4994_, data_stage_2__4993_, data_stage_2__4992_, data_stage_2__4991_, data_stage_2__4990_, data_stage_2__4989_, data_stage_2__4988_, data_stage_2__4987_, data_stage_2__4986_, data_stage_2__4985_, data_stage_2__4984_, data_stage_2__4983_, data_stage_2__4982_, data_stage_2__4981_, data_stage_2__4980_, data_stage_2__4979_, data_stage_2__4978_, data_stage_2__4977_, data_stage_2__4976_, data_stage_2__4975_, data_stage_2__4974_, data_stage_2__4973_, data_stage_2__4972_, data_stage_2__4971_, data_stage_2__4970_, data_stage_2__4969_, data_stage_2__4968_, data_stage_2__4967_, data_stage_2__4966_, data_stage_2__4965_, data_stage_2__4964_, data_stage_2__4963_, data_stage_2__4962_, data_stage_2__4961_, data_stage_2__4960_, data_stage_2__4959_, data_stage_2__4958_, data_stage_2__4957_, data_stage_2__4956_, data_stage_2__4955_, data_stage_2__4954_, data_stage_2__4953_, data_stage_2__4952_, data_stage_2__4951_, data_stage_2__4950_, data_stage_2__4949_, data_stage_2__4948_, data_stage_2__4947_, data_stage_2__4946_, data_stage_2__4945_, data_stage_2__4944_, data_stage_2__4943_, data_stage_2__4942_, data_stage_2__4941_, data_stage_2__4940_, data_stage_2__4939_, data_stage_2__4938_, data_stage_2__4937_, data_stage_2__4936_, data_stage_2__4935_, data_stage_2__4934_, data_stage_2__4933_, data_stage_2__4932_, data_stage_2__4931_, data_stage_2__4930_, data_stage_2__4929_, data_stage_2__4928_, data_stage_2__4927_, data_stage_2__4926_, data_stage_2__4925_, data_stage_2__4924_, data_stage_2__4923_, data_stage_2__4922_, data_stage_2__4921_, data_stage_2__4920_, data_stage_2__4919_, data_stage_2__4918_, data_stage_2__4917_, data_stage_2__4916_, data_stage_2__4915_, data_stage_2__4914_, data_stage_2__4913_, data_stage_2__4912_, data_stage_2__4911_, data_stage_2__4910_, data_stage_2__4909_, data_stage_2__4908_, data_stage_2__4907_, data_stage_2__4906_, data_stage_2__4905_, data_stage_2__4904_, data_stage_2__4903_, data_stage_2__4902_, data_stage_2__4901_, data_stage_2__4900_, data_stage_2__4899_, data_stage_2__4898_, data_stage_2__4897_, data_stage_2__4896_, data_stage_2__4895_, data_stage_2__4894_, data_stage_2__4893_, data_stage_2__4892_, data_stage_2__4891_, data_stage_2__4890_, data_stage_2__4889_, data_stage_2__4888_, data_stage_2__4887_, data_stage_2__4886_, data_stage_2__4885_, data_stage_2__4884_, data_stage_2__4883_, data_stage_2__4882_, data_stage_2__4881_, data_stage_2__4880_, data_stage_2__4879_, data_stage_2__4878_, data_stage_2__4877_, data_stage_2__4876_, data_stage_2__4875_, data_stage_2__4874_, data_stage_2__4873_, data_stage_2__4872_, data_stage_2__4871_, data_stage_2__4870_, data_stage_2__4869_, data_stage_2__4868_, data_stage_2__4867_, data_stage_2__4866_, data_stage_2__4865_, data_stage_2__4864_, data_stage_2__4863_, data_stage_2__4862_, data_stage_2__4861_, data_stage_2__4860_, data_stage_2__4859_, data_stage_2__4858_, data_stage_2__4857_, data_stage_2__4856_, data_stage_2__4855_, data_stage_2__4854_, data_stage_2__4853_, data_stage_2__4852_, data_stage_2__4851_, data_stage_2__4850_, data_stage_2__4849_, data_stage_2__4848_, data_stage_2__4847_, data_stage_2__4846_, data_stage_2__4845_, data_stage_2__4844_, data_stage_2__4843_, data_stage_2__4842_, data_stage_2__4841_, data_stage_2__4840_, data_stage_2__4839_, data_stage_2__4838_, data_stage_2__4837_, data_stage_2__4836_, data_stage_2__4835_, data_stage_2__4834_, data_stage_2__4833_, data_stage_2__4832_, data_stage_2__4831_, data_stage_2__4830_, data_stage_2__4829_, data_stage_2__4828_, data_stage_2__4827_, data_stage_2__4826_, data_stage_2__4825_, data_stage_2__4824_, data_stage_2__4823_, data_stage_2__4822_, data_stage_2__4821_, data_stage_2__4820_, data_stage_2__4819_, data_stage_2__4818_, data_stage_2__4817_, data_stage_2__4816_, data_stage_2__4815_, data_stage_2__4814_, data_stage_2__4813_, data_stage_2__4812_, data_stage_2__4811_, data_stage_2__4810_, data_stage_2__4809_, data_stage_2__4808_, data_stage_2__4807_, data_stage_2__4806_, data_stage_2__4805_, data_stage_2__4804_, data_stage_2__4803_, data_stage_2__4802_, data_stage_2__4801_, data_stage_2__4800_, data_stage_2__4799_, data_stage_2__4798_, data_stage_2__4797_, data_stage_2__4796_, data_stage_2__4795_, data_stage_2__4794_, data_stage_2__4793_, data_stage_2__4792_, data_stage_2__4791_, data_stage_2__4790_, data_stage_2__4789_, data_stage_2__4788_, data_stage_2__4787_, data_stage_2__4786_, data_stage_2__4785_, data_stage_2__4784_, data_stage_2__4783_, data_stage_2__4782_, data_stage_2__4781_, data_stage_2__4780_, data_stage_2__4779_, data_stage_2__4778_, data_stage_2__4777_, data_stage_2__4776_, data_stage_2__4775_, data_stage_2__4774_, data_stage_2__4773_, data_stage_2__4772_, data_stage_2__4771_, data_stage_2__4770_, data_stage_2__4769_, data_stage_2__4768_, data_stage_2__4767_, data_stage_2__4766_, data_stage_2__4765_, data_stage_2__4764_, data_stage_2__4763_, data_stage_2__4762_, data_stage_2__4761_, data_stage_2__4760_, data_stage_2__4759_, data_stage_2__4758_, data_stage_2__4757_, data_stage_2__4756_, data_stage_2__4755_, data_stage_2__4754_, data_stage_2__4753_, data_stage_2__4752_, data_stage_2__4751_, data_stage_2__4750_, data_stage_2__4749_, data_stage_2__4748_, data_stage_2__4747_, data_stage_2__4746_, data_stage_2__4745_, data_stage_2__4744_, data_stage_2__4743_, data_stage_2__4742_, data_stage_2__4741_, data_stage_2__4740_, data_stage_2__4739_, data_stage_2__4738_, data_stage_2__4737_, data_stage_2__4736_, data_stage_2__4735_, data_stage_2__4734_, data_stage_2__4733_, data_stage_2__4732_, data_stage_2__4731_, data_stage_2__4730_, data_stage_2__4729_, data_stage_2__4728_, data_stage_2__4727_, data_stage_2__4726_, data_stage_2__4725_, data_stage_2__4724_, data_stage_2__4723_, data_stage_2__4722_, data_stage_2__4721_, data_stage_2__4720_, data_stage_2__4719_, data_stage_2__4718_, data_stage_2__4717_, data_stage_2__4716_, data_stage_2__4715_, data_stage_2__4714_, data_stage_2__4713_, data_stage_2__4712_, data_stage_2__4711_, data_stage_2__4710_, data_stage_2__4709_, data_stage_2__4708_, data_stage_2__4707_, data_stage_2__4706_, data_stage_2__4705_, data_stage_2__4704_, data_stage_2__4703_, data_stage_2__4702_, data_stage_2__4701_, data_stage_2__4700_, data_stage_2__4699_, data_stage_2__4698_, data_stage_2__4697_, data_stage_2__4696_, data_stage_2__4695_, data_stage_2__4694_, data_stage_2__4693_, data_stage_2__4692_, data_stage_2__4691_, data_stage_2__4690_, data_stage_2__4689_, data_stage_2__4688_, data_stage_2__4687_, data_stage_2__4686_, data_stage_2__4685_, data_stage_2__4684_, data_stage_2__4683_, data_stage_2__4682_, data_stage_2__4681_, data_stage_2__4680_, data_stage_2__4679_, data_stage_2__4678_, data_stage_2__4677_, data_stage_2__4676_, data_stage_2__4675_, data_stage_2__4674_, data_stage_2__4673_, data_stage_2__4672_, data_stage_2__4671_, data_stage_2__4670_, data_stage_2__4669_, data_stage_2__4668_, data_stage_2__4667_, data_stage_2__4666_, data_stage_2__4665_, data_stage_2__4664_, data_stage_2__4663_, data_stage_2__4662_, data_stage_2__4661_, data_stage_2__4660_, data_stage_2__4659_, data_stage_2__4658_, data_stage_2__4657_, data_stage_2__4656_, data_stage_2__4655_, data_stage_2__4654_, data_stage_2__4653_, data_stage_2__4652_, data_stage_2__4651_, data_stage_2__4650_, data_stage_2__4649_, data_stage_2__4648_, data_stage_2__4647_, data_stage_2__4646_, data_stage_2__4645_, data_stage_2__4644_, data_stage_2__4643_, data_stage_2__4642_, data_stage_2__4641_, data_stage_2__4640_, data_stage_2__4639_, data_stage_2__4638_, data_stage_2__4637_, data_stage_2__4636_, data_stage_2__4635_, data_stage_2__4634_, data_stage_2__4633_, data_stage_2__4632_, data_stage_2__4631_, data_stage_2__4630_, data_stage_2__4629_, data_stage_2__4628_, data_stage_2__4627_, data_stage_2__4626_, data_stage_2__4625_, data_stage_2__4624_, data_stage_2__4623_, data_stage_2__4622_, data_stage_2__4621_, data_stage_2__4620_, data_stage_2__4619_, data_stage_2__4618_, data_stage_2__4617_, data_stage_2__4616_, data_stage_2__4615_, data_stage_2__4614_, data_stage_2__4613_, data_stage_2__4612_, data_stage_2__4611_, data_stage_2__4610_, data_stage_2__4609_, data_stage_2__4608_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_10__swap_inst
  (
    .data_i({ data_stage_1__5631_, data_stage_1__5630_, data_stage_1__5629_, data_stage_1__5628_, data_stage_1__5627_, data_stage_1__5626_, data_stage_1__5625_, data_stage_1__5624_, data_stage_1__5623_, data_stage_1__5622_, data_stage_1__5621_, data_stage_1__5620_, data_stage_1__5619_, data_stage_1__5618_, data_stage_1__5617_, data_stage_1__5616_, data_stage_1__5615_, data_stage_1__5614_, data_stage_1__5613_, data_stage_1__5612_, data_stage_1__5611_, data_stage_1__5610_, data_stage_1__5609_, data_stage_1__5608_, data_stage_1__5607_, data_stage_1__5606_, data_stage_1__5605_, data_stage_1__5604_, data_stage_1__5603_, data_stage_1__5602_, data_stage_1__5601_, data_stage_1__5600_, data_stage_1__5599_, data_stage_1__5598_, data_stage_1__5597_, data_stage_1__5596_, data_stage_1__5595_, data_stage_1__5594_, data_stage_1__5593_, data_stage_1__5592_, data_stage_1__5591_, data_stage_1__5590_, data_stage_1__5589_, data_stage_1__5588_, data_stage_1__5587_, data_stage_1__5586_, data_stage_1__5585_, data_stage_1__5584_, data_stage_1__5583_, data_stage_1__5582_, data_stage_1__5581_, data_stage_1__5580_, data_stage_1__5579_, data_stage_1__5578_, data_stage_1__5577_, data_stage_1__5576_, data_stage_1__5575_, data_stage_1__5574_, data_stage_1__5573_, data_stage_1__5572_, data_stage_1__5571_, data_stage_1__5570_, data_stage_1__5569_, data_stage_1__5568_, data_stage_1__5567_, data_stage_1__5566_, data_stage_1__5565_, data_stage_1__5564_, data_stage_1__5563_, data_stage_1__5562_, data_stage_1__5561_, data_stage_1__5560_, data_stage_1__5559_, data_stage_1__5558_, data_stage_1__5557_, data_stage_1__5556_, data_stage_1__5555_, data_stage_1__5554_, data_stage_1__5553_, data_stage_1__5552_, data_stage_1__5551_, data_stage_1__5550_, data_stage_1__5549_, data_stage_1__5548_, data_stage_1__5547_, data_stage_1__5546_, data_stage_1__5545_, data_stage_1__5544_, data_stage_1__5543_, data_stage_1__5542_, data_stage_1__5541_, data_stage_1__5540_, data_stage_1__5539_, data_stage_1__5538_, data_stage_1__5537_, data_stage_1__5536_, data_stage_1__5535_, data_stage_1__5534_, data_stage_1__5533_, data_stage_1__5532_, data_stage_1__5531_, data_stage_1__5530_, data_stage_1__5529_, data_stage_1__5528_, data_stage_1__5527_, data_stage_1__5526_, data_stage_1__5525_, data_stage_1__5524_, data_stage_1__5523_, data_stage_1__5522_, data_stage_1__5521_, data_stage_1__5520_, data_stage_1__5519_, data_stage_1__5518_, data_stage_1__5517_, data_stage_1__5516_, data_stage_1__5515_, data_stage_1__5514_, data_stage_1__5513_, data_stage_1__5512_, data_stage_1__5511_, data_stage_1__5510_, data_stage_1__5509_, data_stage_1__5508_, data_stage_1__5507_, data_stage_1__5506_, data_stage_1__5505_, data_stage_1__5504_, data_stage_1__5503_, data_stage_1__5502_, data_stage_1__5501_, data_stage_1__5500_, data_stage_1__5499_, data_stage_1__5498_, data_stage_1__5497_, data_stage_1__5496_, data_stage_1__5495_, data_stage_1__5494_, data_stage_1__5493_, data_stage_1__5492_, data_stage_1__5491_, data_stage_1__5490_, data_stage_1__5489_, data_stage_1__5488_, data_stage_1__5487_, data_stage_1__5486_, data_stage_1__5485_, data_stage_1__5484_, data_stage_1__5483_, data_stage_1__5482_, data_stage_1__5481_, data_stage_1__5480_, data_stage_1__5479_, data_stage_1__5478_, data_stage_1__5477_, data_stage_1__5476_, data_stage_1__5475_, data_stage_1__5474_, data_stage_1__5473_, data_stage_1__5472_, data_stage_1__5471_, data_stage_1__5470_, data_stage_1__5469_, data_stage_1__5468_, data_stage_1__5467_, data_stage_1__5466_, data_stage_1__5465_, data_stage_1__5464_, data_stage_1__5463_, data_stage_1__5462_, data_stage_1__5461_, data_stage_1__5460_, data_stage_1__5459_, data_stage_1__5458_, data_stage_1__5457_, data_stage_1__5456_, data_stage_1__5455_, data_stage_1__5454_, data_stage_1__5453_, data_stage_1__5452_, data_stage_1__5451_, data_stage_1__5450_, data_stage_1__5449_, data_stage_1__5448_, data_stage_1__5447_, data_stage_1__5446_, data_stage_1__5445_, data_stage_1__5444_, data_stage_1__5443_, data_stage_1__5442_, data_stage_1__5441_, data_stage_1__5440_, data_stage_1__5439_, data_stage_1__5438_, data_stage_1__5437_, data_stage_1__5436_, data_stage_1__5435_, data_stage_1__5434_, data_stage_1__5433_, data_stage_1__5432_, data_stage_1__5431_, data_stage_1__5430_, data_stage_1__5429_, data_stage_1__5428_, data_stage_1__5427_, data_stage_1__5426_, data_stage_1__5425_, data_stage_1__5424_, data_stage_1__5423_, data_stage_1__5422_, data_stage_1__5421_, data_stage_1__5420_, data_stage_1__5419_, data_stage_1__5418_, data_stage_1__5417_, data_stage_1__5416_, data_stage_1__5415_, data_stage_1__5414_, data_stage_1__5413_, data_stage_1__5412_, data_stage_1__5411_, data_stage_1__5410_, data_stage_1__5409_, data_stage_1__5408_, data_stage_1__5407_, data_stage_1__5406_, data_stage_1__5405_, data_stage_1__5404_, data_stage_1__5403_, data_stage_1__5402_, data_stage_1__5401_, data_stage_1__5400_, data_stage_1__5399_, data_stage_1__5398_, data_stage_1__5397_, data_stage_1__5396_, data_stage_1__5395_, data_stage_1__5394_, data_stage_1__5393_, data_stage_1__5392_, data_stage_1__5391_, data_stage_1__5390_, data_stage_1__5389_, data_stage_1__5388_, data_stage_1__5387_, data_stage_1__5386_, data_stage_1__5385_, data_stage_1__5384_, data_stage_1__5383_, data_stage_1__5382_, data_stage_1__5381_, data_stage_1__5380_, data_stage_1__5379_, data_stage_1__5378_, data_stage_1__5377_, data_stage_1__5376_, data_stage_1__5375_, data_stage_1__5374_, data_stage_1__5373_, data_stage_1__5372_, data_stage_1__5371_, data_stage_1__5370_, data_stage_1__5369_, data_stage_1__5368_, data_stage_1__5367_, data_stage_1__5366_, data_stage_1__5365_, data_stage_1__5364_, data_stage_1__5363_, data_stage_1__5362_, data_stage_1__5361_, data_stage_1__5360_, data_stage_1__5359_, data_stage_1__5358_, data_stage_1__5357_, data_stage_1__5356_, data_stage_1__5355_, data_stage_1__5354_, data_stage_1__5353_, data_stage_1__5352_, data_stage_1__5351_, data_stage_1__5350_, data_stage_1__5349_, data_stage_1__5348_, data_stage_1__5347_, data_stage_1__5346_, data_stage_1__5345_, data_stage_1__5344_, data_stage_1__5343_, data_stage_1__5342_, data_stage_1__5341_, data_stage_1__5340_, data_stage_1__5339_, data_stage_1__5338_, data_stage_1__5337_, data_stage_1__5336_, data_stage_1__5335_, data_stage_1__5334_, data_stage_1__5333_, data_stage_1__5332_, data_stage_1__5331_, data_stage_1__5330_, data_stage_1__5329_, data_stage_1__5328_, data_stage_1__5327_, data_stage_1__5326_, data_stage_1__5325_, data_stage_1__5324_, data_stage_1__5323_, data_stage_1__5322_, data_stage_1__5321_, data_stage_1__5320_, data_stage_1__5319_, data_stage_1__5318_, data_stage_1__5317_, data_stage_1__5316_, data_stage_1__5315_, data_stage_1__5314_, data_stage_1__5313_, data_stage_1__5312_, data_stage_1__5311_, data_stage_1__5310_, data_stage_1__5309_, data_stage_1__5308_, data_stage_1__5307_, data_stage_1__5306_, data_stage_1__5305_, data_stage_1__5304_, data_stage_1__5303_, data_stage_1__5302_, data_stage_1__5301_, data_stage_1__5300_, data_stage_1__5299_, data_stage_1__5298_, data_stage_1__5297_, data_stage_1__5296_, data_stage_1__5295_, data_stage_1__5294_, data_stage_1__5293_, data_stage_1__5292_, data_stage_1__5291_, data_stage_1__5290_, data_stage_1__5289_, data_stage_1__5288_, data_stage_1__5287_, data_stage_1__5286_, data_stage_1__5285_, data_stage_1__5284_, data_stage_1__5283_, data_stage_1__5282_, data_stage_1__5281_, data_stage_1__5280_, data_stage_1__5279_, data_stage_1__5278_, data_stage_1__5277_, data_stage_1__5276_, data_stage_1__5275_, data_stage_1__5274_, data_stage_1__5273_, data_stage_1__5272_, data_stage_1__5271_, data_stage_1__5270_, data_stage_1__5269_, data_stage_1__5268_, data_stage_1__5267_, data_stage_1__5266_, data_stage_1__5265_, data_stage_1__5264_, data_stage_1__5263_, data_stage_1__5262_, data_stage_1__5261_, data_stage_1__5260_, data_stage_1__5259_, data_stage_1__5258_, data_stage_1__5257_, data_stage_1__5256_, data_stage_1__5255_, data_stage_1__5254_, data_stage_1__5253_, data_stage_1__5252_, data_stage_1__5251_, data_stage_1__5250_, data_stage_1__5249_, data_stage_1__5248_, data_stage_1__5247_, data_stage_1__5246_, data_stage_1__5245_, data_stage_1__5244_, data_stage_1__5243_, data_stage_1__5242_, data_stage_1__5241_, data_stage_1__5240_, data_stage_1__5239_, data_stage_1__5238_, data_stage_1__5237_, data_stage_1__5236_, data_stage_1__5235_, data_stage_1__5234_, data_stage_1__5233_, data_stage_1__5232_, data_stage_1__5231_, data_stage_1__5230_, data_stage_1__5229_, data_stage_1__5228_, data_stage_1__5227_, data_stage_1__5226_, data_stage_1__5225_, data_stage_1__5224_, data_stage_1__5223_, data_stage_1__5222_, data_stage_1__5221_, data_stage_1__5220_, data_stage_1__5219_, data_stage_1__5218_, data_stage_1__5217_, data_stage_1__5216_, data_stage_1__5215_, data_stage_1__5214_, data_stage_1__5213_, data_stage_1__5212_, data_stage_1__5211_, data_stage_1__5210_, data_stage_1__5209_, data_stage_1__5208_, data_stage_1__5207_, data_stage_1__5206_, data_stage_1__5205_, data_stage_1__5204_, data_stage_1__5203_, data_stage_1__5202_, data_stage_1__5201_, data_stage_1__5200_, data_stage_1__5199_, data_stage_1__5198_, data_stage_1__5197_, data_stage_1__5196_, data_stage_1__5195_, data_stage_1__5194_, data_stage_1__5193_, data_stage_1__5192_, data_stage_1__5191_, data_stage_1__5190_, data_stage_1__5189_, data_stage_1__5188_, data_stage_1__5187_, data_stage_1__5186_, data_stage_1__5185_, data_stage_1__5184_, data_stage_1__5183_, data_stage_1__5182_, data_stage_1__5181_, data_stage_1__5180_, data_stage_1__5179_, data_stage_1__5178_, data_stage_1__5177_, data_stage_1__5176_, data_stage_1__5175_, data_stage_1__5174_, data_stage_1__5173_, data_stage_1__5172_, data_stage_1__5171_, data_stage_1__5170_, data_stage_1__5169_, data_stage_1__5168_, data_stage_1__5167_, data_stage_1__5166_, data_stage_1__5165_, data_stage_1__5164_, data_stage_1__5163_, data_stage_1__5162_, data_stage_1__5161_, data_stage_1__5160_, data_stage_1__5159_, data_stage_1__5158_, data_stage_1__5157_, data_stage_1__5156_, data_stage_1__5155_, data_stage_1__5154_, data_stage_1__5153_, data_stage_1__5152_, data_stage_1__5151_, data_stage_1__5150_, data_stage_1__5149_, data_stage_1__5148_, data_stage_1__5147_, data_stage_1__5146_, data_stage_1__5145_, data_stage_1__5144_, data_stage_1__5143_, data_stage_1__5142_, data_stage_1__5141_, data_stage_1__5140_, data_stage_1__5139_, data_stage_1__5138_, data_stage_1__5137_, data_stage_1__5136_, data_stage_1__5135_, data_stage_1__5134_, data_stage_1__5133_, data_stage_1__5132_, data_stage_1__5131_, data_stage_1__5130_, data_stage_1__5129_, data_stage_1__5128_, data_stage_1__5127_, data_stage_1__5126_, data_stage_1__5125_, data_stage_1__5124_, data_stage_1__5123_, data_stage_1__5122_, data_stage_1__5121_, data_stage_1__5120_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__5631_, data_stage_2__5630_, data_stage_2__5629_, data_stage_2__5628_, data_stage_2__5627_, data_stage_2__5626_, data_stage_2__5625_, data_stage_2__5624_, data_stage_2__5623_, data_stage_2__5622_, data_stage_2__5621_, data_stage_2__5620_, data_stage_2__5619_, data_stage_2__5618_, data_stage_2__5617_, data_stage_2__5616_, data_stage_2__5615_, data_stage_2__5614_, data_stage_2__5613_, data_stage_2__5612_, data_stage_2__5611_, data_stage_2__5610_, data_stage_2__5609_, data_stage_2__5608_, data_stage_2__5607_, data_stage_2__5606_, data_stage_2__5605_, data_stage_2__5604_, data_stage_2__5603_, data_stage_2__5602_, data_stage_2__5601_, data_stage_2__5600_, data_stage_2__5599_, data_stage_2__5598_, data_stage_2__5597_, data_stage_2__5596_, data_stage_2__5595_, data_stage_2__5594_, data_stage_2__5593_, data_stage_2__5592_, data_stage_2__5591_, data_stage_2__5590_, data_stage_2__5589_, data_stage_2__5588_, data_stage_2__5587_, data_stage_2__5586_, data_stage_2__5585_, data_stage_2__5584_, data_stage_2__5583_, data_stage_2__5582_, data_stage_2__5581_, data_stage_2__5580_, data_stage_2__5579_, data_stage_2__5578_, data_stage_2__5577_, data_stage_2__5576_, data_stage_2__5575_, data_stage_2__5574_, data_stage_2__5573_, data_stage_2__5572_, data_stage_2__5571_, data_stage_2__5570_, data_stage_2__5569_, data_stage_2__5568_, data_stage_2__5567_, data_stage_2__5566_, data_stage_2__5565_, data_stage_2__5564_, data_stage_2__5563_, data_stage_2__5562_, data_stage_2__5561_, data_stage_2__5560_, data_stage_2__5559_, data_stage_2__5558_, data_stage_2__5557_, data_stage_2__5556_, data_stage_2__5555_, data_stage_2__5554_, data_stage_2__5553_, data_stage_2__5552_, data_stage_2__5551_, data_stage_2__5550_, data_stage_2__5549_, data_stage_2__5548_, data_stage_2__5547_, data_stage_2__5546_, data_stage_2__5545_, data_stage_2__5544_, data_stage_2__5543_, data_stage_2__5542_, data_stage_2__5541_, data_stage_2__5540_, data_stage_2__5539_, data_stage_2__5538_, data_stage_2__5537_, data_stage_2__5536_, data_stage_2__5535_, data_stage_2__5534_, data_stage_2__5533_, data_stage_2__5532_, data_stage_2__5531_, data_stage_2__5530_, data_stage_2__5529_, data_stage_2__5528_, data_stage_2__5527_, data_stage_2__5526_, data_stage_2__5525_, data_stage_2__5524_, data_stage_2__5523_, data_stage_2__5522_, data_stage_2__5521_, data_stage_2__5520_, data_stage_2__5519_, data_stage_2__5518_, data_stage_2__5517_, data_stage_2__5516_, data_stage_2__5515_, data_stage_2__5514_, data_stage_2__5513_, data_stage_2__5512_, data_stage_2__5511_, data_stage_2__5510_, data_stage_2__5509_, data_stage_2__5508_, data_stage_2__5507_, data_stage_2__5506_, data_stage_2__5505_, data_stage_2__5504_, data_stage_2__5503_, data_stage_2__5502_, data_stage_2__5501_, data_stage_2__5500_, data_stage_2__5499_, data_stage_2__5498_, data_stage_2__5497_, data_stage_2__5496_, data_stage_2__5495_, data_stage_2__5494_, data_stage_2__5493_, data_stage_2__5492_, data_stage_2__5491_, data_stage_2__5490_, data_stage_2__5489_, data_stage_2__5488_, data_stage_2__5487_, data_stage_2__5486_, data_stage_2__5485_, data_stage_2__5484_, data_stage_2__5483_, data_stage_2__5482_, data_stage_2__5481_, data_stage_2__5480_, data_stage_2__5479_, data_stage_2__5478_, data_stage_2__5477_, data_stage_2__5476_, data_stage_2__5475_, data_stage_2__5474_, data_stage_2__5473_, data_stage_2__5472_, data_stage_2__5471_, data_stage_2__5470_, data_stage_2__5469_, data_stage_2__5468_, data_stage_2__5467_, data_stage_2__5466_, data_stage_2__5465_, data_stage_2__5464_, data_stage_2__5463_, data_stage_2__5462_, data_stage_2__5461_, data_stage_2__5460_, data_stage_2__5459_, data_stage_2__5458_, data_stage_2__5457_, data_stage_2__5456_, data_stage_2__5455_, data_stage_2__5454_, data_stage_2__5453_, data_stage_2__5452_, data_stage_2__5451_, data_stage_2__5450_, data_stage_2__5449_, data_stage_2__5448_, data_stage_2__5447_, data_stage_2__5446_, data_stage_2__5445_, data_stage_2__5444_, data_stage_2__5443_, data_stage_2__5442_, data_stage_2__5441_, data_stage_2__5440_, data_stage_2__5439_, data_stage_2__5438_, data_stage_2__5437_, data_stage_2__5436_, data_stage_2__5435_, data_stage_2__5434_, data_stage_2__5433_, data_stage_2__5432_, data_stage_2__5431_, data_stage_2__5430_, data_stage_2__5429_, data_stage_2__5428_, data_stage_2__5427_, data_stage_2__5426_, data_stage_2__5425_, data_stage_2__5424_, data_stage_2__5423_, data_stage_2__5422_, data_stage_2__5421_, data_stage_2__5420_, data_stage_2__5419_, data_stage_2__5418_, data_stage_2__5417_, data_stage_2__5416_, data_stage_2__5415_, data_stage_2__5414_, data_stage_2__5413_, data_stage_2__5412_, data_stage_2__5411_, data_stage_2__5410_, data_stage_2__5409_, data_stage_2__5408_, data_stage_2__5407_, data_stage_2__5406_, data_stage_2__5405_, data_stage_2__5404_, data_stage_2__5403_, data_stage_2__5402_, data_stage_2__5401_, data_stage_2__5400_, data_stage_2__5399_, data_stage_2__5398_, data_stage_2__5397_, data_stage_2__5396_, data_stage_2__5395_, data_stage_2__5394_, data_stage_2__5393_, data_stage_2__5392_, data_stage_2__5391_, data_stage_2__5390_, data_stage_2__5389_, data_stage_2__5388_, data_stage_2__5387_, data_stage_2__5386_, data_stage_2__5385_, data_stage_2__5384_, data_stage_2__5383_, data_stage_2__5382_, data_stage_2__5381_, data_stage_2__5380_, data_stage_2__5379_, data_stage_2__5378_, data_stage_2__5377_, data_stage_2__5376_, data_stage_2__5375_, data_stage_2__5374_, data_stage_2__5373_, data_stage_2__5372_, data_stage_2__5371_, data_stage_2__5370_, data_stage_2__5369_, data_stage_2__5368_, data_stage_2__5367_, data_stage_2__5366_, data_stage_2__5365_, data_stage_2__5364_, data_stage_2__5363_, data_stage_2__5362_, data_stage_2__5361_, data_stage_2__5360_, data_stage_2__5359_, data_stage_2__5358_, data_stage_2__5357_, data_stage_2__5356_, data_stage_2__5355_, data_stage_2__5354_, data_stage_2__5353_, data_stage_2__5352_, data_stage_2__5351_, data_stage_2__5350_, data_stage_2__5349_, data_stage_2__5348_, data_stage_2__5347_, data_stage_2__5346_, data_stage_2__5345_, data_stage_2__5344_, data_stage_2__5343_, data_stage_2__5342_, data_stage_2__5341_, data_stage_2__5340_, data_stage_2__5339_, data_stage_2__5338_, data_stage_2__5337_, data_stage_2__5336_, data_stage_2__5335_, data_stage_2__5334_, data_stage_2__5333_, data_stage_2__5332_, data_stage_2__5331_, data_stage_2__5330_, data_stage_2__5329_, data_stage_2__5328_, data_stage_2__5327_, data_stage_2__5326_, data_stage_2__5325_, data_stage_2__5324_, data_stage_2__5323_, data_stage_2__5322_, data_stage_2__5321_, data_stage_2__5320_, data_stage_2__5319_, data_stage_2__5318_, data_stage_2__5317_, data_stage_2__5316_, data_stage_2__5315_, data_stage_2__5314_, data_stage_2__5313_, data_stage_2__5312_, data_stage_2__5311_, data_stage_2__5310_, data_stage_2__5309_, data_stage_2__5308_, data_stage_2__5307_, data_stage_2__5306_, data_stage_2__5305_, data_stage_2__5304_, data_stage_2__5303_, data_stage_2__5302_, data_stage_2__5301_, data_stage_2__5300_, data_stage_2__5299_, data_stage_2__5298_, data_stage_2__5297_, data_stage_2__5296_, data_stage_2__5295_, data_stage_2__5294_, data_stage_2__5293_, data_stage_2__5292_, data_stage_2__5291_, data_stage_2__5290_, data_stage_2__5289_, data_stage_2__5288_, data_stage_2__5287_, data_stage_2__5286_, data_stage_2__5285_, data_stage_2__5284_, data_stage_2__5283_, data_stage_2__5282_, data_stage_2__5281_, data_stage_2__5280_, data_stage_2__5279_, data_stage_2__5278_, data_stage_2__5277_, data_stage_2__5276_, data_stage_2__5275_, data_stage_2__5274_, data_stage_2__5273_, data_stage_2__5272_, data_stage_2__5271_, data_stage_2__5270_, data_stage_2__5269_, data_stage_2__5268_, data_stage_2__5267_, data_stage_2__5266_, data_stage_2__5265_, data_stage_2__5264_, data_stage_2__5263_, data_stage_2__5262_, data_stage_2__5261_, data_stage_2__5260_, data_stage_2__5259_, data_stage_2__5258_, data_stage_2__5257_, data_stage_2__5256_, data_stage_2__5255_, data_stage_2__5254_, data_stage_2__5253_, data_stage_2__5252_, data_stage_2__5251_, data_stage_2__5250_, data_stage_2__5249_, data_stage_2__5248_, data_stage_2__5247_, data_stage_2__5246_, data_stage_2__5245_, data_stage_2__5244_, data_stage_2__5243_, data_stage_2__5242_, data_stage_2__5241_, data_stage_2__5240_, data_stage_2__5239_, data_stage_2__5238_, data_stage_2__5237_, data_stage_2__5236_, data_stage_2__5235_, data_stage_2__5234_, data_stage_2__5233_, data_stage_2__5232_, data_stage_2__5231_, data_stage_2__5230_, data_stage_2__5229_, data_stage_2__5228_, data_stage_2__5227_, data_stage_2__5226_, data_stage_2__5225_, data_stage_2__5224_, data_stage_2__5223_, data_stage_2__5222_, data_stage_2__5221_, data_stage_2__5220_, data_stage_2__5219_, data_stage_2__5218_, data_stage_2__5217_, data_stage_2__5216_, data_stage_2__5215_, data_stage_2__5214_, data_stage_2__5213_, data_stage_2__5212_, data_stage_2__5211_, data_stage_2__5210_, data_stage_2__5209_, data_stage_2__5208_, data_stage_2__5207_, data_stage_2__5206_, data_stage_2__5205_, data_stage_2__5204_, data_stage_2__5203_, data_stage_2__5202_, data_stage_2__5201_, data_stage_2__5200_, data_stage_2__5199_, data_stage_2__5198_, data_stage_2__5197_, data_stage_2__5196_, data_stage_2__5195_, data_stage_2__5194_, data_stage_2__5193_, data_stage_2__5192_, data_stage_2__5191_, data_stage_2__5190_, data_stage_2__5189_, data_stage_2__5188_, data_stage_2__5187_, data_stage_2__5186_, data_stage_2__5185_, data_stage_2__5184_, data_stage_2__5183_, data_stage_2__5182_, data_stage_2__5181_, data_stage_2__5180_, data_stage_2__5179_, data_stage_2__5178_, data_stage_2__5177_, data_stage_2__5176_, data_stage_2__5175_, data_stage_2__5174_, data_stage_2__5173_, data_stage_2__5172_, data_stage_2__5171_, data_stage_2__5170_, data_stage_2__5169_, data_stage_2__5168_, data_stage_2__5167_, data_stage_2__5166_, data_stage_2__5165_, data_stage_2__5164_, data_stage_2__5163_, data_stage_2__5162_, data_stage_2__5161_, data_stage_2__5160_, data_stage_2__5159_, data_stage_2__5158_, data_stage_2__5157_, data_stage_2__5156_, data_stage_2__5155_, data_stage_2__5154_, data_stage_2__5153_, data_stage_2__5152_, data_stage_2__5151_, data_stage_2__5150_, data_stage_2__5149_, data_stage_2__5148_, data_stage_2__5147_, data_stage_2__5146_, data_stage_2__5145_, data_stage_2__5144_, data_stage_2__5143_, data_stage_2__5142_, data_stage_2__5141_, data_stage_2__5140_, data_stage_2__5139_, data_stage_2__5138_, data_stage_2__5137_, data_stage_2__5136_, data_stage_2__5135_, data_stage_2__5134_, data_stage_2__5133_, data_stage_2__5132_, data_stage_2__5131_, data_stage_2__5130_, data_stage_2__5129_, data_stage_2__5128_, data_stage_2__5127_, data_stage_2__5126_, data_stage_2__5125_, data_stage_2__5124_, data_stage_2__5123_, data_stage_2__5122_, data_stage_2__5121_, data_stage_2__5120_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_11__swap_inst
  (
    .data_i({ data_stage_1__6143_, data_stage_1__6142_, data_stage_1__6141_, data_stage_1__6140_, data_stage_1__6139_, data_stage_1__6138_, data_stage_1__6137_, data_stage_1__6136_, data_stage_1__6135_, data_stage_1__6134_, data_stage_1__6133_, data_stage_1__6132_, data_stage_1__6131_, data_stage_1__6130_, data_stage_1__6129_, data_stage_1__6128_, data_stage_1__6127_, data_stage_1__6126_, data_stage_1__6125_, data_stage_1__6124_, data_stage_1__6123_, data_stage_1__6122_, data_stage_1__6121_, data_stage_1__6120_, data_stage_1__6119_, data_stage_1__6118_, data_stage_1__6117_, data_stage_1__6116_, data_stage_1__6115_, data_stage_1__6114_, data_stage_1__6113_, data_stage_1__6112_, data_stage_1__6111_, data_stage_1__6110_, data_stage_1__6109_, data_stage_1__6108_, data_stage_1__6107_, data_stage_1__6106_, data_stage_1__6105_, data_stage_1__6104_, data_stage_1__6103_, data_stage_1__6102_, data_stage_1__6101_, data_stage_1__6100_, data_stage_1__6099_, data_stage_1__6098_, data_stage_1__6097_, data_stage_1__6096_, data_stage_1__6095_, data_stage_1__6094_, data_stage_1__6093_, data_stage_1__6092_, data_stage_1__6091_, data_stage_1__6090_, data_stage_1__6089_, data_stage_1__6088_, data_stage_1__6087_, data_stage_1__6086_, data_stage_1__6085_, data_stage_1__6084_, data_stage_1__6083_, data_stage_1__6082_, data_stage_1__6081_, data_stage_1__6080_, data_stage_1__6079_, data_stage_1__6078_, data_stage_1__6077_, data_stage_1__6076_, data_stage_1__6075_, data_stage_1__6074_, data_stage_1__6073_, data_stage_1__6072_, data_stage_1__6071_, data_stage_1__6070_, data_stage_1__6069_, data_stage_1__6068_, data_stage_1__6067_, data_stage_1__6066_, data_stage_1__6065_, data_stage_1__6064_, data_stage_1__6063_, data_stage_1__6062_, data_stage_1__6061_, data_stage_1__6060_, data_stage_1__6059_, data_stage_1__6058_, data_stage_1__6057_, data_stage_1__6056_, data_stage_1__6055_, data_stage_1__6054_, data_stage_1__6053_, data_stage_1__6052_, data_stage_1__6051_, data_stage_1__6050_, data_stage_1__6049_, data_stage_1__6048_, data_stage_1__6047_, data_stage_1__6046_, data_stage_1__6045_, data_stage_1__6044_, data_stage_1__6043_, data_stage_1__6042_, data_stage_1__6041_, data_stage_1__6040_, data_stage_1__6039_, data_stage_1__6038_, data_stage_1__6037_, data_stage_1__6036_, data_stage_1__6035_, data_stage_1__6034_, data_stage_1__6033_, data_stage_1__6032_, data_stage_1__6031_, data_stage_1__6030_, data_stage_1__6029_, data_stage_1__6028_, data_stage_1__6027_, data_stage_1__6026_, data_stage_1__6025_, data_stage_1__6024_, data_stage_1__6023_, data_stage_1__6022_, data_stage_1__6021_, data_stage_1__6020_, data_stage_1__6019_, data_stage_1__6018_, data_stage_1__6017_, data_stage_1__6016_, data_stage_1__6015_, data_stage_1__6014_, data_stage_1__6013_, data_stage_1__6012_, data_stage_1__6011_, data_stage_1__6010_, data_stage_1__6009_, data_stage_1__6008_, data_stage_1__6007_, data_stage_1__6006_, data_stage_1__6005_, data_stage_1__6004_, data_stage_1__6003_, data_stage_1__6002_, data_stage_1__6001_, data_stage_1__6000_, data_stage_1__5999_, data_stage_1__5998_, data_stage_1__5997_, data_stage_1__5996_, data_stage_1__5995_, data_stage_1__5994_, data_stage_1__5993_, data_stage_1__5992_, data_stage_1__5991_, data_stage_1__5990_, data_stage_1__5989_, data_stage_1__5988_, data_stage_1__5987_, data_stage_1__5986_, data_stage_1__5985_, data_stage_1__5984_, data_stage_1__5983_, data_stage_1__5982_, data_stage_1__5981_, data_stage_1__5980_, data_stage_1__5979_, data_stage_1__5978_, data_stage_1__5977_, data_stage_1__5976_, data_stage_1__5975_, data_stage_1__5974_, data_stage_1__5973_, data_stage_1__5972_, data_stage_1__5971_, data_stage_1__5970_, data_stage_1__5969_, data_stage_1__5968_, data_stage_1__5967_, data_stage_1__5966_, data_stage_1__5965_, data_stage_1__5964_, data_stage_1__5963_, data_stage_1__5962_, data_stage_1__5961_, data_stage_1__5960_, data_stage_1__5959_, data_stage_1__5958_, data_stage_1__5957_, data_stage_1__5956_, data_stage_1__5955_, data_stage_1__5954_, data_stage_1__5953_, data_stage_1__5952_, data_stage_1__5951_, data_stage_1__5950_, data_stage_1__5949_, data_stage_1__5948_, data_stage_1__5947_, data_stage_1__5946_, data_stage_1__5945_, data_stage_1__5944_, data_stage_1__5943_, data_stage_1__5942_, data_stage_1__5941_, data_stage_1__5940_, data_stage_1__5939_, data_stage_1__5938_, data_stage_1__5937_, data_stage_1__5936_, data_stage_1__5935_, data_stage_1__5934_, data_stage_1__5933_, data_stage_1__5932_, data_stage_1__5931_, data_stage_1__5930_, data_stage_1__5929_, data_stage_1__5928_, data_stage_1__5927_, data_stage_1__5926_, data_stage_1__5925_, data_stage_1__5924_, data_stage_1__5923_, data_stage_1__5922_, data_stage_1__5921_, data_stage_1__5920_, data_stage_1__5919_, data_stage_1__5918_, data_stage_1__5917_, data_stage_1__5916_, data_stage_1__5915_, data_stage_1__5914_, data_stage_1__5913_, data_stage_1__5912_, data_stage_1__5911_, data_stage_1__5910_, data_stage_1__5909_, data_stage_1__5908_, data_stage_1__5907_, data_stage_1__5906_, data_stage_1__5905_, data_stage_1__5904_, data_stage_1__5903_, data_stage_1__5902_, data_stage_1__5901_, data_stage_1__5900_, data_stage_1__5899_, data_stage_1__5898_, data_stage_1__5897_, data_stage_1__5896_, data_stage_1__5895_, data_stage_1__5894_, data_stage_1__5893_, data_stage_1__5892_, data_stage_1__5891_, data_stage_1__5890_, data_stage_1__5889_, data_stage_1__5888_, data_stage_1__5887_, data_stage_1__5886_, data_stage_1__5885_, data_stage_1__5884_, data_stage_1__5883_, data_stage_1__5882_, data_stage_1__5881_, data_stage_1__5880_, data_stage_1__5879_, data_stage_1__5878_, data_stage_1__5877_, data_stage_1__5876_, data_stage_1__5875_, data_stage_1__5874_, data_stage_1__5873_, data_stage_1__5872_, data_stage_1__5871_, data_stage_1__5870_, data_stage_1__5869_, data_stage_1__5868_, data_stage_1__5867_, data_stage_1__5866_, data_stage_1__5865_, data_stage_1__5864_, data_stage_1__5863_, data_stage_1__5862_, data_stage_1__5861_, data_stage_1__5860_, data_stage_1__5859_, data_stage_1__5858_, data_stage_1__5857_, data_stage_1__5856_, data_stage_1__5855_, data_stage_1__5854_, data_stage_1__5853_, data_stage_1__5852_, data_stage_1__5851_, data_stage_1__5850_, data_stage_1__5849_, data_stage_1__5848_, data_stage_1__5847_, data_stage_1__5846_, data_stage_1__5845_, data_stage_1__5844_, data_stage_1__5843_, data_stage_1__5842_, data_stage_1__5841_, data_stage_1__5840_, data_stage_1__5839_, data_stage_1__5838_, data_stage_1__5837_, data_stage_1__5836_, data_stage_1__5835_, data_stage_1__5834_, data_stage_1__5833_, data_stage_1__5832_, data_stage_1__5831_, data_stage_1__5830_, data_stage_1__5829_, data_stage_1__5828_, data_stage_1__5827_, data_stage_1__5826_, data_stage_1__5825_, data_stage_1__5824_, data_stage_1__5823_, data_stage_1__5822_, data_stage_1__5821_, data_stage_1__5820_, data_stage_1__5819_, data_stage_1__5818_, data_stage_1__5817_, data_stage_1__5816_, data_stage_1__5815_, data_stage_1__5814_, data_stage_1__5813_, data_stage_1__5812_, data_stage_1__5811_, data_stage_1__5810_, data_stage_1__5809_, data_stage_1__5808_, data_stage_1__5807_, data_stage_1__5806_, data_stage_1__5805_, data_stage_1__5804_, data_stage_1__5803_, data_stage_1__5802_, data_stage_1__5801_, data_stage_1__5800_, data_stage_1__5799_, data_stage_1__5798_, data_stage_1__5797_, data_stage_1__5796_, data_stage_1__5795_, data_stage_1__5794_, data_stage_1__5793_, data_stage_1__5792_, data_stage_1__5791_, data_stage_1__5790_, data_stage_1__5789_, data_stage_1__5788_, data_stage_1__5787_, data_stage_1__5786_, data_stage_1__5785_, data_stage_1__5784_, data_stage_1__5783_, data_stage_1__5782_, data_stage_1__5781_, data_stage_1__5780_, data_stage_1__5779_, data_stage_1__5778_, data_stage_1__5777_, data_stage_1__5776_, data_stage_1__5775_, data_stage_1__5774_, data_stage_1__5773_, data_stage_1__5772_, data_stage_1__5771_, data_stage_1__5770_, data_stage_1__5769_, data_stage_1__5768_, data_stage_1__5767_, data_stage_1__5766_, data_stage_1__5765_, data_stage_1__5764_, data_stage_1__5763_, data_stage_1__5762_, data_stage_1__5761_, data_stage_1__5760_, data_stage_1__5759_, data_stage_1__5758_, data_stage_1__5757_, data_stage_1__5756_, data_stage_1__5755_, data_stage_1__5754_, data_stage_1__5753_, data_stage_1__5752_, data_stage_1__5751_, data_stage_1__5750_, data_stage_1__5749_, data_stage_1__5748_, data_stage_1__5747_, data_stage_1__5746_, data_stage_1__5745_, data_stage_1__5744_, data_stage_1__5743_, data_stage_1__5742_, data_stage_1__5741_, data_stage_1__5740_, data_stage_1__5739_, data_stage_1__5738_, data_stage_1__5737_, data_stage_1__5736_, data_stage_1__5735_, data_stage_1__5734_, data_stage_1__5733_, data_stage_1__5732_, data_stage_1__5731_, data_stage_1__5730_, data_stage_1__5729_, data_stage_1__5728_, data_stage_1__5727_, data_stage_1__5726_, data_stage_1__5725_, data_stage_1__5724_, data_stage_1__5723_, data_stage_1__5722_, data_stage_1__5721_, data_stage_1__5720_, data_stage_1__5719_, data_stage_1__5718_, data_stage_1__5717_, data_stage_1__5716_, data_stage_1__5715_, data_stage_1__5714_, data_stage_1__5713_, data_stage_1__5712_, data_stage_1__5711_, data_stage_1__5710_, data_stage_1__5709_, data_stage_1__5708_, data_stage_1__5707_, data_stage_1__5706_, data_stage_1__5705_, data_stage_1__5704_, data_stage_1__5703_, data_stage_1__5702_, data_stage_1__5701_, data_stage_1__5700_, data_stage_1__5699_, data_stage_1__5698_, data_stage_1__5697_, data_stage_1__5696_, data_stage_1__5695_, data_stage_1__5694_, data_stage_1__5693_, data_stage_1__5692_, data_stage_1__5691_, data_stage_1__5690_, data_stage_1__5689_, data_stage_1__5688_, data_stage_1__5687_, data_stage_1__5686_, data_stage_1__5685_, data_stage_1__5684_, data_stage_1__5683_, data_stage_1__5682_, data_stage_1__5681_, data_stage_1__5680_, data_stage_1__5679_, data_stage_1__5678_, data_stage_1__5677_, data_stage_1__5676_, data_stage_1__5675_, data_stage_1__5674_, data_stage_1__5673_, data_stage_1__5672_, data_stage_1__5671_, data_stage_1__5670_, data_stage_1__5669_, data_stage_1__5668_, data_stage_1__5667_, data_stage_1__5666_, data_stage_1__5665_, data_stage_1__5664_, data_stage_1__5663_, data_stage_1__5662_, data_stage_1__5661_, data_stage_1__5660_, data_stage_1__5659_, data_stage_1__5658_, data_stage_1__5657_, data_stage_1__5656_, data_stage_1__5655_, data_stage_1__5654_, data_stage_1__5653_, data_stage_1__5652_, data_stage_1__5651_, data_stage_1__5650_, data_stage_1__5649_, data_stage_1__5648_, data_stage_1__5647_, data_stage_1__5646_, data_stage_1__5645_, data_stage_1__5644_, data_stage_1__5643_, data_stage_1__5642_, data_stage_1__5641_, data_stage_1__5640_, data_stage_1__5639_, data_stage_1__5638_, data_stage_1__5637_, data_stage_1__5636_, data_stage_1__5635_, data_stage_1__5634_, data_stage_1__5633_, data_stage_1__5632_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__6143_, data_stage_2__6142_, data_stage_2__6141_, data_stage_2__6140_, data_stage_2__6139_, data_stage_2__6138_, data_stage_2__6137_, data_stage_2__6136_, data_stage_2__6135_, data_stage_2__6134_, data_stage_2__6133_, data_stage_2__6132_, data_stage_2__6131_, data_stage_2__6130_, data_stage_2__6129_, data_stage_2__6128_, data_stage_2__6127_, data_stage_2__6126_, data_stage_2__6125_, data_stage_2__6124_, data_stage_2__6123_, data_stage_2__6122_, data_stage_2__6121_, data_stage_2__6120_, data_stage_2__6119_, data_stage_2__6118_, data_stage_2__6117_, data_stage_2__6116_, data_stage_2__6115_, data_stage_2__6114_, data_stage_2__6113_, data_stage_2__6112_, data_stage_2__6111_, data_stage_2__6110_, data_stage_2__6109_, data_stage_2__6108_, data_stage_2__6107_, data_stage_2__6106_, data_stage_2__6105_, data_stage_2__6104_, data_stage_2__6103_, data_stage_2__6102_, data_stage_2__6101_, data_stage_2__6100_, data_stage_2__6099_, data_stage_2__6098_, data_stage_2__6097_, data_stage_2__6096_, data_stage_2__6095_, data_stage_2__6094_, data_stage_2__6093_, data_stage_2__6092_, data_stage_2__6091_, data_stage_2__6090_, data_stage_2__6089_, data_stage_2__6088_, data_stage_2__6087_, data_stage_2__6086_, data_stage_2__6085_, data_stage_2__6084_, data_stage_2__6083_, data_stage_2__6082_, data_stage_2__6081_, data_stage_2__6080_, data_stage_2__6079_, data_stage_2__6078_, data_stage_2__6077_, data_stage_2__6076_, data_stage_2__6075_, data_stage_2__6074_, data_stage_2__6073_, data_stage_2__6072_, data_stage_2__6071_, data_stage_2__6070_, data_stage_2__6069_, data_stage_2__6068_, data_stage_2__6067_, data_stage_2__6066_, data_stage_2__6065_, data_stage_2__6064_, data_stage_2__6063_, data_stage_2__6062_, data_stage_2__6061_, data_stage_2__6060_, data_stage_2__6059_, data_stage_2__6058_, data_stage_2__6057_, data_stage_2__6056_, data_stage_2__6055_, data_stage_2__6054_, data_stage_2__6053_, data_stage_2__6052_, data_stage_2__6051_, data_stage_2__6050_, data_stage_2__6049_, data_stage_2__6048_, data_stage_2__6047_, data_stage_2__6046_, data_stage_2__6045_, data_stage_2__6044_, data_stage_2__6043_, data_stage_2__6042_, data_stage_2__6041_, data_stage_2__6040_, data_stage_2__6039_, data_stage_2__6038_, data_stage_2__6037_, data_stage_2__6036_, data_stage_2__6035_, data_stage_2__6034_, data_stage_2__6033_, data_stage_2__6032_, data_stage_2__6031_, data_stage_2__6030_, data_stage_2__6029_, data_stage_2__6028_, data_stage_2__6027_, data_stage_2__6026_, data_stage_2__6025_, data_stage_2__6024_, data_stage_2__6023_, data_stage_2__6022_, data_stage_2__6021_, data_stage_2__6020_, data_stage_2__6019_, data_stage_2__6018_, data_stage_2__6017_, data_stage_2__6016_, data_stage_2__6015_, data_stage_2__6014_, data_stage_2__6013_, data_stage_2__6012_, data_stage_2__6011_, data_stage_2__6010_, data_stage_2__6009_, data_stage_2__6008_, data_stage_2__6007_, data_stage_2__6006_, data_stage_2__6005_, data_stage_2__6004_, data_stage_2__6003_, data_stage_2__6002_, data_stage_2__6001_, data_stage_2__6000_, data_stage_2__5999_, data_stage_2__5998_, data_stage_2__5997_, data_stage_2__5996_, data_stage_2__5995_, data_stage_2__5994_, data_stage_2__5993_, data_stage_2__5992_, data_stage_2__5991_, data_stage_2__5990_, data_stage_2__5989_, data_stage_2__5988_, data_stage_2__5987_, data_stage_2__5986_, data_stage_2__5985_, data_stage_2__5984_, data_stage_2__5983_, data_stage_2__5982_, data_stage_2__5981_, data_stage_2__5980_, data_stage_2__5979_, data_stage_2__5978_, data_stage_2__5977_, data_stage_2__5976_, data_stage_2__5975_, data_stage_2__5974_, data_stage_2__5973_, data_stage_2__5972_, data_stage_2__5971_, data_stage_2__5970_, data_stage_2__5969_, data_stage_2__5968_, data_stage_2__5967_, data_stage_2__5966_, data_stage_2__5965_, data_stage_2__5964_, data_stage_2__5963_, data_stage_2__5962_, data_stage_2__5961_, data_stage_2__5960_, data_stage_2__5959_, data_stage_2__5958_, data_stage_2__5957_, data_stage_2__5956_, data_stage_2__5955_, data_stage_2__5954_, data_stage_2__5953_, data_stage_2__5952_, data_stage_2__5951_, data_stage_2__5950_, data_stage_2__5949_, data_stage_2__5948_, data_stage_2__5947_, data_stage_2__5946_, data_stage_2__5945_, data_stage_2__5944_, data_stage_2__5943_, data_stage_2__5942_, data_stage_2__5941_, data_stage_2__5940_, data_stage_2__5939_, data_stage_2__5938_, data_stage_2__5937_, data_stage_2__5936_, data_stage_2__5935_, data_stage_2__5934_, data_stage_2__5933_, data_stage_2__5932_, data_stage_2__5931_, data_stage_2__5930_, data_stage_2__5929_, data_stage_2__5928_, data_stage_2__5927_, data_stage_2__5926_, data_stage_2__5925_, data_stage_2__5924_, data_stage_2__5923_, data_stage_2__5922_, data_stage_2__5921_, data_stage_2__5920_, data_stage_2__5919_, data_stage_2__5918_, data_stage_2__5917_, data_stage_2__5916_, data_stage_2__5915_, data_stage_2__5914_, data_stage_2__5913_, data_stage_2__5912_, data_stage_2__5911_, data_stage_2__5910_, data_stage_2__5909_, data_stage_2__5908_, data_stage_2__5907_, data_stage_2__5906_, data_stage_2__5905_, data_stage_2__5904_, data_stage_2__5903_, data_stage_2__5902_, data_stage_2__5901_, data_stage_2__5900_, data_stage_2__5899_, data_stage_2__5898_, data_stage_2__5897_, data_stage_2__5896_, data_stage_2__5895_, data_stage_2__5894_, data_stage_2__5893_, data_stage_2__5892_, data_stage_2__5891_, data_stage_2__5890_, data_stage_2__5889_, data_stage_2__5888_, data_stage_2__5887_, data_stage_2__5886_, data_stage_2__5885_, data_stage_2__5884_, data_stage_2__5883_, data_stage_2__5882_, data_stage_2__5881_, data_stage_2__5880_, data_stage_2__5879_, data_stage_2__5878_, data_stage_2__5877_, data_stage_2__5876_, data_stage_2__5875_, data_stage_2__5874_, data_stage_2__5873_, data_stage_2__5872_, data_stage_2__5871_, data_stage_2__5870_, data_stage_2__5869_, data_stage_2__5868_, data_stage_2__5867_, data_stage_2__5866_, data_stage_2__5865_, data_stage_2__5864_, data_stage_2__5863_, data_stage_2__5862_, data_stage_2__5861_, data_stage_2__5860_, data_stage_2__5859_, data_stage_2__5858_, data_stage_2__5857_, data_stage_2__5856_, data_stage_2__5855_, data_stage_2__5854_, data_stage_2__5853_, data_stage_2__5852_, data_stage_2__5851_, data_stage_2__5850_, data_stage_2__5849_, data_stage_2__5848_, data_stage_2__5847_, data_stage_2__5846_, data_stage_2__5845_, data_stage_2__5844_, data_stage_2__5843_, data_stage_2__5842_, data_stage_2__5841_, data_stage_2__5840_, data_stage_2__5839_, data_stage_2__5838_, data_stage_2__5837_, data_stage_2__5836_, data_stage_2__5835_, data_stage_2__5834_, data_stage_2__5833_, data_stage_2__5832_, data_stage_2__5831_, data_stage_2__5830_, data_stage_2__5829_, data_stage_2__5828_, data_stage_2__5827_, data_stage_2__5826_, data_stage_2__5825_, data_stage_2__5824_, data_stage_2__5823_, data_stage_2__5822_, data_stage_2__5821_, data_stage_2__5820_, data_stage_2__5819_, data_stage_2__5818_, data_stage_2__5817_, data_stage_2__5816_, data_stage_2__5815_, data_stage_2__5814_, data_stage_2__5813_, data_stage_2__5812_, data_stage_2__5811_, data_stage_2__5810_, data_stage_2__5809_, data_stage_2__5808_, data_stage_2__5807_, data_stage_2__5806_, data_stage_2__5805_, data_stage_2__5804_, data_stage_2__5803_, data_stage_2__5802_, data_stage_2__5801_, data_stage_2__5800_, data_stage_2__5799_, data_stage_2__5798_, data_stage_2__5797_, data_stage_2__5796_, data_stage_2__5795_, data_stage_2__5794_, data_stage_2__5793_, data_stage_2__5792_, data_stage_2__5791_, data_stage_2__5790_, data_stage_2__5789_, data_stage_2__5788_, data_stage_2__5787_, data_stage_2__5786_, data_stage_2__5785_, data_stage_2__5784_, data_stage_2__5783_, data_stage_2__5782_, data_stage_2__5781_, data_stage_2__5780_, data_stage_2__5779_, data_stage_2__5778_, data_stage_2__5777_, data_stage_2__5776_, data_stage_2__5775_, data_stage_2__5774_, data_stage_2__5773_, data_stage_2__5772_, data_stage_2__5771_, data_stage_2__5770_, data_stage_2__5769_, data_stage_2__5768_, data_stage_2__5767_, data_stage_2__5766_, data_stage_2__5765_, data_stage_2__5764_, data_stage_2__5763_, data_stage_2__5762_, data_stage_2__5761_, data_stage_2__5760_, data_stage_2__5759_, data_stage_2__5758_, data_stage_2__5757_, data_stage_2__5756_, data_stage_2__5755_, data_stage_2__5754_, data_stage_2__5753_, data_stage_2__5752_, data_stage_2__5751_, data_stage_2__5750_, data_stage_2__5749_, data_stage_2__5748_, data_stage_2__5747_, data_stage_2__5746_, data_stage_2__5745_, data_stage_2__5744_, data_stage_2__5743_, data_stage_2__5742_, data_stage_2__5741_, data_stage_2__5740_, data_stage_2__5739_, data_stage_2__5738_, data_stage_2__5737_, data_stage_2__5736_, data_stage_2__5735_, data_stage_2__5734_, data_stage_2__5733_, data_stage_2__5732_, data_stage_2__5731_, data_stage_2__5730_, data_stage_2__5729_, data_stage_2__5728_, data_stage_2__5727_, data_stage_2__5726_, data_stage_2__5725_, data_stage_2__5724_, data_stage_2__5723_, data_stage_2__5722_, data_stage_2__5721_, data_stage_2__5720_, data_stage_2__5719_, data_stage_2__5718_, data_stage_2__5717_, data_stage_2__5716_, data_stage_2__5715_, data_stage_2__5714_, data_stage_2__5713_, data_stage_2__5712_, data_stage_2__5711_, data_stage_2__5710_, data_stage_2__5709_, data_stage_2__5708_, data_stage_2__5707_, data_stage_2__5706_, data_stage_2__5705_, data_stage_2__5704_, data_stage_2__5703_, data_stage_2__5702_, data_stage_2__5701_, data_stage_2__5700_, data_stage_2__5699_, data_stage_2__5698_, data_stage_2__5697_, data_stage_2__5696_, data_stage_2__5695_, data_stage_2__5694_, data_stage_2__5693_, data_stage_2__5692_, data_stage_2__5691_, data_stage_2__5690_, data_stage_2__5689_, data_stage_2__5688_, data_stage_2__5687_, data_stage_2__5686_, data_stage_2__5685_, data_stage_2__5684_, data_stage_2__5683_, data_stage_2__5682_, data_stage_2__5681_, data_stage_2__5680_, data_stage_2__5679_, data_stage_2__5678_, data_stage_2__5677_, data_stage_2__5676_, data_stage_2__5675_, data_stage_2__5674_, data_stage_2__5673_, data_stage_2__5672_, data_stage_2__5671_, data_stage_2__5670_, data_stage_2__5669_, data_stage_2__5668_, data_stage_2__5667_, data_stage_2__5666_, data_stage_2__5665_, data_stage_2__5664_, data_stage_2__5663_, data_stage_2__5662_, data_stage_2__5661_, data_stage_2__5660_, data_stage_2__5659_, data_stage_2__5658_, data_stage_2__5657_, data_stage_2__5656_, data_stage_2__5655_, data_stage_2__5654_, data_stage_2__5653_, data_stage_2__5652_, data_stage_2__5651_, data_stage_2__5650_, data_stage_2__5649_, data_stage_2__5648_, data_stage_2__5647_, data_stage_2__5646_, data_stage_2__5645_, data_stage_2__5644_, data_stage_2__5643_, data_stage_2__5642_, data_stage_2__5641_, data_stage_2__5640_, data_stage_2__5639_, data_stage_2__5638_, data_stage_2__5637_, data_stage_2__5636_, data_stage_2__5635_, data_stage_2__5634_, data_stage_2__5633_, data_stage_2__5632_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_12__swap_inst
  (
    .data_i({ data_stage_1__6655_, data_stage_1__6654_, data_stage_1__6653_, data_stage_1__6652_, data_stage_1__6651_, data_stage_1__6650_, data_stage_1__6649_, data_stage_1__6648_, data_stage_1__6647_, data_stage_1__6646_, data_stage_1__6645_, data_stage_1__6644_, data_stage_1__6643_, data_stage_1__6642_, data_stage_1__6641_, data_stage_1__6640_, data_stage_1__6639_, data_stage_1__6638_, data_stage_1__6637_, data_stage_1__6636_, data_stage_1__6635_, data_stage_1__6634_, data_stage_1__6633_, data_stage_1__6632_, data_stage_1__6631_, data_stage_1__6630_, data_stage_1__6629_, data_stage_1__6628_, data_stage_1__6627_, data_stage_1__6626_, data_stage_1__6625_, data_stage_1__6624_, data_stage_1__6623_, data_stage_1__6622_, data_stage_1__6621_, data_stage_1__6620_, data_stage_1__6619_, data_stage_1__6618_, data_stage_1__6617_, data_stage_1__6616_, data_stage_1__6615_, data_stage_1__6614_, data_stage_1__6613_, data_stage_1__6612_, data_stage_1__6611_, data_stage_1__6610_, data_stage_1__6609_, data_stage_1__6608_, data_stage_1__6607_, data_stage_1__6606_, data_stage_1__6605_, data_stage_1__6604_, data_stage_1__6603_, data_stage_1__6602_, data_stage_1__6601_, data_stage_1__6600_, data_stage_1__6599_, data_stage_1__6598_, data_stage_1__6597_, data_stage_1__6596_, data_stage_1__6595_, data_stage_1__6594_, data_stage_1__6593_, data_stage_1__6592_, data_stage_1__6591_, data_stage_1__6590_, data_stage_1__6589_, data_stage_1__6588_, data_stage_1__6587_, data_stage_1__6586_, data_stage_1__6585_, data_stage_1__6584_, data_stage_1__6583_, data_stage_1__6582_, data_stage_1__6581_, data_stage_1__6580_, data_stage_1__6579_, data_stage_1__6578_, data_stage_1__6577_, data_stage_1__6576_, data_stage_1__6575_, data_stage_1__6574_, data_stage_1__6573_, data_stage_1__6572_, data_stage_1__6571_, data_stage_1__6570_, data_stage_1__6569_, data_stage_1__6568_, data_stage_1__6567_, data_stage_1__6566_, data_stage_1__6565_, data_stage_1__6564_, data_stage_1__6563_, data_stage_1__6562_, data_stage_1__6561_, data_stage_1__6560_, data_stage_1__6559_, data_stage_1__6558_, data_stage_1__6557_, data_stage_1__6556_, data_stage_1__6555_, data_stage_1__6554_, data_stage_1__6553_, data_stage_1__6552_, data_stage_1__6551_, data_stage_1__6550_, data_stage_1__6549_, data_stage_1__6548_, data_stage_1__6547_, data_stage_1__6546_, data_stage_1__6545_, data_stage_1__6544_, data_stage_1__6543_, data_stage_1__6542_, data_stage_1__6541_, data_stage_1__6540_, data_stage_1__6539_, data_stage_1__6538_, data_stage_1__6537_, data_stage_1__6536_, data_stage_1__6535_, data_stage_1__6534_, data_stage_1__6533_, data_stage_1__6532_, data_stage_1__6531_, data_stage_1__6530_, data_stage_1__6529_, data_stage_1__6528_, data_stage_1__6527_, data_stage_1__6526_, data_stage_1__6525_, data_stage_1__6524_, data_stage_1__6523_, data_stage_1__6522_, data_stage_1__6521_, data_stage_1__6520_, data_stage_1__6519_, data_stage_1__6518_, data_stage_1__6517_, data_stage_1__6516_, data_stage_1__6515_, data_stage_1__6514_, data_stage_1__6513_, data_stage_1__6512_, data_stage_1__6511_, data_stage_1__6510_, data_stage_1__6509_, data_stage_1__6508_, data_stage_1__6507_, data_stage_1__6506_, data_stage_1__6505_, data_stage_1__6504_, data_stage_1__6503_, data_stage_1__6502_, data_stage_1__6501_, data_stage_1__6500_, data_stage_1__6499_, data_stage_1__6498_, data_stage_1__6497_, data_stage_1__6496_, data_stage_1__6495_, data_stage_1__6494_, data_stage_1__6493_, data_stage_1__6492_, data_stage_1__6491_, data_stage_1__6490_, data_stage_1__6489_, data_stage_1__6488_, data_stage_1__6487_, data_stage_1__6486_, data_stage_1__6485_, data_stage_1__6484_, data_stage_1__6483_, data_stage_1__6482_, data_stage_1__6481_, data_stage_1__6480_, data_stage_1__6479_, data_stage_1__6478_, data_stage_1__6477_, data_stage_1__6476_, data_stage_1__6475_, data_stage_1__6474_, data_stage_1__6473_, data_stage_1__6472_, data_stage_1__6471_, data_stage_1__6470_, data_stage_1__6469_, data_stage_1__6468_, data_stage_1__6467_, data_stage_1__6466_, data_stage_1__6465_, data_stage_1__6464_, data_stage_1__6463_, data_stage_1__6462_, data_stage_1__6461_, data_stage_1__6460_, data_stage_1__6459_, data_stage_1__6458_, data_stage_1__6457_, data_stage_1__6456_, data_stage_1__6455_, data_stage_1__6454_, data_stage_1__6453_, data_stage_1__6452_, data_stage_1__6451_, data_stage_1__6450_, data_stage_1__6449_, data_stage_1__6448_, data_stage_1__6447_, data_stage_1__6446_, data_stage_1__6445_, data_stage_1__6444_, data_stage_1__6443_, data_stage_1__6442_, data_stage_1__6441_, data_stage_1__6440_, data_stage_1__6439_, data_stage_1__6438_, data_stage_1__6437_, data_stage_1__6436_, data_stage_1__6435_, data_stage_1__6434_, data_stage_1__6433_, data_stage_1__6432_, data_stage_1__6431_, data_stage_1__6430_, data_stage_1__6429_, data_stage_1__6428_, data_stage_1__6427_, data_stage_1__6426_, data_stage_1__6425_, data_stage_1__6424_, data_stage_1__6423_, data_stage_1__6422_, data_stage_1__6421_, data_stage_1__6420_, data_stage_1__6419_, data_stage_1__6418_, data_stage_1__6417_, data_stage_1__6416_, data_stage_1__6415_, data_stage_1__6414_, data_stage_1__6413_, data_stage_1__6412_, data_stage_1__6411_, data_stage_1__6410_, data_stage_1__6409_, data_stage_1__6408_, data_stage_1__6407_, data_stage_1__6406_, data_stage_1__6405_, data_stage_1__6404_, data_stage_1__6403_, data_stage_1__6402_, data_stage_1__6401_, data_stage_1__6400_, data_stage_1__6399_, data_stage_1__6398_, data_stage_1__6397_, data_stage_1__6396_, data_stage_1__6395_, data_stage_1__6394_, data_stage_1__6393_, data_stage_1__6392_, data_stage_1__6391_, data_stage_1__6390_, data_stage_1__6389_, data_stage_1__6388_, data_stage_1__6387_, data_stage_1__6386_, data_stage_1__6385_, data_stage_1__6384_, data_stage_1__6383_, data_stage_1__6382_, data_stage_1__6381_, data_stage_1__6380_, data_stage_1__6379_, data_stage_1__6378_, data_stage_1__6377_, data_stage_1__6376_, data_stage_1__6375_, data_stage_1__6374_, data_stage_1__6373_, data_stage_1__6372_, data_stage_1__6371_, data_stage_1__6370_, data_stage_1__6369_, data_stage_1__6368_, data_stage_1__6367_, data_stage_1__6366_, data_stage_1__6365_, data_stage_1__6364_, data_stage_1__6363_, data_stage_1__6362_, data_stage_1__6361_, data_stage_1__6360_, data_stage_1__6359_, data_stage_1__6358_, data_stage_1__6357_, data_stage_1__6356_, data_stage_1__6355_, data_stage_1__6354_, data_stage_1__6353_, data_stage_1__6352_, data_stage_1__6351_, data_stage_1__6350_, data_stage_1__6349_, data_stage_1__6348_, data_stage_1__6347_, data_stage_1__6346_, data_stage_1__6345_, data_stage_1__6344_, data_stage_1__6343_, data_stage_1__6342_, data_stage_1__6341_, data_stage_1__6340_, data_stage_1__6339_, data_stage_1__6338_, data_stage_1__6337_, data_stage_1__6336_, data_stage_1__6335_, data_stage_1__6334_, data_stage_1__6333_, data_stage_1__6332_, data_stage_1__6331_, data_stage_1__6330_, data_stage_1__6329_, data_stage_1__6328_, data_stage_1__6327_, data_stage_1__6326_, data_stage_1__6325_, data_stage_1__6324_, data_stage_1__6323_, data_stage_1__6322_, data_stage_1__6321_, data_stage_1__6320_, data_stage_1__6319_, data_stage_1__6318_, data_stage_1__6317_, data_stage_1__6316_, data_stage_1__6315_, data_stage_1__6314_, data_stage_1__6313_, data_stage_1__6312_, data_stage_1__6311_, data_stage_1__6310_, data_stage_1__6309_, data_stage_1__6308_, data_stage_1__6307_, data_stage_1__6306_, data_stage_1__6305_, data_stage_1__6304_, data_stage_1__6303_, data_stage_1__6302_, data_stage_1__6301_, data_stage_1__6300_, data_stage_1__6299_, data_stage_1__6298_, data_stage_1__6297_, data_stage_1__6296_, data_stage_1__6295_, data_stage_1__6294_, data_stage_1__6293_, data_stage_1__6292_, data_stage_1__6291_, data_stage_1__6290_, data_stage_1__6289_, data_stage_1__6288_, data_stage_1__6287_, data_stage_1__6286_, data_stage_1__6285_, data_stage_1__6284_, data_stage_1__6283_, data_stage_1__6282_, data_stage_1__6281_, data_stage_1__6280_, data_stage_1__6279_, data_stage_1__6278_, data_stage_1__6277_, data_stage_1__6276_, data_stage_1__6275_, data_stage_1__6274_, data_stage_1__6273_, data_stage_1__6272_, data_stage_1__6271_, data_stage_1__6270_, data_stage_1__6269_, data_stage_1__6268_, data_stage_1__6267_, data_stage_1__6266_, data_stage_1__6265_, data_stage_1__6264_, data_stage_1__6263_, data_stage_1__6262_, data_stage_1__6261_, data_stage_1__6260_, data_stage_1__6259_, data_stage_1__6258_, data_stage_1__6257_, data_stage_1__6256_, data_stage_1__6255_, data_stage_1__6254_, data_stage_1__6253_, data_stage_1__6252_, data_stage_1__6251_, data_stage_1__6250_, data_stage_1__6249_, data_stage_1__6248_, data_stage_1__6247_, data_stage_1__6246_, data_stage_1__6245_, data_stage_1__6244_, data_stage_1__6243_, data_stage_1__6242_, data_stage_1__6241_, data_stage_1__6240_, data_stage_1__6239_, data_stage_1__6238_, data_stage_1__6237_, data_stage_1__6236_, data_stage_1__6235_, data_stage_1__6234_, data_stage_1__6233_, data_stage_1__6232_, data_stage_1__6231_, data_stage_1__6230_, data_stage_1__6229_, data_stage_1__6228_, data_stage_1__6227_, data_stage_1__6226_, data_stage_1__6225_, data_stage_1__6224_, data_stage_1__6223_, data_stage_1__6222_, data_stage_1__6221_, data_stage_1__6220_, data_stage_1__6219_, data_stage_1__6218_, data_stage_1__6217_, data_stage_1__6216_, data_stage_1__6215_, data_stage_1__6214_, data_stage_1__6213_, data_stage_1__6212_, data_stage_1__6211_, data_stage_1__6210_, data_stage_1__6209_, data_stage_1__6208_, data_stage_1__6207_, data_stage_1__6206_, data_stage_1__6205_, data_stage_1__6204_, data_stage_1__6203_, data_stage_1__6202_, data_stage_1__6201_, data_stage_1__6200_, data_stage_1__6199_, data_stage_1__6198_, data_stage_1__6197_, data_stage_1__6196_, data_stage_1__6195_, data_stage_1__6194_, data_stage_1__6193_, data_stage_1__6192_, data_stage_1__6191_, data_stage_1__6190_, data_stage_1__6189_, data_stage_1__6188_, data_stage_1__6187_, data_stage_1__6186_, data_stage_1__6185_, data_stage_1__6184_, data_stage_1__6183_, data_stage_1__6182_, data_stage_1__6181_, data_stage_1__6180_, data_stage_1__6179_, data_stage_1__6178_, data_stage_1__6177_, data_stage_1__6176_, data_stage_1__6175_, data_stage_1__6174_, data_stage_1__6173_, data_stage_1__6172_, data_stage_1__6171_, data_stage_1__6170_, data_stage_1__6169_, data_stage_1__6168_, data_stage_1__6167_, data_stage_1__6166_, data_stage_1__6165_, data_stage_1__6164_, data_stage_1__6163_, data_stage_1__6162_, data_stage_1__6161_, data_stage_1__6160_, data_stage_1__6159_, data_stage_1__6158_, data_stage_1__6157_, data_stage_1__6156_, data_stage_1__6155_, data_stage_1__6154_, data_stage_1__6153_, data_stage_1__6152_, data_stage_1__6151_, data_stage_1__6150_, data_stage_1__6149_, data_stage_1__6148_, data_stage_1__6147_, data_stage_1__6146_, data_stage_1__6145_, data_stage_1__6144_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__6655_, data_stage_2__6654_, data_stage_2__6653_, data_stage_2__6652_, data_stage_2__6651_, data_stage_2__6650_, data_stage_2__6649_, data_stage_2__6648_, data_stage_2__6647_, data_stage_2__6646_, data_stage_2__6645_, data_stage_2__6644_, data_stage_2__6643_, data_stage_2__6642_, data_stage_2__6641_, data_stage_2__6640_, data_stage_2__6639_, data_stage_2__6638_, data_stage_2__6637_, data_stage_2__6636_, data_stage_2__6635_, data_stage_2__6634_, data_stage_2__6633_, data_stage_2__6632_, data_stage_2__6631_, data_stage_2__6630_, data_stage_2__6629_, data_stage_2__6628_, data_stage_2__6627_, data_stage_2__6626_, data_stage_2__6625_, data_stage_2__6624_, data_stage_2__6623_, data_stage_2__6622_, data_stage_2__6621_, data_stage_2__6620_, data_stage_2__6619_, data_stage_2__6618_, data_stage_2__6617_, data_stage_2__6616_, data_stage_2__6615_, data_stage_2__6614_, data_stage_2__6613_, data_stage_2__6612_, data_stage_2__6611_, data_stage_2__6610_, data_stage_2__6609_, data_stage_2__6608_, data_stage_2__6607_, data_stage_2__6606_, data_stage_2__6605_, data_stage_2__6604_, data_stage_2__6603_, data_stage_2__6602_, data_stage_2__6601_, data_stage_2__6600_, data_stage_2__6599_, data_stage_2__6598_, data_stage_2__6597_, data_stage_2__6596_, data_stage_2__6595_, data_stage_2__6594_, data_stage_2__6593_, data_stage_2__6592_, data_stage_2__6591_, data_stage_2__6590_, data_stage_2__6589_, data_stage_2__6588_, data_stage_2__6587_, data_stage_2__6586_, data_stage_2__6585_, data_stage_2__6584_, data_stage_2__6583_, data_stage_2__6582_, data_stage_2__6581_, data_stage_2__6580_, data_stage_2__6579_, data_stage_2__6578_, data_stage_2__6577_, data_stage_2__6576_, data_stage_2__6575_, data_stage_2__6574_, data_stage_2__6573_, data_stage_2__6572_, data_stage_2__6571_, data_stage_2__6570_, data_stage_2__6569_, data_stage_2__6568_, data_stage_2__6567_, data_stage_2__6566_, data_stage_2__6565_, data_stage_2__6564_, data_stage_2__6563_, data_stage_2__6562_, data_stage_2__6561_, data_stage_2__6560_, data_stage_2__6559_, data_stage_2__6558_, data_stage_2__6557_, data_stage_2__6556_, data_stage_2__6555_, data_stage_2__6554_, data_stage_2__6553_, data_stage_2__6552_, data_stage_2__6551_, data_stage_2__6550_, data_stage_2__6549_, data_stage_2__6548_, data_stage_2__6547_, data_stage_2__6546_, data_stage_2__6545_, data_stage_2__6544_, data_stage_2__6543_, data_stage_2__6542_, data_stage_2__6541_, data_stage_2__6540_, data_stage_2__6539_, data_stage_2__6538_, data_stage_2__6537_, data_stage_2__6536_, data_stage_2__6535_, data_stage_2__6534_, data_stage_2__6533_, data_stage_2__6532_, data_stage_2__6531_, data_stage_2__6530_, data_stage_2__6529_, data_stage_2__6528_, data_stage_2__6527_, data_stage_2__6526_, data_stage_2__6525_, data_stage_2__6524_, data_stage_2__6523_, data_stage_2__6522_, data_stage_2__6521_, data_stage_2__6520_, data_stage_2__6519_, data_stage_2__6518_, data_stage_2__6517_, data_stage_2__6516_, data_stage_2__6515_, data_stage_2__6514_, data_stage_2__6513_, data_stage_2__6512_, data_stage_2__6511_, data_stage_2__6510_, data_stage_2__6509_, data_stage_2__6508_, data_stage_2__6507_, data_stage_2__6506_, data_stage_2__6505_, data_stage_2__6504_, data_stage_2__6503_, data_stage_2__6502_, data_stage_2__6501_, data_stage_2__6500_, data_stage_2__6499_, data_stage_2__6498_, data_stage_2__6497_, data_stage_2__6496_, data_stage_2__6495_, data_stage_2__6494_, data_stage_2__6493_, data_stage_2__6492_, data_stage_2__6491_, data_stage_2__6490_, data_stage_2__6489_, data_stage_2__6488_, data_stage_2__6487_, data_stage_2__6486_, data_stage_2__6485_, data_stage_2__6484_, data_stage_2__6483_, data_stage_2__6482_, data_stage_2__6481_, data_stage_2__6480_, data_stage_2__6479_, data_stage_2__6478_, data_stage_2__6477_, data_stage_2__6476_, data_stage_2__6475_, data_stage_2__6474_, data_stage_2__6473_, data_stage_2__6472_, data_stage_2__6471_, data_stage_2__6470_, data_stage_2__6469_, data_stage_2__6468_, data_stage_2__6467_, data_stage_2__6466_, data_stage_2__6465_, data_stage_2__6464_, data_stage_2__6463_, data_stage_2__6462_, data_stage_2__6461_, data_stage_2__6460_, data_stage_2__6459_, data_stage_2__6458_, data_stage_2__6457_, data_stage_2__6456_, data_stage_2__6455_, data_stage_2__6454_, data_stage_2__6453_, data_stage_2__6452_, data_stage_2__6451_, data_stage_2__6450_, data_stage_2__6449_, data_stage_2__6448_, data_stage_2__6447_, data_stage_2__6446_, data_stage_2__6445_, data_stage_2__6444_, data_stage_2__6443_, data_stage_2__6442_, data_stage_2__6441_, data_stage_2__6440_, data_stage_2__6439_, data_stage_2__6438_, data_stage_2__6437_, data_stage_2__6436_, data_stage_2__6435_, data_stage_2__6434_, data_stage_2__6433_, data_stage_2__6432_, data_stage_2__6431_, data_stage_2__6430_, data_stage_2__6429_, data_stage_2__6428_, data_stage_2__6427_, data_stage_2__6426_, data_stage_2__6425_, data_stage_2__6424_, data_stage_2__6423_, data_stage_2__6422_, data_stage_2__6421_, data_stage_2__6420_, data_stage_2__6419_, data_stage_2__6418_, data_stage_2__6417_, data_stage_2__6416_, data_stage_2__6415_, data_stage_2__6414_, data_stage_2__6413_, data_stage_2__6412_, data_stage_2__6411_, data_stage_2__6410_, data_stage_2__6409_, data_stage_2__6408_, data_stage_2__6407_, data_stage_2__6406_, data_stage_2__6405_, data_stage_2__6404_, data_stage_2__6403_, data_stage_2__6402_, data_stage_2__6401_, data_stage_2__6400_, data_stage_2__6399_, data_stage_2__6398_, data_stage_2__6397_, data_stage_2__6396_, data_stage_2__6395_, data_stage_2__6394_, data_stage_2__6393_, data_stage_2__6392_, data_stage_2__6391_, data_stage_2__6390_, data_stage_2__6389_, data_stage_2__6388_, data_stage_2__6387_, data_stage_2__6386_, data_stage_2__6385_, data_stage_2__6384_, data_stage_2__6383_, data_stage_2__6382_, data_stage_2__6381_, data_stage_2__6380_, data_stage_2__6379_, data_stage_2__6378_, data_stage_2__6377_, data_stage_2__6376_, data_stage_2__6375_, data_stage_2__6374_, data_stage_2__6373_, data_stage_2__6372_, data_stage_2__6371_, data_stage_2__6370_, data_stage_2__6369_, data_stage_2__6368_, data_stage_2__6367_, data_stage_2__6366_, data_stage_2__6365_, data_stage_2__6364_, data_stage_2__6363_, data_stage_2__6362_, data_stage_2__6361_, data_stage_2__6360_, data_stage_2__6359_, data_stage_2__6358_, data_stage_2__6357_, data_stage_2__6356_, data_stage_2__6355_, data_stage_2__6354_, data_stage_2__6353_, data_stage_2__6352_, data_stage_2__6351_, data_stage_2__6350_, data_stage_2__6349_, data_stage_2__6348_, data_stage_2__6347_, data_stage_2__6346_, data_stage_2__6345_, data_stage_2__6344_, data_stage_2__6343_, data_stage_2__6342_, data_stage_2__6341_, data_stage_2__6340_, data_stage_2__6339_, data_stage_2__6338_, data_stage_2__6337_, data_stage_2__6336_, data_stage_2__6335_, data_stage_2__6334_, data_stage_2__6333_, data_stage_2__6332_, data_stage_2__6331_, data_stage_2__6330_, data_stage_2__6329_, data_stage_2__6328_, data_stage_2__6327_, data_stage_2__6326_, data_stage_2__6325_, data_stage_2__6324_, data_stage_2__6323_, data_stage_2__6322_, data_stage_2__6321_, data_stage_2__6320_, data_stage_2__6319_, data_stage_2__6318_, data_stage_2__6317_, data_stage_2__6316_, data_stage_2__6315_, data_stage_2__6314_, data_stage_2__6313_, data_stage_2__6312_, data_stage_2__6311_, data_stage_2__6310_, data_stage_2__6309_, data_stage_2__6308_, data_stage_2__6307_, data_stage_2__6306_, data_stage_2__6305_, data_stage_2__6304_, data_stage_2__6303_, data_stage_2__6302_, data_stage_2__6301_, data_stage_2__6300_, data_stage_2__6299_, data_stage_2__6298_, data_stage_2__6297_, data_stage_2__6296_, data_stage_2__6295_, data_stage_2__6294_, data_stage_2__6293_, data_stage_2__6292_, data_stage_2__6291_, data_stage_2__6290_, data_stage_2__6289_, data_stage_2__6288_, data_stage_2__6287_, data_stage_2__6286_, data_stage_2__6285_, data_stage_2__6284_, data_stage_2__6283_, data_stage_2__6282_, data_stage_2__6281_, data_stage_2__6280_, data_stage_2__6279_, data_stage_2__6278_, data_stage_2__6277_, data_stage_2__6276_, data_stage_2__6275_, data_stage_2__6274_, data_stage_2__6273_, data_stage_2__6272_, data_stage_2__6271_, data_stage_2__6270_, data_stage_2__6269_, data_stage_2__6268_, data_stage_2__6267_, data_stage_2__6266_, data_stage_2__6265_, data_stage_2__6264_, data_stage_2__6263_, data_stage_2__6262_, data_stage_2__6261_, data_stage_2__6260_, data_stage_2__6259_, data_stage_2__6258_, data_stage_2__6257_, data_stage_2__6256_, data_stage_2__6255_, data_stage_2__6254_, data_stage_2__6253_, data_stage_2__6252_, data_stage_2__6251_, data_stage_2__6250_, data_stage_2__6249_, data_stage_2__6248_, data_stage_2__6247_, data_stage_2__6246_, data_stage_2__6245_, data_stage_2__6244_, data_stage_2__6243_, data_stage_2__6242_, data_stage_2__6241_, data_stage_2__6240_, data_stage_2__6239_, data_stage_2__6238_, data_stage_2__6237_, data_stage_2__6236_, data_stage_2__6235_, data_stage_2__6234_, data_stage_2__6233_, data_stage_2__6232_, data_stage_2__6231_, data_stage_2__6230_, data_stage_2__6229_, data_stage_2__6228_, data_stage_2__6227_, data_stage_2__6226_, data_stage_2__6225_, data_stage_2__6224_, data_stage_2__6223_, data_stage_2__6222_, data_stage_2__6221_, data_stage_2__6220_, data_stage_2__6219_, data_stage_2__6218_, data_stage_2__6217_, data_stage_2__6216_, data_stage_2__6215_, data_stage_2__6214_, data_stage_2__6213_, data_stage_2__6212_, data_stage_2__6211_, data_stage_2__6210_, data_stage_2__6209_, data_stage_2__6208_, data_stage_2__6207_, data_stage_2__6206_, data_stage_2__6205_, data_stage_2__6204_, data_stage_2__6203_, data_stage_2__6202_, data_stage_2__6201_, data_stage_2__6200_, data_stage_2__6199_, data_stage_2__6198_, data_stage_2__6197_, data_stage_2__6196_, data_stage_2__6195_, data_stage_2__6194_, data_stage_2__6193_, data_stage_2__6192_, data_stage_2__6191_, data_stage_2__6190_, data_stage_2__6189_, data_stage_2__6188_, data_stage_2__6187_, data_stage_2__6186_, data_stage_2__6185_, data_stage_2__6184_, data_stage_2__6183_, data_stage_2__6182_, data_stage_2__6181_, data_stage_2__6180_, data_stage_2__6179_, data_stage_2__6178_, data_stage_2__6177_, data_stage_2__6176_, data_stage_2__6175_, data_stage_2__6174_, data_stage_2__6173_, data_stage_2__6172_, data_stage_2__6171_, data_stage_2__6170_, data_stage_2__6169_, data_stage_2__6168_, data_stage_2__6167_, data_stage_2__6166_, data_stage_2__6165_, data_stage_2__6164_, data_stage_2__6163_, data_stage_2__6162_, data_stage_2__6161_, data_stage_2__6160_, data_stage_2__6159_, data_stage_2__6158_, data_stage_2__6157_, data_stage_2__6156_, data_stage_2__6155_, data_stage_2__6154_, data_stage_2__6153_, data_stage_2__6152_, data_stage_2__6151_, data_stage_2__6150_, data_stage_2__6149_, data_stage_2__6148_, data_stage_2__6147_, data_stage_2__6146_, data_stage_2__6145_, data_stage_2__6144_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_13__swap_inst
  (
    .data_i({ data_stage_1__7167_, data_stage_1__7166_, data_stage_1__7165_, data_stage_1__7164_, data_stage_1__7163_, data_stage_1__7162_, data_stage_1__7161_, data_stage_1__7160_, data_stage_1__7159_, data_stage_1__7158_, data_stage_1__7157_, data_stage_1__7156_, data_stage_1__7155_, data_stage_1__7154_, data_stage_1__7153_, data_stage_1__7152_, data_stage_1__7151_, data_stage_1__7150_, data_stage_1__7149_, data_stage_1__7148_, data_stage_1__7147_, data_stage_1__7146_, data_stage_1__7145_, data_stage_1__7144_, data_stage_1__7143_, data_stage_1__7142_, data_stage_1__7141_, data_stage_1__7140_, data_stage_1__7139_, data_stage_1__7138_, data_stage_1__7137_, data_stage_1__7136_, data_stage_1__7135_, data_stage_1__7134_, data_stage_1__7133_, data_stage_1__7132_, data_stage_1__7131_, data_stage_1__7130_, data_stage_1__7129_, data_stage_1__7128_, data_stage_1__7127_, data_stage_1__7126_, data_stage_1__7125_, data_stage_1__7124_, data_stage_1__7123_, data_stage_1__7122_, data_stage_1__7121_, data_stage_1__7120_, data_stage_1__7119_, data_stage_1__7118_, data_stage_1__7117_, data_stage_1__7116_, data_stage_1__7115_, data_stage_1__7114_, data_stage_1__7113_, data_stage_1__7112_, data_stage_1__7111_, data_stage_1__7110_, data_stage_1__7109_, data_stage_1__7108_, data_stage_1__7107_, data_stage_1__7106_, data_stage_1__7105_, data_stage_1__7104_, data_stage_1__7103_, data_stage_1__7102_, data_stage_1__7101_, data_stage_1__7100_, data_stage_1__7099_, data_stage_1__7098_, data_stage_1__7097_, data_stage_1__7096_, data_stage_1__7095_, data_stage_1__7094_, data_stage_1__7093_, data_stage_1__7092_, data_stage_1__7091_, data_stage_1__7090_, data_stage_1__7089_, data_stage_1__7088_, data_stage_1__7087_, data_stage_1__7086_, data_stage_1__7085_, data_stage_1__7084_, data_stage_1__7083_, data_stage_1__7082_, data_stage_1__7081_, data_stage_1__7080_, data_stage_1__7079_, data_stage_1__7078_, data_stage_1__7077_, data_stage_1__7076_, data_stage_1__7075_, data_stage_1__7074_, data_stage_1__7073_, data_stage_1__7072_, data_stage_1__7071_, data_stage_1__7070_, data_stage_1__7069_, data_stage_1__7068_, data_stage_1__7067_, data_stage_1__7066_, data_stage_1__7065_, data_stage_1__7064_, data_stage_1__7063_, data_stage_1__7062_, data_stage_1__7061_, data_stage_1__7060_, data_stage_1__7059_, data_stage_1__7058_, data_stage_1__7057_, data_stage_1__7056_, data_stage_1__7055_, data_stage_1__7054_, data_stage_1__7053_, data_stage_1__7052_, data_stage_1__7051_, data_stage_1__7050_, data_stage_1__7049_, data_stage_1__7048_, data_stage_1__7047_, data_stage_1__7046_, data_stage_1__7045_, data_stage_1__7044_, data_stage_1__7043_, data_stage_1__7042_, data_stage_1__7041_, data_stage_1__7040_, data_stage_1__7039_, data_stage_1__7038_, data_stage_1__7037_, data_stage_1__7036_, data_stage_1__7035_, data_stage_1__7034_, data_stage_1__7033_, data_stage_1__7032_, data_stage_1__7031_, data_stage_1__7030_, data_stage_1__7029_, data_stage_1__7028_, data_stage_1__7027_, data_stage_1__7026_, data_stage_1__7025_, data_stage_1__7024_, data_stage_1__7023_, data_stage_1__7022_, data_stage_1__7021_, data_stage_1__7020_, data_stage_1__7019_, data_stage_1__7018_, data_stage_1__7017_, data_stage_1__7016_, data_stage_1__7015_, data_stage_1__7014_, data_stage_1__7013_, data_stage_1__7012_, data_stage_1__7011_, data_stage_1__7010_, data_stage_1__7009_, data_stage_1__7008_, data_stage_1__7007_, data_stage_1__7006_, data_stage_1__7005_, data_stage_1__7004_, data_stage_1__7003_, data_stage_1__7002_, data_stage_1__7001_, data_stage_1__7000_, data_stage_1__6999_, data_stage_1__6998_, data_stage_1__6997_, data_stage_1__6996_, data_stage_1__6995_, data_stage_1__6994_, data_stage_1__6993_, data_stage_1__6992_, data_stage_1__6991_, data_stage_1__6990_, data_stage_1__6989_, data_stage_1__6988_, data_stage_1__6987_, data_stage_1__6986_, data_stage_1__6985_, data_stage_1__6984_, data_stage_1__6983_, data_stage_1__6982_, data_stage_1__6981_, data_stage_1__6980_, data_stage_1__6979_, data_stage_1__6978_, data_stage_1__6977_, data_stage_1__6976_, data_stage_1__6975_, data_stage_1__6974_, data_stage_1__6973_, data_stage_1__6972_, data_stage_1__6971_, data_stage_1__6970_, data_stage_1__6969_, data_stage_1__6968_, data_stage_1__6967_, data_stage_1__6966_, data_stage_1__6965_, data_stage_1__6964_, data_stage_1__6963_, data_stage_1__6962_, data_stage_1__6961_, data_stage_1__6960_, data_stage_1__6959_, data_stage_1__6958_, data_stage_1__6957_, data_stage_1__6956_, data_stage_1__6955_, data_stage_1__6954_, data_stage_1__6953_, data_stage_1__6952_, data_stage_1__6951_, data_stage_1__6950_, data_stage_1__6949_, data_stage_1__6948_, data_stage_1__6947_, data_stage_1__6946_, data_stage_1__6945_, data_stage_1__6944_, data_stage_1__6943_, data_stage_1__6942_, data_stage_1__6941_, data_stage_1__6940_, data_stage_1__6939_, data_stage_1__6938_, data_stage_1__6937_, data_stage_1__6936_, data_stage_1__6935_, data_stage_1__6934_, data_stage_1__6933_, data_stage_1__6932_, data_stage_1__6931_, data_stage_1__6930_, data_stage_1__6929_, data_stage_1__6928_, data_stage_1__6927_, data_stage_1__6926_, data_stage_1__6925_, data_stage_1__6924_, data_stage_1__6923_, data_stage_1__6922_, data_stage_1__6921_, data_stage_1__6920_, data_stage_1__6919_, data_stage_1__6918_, data_stage_1__6917_, data_stage_1__6916_, data_stage_1__6915_, data_stage_1__6914_, data_stage_1__6913_, data_stage_1__6912_, data_stage_1__6911_, data_stage_1__6910_, data_stage_1__6909_, data_stage_1__6908_, data_stage_1__6907_, data_stage_1__6906_, data_stage_1__6905_, data_stage_1__6904_, data_stage_1__6903_, data_stage_1__6902_, data_stage_1__6901_, data_stage_1__6900_, data_stage_1__6899_, data_stage_1__6898_, data_stage_1__6897_, data_stage_1__6896_, data_stage_1__6895_, data_stage_1__6894_, data_stage_1__6893_, data_stage_1__6892_, data_stage_1__6891_, data_stage_1__6890_, data_stage_1__6889_, data_stage_1__6888_, data_stage_1__6887_, data_stage_1__6886_, data_stage_1__6885_, data_stage_1__6884_, data_stage_1__6883_, data_stage_1__6882_, data_stage_1__6881_, data_stage_1__6880_, data_stage_1__6879_, data_stage_1__6878_, data_stage_1__6877_, data_stage_1__6876_, data_stage_1__6875_, data_stage_1__6874_, data_stage_1__6873_, data_stage_1__6872_, data_stage_1__6871_, data_stage_1__6870_, data_stage_1__6869_, data_stage_1__6868_, data_stage_1__6867_, data_stage_1__6866_, data_stage_1__6865_, data_stage_1__6864_, data_stage_1__6863_, data_stage_1__6862_, data_stage_1__6861_, data_stage_1__6860_, data_stage_1__6859_, data_stage_1__6858_, data_stage_1__6857_, data_stage_1__6856_, data_stage_1__6855_, data_stage_1__6854_, data_stage_1__6853_, data_stage_1__6852_, data_stage_1__6851_, data_stage_1__6850_, data_stage_1__6849_, data_stage_1__6848_, data_stage_1__6847_, data_stage_1__6846_, data_stage_1__6845_, data_stage_1__6844_, data_stage_1__6843_, data_stage_1__6842_, data_stage_1__6841_, data_stage_1__6840_, data_stage_1__6839_, data_stage_1__6838_, data_stage_1__6837_, data_stage_1__6836_, data_stage_1__6835_, data_stage_1__6834_, data_stage_1__6833_, data_stage_1__6832_, data_stage_1__6831_, data_stage_1__6830_, data_stage_1__6829_, data_stage_1__6828_, data_stage_1__6827_, data_stage_1__6826_, data_stage_1__6825_, data_stage_1__6824_, data_stage_1__6823_, data_stage_1__6822_, data_stage_1__6821_, data_stage_1__6820_, data_stage_1__6819_, data_stage_1__6818_, data_stage_1__6817_, data_stage_1__6816_, data_stage_1__6815_, data_stage_1__6814_, data_stage_1__6813_, data_stage_1__6812_, data_stage_1__6811_, data_stage_1__6810_, data_stage_1__6809_, data_stage_1__6808_, data_stage_1__6807_, data_stage_1__6806_, data_stage_1__6805_, data_stage_1__6804_, data_stage_1__6803_, data_stage_1__6802_, data_stage_1__6801_, data_stage_1__6800_, data_stage_1__6799_, data_stage_1__6798_, data_stage_1__6797_, data_stage_1__6796_, data_stage_1__6795_, data_stage_1__6794_, data_stage_1__6793_, data_stage_1__6792_, data_stage_1__6791_, data_stage_1__6790_, data_stage_1__6789_, data_stage_1__6788_, data_stage_1__6787_, data_stage_1__6786_, data_stage_1__6785_, data_stage_1__6784_, data_stage_1__6783_, data_stage_1__6782_, data_stage_1__6781_, data_stage_1__6780_, data_stage_1__6779_, data_stage_1__6778_, data_stage_1__6777_, data_stage_1__6776_, data_stage_1__6775_, data_stage_1__6774_, data_stage_1__6773_, data_stage_1__6772_, data_stage_1__6771_, data_stage_1__6770_, data_stage_1__6769_, data_stage_1__6768_, data_stage_1__6767_, data_stage_1__6766_, data_stage_1__6765_, data_stage_1__6764_, data_stage_1__6763_, data_stage_1__6762_, data_stage_1__6761_, data_stage_1__6760_, data_stage_1__6759_, data_stage_1__6758_, data_stage_1__6757_, data_stage_1__6756_, data_stage_1__6755_, data_stage_1__6754_, data_stage_1__6753_, data_stage_1__6752_, data_stage_1__6751_, data_stage_1__6750_, data_stage_1__6749_, data_stage_1__6748_, data_stage_1__6747_, data_stage_1__6746_, data_stage_1__6745_, data_stage_1__6744_, data_stage_1__6743_, data_stage_1__6742_, data_stage_1__6741_, data_stage_1__6740_, data_stage_1__6739_, data_stage_1__6738_, data_stage_1__6737_, data_stage_1__6736_, data_stage_1__6735_, data_stage_1__6734_, data_stage_1__6733_, data_stage_1__6732_, data_stage_1__6731_, data_stage_1__6730_, data_stage_1__6729_, data_stage_1__6728_, data_stage_1__6727_, data_stage_1__6726_, data_stage_1__6725_, data_stage_1__6724_, data_stage_1__6723_, data_stage_1__6722_, data_stage_1__6721_, data_stage_1__6720_, data_stage_1__6719_, data_stage_1__6718_, data_stage_1__6717_, data_stage_1__6716_, data_stage_1__6715_, data_stage_1__6714_, data_stage_1__6713_, data_stage_1__6712_, data_stage_1__6711_, data_stage_1__6710_, data_stage_1__6709_, data_stage_1__6708_, data_stage_1__6707_, data_stage_1__6706_, data_stage_1__6705_, data_stage_1__6704_, data_stage_1__6703_, data_stage_1__6702_, data_stage_1__6701_, data_stage_1__6700_, data_stage_1__6699_, data_stage_1__6698_, data_stage_1__6697_, data_stage_1__6696_, data_stage_1__6695_, data_stage_1__6694_, data_stage_1__6693_, data_stage_1__6692_, data_stage_1__6691_, data_stage_1__6690_, data_stage_1__6689_, data_stage_1__6688_, data_stage_1__6687_, data_stage_1__6686_, data_stage_1__6685_, data_stage_1__6684_, data_stage_1__6683_, data_stage_1__6682_, data_stage_1__6681_, data_stage_1__6680_, data_stage_1__6679_, data_stage_1__6678_, data_stage_1__6677_, data_stage_1__6676_, data_stage_1__6675_, data_stage_1__6674_, data_stage_1__6673_, data_stage_1__6672_, data_stage_1__6671_, data_stage_1__6670_, data_stage_1__6669_, data_stage_1__6668_, data_stage_1__6667_, data_stage_1__6666_, data_stage_1__6665_, data_stage_1__6664_, data_stage_1__6663_, data_stage_1__6662_, data_stage_1__6661_, data_stage_1__6660_, data_stage_1__6659_, data_stage_1__6658_, data_stage_1__6657_, data_stage_1__6656_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__7167_, data_stage_2__7166_, data_stage_2__7165_, data_stage_2__7164_, data_stage_2__7163_, data_stage_2__7162_, data_stage_2__7161_, data_stage_2__7160_, data_stage_2__7159_, data_stage_2__7158_, data_stage_2__7157_, data_stage_2__7156_, data_stage_2__7155_, data_stage_2__7154_, data_stage_2__7153_, data_stage_2__7152_, data_stage_2__7151_, data_stage_2__7150_, data_stage_2__7149_, data_stage_2__7148_, data_stage_2__7147_, data_stage_2__7146_, data_stage_2__7145_, data_stage_2__7144_, data_stage_2__7143_, data_stage_2__7142_, data_stage_2__7141_, data_stage_2__7140_, data_stage_2__7139_, data_stage_2__7138_, data_stage_2__7137_, data_stage_2__7136_, data_stage_2__7135_, data_stage_2__7134_, data_stage_2__7133_, data_stage_2__7132_, data_stage_2__7131_, data_stage_2__7130_, data_stage_2__7129_, data_stage_2__7128_, data_stage_2__7127_, data_stage_2__7126_, data_stage_2__7125_, data_stage_2__7124_, data_stage_2__7123_, data_stage_2__7122_, data_stage_2__7121_, data_stage_2__7120_, data_stage_2__7119_, data_stage_2__7118_, data_stage_2__7117_, data_stage_2__7116_, data_stage_2__7115_, data_stage_2__7114_, data_stage_2__7113_, data_stage_2__7112_, data_stage_2__7111_, data_stage_2__7110_, data_stage_2__7109_, data_stage_2__7108_, data_stage_2__7107_, data_stage_2__7106_, data_stage_2__7105_, data_stage_2__7104_, data_stage_2__7103_, data_stage_2__7102_, data_stage_2__7101_, data_stage_2__7100_, data_stage_2__7099_, data_stage_2__7098_, data_stage_2__7097_, data_stage_2__7096_, data_stage_2__7095_, data_stage_2__7094_, data_stage_2__7093_, data_stage_2__7092_, data_stage_2__7091_, data_stage_2__7090_, data_stage_2__7089_, data_stage_2__7088_, data_stage_2__7087_, data_stage_2__7086_, data_stage_2__7085_, data_stage_2__7084_, data_stage_2__7083_, data_stage_2__7082_, data_stage_2__7081_, data_stage_2__7080_, data_stage_2__7079_, data_stage_2__7078_, data_stage_2__7077_, data_stage_2__7076_, data_stage_2__7075_, data_stage_2__7074_, data_stage_2__7073_, data_stage_2__7072_, data_stage_2__7071_, data_stage_2__7070_, data_stage_2__7069_, data_stage_2__7068_, data_stage_2__7067_, data_stage_2__7066_, data_stage_2__7065_, data_stage_2__7064_, data_stage_2__7063_, data_stage_2__7062_, data_stage_2__7061_, data_stage_2__7060_, data_stage_2__7059_, data_stage_2__7058_, data_stage_2__7057_, data_stage_2__7056_, data_stage_2__7055_, data_stage_2__7054_, data_stage_2__7053_, data_stage_2__7052_, data_stage_2__7051_, data_stage_2__7050_, data_stage_2__7049_, data_stage_2__7048_, data_stage_2__7047_, data_stage_2__7046_, data_stage_2__7045_, data_stage_2__7044_, data_stage_2__7043_, data_stage_2__7042_, data_stage_2__7041_, data_stage_2__7040_, data_stage_2__7039_, data_stage_2__7038_, data_stage_2__7037_, data_stage_2__7036_, data_stage_2__7035_, data_stage_2__7034_, data_stage_2__7033_, data_stage_2__7032_, data_stage_2__7031_, data_stage_2__7030_, data_stage_2__7029_, data_stage_2__7028_, data_stage_2__7027_, data_stage_2__7026_, data_stage_2__7025_, data_stage_2__7024_, data_stage_2__7023_, data_stage_2__7022_, data_stage_2__7021_, data_stage_2__7020_, data_stage_2__7019_, data_stage_2__7018_, data_stage_2__7017_, data_stage_2__7016_, data_stage_2__7015_, data_stage_2__7014_, data_stage_2__7013_, data_stage_2__7012_, data_stage_2__7011_, data_stage_2__7010_, data_stage_2__7009_, data_stage_2__7008_, data_stage_2__7007_, data_stage_2__7006_, data_stage_2__7005_, data_stage_2__7004_, data_stage_2__7003_, data_stage_2__7002_, data_stage_2__7001_, data_stage_2__7000_, data_stage_2__6999_, data_stage_2__6998_, data_stage_2__6997_, data_stage_2__6996_, data_stage_2__6995_, data_stage_2__6994_, data_stage_2__6993_, data_stage_2__6992_, data_stage_2__6991_, data_stage_2__6990_, data_stage_2__6989_, data_stage_2__6988_, data_stage_2__6987_, data_stage_2__6986_, data_stage_2__6985_, data_stage_2__6984_, data_stage_2__6983_, data_stage_2__6982_, data_stage_2__6981_, data_stage_2__6980_, data_stage_2__6979_, data_stage_2__6978_, data_stage_2__6977_, data_stage_2__6976_, data_stage_2__6975_, data_stage_2__6974_, data_stage_2__6973_, data_stage_2__6972_, data_stage_2__6971_, data_stage_2__6970_, data_stage_2__6969_, data_stage_2__6968_, data_stage_2__6967_, data_stage_2__6966_, data_stage_2__6965_, data_stage_2__6964_, data_stage_2__6963_, data_stage_2__6962_, data_stage_2__6961_, data_stage_2__6960_, data_stage_2__6959_, data_stage_2__6958_, data_stage_2__6957_, data_stage_2__6956_, data_stage_2__6955_, data_stage_2__6954_, data_stage_2__6953_, data_stage_2__6952_, data_stage_2__6951_, data_stage_2__6950_, data_stage_2__6949_, data_stage_2__6948_, data_stage_2__6947_, data_stage_2__6946_, data_stage_2__6945_, data_stage_2__6944_, data_stage_2__6943_, data_stage_2__6942_, data_stage_2__6941_, data_stage_2__6940_, data_stage_2__6939_, data_stage_2__6938_, data_stage_2__6937_, data_stage_2__6936_, data_stage_2__6935_, data_stage_2__6934_, data_stage_2__6933_, data_stage_2__6932_, data_stage_2__6931_, data_stage_2__6930_, data_stage_2__6929_, data_stage_2__6928_, data_stage_2__6927_, data_stage_2__6926_, data_stage_2__6925_, data_stage_2__6924_, data_stage_2__6923_, data_stage_2__6922_, data_stage_2__6921_, data_stage_2__6920_, data_stage_2__6919_, data_stage_2__6918_, data_stage_2__6917_, data_stage_2__6916_, data_stage_2__6915_, data_stage_2__6914_, data_stage_2__6913_, data_stage_2__6912_, data_stage_2__6911_, data_stage_2__6910_, data_stage_2__6909_, data_stage_2__6908_, data_stage_2__6907_, data_stage_2__6906_, data_stage_2__6905_, data_stage_2__6904_, data_stage_2__6903_, data_stage_2__6902_, data_stage_2__6901_, data_stage_2__6900_, data_stage_2__6899_, data_stage_2__6898_, data_stage_2__6897_, data_stage_2__6896_, data_stage_2__6895_, data_stage_2__6894_, data_stage_2__6893_, data_stage_2__6892_, data_stage_2__6891_, data_stage_2__6890_, data_stage_2__6889_, data_stage_2__6888_, data_stage_2__6887_, data_stage_2__6886_, data_stage_2__6885_, data_stage_2__6884_, data_stage_2__6883_, data_stage_2__6882_, data_stage_2__6881_, data_stage_2__6880_, data_stage_2__6879_, data_stage_2__6878_, data_stage_2__6877_, data_stage_2__6876_, data_stage_2__6875_, data_stage_2__6874_, data_stage_2__6873_, data_stage_2__6872_, data_stage_2__6871_, data_stage_2__6870_, data_stage_2__6869_, data_stage_2__6868_, data_stage_2__6867_, data_stage_2__6866_, data_stage_2__6865_, data_stage_2__6864_, data_stage_2__6863_, data_stage_2__6862_, data_stage_2__6861_, data_stage_2__6860_, data_stage_2__6859_, data_stage_2__6858_, data_stage_2__6857_, data_stage_2__6856_, data_stage_2__6855_, data_stage_2__6854_, data_stage_2__6853_, data_stage_2__6852_, data_stage_2__6851_, data_stage_2__6850_, data_stage_2__6849_, data_stage_2__6848_, data_stage_2__6847_, data_stage_2__6846_, data_stage_2__6845_, data_stage_2__6844_, data_stage_2__6843_, data_stage_2__6842_, data_stage_2__6841_, data_stage_2__6840_, data_stage_2__6839_, data_stage_2__6838_, data_stage_2__6837_, data_stage_2__6836_, data_stage_2__6835_, data_stage_2__6834_, data_stage_2__6833_, data_stage_2__6832_, data_stage_2__6831_, data_stage_2__6830_, data_stage_2__6829_, data_stage_2__6828_, data_stage_2__6827_, data_stage_2__6826_, data_stage_2__6825_, data_stage_2__6824_, data_stage_2__6823_, data_stage_2__6822_, data_stage_2__6821_, data_stage_2__6820_, data_stage_2__6819_, data_stage_2__6818_, data_stage_2__6817_, data_stage_2__6816_, data_stage_2__6815_, data_stage_2__6814_, data_stage_2__6813_, data_stage_2__6812_, data_stage_2__6811_, data_stage_2__6810_, data_stage_2__6809_, data_stage_2__6808_, data_stage_2__6807_, data_stage_2__6806_, data_stage_2__6805_, data_stage_2__6804_, data_stage_2__6803_, data_stage_2__6802_, data_stage_2__6801_, data_stage_2__6800_, data_stage_2__6799_, data_stage_2__6798_, data_stage_2__6797_, data_stage_2__6796_, data_stage_2__6795_, data_stage_2__6794_, data_stage_2__6793_, data_stage_2__6792_, data_stage_2__6791_, data_stage_2__6790_, data_stage_2__6789_, data_stage_2__6788_, data_stage_2__6787_, data_stage_2__6786_, data_stage_2__6785_, data_stage_2__6784_, data_stage_2__6783_, data_stage_2__6782_, data_stage_2__6781_, data_stage_2__6780_, data_stage_2__6779_, data_stage_2__6778_, data_stage_2__6777_, data_stage_2__6776_, data_stage_2__6775_, data_stage_2__6774_, data_stage_2__6773_, data_stage_2__6772_, data_stage_2__6771_, data_stage_2__6770_, data_stage_2__6769_, data_stage_2__6768_, data_stage_2__6767_, data_stage_2__6766_, data_stage_2__6765_, data_stage_2__6764_, data_stage_2__6763_, data_stage_2__6762_, data_stage_2__6761_, data_stage_2__6760_, data_stage_2__6759_, data_stage_2__6758_, data_stage_2__6757_, data_stage_2__6756_, data_stage_2__6755_, data_stage_2__6754_, data_stage_2__6753_, data_stage_2__6752_, data_stage_2__6751_, data_stage_2__6750_, data_stage_2__6749_, data_stage_2__6748_, data_stage_2__6747_, data_stage_2__6746_, data_stage_2__6745_, data_stage_2__6744_, data_stage_2__6743_, data_stage_2__6742_, data_stage_2__6741_, data_stage_2__6740_, data_stage_2__6739_, data_stage_2__6738_, data_stage_2__6737_, data_stage_2__6736_, data_stage_2__6735_, data_stage_2__6734_, data_stage_2__6733_, data_stage_2__6732_, data_stage_2__6731_, data_stage_2__6730_, data_stage_2__6729_, data_stage_2__6728_, data_stage_2__6727_, data_stage_2__6726_, data_stage_2__6725_, data_stage_2__6724_, data_stage_2__6723_, data_stage_2__6722_, data_stage_2__6721_, data_stage_2__6720_, data_stage_2__6719_, data_stage_2__6718_, data_stage_2__6717_, data_stage_2__6716_, data_stage_2__6715_, data_stage_2__6714_, data_stage_2__6713_, data_stage_2__6712_, data_stage_2__6711_, data_stage_2__6710_, data_stage_2__6709_, data_stage_2__6708_, data_stage_2__6707_, data_stage_2__6706_, data_stage_2__6705_, data_stage_2__6704_, data_stage_2__6703_, data_stage_2__6702_, data_stage_2__6701_, data_stage_2__6700_, data_stage_2__6699_, data_stage_2__6698_, data_stage_2__6697_, data_stage_2__6696_, data_stage_2__6695_, data_stage_2__6694_, data_stage_2__6693_, data_stage_2__6692_, data_stage_2__6691_, data_stage_2__6690_, data_stage_2__6689_, data_stage_2__6688_, data_stage_2__6687_, data_stage_2__6686_, data_stage_2__6685_, data_stage_2__6684_, data_stage_2__6683_, data_stage_2__6682_, data_stage_2__6681_, data_stage_2__6680_, data_stage_2__6679_, data_stage_2__6678_, data_stage_2__6677_, data_stage_2__6676_, data_stage_2__6675_, data_stage_2__6674_, data_stage_2__6673_, data_stage_2__6672_, data_stage_2__6671_, data_stage_2__6670_, data_stage_2__6669_, data_stage_2__6668_, data_stage_2__6667_, data_stage_2__6666_, data_stage_2__6665_, data_stage_2__6664_, data_stage_2__6663_, data_stage_2__6662_, data_stage_2__6661_, data_stage_2__6660_, data_stage_2__6659_, data_stage_2__6658_, data_stage_2__6657_, data_stage_2__6656_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_14__swap_inst
  (
    .data_i({ data_stage_1__7679_, data_stage_1__7678_, data_stage_1__7677_, data_stage_1__7676_, data_stage_1__7675_, data_stage_1__7674_, data_stage_1__7673_, data_stage_1__7672_, data_stage_1__7671_, data_stage_1__7670_, data_stage_1__7669_, data_stage_1__7668_, data_stage_1__7667_, data_stage_1__7666_, data_stage_1__7665_, data_stage_1__7664_, data_stage_1__7663_, data_stage_1__7662_, data_stage_1__7661_, data_stage_1__7660_, data_stage_1__7659_, data_stage_1__7658_, data_stage_1__7657_, data_stage_1__7656_, data_stage_1__7655_, data_stage_1__7654_, data_stage_1__7653_, data_stage_1__7652_, data_stage_1__7651_, data_stage_1__7650_, data_stage_1__7649_, data_stage_1__7648_, data_stage_1__7647_, data_stage_1__7646_, data_stage_1__7645_, data_stage_1__7644_, data_stage_1__7643_, data_stage_1__7642_, data_stage_1__7641_, data_stage_1__7640_, data_stage_1__7639_, data_stage_1__7638_, data_stage_1__7637_, data_stage_1__7636_, data_stage_1__7635_, data_stage_1__7634_, data_stage_1__7633_, data_stage_1__7632_, data_stage_1__7631_, data_stage_1__7630_, data_stage_1__7629_, data_stage_1__7628_, data_stage_1__7627_, data_stage_1__7626_, data_stage_1__7625_, data_stage_1__7624_, data_stage_1__7623_, data_stage_1__7622_, data_stage_1__7621_, data_stage_1__7620_, data_stage_1__7619_, data_stage_1__7618_, data_stage_1__7617_, data_stage_1__7616_, data_stage_1__7615_, data_stage_1__7614_, data_stage_1__7613_, data_stage_1__7612_, data_stage_1__7611_, data_stage_1__7610_, data_stage_1__7609_, data_stage_1__7608_, data_stage_1__7607_, data_stage_1__7606_, data_stage_1__7605_, data_stage_1__7604_, data_stage_1__7603_, data_stage_1__7602_, data_stage_1__7601_, data_stage_1__7600_, data_stage_1__7599_, data_stage_1__7598_, data_stage_1__7597_, data_stage_1__7596_, data_stage_1__7595_, data_stage_1__7594_, data_stage_1__7593_, data_stage_1__7592_, data_stage_1__7591_, data_stage_1__7590_, data_stage_1__7589_, data_stage_1__7588_, data_stage_1__7587_, data_stage_1__7586_, data_stage_1__7585_, data_stage_1__7584_, data_stage_1__7583_, data_stage_1__7582_, data_stage_1__7581_, data_stage_1__7580_, data_stage_1__7579_, data_stage_1__7578_, data_stage_1__7577_, data_stage_1__7576_, data_stage_1__7575_, data_stage_1__7574_, data_stage_1__7573_, data_stage_1__7572_, data_stage_1__7571_, data_stage_1__7570_, data_stage_1__7569_, data_stage_1__7568_, data_stage_1__7567_, data_stage_1__7566_, data_stage_1__7565_, data_stage_1__7564_, data_stage_1__7563_, data_stage_1__7562_, data_stage_1__7561_, data_stage_1__7560_, data_stage_1__7559_, data_stage_1__7558_, data_stage_1__7557_, data_stage_1__7556_, data_stage_1__7555_, data_stage_1__7554_, data_stage_1__7553_, data_stage_1__7552_, data_stage_1__7551_, data_stage_1__7550_, data_stage_1__7549_, data_stage_1__7548_, data_stage_1__7547_, data_stage_1__7546_, data_stage_1__7545_, data_stage_1__7544_, data_stage_1__7543_, data_stage_1__7542_, data_stage_1__7541_, data_stage_1__7540_, data_stage_1__7539_, data_stage_1__7538_, data_stage_1__7537_, data_stage_1__7536_, data_stage_1__7535_, data_stage_1__7534_, data_stage_1__7533_, data_stage_1__7532_, data_stage_1__7531_, data_stage_1__7530_, data_stage_1__7529_, data_stage_1__7528_, data_stage_1__7527_, data_stage_1__7526_, data_stage_1__7525_, data_stage_1__7524_, data_stage_1__7523_, data_stage_1__7522_, data_stage_1__7521_, data_stage_1__7520_, data_stage_1__7519_, data_stage_1__7518_, data_stage_1__7517_, data_stage_1__7516_, data_stage_1__7515_, data_stage_1__7514_, data_stage_1__7513_, data_stage_1__7512_, data_stage_1__7511_, data_stage_1__7510_, data_stage_1__7509_, data_stage_1__7508_, data_stage_1__7507_, data_stage_1__7506_, data_stage_1__7505_, data_stage_1__7504_, data_stage_1__7503_, data_stage_1__7502_, data_stage_1__7501_, data_stage_1__7500_, data_stage_1__7499_, data_stage_1__7498_, data_stage_1__7497_, data_stage_1__7496_, data_stage_1__7495_, data_stage_1__7494_, data_stage_1__7493_, data_stage_1__7492_, data_stage_1__7491_, data_stage_1__7490_, data_stage_1__7489_, data_stage_1__7488_, data_stage_1__7487_, data_stage_1__7486_, data_stage_1__7485_, data_stage_1__7484_, data_stage_1__7483_, data_stage_1__7482_, data_stage_1__7481_, data_stage_1__7480_, data_stage_1__7479_, data_stage_1__7478_, data_stage_1__7477_, data_stage_1__7476_, data_stage_1__7475_, data_stage_1__7474_, data_stage_1__7473_, data_stage_1__7472_, data_stage_1__7471_, data_stage_1__7470_, data_stage_1__7469_, data_stage_1__7468_, data_stage_1__7467_, data_stage_1__7466_, data_stage_1__7465_, data_stage_1__7464_, data_stage_1__7463_, data_stage_1__7462_, data_stage_1__7461_, data_stage_1__7460_, data_stage_1__7459_, data_stage_1__7458_, data_stage_1__7457_, data_stage_1__7456_, data_stage_1__7455_, data_stage_1__7454_, data_stage_1__7453_, data_stage_1__7452_, data_stage_1__7451_, data_stage_1__7450_, data_stage_1__7449_, data_stage_1__7448_, data_stage_1__7447_, data_stage_1__7446_, data_stage_1__7445_, data_stage_1__7444_, data_stage_1__7443_, data_stage_1__7442_, data_stage_1__7441_, data_stage_1__7440_, data_stage_1__7439_, data_stage_1__7438_, data_stage_1__7437_, data_stage_1__7436_, data_stage_1__7435_, data_stage_1__7434_, data_stage_1__7433_, data_stage_1__7432_, data_stage_1__7431_, data_stage_1__7430_, data_stage_1__7429_, data_stage_1__7428_, data_stage_1__7427_, data_stage_1__7426_, data_stage_1__7425_, data_stage_1__7424_, data_stage_1__7423_, data_stage_1__7422_, data_stage_1__7421_, data_stage_1__7420_, data_stage_1__7419_, data_stage_1__7418_, data_stage_1__7417_, data_stage_1__7416_, data_stage_1__7415_, data_stage_1__7414_, data_stage_1__7413_, data_stage_1__7412_, data_stage_1__7411_, data_stage_1__7410_, data_stage_1__7409_, data_stage_1__7408_, data_stage_1__7407_, data_stage_1__7406_, data_stage_1__7405_, data_stage_1__7404_, data_stage_1__7403_, data_stage_1__7402_, data_stage_1__7401_, data_stage_1__7400_, data_stage_1__7399_, data_stage_1__7398_, data_stage_1__7397_, data_stage_1__7396_, data_stage_1__7395_, data_stage_1__7394_, data_stage_1__7393_, data_stage_1__7392_, data_stage_1__7391_, data_stage_1__7390_, data_stage_1__7389_, data_stage_1__7388_, data_stage_1__7387_, data_stage_1__7386_, data_stage_1__7385_, data_stage_1__7384_, data_stage_1__7383_, data_stage_1__7382_, data_stage_1__7381_, data_stage_1__7380_, data_stage_1__7379_, data_stage_1__7378_, data_stage_1__7377_, data_stage_1__7376_, data_stage_1__7375_, data_stage_1__7374_, data_stage_1__7373_, data_stage_1__7372_, data_stage_1__7371_, data_stage_1__7370_, data_stage_1__7369_, data_stage_1__7368_, data_stage_1__7367_, data_stage_1__7366_, data_stage_1__7365_, data_stage_1__7364_, data_stage_1__7363_, data_stage_1__7362_, data_stage_1__7361_, data_stage_1__7360_, data_stage_1__7359_, data_stage_1__7358_, data_stage_1__7357_, data_stage_1__7356_, data_stage_1__7355_, data_stage_1__7354_, data_stage_1__7353_, data_stage_1__7352_, data_stage_1__7351_, data_stage_1__7350_, data_stage_1__7349_, data_stage_1__7348_, data_stage_1__7347_, data_stage_1__7346_, data_stage_1__7345_, data_stage_1__7344_, data_stage_1__7343_, data_stage_1__7342_, data_stage_1__7341_, data_stage_1__7340_, data_stage_1__7339_, data_stage_1__7338_, data_stage_1__7337_, data_stage_1__7336_, data_stage_1__7335_, data_stage_1__7334_, data_stage_1__7333_, data_stage_1__7332_, data_stage_1__7331_, data_stage_1__7330_, data_stage_1__7329_, data_stage_1__7328_, data_stage_1__7327_, data_stage_1__7326_, data_stage_1__7325_, data_stage_1__7324_, data_stage_1__7323_, data_stage_1__7322_, data_stage_1__7321_, data_stage_1__7320_, data_stage_1__7319_, data_stage_1__7318_, data_stage_1__7317_, data_stage_1__7316_, data_stage_1__7315_, data_stage_1__7314_, data_stage_1__7313_, data_stage_1__7312_, data_stage_1__7311_, data_stage_1__7310_, data_stage_1__7309_, data_stage_1__7308_, data_stage_1__7307_, data_stage_1__7306_, data_stage_1__7305_, data_stage_1__7304_, data_stage_1__7303_, data_stage_1__7302_, data_stage_1__7301_, data_stage_1__7300_, data_stage_1__7299_, data_stage_1__7298_, data_stage_1__7297_, data_stage_1__7296_, data_stage_1__7295_, data_stage_1__7294_, data_stage_1__7293_, data_stage_1__7292_, data_stage_1__7291_, data_stage_1__7290_, data_stage_1__7289_, data_stage_1__7288_, data_stage_1__7287_, data_stage_1__7286_, data_stage_1__7285_, data_stage_1__7284_, data_stage_1__7283_, data_stage_1__7282_, data_stage_1__7281_, data_stage_1__7280_, data_stage_1__7279_, data_stage_1__7278_, data_stage_1__7277_, data_stage_1__7276_, data_stage_1__7275_, data_stage_1__7274_, data_stage_1__7273_, data_stage_1__7272_, data_stage_1__7271_, data_stage_1__7270_, data_stage_1__7269_, data_stage_1__7268_, data_stage_1__7267_, data_stage_1__7266_, data_stage_1__7265_, data_stage_1__7264_, data_stage_1__7263_, data_stage_1__7262_, data_stage_1__7261_, data_stage_1__7260_, data_stage_1__7259_, data_stage_1__7258_, data_stage_1__7257_, data_stage_1__7256_, data_stage_1__7255_, data_stage_1__7254_, data_stage_1__7253_, data_stage_1__7252_, data_stage_1__7251_, data_stage_1__7250_, data_stage_1__7249_, data_stage_1__7248_, data_stage_1__7247_, data_stage_1__7246_, data_stage_1__7245_, data_stage_1__7244_, data_stage_1__7243_, data_stage_1__7242_, data_stage_1__7241_, data_stage_1__7240_, data_stage_1__7239_, data_stage_1__7238_, data_stage_1__7237_, data_stage_1__7236_, data_stage_1__7235_, data_stage_1__7234_, data_stage_1__7233_, data_stage_1__7232_, data_stage_1__7231_, data_stage_1__7230_, data_stage_1__7229_, data_stage_1__7228_, data_stage_1__7227_, data_stage_1__7226_, data_stage_1__7225_, data_stage_1__7224_, data_stage_1__7223_, data_stage_1__7222_, data_stage_1__7221_, data_stage_1__7220_, data_stage_1__7219_, data_stage_1__7218_, data_stage_1__7217_, data_stage_1__7216_, data_stage_1__7215_, data_stage_1__7214_, data_stage_1__7213_, data_stage_1__7212_, data_stage_1__7211_, data_stage_1__7210_, data_stage_1__7209_, data_stage_1__7208_, data_stage_1__7207_, data_stage_1__7206_, data_stage_1__7205_, data_stage_1__7204_, data_stage_1__7203_, data_stage_1__7202_, data_stage_1__7201_, data_stage_1__7200_, data_stage_1__7199_, data_stage_1__7198_, data_stage_1__7197_, data_stage_1__7196_, data_stage_1__7195_, data_stage_1__7194_, data_stage_1__7193_, data_stage_1__7192_, data_stage_1__7191_, data_stage_1__7190_, data_stage_1__7189_, data_stage_1__7188_, data_stage_1__7187_, data_stage_1__7186_, data_stage_1__7185_, data_stage_1__7184_, data_stage_1__7183_, data_stage_1__7182_, data_stage_1__7181_, data_stage_1__7180_, data_stage_1__7179_, data_stage_1__7178_, data_stage_1__7177_, data_stage_1__7176_, data_stage_1__7175_, data_stage_1__7174_, data_stage_1__7173_, data_stage_1__7172_, data_stage_1__7171_, data_stage_1__7170_, data_stage_1__7169_, data_stage_1__7168_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__7679_, data_stage_2__7678_, data_stage_2__7677_, data_stage_2__7676_, data_stage_2__7675_, data_stage_2__7674_, data_stage_2__7673_, data_stage_2__7672_, data_stage_2__7671_, data_stage_2__7670_, data_stage_2__7669_, data_stage_2__7668_, data_stage_2__7667_, data_stage_2__7666_, data_stage_2__7665_, data_stage_2__7664_, data_stage_2__7663_, data_stage_2__7662_, data_stage_2__7661_, data_stage_2__7660_, data_stage_2__7659_, data_stage_2__7658_, data_stage_2__7657_, data_stage_2__7656_, data_stage_2__7655_, data_stage_2__7654_, data_stage_2__7653_, data_stage_2__7652_, data_stage_2__7651_, data_stage_2__7650_, data_stage_2__7649_, data_stage_2__7648_, data_stage_2__7647_, data_stage_2__7646_, data_stage_2__7645_, data_stage_2__7644_, data_stage_2__7643_, data_stage_2__7642_, data_stage_2__7641_, data_stage_2__7640_, data_stage_2__7639_, data_stage_2__7638_, data_stage_2__7637_, data_stage_2__7636_, data_stage_2__7635_, data_stage_2__7634_, data_stage_2__7633_, data_stage_2__7632_, data_stage_2__7631_, data_stage_2__7630_, data_stage_2__7629_, data_stage_2__7628_, data_stage_2__7627_, data_stage_2__7626_, data_stage_2__7625_, data_stage_2__7624_, data_stage_2__7623_, data_stage_2__7622_, data_stage_2__7621_, data_stage_2__7620_, data_stage_2__7619_, data_stage_2__7618_, data_stage_2__7617_, data_stage_2__7616_, data_stage_2__7615_, data_stage_2__7614_, data_stage_2__7613_, data_stage_2__7612_, data_stage_2__7611_, data_stage_2__7610_, data_stage_2__7609_, data_stage_2__7608_, data_stage_2__7607_, data_stage_2__7606_, data_stage_2__7605_, data_stage_2__7604_, data_stage_2__7603_, data_stage_2__7602_, data_stage_2__7601_, data_stage_2__7600_, data_stage_2__7599_, data_stage_2__7598_, data_stage_2__7597_, data_stage_2__7596_, data_stage_2__7595_, data_stage_2__7594_, data_stage_2__7593_, data_stage_2__7592_, data_stage_2__7591_, data_stage_2__7590_, data_stage_2__7589_, data_stage_2__7588_, data_stage_2__7587_, data_stage_2__7586_, data_stage_2__7585_, data_stage_2__7584_, data_stage_2__7583_, data_stage_2__7582_, data_stage_2__7581_, data_stage_2__7580_, data_stage_2__7579_, data_stage_2__7578_, data_stage_2__7577_, data_stage_2__7576_, data_stage_2__7575_, data_stage_2__7574_, data_stage_2__7573_, data_stage_2__7572_, data_stage_2__7571_, data_stage_2__7570_, data_stage_2__7569_, data_stage_2__7568_, data_stage_2__7567_, data_stage_2__7566_, data_stage_2__7565_, data_stage_2__7564_, data_stage_2__7563_, data_stage_2__7562_, data_stage_2__7561_, data_stage_2__7560_, data_stage_2__7559_, data_stage_2__7558_, data_stage_2__7557_, data_stage_2__7556_, data_stage_2__7555_, data_stage_2__7554_, data_stage_2__7553_, data_stage_2__7552_, data_stage_2__7551_, data_stage_2__7550_, data_stage_2__7549_, data_stage_2__7548_, data_stage_2__7547_, data_stage_2__7546_, data_stage_2__7545_, data_stage_2__7544_, data_stage_2__7543_, data_stage_2__7542_, data_stage_2__7541_, data_stage_2__7540_, data_stage_2__7539_, data_stage_2__7538_, data_stage_2__7537_, data_stage_2__7536_, data_stage_2__7535_, data_stage_2__7534_, data_stage_2__7533_, data_stage_2__7532_, data_stage_2__7531_, data_stage_2__7530_, data_stage_2__7529_, data_stage_2__7528_, data_stage_2__7527_, data_stage_2__7526_, data_stage_2__7525_, data_stage_2__7524_, data_stage_2__7523_, data_stage_2__7522_, data_stage_2__7521_, data_stage_2__7520_, data_stage_2__7519_, data_stage_2__7518_, data_stage_2__7517_, data_stage_2__7516_, data_stage_2__7515_, data_stage_2__7514_, data_stage_2__7513_, data_stage_2__7512_, data_stage_2__7511_, data_stage_2__7510_, data_stage_2__7509_, data_stage_2__7508_, data_stage_2__7507_, data_stage_2__7506_, data_stage_2__7505_, data_stage_2__7504_, data_stage_2__7503_, data_stage_2__7502_, data_stage_2__7501_, data_stage_2__7500_, data_stage_2__7499_, data_stage_2__7498_, data_stage_2__7497_, data_stage_2__7496_, data_stage_2__7495_, data_stage_2__7494_, data_stage_2__7493_, data_stage_2__7492_, data_stage_2__7491_, data_stage_2__7490_, data_stage_2__7489_, data_stage_2__7488_, data_stage_2__7487_, data_stage_2__7486_, data_stage_2__7485_, data_stage_2__7484_, data_stage_2__7483_, data_stage_2__7482_, data_stage_2__7481_, data_stage_2__7480_, data_stage_2__7479_, data_stage_2__7478_, data_stage_2__7477_, data_stage_2__7476_, data_stage_2__7475_, data_stage_2__7474_, data_stage_2__7473_, data_stage_2__7472_, data_stage_2__7471_, data_stage_2__7470_, data_stage_2__7469_, data_stage_2__7468_, data_stage_2__7467_, data_stage_2__7466_, data_stage_2__7465_, data_stage_2__7464_, data_stage_2__7463_, data_stage_2__7462_, data_stage_2__7461_, data_stage_2__7460_, data_stage_2__7459_, data_stage_2__7458_, data_stage_2__7457_, data_stage_2__7456_, data_stage_2__7455_, data_stage_2__7454_, data_stage_2__7453_, data_stage_2__7452_, data_stage_2__7451_, data_stage_2__7450_, data_stage_2__7449_, data_stage_2__7448_, data_stage_2__7447_, data_stage_2__7446_, data_stage_2__7445_, data_stage_2__7444_, data_stage_2__7443_, data_stage_2__7442_, data_stage_2__7441_, data_stage_2__7440_, data_stage_2__7439_, data_stage_2__7438_, data_stage_2__7437_, data_stage_2__7436_, data_stage_2__7435_, data_stage_2__7434_, data_stage_2__7433_, data_stage_2__7432_, data_stage_2__7431_, data_stage_2__7430_, data_stage_2__7429_, data_stage_2__7428_, data_stage_2__7427_, data_stage_2__7426_, data_stage_2__7425_, data_stage_2__7424_, data_stage_2__7423_, data_stage_2__7422_, data_stage_2__7421_, data_stage_2__7420_, data_stage_2__7419_, data_stage_2__7418_, data_stage_2__7417_, data_stage_2__7416_, data_stage_2__7415_, data_stage_2__7414_, data_stage_2__7413_, data_stage_2__7412_, data_stage_2__7411_, data_stage_2__7410_, data_stage_2__7409_, data_stage_2__7408_, data_stage_2__7407_, data_stage_2__7406_, data_stage_2__7405_, data_stage_2__7404_, data_stage_2__7403_, data_stage_2__7402_, data_stage_2__7401_, data_stage_2__7400_, data_stage_2__7399_, data_stage_2__7398_, data_stage_2__7397_, data_stage_2__7396_, data_stage_2__7395_, data_stage_2__7394_, data_stage_2__7393_, data_stage_2__7392_, data_stage_2__7391_, data_stage_2__7390_, data_stage_2__7389_, data_stage_2__7388_, data_stage_2__7387_, data_stage_2__7386_, data_stage_2__7385_, data_stage_2__7384_, data_stage_2__7383_, data_stage_2__7382_, data_stage_2__7381_, data_stage_2__7380_, data_stage_2__7379_, data_stage_2__7378_, data_stage_2__7377_, data_stage_2__7376_, data_stage_2__7375_, data_stage_2__7374_, data_stage_2__7373_, data_stage_2__7372_, data_stage_2__7371_, data_stage_2__7370_, data_stage_2__7369_, data_stage_2__7368_, data_stage_2__7367_, data_stage_2__7366_, data_stage_2__7365_, data_stage_2__7364_, data_stage_2__7363_, data_stage_2__7362_, data_stage_2__7361_, data_stage_2__7360_, data_stage_2__7359_, data_stage_2__7358_, data_stage_2__7357_, data_stage_2__7356_, data_stage_2__7355_, data_stage_2__7354_, data_stage_2__7353_, data_stage_2__7352_, data_stage_2__7351_, data_stage_2__7350_, data_stage_2__7349_, data_stage_2__7348_, data_stage_2__7347_, data_stage_2__7346_, data_stage_2__7345_, data_stage_2__7344_, data_stage_2__7343_, data_stage_2__7342_, data_stage_2__7341_, data_stage_2__7340_, data_stage_2__7339_, data_stage_2__7338_, data_stage_2__7337_, data_stage_2__7336_, data_stage_2__7335_, data_stage_2__7334_, data_stage_2__7333_, data_stage_2__7332_, data_stage_2__7331_, data_stage_2__7330_, data_stage_2__7329_, data_stage_2__7328_, data_stage_2__7327_, data_stage_2__7326_, data_stage_2__7325_, data_stage_2__7324_, data_stage_2__7323_, data_stage_2__7322_, data_stage_2__7321_, data_stage_2__7320_, data_stage_2__7319_, data_stage_2__7318_, data_stage_2__7317_, data_stage_2__7316_, data_stage_2__7315_, data_stage_2__7314_, data_stage_2__7313_, data_stage_2__7312_, data_stage_2__7311_, data_stage_2__7310_, data_stage_2__7309_, data_stage_2__7308_, data_stage_2__7307_, data_stage_2__7306_, data_stage_2__7305_, data_stage_2__7304_, data_stage_2__7303_, data_stage_2__7302_, data_stage_2__7301_, data_stage_2__7300_, data_stage_2__7299_, data_stage_2__7298_, data_stage_2__7297_, data_stage_2__7296_, data_stage_2__7295_, data_stage_2__7294_, data_stage_2__7293_, data_stage_2__7292_, data_stage_2__7291_, data_stage_2__7290_, data_stage_2__7289_, data_stage_2__7288_, data_stage_2__7287_, data_stage_2__7286_, data_stage_2__7285_, data_stage_2__7284_, data_stage_2__7283_, data_stage_2__7282_, data_stage_2__7281_, data_stage_2__7280_, data_stage_2__7279_, data_stage_2__7278_, data_stage_2__7277_, data_stage_2__7276_, data_stage_2__7275_, data_stage_2__7274_, data_stage_2__7273_, data_stage_2__7272_, data_stage_2__7271_, data_stage_2__7270_, data_stage_2__7269_, data_stage_2__7268_, data_stage_2__7267_, data_stage_2__7266_, data_stage_2__7265_, data_stage_2__7264_, data_stage_2__7263_, data_stage_2__7262_, data_stage_2__7261_, data_stage_2__7260_, data_stage_2__7259_, data_stage_2__7258_, data_stage_2__7257_, data_stage_2__7256_, data_stage_2__7255_, data_stage_2__7254_, data_stage_2__7253_, data_stage_2__7252_, data_stage_2__7251_, data_stage_2__7250_, data_stage_2__7249_, data_stage_2__7248_, data_stage_2__7247_, data_stage_2__7246_, data_stage_2__7245_, data_stage_2__7244_, data_stage_2__7243_, data_stage_2__7242_, data_stage_2__7241_, data_stage_2__7240_, data_stage_2__7239_, data_stage_2__7238_, data_stage_2__7237_, data_stage_2__7236_, data_stage_2__7235_, data_stage_2__7234_, data_stage_2__7233_, data_stage_2__7232_, data_stage_2__7231_, data_stage_2__7230_, data_stage_2__7229_, data_stage_2__7228_, data_stage_2__7227_, data_stage_2__7226_, data_stage_2__7225_, data_stage_2__7224_, data_stage_2__7223_, data_stage_2__7222_, data_stage_2__7221_, data_stage_2__7220_, data_stage_2__7219_, data_stage_2__7218_, data_stage_2__7217_, data_stage_2__7216_, data_stage_2__7215_, data_stage_2__7214_, data_stage_2__7213_, data_stage_2__7212_, data_stage_2__7211_, data_stage_2__7210_, data_stage_2__7209_, data_stage_2__7208_, data_stage_2__7207_, data_stage_2__7206_, data_stage_2__7205_, data_stage_2__7204_, data_stage_2__7203_, data_stage_2__7202_, data_stage_2__7201_, data_stage_2__7200_, data_stage_2__7199_, data_stage_2__7198_, data_stage_2__7197_, data_stage_2__7196_, data_stage_2__7195_, data_stage_2__7194_, data_stage_2__7193_, data_stage_2__7192_, data_stage_2__7191_, data_stage_2__7190_, data_stage_2__7189_, data_stage_2__7188_, data_stage_2__7187_, data_stage_2__7186_, data_stage_2__7185_, data_stage_2__7184_, data_stage_2__7183_, data_stage_2__7182_, data_stage_2__7181_, data_stage_2__7180_, data_stage_2__7179_, data_stage_2__7178_, data_stage_2__7177_, data_stage_2__7176_, data_stage_2__7175_, data_stage_2__7174_, data_stage_2__7173_, data_stage_2__7172_, data_stage_2__7171_, data_stage_2__7170_, data_stage_2__7169_, data_stage_2__7168_ })
  );


  bsg_swap_width_p256
  mux_stage_1__mux_swap_15__swap_inst
  (
    .data_i({ data_stage_1__8191_, data_stage_1__8190_, data_stage_1__8189_, data_stage_1__8188_, data_stage_1__8187_, data_stage_1__8186_, data_stage_1__8185_, data_stage_1__8184_, data_stage_1__8183_, data_stage_1__8182_, data_stage_1__8181_, data_stage_1__8180_, data_stage_1__8179_, data_stage_1__8178_, data_stage_1__8177_, data_stage_1__8176_, data_stage_1__8175_, data_stage_1__8174_, data_stage_1__8173_, data_stage_1__8172_, data_stage_1__8171_, data_stage_1__8170_, data_stage_1__8169_, data_stage_1__8168_, data_stage_1__8167_, data_stage_1__8166_, data_stage_1__8165_, data_stage_1__8164_, data_stage_1__8163_, data_stage_1__8162_, data_stage_1__8161_, data_stage_1__8160_, data_stage_1__8159_, data_stage_1__8158_, data_stage_1__8157_, data_stage_1__8156_, data_stage_1__8155_, data_stage_1__8154_, data_stage_1__8153_, data_stage_1__8152_, data_stage_1__8151_, data_stage_1__8150_, data_stage_1__8149_, data_stage_1__8148_, data_stage_1__8147_, data_stage_1__8146_, data_stage_1__8145_, data_stage_1__8144_, data_stage_1__8143_, data_stage_1__8142_, data_stage_1__8141_, data_stage_1__8140_, data_stage_1__8139_, data_stage_1__8138_, data_stage_1__8137_, data_stage_1__8136_, data_stage_1__8135_, data_stage_1__8134_, data_stage_1__8133_, data_stage_1__8132_, data_stage_1__8131_, data_stage_1__8130_, data_stage_1__8129_, data_stage_1__8128_, data_stage_1__8127_, data_stage_1__8126_, data_stage_1__8125_, data_stage_1__8124_, data_stage_1__8123_, data_stage_1__8122_, data_stage_1__8121_, data_stage_1__8120_, data_stage_1__8119_, data_stage_1__8118_, data_stage_1__8117_, data_stage_1__8116_, data_stage_1__8115_, data_stage_1__8114_, data_stage_1__8113_, data_stage_1__8112_, data_stage_1__8111_, data_stage_1__8110_, data_stage_1__8109_, data_stage_1__8108_, data_stage_1__8107_, data_stage_1__8106_, data_stage_1__8105_, data_stage_1__8104_, data_stage_1__8103_, data_stage_1__8102_, data_stage_1__8101_, data_stage_1__8100_, data_stage_1__8099_, data_stage_1__8098_, data_stage_1__8097_, data_stage_1__8096_, data_stage_1__8095_, data_stage_1__8094_, data_stage_1__8093_, data_stage_1__8092_, data_stage_1__8091_, data_stage_1__8090_, data_stage_1__8089_, data_stage_1__8088_, data_stage_1__8087_, data_stage_1__8086_, data_stage_1__8085_, data_stage_1__8084_, data_stage_1__8083_, data_stage_1__8082_, data_stage_1__8081_, data_stage_1__8080_, data_stage_1__8079_, data_stage_1__8078_, data_stage_1__8077_, data_stage_1__8076_, data_stage_1__8075_, data_stage_1__8074_, data_stage_1__8073_, data_stage_1__8072_, data_stage_1__8071_, data_stage_1__8070_, data_stage_1__8069_, data_stage_1__8068_, data_stage_1__8067_, data_stage_1__8066_, data_stage_1__8065_, data_stage_1__8064_, data_stage_1__8063_, data_stage_1__8062_, data_stage_1__8061_, data_stage_1__8060_, data_stage_1__8059_, data_stage_1__8058_, data_stage_1__8057_, data_stage_1__8056_, data_stage_1__8055_, data_stage_1__8054_, data_stage_1__8053_, data_stage_1__8052_, data_stage_1__8051_, data_stage_1__8050_, data_stage_1__8049_, data_stage_1__8048_, data_stage_1__8047_, data_stage_1__8046_, data_stage_1__8045_, data_stage_1__8044_, data_stage_1__8043_, data_stage_1__8042_, data_stage_1__8041_, data_stage_1__8040_, data_stage_1__8039_, data_stage_1__8038_, data_stage_1__8037_, data_stage_1__8036_, data_stage_1__8035_, data_stage_1__8034_, data_stage_1__8033_, data_stage_1__8032_, data_stage_1__8031_, data_stage_1__8030_, data_stage_1__8029_, data_stage_1__8028_, data_stage_1__8027_, data_stage_1__8026_, data_stage_1__8025_, data_stage_1__8024_, data_stage_1__8023_, data_stage_1__8022_, data_stage_1__8021_, data_stage_1__8020_, data_stage_1__8019_, data_stage_1__8018_, data_stage_1__8017_, data_stage_1__8016_, data_stage_1__8015_, data_stage_1__8014_, data_stage_1__8013_, data_stage_1__8012_, data_stage_1__8011_, data_stage_1__8010_, data_stage_1__8009_, data_stage_1__8008_, data_stage_1__8007_, data_stage_1__8006_, data_stage_1__8005_, data_stage_1__8004_, data_stage_1__8003_, data_stage_1__8002_, data_stage_1__8001_, data_stage_1__8000_, data_stage_1__7999_, data_stage_1__7998_, data_stage_1__7997_, data_stage_1__7996_, data_stage_1__7995_, data_stage_1__7994_, data_stage_1__7993_, data_stage_1__7992_, data_stage_1__7991_, data_stage_1__7990_, data_stage_1__7989_, data_stage_1__7988_, data_stage_1__7987_, data_stage_1__7986_, data_stage_1__7985_, data_stage_1__7984_, data_stage_1__7983_, data_stage_1__7982_, data_stage_1__7981_, data_stage_1__7980_, data_stage_1__7979_, data_stage_1__7978_, data_stage_1__7977_, data_stage_1__7976_, data_stage_1__7975_, data_stage_1__7974_, data_stage_1__7973_, data_stage_1__7972_, data_stage_1__7971_, data_stage_1__7970_, data_stage_1__7969_, data_stage_1__7968_, data_stage_1__7967_, data_stage_1__7966_, data_stage_1__7965_, data_stage_1__7964_, data_stage_1__7963_, data_stage_1__7962_, data_stage_1__7961_, data_stage_1__7960_, data_stage_1__7959_, data_stage_1__7958_, data_stage_1__7957_, data_stage_1__7956_, data_stage_1__7955_, data_stage_1__7954_, data_stage_1__7953_, data_stage_1__7952_, data_stage_1__7951_, data_stage_1__7950_, data_stage_1__7949_, data_stage_1__7948_, data_stage_1__7947_, data_stage_1__7946_, data_stage_1__7945_, data_stage_1__7944_, data_stage_1__7943_, data_stage_1__7942_, data_stage_1__7941_, data_stage_1__7940_, data_stage_1__7939_, data_stage_1__7938_, data_stage_1__7937_, data_stage_1__7936_, data_stage_1__7935_, data_stage_1__7934_, data_stage_1__7933_, data_stage_1__7932_, data_stage_1__7931_, data_stage_1__7930_, data_stage_1__7929_, data_stage_1__7928_, data_stage_1__7927_, data_stage_1__7926_, data_stage_1__7925_, data_stage_1__7924_, data_stage_1__7923_, data_stage_1__7922_, data_stage_1__7921_, data_stage_1__7920_, data_stage_1__7919_, data_stage_1__7918_, data_stage_1__7917_, data_stage_1__7916_, data_stage_1__7915_, data_stage_1__7914_, data_stage_1__7913_, data_stage_1__7912_, data_stage_1__7911_, data_stage_1__7910_, data_stage_1__7909_, data_stage_1__7908_, data_stage_1__7907_, data_stage_1__7906_, data_stage_1__7905_, data_stage_1__7904_, data_stage_1__7903_, data_stage_1__7902_, data_stage_1__7901_, data_stage_1__7900_, data_stage_1__7899_, data_stage_1__7898_, data_stage_1__7897_, data_stage_1__7896_, data_stage_1__7895_, data_stage_1__7894_, data_stage_1__7893_, data_stage_1__7892_, data_stage_1__7891_, data_stage_1__7890_, data_stage_1__7889_, data_stage_1__7888_, data_stage_1__7887_, data_stage_1__7886_, data_stage_1__7885_, data_stage_1__7884_, data_stage_1__7883_, data_stage_1__7882_, data_stage_1__7881_, data_stage_1__7880_, data_stage_1__7879_, data_stage_1__7878_, data_stage_1__7877_, data_stage_1__7876_, data_stage_1__7875_, data_stage_1__7874_, data_stage_1__7873_, data_stage_1__7872_, data_stage_1__7871_, data_stage_1__7870_, data_stage_1__7869_, data_stage_1__7868_, data_stage_1__7867_, data_stage_1__7866_, data_stage_1__7865_, data_stage_1__7864_, data_stage_1__7863_, data_stage_1__7862_, data_stage_1__7861_, data_stage_1__7860_, data_stage_1__7859_, data_stage_1__7858_, data_stage_1__7857_, data_stage_1__7856_, data_stage_1__7855_, data_stage_1__7854_, data_stage_1__7853_, data_stage_1__7852_, data_stage_1__7851_, data_stage_1__7850_, data_stage_1__7849_, data_stage_1__7848_, data_stage_1__7847_, data_stage_1__7846_, data_stage_1__7845_, data_stage_1__7844_, data_stage_1__7843_, data_stage_1__7842_, data_stage_1__7841_, data_stage_1__7840_, data_stage_1__7839_, data_stage_1__7838_, data_stage_1__7837_, data_stage_1__7836_, data_stage_1__7835_, data_stage_1__7834_, data_stage_1__7833_, data_stage_1__7832_, data_stage_1__7831_, data_stage_1__7830_, data_stage_1__7829_, data_stage_1__7828_, data_stage_1__7827_, data_stage_1__7826_, data_stage_1__7825_, data_stage_1__7824_, data_stage_1__7823_, data_stage_1__7822_, data_stage_1__7821_, data_stage_1__7820_, data_stage_1__7819_, data_stage_1__7818_, data_stage_1__7817_, data_stage_1__7816_, data_stage_1__7815_, data_stage_1__7814_, data_stage_1__7813_, data_stage_1__7812_, data_stage_1__7811_, data_stage_1__7810_, data_stage_1__7809_, data_stage_1__7808_, data_stage_1__7807_, data_stage_1__7806_, data_stage_1__7805_, data_stage_1__7804_, data_stage_1__7803_, data_stage_1__7802_, data_stage_1__7801_, data_stage_1__7800_, data_stage_1__7799_, data_stage_1__7798_, data_stage_1__7797_, data_stage_1__7796_, data_stage_1__7795_, data_stage_1__7794_, data_stage_1__7793_, data_stage_1__7792_, data_stage_1__7791_, data_stage_1__7790_, data_stage_1__7789_, data_stage_1__7788_, data_stage_1__7787_, data_stage_1__7786_, data_stage_1__7785_, data_stage_1__7784_, data_stage_1__7783_, data_stage_1__7782_, data_stage_1__7781_, data_stage_1__7780_, data_stage_1__7779_, data_stage_1__7778_, data_stage_1__7777_, data_stage_1__7776_, data_stage_1__7775_, data_stage_1__7774_, data_stage_1__7773_, data_stage_1__7772_, data_stage_1__7771_, data_stage_1__7770_, data_stage_1__7769_, data_stage_1__7768_, data_stage_1__7767_, data_stage_1__7766_, data_stage_1__7765_, data_stage_1__7764_, data_stage_1__7763_, data_stage_1__7762_, data_stage_1__7761_, data_stage_1__7760_, data_stage_1__7759_, data_stage_1__7758_, data_stage_1__7757_, data_stage_1__7756_, data_stage_1__7755_, data_stage_1__7754_, data_stage_1__7753_, data_stage_1__7752_, data_stage_1__7751_, data_stage_1__7750_, data_stage_1__7749_, data_stage_1__7748_, data_stage_1__7747_, data_stage_1__7746_, data_stage_1__7745_, data_stage_1__7744_, data_stage_1__7743_, data_stage_1__7742_, data_stage_1__7741_, data_stage_1__7740_, data_stage_1__7739_, data_stage_1__7738_, data_stage_1__7737_, data_stage_1__7736_, data_stage_1__7735_, data_stage_1__7734_, data_stage_1__7733_, data_stage_1__7732_, data_stage_1__7731_, data_stage_1__7730_, data_stage_1__7729_, data_stage_1__7728_, data_stage_1__7727_, data_stage_1__7726_, data_stage_1__7725_, data_stage_1__7724_, data_stage_1__7723_, data_stage_1__7722_, data_stage_1__7721_, data_stage_1__7720_, data_stage_1__7719_, data_stage_1__7718_, data_stage_1__7717_, data_stage_1__7716_, data_stage_1__7715_, data_stage_1__7714_, data_stage_1__7713_, data_stage_1__7712_, data_stage_1__7711_, data_stage_1__7710_, data_stage_1__7709_, data_stage_1__7708_, data_stage_1__7707_, data_stage_1__7706_, data_stage_1__7705_, data_stage_1__7704_, data_stage_1__7703_, data_stage_1__7702_, data_stage_1__7701_, data_stage_1__7700_, data_stage_1__7699_, data_stage_1__7698_, data_stage_1__7697_, data_stage_1__7696_, data_stage_1__7695_, data_stage_1__7694_, data_stage_1__7693_, data_stage_1__7692_, data_stage_1__7691_, data_stage_1__7690_, data_stage_1__7689_, data_stage_1__7688_, data_stage_1__7687_, data_stage_1__7686_, data_stage_1__7685_, data_stage_1__7684_, data_stage_1__7683_, data_stage_1__7682_, data_stage_1__7681_, data_stage_1__7680_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__8191_, data_stage_2__8190_, data_stage_2__8189_, data_stage_2__8188_, data_stage_2__8187_, data_stage_2__8186_, data_stage_2__8185_, data_stage_2__8184_, data_stage_2__8183_, data_stage_2__8182_, data_stage_2__8181_, data_stage_2__8180_, data_stage_2__8179_, data_stage_2__8178_, data_stage_2__8177_, data_stage_2__8176_, data_stage_2__8175_, data_stage_2__8174_, data_stage_2__8173_, data_stage_2__8172_, data_stage_2__8171_, data_stage_2__8170_, data_stage_2__8169_, data_stage_2__8168_, data_stage_2__8167_, data_stage_2__8166_, data_stage_2__8165_, data_stage_2__8164_, data_stage_2__8163_, data_stage_2__8162_, data_stage_2__8161_, data_stage_2__8160_, data_stage_2__8159_, data_stage_2__8158_, data_stage_2__8157_, data_stage_2__8156_, data_stage_2__8155_, data_stage_2__8154_, data_stage_2__8153_, data_stage_2__8152_, data_stage_2__8151_, data_stage_2__8150_, data_stage_2__8149_, data_stage_2__8148_, data_stage_2__8147_, data_stage_2__8146_, data_stage_2__8145_, data_stage_2__8144_, data_stage_2__8143_, data_stage_2__8142_, data_stage_2__8141_, data_stage_2__8140_, data_stage_2__8139_, data_stage_2__8138_, data_stage_2__8137_, data_stage_2__8136_, data_stage_2__8135_, data_stage_2__8134_, data_stage_2__8133_, data_stage_2__8132_, data_stage_2__8131_, data_stage_2__8130_, data_stage_2__8129_, data_stage_2__8128_, data_stage_2__8127_, data_stage_2__8126_, data_stage_2__8125_, data_stage_2__8124_, data_stage_2__8123_, data_stage_2__8122_, data_stage_2__8121_, data_stage_2__8120_, data_stage_2__8119_, data_stage_2__8118_, data_stage_2__8117_, data_stage_2__8116_, data_stage_2__8115_, data_stage_2__8114_, data_stage_2__8113_, data_stage_2__8112_, data_stage_2__8111_, data_stage_2__8110_, data_stage_2__8109_, data_stage_2__8108_, data_stage_2__8107_, data_stage_2__8106_, data_stage_2__8105_, data_stage_2__8104_, data_stage_2__8103_, data_stage_2__8102_, data_stage_2__8101_, data_stage_2__8100_, data_stage_2__8099_, data_stage_2__8098_, data_stage_2__8097_, data_stage_2__8096_, data_stage_2__8095_, data_stage_2__8094_, data_stage_2__8093_, data_stage_2__8092_, data_stage_2__8091_, data_stage_2__8090_, data_stage_2__8089_, data_stage_2__8088_, data_stage_2__8087_, data_stage_2__8086_, data_stage_2__8085_, data_stage_2__8084_, data_stage_2__8083_, data_stage_2__8082_, data_stage_2__8081_, data_stage_2__8080_, data_stage_2__8079_, data_stage_2__8078_, data_stage_2__8077_, data_stage_2__8076_, data_stage_2__8075_, data_stage_2__8074_, data_stage_2__8073_, data_stage_2__8072_, data_stage_2__8071_, data_stage_2__8070_, data_stage_2__8069_, data_stage_2__8068_, data_stage_2__8067_, data_stage_2__8066_, data_stage_2__8065_, data_stage_2__8064_, data_stage_2__8063_, data_stage_2__8062_, data_stage_2__8061_, data_stage_2__8060_, data_stage_2__8059_, data_stage_2__8058_, data_stage_2__8057_, data_stage_2__8056_, data_stage_2__8055_, data_stage_2__8054_, data_stage_2__8053_, data_stage_2__8052_, data_stage_2__8051_, data_stage_2__8050_, data_stage_2__8049_, data_stage_2__8048_, data_stage_2__8047_, data_stage_2__8046_, data_stage_2__8045_, data_stage_2__8044_, data_stage_2__8043_, data_stage_2__8042_, data_stage_2__8041_, data_stage_2__8040_, data_stage_2__8039_, data_stage_2__8038_, data_stage_2__8037_, data_stage_2__8036_, data_stage_2__8035_, data_stage_2__8034_, data_stage_2__8033_, data_stage_2__8032_, data_stage_2__8031_, data_stage_2__8030_, data_stage_2__8029_, data_stage_2__8028_, data_stage_2__8027_, data_stage_2__8026_, data_stage_2__8025_, data_stage_2__8024_, data_stage_2__8023_, data_stage_2__8022_, data_stage_2__8021_, data_stage_2__8020_, data_stage_2__8019_, data_stage_2__8018_, data_stage_2__8017_, data_stage_2__8016_, data_stage_2__8015_, data_stage_2__8014_, data_stage_2__8013_, data_stage_2__8012_, data_stage_2__8011_, data_stage_2__8010_, data_stage_2__8009_, data_stage_2__8008_, data_stage_2__8007_, data_stage_2__8006_, data_stage_2__8005_, data_stage_2__8004_, data_stage_2__8003_, data_stage_2__8002_, data_stage_2__8001_, data_stage_2__8000_, data_stage_2__7999_, data_stage_2__7998_, data_stage_2__7997_, data_stage_2__7996_, data_stage_2__7995_, data_stage_2__7994_, data_stage_2__7993_, data_stage_2__7992_, data_stage_2__7991_, data_stage_2__7990_, data_stage_2__7989_, data_stage_2__7988_, data_stage_2__7987_, data_stage_2__7986_, data_stage_2__7985_, data_stage_2__7984_, data_stage_2__7983_, data_stage_2__7982_, data_stage_2__7981_, data_stage_2__7980_, data_stage_2__7979_, data_stage_2__7978_, data_stage_2__7977_, data_stage_2__7976_, data_stage_2__7975_, data_stage_2__7974_, data_stage_2__7973_, data_stage_2__7972_, data_stage_2__7971_, data_stage_2__7970_, data_stage_2__7969_, data_stage_2__7968_, data_stage_2__7967_, data_stage_2__7966_, data_stage_2__7965_, data_stage_2__7964_, data_stage_2__7963_, data_stage_2__7962_, data_stage_2__7961_, data_stage_2__7960_, data_stage_2__7959_, data_stage_2__7958_, data_stage_2__7957_, data_stage_2__7956_, data_stage_2__7955_, data_stage_2__7954_, data_stage_2__7953_, data_stage_2__7952_, data_stage_2__7951_, data_stage_2__7950_, data_stage_2__7949_, data_stage_2__7948_, data_stage_2__7947_, data_stage_2__7946_, data_stage_2__7945_, data_stage_2__7944_, data_stage_2__7943_, data_stage_2__7942_, data_stage_2__7941_, data_stage_2__7940_, data_stage_2__7939_, data_stage_2__7938_, data_stage_2__7937_, data_stage_2__7936_, data_stage_2__7935_, data_stage_2__7934_, data_stage_2__7933_, data_stage_2__7932_, data_stage_2__7931_, data_stage_2__7930_, data_stage_2__7929_, data_stage_2__7928_, data_stage_2__7927_, data_stage_2__7926_, data_stage_2__7925_, data_stage_2__7924_, data_stage_2__7923_, data_stage_2__7922_, data_stage_2__7921_, data_stage_2__7920_, data_stage_2__7919_, data_stage_2__7918_, data_stage_2__7917_, data_stage_2__7916_, data_stage_2__7915_, data_stage_2__7914_, data_stage_2__7913_, data_stage_2__7912_, data_stage_2__7911_, data_stage_2__7910_, data_stage_2__7909_, data_stage_2__7908_, data_stage_2__7907_, data_stage_2__7906_, data_stage_2__7905_, data_stage_2__7904_, data_stage_2__7903_, data_stage_2__7902_, data_stage_2__7901_, data_stage_2__7900_, data_stage_2__7899_, data_stage_2__7898_, data_stage_2__7897_, data_stage_2__7896_, data_stage_2__7895_, data_stage_2__7894_, data_stage_2__7893_, data_stage_2__7892_, data_stage_2__7891_, data_stage_2__7890_, data_stage_2__7889_, data_stage_2__7888_, data_stage_2__7887_, data_stage_2__7886_, data_stage_2__7885_, data_stage_2__7884_, data_stage_2__7883_, data_stage_2__7882_, data_stage_2__7881_, data_stage_2__7880_, data_stage_2__7879_, data_stage_2__7878_, data_stage_2__7877_, data_stage_2__7876_, data_stage_2__7875_, data_stage_2__7874_, data_stage_2__7873_, data_stage_2__7872_, data_stage_2__7871_, data_stage_2__7870_, data_stage_2__7869_, data_stage_2__7868_, data_stage_2__7867_, data_stage_2__7866_, data_stage_2__7865_, data_stage_2__7864_, data_stage_2__7863_, data_stage_2__7862_, data_stage_2__7861_, data_stage_2__7860_, data_stage_2__7859_, data_stage_2__7858_, data_stage_2__7857_, data_stage_2__7856_, data_stage_2__7855_, data_stage_2__7854_, data_stage_2__7853_, data_stage_2__7852_, data_stage_2__7851_, data_stage_2__7850_, data_stage_2__7849_, data_stage_2__7848_, data_stage_2__7847_, data_stage_2__7846_, data_stage_2__7845_, data_stage_2__7844_, data_stage_2__7843_, data_stage_2__7842_, data_stage_2__7841_, data_stage_2__7840_, data_stage_2__7839_, data_stage_2__7838_, data_stage_2__7837_, data_stage_2__7836_, data_stage_2__7835_, data_stage_2__7834_, data_stage_2__7833_, data_stage_2__7832_, data_stage_2__7831_, data_stage_2__7830_, data_stage_2__7829_, data_stage_2__7828_, data_stage_2__7827_, data_stage_2__7826_, data_stage_2__7825_, data_stage_2__7824_, data_stage_2__7823_, data_stage_2__7822_, data_stage_2__7821_, data_stage_2__7820_, data_stage_2__7819_, data_stage_2__7818_, data_stage_2__7817_, data_stage_2__7816_, data_stage_2__7815_, data_stage_2__7814_, data_stage_2__7813_, data_stage_2__7812_, data_stage_2__7811_, data_stage_2__7810_, data_stage_2__7809_, data_stage_2__7808_, data_stage_2__7807_, data_stage_2__7806_, data_stage_2__7805_, data_stage_2__7804_, data_stage_2__7803_, data_stage_2__7802_, data_stage_2__7801_, data_stage_2__7800_, data_stage_2__7799_, data_stage_2__7798_, data_stage_2__7797_, data_stage_2__7796_, data_stage_2__7795_, data_stage_2__7794_, data_stage_2__7793_, data_stage_2__7792_, data_stage_2__7791_, data_stage_2__7790_, data_stage_2__7789_, data_stage_2__7788_, data_stage_2__7787_, data_stage_2__7786_, data_stage_2__7785_, data_stage_2__7784_, data_stage_2__7783_, data_stage_2__7782_, data_stage_2__7781_, data_stage_2__7780_, data_stage_2__7779_, data_stage_2__7778_, data_stage_2__7777_, data_stage_2__7776_, data_stage_2__7775_, data_stage_2__7774_, data_stage_2__7773_, data_stage_2__7772_, data_stage_2__7771_, data_stage_2__7770_, data_stage_2__7769_, data_stage_2__7768_, data_stage_2__7767_, data_stage_2__7766_, data_stage_2__7765_, data_stage_2__7764_, data_stage_2__7763_, data_stage_2__7762_, data_stage_2__7761_, data_stage_2__7760_, data_stage_2__7759_, data_stage_2__7758_, data_stage_2__7757_, data_stage_2__7756_, data_stage_2__7755_, data_stage_2__7754_, data_stage_2__7753_, data_stage_2__7752_, data_stage_2__7751_, data_stage_2__7750_, data_stage_2__7749_, data_stage_2__7748_, data_stage_2__7747_, data_stage_2__7746_, data_stage_2__7745_, data_stage_2__7744_, data_stage_2__7743_, data_stage_2__7742_, data_stage_2__7741_, data_stage_2__7740_, data_stage_2__7739_, data_stage_2__7738_, data_stage_2__7737_, data_stage_2__7736_, data_stage_2__7735_, data_stage_2__7734_, data_stage_2__7733_, data_stage_2__7732_, data_stage_2__7731_, data_stage_2__7730_, data_stage_2__7729_, data_stage_2__7728_, data_stage_2__7727_, data_stage_2__7726_, data_stage_2__7725_, data_stage_2__7724_, data_stage_2__7723_, data_stage_2__7722_, data_stage_2__7721_, data_stage_2__7720_, data_stage_2__7719_, data_stage_2__7718_, data_stage_2__7717_, data_stage_2__7716_, data_stage_2__7715_, data_stage_2__7714_, data_stage_2__7713_, data_stage_2__7712_, data_stage_2__7711_, data_stage_2__7710_, data_stage_2__7709_, data_stage_2__7708_, data_stage_2__7707_, data_stage_2__7706_, data_stage_2__7705_, data_stage_2__7704_, data_stage_2__7703_, data_stage_2__7702_, data_stage_2__7701_, data_stage_2__7700_, data_stage_2__7699_, data_stage_2__7698_, data_stage_2__7697_, data_stage_2__7696_, data_stage_2__7695_, data_stage_2__7694_, data_stage_2__7693_, data_stage_2__7692_, data_stage_2__7691_, data_stage_2__7690_, data_stage_2__7689_, data_stage_2__7688_, data_stage_2__7687_, data_stage_2__7686_, data_stage_2__7685_, data_stage_2__7684_, data_stage_2__7683_, data_stage_2__7682_, data_stage_2__7681_, data_stage_2__7680_ })
  );


  bsg_swap_width_p512
  mux_stage_2__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_2__1023_, data_stage_2__1022_, data_stage_2__1021_, data_stage_2__1020_, data_stage_2__1019_, data_stage_2__1018_, data_stage_2__1017_, data_stage_2__1016_, data_stage_2__1015_, data_stage_2__1014_, data_stage_2__1013_, data_stage_2__1012_, data_stage_2__1011_, data_stage_2__1010_, data_stage_2__1009_, data_stage_2__1008_, data_stage_2__1007_, data_stage_2__1006_, data_stage_2__1005_, data_stage_2__1004_, data_stage_2__1003_, data_stage_2__1002_, data_stage_2__1001_, data_stage_2__1000_, data_stage_2__999_, data_stage_2__998_, data_stage_2__997_, data_stage_2__996_, data_stage_2__995_, data_stage_2__994_, data_stage_2__993_, data_stage_2__992_, data_stage_2__991_, data_stage_2__990_, data_stage_2__989_, data_stage_2__988_, data_stage_2__987_, data_stage_2__986_, data_stage_2__985_, data_stage_2__984_, data_stage_2__983_, data_stage_2__982_, data_stage_2__981_, data_stage_2__980_, data_stage_2__979_, data_stage_2__978_, data_stage_2__977_, data_stage_2__976_, data_stage_2__975_, data_stage_2__974_, data_stage_2__973_, data_stage_2__972_, data_stage_2__971_, data_stage_2__970_, data_stage_2__969_, data_stage_2__968_, data_stage_2__967_, data_stage_2__966_, data_stage_2__965_, data_stage_2__964_, data_stage_2__963_, data_stage_2__962_, data_stage_2__961_, data_stage_2__960_, data_stage_2__959_, data_stage_2__958_, data_stage_2__957_, data_stage_2__956_, data_stage_2__955_, data_stage_2__954_, data_stage_2__953_, data_stage_2__952_, data_stage_2__951_, data_stage_2__950_, data_stage_2__949_, data_stage_2__948_, data_stage_2__947_, data_stage_2__946_, data_stage_2__945_, data_stage_2__944_, data_stage_2__943_, data_stage_2__942_, data_stage_2__941_, data_stage_2__940_, data_stage_2__939_, data_stage_2__938_, data_stage_2__937_, data_stage_2__936_, data_stage_2__935_, data_stage_2__934_, data_stage_2__933_, data_stage_2__932_, data_stage_2__931_, data_stage_2__930_, data_stage_2__929_, data_stage_2__928_, data_stage_2__927_, data_stage_2__926_, data_stage_2__925_, data_stage_2__924_, data_stage_2__923_, data_stage_2__922_, data_stage_2__921_, data_stage_2__920_, data_stage_2__919_, data_stage_2__918_, data_stage_2__917_, data_stage_2__916_, data_stage_2__915_, data_stage_2__914_, data_stage_2__913_, data_stage_2__912_, data_stage_2__911_, data_stage_2__910_, data_stage_2__909_, data_stage_2__908_, data_stage_2__907_, data_stage_2__906_, data_stage_2__905_, data_stage_2__904_, data_stage_2__903_, data_stage_2__902_, data_stage_2__901_, data_stage_2__900_, data_stage_2__899_, data_stage_2__898_, data_stage_2__897_, data_stage_2__896_, data_stage_2__895_, data_stage_2__894_, data_stage_2__893_, data_stage_2__892_, data_stage_2__891_, data_stage_2__890_, data_stage_2__889_, data_stage_2__888_, data_stage_2__887_, data_stage_2__886_, data_stage_2__885_, data_stage_2__884_, data_stage_2__883_, data_stage_2__882_, data_stage_2__881_, data_stage_2__880_, data_stage_2__879_, data_stage_2__878_, data_stage_2__877_, data_stage_2__876_, data_stage_2__875_, data_stage_2__874_, data_stage_2__873_, data_stage_2__872_, data_stage_2__871_, data_stage_2__870_, data_stage_2__869_, data_stage_2__868_, data_stage_2__867_, data_stage_2__866_, data_stage_2__865_, data_stage_2__864_, data_stage_2__863_, data_stage_2__862_, data_stage_2__861_, data_stage_2__860_, data_stage_2__859_, data_stage_2__858_, data_stage_2__857_, data_stage_2__856_, data_stage_2__855_, data_stage_2__854_, data_stage_2__853_, data_stage_2__852_, data_stage_2__851_, data_stage_2__850_, data_stage_2__849_, data_stage_2__848_, data_stage_2__847_, data_stage_2__846_, data_stage_2__845_, data_stage_2__844_, data_stage_2__843_, data_stage_2__842_, data_stage_2__841_, data_stage_2__840_, data_stage_2__839_, data_stage_2__838_, data_stage_2__837_, data_stage_2__836_, data_stage_2__835_, data_stage_2__834_, data_stage_2__833_, data_stage_2__832_, data_stage_2__831_, data_stage_2__830_, data_stage_2__829_, data_stage_2__828_, data_stage_2__827_, data_stage_2__826_, data_stage_2__825_, data_stage_2__824_, data_stage_2__823_, data_stage_2__822_, data_stage_2__821_, data_stage_2__820_, data_stage_2__819_, data_stage_2__818_, data_stage_2__817_, data_stage_2__816_, data_stage_2__815_, data_stage_2__814_, data_stage_2__813_, data_stage_2__812_, data_stage_2__811_, data_stage_2__810_, data_stage_2__809_, data_stage_2__808_, data_stage_2__807_, data_stage_2__806_, data_stage_2__805_, data_stage_2__804_, data_stage_2__803_, data_stage_2__802_, data_stage_2__801_, data_stage_2__800_, data_stage_2__799_, data_stage_2__798_, data_stage_2__797_, data_stage_2__796_, data_stage_2__795_, data_stage_2__794_, data_stage_2__793_, data_stage_2__792_, data_stage_2__791_, data_stage_2__790_, data_stage_2__789_, data_stage_2__788_, data_stage_2__787_, data_stage_2__786_, data_stage_2__785_, data_stage_2__784_, data_stage_2__783_, data_stage_2__782_, data_stage_2__781_, data_stage_2__780_, data_stage_2__779_, data_stage_2__778_, data_stage_2__777_, data_stage_2__776_, data_stage_2__775_, data_stage_2__774_, data_stage_2__773_, data_stage_2__772_, data_stage_2__771_, data_stage_2__770_, data_stage_2__769_, data_stage_2__768_, data_stage_2__767_, data_stage_2__766_, data_stage_2__765_, data_stage_2__764_, data_stage_2__763_, data_stage_2__762_, data_stage_2__761_, data_stage_2__760_, data_stage_2__759_, data_stage_2__758_, data_stage_2__757_, data_stage_2__756_, data_stage_2__755_, data_stage_2__754_, data_stage_2__753_, data_stage_2__752_, data_stage_2__751_, data_stage_2__750_, data_stage_2__749_, data_stage_2__748_, data_stage_2__747_, data_stage_2__746_, data_stage_2__745_, data_stage_2__744_, data_stage_2__743_, data_stage_2__742_, data_stage_2__741_, data_stage_2__740_, data_stage_2__739_, data_stage_2__738_, data_stage_2__737_, data_stage_2__736_, data_stage_2__735_, data_stage_2__734_, data_stage_2__733_, data_stage_2__732_, data_stage_2__731_, data_stage_2__730_, data_stage_2__729_, data_stage_2__728_, data_stage_2__727_, data_stage_2__726_, data_stage_2__725_, data_stage_2__724_, data_stage_2__723_, data_stage_2__722_, data_stage_2__721_, data_stage_2__720_, data_stage_2__719_, data_stage_2__718_, data_stage_2__717_, data_stage_2__716_, data_stage_2__715_, data_stage_2__714_, data_stage_2__713_, data_stage_2__712_, data_stage_2__711_, data_stage_2__710_, data_stage_2__709_, data_stage_2__708_, data_stage_2__707_, data_stage_2__706_, data_stage_2__705_, data_stage_2__704_, data_stage_2__703_, data_stage_2__702_, data_stage_2__701_, data_stage_2__700_, data_stage_2__699_, data_stage_2__698_, data_stage_2__697_, data_stage_2__696_, data_stage_2__695_, data_stage_2__694_, data_stage_2__693_, data_stage_2__692_, data_stage_2__691_, data_stage_2__690_, data_stage_2__689_, data_stage_2__688_, data_stage_2__687_, data_stage_2__686_, data_stage_2__685_, data_stage_2__684_, data_stage_2__683_, data_stage_2__682_, data_stage_2__681_, data_stage_2__680_, data_stage_2__679_, data_stage_2__678_, data_stage_2__677_, data_stage_2__676_, data_stage_2__675_, data_stage_2__674_, data_stage_2__673_, data_stage_2__672_, data_stage_2__671_, data_stage_2__670_, data_stage_2__669_, data_stage_2__668_, data_stage_2__667_, data_stage_2__666_, data_stage_2__665_, data_stage_2__664_, data_stage_2__663_, data_stage_2__662_, data_stage_2__661_, data_stage_2__660_, data_stage_2__659_, data_stage_2__658_, data_stage_2__657_, data_stage_2__656_, data_stage_2__655_, data_stage_2__654_, data_stage_2__653_, data_stage_2__652_, data_stage_2__651_, data_stage_2__650_, data_stage_2__649_, data_stage_2__648_, data_stage_2__647_, data_stage_2__646_, data_stage_2__645_, data_stage_2__644_, data_stage_2__643_, data_stage_2__642_, data_stage_2__641_, data_stage_2__640_, data_stage_2__639_, data_stage_2__638_, data_stage_2__637_, data_stage_2__636_, data_stage_2__635_, data_stage_2__634_, data_stage_2__633_, data_stage_2__632_, data_stage_2__631_, data_stage_2__630_, data_stage_2__629_, data_stage_2__628_, data_stage_2__627_, data_stage_2__626_, data_stage_2__625_, data_stage_2__624_, data_stage_2__623_, data_stage_2__622_, data_stage_2__621_, data_stage_2__620_, data_stage_2__619_, data_stage_2__618_, data_stage_2__617_, data_stage_2__616_, data_stage_2__615_, data_stage_2__614_, data_stage_2__613_, data_stage_2__612_, data_stage_2__611_, data_stage_2__610_, data_stage_2__609_, data_stage_2__608_, data_stage_2__607_, data_stage_2__606_, data_stage_2__605_, data_stage_2__604_, data_stage_2__603_, data_stage_2__602_, data_stage_2__601_, data_stage_2__600_, data_stage_2__599_, data_stage_2__598_, data_stage_2__597_, data_stage_2__596_, data_stage_2__595_, data_stage_2__594_, data_stage_2__593_, data_stage_2__592_, data_stage_2__591_, data_stage_2__590_, data_stage_2__589_, data_stage_2__588_, data_stage_2__587_, data_stage_2__586_, data_stage_2__585_, data_stage_2__584_, data_stage_2__583_, data_stage_2__582_, data_stage_2__581_, data_stage_2__580_, data_stage_2__579_, data_stage_2__578_, data_stage_2__577_, data_stage_2__576_, data_stage_2__575_, data_stage_2__574_, data_stage_2__573_, data_stage_2__572_, data_stage_2__571_, data_stage_2__570_, data_stage_2__569_, data_stage_2__568_, data_stage_2__567_, data_stage_2__566_, data_stage_2__565_, data_stage_2__564_, data_stage_2__563_, data_stage_2__562_, data_stage_2__561_, data_stage_2__560_, data_stage_2__559_, data_stage_2__558_, data_stage_2__557_, data_stage_2__556_, data_stage_2__555_, data_stage_2__554_, data_stage_2__553_, data_stage_2__552_, data_stage_2__551_, data_stage_2__550_, data_stage_2__549_, data_stage_2__548_, data_stage_2__547_, data_stage_2__546_, data_stage_2__545_, data_stage_2__544_, data_stage_2__543_, data_stage_2__542_, data_stage_2__541_, data_stage_2__540_, data_stage_2__539_, data_stage_2__538_, data_stage_2__537_, data_stage_2__536_, data_stage_2__535_, data_stage_2__534_, data_stage_2__533_, data_stage_2__532_, data_stage_2__531_, data_stage_2__530_, data_stage_2__529_, data_stage_2__528_, data_stage_2__527_, data_stage_2__526_, data_stage_2__525_, data_stage_2__524_, data_stage_2__523_, data_stage_2__522_, data_stage_2__521_, data_stage_2__520_, data_stage_2__519_, data_stage_2__518_, data_stage_2__517_, data_stage_2__516_, data_stage_2__515_, data_stage_2__514_, data_stage_2__513_, data_stage_2__512_, data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_, data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_, data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_, data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__1023_, data_stage_3__1022_, data_stage_3__1021_, data_stage_3__1020_, data_stage_3__1019_, data_stage_3__1018_, data_stage_3__1017_, data_stage_3__1016_, data_stage_3__1015_, data_stage_3__1014_, data_stage_3__1013_, data_stage_3__1012_, data_stage_3__1011_, data_stage_3__1010_, data_stage_3__1009_, data_stage_3__1008_, data_stage_3__1007_, data_stage_3__1006_, data_stage_3__1005_, data_stage_3__1004_, data_stage_3__1003_, data_stage_3__1002_, data_stage_3__1001_, data_stage_3__1000_, data_stage_3__999_, data_stage_3__998_, data_stage_3__997_, data_stage_3__996_, data_stage_3__995_, data_stage_3__994_, data_stage_3__993_, data_stage_3__992_, data_stage_3__991_, data_stage_3__990_, data_stage_3__989_, data_stage_3__988_, data_stage_3__987_, data_stage_3__986_, data_stage_3__985_, data_stage_3__984_, data_stage_3__983_, data_stage_3__982_, data_stage_3__981_, data_stage_3__980_, data_stage_3__979_, data_stage_3__978_, data_stage_3__977_, data_stage_3__976_, data_stage_3__975_, data_stage_3__974_, data_stage_3__973_, data_stage_3__972_, data_stage_3__971_, data_stage_3__970_, data_stage_3__969_, data_stage_3__968_, data_stage_3__967_, data_stage_3__966_, data_stage_3__965_, data_stage_3__964_, data_stage_3__963_, data_stage_3__962_, data_stage_3__961_, data_stage_3__960_, data_stage_3__959_, data_stage_3__958_, data_stage_3__957_, data_stage_3__956_, data_stage_3__955_, data_stage_3__954_, data_stage_3__953_, data_stage_3__952_, data_stage_3__951_, data_stage_3__950_, data_stage_3__949_, data_stage_3__948_, data_stage_3__947_, data_stage_3__946_, data_stage_3__945_, data_stage_3__944_, data_stage_3__943_, data_stage_3__942_, data_stage_3__941_, data_stage_3__940_, data_stage_3__939_, data_stage_3__938_, data_stage_3__937_, data_stage_3__936_, data_stage_3__935_, data_stage_3__934_, data_stage_3__933_, data_stage_3__932_, data_stage_3__931_, data_stage_3__930_, data_stage_3__929_, data_stage_3__928_, data_stage_3__927_, data_stage_3__926_, data_stage_3__925_, data_stage_3__924_, data_stage_3__923_, data_stage_3__922_, data_stage_3__921_, data_stage_3__920_, data_stage_3__919_, data_stage_3__918_, data_stage_3__917_, data_stage_3__916_, data_stage_3__915_, data_stage_3__914_, data_stage_3__913_, data_stage_3__912_, data_stage_3__911_, data_stage_3__910_, data_stage_3__909_, data_stage_3__908_, data_stage_3__907_, data_stage_3__906_, data_stage_3__905_, data_stage_3__904_, data_stage_3__903_, data_stage_3__902_, data_stage_3__901_, data_stage_3__900_, data_stage_3__899_, data_stage_3__898_, data_stage_3__897_, data_stage_3__896_, data_stage_3__895_, data_stage_3__894_, data_stage_3__893_, data_stage_3__892_, data_stage_3__891_, data_stage_3__890_, data_stage_3__889_, data_stage_3__888_, data_stage_3__887_, data_stage_3__886_, data_stage_3__885_, data_stage_3__884_, data_stage_3__883_, data_stage_3__882_, data_stage_3__881_, data_stage_3__880_, data_stage_3__879_, data_stage_3__878_, data_stage_3__877_, data_stage_3__876_, data_stage_3__875_, data_stage_3__874_, data_stage_3__873_, data_stage_3__872_, data_stage_3__871_, data_stage_3__870_, data_stage_3__869_, data_stage_3__868_, data_stage_3__867_, data_stage_3__866_, data_stage_3__865_, data_stage_3__864_, data_stage_3__863_, data_stage_3__862_, data_stage_3__861_, data_stage_3__860_, data_stage_3__859_, data_stage_3__858_, data_stage_3__857_, data_stage_3__856_, data_stage_3__855_, data_stage_3__854_, data_stage_3__853_, data_stage_3__852_, data_stage_3__851_, data_stage_3__850_, data_stage_3__849_, data_stage_3__848_, data_stage_3__847_, data_stage_3__846_, data_stage_3__845_, data_stage_3__844_, data_stage_3__843_, data_stage_3__842_, data_stage_3__841_, data_stage_3__840_, data_stage_3__839_, data_stage_3__838_, data_stage_3__837_, data_stage_3__836_, data_stage_3__835_, data_stage_3__834_, data_stage_3__833_, data_stage_3__832_, data_stage_3__831_, data_stage_3__830_, data_stage_3__829_, data_stage_3__828_, data_stage_3__827_, data_stage_3__826_, data_stage_3__825_, data_stage_3__824_, data_stage_3__823_, data_stage_3__822_, data_stage_3__821_, data_stage_3__820_, data_stage_3__819_, data_stage_3__818_, data_stage_3__817_, data_stage_3__816_, data_stage_3__815_, data_stage_3__814_, data_stage_3__813_, data_stage_3__812_, data_stage_3__811_, data_stage_3__810_, data_stage_3__809_, data_stage_3__808_, data_stage_3__807_, data_stage_3__806_, data_stage_3__805_, data_stage_3__804_, data_stage_3__803_, data_stage_3__802_, data_stage_3__801_, data_stage_3__800_, data_stage_3__799_, data_stage_3__798_, data_stage_3__797_, data_stage_3__796_, data_stage_3__795_, data_stage_3__794_, data_stage_3__793_, data_stage_3__792_, data_stage_3__791_, data_stage_3__790_, data_stage_3__789_, data_stage_3__788_, data_stage_3__787_, data_stage_3__786_, data_stage_3__785_, data_stage_3__784_, data_stage_3__783_, data_stage_3__782_, data_stage_3__781_, data_stage_3__780_, data_stage_3__779_, data_stage_3__778_, data_stage_3__777_, data_stage_3__776_, data_stage_3__775_, data_stage_3__774_, data_stage_3__773_, data_stage_3__772_, data_stage_3__771_, data_stage_3__770_, data_stage_3__769_, data_stage_3__768_, data_stage_3__767_, data_stage_3__766_, data_stage_3__765_, data_stage_3__764_, data_stage_3__763_, data_stage_3__762_, data_stage_3__761_, data_stage_3__760_, data_stage_3__759_, data_stage_3__758_, data_stage_3__757_, data_stage_3__756_, data_stage_3__755_, data_stage_3__754_, data_stage_3__753_, data_stage_3__752_, data_stage_3__751_, data_stage_3__750_, data_stage_3__749_, data_stage_3__748_, data_stage_3__747_, data_stage_3__746_, data_stage_3__745_, data_stage_3__744_, data_stage_3__743_, data_stage_3__742_, data_stage_3__741_, data_stage_3__740_, data_stage_3__739_, data_stage_3__738_, data_stage_3__737_, data_stage_3__736_, data_stage_3__735_, data_stage_3__734_, data_stage_3__733_, data_stage_3__732_, data_stage_3__731_, data_stage_3__730_, data_stage_3__729_, data_stage_3__728_, data_stage_3__727_, data_stage_3__726_, data_stage_3__725_, data_stage_3__724_, data_stage_3__723_, data_stage_3__722_, data_stage_3__721_, data_stage_3__720_, data_stage_3__719_, data_stage_3__718_, data_stage_3__717_, data_stage_3__716_, data_stage_3__715_, data_stage_3__714_, data_stage_3__713_, data_stage_3__712_, data_stage_3__711_, data_stage_3__710_, data_stage_3__709_, data_stage_3__708_, data_stage_3__707_, data_stage_3__706_, data_stage_3__705_, data_stage_3__704_, data_stage_3__703_, data_stage_3__702_, data_stage_3__701_, data_stage_3__700_, data_stage_3__699_, data_stage_3__698_, data_stage_3__697_, data_stage_3__696_, data_stage_3__695_, data_stage_3__694_, data_stage_3__693_, data_stage_3__692_, data_stage_3__691_, data_stage_3__690_, data_stage_3__689_, data_stage_3__688_, data_stage_3__687_, data_stage_3__686_, data_stage_3__685_, data_stage_3__684_, data_stage_3__683_, data_stage_3__682_, data_stage_3__681_, data_stage_3__680_, data_stage_3__679_, data_stage_3__678_, data_stage_3__677_, data_stage_3__676_, data_stage_3__675_, data_stage_3__674_, data_stage_3__673_, data_stage_3__672_, data_stage_3__671_, data_stage_3__670_, data_stage_3__669_, data_stage_3__668_, data_stage_3__667_, data_stage_3__666_, data_stage_3__665_, data_stage_3__664_, data_stage_3__663_, data_stage_3__662_, data_stage_3__661_, data_stage_3__660_, data_stage_3__659_, data_stage_3__658_, data_stage_3__657_, data_stage_3__656_, data_stage_3__655_, data_stage_3__654_, data_stage_3__653_, data_stage_3__652_, data_stage_3__651_, data_stage_3__650_, data_stage_3__649_, data_stage_3__648_, data_stage_3__647_, data_stage_3__646_, data_stage_3__645_, data_stage_3__644_, data_stage_3__643_, data_stage_3__642_, data_stage_3__641_, data_stage_3__640_, data_stage_3__639_, data_stage_3__638_, data_stage_3__637_, data_stage_3__636_, data_stage_3__635_, data_stage_3__634_, data_stage_3__633_, data_stage_3__632_, data_stage_3__631_, data_stage_3__630_, data_stage_3__629_, data_stage_3__628_, data_stage_3__627_, data_stage_3__626_, data_stage_3__625_, data_stage_3__624_, data_stage_3__623_, data_stage_3__622_, data_stage_3__621_, data_stage_3__620_, data_stage_3__619_, data_stage_3__618_, data_stage_3__617_, data_stage_3__616_, data_stage_3__615_, data_stage_3__614_, data_stage_3__613_, data_stage_3__612_, data_stage_3__611_, data_stage_3__610_, data_stage_3__609_, data_stage_3__608_, data_stage_3__607_, data_stage_3__606_, data_stage_3__605_, data_stage_3__604_, data_stage_3__603_, data_stage_3__602_, data_stage_3__601_, data_stage_3__600_, data_stage_3__599_, data_stage_3__598_, data_stage_3__597_, data_stage_3__596_, data_stage_3__595_, data_stage_3__594_, data_stage_3__593_, data_stage_3__592_, data_stage_3__591_, data_stage_3__590_, data_stage_3__589_, data_stage_3__588_, data_stage_3__587_, data_stage_3__586_, data_stage_3__585_, data_stage_3__584_, data_stage_3__583_, data_stage_3__582_, data_stage_3__581_, data_stage_3__580_, data_stage_3__579_, data_stage_3__578_, data_stage_3__577_, data_stage_3__576_, data_stage_3__575_, data_stage_3__574_, data_stage_3__573_, data_stage_3__572_, data_stage_3__571_, data_stage_3__570_, data_stage_3__569_, data_stage_3__568_, data_stage_3__567_, data_stage_3__566_, data_stage_3__565_, data_stage_3__564_, data_stage_3__563_, data_stage_3__562_, data_stage_3__561_, data_stage_3__560_, data_stage_3__559_, data_stage_3__558_, data_stage_3__557_, data_stage_3__556_, data_stage_3__555_, data_stage_3__554_, data_stage_3__553_, data_stage_3__552_, data_stage_3__551_, data_stage_3__550_, data_stage_3__549_, data_stage_3__548_, data_stage_3__547_, data_stage_3__546_, data_stage_3__545_, data_stage_3__544_, data_stage_3__543_, data_stage_3__542_, data_stage_3__541_, data_stage_3__540_, data_stage_3__539_, data_stage_3__538_, data_stage_3__537_, data_stage_3__536_, data_stage_3__535_, data_stage_3__534_, data_stage_3__533_, data_stage_3__532_, data_stage_3__531_, data_stage_3__530_, data_stage_3__529_, data_stage_3__528_, data_stage_3__527_, data_stage_3__526_, data_stage_3__525_, data_stage_3__524_, data_stage_3__523_, data_stage_3__522_, data_stage_3__521_, data_stage_3__520_, data_stage_3__519_, data_stage_3__518_, data_stage_3__517_, data_stage_3__516_, data_stage_3__515_, data_stage_3__514_, data_stage_3__513_, data_stage_3__512_, data_stage_3__511_, data_stage_3__510_, data_stage_3__509_, data_stage_3__508_, data_stage_3__507_, data_stage_3__506_, data_stage_3__505_, data_stage_3__504_, data_stage_3__503_, data_stage_3__502_, data_stage_3__501_, data_stage_3__500_, data_stage_3__499_, data_stage_3__498_, data_stage_3__497_, data_stage_3__496_, data_stage_3__495_, data_stage_3__494_, data_stage_3__493_, data_stage_3__492_, data_stage_3__491_, data_stage_3__490_, data_stage_3__489_, data_stage_3__488_, data_stage_3__487_, data_stage_3__486_, data_stage_3__485_, data_stage_3__484_, data_stage_3__483_, data_stage_3__482_, data_stage_3__481_, data_stage_3__480_, data_stage_3__479_, data_stage_3__478_, data_stage_3__477_, data_stage_3__476_, data_stage_3__475_, data_stage_3__474_, data_stage_3__473_, data_stage_3__472_, data_stage_3__471_, data_stage_3__470_, data_stage_3__469_, data_stage_3__468_, data_stage_3__467_, data_stage_3__466_, data_stage_3__465_, data_stage_3__464_, data_stage_3__463_, data_stage_3__462_, data_stage_3__461_, data_stage_3__460_, data_stage_3__459_, data_stage_3__458_, data_stage_3__457_, data_stage_3__456_, data_stage_3__455_, data_stage_3__454_, data_stage_3__453_, data_stage_3__452_, data_stage_3__451_, data_stage_3__450_, data_stage_3__449_, data_stage_3__448_, data_stage_3__447_, data_stage_3__446_, data_stage_3__445_, data_stage_3__444_, data_stage_3__443_, data_stage_3__442_, data_stage_3__441_, data_stage_3__440_, data_stage_3__439_, data_stage_3__438_, data_stage_3__437_, data_stage_3__436_, data_stage_3__435_, data_stage_3__434_, data_stage_3__433_, data_stage_3__432_, data_stage_3__431_, data_stage_3__430_, data_stage_3__429_, data_stage_3__428_, data_stage_3__427_, data_stage_3__426_, data_stage_3__425_, data_stage_3__424_, data_stage_3__423_, data_stage_3__422_, data_stage_3__421_, data_stage_3__420_, data_stage_3__419_, data_stage_3__418_, data_stage_3__417_, data_stage_3__416_, data_stage_3__415_, data_stage_3__414_, data_stage_3__413_, data_stage_3__412_, data_stage_3__411_, data_stage_3__410_, data_stage_3__409_, data_stage_3__408_, data_stage_3__407_, data_stage_3__406_, data_stage_3__405_, data_stage_3__404_, data_stage_3__403_, data_stage_3__402_, data_stage_3__401_, data_stage_3__400_, data_stage_3__399_, data_stage_3__398_, data_stage_3__397_, data_stage_3__396_, data_stage_3__395_, data_stage_3__394_, data_stage_3__393_, data_stage_3__392_, data_stage_3__391_, data_stage_3__390_, data_stage_3__389_, data_stage_3__388_, data_stage_3__387_, data_stage_3__386_, data_stage_3__385_, data_stage_3__384_, data_stage_3__383_, data_stage_3__382_, data_stage_3__381_, data_stage_3__380_, data_stage_3__379_, data_stage_3__378_, data_stage_3__377_, data_stage_3__376_, data_stage_3__375_, data_stage_3__374_, data_stage_3__373_, data_stage_3__372_, data_stage_3__371_, data_stage_3__370_, data_stage_3__369_, data_stage_3__368_, data_stage_3__367_, data_stage_3__366_, data_stage_3__365_, data_stage_3__364_, data_stage_3__363_, data_stage_3__362_, data_stage_3__361_, data_stage_3__360_, data_stage_3__359_, data_stage_3__358_, data_stage_3__357_, data_stage_3__356_, data_stage_3__355_, data_stage_3__354_, data_stage_3__353_, data_stage_3__352_, data_stage_3__351_, data_stage_3__350_, data_stage_3__349_, data_stage_3__348_, data_stage_3__347_, data_stage_3__346_, data_stage_3__345_, data_stage_3__344_, data_stage_3__343_, data_stage_3__342_, data_stage_3__341_, data_stage_3__340_, data_stage_3__339_, data_stage_3__338_, data_stage_3__337_, data_stage_3__336_, data_stage_3__335_, data_stage_3__334_, data_stage_3__333_, data_stage_3__332_, data_stage_3__331_, data_stage_3__330_, data_stage_3__329_, data_stage_3__328_, data_stage_3__327_, data_stage_3__326_, data_stage_3__325_, data_stage_3__324_, data_stage_3__323_, data_stage_3__322_, data_stage_3__321_, data_stage_3__320_, data_stage_3__319_, data_stage_3__318_, data_stage_3__317_, data_stage_3__316_, data_stage_3__315_, data_stage_3__314_, data_stage_3__313_, data_stage_3__312_, data_stage_3__311_, data_stage_3__310_, data_stage_3__309_, data_stage_3__308_, data_stage_3__307_, data_stage_3__306_, data_stage_3__305_, data_stage_3__304_, data_stage_3__303_, data_stage_3__302_, data_stage_3__301_, data_stage_3__300_, data_stage_3__299_, data_stage_3__298_, data_stage_3__297_, data_stage_3__296_, data_stage_3__295_, data_stage_3__294_, data_stage_3__293_, data_stage_3__292_, data_stage_3__291_, data_stage_3__290_, data_stage_3__289_, data_stage_3__288_, data_stage_3__287_, data_stage_3__286_, data_stage_3__285_, data_stage_3__284_, data_stage_3__283_, data_stage_3__282_, data_stage_3__281_, data_stage_3__280_, data_stage_3__279_, data_stage_3__278_, data_stage_3__277_, data_stage_3__276_, data_stage_3__275_, data_stage_3__274_, data_stage_3__273_, data_stage_3__272_, data_stage_3__271_, data_stage_3__270_, data_stage_3__269_, data_stage_3__268_, data_stage_3__267_, data_stage_3__266_, data_stage_3__265_, data_stage_3__264_, data_stage_3__263_, data_stage_3__262_, data_stage_3__261_, data_stage_3__260_, data_stage_3__259_, data_stage_3__258_, data_stage_3__257_, data_stage_3__256_, data_stage_3__255_, data_stage_3__254_, data_stage_3__253_, data_stage_3__252_, data_stage_3__251_, data_stage_3__250_, data_stage_3__249_, data_stage_3__248_, data_stage_3__247_, data_stage_3__246_, data_stage_3__245_, data_stage_3__244_, data_stage_3__243_, data_stage_3__242_, data_stage_3__241_, data_stage_3__240_, data_stage_3__239_, data_stage_3__238_, data_stage_3__237_, data_stage_3__236_, data_stage_3__235_, data_stage_3__234_, data_stage_3__233_, data_stage_3__232_, data_stage_3__231_, data_stage_3__230_, data_stage_3__229_, data_stage_3__228_, data_stage_3__227_, data_stage_3__226_, data_stage_3__225_, data_stage_3__224_, data_stage_3__223_, data_stage_3__222_, data_stage_3__221_, data_stage_3__220_, data_stage_3__219_, data_stage_3__218_, data_stage_3__217_, data_stage_3__216_, data_stage_3__215_, data_stage_3__214_, data_stage_3__213_, data_stage_3__212_, data_stage_3__211_, data_stage_3__210_, data_stage_3__209_, data_stage_3__208_, data_stage_3__207_, data_stage_3__206_, data_stage_3__205_, data_stage_3__204_, data_stage_3__203_, data_stage_3__202_, data_stage_3__201_, data_stage_3__200_, data_stage_3__199_, data_stage_3__198_, data_stage_3__197_, data_stage_3__196_, data_stage_3__195_, data_stage_3__194_, data_stage_3__193_, data_stage_3__192_, data_stage_3__191_, data_stage_3__190_, data_stage_3__189_, data_stage_3__188_, data_stage_3__187_, data_stage_3__186_, data_stage_3__185_, data_stage_3__184_, data_stage_3__183_, data_stage_3__182_, data_stage_3__181_, data_stage_3__180_, data_stage_3__179_, data_stage_3__178_, data_stage_3__177_, data_stage_3__176_, data_stage_3__175_, data_stage_3__174_, data_stage_3__173_, data_stage_3__172_, data_stage_3__171_, data_stage_3__170_, data_stage_3__169_, data_stage_3__168_, data_stage_3__167_, data_stage_3__166_, data_stage_3__165_, data_stage_3__164_, data_stage_3__163_, data_stage_3__162_, data_stage_3__161_, data_stage_3__160_, data_stage_3__159_, data_stage_3__158_, data_stage_3__157_, data_stage_3__156_, data_stage_3__155_, data_stage_3__154_, data_stage_3__153_, data_stage_3__152_, data_stage_3__151_, data_stage_3__150_, data_stage_3__149_, data_stage_3__148_, data_stage_3__147_, data_stage_3__146_, data_stage_3__145_, data_stage_3__144_, data_stage_3__143_, data_stage_3__142_, data_stage_3__141_, data_stage_3__140_, data_stage_3__139_, data_stage_3__138_, data_stage_3__137_, data_stage_3__136_, data_stage_3__135_, data_stage_3__134_, data_stage_3__133_, data_stage_3__132_, data_stage_3__131_, data_stage_3__130_, data_stage_3__129_, data_stage_3__128_, data_stage_3__127_, data_stage_3__126_, data_stage_3__125_, data_stage_3__124_, data_stage_3__123_, data_stage_3__122_, data_stage_3__121_, data_stage_3__120_, data_stage_3__119_, data_stage_3__118_, data_stage_3__117_, data_stage_3__116_, data_stage_3__115_, data_stage_3__114_, data_stage_3__113_, data_stage_3__112_, data_stage_3__111_, data_stage_3__110_, data_stage_3__109_, data_stage_3__108_, data_stage_3__107_, data_stage_3__106_, data_stage_3__105_, data_stage_3__104_, data_stage_3__103_, data_stage_3__102_, data_stage_3__101_, data_stage_3__100_, data_stage_3__99_, data_stage_3__98_, data_stage_3__97_, data_stage_3__96_, data_stage_3__95_, data_stage_3__94_, data_stage_3__93_, data_stage_3__92_, data_stage_3__91_, data_stage_3__90_, data_stage_3__89_, data_stage_3__88_, data_stage_3__87_, data_stage_3__86_, data_stage_3__85_, data_stage_3__84_, data_stage_3__83_, data_stage_3__82_, data_stage_3__81_, data_stage_3__80_, data_stage_3__79_, data_stage_3__78_, data_stage_3__77_, data_stage_3__76_, data_stage_3__75_, data_stage_3__74_, data_stage_3__73_, data_stage_3__72_, data_stage_3__71_, data_stage_3__70_, data_stage_3__69_, data_stage_3__68_, data_stage_3__67_, data_stage_3__66_, data_stage_3__65_, data_stage_3__64_, data_stage_3__63_, data_stage_3__62_, data_stage_3__61_, data_stage_3__60_, data_stage_3__59_, data_stage_3__58_, data_stage_3__57_, data_stage_3__56_, data_stage_3__55_, data_stage_3__54_, data_stage_3__53_, data_stage_3__52_, data_stage_3__51_, data_stage_3__50_, data_stage_3__49_, data_stage_3__48_, data_stage_3__47_, data_stage_3__46_, data_stage_3__45_, data_stage_3__44_, data_stage_3__43_, data_stage_3__42_, data_stage_3__41_, data_stage_3__40_, data_stage_3__39_, data_stage_3__38_, data_stage_3__37_, data_stage_3__36_, data_stage_3__35_, data_stage_3__34_, data_stage_3__33_, data_stage_3__32_, data_stage_3__31_, data_stage_3__30_, data_stage_3__29_, data_stage_3__28_, data_stage_3__27_, data_stage_3__26_, data_stage_3__25_, data_stage_3__24_, data_stage_3__23_, data_stage_3__22_, data_stage_3__21_, data_stage_3__20_, data_stage_3__19_, data_stage_3__18_, data_stage_3__17_, data_stage_3__16_, data_stage_3__15_, data_stage_3__14_, data_stage_3__13_, data_stage_3__12_, data_stage_3__11_, data_stage_3__10_, data_stage_3__9_, data_stage_3__8_, data_stage_3__7_, data_stage_3__6_, data_stage_3__5_, data_stage_3__4_, data_stage_3__3_, data_stage_3__2_, data_stage_3__1_, data_stage_3__0_ })
  );


  bsg_swap_width_p512
  mux_stage_2__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_2__2047_, data_stage_2__2046_, data_stage_2__2045_, data_stage_2__2044_, data_stage_2__2043_, data_stage_2__2042_, data_stage_2__2041_, data_stage_2__2040_, data_stage_2__2039_, data_stage_2__2038_, data_stage_2__2037_, data_stage_2__2036_, data_stage_2__2035_, data_stage_2__2034_, data_stage_2__2033_, data_stage_2__2032_, data_stage_2__2031_, data_stage_2__2030_, data_stage_2__2029_, data_stage_2__2028_, data_stage_2__2027_, data_stage_2__2026_, data_stage_2__2025_, data_stage_2__2024_, data_stage_2__2023_, data_stage_2__2022_, data_stage_2__2021_, data_stage_2__2020_, data_stage_2__2019_, data_stage_2__2018_, data_stage_2__2017_, data_stage_2__2016_, data_stage_2__2015_, data_stage_2__2014_, data_stage_2__2013_, data_stage_2__2012_, data_stage_2__2011_, data_stage_2__2010_, data_stage_2__2009_, data_stage_2__2008_, data_stage_2__2007_, data_stage_2__2006_, data_stage_2__2005_, data_stage_2__2004_, data_stage_2__2003_, data_stage_2__2002_, data_stage_2__2001_, data_stage_2__2000_, data_stage_2__1999_, data_stage_2__1998_, data_stage_2__1997_, data_stage_2__1996_, data_stage_2__1995_, data_stage_2__1994_, data_stage_2__1993_, data_stage_2__1992_, data_stage_2__1991_, data_stage_2__1990_, data_stage_2__1989_, data_stage_2__1988_, data_stage_2__1987_, data_stage_2__1986_, data_stage_2__1985_, data_stage_2__1984_, data_stage_2__1983_, data_stage_2__1982_, data_stage_2__1981_, data_stage_2__1980_, data_stage_2__1979_, data_stage_2__1978_, data_stage_2__1977_, data_stage_2__1976_, data_stage_2__1975_, data_stage_2__1974_, data_stage_2__1973_, data_stage_2__1972_, data_stage_2__1971_, data_stage_2__1970_, data_stage_2__1969_, data_stage_2__1968_, data_stage_2__1967_, data_stage_2__1966_, data_stage_2__1965_, data_stage_2__1964_, data_stage_2__1963_, data_stage_2__1962_, data_stage_2__1961_, data_stage_2__1960_, data_stage_2__1959_, data_stage_2__1958_, data_stage_2__1957_, data_stage_2__1956_, data_stage_2__1955_, data_stage_2__1954_, data_stage_2__1953_, data_stage_2__1952_, data_stage_2__1951_, data_stage_2__1950_, data_stage_2__1949_, data_stage_2__1948_, data_stage_2__1947_, data_stage_2__1946_, data_stage_2__1945_, data_stage_2__1944_, data_stage_2__1943_, data_stage_2__1942_, data_stage_2__1941_, data_stage_2__1940_, data_stage_2__1939_, data_stage_2__1938_, data_stage_2__1937_, data_stage_2__1936_, data_stage_2__1935_, data_stage_2__1934_, data_stage_2__1933_, data_stage_2__1932_, data_stage_2__1931_, data_stage_2__1930_, data_stage_2__1929_, data_stage_2__1928_, data_stage_2__1927_, data_stage_2__1926_, data_stage_2__1925_, data_stage_2__1924_, data_stage_2__1923_, data_stage_2__1922_, data_stage_2__1921_, data_stage_2__1920_, data_stage_2__1919_, data_stage_2__1918_, data_stage_2__1917_, data_stage_2__1916_, data_stage_2__1915_, data_stage_2__1914_, data_stage_2__1913_, data_stage_2__1912_, data_stage_2__1911_, data_stage_2__1910_, data_stage_2__1909_, data_stage_2__1908_, data_stage_2__1907_, data_stage_2__1906_, data_stage_2__1905_, data_stage_2__1904_, data_stage_2__1903_, data_stage_2__1902_, data_stage_2__1901_, data_stage_2__1900_, data_stage_2__1899_, data_stage_2__1898_, data_stage_2__1897_, data_stage_2__1896_, data_stage_2__1895_, data_stage_2__1894_, data_stage_2__1893_, data_stage_2__1892_, data_stage_2__1891_, data_stage_2__1890_, data_stage_2__1889_, data_stage_2__1888_, data_stage_2__1887_, data_stage_2__1886_, data_stage_2__1885_, data_stage_2__1884_, data_stage_2__1883_, data_stage_2__1882_, data_stage_2__1881_, data_stage_2__1880_, data_stage_2__1879_, data_stage_2__1878_, data_stage_2__1877_, data_stage_2__1876_, data_stage_2__1875_, data_stage_2__1874_, data_stage_2__1873_, data_stage_2__1872_, data_stage_2__1871_, data_stage_2__1870_, data_stage_2__1869_, data_stage_2__1868_, data_stage_2__1867_, data_stage_2__1866_, data_stage_2__1865_, data_stage_2__1864_, data_stage_2__1863_, data_stage_2__1862_, data_stage_2__1861_, data_stage_2__1860_, data_stage_2__1859_, data_stage_2__1858_, data_stage_2__1857_, data_stage_2__1856_, data_stage_2__1855_, data_stage_2__1854_, data_stage_2__1853_, data_stage_2__1852_, data_stage_2__1851_, data_stage_2__1850_, data_stage_2__1849_, data_stage_2__1848_, data_stage_2__1847_, data_stage_2__1846_, data_stage_2__1845_, data_stage_2__1844_, data_stage_2__1843_, data_stage_2__1842_, data_stage_2__1841_, data_stage_2__1840_, data_stage_2__1839_, data_stage_2__1838_, data_stage_2__1837_, data_stage_2__1836_, data_stage_2__1835_, data_stage_2__1834_, data_stage_2__1833_, data_stage_2__1832_, data_stage_2__1831_, data_stage_2__1830_, data_stage_2__1829_, data_stage_2__1828_, data_stage_2__1827_, data_stage_2__1826_, data_stage_2__1825_, data_stage_2__1824_, data_stage_2__1823_, data_stage_2__1822_, data_stage_2__1821_, data_stage_2__1820_, data_stage_2__1819_, data_stage_2__1818_, data_stage_2__1817_, data_stage_2__1816_, data_stage_2__1815_, data_stage_2__1814_, data_stage_2__1813_, data_stage_2__1812_, data_stage_2__1811_, data_stage_2__1810_, data_stage_2__1809_, data_stage_2__1808_, data_stage_2__1807_, data_stage_2__1806_, data_stage_2__1805_, data_stage_2__1804_, data_stage_2__1803_, data_stage_2__1802_, data_stage_2__1801_, data_stage_2__1800_, data_stage_2__1799_, data_stage_2__1798_, data_stage_2__1797_, data_stage_2__1796_, data_stage_2__1795_, data_stage_2__1794_, data_stage_2__1793_, data_stage_2__1792_, data_stage_2__1791_, data_stage_2__1790_, data_stage_2__1789_, data_stage_2__1788_, data_stage_2__1787_, data_stage_2__1786_, data_stage_2__1785_, data_stage_2__1784_, data_stage_2__1783_, data_stage_2__1782_, data_stage_2__1781_, data_stage_2__1780_, data_stage_2__1779_, data_stage_2__1778_, data_stage_2__1777_, data_stage_2__1776_, data_stage_2__1775_, data_stage_2__1774_, data_stage_2__1773_, data_stage_2__1772_, data_stage_2__1771_, data_stage_2__1770_, data_stage_2__1769_, data_stage_2__1768_, data_stage_2__1767_, data_stage_2__1766_, data_stage_2__1765_, data_stage_2__1764_, data_stage_2__1763_, data_stage_2__1762_, data_stage_2__1761_, data_stage_2__1760_, data_stage_2__1759_, data_stage_2__1758_, data_stage_2__1757_, data_stage_2__1756_, data_stage_2__1755_, data_stage_2__1754_, data_stage_2__1753_, data_stage_2__1752_, data_stage_2__1751_, data_stage_2__1750_, data_stage_2__1749_, data_stage_2__1748_, data_stage_2__1747_, data_stage_2__1746_, data_stage_2__1745_, data_stage_2__1744_, data_stage_2__1743_, data_stage_2__1742_, data_stage_2__1741_, data_stage_2__1740_, data_stage_2__1739_, data_stage_2__1738_, data_stage_2__1737_, data_stage_2__1736_, data_stage_2__1735_, data_stage_2__1734_, data_stage_2__1733_, data_stage_2__1732_, data_stage_2__1731_, data_stage_2__1730_, data_stage_2__1729_, data_stage_2__1728_, data_stage_2__1727_, data_stage_2__1726_, data_stage_2__1725_, data_stage_2__1724_, data_stage_2__1723_, data_stage_2__1722_, data_stage_2__1721_, data_stage_2__1720_, data_stage_2__1719_, data_stage_2__1718_, data_stage_2__1717_, data_stage_2__1716_, data_stage_2__1715_, data_stage_2__1714_, data_stage_2__1713_, data_stage_2__1712_, data_stage_2__1711_, data_stage_2__1710_, data_stage_2__1709_, data_stage_2__1708_, data_stage_2__1707_, data_stage_2__1706_, data_stage_2__1705_, data_stage_2__1704_, data_stage_2__1703_, data_stage_2__1702_, data_stage_2__1701_, data_stage_2__1700_, data_stage_2__1699_, data_stage_2__1698_, data_stage_2__1697_, data_stage_2__1696_, data_stage_2__1695_, data_stage_2__1694_, data_stage_2__1693_, data_stage_2__1692_, data_stage_2__1691_, data_stage_2__1690_, data_stage_2__1689_, data_stage_2__1688_, data_stage_2__1687_, data_stage_2__1686_, data_stage_2__1685_, data_stage_2__1684_, data_stage_2__1683_, data_stage_2__1682_, data_stage_2__1681_, data_stage_2__1680_, data_stage_2__1679_, data_stage_2__1678_, data_stage_2__1677_, data_stage_2__1676_, data_stage_2__1675_, data_stage_2__1674_, data_stage_2__1673_, data_stage_2__1672_, data_stage_2__1671_, data_stage_2__1670_, data_stage_2__1669_, data_stage_2__1668_, data_stage_2__1667_, data_stage_2__1666_, data_stage_2__1665_, data_stage_2__1664_, data_stage_2__1663_, data_stage_2__1662_, data_stage_2__1661_, data_stage_2__1660_, data_stage_2__1659_, data_stage_2__1658_, data_stage_2__1657_, data_stage_2__1656_, data_stage_2__1655_, data_stage_2__1654_, data_stage_2__1653_, data_stage_2__1652_, data_stage_2__1651_, data_stage_2__1650_, data_stage_2__1649_, data_stage_2__1648_, data_stage_2__1647_, data_stage_2__1646_, data_stage_2__1645_, data_stage_2__1644_, data_stage_2__1643_, data_stage_2__1642_, data_stage_2__1641_, data_stage_2__1640_, data_stage_2__1639_, data_stage_2__1638_, data_stage_2__1637_, data_stage_2__1636_, data_stage_2__1635_, data_stage_2__1634_, data_stage_2__1633_, data_stage_2__1632_, data_stage_2__1631_, data_stage_2__1630_, data_stage_2__1629_, data_stage_2__1628_, data_stage_2__1627_, data_stage_2__1626_, data_stage_2__1625_, data_stage_2__1624_, data_stage_2__1623_, data_stage_2__1622_, data_stage_2__1621_, data_stage_2__1620_, data_stage_2__1619_, data_stage_2__1618_, data_stage_2__1617_, data_stage_2__1616_, data_stage_2__1615_, data_stage_2__1614_, data_stage_2__1613_, data_stage_2__1612_, data_stage_2__1611_, data_stage_2__1610_, data_stage_2__1609_, data_stage_2__1608_, data_stage_2__1607_, data_stage_2__1606_, data_stage_2__1605_, data_stage_2__1604_, data_stage_2__1603_, data_stage_2__1602_, data_stage_2__1601_, data_stage_2__1600_, data_stage_2__1599_, data_stage_2__1598_, data_stage_2__1597_, data_stage_2__1596_, data_stage_2__1595_, data_stage_2__1594_, data_stage_2__1593_, data_stage_2__1592_, data_stage_2__1591_, data_stage_2__1590_, data_stage_2__1589_, data_stage_2__1588_, data_stage_2__1587_, data_stage_2__1586_, data_stage_2__1585_, data_stage_2__1584_, data_stage_2__1583_, data_stage_2__1582_, data_stage_2__1581_, data_stage_2__1580_, data_stage_2__1579_, data_stage_2__1578_, data_stage_2__1577_, data_stage_2__1576_, data_stage_2__1575_, data_stage_2__1574_, data_stage_2__1573_, data_stage_2__1572_, data_stage_2__1571_, data_stage_2__1570_, data_stage_2__1569_, data_stage_2__1568_, data_stage_2__1567_, data_stage_2__1566_, data_stage_2__1565_, data_stage_2__1564_, data_stage_2__1563_, data_stage_2__1562_, data_stage_2__1561_, data_stage_2__1560_, data_stage_2__1559_, data_stage_2__1558_, data_stage_2__1557_, data_stage_2__1556_, data_stage_2__1555_, data_stage_2__1554_, data_stage_2__1553_, data_stage_2__1552_, data_stage_2__1551_, data_stage_2__1550_, data_stage_2__1549_, data_stage_2__1548_, data_stage_2__1547_, data_stage_2__1546_, data_stage_2__1545_, data_stage_2__1544_, data_stage_2__1543_, data_stage_2__1542_, data_stage_2__1541_, data_stage_2__1540_, data_stage_2__1539_, data_stage_2__1538_, data_stage_2__1537_, data_stage_2__1536_, data_stage_2__1535_, data_stage_2__1534_, data_stage_2__1533_, data_stage_2__1532_, data_stage_2__1531_, data_stage_2__1530_, data_stage_2__1529_, data_stage_2__1528_, data_stage_2__1527_, data_stage_2__1526_, data_stage_2__1525_, data_stage_2__1524_, data_stage_2__1523_, data_stage_2__1522_, data_stage_2__1521_, data_stage_2__1520_, data_stage_2__1519_, data_stage_2__1518_, data_stage_2__1517_, data_stage_2__1516_, data_stage_2__1515_, data_stage_2__1514_, data_stage_2__1513_, data_stage_2__1512_, data_stage_2__1511_, data_stage_2__1510_, data_stage_2__1509_, data_stage_2__1508_, data_stage_2__1507_, data_stage_2__1506_, data_stage_2__1505_, data_stage_2__1504_, data_stage_2__1503_, data_stage_2__1502_, data_stage_2__1501_, data_stage_2__1500_, data_stage_2__1499_, data_stage_2__1498_, data_stage_2__1497_, data_stage_2__1496_, data_stage_2__1495_, data_stage_2__1494_, data_stage_2__1493_, data_stage_2__1492_, data_stage_2__1491_, data_stage_2__1490_, data_stage_2__1489_, data_stage_2__1488_, data_stage_2__1487_, data_stage_2__1486_, data_stage_2__1485_, data_stage_2__1484_, data_stage_2__1483_, data_stage_2__1482_, data_stage_2__1481_, data_stage_2__1480_, data_stage_2__1479_, data_stage_2__1478_, data_stage_2__1477_, data_stage_2__1476_, data_stage_2__1475_, data_stage_2__1474_, data_stage_2__1473_, data_stage_2__1472_, data_stage_2__1471_, data_stage_2__1470_, data_stage_2__1469_, data_stage_2__1468_, data_stage_2__1467_, data_stage_2__1466_, data_stage_2__1465_, data_stage_2__1464_, data_stage_2__1463_, data_stage_2__1462_, data_stage_2__1461_, data_stage_2__1460_, data_stage_2__1459_, data_stage_2__1458_, data_stage_2__1457_, data_stage_2__1456_, data_stage_2__1455_, data_stage_2__1454_, data_stage_2__1453_, data_stage_2__1452_, data_stage_2__1451_, data_stage_2__1450_, data_stage_2__1449_, data_stage_2__1448_, data_stage_2__1447_, data_stage_2__1446_, data_stage_2__1445_, data_stage_2__1444_, data_stage_2__1443_, data_stage_2__1442_, data_stage_2__1441_, data_stage_2__1440_, data_stage_2__1439_, data_stage_2__1438_, data_stage_2__1437_, data_stage_2__1436_, data_stage_2__1435_, data_stage_2__1434_, data_stage_2__1433_, data_stage_2__1432_, data_stage_2__1431_, data_stage_2__1430_, data_stage_2__1429_, data_stage_2__1428_, data_stage_2__1427_, data_stage_2__1426_, data_stage_2__1425_, data_stage_2__1424_, data_stage_2__1423_, data_stage_2__1422_, data_stage_2__1421_, data_stage_2__1420_, data_stage_2__1419_, data_stage_2__1418_, data_stage_2__1417_, data_stage_2__1416_, data_stage_2__1415_, data_stage_2__1414_, data_stage_2__1413_, data_stage_2__1412_, data_stage_2__1411_, data_stage_2__1410_, data_stage_2__1409_, data_stage_2__1408_, data_stage_2__1407_, data_stage_2__1406_, data_stage_2__1405_, data_stage_2__1404_, data_stage_2__1403_, data_stage_2__1402_, data_stage_2__1401_, data_stage_2__1400_, data_stage_2__1399_, data_stage_2__1398_, data_stage_2__1397_, data_stage_2__1396_, data_stage_2__1395_, data_stage_2__1394_, data_stage_2__1393_, data_stage_2__1392_, data_stage_2__1391_, data_stage_2__1390_, data_stage_2__1389_, data_stage_2__1388_, data_stage_2__1387_, data_stage_2__1386_, data_stage_2__1385_, data_stage_2__1384_, data_stage_2__1383_, data_stage_2__1382_, data_stage_2__1381_, data_stage_2__1380_, data_stage_2__1379_, data_stage_2__1378_, data_stage_2__1377_, data_stage_2__1376_, data_stage_2__1375_, data_stage_2__1374_, data_stage_2__1373_, data_stage_2__1372_, data_stage_2__1371_, data_stage_2__1370_, data_stage_2__1369_, data_stage_2__1368_, data_stage_2__1367_, data_stage_2__1366_, data_stage_2__1365_, data_stage_2__1364_, data_stage_2__1363_, data_stage_2__1362_, data_stage_2__1361_, data_stage_2__1360_, data_stage_2__1359_, data_stage_2__1358_, data_stage_2__1357_, data_stage_2__1356_, data_stage_2__1355_, data_stage_2__1354_, data_stage_2__1353_, data_stage_2__1352_, data_stage_2__1351_, data_stage_2__1350_, data_stage_2__1349_, data_stage_2__1348_, data_stage_2__1347_, data_stage_2__1346_, data_stage_2__1345_, data_stage_2__1344_, data_stage_2__1343_, data_stage_2__1342_, data_stage_2__1341_, data_stage_2__1340_, data_stage_2__1339_, data_stage_2__1338_, data_stage_2__1337_, data_stage_2__1336_, data_stage_2__1335_, data_stage_2__1334_, data_stage_2__1333_, data_stage_2__1332_, data_stage_2__1331_, data_stage_2__1330_, data_stage_2__1329_, data_stage_2__1328_, data_stage_2__1327_, data_stage_2__1326_, data_stage_2__1325_, data_stage_2__1324_, data_stage_2__1323_, data_stage_2__1322_, data_stage_2__1321_, data_stage_2__1320_, data_stage_2__1319_, data_stage_2__1318_, data_stage_2__1317_, data_stage_2__1316_, data_stage_2__1315_, data_stage_2__1314_, data_stage_2__1313_, data_stage_2__1312_, data_stage_2__1311_, data_stage_2__1310_, data_stage_2__1309_, data_stage_2__1308_, data_stage_2__1307_, data_stage_2__1306_, data_stage_2__1305_, data_stage_2__1304_, data_stage_2__1303_, data_stage_2__1302_, data_stage_2__1301_, data_stage_2__1300_, data_stage_2__1299_, data_stage_2__1298_, data_stage_2__1297_, data_stage_2__1296_, data_stage_2__1295_, data_stage_2__1294_, data_stage_2__1293_, data_stage_2__1292_, data_stage_2__1291_, data_stage_2__1290_, data_stage_2__1289_, data_stage_2__1288_, data_stage_2__1287_, data_stage_2__1286_, data_stage_2__1285_, data_stage_2__1284_, data_stage_2__1283_, data_stage_2__1282_, data_stage_2__1281_, data_stage_2__1280_, data_stage_2__1279_, data_stage_2__1278_, data_stage_2__1277_, data_stage_2__1276_, data_stage_2__1275_, data_stage_2__1274_, data_stage_2__1273_, data_stage_2__1272_, data_stage_2__1271_, data_stage_2__1270_, data_stage_2__1269_, data_stage_2__1268_, data_stage_2__1267_, data_stage_2__1266_, data_stage_2__1265_, data_stage_2__1264_, data_stage_2__1263_, data_stage_2__1262_, data_stage_2__1261_, data_stage_2__1260_, data_stage_2__1259_, data_stage_2__1258_, data_stage_2__1257_, data_stage_2__1256_, data_stage_2__1255_, data_stage_2__1254_, data_stage_2__1253_, data_stage_2__1252_, data_stage_2__1251_, data_stage_2__1250_, data_stage_2__1249_, data_stage_2__1248_, data_stage_2__1247_, data_stage_2__1246_, data_stage_2__1245_, data_stage_2__1244_, data_stage_2__1243_, data_stage_2__1242_, data_stage_2__1241_, data_stage_2__1240_, data_stage_2__1239_, data_stage_2__1238_, data_stage_2__1237_, data_stage_2__1236_, data_stage_2__1235_, data_stage_2__1234_, data_stage_2__1233_, data_stage_2__1232_, data_stage_2__1231_, data_stage_2__1230_, data_stage_2__1229_, data_stage_2__1228_, data_stage_2__1227_, data_stage_2__1226_, data_stage_2__1225_, data_stage_2__1224_, data_stage_2__1223_, data_stage_2__1222_, data_stage_2__1221_, data_stage_2__1220_, data_stage_2__1219_, data_stage_2__1218_, data_stage_2__1217_, data_stage_2__1216_, data_stage_2__1215_, data_stage_2__1214_, data_stage_2__1213_, data_stage_2__1212_, data_stage_2__1211_, data_stage_2__1210_, data_stage_2__1209_, data_stage_2__1208_, data_stage_2__1207_, data_stage_2__1206_, data_stage_2__1205_, data_stage_2__1204_, data_stage_2__1203_, data_stage_2__1202_, data_stage_2__1201_, data_stage_2__1200_, data_stage_2__1199_, data_stage_2__1198_, data_stage_2__1197_, data_stage_2__1196_, data_stage_2__1195_, data_stage_2__1194_, data_stage_2__1193_, data_stage_2__1192_, data_stage_2__1191_, data_stage_2__1190_, data_stage_2__1189_, data_stage_2__1188_, data_stage_2__1187_, data_stage_2__1186_, data_stage_2__1185_, data_stage_2__1184_, data_stage_2__1183_, data_stage_2__1182_, data_stage_2__1181_, data_stage_2__1180_, data_stage_2__1179_, data_stage_2__1178_, data_stage_2__1177_, data_stage_2__1176_, data_stage_2__1175_, data_stage_2__1174_, data_stage_2__1173_, data_stage_2__1172_, data_stage_2__1171_, data_stage_2__1170_, data_stage_2__1169_, data_stage_2__1168_, data_stage_2__1167_, data_stage_2__1166_, data_stage_2__1165_, data_stage_2__1164_, data_stage_2__1163_, data_stage_2__1162_, data_stage_2__1161_, data_stage_2__1160_, data_stage_2__1159_, data_stage_2__1158_, data_stage_2__1157_, data_stage_2__1156_, data_stage_2__1155_, data_stage_2__1154_, data_stage_2__1153_, data_stage_2__1152_, data_stage_2__1151_, data_stage_2__1150_, data_stage_2__1149_, data_stage_2__1148_, data_stage_2__1147_, data_stage_2__1146_, data_stage_2__1145_, data_stage_2__1144_, data_stage_2__1143_, data_stage_2__1142_, data_stage_2__1141_, data_stage_2__1140_, data_stage_2__1139_, data_stage_2__1138_, data_stage_2__1137_, data_stage_2__1136_, data_stage_2__1135_, data_stage_2__1134_, data_stage_2__1133_, data_stage_2__1132_, data_stage_2__1131_, data_stage_2__1130_, data_stage_2__1129_, data_stage_2__1128_, data_stage_2__1127_, data_stage_2__1126_, data_stage_2__1125_, data_stage_2__1124_, data_stage_2__1123_, data_stage_2__1122_, data_stage_2__1121_, data_stage_2__1120_, data_stage_2__1119_, data_stage_2__1118_, data_stage_2__1117_, data_stage_2__1116_, data_stage_2__1115_, data_stage_2__1114_, data_stage_2__1113_, data_stage_2__1112_, data_stage_2__1111_, data_stage_2__1110_, data_stage_2__1109_, data_stage_2__1108_, data_stage_2__1107_, data_stage_2__1106_, data_stage_2__1105_, data_stage_2__1104_, data_stage_2__1103_, data_stage_2__1102_, data_stage_2__1101_, data_stage_2__1100_, data_stage_2__1099_, data_stage_2__1098_, data_stage_2__1097_, data_stage_2__1096_, data_stage_2__1095_, data_stage_2__1094_, data_stage_2__1093_, data_stage_2__1092_, data_stage_2__1091_, data_stage_2__1090_, data_stage_2__1089_, data_stage_2__1088_, data_stage_2__1087_, data_stage_2__1086_, data_stage_2__1085_, data_stage_2__1084_, data_stage_2__1083_, data_stage_2__1082_, data_stage_2__1081_, data_stage_2__1080_, data_stage_2__1079_, data_stage_2__1078_, data_stage_2__1077_, data_stage_2__1076_, data_stage_2__1075_, data_stage_2__1074_, data_stage_2__1073_, data_stage_2__1072_, data_stage_2__1071_, data_stage_2__1070_, data_stage_2__1069_, data_stage_2__1068_, data_stage_2__1067_, data_stage_2__1066_, data_stage_2__1065_, data_stage_2__1064_, data_stage_2__1063_, data_stage_2__1062_, data_stage_2__1061_, data_stage_2__1060_, data_stage_2__1059_, data_stage_2__1058_, data_stage_2__1057_, data_stage_2__1056_, data_stage_2__1055_, data_stage_2__1054_, data_stage_2__1053_, data_stage_2__1052_, data_stage_2__1051_, data_stage_2__1050_, data_stage_2__1049_, data_stage_2__1048_, data_stage_2__1047_, data_stage_2__1046_, data_stage_2__1045_, data_stage_2__1044_, data_stage_2__1043_, data_stage_2__1042_, data_stage_2__1041_, data_stage_2__1040_, data_stage_2__1039_, data_stage_2__1038_, data_stage_2__1037_, data_stage_2__1036_, data_stage_2__1035_, data_stage_2__1034_, data_stage_2__1033_, data_stage_2__1032_, data_stage_2__1031_, data_stage_2__1030_, data_stage_2__1029_, data_stage_2__1028_, data_stage_2__1027_, data_stage_2__1026_, data_stage_2__1025_, data_stage_2__1024_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__2047_, data_stage_3__2046_, data_stage_3__2045_, data_stage_3__2044_, data_stage_3__2043_, data_stage_3__2042_, data_stage_3__2041_, data_stage_3__2040_, data_stage_3__2039_, data_stage_3__2038_, data_stage_3__2037_, data_stage_3__2036_, data_stage_3__2035_, data_stage_3__2034_, data_stage_3__2033_, data_stage_3__2032_, data_stage_3__2031_, data_stage_3__2030_, data_stage_3__2029_, data_stage_3__2028_, data_stage_3__2027_, data_stage_3__2026_, data_stage_3__2025_, data_stage_3__2024_, data_stage_3__2023_, data_stage_3__2022_, data_stage_3__2021_, data_stage_3__2020_, data_stage_3__2019_, data_stage_3__2018_, data_stage_3__2017_, data_stage_3__2016_, data_stage_3__2015_, data_stage_3__2014_, data_stage_3__2013_, data_stage_3__2012_, data_stage_3__2011_, data_stage_3__2010_, data_stage_3__2009_, data_stage_3__2008_, data_stage_3__2007_, data_stage_3__2006_, data_stage_3__2005_, data_stage_3__2004_, data_stage_3__2003_, data_stage_3__2002_, data_stage_3__2001_, data_stage_3__2000_, data_stage_3__1999_, data_stage_3__1998_, data_stage_3__1997_, data_stage_3__1996_, data_stage_3__1995_, data_stage_3__1994_, data_stage_3__1993_, data_stage_3__1992_, data_stage_3__1991_, data_stage_3__1990_, data_stage_3__1989_, data_stage_3__1988_, data_stage_3__1987_, data_stage_3__1986_, data_stage_3__1985_, data_stage_3__1984_, data_stage_3__1983_, data_stage_3__1982_, data_stage_3__1981_, data_stage_3__1980_, data_stage_3__1979_, data_stage_3__1978_, data_stage_3__1977_, data_stage_3__1976_, data_stage_3__1975_, data_stage_3__1974_, data_stage_3__1973_, data_stage_3__1972_, data_stage_3__1971_, data_stage_3__1970_, data_stage_3__1969_, data_stage_3__1968_, data_stage_3__1967_, data_stage_3__1966_, data_stage_3__1965_, data_stage_3__1964_, data_stage_3__1963_, data_stage_3__1962_, data_stage_3__1961_, data_stage_3__1960_, data_stage_3__1959_, data_stage_3__1958_, data_stage_3__1957_, data_stage_3__1956_, data_stage_3__1955_, data_stage_3__1954_, data_stage_3__1953_, data_stage_3__1952_, data_stage_3__1951_, data_stage_3__1950_, data_stage_3__1949_, data_stage_3__1948_, data_stage_3__1947_, data_stage_3__1946_, data_stage_3__1945_, data_stage_3__1944_, data_stage_3__1943_, data_stage_3__1942_, data_stage_3__1941_, data_stage_3__1940_, data_stage_3__1939_, data_stage_3__1938_, data_stage_3__1937_, data_stage_3__1936_, data_stage_3__1935_, data_stage_3__1934_, data_stage_3__1933_, data_stage_3__1932_, data_stage_3__1931_, data_stage_3__1930_, data_stage_3__1929_, data_stage_3__1928_, data_stage_3__1927_, data_stage_3__1926_, data_stage_3__1925_, data_stage_3__1924_, data_stage_3__1923_, data_stage_3__1922_, data_stage_3__1921_, data_stage_3__1920_, data_stage_3__1919_, data_stage_3__1918_, data_stage_3__1917_, data_stage_3__1916_, data_stage_3__1915_, data_stage_3__1914_, data_stage_3__1913_, data_stage_3__1912_, data_stage_3__1911_, data_stage_3__1910_, data_stage_3__1909_, data_stage_3__1908_, data_stage_3__1907_, data_stage_3__1906_, data_stage_3__1905_, data_stage_3__1904_, data_stage_3__1903_, data_stage_3__1902_, data_stage_3__1901_, data_stage_3__1900_, data_stage_3__1899_, data_stage_3__1898_, data_stage_3__1897_, data_stage_3__1896_, data_stage_3__1895_, data_stage_3__1894_, data_stage_3__1893_, data_stage_3__1892_, data_stage_3__1891_, data_stage_3__1890_, data_stage_3__1889_, data_stage_3__1888_, data_stage_3__1887_, data_stage_3__1886_, data_stage_3__1885_, data_stage_3__1884_, data_stage_3__1883_, data_stage_3__1882_, data_stage_3__1881_, data_stage_3__1880_, data_stage_3__1879_, data_stage_3__1878_, data_stage_3__1877_, data_stage_3__1876_, data_stage_3__1875_, data_stage_3__1874_, data_stage_3__1873_, data_stage_3__1872_, data_stage_3__1871_, data_stage_3__1870_, data_stage_3__1869_, data_stage_3__1868_, data_stage_3__1867_, data_stage_3__1866_, data_stage_3__1865_, data_stage_3__1864_, data_stage_3__1863_, data_stage_3__1862_, data_stage_3__1861_, data_stage_3__1860_, data_stage_3__1859_, data_stage_3__1858_, data_stage_3__1857_, data_stage_3__1856_, data_stage_3__1855_, data_stage_3__1854_, data_stage_3__1853_, data_stage_3__1852_, data_stage_3__1851_, data_stage_3__1850_, data_stage_3__1849_, data_stage_3__1848_, data_stage_3__1847_, data_stage_3__1846_, data_stage_3__1845_, data_stage_3__1844_, data_stage_3__1843_, data_stage_3__1842_, data_stage_3__1841_, data_stage_3__1840_, data_stage_3__1839_, data_stage_3__1838_, data_stage_3__1837_, data_stage_3__1836_, data_stage_3__1835_, data_stage_3__1834_, data_stage_3__1833_, data_stage_3__1832_, data_stage_3__1831_, data_stage_3__1830_, data_stage_3__1829_, data_stage_3__1828_, data_stage_3__1827_, data_stage_3__1826_, data_stage_3__1825_, data_stage_3__1824_, data_stage_3__1823_, data_stage_3__1822_, data_stage_3__1821_, data_stage_3__1820_, data_stage_3__1819_, data_stage_3__1818_, data_stage_3__1817_, data_stage_3__1816_, data_stage_3__1815_, data_stage_3__1814_, data_stage_3__1813_, data_stage_3__1812_, data_stage_3__1811_, data_stage_3__1810_, data_stage_3__1809_, data_stage_3__1808_, data_stage_3__1807_, data_stage_3__1806_, data_stage_3__1805_, data_stage_3__1804_, data_stage_3__1803_, data_stage_3__1802_, data_stage_3__1801_, data_stage_3__1800_, data_stage_3__1799_, data_stage_3__1798_, data_stage_3__1797_, data_stage_3__1796_, data_stage_3__1795_, data_stage_3__1794_, data_stage_3__1793_, data_stage_3__1792_, data_stage_3__1791_, data_stage_3__1790_, data_stage_3__1789_, data_stage_3__1788_, data_stage_3__1787_, data_stage_3__1786_, data_stage_3__1785_, data_stage_3__1784_, data_stage_3__1783_, data_stage_3__1782_, data_stage_3__1781_, data_stage_3__1780_, data_stage_3__1779_, data_stage_3__1778_, data_stage_3__1777_, data_stage_3__1776_, data_stage_3__1775_, data_stage_3__1774_, data_stage_3__1773_, data_stage_3__1772_, data_stage_3__1771_, data_stage_3__1770_, data_stage_3__1769_, data_stage_3__1768_, data_stage_3__1767_, data_stage_3__1766_, data_stage_3__1765_, data_stage_3__1764_, data_stage_3__1763_, data_stage_3__1762_, data_stage_3__1761_, data_stage_3__1760_, data_stage_3__1759_, data_stage_3__1758_, data_stage_3__1757_, data_stage_3__1756_, data_stage_3__1755_, data_stage_3__1754_, data_stage_3__1753_, data_stage_3__1752_, data_stage_3__1751_, data_stage_3__1750_, data_stage_3__1749_, data_stage_3__1748_, data_stage_3__1747_, data_stage_3__1746_, data_stage_3__1745_, data_stage_3__1744_, data_stage_3__1743_, data_stage_3__1742_, data_stage_3__1741_, data_stage_3__1740_, data_stage_3__1739_, data_stage_3__1738_, data_stage_3__1737_, data_stage_3__1736_, data_stage_3__1735_, data_stage_3__1734_, data_stage_3__1733_, data_stage_3__1732_, data_stage_3__1731_, data_stage_3__1730_, data_stage_3__1729_, data_stage_3__1728_, data_stage_3__1727_, data_stage_3__1726_, data_stage_3__1725_, data_stage_3__1724_, data_stage_3__1723_, data_stage_3__1722_, data_stage_3__1721_, data_stage_3__1720_, data_stage_3__1719_, data_stage_3__1718_, data_stage_3__1717_, data_stage_3__1716_, data_stage_3__1715_, data_stage_3__1714_, data_stage_3__1713_, data_stage_3__1712_, data_stage_3__1711_, data_stage_3__1710_, data_stage_3__1709_, data_stage_3__1708_, data_stage_3__1707_, data_stage_3__1706_, data_stage_3__1705_, data_stage_3__1704_, data_stage_3__1703_, data_stage_3__1702_, data_stage_3__1701_, data_stage_3__1700_, data_stage_3__1699_, data_stage_3__1698_, data_stage_3__1697_, data_stage_3__1696_, data_stage_3__1695_, data_stage_3__1694_, data_stage_3__1693_, data_stage_3__1692_, data_stage_3__1691_, data_stage_3__1690_, data_stage_3__1689_, data_stage_3__1688_, data_stage_3__1687_, data_stage_3__1686_, data_stage_3__1685_, data_stage_3__1684_, data_stage_3__1683_, data_stage_3__1682_, data_stage_3__1681_, data_stage_3__1680_, data_stage_3__1679_, data_stage_3__1678_, data_stage_3__1677_, data_stage_3__1676_, data_stage_3__1675_, data_stage_3__1674_, data_stage_3__1673_, data_stage_3__1672_, data_stage_3__1671_, data_stage_3__1670_, data_stage_3__1669_, data_stage_3__1668_, data_stage_3__1667_, data_stage_3__1666_, data_stage_3__1665_, data_stage_3__1664_, data_stage_3__1663_, data_stage_3__1662_, data_stage_3__1661_, data_stage_3__1660_, data_stage_3__1659_, data_stage_3__1658_, data_stage_3__1657_, data_stage_3__1656_, data_stage_3__1655_, data_stage_3__1654_, data_stage_3__1653_, data_stage_3__1652_, data_stage_3__1651_, data_stage_3__1650_, data_stage_3__1649_, data_stage_3__1648_, data_stage_3__1647_, data_stage_3__1646_, data_stage_3__1645_, data_stage_3__1644_, data_stage_3__1643_, data_stage_3__1642_, data_stage_3__1641_, data_stage_3__1640_, data_stage_3__1639_, data_stage_3__1638_, data_stage_3__1637_, data_stage_3__1636_, data_stage_3__1635_, data_stage_3__1634_, data_stage_3__1633_, data_stage_3__1632_, data_stage_3__1631_, data_stage_3__1630_, data_stage_3__1629_, data_stage_3__1628_, data_stage_3__1627_, data_stage_3__1626_, data_stage_3__1625_, data_stage_3__1624_, data_stage_3__1623_, data_stage_3__1622_, data_stage_3__1621_, data_stage_3__1620_, data_stage_3__1619_, data_stage_3__1618_, data_stage_3__1617_, data_stage_3__1616_, data_stage_3__1615_, data_stage_3__1614_, data_stage_3__1613_, data_stage_3__1612_, data_stage_3__1611_, data_stage_3__1610_, data_stage_3__1609_, data_stage_3__1608_, data_stage_3__1607_, data_stage_3__1606_, data_stage_3__1605_, data_stage_3__1604_, data_stage_3__1603_, data_stage_3__1602_, data_stage_3__1601_, data_stage_3__1600_, data_stage_3__1599_, data_stage_3__1598_, data_stage_3__1597_, data_stage_3__1596_, data_stage_3__1595_, data_stage_3__1594_, data_stage_3__1593_, data_stage_3__1592_, data_stage_3__1591_, data_stage_3__1590_, data_stage_3__1589_, data_stage_3__1588_, data_stage_3__1587_, data_stage_3__1586_, data_stage_3__1585_, data_stage_3__1584_, data_stage_3__1583_, data_stage_3__1582_, data_stage_3__1581_, data_stage_3__1580_, data_stage_3__1579_, data_stage_3__1578_, data_stage_3__1577_, data_stage_3__1576_, data_stage_3__1575_, data_stage_3__1574_, data_stage_3__1573_, data_stage_3__1572_, data_stage_3__1571_, data_stage_3__1570_, data_stage_3__1569_, data_stage_3__1568_, data_stage_3__1567_, data_stage_3__1566_, data_stage_3__1565_, data_stage_3__1564_, data_stage_3__1563_, data_stage_3__1562_, data_stage_3__1561_, data_stage_3__1560_, data_stage_3__1559_, data_stage_3__1558_, data_stage_3__1557_, data_stage_3__1556_, data_stage_3__1555_, data_stage_3__1554_, data_stage_3__1553_, data_stage_3__1552_, data_stage_3__1551_, data_stage_3__1550_, data_stage_3__1549_, data_stage_3__1548_, data_stage_3__1547_, data_stage_3__1546_, data_stage_3__1545_, data_stage_3__1544_, data_stage_3__1543_, data_stage_3__1542_, data_stage_3__1541_, data_stage_3__1540_, data_stage_3__1539_, data_stage_3__1538_, data_stage_3__1537_, data_stage_3__1536_, data_stage_3__1535_, data_stage_3__1534_, data_stage_3__1533_, data_stage_3__1532_, data_stage_3__1531_, data_stage_3__1530_, data_stage_3__1529_, data_stage_3__1528_, data_stage_3__1527_, data_stage_3__1526_, data_stage_3__1525_, data_stage_3__1524_, data_stage_3__1523_, data_stage_3__1522_, data_stage_3__1521_, data_stage_3__1520_, data_stage_3__1519_, data_stage_3__1518_, data_stage_3__1517_, data_stage_3__1516_, data_stage_3__1515_, data_stage_3__1514_, data_stage_3__1513_, data_stage_3__1512_, data_stage_3__1511_, data_stage_3__1510_, data_stage_3__1509_, data_stage_3__1508_, data_stage_3__1507_, data_stage_3__1506_, data_stage_3__1505_, data_stage_3__1504_, data_stage_3__1503_, data_stage_3__1502_, data_stage_3__1501_, data_stage_3__1500_, data_stage_3__1499_, data_stage_3__1498_, data_stage_3__1497_, data_stage_3__1496_, data_stage_3__1495_, data_stage_3__1494_, data_stage_3__1493_, data_stage_3__1492_, data_stage_3__1491_, data_stage_3__1490_, data_stage_3__1489_, data_stage_3__1488_, data_stage_3__1487_, data_stage_3__1486_, data_stage_3__1485_, data_stage_3__1484_, data_stage_3__1483_, data_stage_3__1482_, data_stage_3__1481_, data_stage_3__1480_, data_stage_3__1479_, data_stage_3__1478_, data_stage_3__1477_, data_stage_3__1476_, data_stage_3__1475_, data_stage_3__1474_, data_stage_3__1473_, data_stage_3__1472_, data_stage_3__1471_, data_stage_3__1470_, data_stage_3__1469_, data_stage_3__1468_, data_stage_3__1467_, data_stage_3__1466_, data_stage_3__1465_, data_stage_3__1464_, data_stage_3__1463_, data_stage_3__1462_, data_stage_3__1461_, data_stage_3__1460_, data_stage_3__1459_, data_stage_3__1458_, data_stage_3__1457_, data_stage_3__1456_, data_stage_3__1455_, data_stage_3__1454_, data_stage_3__1453_, data_stage_3__1452_, data_stage_3__1451_, data_stage_3__1450_, data_stage_3__1449_, data_stage_3__1448_, data_stage_3__1447_, data_stage_3__1446_, data_stage_3__1445_, data_stage_3__1444_, data_stage_3__1443_, data_stage_3__1442_, data_stage_3__1441_, data_stage_3__1440_, data_stage_3__1439_, data_stage_3__1438_, data_stage_3__1437_, data_stage_3__1436_, data_stage_3__1435_, data_stage_3__1434_, data_stage_3__1433_, data_stage_3__1432_, data_stage_3__1431_, data_stage_3__1430_, data_stage_3__1429_, data_stage_3__1428_, data_stage_3__1427_, data_stage_3__1426_, data_stage_3__1425_, data_stage_3__1424_, data_stage_3__1423_, data_stage_3__1422_, data_stage_3__1421_, data_stage_3__1420_, data_stage_3__1419_, data_stage_3__1418_, data_stage_3__1417_, data_stage_3__1416_, data_stage_3__1415_, data_stage_3__1414_, data_stage_3__1413_, data_stage_3__1412_, data_stage_3__1411_, data_stage_3__1410_, data_stage_3__1409_, data_stage_3__1408_, data_stage_3__1407_, data_stage_3__1406_, data_stage_3__1405_, data_stage_3__1404_, data_stage_3__1403_, data_stage_3__1402_, data_stage_3__1401_, data_stage_3__1400_, data_stage_3__1399_, data_stage_3__1398_, data_stage_3__1397_, data_stage_3__1396_, data_stage_3__1395_, data_stage_3__1394_, data_stage_3__1393_, data_stage_3__1392_, data_stage_3__1391_, data_stage_3__1390_, data_stage_3__1389_, data_stage_3__1388_, data_stage_3__1387_, data_stage_3__1386_, data_stage_3__1385_, data_stage_3__1384_, data_stage_3__1383_, data_stage_3__1382_, data_stage_3__1381_, data_stage_3__1380_, data_stage_3__1379_, data_stage_3__1378_, data_stage_3__1377_, data_stage_3__1376_, data_stage_3__1375_, data_stage_3__1374_, data_stage_3__1373_, data_stage_3__1372_, data_stage_3__1371_, data_stage_3__1370_, data_stage_3__1369_, data_stage_3__1368_, data_stage_3__1367_, data_stage_3__1366_, data_stage_3__1365_, data_stage_3__1364_, data_stage_3__1363_, data_stage_3__1362_, data_stage_3__1361_, data_stage_3__1360_, data_stage_3__1359_, data_stage_3__1358_, data_stage_3__1357_, data_stage_3__1356_, data_stage_3__1355_, data_stage_3__1354_, data_stage_3__1353_, data_stage_3__1352_, data_stage_3__1351_, data_stage_3__1350_, data_stage_3__1349_, data_stage_3__1348_, data_stage_3__1347_, data_stage_3__1346_, data_stage_3__1345_, data_stage_3__1344_, data_stage_3__1343_, data_stage_3__1342_, data_stage_3__1341_, data_stage_3__1340_, data_stage_3__1339_, data_stage_3__1338_, data_stage_3__1337_, data_stage_3__1336_, data_stage_3__1335_, data_stage_3__1334_, data_stage_3__1333_, data_stage_3__1332_, data_stage_3__1331_, data_stage_3__1330_, data_stage_3__1329_, data_stage_3__1328_, data_stage_3__1327_, data_stage_3__1326_, data_stage_3__1325_, data_stage_3__1324_, data_stage_3__1323_, data_stage_3__1322_, data_stage_3__1321_, data_stage_3__1320_, data_stage_3__1319_, data_stage_3__1318_, data_stage_3__1317_, data_stage_3__1316_, data_stage_3__1315_, data_stage_3__1314_, data_stage_3__1313_, data_stage_3__1312_, data_stage_3__1311_, data_stage_3__1310_, data_stage_3__1309_, data_stage_3__1308_, data_stage_3__1307_, data_stage_3__1306_, data_stage_3__1305_, data_stage_3__1304_, data_stage_3__1303_, data_stage_3__1302_, data_stage_3__1301_, data_stage_3__1300_, data_stage_3__1299_, data_stage_3__1298_, data_stage_3__1297_, data_stage_3__1296_, data_stage_3__1295_, data_stage_3__1294_, data_stage_3__1293_, data_stage_3__1292_, data_stage_3__1291_, data_stage_3__1290_, data_stage_3__1289_, data_stage_3__1288_, data_stage_3__1287_, data_stage_3__1286_, data_stage_3__1285_, data_stage_3__1284_, data_stage_3__1283_, data_stage_3__1282_, data_stage_3__1281_, data_stage_3__1280_, data_stage_3__1279_, data_stage_3__1278_, data_stage_3__1277_, data_stage_3__1276_, data_stage_3__1275_, data_stage_3__1274_, data_stage_3__1273_, data_stage_3__1272_, data_stage_3__1271_, data_stage_3__1270_, data_stage_3__1269_, data_stage_3__1268_, data_stage_3__1267_, data_stage_3__1266_, data_stage_3__1265_, data_stage_3__1264_, data_stage_3__1263_, data_stage_3__1262_, data_stage_3__1261_, data_stage_3__1260_, data_stage_3__1259_, data_stage_3__1258_, data_stage_3__1257_, data_stage_3__1256_, data_stage_3__1255_, data_stage_3__1254_, data_stage_3__1253_, data_stage_3__1252_, data_stage_3__1251_, data_stage_3__1250_, data_stage_3__1249_, data_stage_3__1248_, data_stage_3__1247_, data_stage_3__1246_, data_stage_3__1245_, data_stage_3__1244_, data_stage_3__1243_, data_stage_3__1242_, data_stage_3__1241_, data_stage_3__1240_, data_stage_3__1239_, data_stage_3__1238_, data_stage_3__1237_, data_stage_3__1236_, data_stage_3__1235_, data_stage_3__1234_, data_stage_3__1233_, data_stage_3__1232_, data_stage_3__1231_, data_stage_3__1230_, data_stage_3__1229_, data_stage_3__1228_, data_stage_3__1227_, data_stage_3__1226_, data_stage_3__1225_, data_stage_3__1224_, data_stage_3__1223_, data_stage_3__1222_, data_stage_3__1221_, data_stage_3__1220_, data_stage_3__1219_, data_stage_3__1218_, data_stage_3__1217_, data_stage_3__1216_, data_stage_3__1215_, data_stage_3__1214_, data_stage_3__1213_, data_stage_3__1212_, data_stage_3__1211_, data_stage_3__1210_, data_stage_3__1209_, data_stage_3__1208_, data_stage_3__1207_, data_stage_3__1206_, data_stage_3__1205_, data_stage_3__1204_, data_stage_3__1203_, data_stage_3__1202_, data_stage_3__1201_, data_stage_3__1200_, data_stage_3__1199_, data_stage_3__1198_, data_stage_3__1197_, data_stage_3__1196_, data_stage_3__1195_, data_stage_3__1194_, data_stage_3__1193_, data_stage_3__1192_, data_stage_3__1191_, data_stage_3__1190_, data_stage_3__1189_, data_stage_3__1188_, data_stage_3__1187_, data_stage_3__1186_, data_stage_3__1185_, data_stage_3__1184_, data_stage_3__1183_, data_stage_3__1182_, data_stage_3__1181_, data_stage_3__1180_, data_stage_3__1179_, data_stage_3__1178_, data_stage_3__1177_, data_stage_3__1176_, data_stage_3__1175_, data_stage_3__1174_, data_stage_3__1173_, data_stage_3__1172_, data_stage_3__1171_, data_stage_3__1170_, data_stage_3__1169_, data_stage_3__1168_, data_stage_3__1167_, data_stage_3__1166_, data_stage_3__1165_, data_stage_3__1164_, data_stage_3__1163_, data_stage_3__1162_, data_stage_3__1161_, data_stage_3__1160_, data_stage_3__1159_, data_stage_3__1158_, data_stage_3__1157_, data_stage_3__1156_, data_stage_3__1155_, data_stage_3__1154_, data_stage_3__1153_, data_stage_3__1152_, data_stage_3__1151_, data_stage_3__1150_, data_stage_3__1149_, data_stage_3__1148_, data_stage_3__1147_, data_stage_3__1146_, data_stage_3__1145_, data_stage_3__1144_, data_stage_3__1143_, data_stage_3__1142_, data_stage_3__1141_, data_stage_3__1140_, data_stage_3__1139_, data_stage_3__1138_, data_stage_3__1137_, data_stage_3__1136_, data_stage_3__1135_, data_stage_3__1134_, data_stage_3__1133_, data_stage_3__1132_, data_stage_3__1131_, data_stage_3__1130_, data_stage_3__1129_, data_stage_3__1128_, data_stage_3__1127_, data_stage_3__1126_, data_stage_3__1125_, data_stage_3__1124_, data_stage_3__1123_, data_stage_3__1122_, data_stage_3__1121_, data_stage_3__1120_, data_stage_3__1119_, data_stage_3__1118_, data_stage_3__1117_, data_stage_3__1116_, data_stage_3__1115_, data_stage_3__1114_, data_stage_3__1113_, data_stage_3__1112_, data_stage_3__1111_, data_stage_3__1110_, data_stage_3__1109_, data_stage_3__1108_, data_stage_3__1107_, data_stage_3__1106_, data_stage_3__1105_, data_stage_3__1104_, data_stage_3__1103_, data_stage_3__1102_, data_stage_3__1101_, data_stage_3__1100_, data_stage_3__1099_, data_stage_3__1098_, data_stage_3__1097_, data_stage_3__1096_, data_stage_3__1095_, data_stage_3__1094_, data_stage_3__1093_, data_stage_3__1092_, data_stage_3__1091_, data_stage_3__1090_, data_stage_3__1089_, data_stage_3__1088_, data_stage_3__1087_, data_stage_3__1086_, data_stage_3__1085_, data_stage_3__1084_, data_stage_3__1083_, data_stage_3__1082_, data_stage_3__1081_, data_stage_3__1080_, data_stage_3__1079_, data_stage_3__1078_, data_stage_3__1077_, data_stage_3__1076_, data_stage_3__1075_, data_stage_3__1074_, data_stage_3__1073_, data_stage_3__1072_, data_stage_3__1071_, data_stage_3__1070_, data_stage_3__1069_, data_stage_3__1068_, data_stage_3__1067_, data_stage_3__1066_, data_stage_3__1065_, data_stage_3__1064_, data_stage_3__1063_, data_stage_3__1062_, data_stage_3__1061_, data_stage_3__1060_, data_stage_3__1059_, data_stage_3__1058_, data_stage_3__1057_, data_stage_3__1056_, data_stage_3__1055_, data_stage_3__1054_, data_stage_3__1053_, data_stage_3__1052_, data_stage_3__1051_, data_stage_3__1050_, data_stage_3__1049_, data_stage_3__1048_, data_stage_3__1047_, data_stage_3__1046_, data_stage_3__1045_, data_stage_3__1044_, data_stage_3__1043_, data_stage_3__1042_, data_stage_3__1041_, data_stage_3__1040_, data_stage_3__1039_, data_stage_3__1038_, data_stage_3__1037_, data_stage_3__1036_, data_stage_3__1035_, data_stage_3__1034_, data_stage_3__1033_, data_stage_3__1032_, data_stage_3__1031_, data_stage_3__1030_, data_stage_3__1029_, data_stage_3__1028_, data_stage_3__1027_, data_stage_3__1026_, data_stage_3__1025_, data_stage_3__1024_ })
  );


  bsg_swap_width_p512
  mux_stage_2__mux_swap_2__swap_inst
  (
    .data_i({ data_stage_2__3071_, data_stage_2__3070_, data_stage_2__3069_, data_stage_2__3068_, data_stage_2__3067_, data_stage_2__3066_, data_stage_2__3065_, data_stage_2__3064_, data_stage_2__3063_, data_stage_2__3062_, data_stage_2__3061_, data_stage_2__3060_, data_stage_2__3059_, data_stage_2__3058_, data_stage_2__3057_, data_stage_2__3056_, data_stage_2__3055_, data_stage_2__3054_, data_stage_2__3053_, data_stage_2__3052_, data_stage_2__3051_, data_stage_2__3050_, data_stage_2__3049_, data_stage_2__3048_, data_stage_2__3047_, data_stage_2__3046_, data_stage_2__3045_, data_stage_2__3044_, data_stage_2__3043_, data_stage_2__3042_, data_stage_2__3041_, data_stage_2__3040_, data_stage_2__3039_, data_stage_2__3038_, data_stage_2__3037_, data_stage_2__3036_, data_stage_2__3035_, data_stage_2__3034_, data_stage_2__3033_, data_stage_2__3032_, data_stage_2__3031_, data_stage_2__3030_, data_stage_2__3029_, data_stage_2__3028_, data_stage_2__3027_, data_stage_2__3026_, data_stage_2__3025_, data_stage_2__3024_, data_stage_2__3023_, data_stage_2__3022_, data_stage_2__3021_, data_stage_2__3020_, data_stage_2__3019_, data_stage_2__3018_, data_stage_2__3017_, data_stage_2__3016_, data_stage_2__3015_, data_stage_2__3014_, data_stage_2__3013_, data_stage_2__3012_, data_stage_2__3011_, data_stage_2__3010_, data_stage_2__3009_, data_stage_2__3008_, data_stage_2__3007_, data_stage_2__3006_, data_stage_2__3005_, data_stage_2__3004_, data_stage_2__3003_, data_stage_2__3002_, data_stage_2__3001_, data_stage_2__3000_, data_stage_2__2999_, data_stage_2__2998_, data_stage_2__2997_, data_stage_2__2996_, data_stage_2__2995_, data_stage_2__2994_, data_stage_2__2993_, data_stage_2__2992_, data_stage_2__2991_, data_stage_2__2990_, data_stage_2__2989_, data_stage_2__2988_, data_stage_2__2987_, data_stage_2__2986_, data_stage_2__2985_, data_stage_2__2984_, data_stage_2__2983_, data_stage_2__2982_, data_stage_2__2981_, data_stage_2__2980_, data_stage_2__2979_, data_stage_2__2978_, data_stage_2__2977_, data_stage_2__2976_, data_stage_2__2975_, data_stage_2__2974_, data_stage_2__2973_, data_stage_2__2972_, data_stage_2__2971_, data_stage_2__2970_, data_stage_2__2969_, data_stage_2__2968_, data_stage_2__2967_, data_stage_2__2966_, data_stage_2__2965_, data_stage_2__2964_, data_stage_2__2963_, data_stage_2__2962_, data_stage_2__2961_, data_stage_2__2960_, data_stage_2__2959_, data_stage_2__2958_, data_stage_2__2957_, data_stage_2__2956_, data_stage_2__2955_, data_stage_2__2954_, data_stage_2__2953_, data_stage_2__2952_, data_stage_2__2951_, data_stage_2__2950_, data_stage_2__2949_, data_stage_2__2948_, data_stage_2__2947_, data_stage_2__2946_, data_stage_2__2945_, data_stage_2__2944_, data_stage_2__2943_, data_stage_2__2942_, data_stage_2__2941_, data_stage_2__2940_, data_stage_2__2939_, data_stage_2__2938_, data_stage_2__2937_, data_stage_2__2936_, data_stage_2__2935_, data_stage_2__2934_, data_stage_2__2933_, data_stage_2__2932_, data_stage_2__2931_, data_stage_2__2930_, data_stage_2__2929_, data_stage_2__2928_, data_stage_2__2927_, data_stage_2__2926_, data_stage_2__2925_, data_stage_2__2924_, data_stage_2__2923_, data_stage_2__2922_, data_stage_2__2921_, data_stage_2__2920_, data_stage_2__2919_, data_stage_2__2918_, data_stage_2__2917_, data_stage_2__2916_, data_stage_2__2915_, data_stage_2__2914_, data_stage_2__2913_, data_stage_2__2912_, data_stage_2__2911_, data_stage_2__2910_, data_stage_2__2909_, data_stage_2__2908_, data_stage_2__2907_, data_stage_2__2906_, data_stage_2__2905_, data_stage_2__2904_, data_stage_2__2903_, data_stage_2__2902_, data_stage_2__2901_, data_stage_2__2900_, data_stage_2__2899_, data_stage_2__2898_, data_stage_2__2897_, data_stage_2__2896_, data_stage_2__2895_, data_stage_2__2894_, data_stage_2__2893_, data_stage_2__2892_, data_stage_2__2891_, data_stage_2__2890_, data_stage_2__2889_, data_stage_2__2888_, data_stage_2__2887_, data_stage_2__2886_, data_stage_2__2885_, data_stage_2__2884_, data_stage_2__2883_, data_stage_2__2882_, data_stage_2__2881_, data_stage_2__2880_, data_stage_2__2879_, data_stage_2__2878_, data_stage_2__2877_, data_stage_2__2876_, data_stage_2__2875_, data_stage_2__2874_, data_stage_2__2873_, data_stage_2__2872_, data_stage_2__2871_, data_stage_2__2870_, data_stage_2__2869_, data_stage_2__2868_, data_stage_2__2867_, data_stage_2__2866_, data_stage_2__2865_, data_stage_2__2864_, data_stage_2__2863_, data_stage_2__2862_, data_stage_2__2861_, data_stage_2__2860_, data_stage_2__2859_, data_stage_2__2858_, data_stage_2__2857_, data_stage_2__2856_, data_stage_2__2855_, data_stage_2__2854_, data_stage_2__2853_, data_stage_2__2852_, data_stage_2__2851_, data_stage_2__2850_, data_stage_2__2849_, data_stage_2__2848_, data_stage_2__2847_, data_stage_2__2846_, data_stage_2__2845_, data_stage_2__2844_, data_stage_2__2843_, data_stage_2__2842_, data_stage_2__2841_, data_stage_2__2840_, data_stage_2__2839_, data_stage_2__2838_, data_stage_2__2837_, data_stage_2__2836_, data_stage_2__2835_, data_stage_2__2834_, data_stage_2__2833_, data_stage_2__2832_, data_stage_2__2831_, data_stage_2__2830_, data_stage_2__2829_, data_stage_2__2828_, data_stage_2__2827_, data_stage_2__2826_, data_stage_2__2825_, data_stage_2__2824_, data_stage_2__2823_, data_stage_2__2822_, data_stage_2__2821_, data_stage_2__2820_, data_stage_2__2819_, data_stage_2__2818_, data_stage_2__2817_, data_stage_2__2816_, data_stage_2__2815_, data_stage_2__2814_, data_stage_2__2813_, data_stage_2__2812_, data_stage_2__2811_, data_stage_2__2810_, data_stage_2__2809_, data_stage_2__2808_, data_stage_2__2807_, data_stage_2__2806_, data_stage_2__2805_, data_stage_2__2804_, data_stage_2__2803_, data_stage_2__2802_, data_stage_2__2801_, data_stage_2__2800_, data_stage_2__2799_, data_stage_2__2798_, data_stage_2__2797_, data_stage_2__2796_, data_stage_2__2795_, data_stage_2__2794_, data_stage_2__2793_, data_stage_2__2792_, data_stage_2__2791_, data_stage_2__2790_, data_stage_2__2789_, data_stage_2__2788_, data_stage_2__2787_, data_stage_2__2786_, data_stage_2__2785_, data_stage_2__2784_, data_stage_2__2783_, data_stage_2__2782_, data_stage_2__2781_, data_stage_2__2780_, data_stage_2__2779_, data_stage_2__2778_, data_stage_2__2777_, data_stage_2__2776_, data_stage_2__2775_, data_stage_2__2774_, data_stage_2__2773_, data_stage_2__2772_, data_stage_2__2771_, data_stage_2__2770_, data_stage_2__2769_, data_stage_2__2768_, data_stage_2__2767_, data_stage_2__2766_, data_stage_2__2765_, data_stage_2__2764_, data_stage_2__2763_, data_stage_2__2762_, data_stage_2__2761_, data_stage_2__2760_, data_stage_2__2759_, data_stage_2__2758_, data_stage_2__2757_, data_stage_2__2756_, data_stage_2__2755_, data_stage_2__2754_, data_stage_2__2753_, data_stage_2__2752_, data_stage_2__2751_, data_stage_2__2750_, data_stage_2__2749_, data_stage_2__2748_, data_stage_2__2747_, data_stage_2__2746_, data_stage_2__2745_, data_stage_2__2744_, data_stage_2__2743_, data_stage_2__2742_, data_stage_2__2741_, data_stage_2__2740_, data_stage_2__2739_, data_stage_2__2738_, data_stage_2__2737_, data_stage_2__2736_, data_stage_2__2735_, data_stage_2__2734_, data_stage_2__2733_, data_stage_2__2732_, data_stage_2__2731_, data_stage_2__2730_, data_stage_2__2729_, data_stage_2__2728_, data_stage_2__2727_, data_stage_2__2726_, data_stage_2__2725_, data_stage_2__2724_, data_stage_2__2723_, data_stage_2__2722_, data_stage_2__2721_, data_stage_2__2720_, data_stage_2__2719_, data_stage_2__2718_, data_stage_2__2717_, data_stage_2__2716_, data_stage_2__2715_, data_stage_2__2714_, data_stage_2__2713_, data_stage_2__2712_, data_stage_2__2711_, data_stage_2__2710_, data_stage_2__2709_, data_stage_2__2708_, data_stage_2__2707_, data_stage_2__2706_, data_stage_2__2705_, data_stage_2__2704_, data_stage_2__2703_, data_stage_2__2702_, data_stage_2__2701_, data_stage_2__2700_, data_stage_2__2699_, data_stage_2__2698_, data_stage_2__2697_, data_stage_2__2696_, data_stage_2__2695_, data_stage_2__2694_, data_stage_2__2693_, data_stage_2__2692_, data_stage_2__2691_, data_stage_2__2690_, data_stage_2__2689_, data_stage_2__2688_, data_stage_2__2687_, data_stage_2__2686_, data_stage_2__2685_, data_stage_2__2684_, data_stage_2__2683_, data_stage_2__2682_, data_stage_2__2681_, data_stage_2__2680_, data_stage_2__2679_, data_stage_2__2678_, data_stage_2__2677_, data_stage_2__2676_, data_stage_2__2675_, data_stage_2__2674_, data_stage_2__2673_, data_stage_2__2672_, data_stage_2__2671_, data_stage_2__2670_, data_stage_2__2669_, data_stage_2__2668_, data_stage_2__2667_, data_stage_2__2666_, data_stage_2__2665_, data_stage_2__2664_, data_stage_2__2663_, data_stage_2__2662_, data_stage_2__2661_, data_stage_2__2660_, data_stage_2__2659_, data_stage_2__2658_, data_stage_2__2657_, data_stage_2__2656_, data_stage_2__2655_, data_stage_2__2654_, data_stage_2__2653_, data_stage_2__2652_, data_stage_2__2651_, data_stage_2__2650_, data_stage_2__2649_, data_stage_2__2648_, data_stage_2__2647_, data_stage_2__2646_, data_stage_2__2645_, data_stage_2__2644_, data_stage_2__2643_, data_stage_2__2642_, data_stage_2__2641_, data_stage_2__2640_, data_stage_2__2639_, data_stage_2__2638_, data_stage_2__2637_, data_stage_2__2636_, data_stage_2__2635_, data_stage_2__2634_, data_stage_2__2633_, data_stage_2__2632_, data_stage_2__2631_, data_stage_2__2630_, data_stage_2__2629_, data_stage_2__2628_, data_stage_2__2627_, data_stage_2__2626_, data_stage_2__2625_, data_stage_2__2624_, data_stage_2__2623_, data_stage_2__2622_, data_stage_2__2621_, data_stage_2__2620_, data_stage_2__2619_, data_stage_2__2618_, data_stage_2__2617_, data_stage_2__2616_, data_stage_2__2615_, data_stage_2__2614_, data_stage_2__2613_, data_stage_2__2612_, data_stage_2__2611_, data_stage_2__2610_, data_stage_2__2609_, data_stage_2__2608_, data_stage_2__2607_, data_stage_2__2606_, data_stage_2__2605_, data_stage_2__2604_, data_stage_2__2603_, data_stage_2__2602_, data_stage_2__2601_, data_stage_2__2600_, data_stage_2__2599_, data_stage_2__2598_, data_stage_2__2597_, data_stage_2__2596_, data_stage_2__2595_, data_stage_2__2594_, data_stage_2__2593_, data_stage_2__2592_, data_stage_2__2591_, data_stage_2__2590_, data_stage_2__2589_, data_stage_2__2588_, data_stage_2__2587_, data_stage_2__2586_, data_stage_2__2585_, data_stage_2__2584_, data_stage_2__2583_, data_stage_2__2582_, data_stage_2__2581_, data_stage_2__2580_, data_stage_2__2579_, data_stage_2__2578_, data_stage_2__2577_, data_stage_2__2576_, data_stage_2__2575_, data_stage_2__2574_, data_stage_2__2573_, data_stage_2__2572_, data_stage_2__2571_, data_stage_2__2570_, data_stage_2__2569_, data_stage_2__2568_, data_stage_2__2567_, data_stage_2__2566_, data_stage_2__2565_, data_stage_2__2564_, data_stage_2__2563_, data_stage_2__2562_, data_stage_2__2561_, data_stage_2__2560_, data_stage_2__2559_, data_stage_2__2558_, data_stage_2__2557_, data_stage_2__2556_, data_stage_2__2555_, data_stage_2__2554_, data_stage_2__2553_, data_stage_2__2552_, data_stage_2__2551_, data_stage_2__2550_, data_stage_2__2549_, data_stage_2__2548_, data_stage_2__2547_, data_stage_2__2546_, data_stage_2__2545_, data_stage_2__2544_, data_stage_2__2543_, data_stage_2__2542_, data_stage_2__2541_, data_stage_2__2540_, data_stage_2__2539_, data_stage_2__2538_, data_stage_2__2537_, data_stage_2__2536_, data_stage_2__2535_, data_stage_2__2534_, data_stage_2__2533_, data_stage_2__2532_, data_stage_2__2531_, data_stage_2__2530_, data_stage_2__2529_, data_stage_2__2528_, data_stage_2__2527_, data_stage_2__2526_, data_stage_2__2525_, data_stage_2__2524_, data_stage_2__2523_, data_stage_2__2522_, data_stage_2__2521_, data_stage_2__2520_, data_stage_2__2519_, data_stage_2__2518_, data_stage_2__2517_, data_stage_2__2516_, data_stage_2__2515_, data_stage_2__2514_, data_stage_2__2513_, data_stage_2__2512_, data_stage_2__2511_, data_stage_2__2510_, data_stage_2__2509_, data_stage_2__2508_, data_stage_2__2507_, data_stage_2__2506_, data_stage_2__2505_, data_stage_2__2504_, data_stage_2__2503_, data_stage_2__2502_, data_stage_2__2501_, data_stage_2__2500_, data_stage_2__2499_, data_stage_2__2498_, data_stage_2__2497_, data_stage_2__2496_, data_stage_2__2495_, data_stage_2__2494_, data_stage_2__2493_, data_stage_2__2492_, data_stage_2__2491_, data_stage_2__2490_, data_stage_2__2489_, data_stage_2__2488_, data_stage_2__2487_, data_stage_2__2486_, data_stage_2__2485_, data_stage_2__2484_, data_stage_2__2483_, data_stage_2__2482_, data_stage_2__2481_, data_stage_2__2480_, data_stage_2__2479_, data_stage_2__2478_, data_stage_2__2477_, data_stage_2__2476_, data_stage_2__2475_, data_stage_2__2474_, data_stage_2__2473_, data_stage_2__2472_, data_stage_2__2471_, data_stage_2__2470_, data_stage_2__2469_, data_stage_2__2468_, data_stage_2__2467_, data_stage_2__2466_, data_stage_2__2465_, data_stage_2__2464_, data_stage_2__2463_, data_stage_2__2462_, data_stage_2__2461_, data_stage_2__2460_, data_stage_2__2459_, data_stage_2__2458_, data_stage_2__2457_, data_stage_2__2456_, data_stage_2__2455_, data_stage_2__2454_, data_stage_2__2453_, data_stage_2__2452_, data_stage_2__2451_, data_stage_2__2450_, data_stage_2__2449_, data_stage_2__2448_, data_stage_2__2447_, data_stage_2__2446_, data_stage_2__2445_, data_stage_2__2444_, data_stage_2__2443_, data_stage_2__2442_, data_stage_2__2441_, data_stage_2__2440_, data_stage_2__2439_, data_stage_2__2438_, data_stage_2__2437_, data_stage_2__2436_, data_stage_2__2435_, data_stage_2__2434_, data_stage_2__2433_, data_stage_2__2432_, data_stage_2__2431_, data_stage_2__2430_, data_stage_2__2429_, data_stage_2__2428_, data_stage_2__2427_, data_stage_2__2426_, data_stage_2__2425_, data_stage_2__2424_, data_stage_2__2423_, data_stage_2__2422_, data_stage_2__2421_, data_stage_2__2420_, data_stage_2__2419_, data_stage_2__2418_, data_stage_2__2417_, data_stage_2__2416_, data_stage_2__2415_, data_stage_2__2414_, data_stage_2__2413_, data_stage_2__2412_, data_stage_2__2411_, data_stage_2__2410_, data_stage_2__2409_, data_stage_2__2408_, data_stage_2__2407_, data_stage_2__2406_, data_stage_2__2405_, data_stage_2__2404_, data_stage_2__2403_, data_stage_2__2402_, data_stage_2__2401_, data_stage_2__2400_, data_stage_2__2399_, data_stage_2__2398_, data_stage_2__2397_, data_stage_2__2396_, data_stage_2__2395_, data_stage_2__2394_, data_stage_2__2393_, data_stage_2__2392_, data_stage_2__2391_, data_stage_2__2390_, data_stage_2__2389_, data_stage_2__2388_, data_stage_2__2387_, data_stage_2__2386_, data_stage_2__2385_, data_stage_2__2384_, data_stage_2__2383_, data_stage_2__2382_, data_stage_2__2381_, data_stage_2__2380_, data_stage_2__2379_, data_stage_2__2378_, data_stage_2__2377_, data_stage_2__2376_, data_stage_2__2375_, data_stage_2__2374_, data_stage_2__2373_, data_stage_2__2372_, data_stage_2__2371_, data_stage_2__2370_, data_stage_2__2369_, data_stage_2__2368_, data_stage_2__2367_, data_stage_2__2366_, data_stage_2__2365_, data_stage_2__2364_, data_stage_2__2363_, data_stage_2__2362_, data_stage_2__2361_, data_stage_2__2360_, data_stage_2__2359_, data_stage_2__2358_, data_stage_2__2357_, data_stage_2__2356_, data_stage_2__2355_, data_stage_2__2354_, data_stage_2__2353_, data_stage_2__2352_, data_stage_2__2351_, data_stage_2__2350_, data_stage_2__2349_, data_stage_2__2348_, data_stage_2__2347_, data_stage_2__2346_, data_stage_2__2345_, data_stage_2__2344_, data_stage_2__2343_, data_stage_2__2342_, data_stage_2__2341_, data_stage_2__2340_, data_stage_2__2339_, data_stage_2__2338_, data_stage_2__2337_, data_stage_2__2336_, data_stage_2__2335_, data_stage_2__2334_, data_stage_2__2333_, data_stage_2__2332_, data_stage_2__2331_, data_stage_2__2330_, data_stage_2__2329_, data_stage_2__2328_, data_stage_2__2327_, data_stage_2__2326_, data_stage_2__2325_, data_stage_2__2324_, data_stage_2__2323_, data_stage_2__2322_, data_stage_2__2321_, data_stage_2__2320_, data_stage_2__2319_, data_stage_2__2318_, data_stage_2__2317_, data_stage_2__2316_, data_stage_2__2315_, data_stage_2__2314_, data_stage_2__2313_, data_stage_2__2312_, data_stage_2__2311_, data_stage_2__2310_, data_stage_2__2309_, data_stage_2__2308_, data_stage_2__2307_, data_stage_2__2306_, data_stage_2__2305_, data_stage_2__2304_, data_stage_2__2303_, data_stage_2__2302_, data_stage_2__2301_, data_stage_2__2300_, data_stage_2__2299_, data_stage_2__2298_, data_stage_2__2297_, data_stage_2__2296_, data_stage_2__2295_, data_stage_2__2294_, data_stage_2__2293_, data_stage_2__2292_, data_stage_2__2291_, data_stage_2__2290_, data_stage_2__2289_, data_stage_2__2288_, data_stage_2__2287_, data_stage_2__2286_, data_stage_2__2285_, data_stage_2__2284_, data_stage_2__2283_, data_stage_2__2282_, data_stage_2__2281_, data_stage_2__2280_, data_stage_2__2279_, data_stage_2__2278_, data_stage_2__2277_, data_stage_2__2276_, data_stage_2__2275_, data_stage_2__2274_, data_stage_2__2273_, data_stage_2__2272_, data_stage_2__2271_, data_stage_2__2270_, data_stage_2__2269_, data_stage_2__2268_, data_stage_2__2267_, data_stage_2__2266_, data_stage_2__2265_, data_stage_2__2264_, data_stage_2__2263_, data_stage_2__2262_, data_stage_2__2261_, data_stage_2__2260_, data_stage_2__2259_, data_stage_2__2258_, data_stage_2__2257_, data_stage_2__2256_, data_stage_2__2255_, data_stage_2__2254_, data_stage_2__2253_, data_stage_2__2252_, data_stage_2__2251_, data_stage_2__2250_, data_stage_2__2249_, data_stage_2__2248_, data_stage_2__2247_, data_stage_2__2246_, data_stage_2__2245_, data_stage_2__2244_, data_stage_2__2243_, data_stage_2__2242_, data_stage_2__2241_, data_stage_2__2240_, data_stage_2__2239_, data_stage_2__2238_, data_stage_2__2237_, data_stage_2__2236_, data_stage_2__2235_, data_stage_2__2234_, data_stage_2__2233_, data_stage_2__2232_, data_stage_2__2231_, data_stage_2__2230_, data_stage_2__2229_, data_stage_2__2228_, data_stage_2__2227_, data_stage_2__2226_, data_stage_2__2225_, data_stage_2__2224_, data_stage_2__2223_, data_stage_2__2222_, data_stage_2__2221_, data_stage_2__2220_, data_stage_2__2219_, data_stage_2__2218_, data_stage_2__2217_, data_stage_2__2216_, data_stage_2__2215_, data_stage_2__2214_, data_stage_2__2213_, data_stage_2__2212_, data_stage_2__2211_, data_stage_2__2210_, data_stage_2__2209_, data_stage_2__2208_, data_stage_2__2207_, data_stage_2__2206_, data_stage_2__2205_, data_stage_2__2204_, data_stage_2__2203_, data_stage_2__2202_, data_stage_2__2201_, data_stage_2__2200_, data_stage_2__2199_, data_stage_2__2198_, data_stage_2__2197_, data_stage_2__2196_, data_stage_2__2195_, data_stage_2__2194_, data_stage_2__2193_, data_stage_2__2192_, data_stage_2__2191_, data_stage_2__2190_, data_stage_2__2189_, data_stage_2__2188_, data_stage_2__2187_, data_stage_2__2186_, data_stage_2__2185_, data_stage_2__2184_, data_stage_2__2183_, data_stage_2__2182_, data_stage_2__2181_, data_stage_2__2180_, data_stage_2__2179_, data_stage_2__2178_, data_stage_2__2177_, data_stage_2__2176_, data_stage_2__2175_, data_stage_2__2174_, data_stage_2__2173_, data_stage_2__2172_, data_stage_2__2171_, data_stage_2__2170_, data_stage_2__2169_, data_stage_2__2168_, data_stage_2__2167_, data_stage_2__2166_, data_stage_2__2165_, data_stage_2__2164_, data_stage_2__2163_, data_stage_2__2162_, data_stage_2__2161_, data_stage_2__2160_, data_stage_2__2159_, data_stage_2__2158_, data_stage_2__2157_, data_stage_2__2156_, data_stage_2__2155_, data_stage_2__2154_, data_stage_2__2153_, data_stage_2__2152_, data_stage_2__2151_, data_stage_2__2150_, data_stage_2__2149_, data_stage_2__2148_, data_stage_2__2147_, data_stage_2__2146_, data_stage_2__2145_, data_stage_2__2144_, data_stage_2__2143_, data_stage_2__2142_, data_stage_2__2141_, data_stage_2__2140_, data_stage_2__2139_, data_stage_2__2138_, data_stage_2__2137_, data_stage_2__2136_, data_stage_2__2135_, data_stage_2__2134_, data_stage_2__2133_, data_stage_2__2132_, data_stage_2__2131_, data_stage_2__2130_, data_stage_2__2129_, data_stage_2__2128_, data_stage_2__2127_, data_stage_2__2126_, data_stage_2__2125_, data_stage_2__2124_, data_stage_2__2123_, data_stage_2__2122_, data_stage_2__2121_, data_stage_2__2120_, data_stage_2__2119_, data_stage_2__2118_, data_stage_2__2117_, data_stage_2__2116_, data_stage_2__2115_, data_stage_2__2114_, data_stage_2__2113_, data_stage_2__2112_, data_stage_2__2111_, data_stage_2__2110_, data_stage_2__2109_, data_stage_2__2108_, data_stage_2__2107_, data_stage_2__2106_, data_stage_2__2105_, data_stage_2__2104_, data_stage_2__2103_, data_stage_2__2102_, data_stage_2__2101_, data_stage_2__2100_, data_stage_2__2099_, data_stage_2__2098_, data_stage_2__2097_, data_stage_2__2096_, data_stage_2__2095_, data_stage_2__2094_, data_stage_2__2093_, data_stage_2__2092_, data_stage_2__2091_, data_stage_2__2090_, data_stage_2__2089_, data_stage_2__2088_, data_stage_2__2087_, data_stage_2__2086_, data_stage_2__2085_, data_stage_2__2084_, data_stage_2__2083_, data_stage_2__2082_, data_stage_2__2081_, data_stage_2__2080_, data_stage_2__2079_, data_stage_2__2078_, data_stage_2__2077_, data_stage_2__2076_, data_stage_2__2075_, data_stage_2__2074_, data_stage_2__2073_, data_stage_2__2072_, data_stage_2__2071_, data_stage_2__2070_, data_stage_2__2069_, data_stage_2__2068_, data_stage_2__2067_, data_stage_2__2066_, data_stage_2__2065_, data_stage_2__2064_, data_stage_2__2063_, data_stage_2__2062_, data_stage_2__2061_, data_stage_2__2060_, data_stage_2__2059_, data_stage_2__2058_, data_stage_2__2057_, data_stage_2__2056_, data_stage_2__2055_, data_stage_2__2054_, data_stage_2__2053_, data_stage_2__2052_, data_stage_2__2051_, data_stage_2__2050_, data_stage_2__2049_, data_stage_2__2048_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__3071_, data_stage_3__3070_, data_stage_3__3069_, data_stage_3__3068_, data_stage_3__3067_, data_stage_3__3066_, data_stage_3__3065_, data_stage_3__3064_, data_stage_3__3063_, data_stage_3__3062_, data_stage_3__3061_, data_stage_3__3060_, data_stage_3__3059_, data_stage_3__3058_, data_stage_3__3057_, data_stage_3__3056_, data_stage_3__3055_, data_stage_3__3054_, data_stage_3__3053_, data_stage_3__3052_, data_stage_3__3051_, data_stage_3__3050_, data_stage_3__3049_, data_stage_3__3048_, data_stage_3__3047_, data_stage_3__3046_, data_stage_3__3045_, data_stage_3__3044_, data_stage_3__3043_, data_stage_3__3042_, data_stage_3__3041_, data_stage_3__3040_, data_stage_3__3039_, data_stage_3__3038_, data_stage_3__3037_, data_stage_3__3036_, data_stage_3__3035_, data_stage_3__3034_, data_stage_3__3033_, data_stage_3__3032_, data_stage_3__3031_, data_stage_3__3030_, data_stage_3__3029_, data_stage_3__3028_, data_stage_3__3027_, data_stage_3__3026_, data_stage_3__3025_, data_stage_3__3024_, data_stage_3__3023_, data_stage_3__3022_, data_stage_3__3021_, data_stage_3__3020_, data_stage_3__3019_, data_stage_3__3018_, data_stage_3__3017_, data_stage_3__3016_, data_stage_3__3015_, data_stage_3__3014_, data_stage_3__3013_, data_stage_3__3012_, data_stage_3__3011_, data_stage_3__3010_, data_stage_3__3009_, data_stage_3__3008_, data_stage_3__3007_, data_stage_3__3006_, data_stage_3__3005_, data_stage_3__3004_, data_stage_3__3003_, data_stage_3__3002_, data_stage_3__3001_, data_stage_3__3000_, data_stage_3__2999_, data_stage_3__2998_, data_stage_3__2997_, data_stage_3__2996_, data_stage_3__2995_, data_stage_3__2994_, data_stage_3__2993_, data_stage_3__2992_, data_stage_3__2991_, data_stage_3__2990_, data_stage_3__2989_, data_stage_3__2988_, data_stage_3__2987_, data_stage_3__2986_, data_stage_3__2985_, data_stage_3__2984_, data_stage_3__2983_, data_stage_3__2982_, data_stage_3__2981_, data_stage_3__2980_, data_stage_3__2979_, data_stage_3__2978_, data_stage_3__2977_, data_stage_3__2976_, data_stage_3__2975_, data_stage_3__2974_, data_stage_3__2973_, data_stage_3__2972_, data_stage_3__2971_, data_stage_3__2970_, data_stage_3__2969_, data_stage_3__2968_, data_stage_3__2967_, data_stage_3__2966_, data_stage_3__2965_, data_stage_3__2964_, data_stage_3__2963_, data_stage_3__2962_, data_stage_3__2961_, data_stage_3__2960_, data_stage_3__2959_, data_stage_3__2958_, data_stage_3__2957_, data_stage_3__2956_, data_stage_3__2955_, data_stage_3__2954_, data_stage_3__2953_, data_stage_3__2952_, data_stage_3__2951_, data_stage_3__2950_, data_stage_3__2949_, data_stage_3__2948_, data_stage_3__2947_, data_stage_3__2946_, data_stage_3__2945_, data_stage_3__2944_, data_stage_3__2943_, data_stage_3__2942_, data_stage_3__2941_, data_stage_3__2940_, data_stage_3__2939_, data_stage_3__2938_, data_stage_3__2937_, data_stage_3__2936_, data_stage_3__2935_, data_stage_3__2934_, data_stage_3__2933_, data_stage_3__2932_, data_stage_3__2931_, data_stage_3__2930_, data_stage_3__2929_, data_stage_3__2928_, data_stage_3__2927_, data_stage_3__2926_, data_stage_3__2925_, data_stage_3__2924_, data_stage_3__2923_, data_stage_3__2922_, data_stage_3__2921_, data_stage_3__2920_, data_stage_3__2919_, data_stage_3__2918_, data_stage_3__2917_, data_stage_3__2916_, data_stage_3__2915_, data_stage_3__2914_, data_stage_3__2913_, data_stage_3__2912_, data_stage_3__2911_, data_stage_3__2910_, data_stage_3__2909_, data_stage_3__2908_, data_stage_3__2907_, data_stage_3__2906_, data_stage_3__2905_, data_stage_3__2904_, data_stage_3__2903_, data_stage_3__2902_, data_stage_3__2901_, data_stage_3__2900_, data_stage_3__2899_, data_stage_3__2898_, data_stage_3__2897_, data_stage_3__2896_, data_stage_3__2895_, data_stage_3__2894_, data_stage_3__2893_, data_stage_3__2892_, data_stage_3__2891_, data_stage_3__2890_, data_stage_3__2889_, data_stage_3__2888_, data_stage_3__2887_, data_stage_3__2886_, data_stage_3__2885_, data_stage_3__2884_, data_stage_3__2883_, data_stage_3__2882_, data_stage_3__2881_, data_stage_3__2880_, data_stage_3__2879_, data_stage_3__2878_, data_stage_3__2877_, data_stage_3__2876_, data_stage_3__2875_, data_stage_3__2874_, data_stage_3__2873_, data_stage_3__2872_, data_stage_3__2871_, data_stage_3__2870_, data_stage_3__2869_, data_stage_3__2868_, data_stage_3__2867_, data_stage_3__2866_, data_stage_3__2865_, data_stage_3__2864_, data_stage_3__2863_, data_stage_3__2862_, data_stage_3__2861_, data_stage_3__2860_, data_stage_3__2859_, data_stage_3__2858_, data_stage_3__2857_, data_stage_3__2856_, data_stage_3__2855_, data_stage_3__2854_, data_stage_3__2853_, data_stage_3__2852_, data_stage_3__2851_, data_stage_3__2850_, data_stage_3__2849_, data_stage_3__2848_, data_stage_3__2847_, data_stage_3__2846_, data_stage_3__2845_, data_stage_3__2844_, data_stage_3__2843_, data_stage_3__2842_, data_stage_3__2841_, data_stage_3__2840_, data_stage_3__2839_, data_stage_3__2838_, data_stage_3__2837_, data_stage_3__2836_, data_stage_3__2835_, data_stage_3__2834_, data_stage_3__2833_, data_stage_3__2832_, data_stage_3__2831_, data_stage_3__2830_, data_stage_3__2829_, data_stage_3__2828_, data_stage_3__2827_, data_stage_3__2826_, data_stage_3__2825_, data_stage_3__2824_, data_stage_3__2823_, data_stage_3__2822_, data_stage_3__2821_, data_stage_3__2820_, data_stage_3__2819_, data_stage_3__2818_, data_stage_3__2817_, data_stage_3__2816_, data_stage_3__2815_, data_stage_3__2814_, data_stage_3__2813_, data_stage_3__2812_, data_stage_3__2811_, data_stage_3__2810_, data_stage_3__2809_, data_stage_3__2808_, data_stage_3__2807_, data_stage_3__2806_, data_stage_3__2805_, data_stage_3__2804_, data_stage_3__2803_, data_stage_3__2802_, data_stage_3__2801_, data_stage_3__2800_, data_stage_3__2799_, data_stage_3__2798_, data_stage_3__2797_, data_stage_3__2796_, data_stage_3__2795_, data_stage_3__2794_, data_stage_3__2793_, data_stage_3__2792_, data_stage_3__2791_, data_stage_3__2790_, data_stage_3__2789_, data_stage_3__2788_, data_stage_3__2787_, data_stage_3__2786_, data_stage_3__2785_, data_stage_3__2784_, data_stage_3__2783_, data_stage_3__2782_, data_stage_3__2781_, data_stage_3__2780_, data_stage_3__2779_, data_stage_3__2778_, data_stage_3__2777_, data_stage_3__2776_, data_stage_3__2775_, data_stage_3__2774_, data_stage_3__2773_, data_stage_3__2772_, data_stage_3__2771_, data_stage_3__2770_, data_stage_3__2769_, data_stage_3__2768_, data_stage_3__2767_, data_stage_3__2766_, data_stage_3__2765_, data_stage_3__2764_, data_stage_3__2763_, data_stage_3__2762_, data_stage_3__2761_, data_stage_3__2760_, data_stage_3__2759_, data_stage_3__2758_, data_stage_3__2757_, data_stage_3__2756_, data_stage_3__2755_, data_stage_3__2754_, data_stage_3__2753_, data_stage_3__2752_, data_stage_3__2751_, data_stage_3__2750_, data_stage_3__2749_, data_stage_3__2748_, data_stage_3__2747_, data_stage_3__2746_, data_stage_3__2745_, data_stage_3__2744_, data_stage_3__2743_, data_stage_3__2742_, data_stage_3__2741_, data_stage_3__2740_, data_stage_3__2739_, data_stage_3__2738_, data_stage_3__2737_, data_stage_3__2736_, data_stage_3__2735_, data_stage_3__2734_, data_stage_3__2733_, data_stage_3__2732_, data_stage_3__2731_, data_stage_3__2730_, data_stage_3__2729_, data_stage_3__2728_, data_stage_3__2727_, data_stage_3__2726_, data_stage_3__2725_, data_stage_3__2724_, data_stage_3__2723_, data_stage_3__2722_, data_stage_3__2721_, data_stage_3__2720_, data_stage_3__2719_, data_stage_3__2718_, data_stage_3__2717_, data_stage_3__2716_, data_stage_3__2715_, data_stage_3__2714_, data_stage_3__2713_, data_stage_3__2712_, data_stage_3__2711_, data_stage_3__2710_, data_stage_3__2709_, data_stage_3__2708_, data_stage_3__2707_, data_stage_3__2706_, data_stage_3__2705_, data_stage_3__2704_, data_stage_3__2703_, data_stage_3__2702_, data_stage_3__2701_, data_stage_3__2700_, data_stage_3__2699_, data_stage_3__2698_, data_stage_3__2697_, data_stage_3__2696_, data_stage_3__2695_, data_stage_3__2694_, data_stage_3__2693_, data_stage_3__2692_, data_stage_3__2691_, data_stage_3__2690_, data_stage_3__2689_, data_stage_3__2688_, data_stage_3__2687_, data_stage_3__2686_, data_stage_3__2685_, data_stage_3__2684_, data_stage_3__2683_, data_stage_3__2682_, data_stage_3__2681_, data_stage_3__2680_, data_stage_3__2679_, data_stage_3__2678_, data_stage_3__2677_, data_stage_3__2676_, data_stage_3__2675_, data_stage_3__2674_, data_stage_3__2673_, data_stage_3__2672_, data_stage_3__2671_, data_stage_3__2670_, data_stage_3__2669_, data_stage_3__2668_, data_stage_3__2667_, data_stage_3__2666_, data_stage_3__2665_, data_stage_3__2664_, data_stage_3__2663_, data_stage_3__2662_, data_stage_3__2661_, data_stage_3__2660_, data_stage_3__2659_, data_stage_3__2658_, data_stage_3__2657_, data_stage_3__2656_, data_stage_3__2655_, data_stage_3__2654_, data_stage_3__2653_, data_stage_3__2652_, data_stage_3__2651_, data_stage_3__2650_, data_stage_3__2649_, data_stage_3__2648_, data_stage_3__2647_, data_stage_3__2646_, data_stage_3__2645_, data_stage_3__2644_, data_stage_3__2643_, data_stage_3__2642_, data_stage_3__2641_, data_stage_3__2640_, data_stage_3__2639_, data_stage_3__2638_, data_stage_3__2637_, data_stage_3__2636_, data_stage_3__2635_, data_stage_3__2634_, data_stage_3__2633_, data_stage_3__2632_, data_stage_3__2631_, data_stage_3__2630_, data_stage_3__2629_, data_stage_3__2628_, data_stage_3__2627_, data_stage_3__2626_, data_stage_3__2625_, data_stage_3__2624_, data_stage_3__2623_, data_stage_3__2622_, data_stage_3__2621_, data_stage_3__2620_, data_stage_3__2619_, data_stage_3__2618_, data_stage_3__2617_, data_stage_3__2616_, data_stage_3__2615_, data_stage_3__2614_, data_stage_3__2613_, data_stage_3__2612_, data_stage_3__2611_, data_stage_3__2610_, data_stage_3__2609_, data_stage_3__2608_, data_stage_3__2607_, data_stage_3__2606_, data_stage_3__2605_, data_stage_3__2604_, data_stage_3__2603_, data_stage_3__2602_, data_stage_3__2601_, data_stage_3__2600_, data_stage_3__2599_, data_stage_3__2598_, data_stage_3__2597_, data_stage_3__2596_, data_stage_3__2595_, data_stage_3__2594_, data_stage_3__2593_, data_stage_3__2592_, data_stage_3__2591_, data_stage_3__2590_, data_stage_3__2589_, data_stage_3__2588_, data_stage_3__2587_, data_stage_3__2586_, data_stage_3__2585_, data_stage_3__2584_, data_stage_3__2583_, data_stage_3__2582_, data_stage_3__2581_, data_stage_3__2580_, data_stage_3__2579_, data_stage_3__2578_, data_stage_3__2577_, data_stage_3__2576_, data_stage_3__2575_, data_stage_3__2574_, data_stage_3__2573_, data_stage_3__2572_, data_stage_3__2571_, data_stage_3__2570_, data_stage_3__2569_, data_stage_3__2568_, data_stage_3__2567_, data_stage_3__2566_, data_stage_3__2565_, data_stage_3__2564_, data_stage_3__2563_, data_stage_3__2562_, data_stage_3__2561_, data_stage_3__2560_, data_stage_3__2559_, data_stage_3__2558_, data_stage_3__2557_, data_stage_3__2556_, data_stage_3__2555_, data_stage_3__2554_, data_stage_3__2553_, data_stage_3__2552_, data_stage_3__2551_, data_stage_3__2550_, data_stage_3__2549_, data_stage_3__2548_, data_stage_3__2547_, data_stage_3__2546_, data_stage_3__2545_, data_stage_3__2544_, data_stage_3__2543_, data_stage_3__2542_, data_stage_3__2541_, data_stage_3__2540_, data_stage_3__2539_, data_stage_3__2538_, data_stage_3__2537_, data_stage_3__2536_, data_stage_3__2535_, data_stage_3__2534_, data_stage_3__2533_, data_stage_3__2532_, data_stage_3__2531_, data_stage_3__2530_, data_stage_3__2529_, data_stage_3__2528_, data_stage_3__2527_, data_stage_3__2526_, data_stage_3__2525_, data_stage_3__2524_, data_stage_3__2523_, data_stage_3__2522_, data_stage_3__2521_, data_stage_3__2520_, data_stage_3__2519_, data_stage_3__2518_, data_stage_3__2517_, data_stage_3__2516_, data_stage_3__2515_, data_stage_3__2514_, data_stage_3__2513_, data_stage_3__2512_, data_stage_3__2511_, data_stage_3__2510_, data_stage_3__2509_, data_stage_3__2508_, data_stage_3__2507_, data_stage_3__2506_, data_stage_3__2505_, data_stage_3__2504_, data_stage_3__2503_, data_stage_3__2502_, data_stage_3__2501_, data_stage_3__2500_, data_stage_3__2499_, data_stage_3__2498_, data_stage_3__2497_, data_stage_3__2496_, data_stage_3__2495_, data_stage_3__2494_, data_stage_3__2493_, data_stage_3__2492_, data_stage_3__2491_, data_stage_3__2490_, data_stage_3__2489_, data_stage_3__2488_, data_stage_3__2487_, data_stage_3__2486_, data_stage_3__2485_, data_stage_3__2484_, data_stage_3__2483_, data_stage_3__2482_, data_stage_3__2481_, data_stage_3__2480_, data_stage_3__2479_, data_stage_3__2478_, data_stage_3__2477_, data_stage_3__2476_, data_stage_3__2475_, data_stage_3__2474_, data_stage_3__2473_, data_stage_3__2472_, data_stage_3__2471_, data_stage_3__2470_, data_stage_3__2469_, data_stage_3__2468_, data_stage_3__2467_, data_stage_3__2466_, data_stage_3__2465_, data_stage_3__2464_, data_stage_3__2463_, data_stage_3__2462_, data_stage_3__2461_, data_stage_3__2460_, data_stage_3__2459_, data_stage_3__2458_, data_stage_3__2457_, data_stage_3__2456_, data_stage_3__2455_, data_stage_3__2454_, data_stage_3__2453_, data_stage_3__2452_, data_stage_3__2451_, data_stage_3__2450_, data_stage_3__2449_, data_stage_3__2448_, data_stage_3__2447_, data_stage_3__2446_, data_stage_3__2445_, data_stage_3__2444_, data_stage_3__2443_, data_stage_3__2442_, data_stage_3__2441_, data_stage_3__2440_, data_stage_3__2439_, data_stage_3__2438_, data_stage_3__2437_, data_stage_3__2436_, data_stage_3__2435_, data_stage_3__2434_, data_stage_3__2433_, data_stage_3__2432_, data_stage_3__2431_, data_stage_3__2430_, data_stage_3__2429_, data_stage_3__2428_, data_stage_3__2427_, data_stage_3__2426_, data_stage_3__2425_, data_stage_3__2424_, data_stage_3__2423_, data_stage_3__2422_, data_stage_3__2421_, data_stage_3__2420_, data_stage_3__2419_, data_stage_3__2418_, data_stage_3__2417_, data_stage_3__2416_, data_stage_3__2415_, data_stage_3__2414_, data_stage_3__2413_, data_stage_3__2412_, data_stage_3__2411_, data_stage_3__2410_, data_stage_3__2409_, data_stage_3__2408_, data_stage_3__2407_, data_stage_3__2406_, data_stage_3__2405_, data_stage_3__2404_, data_stage_3__2403_, data_stage_3__2402_, data_stage_3__2401_, data_stage_3__2400_, data_stage_3__2399_, data_stage_3__2398_, data_stage_3__2397_, data_stage_3__2396_, data_stage_3__2395_, data_stage_3__2394_, data_stage_3__2393_, data_stage_3__2392_, data_stage_3__2391_, data_stage_3__2390_, data_stage_3__2389_, data_stage_3__2388_, data_stage_3__2387_, data_stage_3__2386_, data_stage_3__2385_, data_stage_3__2384_, data_stage_3__2383_, data_stage_3__2382_, data_stage_3__2381_, data_stage_3__2380_, data_stage_3__2379_, data_stage_3__2378_, data_stage_3__2377_, data_stage_3__2376_, data_stage_3__2375_, data_stage_3__2374_, data_stage_3__2373_, data_stage_3__2372_, data_stage_3__2371_, data_stage_3__2370_, data_stage_3__2369_, data_stage_3__2368_, data_stage_3__2367_, data_stage_3__2366_, data_stage_3__2365_, data_stage_3__2364_, data_stage_3__2363_, data_stage_3__2362_, data_stage_3__2361_, data_stage_3__2360_, data_stage_3__2359_, data_stage_3__2358_, data_stage_3__2357_, data_stage_3__2356_, data_stage_3__2355_, data_stage_3__2354_, data_stage_3__2353_, data_stage_3__2352_, data_stage_3__2351_, data_stage_3__2350_, data_stage_3__2349_, data_stage_3__2348_, data_stage_3__2347_, data_stage_3__2346_, data_stage_3__2345_, data_stage_3__2344_, data_stage_3__2343_, data_stage_3__2342_, data_stage_3__2341_, data_stage_3__2340_, data_stage_3__2339_, data_stage_3__2338_, data_stage_3__2337_, data_stage_3__2336_, data_stage_3__2335_, data_stage_3__2334_, data_stage_3__2333_, data_stage_3__2332_, data_stage_3__2331_, data_stage_3__2330_, data_stage_3__2329_, data_stage_3__2328_, data_stage_3__2327_, data_stage_3__2326_, data_stage_3__2325_, data_stage_3__2324_, data_stage_3__2323_, data_stage_3__2322_, data_stage_3__2321_, data_stage_3__2320_, data_stage_3__2319_, data_stage_3__2318_, data_stage_3__2317_, data_stage_3__2316_, data_stage_3__2315_, data_stage_3__2314_, data_stage_3__2313_, data_stage_3__2312_, data_stage_3__2311_, data_stage_3__2310_, data_stage_3__2309_, data_stage_3__2308_, data_stage_3__2307_, data_stage_3__2306_, data_stage_3__2305_, data_stage_3__2304_, data_stage_3__2303_, data_stage_3__2302_, data_stage_3__2301_, data_stage_3__2300_, data_stage_3__2299_, data_stage_3__2298_, data_stage_3__2297_, data_stage_3__2296_, data_stage_3__2295_, data_stage_3__2294_, data_stage_3__2293_, data_stage_3__2292_, data_stage_3__2291_, data_stage_3__2290_, data_stage_3__2289_, data_stage_3__2288_, data_stage_3__2287_, data_stage_3__2286_, data_stage_3__2285_, data_stage_3__2284_, data_stage_3__2283_, data_stage_3__2282_, data_stage_3__2281_, data_stage_3__2280_, data_stage_3__2279_, data_stage_3__2278_, data_stage_3__2277_, data_stage_3__2276_, data_stage_3__2275_, data_stage_3__2274_, data_stage_3__2273_, data_stage_3__2272_, data_stage_3__2271_, data_stage_3__2270_, data_stage_3__2269_, data_stage_3__2268_, data_stage_3__2267_, data_stage_3__2266_, data_stage_3__2265_, data_stage_3__2264_, data_stage_3__2263_, data_stage_3__2262_, data_stage_3__2261_, data_stage_3__2260_, data_stage_3__2259_, data_stage_3__2258_, data_stage_3__2257_, data_stage_3__2256_, data_stage_3__2255_, data_stage_3__2254_, data_stage_3__2253_, data_stage_3__2252_, data_stage_3__2251_, data_stage_3__2250_, data_stage_3__2249_, data_stage_3__2248_, data_stage_3__2247_, data_stage_3__2246_, data_stage_3__2245_, data_stage_3__2244_, data_stage_3__2243_, data_stage_3__2242_, data_stage_3__2241_, data_stage_3__2240_, data_stage_3__2239_, data_stage_3__2238_, data_stage_3__2237_, data_stage_3__2236_, data_stage_3__2235_, data_stage_3__2234_, data_stage_3__2233_, data_stage_3__2232_, data_stage_3__2231_, data_stage_3__2230_, data_stage_3__2229_, data_stage_3__2228_, data_stage_3__2227_, data_stage_3__2226_, data_stage_3__2225_, data_stage_3__2224_, data_stage_3__2223_, data_stage_3__2222_, data_stage_3__2221_, data_stage_3__2220_, data_stage_3__2219_, data_stage_3__2218_, data_stage_3__2217_, data_stage_3__2216_, data_stage_3__2215_, data_stage_3__2214_, data_stage_3__2213_, data_stage_3__2212_, data_stage_3__2211_, data_stage_3__2210_, data_stage_3__2209_, data_stage_3__2208_, data_stage_3__2207_, data_stage_3__2206_, data_stage_3__2205_, data_stage_3__2204_, data_stage_3__2203_, data_stage_3__2202_, data_stage_3__2201_, data_stage_3__2200_, data_stage_3__2199_, data_stage_3__2198_, data_stage_3__2197_, data_stage_3__2196_, data_stage_3__2195_, data_stage_3__2194_, data_stage_3__2193_, data_stage_3__2192_, data_stage_3__2191_, data_stage_3__2190_, data_stage_3__2189_, data_stage_3__2188_, data_stage_3__2187_, data_stage_3__2186_, data_stage_3__2185_, data_stage_3__2184_, data_stage_3__2183_, data_stage_3__2182_, data_stage_3__2181_, data_stage_3__2180_, data_stage_3__2179_, data_stage_3__2178_, data_stage_3__2177_, data_stage_3__2176_, data_stage_3__2175_, data_stage_3__2174_, data_stage_3__2173_, data_stage_3__2172_, data_stage_3__2171_, data_stage_3__2170_, data_stage_3__2169_, data_stage_3__2168_, data_stage_3__2167_, data_stage_3__2166_, data_stage_3__2165_, data_stage_3__2164_, data_stage_3__2163_, data_stage_3__2162_, data_stage_3__2161_, data_stage_3__2160_, data_stage_3__2159_, data_stage_3__2158_, data_stage_3__2157_, data_stage_3__2156_, data_stage_3__2155_, data_stage_3__2154_, data_stage_3__2153_, data_stage_3__2152_, data_stage_3__2151_, data_stage_3__2150_, data_stage_3__2149_, data_stage_3__2148_, data_stage_3__2147_, data_stage_3__2146_, data_stage_3__2145_, data_stage_3__2144_, data_stage_3__2143_, data_stage_3__2142_, data_stage_3__2141_, data_stage_3__2140_, data_stage_3__2139_, data_stage_3__2138_, data_stage_3__2137_, data_stage_3__2136_, data_stage_3__2135_, data_stage_3__2134_, data_stage_3__2133_, data_stage_3__2132_, data_stage_3__2131_, data_stage_3__2130_, data_stage_3__2129_, data_stage_3__2128_, data_stage_3__2127_, data_stage_3__2126_, data_stage_3__2125_, data_stage_3__2124_, data_stage_3__2123_, data_stage_3__2122_, data_stage_3__2121_, data_stage_3__2120_, data_stage_3__2119_, data_stage_3__2118_, data_stage_3__2117_, data_stage_3__2116_, data_stage_3__2115_, data_stage_3__2114_, data_stage_3__2113_, data_stage_3__2112_, data_stage_3__2111_, data_stage_3__2110_, data_stage_3__2109_, data_stage_3__2108_, data_stage_3__2107_, data_stage_3__2106_, data_stage_3__2105_, data_stage_3__2104_, data_stage_3__2103_, data_stage_3__2102_, data_stage_3__2101_, data_stage_3__2100_, data_stage_3__2099_, data_stage_3__2098_, data_stage_3__2097_, data_stage_3__2096_, data_stage_3__2095_, data_stage_3__2094_, data_stage_3__2093_, data_stage_3__2092_, data_stage_3__2091_, data_stage_3__2090_, data_stage_3__2089_, data_stage_3__2088_, data_stage_3__2087_, data_stage_3__2086_, data_stage_3__2085_, data_stage_3__2084_, data_stage_3__2083_, data_stage_3__2082_, data_stage_3__2081_, data_stage_3__2080_, data_stage_3__2079_, data_stage_3__2078_, data_stage_3__2077_, data_stage_3__2076_, data_stage_3__2075_, data_stage_3__2074_, data_stage_3__2073_, data_stage_3__2072_, data_stage_3__2071_, data_stage_3__2070_, data_stage_3__2069_, data_stage_3__2068_, data_stage_3__2067_, data_stage_3__2066_, data_stage_3__2065_, data_stage_3__2064_, data_stage_3__2063_, data_stage_3__2062_, data_stage_3__2061_, data_stage_3__2060_, data_stage_3__2059_, data_stage_3__2058_, data_stage_3__2057_, data_stage_3__2056_, data_stage_3__2055_, data_stage_3__2054_, data_stage_3__2053_, data_stage_3__2052_, data_stage_3__2051_, data_stage_3__2050_, data_stage_3__2049_, data_stage_3__2048_ })
  );


  bsg_swap_width_p512
  mux_stage_2__mux_swap_3__swap_inst
  (
    .data_i({ data_stage_2__4095_, data_stage_2__4094_, data_stage_2__4093_, data_stage_2__4092_, data_stage_2__4091_, data_stage_2__4090_, data_stage_2__4089_, data_stage_2__4088_, data_stage_2__4087_, data_stage_2__4086_, data_stage_2__4085_, data_stage_2__4084_, data_stage_2__4083_, data_stage_2__4082_, data_stage_2__4081_, data_stage_2__4080_, data_stage_2__4079_, data_stage_2__4078_, data_stage_2__4077_, data_stage_2__4076_, data_stage_2__4075_, data_stage_2__4074_, data_stage_2__4073_, data_stage_2__4072_, data_stage_2__4071_, data_stage_2__4070_, data_stage_2__4069_, data_stage_2__4068_, data_stage_2__4067_, data_stage_2__4066_, data_stage_2__4065_, data_stage_2__4064_, data_stage_2__4063_, data_stage_2__4062_, data_stage_2__4061_, data_stage_2__4060_, data_stage_2__4059_, data_stage_2__4058_, data_stage_2__4057_, data_stage_2__4056_, data_stage_2__4055_, data_stage_2__4054_, data_stage_2__4053_, data_stage_2__4052_, data_stage_2__4051_, data_stage_2__4050_, data_stage_2__4049_, data_stage_2__4048_, data_stage_2__4047_, data_stage_2__4046_, data_stage_2__4045_, data_stage_2__4044_, data_stage_2__4043_, data_stage_2__4042_, data_stage_2__4041_, data_stage_2__4040_, data_stage_2__4039_, data_stage_2__4038_, data_stage_2__4037_, data_stage_2__4036_, data_stage_2__4035_, data_stage_2__4034_, data_stage_2__4033_, data_stage_2__4032_, data_stage_2__4031_, data_stage_2__4030_, data_stage_2__4029_, data_stage_2__4028_, data_stage_2__4027_, data_stage_2__4026_, data_stage_2__4025_, data_stage_2__4024_, data_stage_2__4023_, data_stage_2__4022_, data_stage_2__4021_, data_stage_2__4020_, data_stage_2__4019_, data_stage_2__4018_, data_stage_2__4017_, data_stage_2__4016_, data_stage_2__4015_, data_stage_2__4014_, data_stage_2__4013_, data_stage_2__4012_, data_stage_2__4011_, data_stage_2__4010_, data_stage_2__4009_, data_stage_2__4008_, data_stage_2__4007_, data_stage_2__4006_, data_stage_2__4005_, data_stage_2__4004_, data_stage_2__4003_, data_stage_2__4002_, data_stage_2__4001_, data_stage_2__4000_, data_stage_2__3999_, data_stage_2__3998_, data_stage_2__3997_, data_stage_2__3996_, data_stage_2__3995_, data_stage_2__3994_, data_stage_2__3993_, data_stage_2__3992_, data_stage_2__3991_, data_stage_2__3990_, data_stage_2__3989_, data_stage_2__3988_, data_stage_2__3987_, data_stage_2__3986_, data_stage_2__3985_, data_stage_2__3984_, data_stage_2__3983_, data_stage_2__3982_, data_stage_2__3981_, data_stage_2__3980_, data_stage_2__3979_, data_stage_2__3978_, data_stage_2__3977_, data_stage_2__3976_, data_stage_2__3975_, data_stage_2__3974_, data_stage_2__3973_, data_stage_2__3972_, data_stage_2__3971_, data_stage_2__3970_, data_stage_2__3969_, data_stage_2__3968_, data_stage_2__3967_, data_stage_2__3966_, data_stage_2__3965_, data_stage_2__3964_, data_stage_2__3963_, data_stage_2__3962_, data_stage_2__3961_, data_stage_2__3960_, data_stage_2__3959_, data_stage_2__3958_, data_stage_2__3957_, data_stage_2__3956_, data_stage_2__3955_, data_stage_2__3954_, data_stage_2__3953_, data_stage_2__3952_, data_stage_2__3951_, data_stage_2__3950_, data_stage_2__3949_, data_stage_2__3948_, data_stage_2__3947_, data_stage_2__3946_, data_stage_2__3945_, data_stage_2__3944_, data_stage_2__3943_, data_stage_2__3942_, data_stage_2__3941_, data_stage_2__3940_, data_stage_2__3939_, data_stage_2__3938_, data_stage_2__3937_, data_stage_2__3936_, data_stage_2__3935_, data_stage_2__3934_, data_stage_2__3933_, data_stage_2__3932_, data_stage_2__3931_, data_stage_2__3930_, data_stage_2__3929_, data_stage_2__3928_, data_stage_2__3927_, data_stage_2__3926_, data_stage_2__3925_, data_stage_2__3924_, data_stage_2__3923_, data_stage_2__3922_, data_stage_2__3921_, data_stage_2__3920_, data_stage_2__3919_, data_stage_2__3918_, data_stage_2__3917_, data_stage_2__3916_, data_stage_2__3915_, data_stage_2__3914_, data_stage_2__3913_, data_stage_2__3912_, data_stage_2__3911_, data_stage_2__3910_, data_stage_2__3909_, data_stage_2__3908_, data_stage_2__3907_, data_stage_2__3906_, data_stage_2__3905_, data_stage_2__3904_, data_stage_2__3903_, data_stage_2__3902_, data_stage_2__3901_, data_stage_2__3900_, data_stage_2__3899_, data_stage_2__3898_, data_stage_2__3897_, data_stage_2__3896_, data_stage_2__3895_, data_stage_2__3894_, data_stage_2__3893_, data_stage_2__3892_, data_stage_2__3891_, data_stage_2__3890_, data_stage_2__3889_, data_stage_2__3888_, data_stage_2__3887_, data_stage_2__3886_, data_stage_2__3885_, data_stage_2__3884_, data_stage_2__3883_, data_stage_2__3882_, data_stage_2__3881_, data_stage_2__3880_, data_stage_2__3879_, data_stage_2__3878_, data_stage_2__3877_, data_stage_2__3876_, data_stage_2__3875_, data_stage_2__3874_, data_stage_2__3873_, data_stage_2__3872_, data_stage_2__3871_, data_stage_2__3870_, data_stage_2__3869_, data_stage_2__3868_, data_stage_2__3867_, data_stage_2__3866_, data_stage_2__3865_, data_stage_2__3864_, data_stage_2__3863_, data_stage_2__3862_, data_stage_2__3861_, data_stage_2__3860_, data_stage_2__3859_, data_stage_2__3858_, data_stage_2__3857_, data_stage_2__3856_, data_stage_2__3855_, data_stage_2__3854_, data_stage_2__3853_, data_stage_2__3852_, data_stage_2__3851_, data_stage_2__3850_, data_stage_2__3849_, data_stage_2__3848_, data_stage_2__3847_, data_stage_2__3846_, data_stage_2__3845_, data_stage_2__3844_, data_stage_2__3843_, data_stage_2__3842_, data_stage_2__3841_, data_stage_2__3840_, data_stage_2__3839_, data_stage_2__3838_, data_stage_2__3837_, data_stage_2__3836_, data_stage_2__3835_, data_stage_2__3834_, data_stage_2__3833_, data_stage_2__3832_, data_stage_2__3831_, data_stage_2__3830_, data_stage_2__3829_, data_stage_2__3828_, data_stage_2__3827_, data_stage_2__3826_, data_stage_2__3825_, data_stage_2__3824_, data_stage_2__3823_, data_stage_2__3822_, data_stage_2__3821_, data_stage_2__3820_, data_stage_2__3819_, data_stage_2__3818_, data_stage_2__3817_, data_stage_2__3816_, data_stage_2__3815_, data_stage_2__3814_, data_stage_2__3813_, data_stage_2__3812_, data_stage_2__3811_, data_stage_2__3810_, data_stage_2__3809_, data_stage_2__3808_, data_stage_2__3807_, data_stage_2__3806_, data_stage_2__3805_, data_stage_2__3804_, data_stage_2__3803_, data_stage_2__3802_, data_stage_2__3801_, data_stage_2__3800_, data_stage_2__3799_, data_stage_2__3798_, data_stage_2__3797_, data_stage_2__3796_, data_stage_2__3795_, data_stage_2__3794_, data_stage_2__3793_, data_stage_2__3792_, data_stage_2__3791_, data_stage_2__3790_, data_stage_2__3789_, data_stage_2__3788_, data_stage_2__3787_, data_stage_2__3786_, data_stage_2__3785_, data_stage_2__3784_, data_stage_2__3783_, data_stage_2__3782_, data_stage_2__3781_, data_stage_2__3780_, data_stage_2__3779_, data_stage_2__3778_, data_stage_2__3777_, data_stage_2__3776_, data_stage_2__3775_, data_stage_2__3774_, data_stage_2__3773_, data_stage_2__3772_, data_stage_2__3771_, data_stage_2__3770_, data_stage_2__3769_, data_stage_2__3768_, data_stage_2__3767_, data_stage_2__3766_, data_stage_2__3765_, data_stage_2__3764_, data_stage_2__3763_, data_stage_2__3762_, data_stage_2__3761_, data_stage_2__3760_, data_stage_2__3759_, data_stage_2__3758_, data_stage_2__3757_, data_stage_2__3756_, data_stage_2__3755_, data_stage_2__3754_, data_stage_2__3753_, data_stage_2__3752_, data_stage_2__3751_, data_stage_2__3750_, data_stage_2__3749_, data_stage_2__3748_, data_stage_2__3747_, data_stage_2__3746_, data_stage_2__3745_, data_stage_2__3744_, data_stage_2__3743_, data_stage_2__3742_, data_stage_2__3741_, data_stage_2__3740_, data_stage_2__3739_, data_stage_2__3738_, data_stage_2__3737_, data_stage_2__3736_, data_stage_2__3735_, data_stage_2__3734_, data_stage_2__3733_, data_stage_2__3732_, data_stage_2__3731_, data_stage_2__3730_, data_stage_2__3729_, data_stage_2__3728_, data_stage_2__3727_, data_stage_2__3726_, data_stage_2__3725_, data_stage_2__3724_, data_stage_2__3723_, data_stage_2__3722_, data_stage_2__3721_, data_stage_2__3720_, data_stage_2__3719_, data_stage_2__3718_, data_stage_2__3717_, data_stage_2__3716_, data_stage_2__3715_, data_stage_2__3714_, data_stage_2__3713_, data_stage_2__3712_, data_stage_2__3711_, data_stage_2__3710_, data_stage_2__3709_, data_stage_2__3708_, data_stage_2__3707_, data_stage_2__3706_, data_stage_2__3705_, data_stage_2__3704_, data_stage_2__3703_, data_stage_2__3702_, data_stage_2__3701_, data_stage_2__3700_, data_stage_2__3699_, data_stage_2__3698_, data_stage_2__3697_, data_stage_2__3696_, data_stage_2__3695_, data_stage_2__3694_, data_stage_2__3693_, data_stage_2__3692_, data_stage_2__3691_, data_stage_2__3690_, data_stage_2__3689_, data_stage_2__3688_, data_stage_2__3687_, data_stage_2__3686_, data_stage_2__3685_, data_stage_2__3684_, data_stage_2__3683_, data_stage_2__3682_, data_stage_2__3681_, data_stage_2__3680_, data_stage_2__3679_, data_stage_2__3678_, data_stage_2__3677_, data_stage_2__3676_, data_stage_2__3675_, data_stage_2__3674_, data_stage_2__3673_, data_stage_2__3672_, data_stage_2__3671_, data_stage_2__3670_, data_stage_2__3669_, data_stage_2__3668_, data_stage_2__3667_, data_stage_2__3666_, data_stage_2__3665_, data_stage_2__3664_, data_stage_2__3663_, data_stage_2__3662_, data_stage_2__3661_, data_stage_2__3660_, data_stage_2__3659_, data_stage_2__3658_, data_stage_2__3657_, data_stage_2__3656_, data_stage_2__3655_, data_stage_2__3654_, data_stage_2__3653_, data_stage_2__3652_, data_stage_2__3651_, data_stage_2__3650_, data_stage_2__3649_, data_stage_2__3648_, data_stage_2__3647_, data_stage_2__3646_, data_stage_2__3645_, data_stage_2__3644_, data_stage_2__3643_, data_stage_2__3642_, data_stage_2__3641_, data_stage_2__3640_, data_stage_2__3639_, data_stage_2__3638_, data_stage_2__3637_, data_stage_2__3636_, data_stage_2__3635_, data_stage_2__3634_, data_stage_2__3633_, data_stage_2__3632_, data_stage_2__3631_, data_stage_2__3630_, data_stage_2__3629_, data_stage_2__3628_, data_stage_2__3627_, data_stage_2__3626_, data_stage_2__3625_, data_stage_2__3624_, data_stage_2__3623_, data_stage_2__3622_, data_stage_2__3621_, data_stage_2__3620_, data_stage_2__3619_, data_stage_2__3618_, data_stage_2__3617_, data_stage_2__3616_, data_stage_2__3615_, data_stage_2__3614_, data_stage_2__3613_, data_stage_2__3612_, data_stage_2__3611_, data_stage_2__3610_, data_stage_2__3609_, data_stage_2__3608_, data_stage_2__3607_, data_stage_2__3606_, data_stage_2__3605_, data_stage_2__3604_, data_stage_2__3603_, data_stage_2__3602_, data_stage_2__3601_, data_stage_2__3600_, data_stage_2__3599_, data_stage_2__3598_, data_stage_2__3597_, data_stage_2__3596_, data_stage_2__3595_, data_stage_2__3594_, data_stage_2__3593_, data_stage_2__3592_, data_stage_2__3591_, data_stage_2__3590_, data_stage_2__3589_, data_stage_2__3588_, data_stage_2__3587_, data_stage_2__3586_, data_stage_2__3585_, data_stage_2__3584_, data_stage_2__3583_, data_stage_2__3582_, data_stage_2__3581_, data_stage_2__3580_, data_stage_2__3579_, data_stage_2__3578_, data_stage_2__3577_, data_stage_2__3576_, data_stage_2__3575_, data_stage_2__3574_, data_stage_2__3573_, data_stage_2__3572_, data_stage_2__3571_, data_stage_2__3570_, data_stage_2__3569_, data_stage_2__3568_, data_stage_2__3567_, data_stage_2__3566_, data_stage_2__3565_, data_stage_2__3564_, data_stage_2__3563_, data_stage_2__3562_, data_stage_2__3561_, data_stage_2__3560_, data_stage_2__3559_, data_stage_2__3558_, data_stage_2__3557_, data_stage_2__3556_, data_stage_2__3555_, data_stage_2__3554_, data_stage_2__3553_, data_stage_2__3552_, data_stage_2__3551_, data_stage_2__3550_, data_stage_2__3549_, data_stage_2__3548_, data_stage_2__3547_, data_stage_2__3546_, data_stage_2__3545_, data_stage_2__3544_, data_stage_2__3543_, data_stage_2__3542_, data_stage_2__3541_, data_stage_2__3540_, data_stage_2__3539_, data_stage_2__3538_, data_stage_2__3537_, data_stage_2__3536_, data_stage_2__3535_, data_stage_2__3534_, data_stage_2__3533_, data_stage_2__3532_, data_stage_2__3531_, data_stage_2__3530_, data_stage_2__3529_, data_stage_2__3528_, data_stage_2__3527_, data_stage_2__3526_, data_stage_2__3525_, data_stage_2__3524_, data_stage_2__3523_, data_stage_2__3522_, data_stage_2__3521_, data_stage_2__3520_, data_stage_2__3519_, data_stage_2__3518_, data_stage_2__3517_, data_stage_2__3516_, data_stage_2__3515_, data_stage_2__3514_, data_stage_2__3513_, data_stage_2__3512_, data_stage_2__3511_, data_stage_2__3510_, data_stage_2__3509_, data_stage_2__3508_, data_stage_2__3507_, data_stage_2__3506_, data_stage_2__3505_, data_stage_2__3504_, data_stage_2__3503_, data_stage_2__3502_, data_stage_2__3501_, data_stage_2__3500_, data_stage_2__3499_, data_stage_2__3498_, data_stage_2__3497_, data_stage_2__3496_, data_stage_2__3495_, data_stage_2__3494_, data_stage_2__3493_, data_stage_2__3492_, data_stage_2__3491_, data_stage_2__3490_, data_stage_2__3489_, data_stage_2__3488_, data_stage_2__3487_, data_stage_2__3486_, data_stage_2__3485_, data_stage_2__3484_, data_stage_2__3483_, data_stage_2__3482_, data_stage_2__3481_, data_stage_2__3480_, data_stage_2__3479_, data_stage_2__3478_, data_stage_2__3477_, data_stage_2__3476_, data_stage_2__3475_, data_stage_2__3474_, data_stage_2__3473_, data_stage_2__3472_, data_stage_2__3471_, data_stage_2__3470_, data_stage_2__3469_, data_stage_2__3468_, data_stage_2__3467_, data_stage_2__3466_, data_stage_2__3465_, data_stage_2__3464_, data_stage_2__3463_, data_stage_2__3462_, data_stage_2__3461_, data_stage_2__3460_, data_stage_2__3459_, data_stage_2__3458_, data_stage_2__3457_, data_stage_2__3456_, data_stage_2__3455_, data_stage_2__3454_, data_stage_2__3453_, data_stage_2__3452_, data_stage_2__3451_, data_stage_2__3450_, data_stage_2__3449_, data_stage_2__3448_, data_stage_2__3447_, data_stage_2__3446_, data_stage_2__3445_, data_stage_2__3444_, data_stage_2__3443_, data_stage_2__3442_, data_stage_2__3441_, data_stage_2__3440_, data_stage_2__3439_, data_stage_2__3438_, data_stage_2__3437_, data_stage_2__3436_, data_stage_2__3435_, data_stage_2__3434_, data_stage_2__3433_, data_stage_2__3432_, data_stage_2__3431_, data_stage_2__3430_, data_stage_2__3429_, data_stage_2__3428_, data_stage_2__3427_, data_stage_2__3426_, data_stage_2__3425_, data_stage_2__3424_, data_stage_2__3423_, data_stage_2__3422_, data_stage_2__3421_, data_stage_2__3420_, data_stage_2__3419_, data_stage_2__3418_, data_stage_2__3417_, data_stage_2__3416_, data_stage_2__3415_, data_stage_2__3414_, data_stage_2__3413_, data_stage_2__3412_, data_stage_2__3411_, data_stage_2__3410_, data_stage_2__3409_, data_stage_2__3408_, data_stage_2__3407_, data_stage_2__3406_, data_stage_2__3405_, data_stage_2__3404_, data_stage_2__3403_, data_stage_2__3402_, data_stage_2__3401_, data_stage_2__3400_, data_stage_2__3399_, data_stage_2__3398_, data_stage_2__3397_, data_stage_2__3396_, data_stage_2__3395_, data_stage_2__3394_, data_stage_2__3393_, data_stage_2__3392_, data_stage_2__3391_, data_stage_2__3390_, data_stage_2__3389_, data_stage_2__3388_, data_stage_2__3387_, data_stage_2__3386_, data_stage_2__3385_, data_stage_2__3384_, data_stage_2__3383_, data_stage_2__3382_, data_stage_2__3381_, data_stage_2__3380_, data_stage_2__3379_, data_stage_2__3378_, data_stage_2__3377_, data_stage_2__3376_, data_stage_2__3375_, data_stage_2__3374_, data_stage_2__3373_, data_stage_2__3372_, data_stage_2__3371_, data_stage_2__3370_, data_stage_2__3369_, data_stage_2__3368_, data_stage_2__3367_, data_stage_2__3366_, data_stage_2__3365_, data_stage_2__3364_, data_stage_2__3363_, data_stage_2__3362_, data_stage_2__3361_, data_stage_2__3360_, data_stage_2__3359_, data_stage_2__3358_, data_stage_2__3357_, data_stage_2__3356_, data_stage_2__3355_, data_stage_2__3354_, data_stage_2__3353_, data_stage_2__3352_, data_stage_2__3351_, data_stage_2__3350_, data_stage_2__3349_, data_stage_2__3348_, data_stage_2__3347_, data_stage_2__3346_, data_stage_2__3345_, data_stage_2__3344_, data_stage_2__3343_, data_stage_2__3342_, data_stage_2__3341_, data_stage_2__3340_, data_stage_2__3339_, data_stage_2__3338_, data_stage_2__3337_, data_stage_2__3336_, data_stage_2__3335_, data_stage_2__3334_, data_stage_2__3333_, data_stage_2__3332_, data_stage_2__3331_, data_stage_2__3330_, data_stage_2__3329_, data_stage_2__3328_, data_stage_2__3327_, data_stage_2__3326_, data_stage_2__3325_, data_stage_2__3324_, data_stage_2__3323_, data_stage_2__3322_, data_stage_2__3321_, data_stage_2__3320_, data_stage_2__3319_, data_stage_2__3318_, data_stage_2__3317_, data_stage_2__3316_, data_stage_2__3315_, data_stage_2__3314_, data_stage_2__3313_, data_stage_2__3312_, data_stage_2__3311_, data_stage_2__3310_, data_stage_2__3309_, data_stage_2__3308_, data_stage_2__3307_, data_stage_2__3306_, data_stage_2__3305_, data_stage_2__3304_, data_stage_2__3303_, data_stage_2__3302_, data_stage_2__3301_, data_stage_2__3300_, data_stage_2__3299_, data_stage_2__3298_, data_stage_2__3297_, data_stage_2__3296_, data_stage_2__3295_, data_stage_2__3294_, data_stage_2__3293_, data_stage_2__3292_, data_stage_2__3291_, data_stage_2__3290_, data_stage_2__3289_, data_stage_2__3288_, data_stage_2__3287_, data_stage_2__3286_, data_stage_2__3285_, data_stage_2__3284_, data_stage_2__3283_, data_stage_2__3282_, data_stage_2__3281_, data_stage_2__3280_, data_stage_2__3279_, data_stage_2__3278_, data_stage_2__3277_, data_stage_2__3276_, data_stage_2__3275_, data_stage_2__3274_, data_stage_2__3273_, data_stage_2__3272_, data_stage_2__3271_, data_stage_2__3270_, data_stage_2__3269_, data_stage_2__3268_, data_stage_2__3267_, data_stage_2__3266_, data_stage_2__3265_, data_stage_2__3264_, data_stage_2__3263_, data_stage_2__3262_, data_stage_2__3261_, data_stage_2__3260_, data_stage_2__3259_, data_stage_2__3258_, data_stage_2__3257_, data_stage_2__3256_, data_stage_2__3255_, data_stage_2__3254_, data_stage_2__3253_, data_stage_2__3252_, data_stage_2__3251_, data_stage_2__3250_, data_stage_2__3249_, data_stage_2__3248_, data_stage_2__3247_, data_stage_2__3246_, data_stage_2__3245_, data_stage_2__3244_, data_stage_2__3243_, data_stage_2__3242_, data_stage_2__3241_, data_stage_2__3240_, data_stage_2__3239_, data_stage_2__3238_, data_stage_2__3237_, data_stage_2__3236_, data_stage_2__3235_, data_stage_2__3234_, data_stage_2__3233_, data_stage_2__3232_, data_stage_2__3231_, data_stage_2__3230_, data_stage_2__3229_, data_stage_2__3228_, data_stage_2__3227_, data_stage_2__3226_, data_stage_2__3225_, data_stage_2__3224_, data_stage_2__3223_, data_stage_2__3222_, data_stage_2__3221_, data_stage_2__3220_, data_stage_2__3219_, data_stage_2__3218_, data_stage_2__3217_, data_stage_2__3216_, data_stage_2__3215_, data_stage_2__3214_, data_stage_2__3213_, data_stage_2__3212_, data_stage_2__3211_, data_stage_2__3210_, data_stage_2__3209_, data_stage_2__3208_, data_stage_2__3207_, data_stage_2__3206_, data_stage_2__3205_, data_stage_2__3204_, data_stage_2__3203_, data_stage_2__3202_, data_stage_2__3201_, data_stage_2__3200_, data_stage_2__3199_, data_stage_2__3198_, data_stage_2__3197_, data_stage_2__3196_, data_stage_2__3195_, data_stage_2__3194_, data_stage_2__3193_, data_stage_2__3192_, data_stage_2__3191_, data_stage_2__3190_, data_stage_2__3189_, data_stage_2__3188_, data_stage_2__3187_, data_stage_2__3186_, data_stage_2__3185_, data_stage_2__3184_, data_stage_2__3183_, data_stage_2__3182_, data_stage_2__3181_, data_stage_2__3180_, data_stage_2__3179_, data_stage_2__3178_, data_stage_2__3177_, data_stage_2__3176_, data_stage_2__3175_, data_stage_2__3174_, data_stage_2__3173_, data_stage_2__3172_, data_stage_2__3171_, data_stage_2__3170_, data_stage_2__3169_, data_stage_2__3168_, data_stage_2__3167_, data_stage_2__3166_, data_stage_2__3165_, data_stage_2__3164_, data_stage_2__3163_, data_stage_2__3162_, data_stage_2__3161_, data_stage_2__3160_, data_stage_2__3159_, data_stage_2__3158_, data_stage_2__3157_, data_stage_2__3156_, data_stage_2__3155_, data_stage_2__3154_, data_stage_2__3153_, data_stage_2__3152_, data_stage_2__3151_, data_stage_2__3150_, data_stage_2__3149_, data_stage_2__3148_, data_stage_2__3147_, data_stage_2__3146_, data_stage_2__3145_, data_stage_2__3144_, data_stage_2__3143_, data_stage_2__3142_, data_stage_2__3141_, data_stage_2__3140_, data_stage_2__3139_, data_stage_2__3138_, data_stage_2__3137_, data_stage_2__3136_, data_stage_2__3135_, data_stage_2__3134_, data_stage_2__3133_, data_stage_2__3132_, data_stage_2__3131_, data_stage_2__3130_, data_stage_2__3129_, data_stage_2__3128_, data_stage_2__3127_, data_stage_2__3126_, data_stage_2__3125_, data_stage_2__3124_, data_stage_2__3123_, data_stage_2__3122_, data_stage_2__3121_, data_stage_2__3120_, data_stage_2__3119_, data_stage_2__3118_, data_stage_2__3117_, data_stage_2__3116_, data_stage_2__3115_, data_stage_2__3114_, data_stage_2__3113_, data_stage_2__3112_, data_stage_2__3111_, data_stage_2__3110_, data_stage_2__3109_, data_stage_2__3108_, data_stage_2__3107_, data_stage_2__3106_, data_stage_2__3105_, data_stage_2__3104_, data_stage_2__3103_, data_stage_2__3102_, data_stage_2__3101_, data_stage_2__3100_, data_stage_2__3099_, data_stage_2__3098_, data_stage_2__3097_, data_stage_2__3096_, data_stage_2__3095_, data_stage_2__3094_, data_stage_2__3093_, data_stage_2__3092_, data_stage_2__3091_, data_stage_2__3090_, data_stage_2__3089_, data_stage_2__3088_, data_stage_2__3087_, data_stage_2__3086_, data_stage_2__3085_, data_stage_2__3084_, data_stage_2__3083_, data_stage_2__3082_, data_stage_2__3081_, data_stage_2__3080_, data_stage_2__3079_, data_stage_2__3078_, data_stage_2__3077_, data_stage_2__3076_, data_stage_2__3075_, data_stage_2__3074_, data_stage_2__3073_, data_stage_2__3072_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__4095_, data_stage_3__4094_, data_stage_3__4093_, data_stage_3__4092_, data_stage_3__4091_, data_stage_3__4090_, data_stage_3__4089_, data_stage_3__4088_, data_stage_3__4087_, data_stage_3__4086_, data_stage_3__4085_, data_stage_3__4084_, data_stage_3__4083_, data_stage_3__4082_, data_stage_3__4081_, data_stage_3__4080_, data_stage_3__4079_, data_stage_3__4078_, data_stage_3__4077_, data_stage_3__4076_, data_stage_3__4075_, data_stage_3__4074_, data_stage_3__4073_, data_stage_3__4072_, data_stage_3__4071_, data_stage_3__4070_, data_stage_3__4069_, data_stage_3__4068_, data_stage_3__4067_, data_stage_3__4066_, data_stage_3__4065_, data_stage_3__4064_, data_stage_3__4063_, data_stage_3__4062_, data_stage_3__4061_, data_stage_3__4060_, data_stage_3__4059_, data_stage_3__4058_, data_stage_3__4057_, data_stage_3__4056_, data_stage_3__4055_, data_stage_3__4054_, data_stage_3__4053_, data_stage_3__4052_, data_stage_3__4051_, data_stage_3__4050_, data_stage_3__4049_, data_stage_3__4048_, data_stage_3__4047_, data_stage_3__4046_, data_stage_3__4045_, data_stage_3__4044_, data_stage_3__4043_, data_stage_3__4042_, data_stage_3__4041_, data_stage_3__4040_, data_stage_3__4039_, data_stage_3__4038_, data_stage_3__4037_, data_stage_3__4036_, data_stage_3__4035_, data_stage_3__4034_, data_stage_3__4033_, data_stage_3__4032_, data_stage_3__4031_, data_stage_3__4030_, data_stage_3__4029_, data_stage_3__4028_, data_stage_3__4027_, data_stage_3__4026_, data_stage_3__4025_, data_stage_3__4024_, data_stage_3__4023_, data_stage_3__4022_, data_stage_3__4021_, data_stage_3__4020_, data_stage_3__4019_, data_stage_3__4018_, data_stage_3__4017_, data_stage_3__4016_, data_stage_3__4015_, data_stage_3__4014_, data_stage_3__4013_, data_stage_3__4012_, data_stage_3__4011_, data_stage_3__4010_, data_stage_3__4009_, data_stage_3__4008_, data_stage_3__4007_, data_stage_3__4006_, data_stage_3__4005_, data_stage_3__4004_, data_stage_3__4003_, data_stage_3__4002_, data_stage_3__4001_, data_stage_3__4000_, data_stage_3__3999_, data_stage_3__3998_, data_stage_3__3997_, data_stage_3__3996_, data_stage_3__3995_, data_stage_3__3994_, data_stage_3__3993_, data_stage_3__3992_, data_stage_3__3991_, data_stage_3__3990_, data_stage_3__3989_, data_stage_3__3988_, data_stage_3__3987_, data_stage_3__3986_, data_stage_3__3985_, data_stage_3__3984_, data_stage_3__3983_, data_stage_3__3982_, data_stage_3__3981_, data_stage_3__3980_, data_stage_3__3979_, data_stage_3__3978_, data_stage_3__3977_, data_stage_3__3976_, data_stage_3__3975_, data_stage_3__3974_, data_stage_3__3973_, data_stage_3__3972_, data_stage_3__3971_, data_stage_3__3970_, data_stage_3__3969_, data_stage_3__3968_, data_stage_3__3967_, data_stage_3__3966_, data_stage_3__3965_, data_stage_3__3964_, data_stage_3__3963_, data_stage_3__3962_, data_stage_3__3961_, data_stage_3__3960_, data_stage_3__3959_, data_stage_3__3958_, data_stage_3__3957_, data_stage_3__3956_, data_stage_3__3955_, data_stage_3__3954_, data_stage_3__3953_, data_stage_3__3952_, data_stage_3__3951_, data_stage_3__3950_, data_stage_3__3949_, data_stage_3__3948_, data_stage_3__3947_, data_stage_3__3946_, data_stage_3__3945_, data_stage_3__3944_, data_stage_3__3943_, data_stage_3__3942_, data_stage_3__3941_, data_stage_3__3940_, data_stage_3__3939_, data_stage_3__3938_, data_stage_3__3937_, data_stage_3__3936_, data_stage_3__3935_, data_stage_3__3934_, data_stage_3__3933_, data_stage_3__3932_, data_stage_3__3931_, data_stage_3__3930_, data_stage_3__3929_, data_stage_3__3928_, data_stage_3__3927_, data_stage_3__3926_, data_stage_3__3925_, data_stage_3__3924_, data_stage_3__3923_, data_stage_3__3922_, data_stage_3__3921_, data_stage_3__3920_, data_stage_3__3919_, data_stage_3__3918_, data_stage_3__3917_, data_stage_3__3916_, data_stage_3__3915_, data_stage_3__3914_, data_stage_3__3913_, data_stage_3__3912_, data_stage_3__3911_, data_stage_3__3910_, data_stage_3__3909_, data_stage_3__3908_, data_stage_3__3907_, data_stage_3__3906_, data_stage_3__3905_, data_stage_3__3904_, data_stage_3__3903_, data_stage_3__3902_, data_stage_3__3901_, data_stage_3__3900_, data_stage_3__3899_, data_stage_3__3898_, data_stage_3__3897_, data_stage_3__3896_, data_stage_3__3895_, data_stage_3__3894_, data_stage_3__3893_, data_stage_3__3892_, data_stage_3__3891_, data_stage_3__3890_, data_stage_3__3889_, data_stage_3__3888_, data_stage_3__3887_, data_stage_3__3886_, data_stage_3__3885_, data_stage_3__3884_, data_stage_3__3883_, data_stage_3__3882_, data_stage_3__3881_, data_stage_3__3880_, data_stage_3__3879_, data_stage_3__3878_, data_stage_3__3877_, data_stage_3__3876_, data_stage_3__3875_, data_stage_3__3874_, data_stage_3__3873_, data_stage_3__3872_, data_stage_3__3871_, data_stage_3__3870_, data_stage_3__3869_, data_stage_3__3868_, data_stage_3__3867_, data_stage_3__3866_, data_stage_3__3865_, data_stage_3__3864_, data_stage_3__3863_, data_stage_3__3862_, data_stage_3__3861_, data_stage_3__3860_, data_stage_3__3859_, data_stage_3__3858_, data_stage_3__3857_, data_stage_3__3856_, data_stage_3__3855_, data_stage_3__3854_, data_stage_3__3853_, data_stage_3__3852_, data_stage_3__3851_, data_stage_3__3850_, data_stage_3__3849_, data_stage_3__3848_, data_stage_3__3847_, data_stage_3__3846_, data_stage_3__3845_, data_stage_3__3844_, data_stage_3__3843_, data_stage_3__3842_, data_stage_3__3841_, data_stage_3__3840_, data_stage_3__3839_, data_stage_3__3838_, data_stage_3__3837_, data_stage_3__3836_, data_stage_3__3835_, data_stage_3__3834_, data_stage_3__3833_, data_stage_3__3832_, data_stage_3__3831_, data_stage_3__3830_, data_stage_3__3829_, data_stage_3__3828_, data_stage_3__3827_, data_stage_3__3826_, data_stage_3__3825_, data_stage_3__3824_, data_stage_3__3823_, data_stage_3__3822_, data_stage_3__3821_, data_stage_3__3820_, data_stage_3__3819_, data_stage_3__3818_, data_stage_3__3817_, data_stage_3__3816_, data_stage_3__3815_, data_stage_3__3814_, data_stage_3__3813_, data_stage_3__3812_, data_stage_3__3811_, data_stage_3__3810_, data_stage_3__3809_, data_stage_3__3808_, data_stage_3__3807_, data_stage_3__3806_, data_stage_3__3805_, data_stage_3__3804_, data_stage_3__3803_, data_stage_3__3802_, data_stage_3__3801_, data_stage_3__3800_, data_stage_3__3799_, data_stage_3__3798_, data_stage_3__3797_, data_stage_3__3796_, data_stage_3__3795_, data_stage_3__3794_, data_stage_3__3793_, data_stage_3__3792_, data_stage_3__3791_, data_stage_3__3790_, data_stage_3__3789_, data_stage_3__3788_, data_stage_3__3787_, data_stage_3__3786_, data_stage_3__3785_, data_stage_3__3784_, data_stage_3__3783_, data_stage_3__3782_, data_stage_3__3781_, data_stage_3__3780_, data_stage_3__3779_, data_stage_3__3778_, data_stage_3__3777_, data_stage_3__3776_, data_stage_3__3775_, data_stage_3__3774_, data_stage_3__3773_, data_stage_3__3772_, data_stage_3__3771_, data_stage_3__3770_, data_stage_3__3769_, data_stage_3__3768_, data_stage_3__3767_, data_stage_3__3766_, data_stage_3__3765_, data_stage_3__3764_, data_stage_3__3763_, data_stage_3__3762_, data_stage_3__3761_, data_stage_3__3760_, data_stage_3__3759_, data_stage_3__3758_, data_stage_3__3757_, data_stage_3__3756_, data_stage_3__3755_, data_stage_3__3754_, data_stage_3__3753_, data_stage_3__3752_, data_stage_3__3751_, data_stage_3__3750_, data_stage_3__3749_, data_stage_3__3748_, data_stage_3__3747_, data_stage_3__3746_, data_stage_3__3745_, data_stage_3__3744_, data_stage_3__3743_, data_stage_3__3742_, data_stage_3__3741_, data_stage_3__3740_, data_stage_3__3739_, data_stage_3__3738_, data_stage_3__3737_, data_stage_3__3736_, data_stage_3__3735_, data_stage_3__3734_, data_stage_3__3733_, data_stage_3__3732_, data_stage_3__3731_, data_stage_3__3730_, data_stage_3__3729_, data_stage_3__3728_, data_stage_3__3727_, data_stage_3__3726_, data_stage_3__3725_, data_stage_3__3724_, data_stage_3__3723_, data_stage_3__3722_, data_stage_3__3721_, data_stage_3__3720_, data_stage_3__3719_, data_stage_3__3718_, data_stage_3__3717_, data_stage_3__3716_, data_stage_3__3715_, data_stage_3__3714_, data_stage_3__3713_, data_stage_3__3712_, data_stage_3__3711_, data_stage_3__3710_, data_stage_3__3709_, data_stage_3__3708_, data_stage_3__3707_, data_stage_3__3706_, data_stage_3__3705_, data_stage_3__3704_, data_stage_3__3703_, data_stage_3__3702_, data_stage_3__3701_, data_stage_3__3700_, data_stage_3__3699_, data_stage_3__3698_, data_stage_3__3697_, data_stage_3__3696_, data_stage_3__3695_, data_stage_3__3694_, data_stage_3__3693_, data_stage_3__3692_, data_stage_3__3691_, data_stage_3__3690_, data_stage_3__3689_, data_stage_3__3688_, data_stage_3__3687_, data_stage_3__3686_, data_stage_3__3685_, data_stage_3__3684_, data_stage_3__3683_, data_stage_3__3682_, data_stage_3__3681_, data_stage_3__3680_, data_stage_3__3679_, data_stage_3__3678_, data_stage_3__3677_, data_stage_3__3676_, data_stage_3__3675_, data_stage_3__3674_, data_stage_3__3673_, data_stage_3__3672_, data_stage_3__3671_, data_stage_3__3670_, data_stage_3__3669_, data_stage_3__3668_, data_stage_3__3667_, data_stage_3__3666_, data_stage_3__3665_, data_stage_3__3664_, data_stage_3__3663_, data_stage_3__3662_, data_stage_3__3661_, data_stage_3__3660_, data_stage_3__3659_, data_stage_3__3658_, data_stage_3__3657_, data_stage_3__3656_, data_stage_3__3655_, data_stage_3__3654_, data_stage_3__3653_, data_stage_3__3652_, data_stage_3__3651_, data_stage_3__3650_, data_stage_3__3649_, data_stage_3__3648_, data_stage_3__3647_, data_stage_3__3646_, data_stage_3__3645_, data_stage_3__3644_, data_stage_3__3643_, data_stage_3__3642_, data_stage_3__3641_, data_stage_3__3640_, data_stage_3__3639_, data_stage_3__3638_, data_stage_3__3637_, data_stage_3__3636_, data_stage_3__3635_, data_stage_3__3634_, data_stage_3__3633_, data_stage_3__3632_, data_stage_3__3631_, data_stage_3__3630_, data_stage_3__3629_, data_stage_3__3628_, data_stage_3__3627_, data_stage_3__3626_, data_stage_3__3625_, data_stage_3__3624_, data_stage_3__3623_, data_stage_3__3622_, data_stage_3__3621_, data_stage_3__3620_, data_stage_3__3619_, data_stage_3__3618_, data_stage_3__3617_, data_stage_3__3616_, data_stage_3__3615_, data_stage_3__3614_, data_stage_3__3613_, data_stage_3__3612_, data_stage_3__3611_, data_stage_3__3610_, data_stage_3__3609_, data_stage_3__3608_, data_stage_3__3607_, data_stage_3__3606_, data_stage_3__3605_, data_stage_3__3604_, data_stage_3__3603_, data_stage_3__3602_, data_stage_3__3601_, data_stage_3__3600_, data_stage_3__3599_, data_stage_3__3598_, data_stage_3__3597_, data_stage_3__3596_, data_stage_3__3595_, data_stage_3__3594_, data_stage_3__3593_, data_stage_3__3592_, data_stage_3__3591_, data_stage_3__3590_, data_stage_3__3589_, data_stage_3__3588_, data_stage_3__3587_, data_stage_3__3586_, data_stage_3__3585_, data_stage_3__3584_, data_stage_3__3583_, data_stage_3__3582_, data_stage_3__3581_, data_stage_3__3580_, data_stage_3__3579_, data_stage_3__3578_, data_stage_3__3577_, data_stage_3__3576_, data_stage_3__3575_, data_stage_3__3574_, data_stage_3__3573_, data_stage_3__3572_, data_stage_3__3571_, data_stage_3__3570_, data_stage_3__3569_, data_stage_3__3568_, data_stage_3__3567_, data_stage_3__3566_, data_stage_3__3565_, data_stage_3__3564_, data_stage_3__3563_, data_stage_3__3562_, data_stage_3__3561_, data_stage_3__3560_, data_stage_3__3559_, data_stage_3__3558_, data_stage_3__3557_, data_stage_3__3556_, data_stage_3__3555_, data_stage_3__3554_, data_stage_3__3553_, data_stage_3__3552_, data_stage_3__3551_, data_stage_3__3550_, data_stage_3__3549_, data_stage_3__3548_, data_stage_3__3547_, data_stage_3__3546_, data_stage_3__3545_, data_stage_3__3544_, data_stage_3__3543_, data_stage_3__3542_, data_stage_3__3541_, data_stage_3__3540_, data_stage_3__3539_, data_stage_3__3538_, data_stage_3__3537_, data_stage_3__3536_, data_stage_3__3535_, data_stage_3__3534_, data_stage_3__3533_, data_stage_3__3532_, data_stage_3__3531_, data_stage_3__3530_, data_stage_3__3529_, data_stage_3__3528_, data_stage_3__3527_, data_stage_3__3526_, data_stage_3__3525_, data_stage_3__3524_, data_stage_3__3523_, data_stage_3__3522_, data_stage_3__3521_, data_stage_3__3520_, data_stage_3__3519_, data_stage_3__3518_, data_stage_3__3517_, data_stage_3__3516_, data_stage_3__3515_, data_stage_3__3514_, data_stage_3__3513_, data_stage_3__3512_, data_stage_3__3511_, data_stage_3__3510_, data_stage_3__3509_, data_stage_3__3508_, data_stage_3__3507_, data_stage_3__3506_, data_stage_3__3505_, data_stage_3__3504_, data_stage_3__3503_, data_stage_3__3502_, data_stage_3__3501_, data_stage_3__3500_, data_stage_3__3499_, data_stage_3__3498_, data_stage_3__3497_, data_stage_3__3496_, data_stage_3__3495_, data_stage_3__3494_, data_stage_3__3493_, data_stage_3__3492_, data_stage_3__3491_, data_stage_3__3490_, data_stage_3__3489_, data_stage_3__3488_, data_stage_3__3487_, data_stage_3__3486_, data_stage_3__3485_, data_stage_3__3484_, data_stage_3__3483_, data_stage_3__3482_, data_stage_3__3481_, data_stage_3__3480_, data_stage_3__3479_, data_stage_3__3478_, data_stage_3__3477_, data_stage_3__3476_, data_stage_3__3475_, data_stage_3__3474_, data_stage_3__3473_, data_stage_3__3472_, data_stage_3__3471_, data_stage_3__3470_, data_stage_3__3469_, data_stage_3__3468_, data_stage_3__3467_, data_stage_3__3466_, data_stage_3__3465_, data_stage_3__3464_, data_stage_3__3463_, data_stage_3__3462_, data_stage_3__3461_, data_stage_3__3460_, data_stage_3__3459_, data_stage_3__3458_, data_stage_3__3457_, data_stage_3__3456_, data_stage_3__3455_, data_stage_3__3454_, data_stage_3__3453_, data_stage_3__3452_, data_stage_3__3451_, data_stage_3__3450_, data_stage_3__3449_, data_stage_3__3448_, data_stage_3__3447_, data_stage_3__3446_, data_stage_3__3445_, data_stage_3__3444_, data_stage_3__3443_, data_stage_3__3442_, data_stage_3__3441_, data_stage_3__3440_, data_stage_3__3439_, data_stage_3__3438_, data_stage_3__3437_, data_stage_3__3436_, data_stage_3__3435_, data_stage_3__3434_, data_stage_3__3433_, data_stage_3__3432_, data_stage_3__3431_, data_stage_3__3430_, data_stage_3__3429_, data_stage_3__3428_, data_stage_3__3427_, data_stage_3__3426_, data_stage_3__3425_, data_stage_3__3424_, data_stage_3__3423_, data_stage_3__3422_, data_stage_3__3421_, data_stage_3__3420_, data_stage_3__3419_, data_stage_3__3418_, data_stage_3__3417_, data_stage_3__3416_, data_stage_3__3415_, data_stage_3__3414_, data_stage_3__3413_, data_stage_3__3412_, data_stage_3__3411_, data_stage_3__3410_, data_stage_3__3409_, data_stage_3__3408_, data_stage_3__3407_, data_stage_3__3406_, data_stage_3__3405_, data_stage_3__3404_, data_stage_3__3403_, data_stage_3__3402_, data_stage_3__3401_, data_stage_3__3400_, data_stage_3__3399_, data_stage_3__3398_, data_stage_3__3397_, data_stage_3__3396_, data_stage_3__3395_, data_stage_3__3394_, data_stage_3__3393_, data_stage_3__3392_, data_stage_3__3391_, data_stage_3__3390_, data_stage_3__3389_, data_stage_3__3388_, data_stage_3__3387_, data_stage_3__3386_, data_stage_3__3385_, data_stage_3__3384_, data_stage_3__3383_, data_stage_3__3382_, data_stage_3__3381_, data_stage_3__3380_, data_stage_3__3379_, data_stage_3__3378_, data_stage_3__3377_, data_stage_3__3376_, data_stage_3__3375_, data_stage_3__3374_, data_stage_3__3373_, data_stage_3__3372_, data_stage_3__3371_, data_stage_3__3370_, data_stage_3__3369_, data_stage_3__3368_, data_stage_3__3367_, data_stage_3__3366_, data_stage_3__3365_, data_stage_3__3364_, data_stage_3__3363_, data_stage_3__3362_, data_stage_3__3361_, data_stage_3__3360_, data_stage_3__3359_, data_stage_3__3358_, data_stage_3__3357_, data_stage_3__3356_, data_stage_3__3355_, data_stage_3__3354_, data_stage_3__3353_, data_stage_3__3352_, data_stage_3__3351_, data_stage_3__3350_, data_stage_3__3349_, data_stage_3__3348_, data_stage_3__3347_, data_stage_3__3346_, data_stage_3__3345_, data_stage_3__3344_, data_stage_3__3343_, data_stage_3__3342_, data_stage_3__3341_, data_stage_3__3340_, data_stage_3__3339_, data_stage_3__3338_, data_stage_3__3337_, data_stage_3__3336_, data_stage_3__3335_, data_stage_3__3334_, data_stage_3__3333_, data_stage_3__3332_, data_stage_3__3331_, data_stage_3__3330_, data_stage_3__3329_, data_stage_3__3328_, data_stage_3__3327_, data_stage_3__3326_, data_stage_3__3325_, data_stage_3__3324_, data_stage_3__3323_, data_stage_3__3322_, data_stage_3__3321_, data_stage_3__3320_, data_stage_3__3319_, data_stage_3__3318_, data_stage_3__3317_, data_stage_3__3316_, data_stage_3__3315_, data_stage_3__3314_, data_stage_3__3313_, data_stage_3__3312_, data_stage_3__3311_, data_stage_3__3310_, data_stage_3__3309_, data_stage_3__3308_, data_stage_3__3307_, data_stage_3__3306_, data_stage_3__3305_, data_stage_3__3304_, data_stage_3__3303_, data_stage_3__3302_, data_stage_3__3301_, data_stage_3__3300_, data_stage_3__3299_, data_stage_3__3298_, data_stage_3__3297_, data_stage_3__3296_, data_stage_3__3295_, data_stage_3__3294_, data_stage_3__3293_, data_stage_3__3292_, data_stage_3__3291_, data_stage_3__3290_, data_stage_3__3289_, data_stage_3__3288_, data_stage_3__3287_, data_stage_3__3286_, data_stage_3__3285_, data_stage_3__3284_, data_stage_3__3283_, data_stage_3__3282_, data_stage_3__3281_, data_stage_3__3280_, data_stage_3__3279_, data_stage_3__3278_, data_stage_3__3277_, data_stage_3__3276_, data_stage_3__3275_, data_stage_3__3274_, data_stage_3__3273_, data_stage_3__3272_, data_stage_3__3271_, data_stage_3__3270_, data_stage_3__3269_, data_stage_3__3268_, data_stage_3__3267_, data_stage_3__3266_, data_stage_3__3265_, data_stage_3__3264_, data_stage_3__3263_, data_stage_3__3262_, data_stage_3__3261_, data_stage_3__3260_, data_stage_3__3259_, data_stage_3__3258_, data_stage_3__3257_, data_stage_3__3256_, data_stage_3__3255_, data_stage_3__3254_, data_stage_3__3253_, data_stage_3__3252_, data_stage_3__3251_, data_stage_3__3250_, data_stage_3__3249_, data_stage_3__3248_, data_stage_3__3247_, data_stage_3__3246_, data_stage_3__3245_, data_stage_3__3244_, data_stage_3__3243_, data_stage_3__3242_, data_stage_3__3241_, data_stage_3__3240_, data_stage_3__3239_, data_stage_3__3238_, data_stage_3__3237_, data_stage_3__3236_, data_stage_3__3235_, data_stage_3__3234_, data_stage_3__3233_, data_stage_3__3232_, data_stage_3__3231_, data_stage_3__3230_, data_stage_3__3229_, data_stage_3__3228_, data_stage_3__3227_, data_stage_3__3226_, data_stage_3__3225_, data_stage_3__3224_, data_stage_3__3223_, data_stage_3__3222_, data_stage_3__3221_, data_stage_3__3220_, data_stage_3__3219_, data_stage_3__3218_, data_stage_3__3217_, data_stage_3__3216_, data_stage_3__3215_, data_stage_3__3214_, data_stage_3__3213_, data_stage_3__3212_, data_stage_3__3211_, data_stage_3__3210_, data_stage_3__3209_, data_stage_3__3208_, data_stage_3__3207_, data_stage_3__3206_, data_stage_3__3205_, data_stage_3__3204_, data_stage_3__3203_, data_stage_3__3202_, data_stage_3__3201_, data_stage_3__3200_, data_stage_3__3199_, data_stage_3__3198_, data_stage_3__3197_, data_stage_3__3196_, data_stage_3__3195_, data_stage_3__3194_, data_stage_3__3193_, data_stage_3__3192_, data_stage_3__3191_, data_stage_3__3190_, data_stage_3__3189_, data_stage_3__3188_, data_stage_3__3187_, data_stage_3__3186_, data_stage_3__3185_, data_stage_3__3184_, data_stage_3__3183_, data_stage_3__3182_, data_stage_3__3181_, data_stage_3__3180_, data_stage_3__3179_, data_stage_3__3178_, data_stage_3__3177_, data_stage_3__3176_, data_stage_3__3175_, data_stage_3__3174_, data_stage_3__3173_, data_stage_3__3172_, data_stage_3__3171_, data_stage_3__3170_, data_stage_3__3169_, data_stage_3__3168_, data_stage_3__3167_, data_stage_3__3166_, data_stage_3__3165_, data_stage_3__3164_, data_stage_3__3163_, data_stage_3__3162_, data_stage_3__3161_, data_stage_3__3160_, data_stage_3__3159_, data_stage_3__3158_, data_stage_3__3157_, data_stage_3__3156_, data_stage_3__3155_, data_stage_3__3154_, data_stage_3__3153_, data_stage_3__3152_, data_stage_3__3151_, data_stage_3__3150_, data_stage_3__3149_, data_stage_3__3148_, data_stage_3__3147_, data_stage_3__3146_, data_stage_3__3145_, data_stage_3__3144_, data_stage_3__3143_, data_stage_3__3142_, data_stage_3__3141_, data_stage_3__3140_, data_stage_3__3139_, data_stage_3__3138_, data_stage_3__3137_, data_stage_3__3136_, data_stage_3__3135_, data_stage_3__3134_, data_stage_3__3133_, data_stage_3__3132_, data_stage_3__3131_, data_stage_3__3130_, data_stage_3__3129_, data_stage_3__3128_, data_stage_3__3127_, data_stage_3__3126_, data_stage_3__3125_, data_stage_3__3124_, data_stage_3__3123_, data_stage_3__3122_, data_stage_3__3121_, data_stage_3__3120_, data_stage_3__3119_, data_stage_3__3118_, data_stage_3__3117_, data_stage_3__3116_, data_stage_3__3115_, data_stage_3__3114_, data_stage_3__3113_, data_stage_3__3112_, data_stage_3__3111_, data_stage_3__3110_, data_stage_3__3109_, data_stage_3__3108_, data_stage_3__3107_, data_stage_3__3106_, data_stage_3__3105_, data_stage_3__3104_, data_stage_3__3103_, data_stage_3__3102_, data_stage_3__3101_, data_stage_3__3100_, data_stage_3__3099_, data_stage_3__3098_, data_stage_3__3097_, data_stage_3__3096_, data_stage_3__3095_, data_stage_3__3094_, data_stage_3__3093_, data_stage_3__3092_, data_stage_3__3091_, data_stage_3__3090_, data_stage_3__3089_, data_stage_3__3088_, data_stage_3__3087_, data_stage_3__3086_, data_stage_3__3085_, data_stage_3__3084_, data_stage_3__3083_, data_stage_3__3082_, data_stage_3__3081_, data_stage_3__3080_, data_stage_3__3079_, data_stage_3__3078_, data_stage_3__3077_, data_stage_3__3076_, data_stage_3__3075_, data_stage_3__3074_, data_stage_3__3073_, data_stage_3__3072_ })
  );


  bsg_swap_width_p512
  mux_stage_2__mux_swap_4__swap_inst
  (
    .data_i({ data_stage_2__5119_, data_stage_2__5118_, data_stage_2__5117_, data_stage_2__5116_, data_stage_2__5115_, data_stage_2__5114_, data_stage_2__5113_, data_stage_2__5112_, data_stage_2__5111_, data_stage_2__5110_, data_stage_2__5109_, data_stage_2__5108_, data_stage_2__5107_, data_stage_2__5106_, data_stage_2__5105_, data_stage_2__5104_, data_stage_2__5103_, data_stage_2__5102_, data_stage_2__5101_, data_stage_2__5100_, data_stage_2__5099_, data_stage_2__5098_, data_stage_2__5097_, data_stage_2__5096_, data_stage_2__5095_, data_stage_2__5094_, data_stage_2__5093_, data_stage_2__5092_, data_stage_2__5091_, data_stage_2__5090_, data_stage_2__5089_, data_stage_2__5088_, data_stage_2__5087_, data_stage_2__5086_, data_stage_2__5085_, data_stage_2__5084_, data_stage_2__5083_, data_stage_2__5082_, data_stage_2__5081_, data_stage_2__5080_, data_stage_2__5079_, data_stage_2__5078_, data_stage_2__5077_, data_stage_2__5076_, data_stage_2__5075_, data_stage_2__5074_, data_stage_2__5073_, data_stage_2__5072_, data_stage_2__5071_, data_stage_2__5070_, data_stage_2__5069_, data_stage_2__5068_, data_stage_2__5067_, data_stage_2__5066_, data_stage_2__5065_, data_stage_2__5064_, data_stage_2__5063_, data_stage_2__5062_, data_stage_2__5061_, data_stage_2__5060_, data_stage_2__5059_, data_stage_2__5058_, data_stage_2__5057_, data_stage_2__5056_, data_stage_2__5055_, data_stage_2__5054_, data_stage_2__5053_, data_stage_2__5052_, data_stage_2__5051_, data_stage_2__5050_, data_stage_2__5049_, data_stage_2__5048_, data_stage_2__5047_, data_stage_2__5046_, data_stage_2__5045_, data_stage_2__5044_, data_stage_2__5043_, data_stage_2__5042_, data_stage_2__5041_, data_stage_2__5040_, data_stage_2__5039_, data_stage_2__5038_, data_stage_2__5037_, data_stage_2__5036_, data_stage_2__5035_, data_stage_2__5034_, data_stage_2__5033_, data_stage_2__5032_, data_stage_2__5031_, data_stage_2__5030_, data_stage_2__5029_, data_stage_2__5028_, data_stage_2__5027_, data_stage_2__5026_, data_stage_2__5025_, data_stage_2__5024_, data_stage_2__5023_, data_stage_2__5022_, data_stage_2__5021_, data_stage_2__5020_, data_stage_2__5019_, data_stage_2__5018_, data_stage_2__5017_, data_stage_2__5016_, data_stage_2__5015_, data_stage_2__5014_, data_stage_2__5013_, data_stage_2__5012_, data_stage_2__5011_, data_stage_2__5010_, data_stage_2__5009_, data_stage_2__5008_, data_stage_2__5007_, data_stage_2__5006_, data_stage_2__5005_, data_stage_2__5004_, data_stage_2__5003_, data_stage_2__5002_, data_stage_2__5001_, data_stage_2__5000_, data_stage_2__4999_, data_stage_2__4998_, data_stage_2__4997_, data_stage_2__4996_, data_stage_2__4995_, data_stage_2__4994_, data_stage_2__4993_, data_stage_2__4992_, data_stage_2__4991_, data_stage_2__4990_, data_stage_2__4989_, data_stage_2__4988_, data_stage_2__4987_, data_stage_2__4986_, data_stage_2__4985_, data_stage_2__4984_, data_stage_2__4983_, data_stage_2__4982_, data_stage_2__4981_, data_stage_2__4980_, data_stage_2__4979_, data_stage_2__4978_, data_stage_2__4977_, data_stage_2__4976_, data_stage_2__4975_, data_stage_2__4974_, data_stage_2__4973_, data_stage_2__4972_, data_stage_2__4971_, data_stage_2__4970_, data_stage_2__4969_, data_stage_2__4968_, data_stage_2__4967_, data_stage_2__4966_, data_stage_2__4965_, data_stage_2__4964_, data_stage_2__4963_, data_stage_2__4962_, data_stage_2__4961_, data_stage_2__4960_, data_stage_2__4959_, data_stage_2__4958_, data_stage_2__4957_, data_stage_2__4956_, data_stage_2__4955_, data_stage_2__4954_, data_stage_2__4953_, data_stage_2__4952_, data_stage_2__4951_, data_stage_2__4950_, data_stage_2__4949_, data_stage_2__4948_, data_stage_2__4947_, data_stage_2__4946_, data_stage_2__4945_, data_stage_2__4944_, data_stage_2__4943_, data_stage_2__4942_, data_stage_2__4941_, data_stage_2__4940_, data_stage_2__4939_, data_stage_2__4938_, data_stage_2__4937_, data_stage_2__4936_, data_stage_2__4935_, data_stage_2__4934_, data_stage_2__4933_, data_stage_2__4932_, data_stage_2__4931_, data_stage_2__4930_, data_stage_2__4929_, data_stage_2__4928_, data_stage_2__4927_, data_stage_2__4926_, data_stage_2__4925_, data_stage_2__4924_, data_stage_2__4923_, data_stage_2__4922_, data_stage_2__4921_, data_stage_2__4920_, data_stage_2__4919_, data_stage_2__4918_, data_stage_2__4917_, data_stage_2__4916_, data_stage_2__4915_, data_stage_2__4914_, data_stage_2__4913_, data_stage_2__4912_, data_stage_2__4911_, data_stage_2__4910_, data_stage_2__4909_, data_stage_2__4908_, data_stage_2__4907_, data_stage_2__4906_, data_stage_2__4905_, data_stage_2__4904_, data_stage_2__4903_, data_stage_2__4902_, data_stage_2__4901_, data_stage_2__4900_, data_stage_2__4899_, data_stage_2__4898_, data_stage_2__4897_, data_stage_2__4896_, data_stage_2__4895_, data_stage_2__4894_, data_stage_2__4893_, data_stage_2__4892_, data_stage_2__4891_, data_stage_2__4890_, data_stage_2__4889_, data_stage_2__4888_, data_stage_2__4887_, data_stage_2__4886_, data_stage_2__4885_, data_stage_2__4884_, data_stage_2__4883_, data_stage_2__4882_, data_stage_2__4881_, data_stage_2__4880_, data_stage_2__4879_, data_stage_2__4878_, data_stage_2__4877_, data_stage_2__4876_, data_stage_2__4875_, data_stage_2__4874_, data_stage_2__4873_, data_stage_2__4872_, data_stage_2__4871_, data_stage_2__4870_, data_stage_2__4869_, data_stage_2__4868_, data_stage_2__4867_, data_stage_2__4866_, data_stage_2__4865_, data_stage_2__4864_, data_stage_2__4863_, data_stage_2__4862_, data_stage_2__4861_, data_stage_2__4860_, data_stage_2__4859_, data_stage_2__4858_, data_stage_2__4857_, data_stage_2__4856_, data_stage_2__4855_, data_stage_2__4854_, data_stage_2__4853_, data_stage_2__4852_, data_stage_2__4851_, data_stage_2__4850_, data_stage_2__4849_, data_stage_2__4848_, data_stage_2__4847_, data_stage_2__4846_, data_stage_2__4845_, data_stage_2__4844_, data_stage_2__4843_, data_stage_2__4842_, data_stage_2__4841_, data_stage_2__4840_, data_stage_2__4839_, data_stage_2__4838_, data_stage_2__4837_, data_stage_2__4836_, data_stage_2__4835_, data_stage_2__4834_, data_stage_2__4833_, data_stage_2__4832_, data_stage_2__4831_, data_stage_2__4830_, data_stage_2__4829_, data_stage_2__4828_, data_stage_2__4827_, data_stage_2__4826_, data_stage_2__4825_, data_stage_2__4824_, data_stage_2__4823_, data_stage_2__4822_, data_stage_2__4821_, data_stage_2__4820_, data_stage_2__4819_, data_stage_2__4818_, data_stage_2__4817_, data_stage_2__4816_, data_stage_2__4815_, data_stage_2__4814_, data_stage_2__4813_, data_stage_2__4812_, data_stage_2__4811_, data_stage_2__4810_, data_stage_2__4809_, data_stage_2__4808_, data_stage_2__4807_, data_stage_2__4806_, data_stage_2__4805_, data_stage_2__4804_, data_stage_2__4803_, data_stage_2__4802_, data_stage_2__4801_, data_stage_2__4800_, data_stage_2__4799_, data_stage_2__4798_, data_stage_2__4797_, data_stage_2__4796_, data_stage_2__4795_, data_stage_2__4794_, data_stage_2__4793_, data_stage_2__4792_, data_stage_2__4791_, data_stage_2__4790_, data_stage_2__4789_, data_stage_2__4788_, data_stage_2__4787_, data_stage_2__4786_, data_stage_2__4785_, data_stage_2__4784_, data_stage_2__4783_, data_stage_2__4782_, data_stage_2__4781_, data_stage_2__4780_, data_stage_2__4779_, data_stage_2__4778_, data_stage_2__4777_, data_stage_2__4776_, data_stage_2__4775_, data_stage_2__4774_, data_stage_2__4773_, data_stage_2__4772_, data_stage_2__4771_, data_stage_2__4770_, data_stage_2__4769_, data_stage_2__4768_, data_stage_2__4767_, data_stage_2__4766_, data_stage_2__4765_, data_stage_2__4764_, data_stage_2__4763_, data_stage_2__4762_, data_stage_2__4761_, data_stage_2__4760_, data_stage_2__4759_, data_stage_2__4758_, data_stage_2__4757_, data_stage_2__4756_, data_stage_2__4755_, data_stage_2__4754_, data_stage_2__4753_, data_stage_2__4752_, data_stage_2__4751_, data_stage_2__4750_, data_stage_2__4749_, data_stage_2__4748_, data_stage_2__4747_, data_stage_2__4746_, data_stage_2__4745_, data_stage_2__4744_, data_stage_2__4743_, data_stage_2__4742_, data_stage_2__4741_, data_stage_2__4740_, data_stage_2__4739_, data_stage_2__4738_, data_stage_2__4737_, data_stage_2__4736_, data_stage_2__4735_, data_stage_2__4734_, data_stage_2__4733_, data_stage_2__4732_, data_stage_2__4731_, data_stage_2__4730_, data_stage_2__4729_, data_stage_2__4728_, data_stage_2__4727_, data_stage_2__4726_, data_stage_2__4725_, data_stage_2__4724_, data_stage_2__4723_, data_stage_2__4722_, data_stage_2__4721_, data_stage_2__4720_, data_stage_2__4719_, data_stage_2__4718_, data_stage_2__4717_, data_stage_2__4716_, data_stage_2__4715_, data_stage_2__4714_, data_stage_2__4713_, data_stage_2__4712_, data_stage_2__4711_, data_stage_2__4710_, data_stage_2__4709_, data_stage_2__4708_, data_stage_2__4707_, data_stage_2__4706_, data_stage_2__4705_, data_stage_2__4704_, data_stage_2__4703_, data_stage_2__4702_, data_stage_2__4701_, data_stage_2__4700_, data_stage_2__4699_, data_stage_2__4698_, data_stage_2__4697_, data_stage_2__4696_, data_stage_2__4695_, data_stage_2__4694_, data_stage_2__4693_, data_stage_2__4692_, data_stage_2__4691_, data_stage_2__4690_, data_stage_2__4689_, data_stage_2__4688_, data_stage_2__4687_, data_stage_2__4686_, data_stage_2__4685_, data_stage_2__4684_, data_stage_2__4683_, data_stage_2__4682_, data_stage_2__4681_, data_stage_2__4680_, data_stage_2__4679_, data_stage_2__4678_, data_stage_2__4677_, data_stage_2__4676_, data_stage_2__4675_, data_stage_2__4674_, data_stage_2__4673_, data_stage_2__4672_, data_stage_2__4671_, data_stage_2__4670_, data_stage_2__4669_, data_stage_2__4668_, data_stage_2__4667_, data_stage_2__4666_, data_stage_2__4665_, data_stage_2__4664_, data_stage_2__4663_, data_stage_2__4662_, data_stage_2__4661_, data_stage_2__4660_, data_stage_2__4659_, data_stage_2__4658_, data_stage_2__4657_, data_stage_2__4656_, data_stage_2__4655_, data_stage_2__4654_, data_stage_2__4653_, data_stage_2__4652_, data_stage_2__4651_, data_stage_2__4650_, data_stage_2__4649_, data_stage_2__4648_, data_stage_2__4647_, data_stage_2__4646_, data_stage_2__4645_, data_stage_2__4644_, data_stage_2__4643_, data_stage_2__4642_, data_stage_2__4641_, data_stage_2__4640_, data_stage_2__4639_, data_stage_2__4638_, data_stage_2__4637_, data_stage_2__4636_, data_stage_2__4635_, data_stage_2__4634_, data_stage_2__4633_, data_stage_2__4632_, data_stage_2__4631_, data_stage_2__4630_, data_stage_2__4629_, data_stage_2__4628_, data_stage_2__4627_, data_stage_2__4626_, data_stage_2__4625_, data_stage_2__4624_, data_stage_2__4623_, data_stage_2__4622_, data_stage_2__4621_, data_stage_2__4620_, data_stage_2__4619_, data_stage_2__4618_, data_stage_2__4617_, data_stage_2__4616_, data_stage_2__4615_, data_stage_2__4614_, data_stage_2__4613_, data_stage_2__4612_, data_stage_2__4611_, data_stage_2__4610_, data_stage_2__4609_, data_stage_2__4608_, data_stage_2__4607_, data_stage_2__4606_, data_stage_2__4605_, data_stage_2__4604_, data_stage_2__4603_, data_stage_2__4602_, data_stage_2__4601_, data_stage_2__4600_, data_stage_2__4599_, data_stage_2__4598_, data_stage_2__4597_, data_stage_2__4596_, data_stage_2__4595_, data_stage_2__4594_, data_stage_2__4593_, data_stage_2__4592_, data_stage_2__4591_, data_stage_2__4590_, data_stage_2__4589_, data_stage_2__4588_, data_stage_2__4587_, data_stage_2__4586_, data_stage_2__4585_, data_stage_2__4584_, data_stage_2__4583_, data_stage_2__4582_, data_stage_2__4581_, data_stage_2__4580_, data_stage_2__4579_, data_stage_2__4578_, data_stage_2__4577_, data_stage_2__4576_, data_stage_2__4575_, data_stage_2__4574_, data_stage_2__4573_, data_stage_2__4572_, data_stage_2__4571_, data_stage_2__4570_, data_stage_2__4569_, data_stage_2__4568_, data_stage_2__4567_, data_stage_2__4566_, data_stage_2__4565_, data_stage_2__4564_, data_stage_2__4563_, data_stage_2__4562_, data_stage_2__4561_, data_stage_2__4560_, data_stage_2__4559_, data_stage_2__4558_, data_stage_2__4557_, data_stage_2__4556_, data_stage_2__4555_, data_stage_2__4554_, data_stage_2__4553_, data_stage_2__4552_, data_stage_2__4551_, data_stage_2__4550_, data_stage_2__4549_, data_stage_2__4548_, data_stage_2__4547_, data_stage_2__4546_, data_stage_2__4545_, data_stage_2__4544_, data_stage_2__4543_, data_stage_2__4542_, data_stage_2__4541_, data_stage_2__4540_, data_stage_2__4539_, data_stage_2__4538_, data_stage_2__4537_, data_stage_2__4536_, data_stage_2__4535_, data_stage_2__4534_, data_stage_2__4533_, data_stage_2__4532_, data_stage_2__4531_, data_stage_2__4530_, data_stage_2__4529_, data_stage_2__4528_, data_stage_2__4527_, data_stage_2__4526_, data_stage_2__4525_, data_stage_2__4524_, data_stage_2__4523_, data_stage_2__4522_, data_stage_2__4521_, data_stage_2__4520_, data_stage_2__4519_, data_stage_2__4518_, data_stage_2__4517_, data_stage_2__4516_, data_stage_2__4515_, data_stage_2__4514_, data_stage_2__4513_, data_stage_2__4512_, data_stage_2__4511_, data_stage_2__4510_, data_stage_2__4509_, data_stage_2__4508_, data_stage_2__4507_, data_stage_2__4506_, data_stage_2__4505_, data_stage_2__4504_, data_stage_2__4503_, data_stage_2__4502_, data_stage_2__4501_, data_stage_2__4500_, data_stage_2__4499_, data_stage_2__4498_, data_stage_2__4497_, data_stage_2__4496_, data_stage_2__4495_, data_stage_2__4494_, data_stage_2__4493_, data_stage_2__4492_, data_stage_2__4491_, data_stage_2__4490_, data_stage_2__4489_, data_stage_2__4488_, data_stage_2__4487_, data_stage_2__4486_, data_stage_2__4485_, data_stage_2__4484_, data_stage_2__4483_, data_stage_2__4482_, data_stage_2__4481_, data_stage_2__4480_, data_stage_2__4479_, data_stage_2__4478_, data_stage_2__4477_, data_stage_2__4476_, data_stage_2__4475_, data_stage_2__4474_, data_stage_2__4473_, data_stage_2__4472_, data_stage_2__4471_, data_stage_2__4470_, data_stage_2__4469_, data_stage_2__4468_, data_stage_2__4467_, data_stage_2__4466_, data_stage_2__4465_, data_stage_2__4464_, data_stage_2__4463_, data_stage_2__4462_, data_stage_2__4461_, data_stage_2__4460_, data_stage_2__4459_, data_stage_2__4458_, data_stage_2__4457_, data_stage_2__4456_, data_stage_2__4455_, data_stage_2__4454_, data_stage_2__4453_, data_stage_2__4452_, data_stage_2__4451_, data_stage_2__4450_, data_stage_2__4449_, data_stage_2__4448_, data_stage_2__4447_, data_stage_2__4446_, data_stage_2__4445_, data_stage_2__4444_, data_stage_2__4443_, data_stage_2__4442_, data_stage_2__4441_, data_stage_2__4440_, data_stage_2__4439_, data_stage_2__4438_, data_stage_2__4437_, data_stage_2__4436_, data_stage_2__4435_, data_stage_2__4434_, data_stage_2__4433_, data_stage_2__4432_, data_stage_2__4431_, data_stage_2__4430_, data_stage_2__4429_, data_stage_2__4428_, data_stage_2__4427_, data_stage_2__4426_, data_stage_2__4425_, data_stage_2__4424_, data_stage_2__4423_, data_stage_2__4422_, data_stage_2__4421_, data_stage_2__4420_, data_stage_2__4419_, data_stage_2__4418_, data_stage_2__4417_, data_stage_2__4416_, data_stage_2__4415_, data_stage_2__4414_, data_stage_2__4413_, data_stage_2__4412_, data_stage_2__4411_, data_stage_2__4410_, data_stage_2__4409_, data_stage_2__4408_, data_stage_2__4407_, data_stage_2__4406_, data_stage_2__4405_, data_stage_2__4404_, data_stage_2__4403_, data_stage_2__4402_, data_stage_2__4401_, data_stage_2__4400_, data_stage_2__4399_, data_stage_2__4398_, data_stage_2__4397_, data_stage_2__4396_, data_stage_2__4395_, data_stage_2__4394_, data_stage_2__4393_, data_stage_2__4392_, data_stage_2__4391_, data_stage_2__4390_, data_stage_2__4389_, data_stage_2__4388_, data_stage_2__4387_, data_stage_2__4386_, data_stage_2__4385_, data_stage_2__4384_, data_stage_2__4383_, data_stage_2__4382_, data_stage_2__4381_, data_stage_2__4380_, data_stage_2__4379_, data_stage_2__4378_, data_stage_2__4377_, data_stage_2__4376_, data_stage_2__4375_, data_stage_2__4374_, data_stage_2__4373_, data_stage_2__4372_, data_stage_2__4371_, data_stage_2__4370_, data_stage_2__4369_, data_stage_2__4368_, data_stage_2__4367_, data_stage_2__4366_, data_stage_2__4365_, data_stage_2__4364_, data_stage_2__4363_, data_stage_2__4362_, data_stage_2__4361_, data_stage_2__4360_, data_stage_2__4359_, data_stage_2__4358_, data_stage_2__4357_, data_stage_2__4356_, data_stage_2__4355_, data_stage_2__4354_, data_stage_2__4353_, data_stage_2__4352_, data_stage_2__4351_, data_stage_2__4350_, data_stage_2__4349_, data_stage_2__4348_, data_stage_2__4347_, data_stage_2__4346_, data_stage_2__4345_, data_stage_2__4344_, data_stage_2__4343_, data_stage_2__4342_, data_stage_2__4341_, data_stage_2__4340_, data_stage_2__4339_, data_stage_2__4338_, data_stage_2__4337_, data_stage_2__4336_, data_stage_2__4335_, data_stage_2__4334_, data_stage_2__4333_, data_stage_2__4332_, data_stage_2__4331_, data_stage_2__4330_, data_stage_2__4329_, data_stage_2__4328_, data_stage_2__4327_, data_stage_2__4326_, data_stage_2__4325_, data_stage_2__4324_, data_stage_2__4323_, data_stage_2__4322_, data_stage_2__4321_, data_stage_2__4320_, data_stage_2__4319_, data_stage_2__4318_, data_stage_2__4317_, data_stage_2__4316_, data_stage_2__4315_, data_stage_2__4314_, data_stage_2__4313_, data_stage_2__4312_, data_stage_2__4311_, data_stage_2__4310_, data_stage_2__4309_, data_stage_2__4308_, data_stage_2__4307_, data_stage_2__4306_, data_stage_2__4305_, data_stage_2__4304_, data_stage_2__4303_, data_stage_2__4302_, data_stage_2__4301_, data_stage_2__4300_, data_stage_2__4299_, data_stage_2__4298_, data_stage_2__4297_, data_stage_2__4296_, data_stage_2__4295_, data_stage_2__4294_, data_stage_2__4293_, data_stage_2__4292_, data_stage_2__4291_, data_stage_2__4290_, data_stage_2__4289_, data_stage_2__4288_, data_stage_2__4287_, data_stage_2__4286_, data_stage_2__4285_, data_stage_2__4284_, data_stage_2__4283_, data_stage_2__4282_, data_stage_2__4281_, data_stage_2__4280_, data_stage_2__4279_, data_stage_2__4278_, data_stage_2__4277_, data_stage_2__4276_, data_stage_2__4275_, data_stage_2__4274_, data_stage_2__4273_, data_stage_2__4272_, data_stage_2__4271_, data_stage_2__4270_, data_stage_2__4269_, data_stage_2__4268_, data_stage_2__4267_, data_stage_2__4266_, data_stage_2__4265_, data_stage_2__4264_, data_stage_2__4263_, data_stage_2__4262_, data_stage_2__4261_, data_stage_2__4260_, data_stage_2__4259_, data_stage_2__4258_, data_stage_2__4257_, data_stage_2__4256_, data_stage_2__4255_, data_stage_2__4254_, data_stage_2__4253_, data_stage_2__4252_, data_stage_2__4251_, data_stage_2__4250_, data_stage_2__4249_, data_stage_2__4248_, data_stage_2__4247_, data_stage_2__4246_, data_stage_2__4245_, data_stage_2__4244_, data_stage_2__4243_, data_stage_2__4242_, data_stage_2__4241_, data_stage_2__4240_, data_stage_2__4239_, data_stage_2__4238_, data_stage_2__4237_, data_stage_2__4236_, data_stage_2__4235_, data_stage_2__4234_, data_stage_2__4233_, data_stage_2__4232_, data_stage_2__4231_, data_stage_2__4230_, data_stage_2__4229_, data_stage_2__4228_, data_stage_2__4227_, data_stage_2__4226_, data_stage_2__4225_, data_stage_2__4224_, data_stage_2__4223_, data_stage_2__4222_, data_stage_2__4221_, data_stage_2__4220_, data_stage_2__4219_, data_stage_2__4218_, data_stage_2__4217_, data_stage_2__4216_, data_stage_2__4215_, data_stage_2__4214_, data_stage_2__4213_, data_stage_2__4212_, data_stage_2__4211_, data_stage_2__4210_, data_stage_2__4209_, data_stage_2__4208_, data_stage_2__4207_, data_stage_2__4206_, data_stage_2__4205_, data_stage_2__4204_, data_stage_2__4203_, data_stage_2__4202_, data_stage_2__4201_, data_stage_2__4200_, data_stage_2__4199_, data_stage_2__4198_, data_stage_2__4197_, data_stage_2__4196_, data_stage_2__4195_, data_stage_2__4194_, data_stage_2__4193_, data_stage_2__4192_, data_stage_2__4191_, data_stage_2__4190_, data_stage_2__4189_, data_stage_2__4188_, data_stage_2__4187_, data_stage_2__4186_, data_stage_2__4185_, data_stage_2__4184_, data_stage_2__4183_, data_stage_2__4182_, data_stage_2__4181_, data_stage_2__4180_, data_stage_2__4179_, data_stage_2__4178_, data_stage_2__4177_, data_stage_2__4176_, data_stage_2__4175_, data_stage_2__4174_, data_stage_2__4173_, data_stage_2__4172_, data_stage_2__4171_, data_stage_2__4170_, data_stage_2__4169_, data_stage_2__4168_, data_stage_2__4167_, data_stage_2__4166_, data_stage_2__4165_, data_stage_2__4164_, data_stage_2__4163_, data_stage_2__4162_, data_stage_2__4161_, data_stage_2__4160_, data_stage_2__4159_, data_stage_2__4158_, data_stage_2__4157_, data_stage_2__4156_, data_stage_2__4155_, data_stage_2__4154_, data_stage_2__4153_, data_stage_2__4152_, data_stage_2__4151_, data_stage_2__4150_, data_stage_2__4149_, data_stage_2__4148_, data_stage_2__4147_, data_stage_2__4146_, data_stage_2__4145_, data_stage_2__4144_, data_stage_2__4143_, data_stage_2__4142_, data_stage_2__4141_, data_stage_2__4140_, data_stage_2__4139_, data_stage_2__4138_, data_stage_2__4137_, data_stage_2__4136_, data_stage_2__4135_, data_stage_2__4134_, data_stage_2__4133_, data_stage_2__4132_, data_stage_2__4131_, data_stage_2__4130_, data_stage_2__4129_, data_stage_2__4128_, data_stage_2__4127_, data_stage_2__4126_, data_stage_2__4125_, data_stage_2__4124_, data_stage_2__4123_, data_stage_2__4122_, data_stage_2__4121_, data_stage_2__4120_, data_stage_2__4119_, data_stage_2__4118_, data_stage_2__4117_, data_stage_2__4116_, data_stage_2__4115_, data_stage_2__4114_, data_stage_2__4113_, data_stage_2__4112_, data_stage_2__4111_, data_stage_2__4110_, data_stage_2__4109_, data_stage_2__4108_, data_stage_2__4107_, data_stage_2__4106_, data_stage_2__4105_, data_stage_2__4104_, data_stage_2__4103_, data_stage_2__4102_, data_stage_2__4101_, data_stage_2__4100_, data_stage_2__4099_, data_stage_2__4098_, data_stage_2__4097_, data_stage_2__4096_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__5119_, data_stage_3__5118_, data_stage_3__5117_, data_stage_3__5116_, data_stage_3__5115_, data_stage_3__5114_, data_stage_3__5113_, data_stage_3__5112_, data_stage_3__5111_, data_stage_3__5110_, data_stage_3__5109_, data_stage_3__5108_, data_stage_3__5107_, data_stage_3__5106_, data_stage_3__5105_, data_stage_3__5104_, data_stage_3__5103_, data_stage_3__5102_, data_stage_3__5101_, data_stage_3__5100_, data_stage_3__5099_, data_stage_3__5098_, data_stage_3__5097_, data_stage_3__5096_, data_stage_3__5095_, data_stage_3__5094_, data_stage_3__5093_, data_stage_3__5092_, data_stage_3__5091_, data_stage_3__5090_, data_stage_3__5089_, data_stage_3__5088_, data_stage_3__5087_, data_stage_3__5086_, data_stage_3__5085_, data_stage_3__5084_, data_stage_3__5083_, data_stage_3__5082_, data_stage_3__5081_, data_stage_3__5080_, data_stage_3__5079_, data_stage_3__5078_, data_stage_3__5077_, data_stage_3__5076_, data_stage_3__5075_, data_stage_3__5074_, data_stage_3__5073_, data_stage_3__5072_, data_stage_3__5071_, data_stage_3__5070_, data_stage_3__5069_, data_stage_3__5068_, data_stage_3__5067_, data_stage_3__5066_, data_stage_3__5065_, data_stage_3__5064_, data_stage_3__5063_, data_stage_3__5062_, data_stage_3__5061_, data_stage_3__5060_, data_stage_3__5059_, data_stage_3__5058_, data_stage_3__5057_, data_stage_3__5056_, data_stage_3__5055_, data_stage_3__5054_, data_stage_3__5053_, data_stage_3__5052_, data_stage_3__5051_, data_stage_3__5050_, data_stage_3__5049_, data_stage_3__5048_, data_stage_3__5047_, data_stage_3__5046_, data_stage_3__5045_, data_stage_3__5044_, data_stage_3__5043_, data_stage_3__5042_, data_stage_3__5041_, data_stage_3__5040_, data_stage_3__5039_, data_stage_3__5038_, data_stage_3__5037_, data_stage_3__5036_, data_stage_3__5035_, data_stage_3__5034_, data_stage_3__5033_, data_stage_3__5032_, data_stage_3__5031_, data_stage_3__5030_, data_stage_3__5029_, data_stage_3__5028_, data_stage_3__5027_, data_stage_3__5026_, data_stage_3__5025_, data_stage_3__5024_, data_stage_3__5023_, data_stage_3__5022_, data_stage_3__5021_, data_stage_3__5020_, data_stage_3__5019_, data_stage_3__5018_, data_stage_3__5017_, data_stage_3__5016_, data_stage_3__5015_, data_stage_3__5014_, data_stage_3__5013_, data_stage_3__5012_, data_stage_3__5011_, data_stage_3__5010_, data_stage_3__5009_, data_stage_3__5008_, data_stage_3__5007_, data_stage_3__5006_, data_stage_3__5005_, data_stage_3__5004_, data_stage_3__5003_, data_stage_3__5002_, data_stage_3__5001_, data_stage_3__5000_, data_stage_3__4999_, data_stage_3__4998_, data_stage_3__4997_, data_stage_3__4996_, data_stage_3__4995_, data_stage_3__4994_, data_stage_3__4993_, data_stage_3__4992_, data_stage_3__4991_, data_stage_3__4990_, data_stage_3__4989_, data_stage_3__4988_, data_stage_3__4987_, data_stage_3__4986_, data_stage_3__4985_, data_stage_3__4984_, data_stage_3__4983_, data_stage_3__4982_, data_stage_3__4981_, data_stage_3__4980_, data_stage_3__4979_, data_stage_3__4978_, data_stage_3__4977_, data_stage_3__4976_, data_stage_3__4975_, data_stage_3__4974_, data_stage_3__4973_, data_stage_3__4972_, data_stage_3__4971_, data_stage_3__4970_, data_stage_3__4969_, data_stage_3__4968_, data_stage_3__4967_, data_stage_3__4966_, data_stage_3__4965_, data_stage_3__4964_, data_stage_3__4963_, data_stage_3__4962_, data_stage_3__4961_, data_stage_3__4960_, data_stage_3__4959_, data_stage_3__4958_, data_stage_3__4957_, data_stage_3__4956_, data_stage_3__4955_, data_stage_3__4954_, data_stage_3__4953_, data_stage_3__4952_, data_stage_3__4951_, data_stage_3__4950_, data_stage_3__4949_, data_stage_3__4948_, data_stage_3__4947_, data_stage_3__4946_, data_stage_3__4945_, data_stage_3__4944_, data_stage_3__4943_, data_stage_3__4942_, data_stage_3__4941_, data_stage_3__4940_, data_stage_3__4939_, data_stage_3__4938_, data_stage_3__4937_, data_stage_3__4936_, data_stage_3__4935_, data_stage_3__4934_, data_stage_3__4933_, data_stage_3__4932_, data_stage_3__4931_, data_stage_3__4930_, data_stage_3__4929_, data_stage_3__4928_, data_stage_3__4927_, data_stage_3__4926_, data_stage_3__4925_, data_stage_3__4924_, data_stage_3__4923_, data_stage_3__4922_, data_stage_3__4921_, data_stage_3__4920_, data_stage_3__4919_, data_stage_3__4918_, data_stage_3__4917_, data_stage_3__4916_, data_stage_3__4915_, data_stage_3__4914_, data_stage_3__4913_, data_stage_3__4912_, data_stage_3__4911_, data_stage_3__4910_, data_stage_3__4909_, data_stage_3__4908_, data_stage_3__4907_, data_stage_3__4906_, data_stage_3__4905_, data_stage_3__4904_, data_stage_3__4903_, data_stage_3__4902_, data_stage_3__4901_, data_stage_3__4900_, data_stage_3__4899_, data_stage_3__4898_, data_stage_3__4897_, data_stage_3__4896_, data_stage_3__4895_, data_stage_3__4894_, data_stage_3__4893_, data_stage_3__4892_, data_stage_3__4891_, data_stage_3__4890_, data_stage_3__4889_, data_stage_3__4888_, data_stage_3__4887_, data_stage_3__4886_, data_stage_3__4885_, data_stage_3__4884_, data_stage_3__4883_, data_stage_3__4882_, data_stage_3__4881_, data_stage_3__4880_, data_stage_3__4879_, data_stage_3__4878_, data_stage_3__4877_, data_stage_3__4876_, data_stage_3__4875_, data_stage_3__4874_, data_stage_3__4873_, data_stage_3__4872_, data_stage_3__4871_, data_stage_3__4870_, data_stage_3__4869_, data_stage_3__4868_, data_stage_3__4867_, data_stage_3__4866_, data_stage_3__4865_, data_stage_3__4864_, data_stage_3__4863_, data_stage_3__4862_, data_stage_3__4861_, data_stage_3__4860_, data_stage_3__4859_, data_stage_3__4858_, data_stage_3__4857_, data_stage_3__4856_, data_stage_3__4855_, data_stage_3__4854_, data_stage_3__4853_, data_stage_3__4852_, data_stage_3__4851_, data_stage_3__4850_, data_stage_3__4849_, data_stage_3__4848_, data_stage_3__4847_, data_stage_3__4846_, data_stage_3__4845_, data_stage_3__4844_, data_stage_3__4843_, data_stage_3__4842_, data_stage_3__4841_, data_stage_3__4840_, data_stage_3__4839_, data_stage_3__4838_, data_stage_3__4837_, data_stage_3__4836_, data_stage_3__4835_, data_stage_3__4834_, data_stage_3__4833_, data_stage_3__4832_, data_stage_3__4831_, data_stage_3__4830_, data_stage_3__4829_, data_stage_3__4828_, data_stage_3__4827_, data_stage_3__4826_, data_stage_3__4825_, data_stage_3__4824_, data_stage_3__4823_, data_stage_3__4822_, data_stage_3__4821_, data_stage_3__4820_, data_stage_3__4819_, data_stage_3__4818_, data_stage_3__4817_, data_stage_3__4816_, data_stage_3__4815_, data_stage_3__4814_, data_stage_3__4813_, data_stage_3__4812_, data_stage_3__4811_, data_stage_3__4810_, data_stage_3__4809_, data_stage_3__4808_, data_stage_3__4807_, data_stage_3__4806_, data_stage_3__4805_, data_stage_3__4804_, data_stage_3__4803_, data_stage_3__4802_, data_stage_3__4801_, data_stage_3__4800_, data_stage_3__4799_, data_stage_3__4798_, data_stage_3__4797_, data_stage_3__4796_, data_stage_3__4795_, data_stage_3__4794_, data_stage_3__4793_, data_stage_3__4792_, data_stage_3__4791_, data_stage_3__4790_, data_stage_3__4789_, data_stage_3__4788_, data_stage_3__4787_, data_stage_3__4786_, data_stage_3__4785_, data_stage_3__4784_, data_stage_3__4783_, data_stage_3__4782_, data_stage_3__4781_, data_stage_3__4780_, data_stage_3__4779_, data_stage_3__4778_, data_stage_3__4777_, data_stage_3__4776_, data_stage_3__4775_, data_stage_3__4774_, data_stage_3__4773_, data_stage_3__4772_, data_stage_3__4771_, data_stage_3__4770_, data_stage_3__4769_, data_stage_3__4768_, data_stage_3__4767_, data_stage_3__4766_, data_stage_3__4765_, data_stage_3__4764_, data_stage_3__4763_, data_stage_3__4762_, data_stage_3__4761_, data_stage_3__4760_, data_stage_3__4759_, data_stage_3__4758_, data_stage_3__4757_, data_stage_3__4756_, data_stage_3__4755_, data_stage_3__4754_, data_stage_3__4753_, data_stage_3__4752_, data_stage_3__4751_, data_stage_3__4750_, data_stage_3__4749_, data_stage_3__4748_, data_stage_3__4747_, data_stage_3__4746_, data_stage_3__4745_, data_stage_3__4744_, data_stage_3__4743_, data_stage_3__4742_, data_stage_3__4741_, data_stage_3__4740_, data_stage_3__4739_, data_stage_3__4738_, data_stage_3__4737_, data_stage_3__4736_, data_stage_3__4735_, data_stage_3__4734_, data_stage_3__4733_, data_stage_3__4732_, data_stage_3__4731_, data_stage_3__4730_, data_stage_3__4729_, data_stage_3__4728_, data_stage_3__4727_, data_stage_3__4726_, data_stage_3__4725_, data_stage_3__4724_, data_stage_3__4723_, data_stage_3__4722_, data_stage_3__4721_, data_stage_3__4720_, data_stage_3__4719_, data_stage_3__4718_, data_stage_3__4717_, data_stage_3__4716_, data_stage_3__4715_, data_stage_3__4714_, data_stage_3__4713_, data_stage_3__4712_, data_stage_3__4711_, data_stage_3__4710_, data_stage_3__4709_, data_stage_3__4708_, data_stage_3__4707_, data_stage_3__4706_, data_stage_3__4705_, data_stage_3__4704_, data_stage_3__4703_, data_stage_3__4702_, data_stage_3__4701_, data_stage_3__4700_, data_stage_3__4699_, data_stage_3__4698_, data_stage_3__4697_, data_stage_3__4696_, data_stage_3__4695_, data_stage_3__4694_, data_stage_3__4693_, data_stage_3__4692_, data_stage_3__4691_, data_stage_3__4690_, data_stage_3__4689_, data_stage_3__4688_, data_stage_3__4687_, data_stage_3__4686_, data_stage_3__4685_, data_stage_3__4684_, data_stage_3__4683_, data_stage_3__4682_, data_stage_3__4681_, data_stage_3__4680_, data_stage_3__4679_, data_stage_3__4678_, data_stage_3__4677_, data_stage_3__4676_, data_stage_3__4675_, data_stage_3__4674_, data_stage_3__4673_, data_stage_3__4672_, data_stage_3__4671_, data_stage_3__4670_, data_stage_3__4669_, data_stage_3__4668_, data_stage_3__4667_, data_stage_3__4666_, data_stage_3__4665_, data_stage_3__4664_, data_stage_3__4663_, data_stage_3__4662_, data_stage_3__4661_, data_stage_3__4660_, data_stage_3__4659_, data_stage_3__4658_, data_stage_3__4657_, data_stage_3__4656_, data_stage_3__4655_, data_stage_3__4654_, data_stage_3__4653_, data_stage_3__4652_, data_stage_3__4651_, data_stage_3__4650_, data_stage_3__4649_, data_stage_3__4648_, data_stage_3__4647_, data_stage_3__4646_, data_stage_3__4645_, data_stage_3__4644_, data_stage_3__4643_, data_stage_3__4642_, data_stage_3__4641_, data_stage_3__4640_, data_stage_3__4639_, data_stage_3__4638_, data_stage_3__4637_, data_stage_3__4636_, data_stage_3__4635_, data_stage_3__4634_, data_stage_3__4633_, data_stage_3__4632_, data_stage_3__4631_, data_stage_3__4630_, data_stage_3__4629_, data_stage_3__4628_, data_stage_3__4627_, data_stage_3__4626_, data_stage_3__4625_, data_stage_3__4624_, data_stage_3__4623_, data_stage_3__4622_, data_stage_3__4621_, data_stage_3__4620_, data_stage_3__4619_, data_stage_3__4618_, data_stage_3__4617_, data_stage_3__4616_, data_stage_3__4615_, data_stage_3__4614_, data_stage_3__4613_, data_stage_3__4612_, data_stage_3__4611_, data_stage_3__4610_, data_stage_3__4609_, data_stage_3__4608_, data_stage_3__4607_, data_stage_3__4606_, data_stage_3__4605_, data_stage_3__4604_, data_stage_3__4603_, data_stage_3__4602_, data_stage_3__4601_, data_stage_3__4600_, data_stage_3__4599_, data_stage_3__4598_, data_stage_3__4597_, data_stage_3__4596_, data_stage_3__4595_, data_stage_3__4594_, data_stage_3__4593_, data_stage_3__4592_, data_stage_3__4591_, data_stage_3__4590_, data_stage_3__4589_, data_stage_3__4588_, data_stage_3__4587_, data_stage_3__4586_, data_stage_3__4585_, data_stage_3__4584_, data_stage_3__4583_, data_stage_3__4582_, data_stage_3__4581_, data_stage_3__4580_, data_stage_3__4579_, data_stage_3__4578_, data_stage_3__4577_, data_stage_3__4576_, data_stage_3__4575_, data_stage_3__4574_, data_stage_3__4573_, data_stage_3__4572_, data_stage_3__4571_, data_stage_3__4570_, data_stage_3__4569_, data_stage_3__4568_, data_stage_3__4567_, data_stage_3__4566_, data_stage_3__4565_, data_stage_3__4564_, data_stage_3__4563_, data_stage_3__4562_, data_stage_3__4561_, data_stage_3__4560_, data_stage_3__4559_, data_stage_3__4558_, data_stage_3__4557_, data_stage_3__4556_, data_stage_3__4555_, data_stage_3__4554_, data_stage_3__4553_, data_stage_3__4552_, data_stage_3__4551_, data_stage_3__4550_, data_stage_3__4549_, data_stage_3__4548_, data_stage_3__4547_, data_stage_3__4546_, data_stage_3__4545_, data_stage_3__4544_, data_stage_3__4543_, data_stage_3__4542_, data_stage_3__4541_, data_stage_3__4540_, data_stage_3__4539_, data_stage_3__4538_, data_stage_3__4537_, data_stage_3__4536_, data_stage_3__4535_, data_stage_3__4534_, data_stage_3__4533_, data_stage_3__4532_, data_stage_3__4531_, data_stage_3__4530_, data_stage_3__4529_, data_stage_3__4528_, data_stage_3__4527_, data_stage_3__4526_, data_stage_3__4525_, data_stage_3__4524_, data_stage_3__4523_, data_stage_3__4522_, data_stage_3__4521_, data_stage_3__4520_, data_stage_3__4519_, data_stage_3__4518_, data_stage_3__4517_, data_stage_3__4516_, data_stage_3__4515_, data_stage_3__4514_, data_stage_3__4513_, data_stage_3__4512_, data_stage_3__4511_, data_stage_3__4510_, data_stage_3__4509_, data_stage_3__4508_, data_stage_3__4507_, data_stage_3__4506_, data_stage_3__4505_, data_stage_3__4504_, data_stage_3__4503_, data_stage_3__4502_, data_stage_3__4501_, data_stage_3__4500_, data_stage_3__4499_, data_stage_3__4498_, data_stage_3__4497_, data_stage_3__4496_, data_stage_3__4495_, data_stage_3__4494_, data_stage_3__4493_, data_stage_3__4492_, data_stage_3__4491_, data_stage_3__4490_, data_stage_3__4489_, data_stage_3__4488_, data_stage_3__4487_, data_stage_3__4486_, data_stage_3__4485_, data_stage_3__4484_, data_stage_3__4483_, data_stage_3__4482_, data_stage_3__4481_, data_stage_3__4480_, data_stage_3__4479_, data_stage_3__4478_, data_stage_3__4477_, data_stage_3__4476_, data_stage_3__4475_, data_stage_3__4474_, data_stage_3__4473_, data_stage_3__4472_, data_stage_3__4471_, data_stage_3__4470_, data_stage_3__4469_, data_stage_3__4468_, data_stage_3__4467_, data_stage_3__4466_, data_stage_3__4465_, data_stage_3__4464_, data_stage_3__4463_, data_stage_3__4462_, data_stage_3__4461_, data_stage_3__4460_, data_stage_3__4459_, data_stage_3__4458_, data_stage_3__4457_, data_stage_3__4456_, data_stage_3__4455_, data_stage_3__4454_, data_stage_3__4453_, data_stage_3__4452_, data_stage_3__4451_, data_stage_3__4450_, data_stage_3__4449_, data_stage_3__4448_, data_stage_3__4447_, data_stage_3__4446_, data_stage_3__4445_, data_stage_3__4444_, data_stage_3__4443_, data_stage_3__4442_, data_stage_3__4441_, data_stage_3__4440_, data_stage_3__4439_, data_stage_3__4438_, data_stage_3__4437_, data_stage_3__4436_, data_stage_3__4435_, data_stage_3__4434_, data_stage_3__4433_, data_stage_3__4432_, data_stage_3__4431_, data_stage_3__4430_, data_stage_3__4429_, data_stage_3__4428_, data_stage_3__4427_, data_stage_3__4426_, data_stage_3__4425_, data_stage_3__4424_, data_stage_3__4423_, data_stage_3__4422_, data_stage_3__4421_, data_stage_3__4420_, data_stage_3__4419_, data_stage_3__4418_, data_stage_3__4417_, data_stage_3__4416_, data_stage_3__4415_, data_stage_3__4414_, data_stage_3__4413_, data_stage_3__4412_, data_stage_3__4411_, data_stage_3__4410_, data_stage_3__4409_, data_stage_3__4408_, data_stage_3__4407_, data_stage_3__4406_, data_stage_3__4405_, data_stage_3__4404_, data_stage_3__4403_, data_stage_3__4402_, data_stage_3__4401_, data_stage_3__4400_, data_stage_3__4399_, data_stage_3__4398_, data_stage_3__4397_, data_stage_3__4396_, data_stage_3__4395_, data_stage_3__4394_, data_stage_3__4393_, data_stage_3__4392_, data_stage_3__4391_, data_stage_3__4390_, data_stage_3__4389_, data_stage_3__4388_, data_stage_3__4387_, data_stage_3__4386_, data_stage_3__4385_, data_stage_3__4384_, data_stage_3__4383_, data_stage_3__4382_, data_stage_3__4381_, data_stage_3__4380_, data_stage_3__4379_, data_stage_3__4378_, data_stage_3__4377_, data_stage_3__4376_, data_stage_3__4375_, data_stage_3__4374_, data_stage_3__4373_, data_stage_3__4372_, data_stage_3__4371_, data_stage_3__4370_, data_stage_3__4369_, data_stage_3__4368_, data_stage_3__4367_, data_stage_3__4366_, data_stage_3__4365_, data_stage_3__4364_, data_stage_3__4363_, data_stage_3__4362_, data_stage_3__4361_, data_stage_3__4360_, data_stage_3__4359_, data_stage_3__4358_, data_stage_3__4357_, data_stage_3__4356_, data_stage_3__4355_, data_stage_3__4354_, data_stage_3__4353_, data_stage_3__4352_, data_stage_3__4351_, data_stage_3__4350_, data_stage_3__4349_, data_stage_3__4348_, data_stage_3__4347_, data_stage_3__4346_, data_stage_3__4345_, data_stage_3__4344_, data_stage_3__4343_, data_stage_3__4342_, data_stage_3__4341_, data_stage_3__4340_, data_stage_3__4339_, data_stage_3__4338_, data_stage_3__4337_, data_stage_3__4336_, data_stage_3__4335_, data_stage_3__4334_, data_stage_3__4333_, data_stage_3__4332_, data_stage_3__4331_, data_stage_3__4330_, data_stage_3__4329_, data_stage_3__4328_, data_stage_3__4327_, data_stage_3__4326_, data_stage_3__4325_, data_stage_3__4324_, data_stage_3__4323_, data_stage_3__4322_, data_stage_3__4321_, data_stage_3__4320_, data_stage_3__4319_, data_stage_3__4318_, data_stage_3__4317_, data_stage_3__4316_, data_stage_3__4315_, data_stage_3__4314_, data_stage_3__4313_, data_stage_3__4312_, data_stage_3__4311_, data_stage_3__4310_, data_stage_3__4309_, data_stage_3__4308_, data_stage_3__4307_, data_stage_3__4306_, data_stage_3__4305_, data_stage_3__4304_, data_stage_3__4303_, data_stage_3__4302_, data_stage_3__4301_, data_stage_3__4300_, data_stage_3__4299_, data_stage_3__4298_, data_stage_3__4297_, data_stage_3__4296_, data_stage_3__4295_, data_stage_3__4294_, data_stage_3__4293_, data_stage_3__4292_, data_stage_3__4291_, data_stage_3__4290_, data_stage_3__4289_, data_stage_3__4288_, data_stage_3__4287_, data_stage_3__4286_, data_stage_3__4285_, data_stage_3__4284_, data_stage_3__4283_, data_stage_3__4282_, data_stage_3__4281_, data_stage_3__4280_, data_stage_3__4279_, data_stage_3__4278_, data_stage_3__4277_, data_stage_3__4276_, data_stage_3__4275_, data_stage_3__4274_, data_stage_3__4273_, data_stage_3__4272_, data_stage_3__4271_, data_stage_3__4270_, data_stage_3__4269_, data_stage_3__4268_, data_stage_3__4267_, data_stage_3__4266_, data_stage_3__4265_, data_stage_3__4264_, data_stage_3__4263_, data_stage_3__4262_, data_stage_3__4261_, data_stage_3__4260_, data_stage_3__4259_, data_stage_3__4258_, data_stage_3__4257_, data_stage_3__4256_, data_stage_3__4255_, data_stage_3__4254_, data_stage_3__4253_, data_stage_3__4252_, data_stage_3__4251_, data_stage_3__4250_, data_stage_3__4249_, data_stage_3__4248_, data_stage_3__4247_, data_stage_3__4246_, data_stage_3__4245_, data_stage_3__4244_, data_stage_3__4243_, data_stage_3__4242_, data_stage_3__4241_, data_stage_3__4240_, data_stage_3__4239_, data_stage_3__4238_, data_stage_3__4237_, data_stage_3__4236_, data_stage_3__4235_, data_stage_3__4234_, data_stage_3__4233_, data_stage_3__4232_, data_stage_3__4231_, data_stage_3__4230_, data_stage_3__4229_, data_stage_3__4228_, data_stage_3__4227_, data_stage_3__4226_, data_stage_3__4225_, data_stage_3__4224_, data_stage_3__4223_, data_stage_3__4222_, data_stage_3__4221_, data_stage_3__4220_, data_stage_3__4219_, data_stage_3__4218_, data_stage_3__4217_, data_stage_3__4216_, data_stage_3__4215_, data_stage_3__4214_, data_stage_3__4213_, data_stage_3__4212_, data_stage_3__4211_, data_stage_3__4210_, data_stage_3__4209_, data_stage_3__4208_, data_stage_3__4207_, data_stage_3__4206_, data_stage_3__4205_, data_stage_3__4204_, data_stage_3__4203_, data_stage_3__4202_, data_stage_3__4201_, data_stage_3__4200_, data_stage_3__4199_, data_stage_3__4198_, data_stage_3__4197_, data_stage_3__4196_, data_stage_3__4195_, data_stage_3__4194_, data_stage_3__4193_, data_stage_3__4192_, data_stage_3__4191_, data_stage_3__4190_, data_stage_3__4189_, data_stage_3__4188_, data_stage_3__4187_, data_stage_3__4186_, data_stage_3__4185_, data_stage_3__4184_, data_stage_3__4183_, data_stage_3__4182_, data_stage_3__4181_, data_stage_3__4180_, data_stage_3__4179_, data_stage_3__4178_, data_stage_3__4177_, data_stage_3__4176_, data_stage_3__4175_, data_stage_3__4174_, data_stage_3__4173_, data_stage_3__4172_, data_stage_3__4171_, data_stage_3__4170_, data_stage_3__4169_, data_stage_3__4168_, data_stage_3__4167_, data_stage_3__4166_, data_stage_3__4165_, data_stage_3__4164_, data_stage_3__4163_, data_stage_3__4162_, data_stage_3__4161_, data_stage_3__4160_, data_stage_3__4159_, data_stage_3__4158_, data_stage_3__4157_, data_stage_3__4156_, data_stage_3__4155_, data_stage_3__4154_, data_stage_3__4153_, data_stage_3__4152_, data_stage_3__4151_, data_stage_3__4150_, data_stage_3__4149_, data_stage_3__4148_, data_stage_3__4147_, data_stage_3__4146_, data_stage_3__4145_, data_stage_3__4144_, data_stage_3__4143_, data_stage_3__4142_, data_stage_3__4141_, data_stage_3__4140_, data_stage_3__4139_, data_stage_3__4138_, data_stage_3__4137_, data_stage_3__4136_, data_stage_3__4135_, data_stage_3__4134_, data_stage_3__4133_, data_stage_3__4132_, data_stage_3__4131_, data_stage_3__4130_, data_stage_3__4129_, data_stage_3__4128_, data_stage_3__4127_, data_stage_3__4126_, data_stage_3__4125_, data_stage_3__4124_, data_stage_3__4123_, data_stage_3__4122_, data_stage_3__4121_, data_stage_3__4120_, data_stage_3__4119_, data_stage_3__4118_, data_stage_3__4117_, data_stage_3__4116_, data_stage_3__4115_, data_stage_3__4114_, data_stage_3__4113_, data_stage_3__4112_, data_stage_3__4111_, data_stage_3__4110_, data_stage_3__4109_, data_stage_3__4108_, data_stage_3__4107_, data_stage_3__4106_, data_stage_3__4105_, data_stage_3__4104_, data_stage_3__4103_, data_stage_3__4102_, data_stage_3__4101_, data_stage_3__4100_, data_stage_3__4099_, data_stage_3__4098_, data_stage_3__4097_, data_stage_3__4096_ })
  );


  bsg_swap_width_p512
  mux_stage_2__mux_swap_5__swap_inst
  (
    .data_i({ data_stage_2__6143_, data_stage_2__6142_, data_stage_2__6141_, data_stage_2__6140_, data_stage_2__6139_, data_stage_2__6138_, data_stage_2__6137_, data_stage_2__6136_, data_stage_2__6135_, data_stage_2__6134_, data_stage_2__6133_, data_stage_2__6132_, data_stage_2__6131_, data_stage_2__6130_, data_stage_2__6129_, data_stage_2__6128_, data_stage_2__6127_, data_stage_2__6126_, data_stage_2__6125_, data_stage_2__6124_, data_stage_2__6123_, data_stage_2__6122_, data_stage_2__6121_, data_stage_2__6120_, data_stage_2__6119_, data_stage_2__6118_, data_stage_2__6117_, data_stage_2__6116_, data_stage_2__6115_, data_stage_2__6114_, data_stage_2__6113_, data_stage_2__6112_, data_stage_2__6111_, data_stage_2__6110_, data_stage_2__6109_, data_stage_2__6108_, data_stage_2__6107_, data_stage_2__6106_, data_stage_2__6105_, data_stage_2__6104_, data_stage_2__6103_, data_stage_2__6102_, data_stage_2__6101_, data_stage_2__6100_, data_stage_2__6099_, data_stage_2__6098_, data_stage_2__6097_, data_stage_2__6096_, data_stage_2__6095_, data_stage_2__6094_, data_stage_2__6093_, data_stage_2__6092_, data_stage_2__6091_, data_stage_2__6090_, data_stage_2__6089_, data_stage_2__6088_, data_stage_2__6087_, data_stage_2__6086_, data_stage_2__6085_, data_stage_2__6084_, data_stage_2__6083_, data_stage_2__6082_, data_stage_2__6081_, data_stage_2__6080_, data_stage_2__6079_, data_stage_2__6078_, data_stage_2__6077_, data_stage_2__6076_, data_stage_2__6075_, data_stage_2__6074_, data_stage_2__6073_, data_stage_2__6072_, data_stage_2__6071_, data_stage_2__6070_, data_stage_2__6069_, data_stage_2__6068_, data_stage_2__6067_, data_stage_2__6066_, data_stage_2__6065_, data_stage_2__6064_, data_stage_2__6063_, data_stage_2__6062_, data_stage_2__6061_, data_stage_2__6060_, data_stage_2__6059_, data_stage_2__6058_, data_stage_2__6057_, data_stage_2__6056_, data_stage_2__6055_, data_stage_2__6054_, data_stage_2__6053_, data_stage_2__6052_, data_stage_2__6051_, data_stage_2__6050_, data_stage_2__6049_, data_stage_2__6048_, data_stage_2__6047_, data_stage_2__6046_, data_stage_2__6045_, data_stage_2__6044_, data_stage_2__6043_, data_stage_2__6042_, data_stage_2__6041_, data_stage_2__6040_, data_stage_2__6039_, data_stage_2__6038_, data_stage_2__6037_, data_stage_2__6036_, data_stage_2__6035_, data_stage_2__6034_, data_stage_2__6033_, data_stage_2__6032_, data_stage_2__6031_, data_stage_2__6030_, data_stage_2__6029_, data_stage_2__6028_, data_stage_2__6027_, data_stage_2__6026_, data_stage_2__6025_, data_stage_2__6024_, data_stage_2__6023_, data_stage_2__6022_, data_stage_2__6021_, data_stage_2__6020_, data_stage_2__6019_, data_stage_2__6018_, data_stage_2__6017_, data_stage_2__6016_, data_stage_2__6015_, data_stage_2__6014_, data_stage_2__6013_, data_stage_2__6012_, data_stage_2__6011_, data_stage_2__6010_, data_stage_2__6009_, data_stage_2__6008_, data_stage_2__6007_, data_stage_2__6006_, data_stage_2__6005_, data_stage_2__6004_, data_stage_2__6003_, data_stage_2__6002_, data_stage_2__6001_, data_stage_2__6000_, data_stage_2__5999_, data_stage_2__5998_, data_stage_2__5997_, data_stage_2__5996_, data_stage_2__5995_, data_stage_2__5994_, data_stage_2__5993_, data_stage_2__5992_, data_stage_2__5991_, data_stage_2__5990_, data_stage_2__5989_, data_stage_2__5988_, data_stage_2__5987_, data_stage_2__5986_, data_stage_2__5985_, data_stage_2__5984_, data_stage_2__5983_, data_stage_2__5982_, data_stage_2__5981_, data_stage_2__5980_, data_stage_2__5979_, data_stage_2__5978_, data_stage_2__5977_, data_stage_2__5976_, data_stage_2__5975_, data_stage_2__5974_, data_stage_2__5973_, data_stage_2__5972_, data_stage_2__5971_, data_stage_2__5970_, data_stage_2__5969_, data_stage_2__5968_, data_stage_2__5967_, data_stage_2__5966_, data_stage_2__5965_, data_stage_2__5964_, data_stage_2__5963_, data_stage_2__5962_, data_stage_2__5961_, data_stage_2__5960_, data_stage_2__5959_, data_stage_2__5958_, data_stage_2__5957_, data_stage_2__5956_, data_stage_2__5955_, data_stage_2__5954_, data_stage_2__5953_, data_stage_2__5952_, data_stage_2__5951_, data_stage_2__5950_, data_stage_2__5949_, data_stage_2__5948_, data_stage_2__5947_, data_stage_2__5946_, data_stage_2__5945_, data_stage_2__5944_, data_stage_2__5943_, data_stage_2__5942_, data_stage_2__5941_, data_stage_2__5940_, data_stage_2__5939_, data_stage_2__5938_, data_stage_2__5937_, data_stage_2__5936_, data_stage_2__5935_, data_stage_2__5934_, data_stage_2__5933_, data_stage_2__5932_, data_stage_2__5931_, data_stage_2__5930_, data_stage_2__5929_, data_stage_2__5928_, data_stage_2__5927_, data_stage_2__5926_, data_stage_2__5925_, data_stage_2__5924_, data_stage_2__5923_, data_stage_2__5922_, data_stage_2__5921_, data_stage_2__5920_, data_stage_2__5919_, data_stage_2__5918_, data_stage_2__5917_, data_stage_2__5916_, data_stage_2__5915_, data_stage_2__5914_, data_stage_2__5913_, data_stage_2__5912_, data_stage_2__5911_, data_stage_2__5910_, data_stage_2__5909_, data_stage_2__5908_, data_stage_2__5907_, data_stage_2__5906_, data_stage_2__5905_, data_stage_2__5904_, data_stage_2__5903_, data_stage_2__5902_, data_stage_2__5901_, data_stage_2__5900_, data_stage_2__5899_, data_stage_2__5898_, data_stage_2__5897_, data_stage_2__5896_, data_stage_2__5895_, data_stage_2__5894_, data_stage_2__5893_, data_stage_2__5892_, data_stage_2__5891_, data_stage_2__5890_, data_stage_2__5889_, data_stage_2__5888_, data_stage_2__5887_, data_stage_2__5886_, data_stage_2__5885_, data_stage_2__5884_, data_stage_2__5883_, data_stage_2__5882_, data_stage_2__5881_, data_stage_2__5880_, data_stage_2__5879_, data_stage_2__5878_, data_stage_2__5877_, data_stage_2__5876_, data_stage_2__5875_, data_stage_2__5874_, data_stage_2__5873_, data_stage_2__5872_, data_stage_2__5871_, data_stage_2__5870_, data_stage_2__5869_, data_stage_2__5868_, data_stage_2__5867_, data_stage_2__5866_, data_stage_2__5865_, data_stage_2__5864_, data_stage_2__5863_, data_stage_2__5862_, data_stage_2__5861_, data_stage_2__5860_, data_stage_2__5859_, data_stage_2__5858_, data_stage_2__5857_, data_stage_2__5856_, data_stage_2__5855_, data_stage_2__5854_, data_stage_2__5853_, data_stage_2__5852_, data_stage_2__5851_, data_stage_2__5850_, data_stage_2__5849_, data_stage_2__5848_, data_stage_2__5847_, data_stage_2__5846_, data_stage_2__5845_, data_stage_2__5844_, data_stage_2__5843_, data_stage_2__5842_, data_stage_2__5841_, data_stage_2__5840_, data_stage_2__5839_, data_stage_2__5838_, data_stage_2__5837_, data_stage_2__5836_, data_stage_2__5835_, data_stage_2__5834_, data_stage_2__5833_, data_stage_2__5832_, data_stage_2__5831_, data_stage_2__5830_, data_stage_2__5829_, data_stage_2__5828_, data_stage_2__5827_, data_stage_2__5826_, data_stage_2__5825_, data_stage_2__5824_, data_stage_2__5823_, data_stage_2__5822_, data_stage_2__5821_, data_stage_2__5820_, data_stage_2__5819_, data_stage_2__5818_, data_stage_2__5817_, data_stage_2__5816_, data_stage_2__5815_, data_stage_2__5814_, data_stage_2__5813_, data_stage_2__5812_, data_stage_2__5811_, data_stage_2__5810_, data_stage_2__5809_, data_stage_2__5808_, data_stage_2__5807_, data_stage_2__5806_, data_stage_2__5805_, data_stage_2__5804_, data_stage_2__5803_, data_stage_2__5802_, data_stage_2__5801_, data_stage_2__5800_, data_stage_2__5799_, data_stage_2__5798_, data_stage_2__5797_, data_stage_2__5796_, data_stage_2__5795_, data_stage_2__5794_, data_stage_2__5793_, data_stage_2__5792_, data_stage_2__5791_, data_stage_2__5790_, data_stage_2__5789_, data_stage_2__5788_, data_stage_2__5787_, data_stage_2__5786_, data_stage_2__5785_, data_stage_2__5784_, data_stage_2__5783_, data_stage_2__5782_, data_stage_2__5781_, data_stage_2__5780_, data_stage_2__5779_, data_stage_2__5778_, data_stage_2__5777_, data_stage_2__5776_, data_stage_2__5775_, data_stage_2__5774_, data_stage_2__5773_, data_stage_2__5772_, data_stage_2__5771_, data_stage_2__5770_, data_stage_2__5769_, data_stage_2__5768_, data_stage_2__5767_, data_stage_2__5766_, data_stage_2__5765_, data_stage_2__5764_, data_stage_2__5763_, data_stage_2__5762_, data_stage_2__5761_, data_stage_2__5760_, data_stage_2__5759_, data_stage_2__5758_, data_stage_2__5757_, data_stage_2__5756_, data_stage_2__5755_, data_stage_2__5754_, data_stage_2__5753_, data_stage_2__5752_, data_stage_2__5751_, data_stage_2__5750_, data_stage_2__5749_, data_stage_2__5748_, data_stage_2__5747_, data_stage_2__5746_, data_stage_2__5745_, data_stage_2__5744_, data_stage_2__5743_, data_stage_2__5742_, data_stage_2__5741_, data_stage_2__5740_, data_stage_2__5739_, data_stage_2__5738_, data_stage_2__5737_, data_stage_2__5736_, data_stage_2__5735_, data_stage_2__5734_, data_stage_2__5733_, data_stage_2__5732_, data_stage_2__5731_, data_stage_2__5730_, data_stage_2__5729_, data_stage_2__5728_, data_stage_2__5727_, data_stage_2__5726_, data_stage_2__5725_, data_stage_2__5724_, data_stage_2__5723_, data_stage_2__5722_, data_stage_2__5721_, data_stage_2__5720_, data_stage_2__5719_, data_stage_2__5718_, data_stage_2__5717_, data_stage_2__5716_, data_stage_2__5715_, data_stage_2__5714_, data_stage_2__5713_, data_stage_2__5712_, data_stage_2__5711_, data_stage_2__5710_, data_stage_2__5709_, data_stage_2__5708_, data_stage_2__5707_, data_stage_2__5706_, data_stage_2__5705_, data_stage_2__5704_, data_stage_2__5703_, data_stage_2__5702_, data_stage_2__5701_, data_stage_2__5700_, data_stage_2__5699_, data_stage_2__5698_, data_stage_2__5697_, data_stage_2__5696_, data_stage_2__5695_, data_stage_2__5694_, data_stage_2__5693_, data_stage_2__5692_, data_stage_2__5691_, data_stage_2__5690_, data_stage_2__5689_, data_stage_2__5688_, data_stage_2__5687_, data_stage_2__5686_, data_stage_2__5685_, data_stage_2__5684_, data_stage_2__5683_, data_stage_2__5682_, data_stage_2__5681_, data_stage_2__5680_, data_stage_2__5679_, data_stage_2__5678_, data_stage_2__5677_, data_stage_2__5676_, data_stage_2__5675_, data_stage_2__5674_, data_stage_2__5673_, data_stage_2__5672_, data_stage_2__5671_, data_stage_2__5670_, data_stage_2__5669_, data_stage_2__5668_, data_stage_2__5667_, data_stage_2__5666_, data_stage_2__5665_, data_stage_2__5664_, data_stage_2__5663_, data_stage_2__5662_, data_stage_2__5661_, data_stage_2__5660_, data_stage_2__5659_, data_stage_2__5658_, data_stage_2__5657_, data_stage_2__5656_, data_stage_2__5655_, data_stage_2__5654_, data_stage_2__5653_, data_stage_2__5652_, data_stage_2__5651_, data_stage_2__5650_, data_stage_2__5649_, data_stage_2__5648_, data_stage_2__5647_, data_stage_2__5646_, data_stage_2__5645_, data_stage_2__5644_, data_stage_2__5643_, data_stage_2__5642_, data_stage_2__5641_, data_stage_2__5640_, data_stage_2__5639_, data_stage_2__5638_, data_stage_2__5637_, data_stage_2__5636_, data_stage_2__5635_, data_stage_2__5634_, data_stage_2__5633_, data_stage_2__5632_, data_stage_2__5631_, data_stage_2__5630_, data_stage_2__5629_, data_stage_2__5628_, data_stage_2__5627_, data_stage_2__5626_, data_stage_2__5625_, data_stage_2__5624_, data_stage_2__5623_, data_stage_2__5622_, data_stage_2__5621_, data_stage_2__5620_, data_stage_2__5619_, data_stage_2__5618_, data_stage_2__5617_, data_stage_2__5616_, data_stage_2__5615_, data_stage_2__5614_, data_stage_2__5613_, data_stage_2__5612_, data_stage_2__5611_, data_stage_2__5610_, data_stage_2__5609_, data_stage_2__5608_, data_stage_2__5607_, data_stage_2__5606_, data_stage_2__5605_, data_stage_2__5604_, data_stage_2__5603_, data_stage_2__5602_, data_stage_2__5601_, data_stage_2__5600_, data_stage_2__5599_, data_stage_2__5598_, data_stage_2__5597_, data_stage_2__5596_, data_stage_2__5595_, data_stage_2__5594_, data_stage_2__5593_, data_stage_2__5592_, data_stage_2__5591_, data_stage_2__5590_, data_stage_2__5589_, data_stage_2__5588_, data_stage_2__5587_, data_stage_2__5586_, data_stage_2__5585_, data_stage_2__5584_, data_stage_2__5583_, data_stage_2__5582_, data_stage_2__5581_, data_stage_2__5580_, data_stage_2__5579_, data_stage_2__5578_, data_stage_2__5577_, data_stage_2__5576_, data_stage_2__5575_, data_stage_2__5574_, data_stage_2__5573_, data_stage_2__5572_, data_stage_2__5571_, data_stage_2__5570_, data_stage_2__5569_, data_stage_2__5568_, data_stage_2__5567_, data_stage_2__5566_, data_stage_2__5565_, data_stage_2__5564_, data_stage_2__5563_, data_stage_2__5562_, data_stage_2__5561_, data_stage_2__5560_, data_stage_2__5559_, data_stage_2__5558_, data_stage_2__5557_, data_stage_2__5556_, data_stage_2__5555_, data_stage_2__5554_, data_stage_2__5553_, data_stage_2__5552_, data_stage_2__5551_, data_stage_2__5550_, data_stage_2__5549_, data_stage_2__5548_, data_stage_2__5547_, data_stage_2__5546_, data_stage_2__5545_, data_stage_2__5544_, data_stage_2__5543_, data_stage_2__5542_, data_stage_2__5541_, data_stage_2__5540_, data_stage_2__5539_, data_stage_2__5538_, data_stage_2__5537_, data_stage_2__5536_, data_stage_2__5535_, data_stage_2__5534_, data_stage_2__5533_, data_stage_2__5532_, data_stage_2__5531_, data_stage_2__5530_, data_stage_2__5529_, data_stage_2__5528_, data_stage_2__5527_, data_stage_2__5526_, data_stage_2__5525_, data_stage_2__5524_, data_stage_2__5523_, data_stage_2__5522_, data_stage_2__5521_, data_stage_2__5520_, data_stage_2__5519_, data_stage_2__5518_, data_stage_2__5517_, data_stage_2__5516_, data_stage_2__5515_, data_stage_2__5514_, data_stage_2__5513_, data_stage_2__5512_, data_stage_2__5511_, data_stage_2__5510_, data_stage_2__5509_, data_stage_2__5508_, data_stage_2__5507_, data_stage_2__5506_, data_stage_2__5505_, data_stage_2__5504_, data_stage_2__5503_, data_stage_2__5502_, data_stage_2__5501_, data_stage_2__5500_, data_stage_2__5499_, data_stage_2__5498_, data_stage_2__5497_, data_stage_2__5496_, data_stage_2__5495_, data_stage_2__5494_, data_stage_2__5493_, data_stage_2__5492_, data_stage_2__5491_, data_stage_2__5490_, data_stage_2__5489_, data_stage_2__5488_, data_stage_2__5487_, data_stage_2__5486_, data_stage_2__5485_, data_stage_2__5484_, data_stage_2__5483_, data_stage_2__5482_, data_stage_2__5481_, data_stage_2__5480_, data_stage_2__5479_, data_stage_2__5478_, data_stage_2__5477_, data_stage_2__5476_, data_stage_2__5475_, data_stage_2__5474_, data_stage_2__5473_, data_stage_2__5472_, data_stage_2__5471_, data_stage_2__5470_, data_stage_2__5469_, data_stage_2__5468_, data_stage_2__5467_, data_stage_2__5466_, data_stage_2__5465_, data_stage_2__5464_, data_stage_2__5463_, data_stage_2__5462_, data_stage_2__5461_, data_stage_2__5460_, data_stage_2__5459_, data_stage_2__5458_, data_stage_2__5457_, data_stage_2__5456_, data_stage_2__5455_, data_stage_2__5454_, data_stage_2__5453_, data_stage_2__5452_, data_stage_2__5451_, data_stage_2__5450_, data_stage_2__5449_, data_stage_2__5448_, data_stage_2__5447_, data_stage_2__5446_, data_stage_2__5445_, data_stage_2__5444_, data_stage_2__5443_, data_stage_2__5442_, data_stage_2__5441_, data_stage_2__5440_, data_stage_2__5439_, data_stage_2__5438_, data_stage_2__5437_, data_stage_2__5436_, data_stage_2__5435_, data_stage_2__5434_, data_stage_2__5433_, data_stage_2__5432_, data_stage_2__5431_, data_stage_2__5430_, data_stage_2__5429_, data_stage_2__5428_, data_stage_2__5427_, data_stage_2__5426_, data_stage_2__5425_, data_stage_2__5424_, data_stage_2__5423_, data_stage_2__5422_, data_stage_2__5421_, data_stage_2__5420_, data_stage_2__5419_, data_stage_2__5418_, data_stage_2__5417_, data_stage_2__5416_, data_stage_2__5415_, data_stage_2__5414_, data_stage_2__5413_, data_stage_2__5412_, data_stage_2__5411_, data_stage_2__5410_, data_stage_2__5409_, data_stage_2__5408_, data_stage_2__5407_, data_stage_2__5406_, data_stage_2__5405_, data_stage_2__5404_, data_stage_2__5403_, data_stage_2__5402_, data_stage_2__5401_, data_stage_2__5400_, data_stage_2__5399_, data_stage_2__5398_, data_stage_2__5397_, data_stage_2__5396_, data_stage_2__5395_, data_stage_2__5394_, data_stage_2__5393_, data_stage_2__5392_, data_stage_2__5391_, data_stage_2__5390_, data_stage_2__5389_, data_stage_2__5388_, data_stage_2__5387_, data_stage_2__5386_, data_stage_2__5385_, data_stage_2__5384_, data_stage_2__5383_, data_stage_2__5382_, data_stage_2__5381_, data_stage_2__5380_, data_stage_2__5379_, data_stage_2__5378_, data_stage_2__5377_, data_stage_2__5376_, data_stage_2__5375_, data_stage_2__5374_, data_stage_2__5373_, data_stage_2__5372_, data_stage_2__5371_, data_stage_2__5370_, data_stage_2__5369_, data_stage_2__5368_, data_stage_2__5367_, data_stage_2__5366_, data_stage_2__5365_, data_stage_2__5364_, data_stage_2__5363_, data_stage_2__5362_, data_stage_2__5361_, data_stage_2__5360_, data_stage_2__5359_, data_stage_2__5358_, data_stage_2__5357_, data_stage_2__5356_, data_stage_2__5355_, data_stage_2__5354_, data_stage_2__5353_, data_stage_2__5352_, data_stage_2__5351_, data_stage_2__5350_, data_stage_2__5349_, data_stage_2__5348_, data_stage_2__5347_, data_stage_2__5346_, data_stage_2__5345_, data_stage_2__5344_, data_stage_2__5343_, data_stage_2__5342_, data_stage_2__5341_, data_stage_2__5340_, data_stage_2__5339_, data_stage_2__5338_, data_stage_2__5337_, data_stage_2__5336_, data_stage_2__5335_, data_stage_2__5334_, data_stage_2__5333_, data_stage_2__5332_, data_stage_2__5331_, data_stage_2__5330_, data_stage_2__5329_, data_stage_2__5328_, data_stage_2__5327_, data_stage_2__5326_, data_stage_2__5325_, data_stage_2__5324_, data_stage_2__5323_, data_stage_2__5322_, data_stage_2__5321_, data_stage_2__5320_, data_stage_2__5319_, data_stage_2__5318_, data_stage_2__5317_, data_stage_2__5316_, data_stage_2__5315_, data_stage_2__5314_, data_stage_2__5313_, data_stage_2__5312_, data_stage_2__5311_, data_stage_2__5310_, data_stage_2__5309_, data_stage_2__5308_, data_stage_2__5307_, data_stage_2__5306_, data_stage_2__5305_, data_stage_2__5304_, data_stage_2__5303_, data_stage_2__5302_, data_stage_2__5301_, data_stage_2__5300_, data_stage_2__5299_, data_stage_2__5298_, data_stage_2__5297_, data_stage_2__5296_, data_stage_2__5295_, data_stage_2__5294_, data_stage_2__5293_, data_stage_2__5292_, data_stage_2__5291_, data_stage_2__5290_, data_stage_2__5289_, data_stage_2__5288_, data_stage_2__5287_, data_stage_2__5286_, data_stage_2__5285_, data_stage_2__5284_, data_stage_2__5283_, data_stage_2__5282_, data_stage_2__5281_, data_stage_2__5280_, data_stage_2__5279_, data_stage_2__5278_, data_stage_2__5277_, data_stage_2__5276_, data_stage_2__5275_, data_stage_2__5274_, data_stage_2__5273_, data_stage_2__5272_, data_stage_2__5271_, data_stage_2__5270_, data_stage_2__5269_, data_stage_2__5268_, data_stage_2__5267_, data_stage_2__5266_, data_stage_2__5265_, data_stage_2__5264_, data_stage_2__5263_, data_stage_2__5262_, data_stage_2__5261_, data_stage_2__5260_, data_stage_2__5259_, data_stage_2__5258_, data_stage_2__5257_, data_stage_2__5256_, data_stage_2__5255_, data_stage_2__5254_, data_stage_2__5253_, data_stage_2__5252_, data_stage_2__5251_, data_stage_2__5250_, data_stage_2__5249_, data_stage_2__5248_, data_stage_2__5247_, data_stage_2__5246_, data_stage_2__5245_, data_stage_2__5244_, data_stage_2__5243_, data_stage_2__5242_, data_stage_2__5241_, data_stage_2__5240_, data_stage_2__5239_, data_stage_2__5238_, data_stage_2__5237_, data_stage_2__5236_, data_stage_2__5235_, data_stage_2__5234_, data_stage_2__5233_, data_stage_2__5232_, data_stage_2__5231_, data_stage_2__5230_, data_stage_2__5229_, data_stage_2__5228_, data_stage_2__5227_, data_stage_2__5226_, data_stage_2__5225_, data_stage_2__5224_, data_stage_2__5223_, data_stage_2__5222_, data_stage_2__5221_, data_stage_2__5220_, data_stage_2__5219_, data_stage_2__5218_, data_stage_2__5217_, data_stage_2__5216_, data_stage_2__5215_, data_stage_2__5214_, data_stage_2__5213_, data_stage_2__5212_, data_stage_2__5211_, data_stage_2__5210_, data_stage_2__5209_, data_stage_2__5208_, data_stage_2__5207_, data_stage_2__5206_, data_stage_2__5205_, data_stage_2__5204_, data_stage_2__5203_, data_stage_2__5202_, data_stage_2__5201_, data_stage_2__5200_, data_stage_2__5199_, data_stage_2__5198_, data_stage_2__5197_, data_stage_2__5196_, data_stage_2__5195_, data_stage_2__5194_, data_stage_2__5193_, data_stage_2__5192_, data_stage_2__5191_, data_stage_2__5190_, data_stage_2__5189_, data_stage_2__5188_, data_stage_2__5187_, data_stage_2__5186_, data_stage_2__5185_, data_stage_2__5184_, data_stage_2__5183_, data_stage_2__5182_, data_stage_2__5181_, data_stage_2__5180_, data_stage_2__5179_, data_stage_2__5178_, data_stage_2__5177_, data_stage_2__5176_, data_stage_2__5175_, data_stage_2__5174_, data_stage_2__5173_, data_stage_2__5172_, data_stage_2__5171_, data_stage_2__5170_, data_stage_2__5169_, data_stage_2__5168_, data_stage_2__5167_, data_stage_2__5166_, data_stage_2__5165_, data_stage_2__5164_, data_stage_2__5163_, data_stage_2__5162_, data_stage_2__5161_, data_stage_2__5160_, data_stage_2__5159_, data_stage_2__5158_, data_stage_2__5157_, data_stage_2__5156_, data_stage_2__5155_, data_stage_2__5154_, data_stage_2__5153_, data_stage_2__5152_, data_stage_2__5151_, data_stage_2__5150_, data_stage_2__5149_, data_stage_2__5148_, data_stage_2__5147_, data_stage_2__5146_, data_stage_2__5145_, data_stage_2__5144_, data_stage_2__5143_, data_stage_2__5142_, data_stage_2__5141_, data_stage_2__5140_, data_stage_2__5139_, data_stage_2__5138_, data_stage_2__5137_, data_stage_2__5136_, data_stage_2__5135_, data_stage_2__5134_, data_stage_2__5133_, data_stage_2__5132_, data_stage_2__5131_, data_stage_2__5130_, data_stage_2__5129_, data_stage_2__5128_, data_stage_2__5127_, data_stage_2__5126_, data_stage_2__5125_, data_stage_2__5124_, data_stage_2__5123_, data_stage_2__5122_, data_stage_2__5121_, data_stage_2__5120_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__6143_, data_stage_3__6142_, data_stage_3__6141_, data_stage_3__6140_, data_stage_3__6139_, data_stage_3__6138_, data_stage_3__6137_, data_stage_3__6136_, data_stage_3__6135_, data_stage_3__6134_, data_stage_3__6133_, data_stage_3__6132_, data_stage_3__6131_, data_stage_3__6130_, data_stage_3__6129_, data_stage_3__6128_, data_stage_3__6127_, data_stage_3__6126_, data_stage_3__6125_, data_stage_3__6124_, data_stage_3__6123_, data_stage_3__6122_, data_stage_3__6121_, data_stage_3__6120_, data_stage_3__6119_, data_stage_3__6118_, data_stage_3__6117_, data_stage_3__6116_, data_stage_3__6115_, data_stage_3__6114_, data_stage_3__6113_, data_stage_3__6112_, data_stage_3__6111_, data_stage_3__6110_, data_stage_3__6109_, data_stage_3__6108_, data_stage_3__6107_, data_stage_3__6106_, data_stage_3__6105_, data_stage_3__6104_, data_stage_3__6103_, data_stage_3__6102_, data_stage_3__6101_, data_stage_3__6100_, data_stage_3__6099_, data_stage_3__6098_, data_stage_3__6097_, data_stage_3__6096_, data_stage_3__6095_, data_stage_3__6094_, data_stage_3__6093_, data_stage_3__6092_, data_stage_3__6091_, data_stage_3__6090_, data_stage_3__6089_, data_stage_3__6088_, data_stage_3__6087_, data_stage_3__6086_, data_stage_3__6085_, data_stage_3__6084_, data_stage_3__6083_, data_stage_3__6082_, data_stage_3__6081_, data_stage_3__6080_, data_stage_3__6079_, data_stage_3__6078_, data_stage_3__6077_, data_stage_3__6076_, data_stage_3__6075_, data_stage_3__6074_, data_stage_3__6073_, data_stage_3__6072_, data_stage_3__6071_, data_stage_3__6070_, data_stage_3__6069_, data_stage_3__6068_, data_stage_3__6067_, data_stage_3__6066_, data_stage_3__6065_, data_stage_3__6064_, data_stage_3__6063_, data_stage_3__6062_, data_stage_3__6061_, data_stage_3__6060_, data_stage_3__6059_, data_stage_3__6058_, data_stage_3__6057_, data_stage_3__6056_, data_stage_3__6055_, data_stage_3__6054_, data_stage_3__6053_, data_stage_3__6052_, data_stage_3__6051_, data_stage_3__6050_, data_stage_3__6049_, data_stage_3__6048_, data_stage_3__6047_, data_stage_3__6046_, data_stage_3__6045_, data_stage_3__6044_, data_stage_3__6043_, data_stage_3__6042_, data_stage_3__6041_, data_stage_3__6040_, data_stage_3__6039_, data_stage_3__6038_, data_stage_3__6037_, data_stage_3__6036_, data_stage_3__6035_, data_stage_3__6034_, data_stage_3__6033_, data_stage_3__6032_, data_stage_3__6031_, data_stage_3__6030_, data_stage_3__6029_, data_stage_3__6028_, data_stage_3__6027_, data_stage_3__6026_, data_stage_3__6025_, data_stage_3__6024_, data_stage_3__6023_, data_stage_3__6022_, data_stage_3__6021_, data_stage_3__6020_, data_stage_3__6019_, data_stage_3__6018_, data_stage_3__6017_, data_stage_3__6016_, data_stage_3__6015_, data_stage_3__6014_, data_stage_3__6013_, data_stage_3__6012_, data_stage_3__6011_, data_stage_3__6010_, data_stage_3__6009_, data_stage_3__6008_, data_stage_3__6007_, data_stage_3__6006_, data_stage_3__6005_, data_stage_3__6004_, data_stage_3__6003_, data_stage_3__6002_, data_stage_3__6001_, data_stage_3__6000_, data_stage_3__5999_, data_stage_3__5998_, data_stage_3__5997_, data_stage_3__5996_, data_stage_3__5995_, data_stage_3__5994_, data_stage_3__5993_, data_stage_3__5992_, data_stage_3__5991_, data_stage_3__5990_, data_stage_3__5989_, data_stage_3__5988_, data_stage_3__5987_, data_stage_3__5986_, data_stage_3__5985_, data_stage_3__5984_, data_stage_3__5983_, data_stage_3__5982_, data_stage_3__5981_, data_stage_3__5980_, data_stage_3__5979_, data_stage_3__5978_, data_stage_3__5977_, data_stage_3__5976_, data_stage_3__5975_, data_stage_3__5974_, data_stage_3__5973_, data_stage_3__5972_, data_stage_3__5971_, data_stage_3__5970_, data_stage_3__5969_, data_stage_3__5968_, data_stage_3__5967_, data_stage_3__5966_, data_stage_3__5965_, data_stage_3__5964_, data_stage_3__5963_, data_stage_3__5962_, data_stage_3__5961_, data_stage_3__5960_, data_stage_3__5959_, data_stage_3__5958_, data_stage_3__5957_, data_stage_3__5956_, data_stage_3__5955_, data_stage_3__5954_, data_stage_3__5953_, data_stage_3__5952_, data_stage_3__5951_, data_stage_3__5950_, data_stage_3__5949_, data_stage_3__5948_, data_stage_3__5947_, data_stage_3__5946_, data_stage_3__5945_, data_stage_3__5944_, data_stage_3__5943_, data_stage_3__5942_, data_stage_3__5941_, data_stage_3__5940_, data_stage_3__5939_, data_stage_3__5938_, data_stage_3__5937_, data_stage_3__5936_, data_stage_3__5935_, data_stage_3__5934_, data_stage_3__5933_, data_stage_3__5932_, data_stage_3__5931_, data_stage_3__5930_, data_stage_3__5929_, data_stage_3__5928_, data_stage_3__5927_, data_stage_3__5926_, data_stage_3__5925_, data_stage_3__5924_, data_stage_3__5923_, data_stage_3__5922_, data_stage_3__5921_, data_stage_3__5920_, data_stage_3__5919_, data_stage_3__5918_, data_stage_3__5917_, data_stage_3__5916_, data_stage_3__5915_, data_stage_3__5914_, data_stage_3__5913_, data_stage_3__5912_, data_stage_3__5911_, data_stage_3__5910_, data_stage_3__5909_, data_stage_3__5908_, data_stage_3__5907_, data_stage_3__5906_, data_stage_3__5905_, data_stage_3__5904_, data_stage_3__5903_, data_stage_3__5902_, data_stage_3__5901_, data_stage_3__5900_, data_stage_3__5899_, data_stage_3__5898_, data_stage_3__5897_, data_stage_3__5896_, data_stage_3__5895_, data_stage_3__5894_, data_stage_3__5893_, data_stage_3__5892_, data_stage_3__5891_, data_stage_3__5890_, data_stage_3__5889_, data_stage_3__5888_, data_stage_3__5887_, data_stage_3__5886_, data_stage_3__5885_, data_stage_3__5884_, data_stage_3__5883_, data_stage_3__5882_, data_stage_3__5881_, data_stage_3__5880_, data_stage_3__5879_, data_stage_3__5878_, data_stage_3__5877_, data_stage_3__5876_, data_stage_3__5875_, data_stage_3__5874_, data_stage_3__5873_, data_stage_3__5872_, data_stage_3__5871_, data_stage_3__5870_, data_stage_3__5869_, data_stage_3__5868_, data_stage_3__5867_, data_stage_3__5866_, data_stage_3__5865_, data_stage_3__5864_, data_stage_3__5863_, data_stage_3__5862_, data_stage_3__5861_, data_stage_3__5860_, data_stage_3__5859_, data_stage_3__5858_, data_stage_3__5857_, data_stage_3__5856_, data_stage_3__5855_, data_stage_3__5854_, data_stage_3__5853_, data_stage_3__5852_, data_stage_3__5851_, data_stage_3__5850_, data_stage_3__5849_, data_stage_3__5848_, data_stage_3__5847_, data_stage_3__5846_, data_stage_3__5845_, data_stage_3__5844_, data_stage_3__5843_, data_stage_3__5842_, data_stage_3__5841_, data_stage_3__5840_, data_stage_3__5839_, data_stage_3__5838_, data_stage_3__5837_, data_stage_3__5836_, data_stage_3__5835_, data_stage_3__5834_, data_stage_3__5833_, data_stage_3__5832_, data_stage_3__5831_, data_stage_3__5830_, data_stage_3__5829_, data_stage_3__5828_, data_stage_3__5827_, data_stage_3__5826_, data_stage_3__5825_, data_stage_3__5824_, data_stage_3__5823_, data_stage_3__5822_, data_stage_3__5821_, data_stage_3__5820_, data_stage_3__5819_, data_stage_3__5818_, data_stage_3__5817_, data_stage_3__5816_, data_stage_3__5815_, data_stage_3__5814_, data_stage_3__5813_, data_stage_3__5812_, data_stage_3__5811_, data_stage_3__5810_, data_stage_3__5809_, data_stage_3__5808_, data_stage_3__5807_, data_stage_3__5806_, data_stage_3__5805_, data_stage_3__5804_, data_stage_3__5803_, data_stage_3__5802_, data_stage_3__5801_, data_stage_3__5800_, data_stage_3__5799_, data_stage_3__5798_, data_stage_3__5797_, data_stage_3__5796_, data_stage_3__5795_, data_stage_3__5794_, data_stage_3__5793_, data_stage_3__5792_, data_stage_3__5791_, data_stage_3__5790_, data_stage_3__5789_, data_stage_3__5788_, data_stage_3__5787_, data_stage_3__5786_, data_stage_3__5785_, data_stage_3__5784_, data_stage_3__5783_, data_stage_3__5782_, data_stage_3__5781_, data_stage_3__5780_, data_stage_3__5779_, data_stage_3__5778_, data_stage_3__5777_, data_stage_3__5776_, data_stage_3__5775_, data_stage_3__5774_, data_stage_3__5773_, data_stage_3__5772_, data_stage_3__5771_, data_stage_3__5770_, data_stage_3__5769_, data_stage_3__5768_, data_stage_3__5767_, data_stage_3__5766_, data_stage_3__5765_, data_stage_3__5764_, data_stage_3__5763_, data_stage_3__5762_, data_stage_3__5761_, data_stage_3__5760_, data_stage_3__5759_, data_stage_3__5758_, data_stage_3__5757_, data_stage_3__5756_, data_stage_3__5755_, data_stage_3__5754_, data_stage_3__5753_, data_stage_3__5752_, data_stage_3__5751_, data_stage_3__5750_, data_stage_3__5749_, data_stage_3__5748_, data_stage_3__5747_, data_stage_3__5746_, data_stage_3__5745_, data_stage_3__5744_, data_stage_3__5743_, data_stage_3__5742_, data_stage_3__5741_, data_stage_3__5740_, data_stage_3__5739_, data_stage_3__5738_, data_stage_3__5737_, data_stage_3__5736_, data_stage_3__5735_, data_stage_3__5734_, data_stage_3__5733_, data_stage_3__5732_, data_stage_3__5731_, data_stage_3__5730_, data_stage_3__5729_, data_stage_3__5728_, data_stage_3__5727_, data_stage_3__5726_, data_stage_3__5725_, data_stage_3__5724_, data_stage_3__5723_, data_stage_3__5722_, data_stage_3__5721_, data_stage_3__5720_, data_stage_3__5719_, data_stage_3__5718_, data_stage_3__5717_, data_stage_3__5716_, data_stage_3__5715_, data_stage_3__5714_, data_stage_3__5713_, data_stage_3__5712_, data_stage_3__5711_, data_stage_3__5710_, data_stage_3__5709_, data_stage_3__5708_, data_stage_3__5707_, data_stage_3__5706_, data_stage_3__5705_, data_stage_3__5704_, data_stage_3__5703_, data_stage_3__5702_, data_stage_3__5701_, data_stage_3__5700_, data_stage_3__5699_, data_stage_3__5698_, data_stage_3__5697_, data_stage_3__5696_, data_stage_3__5695_, data_stage_3__5694_, data_stage_3__5693_, data_stage_3__5692_, data_stage_3__5691_, data_stage_3__5690_, data_stage_3__5689_, data_stage_3__5688_, data_stage_3__5687_, data_stage_3__5686_, data_stage_3__5685_, data_stage_3__5684_, data_stage_3__5683_, data_stage_3__5682_, data_stage_3__5681_, data_stage_3__5680_, data_stage_3__5679_, data_stage_3__5678_, data_stage_3__5677_, data_stage_3__5676_, data_stage_3__5675_, data_stage_3__5674_, data_stage_3__5673_, data_stage_3__5672_, data_stage_3__5671_, data_stage_3__5670_, data_stage_3__5669_, data_stage_3__5668_, data_stage_3__5667_, data_stage_3__5666_, data_stage_3__5665_, data_stage_3__5664_, data_stage_3__5663_, data_stage_3__5662_, data_stage_3__5661_, data_stage_3__5660_, data_stage_3__5659_, data_stage_3__5658_, data_stage_3__5657_, data_stage_3__5656_, data_stage_3__5655_, data_stage_3__5654_, data_stage_3__5653_, data_stage_3__5652_, data_stage_3__5651_, data_stage_3__5650_, data_stage_3__5649_, data_stage_3__5648_, data_stage_3__5647_, data_stage_3__5646_, data_stage_3__5645_, data_stage_3__5644_, data_stage_3__5643_, data_stage_3__5642_, data_stage_3__5641_, data_stage_3__5640_, data_stage_3__5639_, data_stage_3__5638_, data_stage_3__5637_, data_stage_3__5636_, data_stage_3__5635_, data_stage_3__5634_, data_stage_3__5633_, data_stage_3__5632_, data_stage_3__5631_, data_stage_3__5630_, data_stage_3__5629_, data_stage_3__5628_, data_stage_3__5627_, data_stage_3__5626_, data_stage_3__5625_, data_stage_3__5624_, data_stage_3__5623_, data_stage_3__5622_, data_stage_3__5621_, data_stage_3__5620_, data_stage_3__5619_, data_stage_3__5618_, data_stage_3__5617_, data_stage_3__5616_, data_stage_3__5615_, data_stage_3__5614_, data_stage_3__5613_, data_stage_3__5612_, data_stage_3__5611_, data_stage_3__5610_, data_stage_3__5609_, data_stage_3__5608_, data_stage_3__5607_, data_stage_3__5606_, data_stage_3__5605_, data_stage_3__5604_, data_stage_3__5603_, data_stage_3__5602_, data_stage_3__5601_, data_stage_3__5600_, data_stage_3__5599_, data_stage_3__5598_, data_stage_3__5597_, data_stage_3__5596_, data_stage_3__5595_, data_stage_3__5594_, data_stage_3__5593_, data_stage_3__5592_, data_stage_3__5591_, data_stage_3__5590_, data_stage_3__5589_, data_stage_3__5588_, data_stage_3__5587_, data_stage_3__5586_, data_stage_3__5585_, data_stage_3__5584_, data_stage_3__5583_, data_stage_3__5582_, data_stage_3__5581_, data_stage_3__5580_, data_stage_3__5579_, data_stage_3__5578_, data_stage_3__5577_, data_stage_3__5576_, data_stage_3__5575_, data_stage_3__5574_, data_stage_3__5573_, data_stage_3__5572_, data_stage_3__5571_, data_stage_3__5570_, data_stage_3__5569_, data_stage_3__5568_, data_stage_3__5567_, data_stage_3__5566_, data_stage_3__5565_, data_stage_3__5564_, data_stage_3__5563_, data_stage_3__5562_, data_stage_3__5561_, data_stage_3__5560_, data_stage_3__5559_, data_stage_3__5558_, data_stage_3__5557_, data_stage_3__5556_, data_stage_3__5555_, data_stage_3__5554_, data_stage_3__5553_, data_stage_3__5552_, data_stage_3__5551_, data_stage_3__5550_, data_stage_3__5549_, data_stage_3__5548_, data_stage_3__5547_, data_stage_3__5546_, data_stage_3__5545_, data_stage_3__5544_, data_stage_3__5543_, data_stage_3__5542_, data_stage_3__5541_, data_stage_3__5540_, data_stage_3__5539_, data_stage_3__5538_, data_stage_3__5537_, data_stage_3__5536_, data_stage_3__5535_, data_stage_3__5534_, data_stage_3__5533_, data_stage_3__5532_, data_stage_3__5531_, data_stage_3__5530_, data_stage_3__5529_, data_stage_3__5528_, data_stage_3__5527_, data_stage_3__5526_, data_stage_3__5525_, data_stage_3__5524_, data_stage_3__5523_, data_stage_3__5522_, data_stage_3__5521_, data_stage_3__5520_, data_stage_3__5519_, data_stage_3__5518_, data_stage_3__5517_, data_stage_3__5516_, data_stage_3__5515_, data_stage_3__5514_, data_stage_3__5513_, data_stage_3__5512_, data_stage_3__5511_, data_stage_3__5510_, data_stage_3__5509_, data_stage_3__5508_, data_stage_3__5507_, data_stage_3__5506_, data_stage_3__5505_, data_stage_3__5504_, data_stage_3__5503_, data_stage_3__5502_, data_stage_3__5501_, data_stage_3__5500_, data_stage_3__5499_, data_stage_3__5498_, data_stage_3__5497_, data_stage_3__5496_, data_stage_3__5495_, data_stage_3__5494_, data_stage_3__5493_, data_stage_3__5492_, data_stage_3__5491_, data_stage_3__5490_, data_stage_3__5489_, data_stage_3__5488_, data_stage_3__5487_, data_stage_3__5486_, data_stage_3__5485_, data_stage_3__5484_, data_stage_3__5483_, data_stage_3__5482_, data_stage_3__5481_, data_stage_3__5480_, data_stage_3__5479_, data_stage_3__5478_, data_stage_3__5477_, data_stage_3__5476_, data_stage_3__5475_, data_stage_3__5474_, data_stage_3__5473_, data_stage_3__5472_, data_stage_3__5471_, data_stage_3__5470_, data_stage_3__5469_, data_stage_3__5468_, data_stage_3__5467_, data_stage_3__5466_, data_stage_3__5465_, data_stage_3__5464_, data_stage_3__5463_, data_stage_3__5462_, data_stage_3__5461_, data_stage_3__5460_, data_stage_3__5459_, data_stage_3__5458_, data_stage_3__5457_, data_stage_3__5456_, data_stage_3__5455_, data_stage_3__5454_, data_stage_3__5453_, data_stage_3__5452_, data_stage_3__5451_, data_stage_3__5450_, data_stage_3__5449_, data_stage_3__5448_, data_stage_3__5447_, data_stage_3__5446_, data_stage_3__5445_, data_stage_3__5444_, data_stage_3__5443_, data_stage_3__5442_, data_stage_3__5441_, data_stage_3__5440_, data_stage_3__5439_, data_stage_3__5438_, data_stage_3__5437_, data_stage_3__5436_, data_stage_3__5435_, data_stage_3__5434_, data_stage_3__5433_, data_stage_3__5432_, data_stage_3__5431_, data_stage_3__5430_, data_stage_3__5429_, data_stage_3__5428_, data_stage_3__5427_, data_stage_3__5426_, data_stage_3__5425_, data_stage_3__5424_, data_stage_3__5423_, data_stage_3__5422_, data_stage_3__5421_, data_stage_3__5420_, data_stage_3__5419_, data_stage_3__5418_, data_stage_3__5417_, data_stage_3__5416_, data_stage_3__5415_, data_stage_3__5414_, data_stage_3__5413_, data_stage_3__5412_, data_stage_3__5411_, data_stage_3__5410_, data_stage_3__5409_, data_stage_3__5408_, data_stage_3__5407_, data_stage_3__5406_, data_stage_3__5405_, data_stage_3__5404_, data_stage_3__5403_, data_stage_3__5402_, data_stage_3__5401_, data_stage_3__5400_, data_stage_3__5399_, data_stage_3__5398_, data_stage_3__5397_, data_stage_3__5396_, data_stage_3__5395_, data_stage_3__5394_, data_stage_3__5393_, data_stage_3__5392_, data_stage_3__5391_, data_stage_3__5390_, data_stage_3__5389_, data_stage_3__5388_, data_stage_3__5387_, data_stage_3__5386_, data_stage_3__5385_, data_stage_3__5384_, data_stage_3__5383_, data_stage_3__5382_, data_stage_3__5381_, data_stage_3__5380_, data_stage_3__5379_, data_stage_3__5378_, data_stage_3__5377_, data_stage_3__5376_, data_stage_3__5375_, data_stage_3__5374_, data_stage_3__5373_, data_stage_3__5372_, data_stage_3__5371_, data_stage_3__5370_, data_stage_3__5369_, data_stage_3__5368_, data_stage_3__5367_, data_stage_3__5366_, data_stage_3__5365_, data_stage_3__5364_, data_stage_3__5363_, data_stage_3__5362_, data_stage_3__5361_, data_stage_3__5360_, data_stage_3__5359_, data_stage_3__5358_, data_stage_3__5357_, data_stage_3__5356_, data_stage_3__5355_, data_stage_3__5354_, data_stage_3__5353_, data_stage_3__5352_, data_stage_3__5351_, data_stage_3__5350_, data_stage_3__5349_, data_stage_3__5348_, data_stage_3__5347_, data_stage_3__5346_, data_stage_3__5345_, data_stage_3__5344_, data_stage_3__5343_, data_stage_3__5342_, data_stage_3__5341_, data_stage_3__5340_, data_stage_3__5339_, data_stage_3__5338_, data_stage_3__5337_, data_stage_3__5336_, data_stage_3__5335_, data_stage_3__5334_, data_stage_3__5333_, data_stage_3__5332_, data_stage_3__5331_, data_stage_3__5330_, data_stage_3__5329_, data_stage_3__5328_, data_stage_3__5327_, data_stage_3__5326_, data_stage_3__5325_, data_stage_3__5324_, data_stage_3__5323_, data_stage_3__5322_, data_stage_3__5321_, data_stage_3__5320_, data_stage_3__5319_, data_stage_3__5318_, data_stage_3__5317_, data_stage_3__5316_, data_stage_3__5315_, data_stage_3__5314_, data_stage_3__5313_, data_stage_3__5312_, data_stage_3__5311_, data_stage_3__5310_, data_stage_3__5309_, data_stage_3__5308_, data_stage_3__5307_, data_stage_3__5306_, data_stage_3__5305_, data_stage_3__5304_, data_stage_3__5303_, data_stage_3__5302_, data_stage_3__5301_, data_stage_3__5300_, data_stage_3__5299_, data_stage_3__5298_, data_stage_3__5297_, data_stage_3__5296_, data_stage_3__5295_, data_stage_3__5294_, data_stage_3__5293_, data_stage_3__5292_, data_stage_3__5291_, data_stage_3__5290_, data_stage_3__5289_, data_stage_3__5288_, data_stage_3__5287_, data_stage_3__5286_, data_stage_3__5285_, data_stage_3__5284_, data_stage_3__5283_, data_stage_3__5282_, data_stage_3__5281_, data_stage_3__5280_, data_stage_3__5279_, data_stage_3__5278_, data_stage_3__5277_, data_stage_3__5276_, data_stage_3__5275_, data_stage_3__5274_, data_stage_3__5273_, data_stage_3__5272_, data_stage_3__5271_, data_stage_3__5270_, data_stage_3__5269_, data_stage_3__5268_, data_stage_3__5267_, data_stage_3__5266_, data_stage_3__5265_, data_stage_3__5264_, data_stage_3__5263_, data_stage_3__5262_, data_stage_3__5261_, data_stage_3__5260_, data_stage_3__5259_, data_stage_3__5258_, data_stage_3__5257_, data_stage_3__5256_, data_stage_3__5255_, data_stage_3__5254_, data_stage_3__5253_, data_stage_3__5252_, data_stage_3__5251_, data_stage_3__5250_, data_stage_3__5249_, data_stage_3__5248_, data_stage_3__5247_, data_stage_3__5246_, data_stage_3__5245_, data_stage_3__5244_, data_stage_3__5243_, data_stage_3__5242_, data_stage_3__5241_, data_stage_3__5240_, data_stage_3__5239_, data_stage_3__5238_, data_stage_3__5237_, data_stage_3__5236_, data_stage_3__5235_, data_stage_3__5234_, data_stage_3__5233_, data_stage_3__5232_, data_stage_3__5231_, data_stage_3__5230_, data_stage_3__5229_, data_stage_3__5228_, data_stage_3__5227_, data_stage_3__5226_, data_stage_3__5225_, data_stage_3__5224_, data_stage_3__5223_, data_stage_3__5222_, data_stage_3__5221_, data_stage_3__5220_, data_stage_3__5219_, data_stage_3__5218_, data_stage_3__5217_, data_stage_3__5216_, data_stage_3__5215_, data_stage_3__5214_, data_stage_3__5213_, data_stage_3__5212_, data_stage_3__5211_, data_stage_3__5210_, data_stage_3__5209_, data_stage_3__5208_, data_stage_3__5207_, data_stage_3__5206_, data_stage_3__5205_, data_stage_3__5204_, data_stage_3__5203_, data_stage_3__5202_, data_stage_3__5201_, data_stage_3__5200_, data_stage_3__5199_, data_stage_3__5198_, data_stage_3__5197_, data_stage_3__5196_, data_stage_3__5195_, data_stage_3__5194_, data_stage_3__5193_, data_stage_3__5192_, data_stage_3__5191_, data_stage_3__5190_, data_stage_3__5189_, data_stage_3__5188_, data_stage_3__5187_, data_stage_3__5186_, data_stage_3__5185_, data_stage_3__5184_, data_stage_3__5183_, data_stage_3__5182_, data_stage_3__5181_, data_stage_3__5180_, data_stage_3__5179_, data_stage_3__5178_, data_stage_3__5177_, data_stage_3__5176_, data_stage_3__5175_, data_stage_3__5174_, data_stage_3__5173_, data_stage_3__5172_, data_stage_3__5171_, data_stage_3__5170_, data_stage_3__5169_, data_stage_3__5168_, data_stage_3__5167_, data_stage_3__5166_, data_stage_3__5165_, data_stage_3__5164_, data_stage_3__5163_, data_stage_3__5162_, data_stage_3__5161_, data_stage_3__5160_, data_stage_3__5159_, data_stage_3__5158_, data_stage_3__5157_, data_stage_3__5156_, data_stage_3__5155_, data_stage_3__5154_, data_stage_3__5153_, data_stage_3__5152_, data_stage_3__5151_, data_stage_3__5150_, data_stage_3__5149_, data_stage_3__5148_, data_stage_3__5147_, data_stage_3__5146_, data_stage_3__5145_, data_stage_3__5144_, data_stage_3__5143_, data_stage_3__5142_, data_stage_3__5141_, data_stage_3__5140_, data_stage_3__5139_, data_stage_3__5138_, data_stage_3__5137_, data_stage_3__5136_, data_stage_3__5135_, data_stage_3__5134_, data_stage_3__5133_, data_stage_3__5132_, data_stage_3__5131_, data_stage_3__5130_, data_stage_3__5129_, data_stage_3__5128_, data_stage_3__5127_, data_stage_3__5126_, data_stage_3__5125_, data_stage_3__5124_, data_stage_3__5123_, data_stage_3__5122_, data_stage_3__5121_, data_stage_3__5120_ })
  );


  bsg_swap_width_p512
  mux_stage_2__mux_swap_6__swap_inst
  (
    .data_i({ data_stage_2__7167_, data_stage_2__7166_, data_stage_2__7165_, data_stage_2__7164_, data_stage_2__7163_, data_stage_2__7162_, data_stage_2__7161_, data_stage_2__7160_, data_stage_2__7159_, data_stage_2__7158_, data_stage_2__7157_, data_stage_2__7156_, data_stage_2__7155_, data_stage_2__7154_, data_stage_2__7153_, data_stage_2__7152_, data_stage_2__7151_, data_stage_2__7150_, data_stage_2__7149_, data_stage_2__7148_, data_stage_2__7147_, data_stage_2__7146_, data_stage_2__7145_, data_stage_2__7144_, data_stage_2__7143_, data_stage_2__7142_, data_stage_2__7141_, data_stage_2__7140_, data_stage_2__7139_, data_stage_2__7138_, data_stage_2__7137_, data_stage_2__7136_, data_stage_2__7135_, data_stage_2__7134_, data_stage_2__7133_, data_stage_2__7132_, data_stage_2__7131_, data_stage_2__7130_, data_stage_2__7129_, data_stage_2__7128_, data_stage_2__7127_, data_stage_2__7126_, data_stage_2__7125_, data_stage_2__7124_, data_stage_2__7123_, data_stage_2__7122_, data_stage_2__7121_, data_stage_2__7120_, data_stage_2__7119_, data_stage_2__7118_, data_stage_2__7117_, data_stage_2__7116_, data_stage_2__7115_, data_stage_2__7114_, data_stage_2__7113_, data_stage_2__7112_, data_stage_2__7111_, data_stage_2__7110_, data_stage_2__7109_, data_stage_2__7108_, data_stage_2__7107_, data_stage_2__7106_, data_stage_2__7105_, data_stage_2__7104_, data_stage_2__7103_, data_stage_2__7102_, data_stage_2__7101_, data_stage_2__7100_, data_stage_2__7099_, data_stage_2__7098_, data_stage_2__7097_, data_stage_2__7096_, data_stage_2__7095_, data_stage_2__7094_, data_stage_2__7093_, data_stage_2__7092_, data_stage_2__7091_, data_stage_2__7090_, data_stage_2__7089_, data_stage_2__7088_, data_stage_2__7087_, data_stage_2__7086_, data_stage_2__7085_, data_stage_2__7084_, data_stage_2__7083_, data_stage_2__7082_, data_stage_2__7081_, data_stage_2__7080_, data_stage_2__7079_, data_stage_2__7078_, data_stage_2__7077_, data_stage_2__7076_, data_stage_2__7075_, data_stage_2__7074_, data_stage_2__7073_, data_stage_2__7072_, data_stage_2__7071_, data_stage_2__7070_, data_stage_2__7069_, data_stage_2__7068_, data_stage_2__7067_, data_stage_2__7066_, data_stage_2__7065_, data_stage_2__7064_, data_stage_2__7063_, data_stage_2__7062_, data_stage_2__7061_, data_stage_2__7060_, data_stage_2__7059_, data_stage_2__7058_, data_stage_2__7057_, data_stage_2__7056_, data_stage_2__7055_, data_stage_2__7054_, data_stage_2__7053_, data_stage_2__7052_, data_stage_2__7051_, data_stage_2__7050_, data_stage_2__7049_, data_stage_2__7048_, data_stage_2__7047_, data_stage_2__7046_, data_stage_2__7045_, data_stage_2__7044_, data_stage_2__7043_, data_stage_2__7042_, data_stage_2__7041_, data_stage_2__7040_, data_stage_2__7039_, data_stage_2__7038_, data_stage_2__7037_, data_stage_2__7036_, data_stage_2__7035_, data_stage_2__7034_, data_stage_2__7033_, data_stage_2__7032_, data_stage_2__7031_, data_stage_2__7030_, data_stage_2__7029_, data_stage_2__7028_, data_stage_2__7027_, data_stage_2__7026_, data_stage_2__7025_, data_stage_2__7024_, data_stage_2__7023_, data_stage_2__7022_, data_stage_2__7021_, data_stage_2__7020_, data_stage_2__7019_, data_stage_2__7018_, data_stage_2__7017_, data_stage_2__7016_, data_stage_2__7015_, data_stage_2__7014_, data_stage_2__7013_, data_stage_2__7012_, data_stage_2__7011_, data_stage_2__7010_, data_stage_2__7009_, data_stage_2__7008_, data_stage_2__7007_, data_stage_2__7006_, data_stage_2__7005_, data_stage_2__7004_, data_stage_2__7003_, data_stage_2__7002_, data_stage_2__7001_, data_stage_2__7000_, data_stage_2__6999_, data_stage_2__6998_, data_stage_2__6997_, data_stage_2__6996_, data_stage_2__6995_, data_stage_2__6994_, data_stage_2__6993_, data_stage_2__6992_, data_stage_2__6991_, data_stage_2__6990_, data_stage_2__6989_, data_stage_2__6988_, data_stage_2__6987_, data_stage_2__6986_, data_stage_2__6985_, data_stage_2__6984_, data_stage_2__6983_, data_stage_2__6982_, data_stage_2__6981_, data_stage_2__6980_, data_stage_2__6979_, data_stage_2__6978_, data_stage_2__6977_, data_stage_2__6976_, data_stage_2__6975_, data_stage_2__6974_, data_stage_2__6973_, data_stage_2__6972_, data_stage_2__6971_, data_stage_2__6970_, data_stage_2__6969_, data_stage_2__6968_, data_stage_2__6967_, data_stage_2__6966_, data_stage_2__6965_, data_stage_2__6964_, data_stage_2__6963_, data_stage_2__6962_, data_stage_2__6961_, data_stage_2__6960_, data_stage_2__6959_, data_stage_2__6958_, data_stage_2__6957_, data_stage_2__6956_, data_stage_2__6955_, data_stage_2__6954_, data_stage_2__6953_, data_stage_2__6952_, data_stage_2__6951_, data_stage_2__6950_, data_stage_2__6949_, data_stage_2__6948_, data_stage_2__6947_, data_stage_2__6946_, data_stage_2__6945_, data_stage_2__6944_, data_stage_2__6943_, data_stage_2__6942_, data_stage_2__6941_, data_stage_2__6940_, data_stage_2__6939_, data_stage_2__6938_, data_stage_2__6937_, data_stage_2__6936_, data_stage_2__6935_, data_stage_2__6934_, data_stage_2__6933_, data_stage_2__6932_, data_stage_2__6931_, data_stage_2__6930_, data_stage_2__6929_, data_stage_2__6928_, data_stage_2__6927_, data_stage_2__6926_, data_stage_2__6925_, data_stage_2__6924_, data_stage_2__6923_, data_stage_2__6922_, data_stage_2__6921_, data_stage_2__6920_, data_stage_2__6919_, data_stage_2__6918_, data_stage_2__6917_, data_stage_2__6916_, data_stage_2__6915_, data_stage_2__6914_, data_stage_2__6913_, data_stage_2__6912_, data_stage_2__6911_, data_stage_2__6910_, data_stage_2__6909_, data_stage_2__6908_, data_stage_2__6907_, data_stage_2__6906_, data_stage_2__6905_, data_stage_2__6904_, data_stage_2__6903_, data_stage_2__6902_, data_stage_2__6901_, data_stage_2__6900_, data_stage_2__6899_, data_stage_2__6898_, data_stage_2__6897_, data_stage_2__6896_, data_stage_2__6895_, data_stage_2__6894_, data_stage_2__6893_, data_stage_2__6892_, data_stage_2__6891_, data_stage_2__6890_, data_stage_2__6889_, data_stage_2__6888_, data_stage_2__6887_, data_stage_2__6886_, data_stage_2__6885_, data_stage_2__6884_, data_stage_2__6883_, data_stage_2__6882_, data_stage_2__6881_, data_stage_2__6880_, data_stage_2__6879_, data_stage_2__6878_, data_stage_2__6877_, data_stage_2__6876_, data_stage_2__6875_, data_stage_2__6874_, data_stage_2__6873_, data_stage_2__6872_, data_stage_2__6871_, data_stage_2__6870_, data_stage_2__6869_, data_stage_2__6868_, data_stage_2__6867_, data_stage_2__6866_, data_stage_2__6865_, data_stage_2__6864_, data_stage_2__6863_, data_stage_2__6862_, data_stage_2__6861_, data_stage_2__6860_, data_stage_2__6859_, data_stage_2__6858_, data_stage_2__6857_, data_stage_2__6856_, data_stage_2__6855_, data_stage_2__6854_, data_stage_2__6853_, data_stage_2__6852_, data_stage_2__6851_, data_stage_2__6850_, data_stage_2__6849_, data_stage_2__6848_, data_stage_2__6847_, data_stage_2__6846_, data_stage_2__6845_, data_stage_2__6844_, data_stage_2__6843_, data_stage_2__6842_, data_stage_2__6841_, data_stage_2__6840_, data_stage_2__6839_, data_stage_2__6838_, data_stage_2__6837_, data_stage_2__6836_, data_stage_2__6835_, data_stage_2__6834_, data_stage_2__6833_, data_stage_2__6832_, data_stage_2__6831_, data_stage_2__6830_, data_stage_2__6829_, data_stage_2__6828_, data_stage_2__6827_, data_stage_2__6826_, data_stage_2__6825_, data_stage_2__6824_, data_stage_2__6823_, data_stage_2__6822_, data_stage_2__6821_, data_stage_2__6820_, data_stage_2__6819_, data_stage_2__6818_, data_stage_2__6817_, data_stage_2__6816_, data_stage_2__6815_, data_stage_2__6814_, data_stage_2__6813_, data_stage_2__6812_, data_stage_2__6811_, data_stage_2__6810_, data_stage_2__6809_, data_stage_2__6808_, data_stage_2__6807_, data_stage_2__6806_, data_stage_2__6805_, data_stage_2__6804_, data_stage_2__6803_, data_stage_2__6802_, data_stage_2__6801_, data_stage_2__6800_, data_stage_2__6799_, data_stage_2__6798_, data_stage_2__6797_, data_stage_2__6796_, data_stage_2__6795_, data_stage_2__6794_, data_stage_2__6793_, data_stage_2__6792_, data_stage_2__6791_, data_stage_2__6790_, data_stage_2__6789_, data_stage_2__6788_, data_stage_2__6787_, data_stage_2__6786_, data_stage_2__6785_, data_stage_2__6784_, data_stage_2__6783_, data_stage_2__6782_, data_stage_2__6781_, data_stage_2__6780_, data_stage_2__6779_, data_stage_2__6778_, data_stage_2__6777_, data_stage_2__6776_, data_stage_2__6775_, data_stage_2__6774_, data_stage_2__6773_, data_stage_2__6772_, data_stage_2__6771_, data_stage_2__6770_, data_stage_2__6769_, data_stage_2__6768_, data_stage_2__6767_, data_stage_2__6766_, data_stage_2__6765_, data_stage_2__6764_, data_stage_2__6763_, data_stage_2__6762_, data_stage_2__6761_, data_stage_2__6760_, data_stage_2__6759_, data_stage_2__6758_, data_stage_2__6757_, data_stage_2__6756_, data_stage_2__6755_, data_stage_2__6754_, data_stage_2__6753_, data_stage_2__6752_, data_stage_2__6751_, data_stage_2__6750_, data_stage_2__6749_, data_stage_2__6748_, data_stage_2__6747_, data_stage_2__6746_, data_stage_2__6745_, data_stage_2__6744_, data_stage_2__6743_, data_stage_2__6742_, data_stage_2__6741_, data_stage_2__6740_, data_stage_2__6739_, data_stage_2__6738_, data_stage_2__6737_, data_stage_2__6736_, data_stage_2__6735_, data_stage_2__6734_, data_stage_2__6733_, data_stage_2__6732_, data_stage_2__6731_, data_stage_2__6730_, data_stage_2__6729_, data_stage_2__6728_, data_stage_2__6727_, data_stage_2__6726_, data_stage_2__6725_, data_stage_2__6724_, data_stage_2__6723_, data_stage_2__6722_, data_stage_2__6721_, data_stage_2__6720_, data_stage_2__6719_, data_stage_2__6718_, data_stage_2__6717_, data_stage_2__6716_, data_stage_2__6715_, data_stage_2__6714_, data_stage_2__6713_, data_stage_2__6712_, data_stage_2__6711_, data_stage_2__6710_, data_stage_2__6709_, data_stage_2__6708_, data_stage_2__6707_, data_stage_2__6706_, data_stage_2__6705_, data_stage_2__6704_, data_stage_2__6703_, data_stage_2__6702_, data_stage_2__6701_, data_stage_2__6700_, data_stage_2__6699_, data_stage_2__6698_, data_stage_2__6697_, data_stage_2__6696_, data_stage_2__6695_, data_stage_2__6694_, data_stage_2__6693_, data_stage_2__6692_, data_stage_2__6691_, data_stage_2__6690_, data_stage_2__6689_, data_stage_2__6688_, data_stage_2__6687_, data_stage_2__6686_, data_stage_2__6685_, data_stage_2__6684_, data_stage_2__6683_, data_stage_2__6682_, data_stage_2__6681_, data_stage_2__6680_, data_stage_2__6679_, data_stage_2__6678_, data_stage_2__6677_, data_stage_2__6676_, data_stage_2__6675_, data_stage_2__6674_, data_stage_2__6673_, data_stage_2__6672_, data_stage_2__6671_, data_stage_2__6670_, data_stage_2__6669_, data_stage_2__6668_, data_stage_2__6667_, data_stage_2__6666_, data_stage_2__6665_, data_stage_2__6664_, data_stage_2__6663_, data_stage_2__6662_, data_stage_2__6661_, data_stage_2__6660_, data_stage_2__6659_, data_stage_2__6658_, data_stage_2__6657_, data_stage_2__6656_, data_stage_2__6655_, data_stage_2__6654_, data_stage_2__6653_, data_stage_2__6652_, data_stage_2__6651_, data_stage_2__6650_, data_stage_2__6649_, data_stage_2__6648_, data_stage_2__6647_, data_stage_2__6646_, data_stage_2__6645_, data_stage_2__6644_, data_stage_2__6643_, data_stage_2__6642_, data_stage_2__6641_, data_stage_2__6640_, data_stage_2__6639_, data_stage_2__6638_, data_stage_2__6637_, data_stage_2__6636_, data_stage_2__6635_, data_stage_2__6634_, data_stage_2__6633_, data_stage_2__6632_, data_stage_2__6631_, data_stage_2__6630_, data_stage_2__6629_, data_stage_2__6628_, data_stage_2__6627_, data_stage_2__6626_, data_stage_2__6625_, data_stage_2__6624_, data_stage_2__6623_, data_stage_2__6622_, data_stage_2__6621_, data_stage_2__6620_, data_stage_2__6619_, data_stage_2__6618_, data_stage_2__6617_, data_stage_2__6616_, data_stage_2__6615_, data_stage_2__6614_, data_stage_2__6613_, data_stage_2__6612_, data_stage_2__6611_, data_stage_2__6610_, data_stage_2__6609_, data_stage_2__6608_, data_stage_2__6607_, data_stage_2__6606_, data_stage_2__6605_, data_stage_2__6604_, data_stage_2__6603_, data_stage_2__6602_, data_stage_2__6601_, data_stage_2__6600_, data_stage_2__6599_, data_stage_2__6598_, data_stage_2__6597_, data_stage_2__6596_, data_stage_2__6595_, data_stage_2__6594_, data_stage_2__6593_, data_stage_2__6592_, data_stage_2__6591_, data_stage_2__6590_, data_stage_2__6589_, data_stage_2__6588_, data_stage_2__6587_, data_stage_2__6586_, data_stage_2__6585_, data_stage_2__6584_, data_stage_2__6583_, data_stage_2__6582_, data_stage_2__6581_, data_stage_2__6580_, data_stage_2__6579_, data_stage_2__6578_, data_stage_2__6577_, data_stage_2__6576_, data_stage_2__6575_, data_stage_2__6574_, data_stage_2__6573_, data_stage_2__6572_, data_stage_2__6571_, data_stage_2__6570_, data_stage_2__6569_, data_stage_2__6568_, data_stage_2__6567_, data_stage_2__6566_, data_stage_2__6565_, data_stage_2__6564_, data_stage_2__6563_, data_stage_2__6562_, data_stage_2__6561_, data_stage_2__6560_, data_stage_2__6559_, data_stage_2__6558_, data_stage_2__6557_, data_stage_2__6556_, data_stage_2__6555_, data_stage_2__6554_, data_stage_2__6553_, data_stage_2__6552_, data_stage_2__6551_, data_stage_2__6550_, data_stage_2__6549_, data_stage_2__6548_, data_stage_2__6547_, data_stage_2__6546_, data_stage_2__6545_, data_stage_2__6544_, data_stage_2__6543_, data_stage_2__6542_, data_stage_2__6541_, data_stage_2__6540_, data_stage_2__6539_, data_stage_2__6538_, data_stage_2__6537_, data_stage_2__6536_, data_stage_2__6535_, data_stage_2__6534_, data_stage_2__6533_, data_stage_2__6532_, data_stage_2__6531_, data_stage_2__6530_, data_stage_2__6529_, data_stage_2__6528_, data_stage_2__6527_, data_stage_2__6526_, data_stage_2__6525_, data_stage_2__6524_, data_stage_2__6523_, data_stage_2__6522_, data_stage_2__6521_, data_stage_2__6520_, data_stage_2__6519_, data_stage_2__6518_, data_stage_2__6517_, data_stage_2__6516_, data_stage_2__6515_, data_stage_2__6514_, data_stage_2__6513_, data_stage_2__6512_, data_stage_2__6511_, data_stage_2__6510_, data_stage_2__6509_, data_stage_2__6508_, data_stage_2__6507_, data_stage_2__6506_, data_stage_2__6505_, data_stage_2__6504_, data_stage_2__6503_, data_stage_2__6502_, data_stage_2__6501_, data_stage_2__6500_, data_stage_2__6499_, data_stage_2__6498_, data_stage_2__6497_, data_stage_2__6496_, data_stage_2__6495_, data_stage_2__6494_, data_stage_2__6493_, data_stage_2__6492_, data_stage_2__6491_, data_stage_2__6490_, data_stage_2__6489_, data_stage_2__6488_, data_stage_2__6487_, data_stage_2__6486_, data_stage_2__6485_, data_stage_2__6484_, data_stage_2__6483_, data_stage_2__6482_, data_stage_2__6481_, data_stage_2__6480_, data_stage_2__6479_, data_stage_2__6478_, data_stage_2__6477_, data_stage_2__6476_, data_stage_2__6475_, data_stage_2__6474_, data_stage_2__6473_, data_stage_2__6472_, data_stage_2__6471_, data_stage_2__6470_, data_stage_2__6469_, data_stage_2__6468_, data_stage_2__6467_, data_stage_2__6466_, data_stage_2__6465_, data_stage_2__6464_, data_stage_2__6463_, data_stage_2__6462_, data_stage_2__6461_, data_stage_2__6460_, data_stage_2__6459_, data_stage_2__6458_, data_stage_2__6457_, data_stage_2__6456_, data_stage_2__6455_, data_stage_2__6454_, data_stage_2__6453_, data_stage_2__6452_, data_stage_2__6451_, data_stage_2__6450_, data_stage_2__6449_, data_stage_2__6448_, data_stage_2__6447_, data_stage_2__6446_, data_stage_2__6445_, data_stage_2__6444_, data_stage_2__6443_, data_stage_2__6442_, data_stage_2__6441_, data_stage_2__6440_, data_stage_2__6439_, data_stage_2__6438_, data_stage_2__6437_, data_stage_2__6436_, data_stage_2__6435_, data_stage_2__6434_, data_stage_2__6433_, data_stage_2__6432_, data_stage_2__6431_, data_stage_2__6430_, data_stage_2__6429_, data_stage_2__6428_, data_stage_2__6427_, data_stage_2__6426_, data_stage_2__6425_, data_stage_2__6424_, data_stage_2__6423_, data_stage_2__6422_, data_stage_2__6421_, data_stage_2__6420_, data_stage_2__6419_, data_stage_2__6418_, data_stage_2__6417_, data_stage_2__6416_, data_stage_2__6415_, data_stage_2__6414_, data_stage_2__6413_, data_stage_2__6412_, data_stage_2__6411_, data_stage_2__6410_, data_stage_2__6409_, data_stage_2__6408_, data_stage_2__6407_, data_stage_2__6406_, data_stage_2__6405_, data_stage_2__6404_, data_stage_2__6403_, data_stage_2__6402_, data_stage_2__6401_, data_stage_2__6400_, data_stage_2__6399_, data_stage_2__6398_, data_stage_2__6397_, data_stage_2__6396_, data_stage_2__6395_, data_stage_2__6394_, data_stage_2__6393_, data_stage_2__6392_, data_stage_2__6391_, data_stage_2__6390_, data_stage_2__6389_, data_stage_2__6388_, data_stage_2__6387_, data_stage_2__6386_, data_stage_2__6385_, data_stage_2__6384_, data_stage_2__6383_, data_stage_2__6382_, data_stage_2__6381_, data_stage_2__6380_, data_stage_2__6379_, data_stage_2__6378_, data_stage_2__6377_, data_stage_2__6376_, data_stage_2__6375_, data_stage_2__6374_, data_stage_2__6373_, data_stage_2__6372_, data_stage_2__6371_, data_stage_2__6370_, data_stage_2__6369_, data_stage_2__6368_, data_stage_2__6367_, data_stage_2__6366_, data_stage_2__6365_, data_stage_2__6364_, data_stage_2__6363_, data_stage_2__6362_, data_stage_2__6361_, data_stage_2__6360_, data_stage_2__6359_, data_stage_2__6358_, data_stage_2__6357_, data_stage_2__6356_, data_stage_2__6355_, data_stage_2__6354_, data_stage_2__6353_, data_stage_2__6352_, data_stage_2__6351_, data_stage_2__6350_, data_stage_2__6349_, data_stage_2__6348_, data_stage_2__6347_, data_stage_2__6346_, data_stage_2__6345_, data_stage_2__6344_, data_stage_2__6343_, data_stage_2__6342_, data_stage_2__6341_, data_stage_2__6340_, data_stage_2__6339_, data_stage_2__6338_, data_stage_2__6337_, data_stage_2__6336_, data_stage_2__6335_, data_stage_2__6334_, data_stage_2__6333_, data_stage_2__6332_, data_stage_2__6331_, data_stage_2__6330_, data_stage_2__6329_, data_stage_2__6328_, data_stage_2__6327_, data_stage_2__6326_, data_stage_2__6325_, data_stage_2__6324_, data_stage_2__6323_, data_stage_2__6322_, data_stage_2__6321_, data_stage_2__6320_, data_stage_2__6319_, data_stage_2__6318_, data_stage_2__6317_, data_stage_2__6316_, data_stage_2__6315_, data_stage_2__6314_, data_stage_2__6313_, data_stage_2__6312_, data_stage_2__6311_, data_stage_2__6310_, data_stage_2__6309_, data_stage_2__6308_, data_stage_2__6307_, data_stage_2__6306_, data_stage_2__6305_, data_stage_2__6304_, data_stage_2__6303_, data_stage_2__6302_, data_stage_2__6301_, data_stage_2__6300_, data_stage_2__6299_, data_stage_2__6298_, data_stage_2__6297_, data_stage_2__6296_, data_stage_2__6295_, data_stage_2__6294_, data_stage_2__6293_, data_stage_2__6292_, data_stage_2__6291_, data_stage_2__6290_, data_stage_2__6289_, data_stage_2__6288_, data_stage_2__6287_, data_stage_2__6286_, data_stage_2__6285_, data_stage_2__6284_, data_stage_2__6283_, data_stage_2__6282_, data_stage_2__6281_, data_stage_2__6280_, data_stage_2__6279_, data_stage_2__6278_, data_stage_2__6277_, data_stage_2__6276_, data_stage_2__6275_, data_stage_2__6274_, data_stage_2__6273_, data_stage_2__6272_, data_stage_2__6271_, data_stage_2__6270_, data_stage_2__6269_, data_stage_2__6268_, data_stage_2__6267_, data_stage_2__6266_, data_stage_2__6265_, data_stage_2__6264_, data_stage_2__6263_, data_stage_2__6262_, data_stage_2__6261_, data_stage_2__6260_, data_stage_2__6259_, data_stage_2__6258_, data_stage_2__6257_, data_stage_2__6256_, data_stage_2__6255_, data_stage_2__6254_, data_stage_2__6253_, data_stage_2__6252_, data_stage_2__6251_, data_stage_2__6250_, data_stage_2__6249_, data_stage_2__6248_, data_stage_2__6247_, data_stage_2__6246_, data_stage_2__6245_, data_stage_2__6244_, data_stage_2__6243_, data_stage_2__6242_, data_stage_2__6241_, data_stage_2__6240_, data_stage_2__6239_, data_stage_2__6238_, data_stage_2__6237_, data_stage_2__6236_, data_stage_2__6235_, data_stage_2__6234_, data_stage_2__6233_, data_stage_2__6232_, data_stage_2__6231_, data_stage_2__6230_, data_stage_2__6229_, data_stage_2__6228_, data_stage_2__6227_, data_stage_2__6226_, data_stage_2__6225_, data_stage_2__6224_, data_stage_2__6223_, data_stage_2__6222_, data_stage_2__6221_, data_stage_2__6220_, data_stage_2__6219_, data_stage_2__6218_, data_stage_2__6217_, data_stage_2__6216_, data_stage_2__6215_, data_stage_2__6214_, data_stage_2__6213_, data_stage_2__6212_, data_stage_2__6211_, data_stage_2__6210_, data_stage_2__6209_, data_stage_2__6208_, data_stage_2__6207_, data_stage_2__6206_, data_stage_2__6205_, data_stage_2__6204_, data_stage_2__6203_, data_stage_2__6202_, data_stage_2__6201_, data_stage_2__6200_, data_stage_2__6199_, data_stage_2__6198_, data_stage_2__6197_, data_stage_2__6196_, data_stage_2__6195_, data_stage_2__6194_, data_stage_2__6193_, data_stage_2__6192_, data_stage_2__6191_, data_stage_2__6190_, data_stage_2__6189_, data_stage_2__6188_, data_stage_2__6187_, data_stage_2__6186_, data_stage_2__6185_, data_stage_2__6184_, data_stage_2__6183_, data_stage_2__6182_, data_stage_2__6181_, data_stage_2__6180_, data_stage_2__6179_, data_stage_2__6178_, data_stage_2__6177_, data_stage_2__6176_, data_stage_2__6175_, data_stage_2__6174_, data_stage_2__6173_, data_stage_2__6172_, data_stage_2__6171_, data_stage_2__6170_, data_stage_2__6169_, data_stage_2__6168_, data_stage_2__6167_, data_stage_2__6166_, data_stage_2__6165_, data_stage_2__6164_, data_stage_2__6163_, data_stage_2__6162_, data_stage_2__6161_, data_stage_2__6160_, data_stage_2__6159_, data_stage_2__6158_, data_stage_2__6157_, data_stage_2__6156_, data_stage_2__6155_, data_stage_2__6154_, data_stage_2__6153_, data_stage_2__6152_, data_stage_2__6151_, data_stage_2__6150_, data_stage_2__6149_, data_stage_2__6148_, data_stage_2__6147_, data_stage_2__6146_, data_stage_2__6145_, data_stage_2__6144_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__7167_, data_stage_3__7166_, data_stage_3__7165_, data_stage_3__7164_, data_stage_3__7163_, data_stage_3__7162_, data_stage_3__7161_, data_stage_3__7160_, data_stage_3__7159_, data_stage_3__7158_, data_stage_3__7157_, data_stage_3__7156_, data_stage_3__7155_, data_stage_3__7154_, data_stage_3__7153_, data_stage_3__7152_, data_stage_3__7151_, data_stage_3__7150_, data_stage_3__7149_, data_stage_3__7148_, data_stage_3__7147_, data_stage_3__7146_, data_stage_3__7145_, data_stage_3__7144_, data_stage_3__7143_, data_stage_3__7142_, data_stage_3__7141_, data_stage_3__7140_, data_stage_3__7139_, data_stage_3__7138_, data_stage_3__7137_, data_stage_3__7136_, data_stage_3__7135_, data_stage_3__7134_, data_stage_3__7133_, data_stage_3__7132_, data_stage_3__7131_, data_stage_3__7130_, data_stage_3__7129_, data_stage_3__7128_, data_stage_3__7127_, data_stage_3__7126_, data_stage_3__7125_, data_stage_3__7124_, data_stage_3__7123_, data_stage_3__7122_, data_stage_3__7121_, data_stage_3__7120_, data_stage_3__7119_, data_stage_3__7118_, data_stage_3__7117_, data_stage_3__7116_, data_stage_3__7115_, data_stage_3__7114_, data_stage_3__7113_, data_stage_3__7112_, data_stage_3__7111_, data_stage_3__7110_, data_stage_3__7109_, data_stage_3__7108_, data_stage_3__7107_, data_stage_3__7106_, data_stage_3__7105_, data_stage_3__7104_, data_stage_3__7103_, data_stage_3__7102_, data_stage_3__7101_, data_stage_3__7100_, data_stage_3__7099_, data_stage_3__7098_, data_stage_3__7097_, data_stage_3__7096_, data_stage_3__7095_, data_stage_3__7094_, data_stage_3__7093_, data_stage_3__7092_, data_stage_3__7091_, data_stage_3__7090_, data_stage_3__7089_, data_stage_3__7088_, data_stage_3__7087_, data_stage_3__7086_, data_stage_3__7085_, data_stage_3__7084_, data_stage_3__7083_, data_stage_3__7082_, data_stage_3__7081_, data_stage_3__7080_, data_stage_3__7079_, data_stage_3__7078_, data_stage_3__7077_, data_stage_3__7076_, data_stage_3__7075_, data_stage_3__7074_, data_stage_3__7073_, data_stage_3__7072_, data_stage_3__7071_, data_stage_3__7070_, data_stage_3__7069_, data_stage_3__7068_, data_stage_3__7067_, data_stage_3__7066_, data_stage_3__7065_, data_stage_3__7064_, data_stage_3__7063_, data_stage_3__7062_, data_stage_3__7061_, data_stage_3__7060_, data_stage_3__7059_, data_stage_3__7058_, data_stage_3__7057_, data_stage_3__7056_, data_stage_3__7055_, data_stage_3__7054_, data_stage_3__7053_, data_stage_3__7052_, data_stage_3__7051_, data_stage_3__7050_, data_stage_3__7049_, data_stage_3__7048_, data_stage_3__7047_, data_stage_3__7046_, data_stage_3__7045_, data_stage_3__7044_, data_stage_3__7043_, data_stage_3__7042_, data_stage_3__7041_, data_stage_3__7040_, data_stage_3__7039_, data_stage_3__7038_, data_stage_3__7037_, data_stage_3__7036_, data_stage_3__7035_, data_stage_3__7034_, data_stage_3__7033_, data_stage_3__7032_, data_stage_3__7031_, data_stage_3__7030_, data_stage_3__7029_, data_stage_3__7028_, data_stage_3__7027_, data_stage_3__7026_, data_stage_3__7025_, data_stage_3__7024_, data_stage_3__7023_, data_stage_3__7022_, data_stage_3__7021_, data_stage_3__7020_, data_stage_3__7019_, data_stage_3__7018_, data_stage_3__7017_, data_stage_3__7016_, data_stage_3__7015_, data_stage_3__7014_, data_stage_3__7013_, data_stage_3__7012_, data_stage_3__7011_, data_stage_3__7010_, data_stage_3__7009_, data_stage_3__7008_, data_stage_3__7007_, data_stage_3__7006_, data_stage_3__7005_, data_stage_3__7004_, data_stage_3__7003_, data_stage_3__7002_, data_stage_3__7001_, data_stage_3__7000_, data_stage_3__6999_, data_stage_3__6998_, data_stage_3__6997_, data_stage_3__6996_, data_stage_3__6995_, data_stage_3__6994_, data_stage_3__6993_, data_stage_3__6992_, data_stage_3__6991_, data_stage_3__6990_, data_stage_3__6989_, data_stage_3__6988_, data_stage_3__6987_, data_stage_3__6986_, data_stage_3__6985_, data_stage_3__6984_, data_stage_3__6983_, data_stage_3__6982_, data_stage_3__6981_, data_stage_3__6980_, data_stage_3__6979_, data_stage_3__6978_, data_stage_3__6977_, data_stage_3__6976_, data_stage_3__6975_, data_stage_3__6974_, data_stage_3__6973_, data_stage_3__6972_, data_stage_3__6971_, data_stage_3__6970_, data_stage_3__6969_, data_stage_3__6968_, data_stage_3__6967_, data_stage_3__6966_, data_stage_3__6965_, data_stage_3__6964_, data_stage_3__6963_, data_stage_3__6962_, data_stage_3__6961_, data_stage_3__6960_, data_stage_3__6959_, data_stage_3__6958_, data_stage_3__6957_, data_stage_3__6956_, data_stage_3__6955_, data_stage_3__6954_, data_stage_3__6953_, data_stage_3__6952_, data_stage_3__6951_, data_stage_3__6950_, data_stage_3__6949_, data_stage_3__6948_, data_stage_3__6947_, data_stage_3__6946_, data_stage_3__6945_, data_stage_3__6944_, data_stage_3__6943_, data_stage_3__6942_, data_stage_3__6941_, data_stage_3__6940_, data_stage_3__6939_, data_stage_3__6938_, data_stage_3__6937_, data_stage_3__6936_, data_stage_3__6935_, data_stage_3__6934_, data_stage_3__6933_, data_stage_3__6932_, data_stage_3__6931_, data_stage_3__6930_, data_stage_3__6929_, data_stage_3__6928_, data_stage_3__6927_, data_stage_3__6926_, data_stage_3__6925_, data_stage_3__6924_, data_stage_3__6923_, data_stage_3__6922_, data_stage_3__6921_, data_stage_3__6920_, data_stage_3__6919_, data_stage_3__6918_, data_stage_3__6917_, data_stage_3__6916_, data_stage_3__6915_, data_stage_3__6914_, data_stage_3__6913_, data_stage_3__6912_, data_stage_3__6911_, data_stage_3__6910_, data_stage_3__6909_, data_stage_3__6908_, data_stage_3__6907_, data_stage_3__6906_, data_stage_3__6905_, data_stage_3__6904_, data_stage_3__6903_, data_stage_3__6902_, data_stage_3__6901_, data_stage_3__6900_, data_stage_3__6899_, data_stage_3__6898_, data_stage_3__6897_, data_stage_3__6896_, data_stage_3__6895_, data_stage_3__6894_, data_stage_3__6893_, data_stage_3__6892_, data_stage_3__6891_, data_stage_3__6890_, data_stage_3__6889_, data_stage_3__6888_, data_stage_3__6887_, data_stage_3__6886_, data_stage_3__6885_, data_stage_3__6884_, data_stage_3__6883_, data_stage_3__6882_, data_stage_3__6881_, data_stage_3__6880_, data_stage_3__6879_, data_stage_3__6878_, data_stage_3__6877_, data_stage_3__6876_, data_stage_3__6875_, data_stage_3__6874_, data_stage_3__6873_, data_stage_3__6872_, data_stage_3__6871_, data_stage_3__6870_, data_stage_3__6869_, data_stage_3__6868_, data_stage_3__6867_, data_stage_3__6866_, data_stage_3__6865_, data_stage_3__6864_, data_stage_3__6863_, data_stage_3__6862_, data_stage_3__6861_, data_stage_3__6860_, data_stage_3__6859_, data_stage_3__6858_, data_stage_3__6857_, data_stage_3__6856_, data_stage_3__6855_, data_stage_3__6854_, data_stage_3__6853_, data_stage_3__6852_, data_stage_3__6851_, data_stage_3__6850_, data_stage_3__6849_, data_stage_3__6848_, data_stage_3__6847_, data_stage_3__6846_, data_stage_3__6845_, data_stage_3__6844_, data_stage_3__6843_, data_stage_3__6842_, data_stage_3__6841_, data_stage_3__6840_, data_stage_3__6839_, data_stage_3__6838_, data_stage_3__6837_, data_stage_3__6836_, data_stage_3__6835_, data_stage_3__6834_, data_stage_3__6833_, data_stage_3__6832_, data_stage_3__6831_, data_stage_3__6830_, data_stage_3__6829_, data_stage_3__6828_, data_stage_3__6827_, data_stage_3__6826_, data_stage_3__6825_, data_stage_3__6824_, data_stage_3__6823_, data_stage_3__6822_, data_stage_3__6821_, data_stage_3__6820_, data_stage_3__6819_, data_stage_3__6818_, data_stage_3__6817_, data_stage_3__6816_, data_stage_3__6815_, data_stage_3__6814_, data_stage_3__6813_, data_stage_3__6812_, data_stage_3__6811_, data_stage_3__6810_, data_stage_3__6809_, data_stage_3__6808_, data_stage_3__6807_, data_stage_3__6806_, data_stage_3__6805_, data_stage_3__6804_, data_stage_3__6803_, data_stage_3__6802_, data_stage_3__6801_, data_stage_3__6800_, data_stage_3__6799_, data_stage_3__6798_, data_stage_3__6797_, data_stage_3__6796_, data_stage_3__6795_, data_stage_3__6794_, data_stage_3__6793_, data_stage_3__6792_, data_stage_3__6791_, data_stage_3__6790_, data_stage_3__6789_, data_stage_3__6788_, data_stage_3__6787_, data_stage_3__6786_, data_stage_3__6785_, data_stage_3__6784_, data_stage_3__6783_, data_stage_3__6782_, data_stage_3__6781_, data_stage_3__6780_, data_stage_3__6779_, data_stage_3__6778_, data_stage_3__6777_, data_stage_3__6776_, data_stage_3__6775_, data_stage_3__6774_, data_stage_3__6773_, data_stage_3__6772_, data_stage_3__6771_, data_stage_3__6770_, data_stage_3__6769_, data_stage_3__6768_, data_stage_3__6767_, data_stage_3__6766_, data_stage_3__6765_, data_stage_3__6764_, data_stage_3__6763_, data_stage_3__6762_, data_stage_3__6761_, data_stage_3__6760_, data_stage_3__6759_, data_stage_3__6758_, data_stage_3__6757_, data_stage_3__6756_, data_stage_3__6755_, data_stage_3__6754_, data_stage_3__6753_, data_stage_3__6752_, data_stage_3__6751_, data_stage_3__6750_, data_stage_3__6749_, data_stage_3__6748_, data_stage_3__6747_, data_stage_3__6746_, data_stage_3__6745_, data_stage_3__6744_, data_stage_3__6743_, data_stage_3__6742_, data_stage_3__6741_, data_stage_3__6740_, data_stage_3__6739_, data_stage_3__6738_, data_stage_3__6737_, data_stage_3__6736_, data_stage_3__6735_, data_stage_3__6734_, data_stage_3__6733_, data_stage_3__6732_, data_stage_3__6731_, data_stage_3__6730_, data_stage_3__6729_, data_stage_3__6728_, data_stage_3__6727_, data_stage_3__6726_, data_stage_3__6725_, data_stage_3__6724_, data_stage_3__6723_, data_stage_3__6722_, data_stage_3__6721_, data_stage_3__6720_, data_stage_3__6719_, data_stage_3__6718_, data_stage_3__6717_, data_stage_3__6716_, data_stage_3__6715_, data_stage_3__6714_, data_stage_3__6713_, data_stage_3__6712_, data_stage_3__6711_, data_stage_3__6710_, data_stage_3__6709_, data_stage_3__6708_, data_stage_3__6707_, data_stage_3__6706_, data_stage_3__6705_, data_stage_3__6704_, data_stage_3__6703_, data_stage_3__6702_, data_stage_3__6701_, data_stage_3__6700_, data_stage_3__6699_, data_stage_3__6698_, data_stage_3__6697_, data_stage_3__6696_, data_stage_3__6695_, data_stage_3__6694_, data_stage_3__6693_, data_stage_3__6692_, data_stage_3__6691_, data_stage_3__6690_, data_stage_3__6689_, data_stage_3__6688_, data_stage_3__6687_, data_stage_3__6686_, data_stage_3__6685_, data_stage_3__6684_, data_stage_3__6683_, data_stage_3__6682_, data_stage_3__6681_, data_stage_3__6680_, data_stage_3__6679_, data_stage_3__6678_, data_stage_3__6677_, data_stage_3__6676_, data_stage_3__6675_, data_stage_3__6674_, data_stage_3__6673_, data_stage_3__6672_, data_stage_3__6671_, data_stage_3__6670_, data_stage_3__6669_, data_stage_3__6668_, data_stage_3__6667_, data_stage_3__6666_, data_stage_3__6665_, data_stage_3__6664_, data_stage_3__6663_, data_stage_3__6662_, data_stage_3__6661_, data_stage_3__6660_, data_stage_3__6659_, data_stage_3__6658_, data_stage_3__6657_, data_stage_3__6656_, data_stage_3__6655_, data_stage_3__6654_, data_stage_3__6653_, data_stage_3__6652_, data_stage_3__6651_, data_stage_3__6650_, data_stage_3__6649_, data_stage_3__6648_, data_stage_3__6647_, data_stage_3__6646_, data_stage_3__6645_, data_stage_3__6644_, data_stage_3__6643_, data_stage_3__6642_, data_stage_3__6641_, data_stage_3__6640_, data_stage_3__6639_, data_stage_3__6638_, data_stage_3__6637_, data_stage_3__6636_, data_stage_3__6635_, data_stage_3__6634_, data_stage_3__6633_, data_stage_3__6632_, data_stage_3__6631_, data_stage_3__6630_, data_stage_3__6629_, data_stage_3__6628_, data_stage_3__6627_, data_stage_3__6626_, data_stage_3__6625_, data_stage_3__6624_, data_stage_3__6623_, data_stage_3__6622_, data_stage_3__6621_, data_stage_3__6620_, data_stage_3__6619_, data_stage_3__6618_, data_stage_3__6617_, data_stage_3__6616_, data_stage_3__6615_, data_stage_3__6614_, data_stage_3__6613_, data_stage_3__6612_, data_stage_3__6611_, data_stage_3__6610_, data_stage_3__6609_, data_stage_3__6608_, data_stage_3__6607_, data_stage_3__6606_, data_stage_3__6605_, data_stage_3__6604_, data_stage_3__6603_, data_stage_3__6602_, data_stage_3__6601_, data_stage_3__6600_, data_stage_3__6599_, data_stage_3__6598_, data_stage_3__6597_, data_stage_3__6596_, data_stage_3__6595_, data_stage_3__6594_, data_stage_3__6593_, data_stage_3__6592_, data_stage_3__6591_, data_stage_3__6590_, data_stage_3__6589_, data_stage_3__6588_, data_stage_3__6587_, data_stage_3__6586_, data_stage_3__6585_, data_stage_3__6584_, data_stage_3__6583_, data_stage_3__6582_, data_stage_3__6581_, data_stage_3__6580_, data_stage_3__6579_, data_stage_3__6578_, data_stage_3__6577_, data_stage_3__6576_, data_stage_3__6575_, data_stage_3__6574_, data_stage_3__6573_, data_stage_3__6572_, data_stage_3__6571_, data_stage_3__6570_, data_stage_3__6569_, data_stage_3__6568_, data_stage_3__6567_, data_stage_3__6566_, data_stage_3__6565_, data_stage_3__6564_, data_stage_3__6563_, data_stage_3__6562_, data_stage_3__6561_, data_stage_3__6560_, data_stage_3__6559_, data_stage_3__6558_, data_stage_3__6557_, data_stage_3__6556_, data_stage_3__6555_, data_stage_3__6554_, data_stage_3__6553_, data_stage_3__6552_, data_stage_3__6551_, data_stage_3__6550_, data_stage_3__6549_, data_stage_3__6548_, data_stage_3__6547_, data_stage_3__6546_, data_stage_3__6545_, data_stage_3__6544_, data_stage_3__6543_, data_stage_3__6542_, data_stage_3__6541_, data_stage_3__6540_, data_stage_3__6539_, data_stage_3__6538_, data_stage_3__6537_, data_stage_3__6536_, data_stage_3__6535_, data_stage_3__6534_, data_stage_3__6533_, data_stage_3__6532_, data_stage_3__6531_, data_stage_3__6530_, data_stage_3__6529_, data_stage_3__6528_, data_stage_3__6527_, data_stage_3__6526_, data_stage_3__6525_, data_stage_3__6524_, data_stage_3__6523_, data_stage_3__6522_, data_stage_3__6521_, data_stage_3__6520_, data_stage_3__6519_, data_stage_3__6518_, data_stage_3__6517_, data_stage_3__6516_, data_stage_3__6515_, data_stage_3__6514_, data_stage_3__6513_, data_stage_3__6512_, data_stage_3__6511_, data_stage_3__6510_, data_stage_3__6509_, data_stage_3__6508_, data_stage_3__6507_, data_stage_3__6506_, data_stage_3__6505_, data_stage_3__6504_, data_stage_3__6503_, data_stage_3__6502_, data_stage_3__6501_, data_stage_3__6500_, data_stage_3__6499_, data_stage_3__6498_, data_stage_3__6497_, data_stage_3__6496_, data_stage_3__6495_, data_stage_3__6494_, data_stage_3__6493_, data_stage_3__6492_, data_stage_3__6491_, data_stage_3__6490_, data_stage_3__6489_, data_stage_3__6488_, data_stage_3__6487_, data_stage_3__6486_, data_stage_3__6485_, data_stage_3__6484_, data_stage_3__6483_, data_stage_3__6482_, data_stage_3__6481_, data_stage_3__6480_, data_stage_3__6479_, data_stage_3__6478_, data_stage_3__6477_, data_stage_3__6476_, data_stage_3__6475_, data_stage_3__6474_, data_stage_3__6473_, data_stage_3__6472_, data_stage_3__6471_, data_stage_3__6470_, data_stage_3__6469_, data_stage_3__6468_, data_stage_3__6467_, data_stage_3__6466_, data_stage_3__6465_, data_stage_3__6464_, data_stage_3__6463_, data_stage_3__6462_, data_stage_3__6461_, data_stage_3__6460_, data_stage_3__6459_, data_stage_3__6458_, data_stage_3__6457_, data_stage_3__6456_, data_stage_3__6455_, data_stage_3__6454_, data_stage_3__6453_, data_stage_3__6452_, data_stage_3__6451_, data_stage_3__6450_, data_stage_3__6449_, data_stage_3__6448_, data_stage_3__6447_, data_stage_3__6446_, data_stage_3__6445_, data_stage_3__6444_, data_stage_3__6443_, data_stage_3__6442_, data_stage_3__6441_, data_stage_3__6440_, data_stage_3__6439_, data_stage_3__6438_, data_stage_3__6437_, data_stage_3__6436_, data_stage_3__6435_, data_stage_3__6434_, data_stage_3__6433_, data_stage_3__6432_, data_stage_3__6431_, data_stage_3__6430_, data_stage_3__6429_, data_stage_3__6428_, data_stage_3__6427_, data_stage_3__6426_, data_stage_3__6425_, data_stage_3__6424_, data_stage_3__6423_, data_stage_3__6422_, data_stage_3__6421_, data_stage_3__6420_, data_stage_3__6419_, data_stage_3__6418_, data_stage_3__6417_, data_stage_3__6416_, data_stage_3__6415_, data_stage_3__6414_, data_stage_3__6413_, data_stage_3__6412_, data_stage_3__6411_, data_stage_3__6410_, data_stage_3__6409_, data_stage_3__6408_, data_stage_3__6407_, data_stage_3__6406_, data_stage_3__6405_, data_stage_3__6404_, data_stage_3__6403_, data_stage_3__6402_, data_stage_3__6401_, data_stage_3__6400_, data_stage_3__6399_, data_stage_3__6398_, data_stage_3__6397_, data_stage_3__6396_, data_stage_3__6395_, data_stage_3__6394_, data_stage_3__6393_, data_stage_3__6392_, data_stage_3__6391_, data_stage_3__6390_, data_stage_3__6389_, data_stage_3__6388_, data_stage_3__6387_, data_stage_3__6386_, data_stage_3__6385_, data_stage_3__6384_, data_stage_3__6383_, data_stage_3__6382_, data_stage_3__6381_, data_stage_3__6380_, data_stage_3__6379_, data_stage_3__6378_, data_stage_3__6377_, data_stage_3__6376_, data_stage_3__6375_, data_stage_3__6374_, data_stage_3__6373_, data_stage_3__6372_, data_stage_3__6371_, data_stage_3__6370_, data_stage_3__6369_, data_stage_3__6368_, data_stage_3__6367_, data_stage_3__6366_, data_stage_3__6365_, data_stage_3__6364_, data_stage_3__6363_, data_stage_3__6362_, data_stage_3__6361_, data_stage_3__6360_, data_stage_3__6359_, data_stage_3__6358_, data_stage_3__6357_, data_stage_3__6356_, data_stage_3__6355_, data_stage_3__6354_, data_stage_3__6353_, data_stage_3__6352_, data_stage_3__6351_, data_stage_3__6350_, data_stage_3__6349_, data_stage_3__6348_, data_stage_3__6347_, data_stage_3__6346_, data_stage_3__6345_, data_stage_3__6344_, data_stage_3__6343_, data_stage_3__6342_, data_stage_3__6341_, data_stage_3__6340_, data_stage_3__6339_, data_stage_3__6338_, data_stage_3__6337_, data_stage_3__6336_, data_stage_3__6335_, data_stage_3__6334_, data_stage_3__6333_, data_stage_3__6332_, data_stage_3__6331_, data_stage_3__6330_, data_stage_3__6329_, data_stage_3__6328_, data_stage_3__6327_, data_stage_3__6326_, data_stage_3__6325_, data_stage_3__6324_, data_stage_3__6323_, data_stage_3__6322_, data_stage_3__6321_, data_stage_3__6320_, data_stage_3__6319_, data_stage_3__6318_, data_stage_3__6317_, data_stage_3__6316_, data_stage_3__6315_, data_stage_3__6314_, data_stage_3__6313_, data_stage_3__6312_, data_stage_3__6311_, data_stage_3__6310_, data_stage_3__6309_, data_stage_3__6308_, data_stage_3__6307_, data_stage_3__6306_, data_stage_3__6305_, data_stage_3__6304_, data_stage_3__6303_, data_stage_3__6302_, data_stage_3__6301_, data_stage_3__6300_, data_stage_3__6299_, data_stage_3__6298_, data_stage_3__6297_, data_stage_3__6296_, data_stage_3__6295_, data_stage_3__6294_, data_stage_3__6293_, data_stage_3__6292_, data_stage_3__6291_, data_stage_3__6290_, data_stage_3__6289_, data_stage_3__6288_, data_stage_3__6287_, data_stage_3__6286_, data_stage_3__6285_, data_stage_3__6284_, data_stage_3__6283_, data_stage_3__6282_, data_stage_3__6281_, data_stage_3__6280_, data_stage_3__6279_, data_stage_3__6278_, data_stage_3__6277_, data_stage_3__6276_, data_stage_3__6275_, data_stage_3__6274_, data_stage_3__6273_, data_stage_3__6272_, data_stage_3__6271_, data_stage_3__6270_, data_stage_3__6269_, data_stage_3__6268_, data_stage_3__6267_, data_stage_3__6266_, data_stage_3__6265_, data_stage_3__6264_, data_stage_3__6263_, data_stage_3__6262_, data_stage_3__6261_, data_stage_3__6260_, data_stage_3__6259_, data_stage_3__6258_, data_stage_3__6257_, data_stage_3__6256_, data_stage_3__6255_, data_stage_3__6254_, data_stage_3__6253_, data_stage_3__6252_, data_stage_3__6251_, data_stage_3__6250_, data_stage_3__6249_, data_stage_3__6248_, data_stage_3__6247_, data_stage_3__6246_, data_stage_3__6245_, data_stage_3__6244_, data_stage_3__6243_, data_stage_3__6242_, data_stage_3__6241_, data_stage_3__6240_, data_stage_3__6239_, data_stage_3__6238_, data_stage_3__6237_, data_stage_3__6236_, data_stage_3__6235_, data_stage_3__6234_, data_stage_3__6233_, data_stage_3__6232_, data_stage_3__6231_, data_stage_3__6230_, data_stage_3__6229_, data_stage_3__6228_, data_stage_3__6227_, data_stage_3__6226_, data_stage_3__6225_, data_stage_3__6224_, data_stage_3__6223_, data_stage_3__6222_, data_stage_3__6221_, data_stage_3__6220_, data_stage_3__6219_, data_stage_3__6218_, data_stage_3__6217_, data_stage_3__6216_, data_stage_3__6215_, data_stage_3__6214_, data_stage_3__6213_, data_stage_3__6212_, data_stage_3__6211_, data_stage_3__6210_, data_stage_3__6209_, data_stage_3__6208_, data_stage_3__6207_, data_stage_3__6206_, data_stage_3__6205_, data_stage_3__6204_, data_stage_3__6203_, data_stage_3__6202_, data_stage_3__6201_, data_stage_3__6200_, data_stage_3__6199_, data_stage_3__6198_, data_stage_3__6197_, data_stage_3__6196_, data_stage_3__6195_, data_stage_3__6194_, data_stage_3__6193_, data_stage_3__6192_, data_stage_3__6191_, data_stage_3__6190_, data_stage_3__6189_, data_stage_3__6188_, data_stage_3__6187_, data_stage_3__6186_, data_stage_3__6185_, data_stage_3__6184_, data_stage_3__6183_, data_stage_3__6182_, data_stage_3__6181_, data_stage_3__6180_, data_stage_3__6179_, data_stage_3__6178_, data_stage_3__6177_, data_stage_3__6176_, data_stage_3__6175_, data_stage_3__6174_, data_stage_3__6173_, data_stage_3__6172_, data_stage_3__6171_, data_stage_3__6170_, data_stage_3__6169_, data_stage_3__6168_, data_stage_3__6167_, data_stage_3__6166_, data_stage_3__6165_, data_stage_3__6164_, data_stage_3__6163_, data_stage_3__6162_, data_stage_3__6161_, data_stage_3__6160_, data_stage_3__6159_, data_stage_3__6158_, data_stage_3__6157_, data_stage_3__6156_, data_stage_3__6155_, data_stage_3__6154_, data_stage_3__6153_, data_stage_3__6152_, data_stage_3__6151_, data_stage_3__6150_, data_stage_3__6149_, data_stage_3__6148_, data_stage_3__6147_, data_stage_3__6146_, data_stage_3__6145_, data_stage_3__6144_ })
  );


  bsg_swap_width_p512
  mux_stage_2__mux_swap_7__swap_inst
  (
    .data_i({ data_stage_2__8191_, data_stage_2__8190_, data_stage_2__8189_, data_stage_2__8188_, data_stage_2__8187_, data_stage_2__8186_, data_stage_2__8185_, data_stage_2__8184_, data_stage_2__8183_, data_stage_2__8182_, data_stage_2__8181_, data_stage_2__8180_, data_stage_2__8179_, data_stage_2__8178_, data_stage_2__8177_, data_stage_2__8176_, data_stage_2__8175_, data_stage_2__8174_, data_stage_2__8173_, data_stage_2__8172_, data_stage_2__8171_, data_stage_2__8170_, data_stage_2__8169_, data_stage_2__8168_, data_stage_2__8167_, data_stage_2__8166_, data_stage_2__8165_, data_stage_2__8164_, data_stage_2__8163_, data_stage_2__8162_, data_stage_2__8161_, data_stage_2__8160_, data_stage_2__8159_, data_stage_2__8158_, data_stage_2__8157_, data_stage_2__8156_, data_stage_2__8155_, data_stage_2__8154_, data_stage_2__8153_, data_stage_2__8152_, data_stage_2__8151_, data_stage_2__8150_, data_stage_2__8149_, data_stage_2__8148_, data_stage_2__8147_, data_stage_2__8146_, data_stage_2__8145_, data_stage_2__8144_, data_stage_2__8143_, data_stage_2__8142_, data_stage_2__8141_, data_stage_2__8140_, data_stage_2__8139_, data_stage_2__8138_, data_stage_2__8137_, data_stage_2__8136_, data_stage_2__8135_, data_stage_2__8134_, data_stage_2__8133_, data_stage_2__8132_, data_stage_2__8131_, data_stage_2__8130_, data_stage_2__8129_, data_stage_2__8128_, data_stage_2__8127_, data_stage_2__8126_, data_stage_2__8125_, data_stage_2__8124_, data_stage_2__8123_, data_stage_2__8122_, data_stage_2__8121_, data_stage_2__8120_, data_stage_2__8119_, data_stage_2__8118_, data_stage_2__8117_, data_stage_2__8116_, data_stage_2__8115_, data_stage_2__8114_, data_stage_2__8113_, data_stage_2__8112_, data_stage_2__8111_, data_stage_2__8110_, data_stage_2__8109_, data_stage_2__8108_, data_stage_2__8107_, data_stage_2__8106_, data_stage_2__8105_, data_stage_2__8104_, data_stage_2__8103_, data_stage_2__8102_, data_stage_2__8101_, data_stage_2__8100_, data_stage_2__8099_, data_stage_2__8098_, data_stage_2__8097_, data_stage_2__8096_, data_stage_2__8095_, data_stage_2__8094_, data_stage_2__8093_, data_stage_2__8092_, data_stage_2__8091_, data_stage_2__8090_, data_stage_2__8089_, data_stage_2__8088_, data_stage_2__8087_, data_stage_2__8086_, data_stage_2__8085_, data_stage_2__8084_, data_stage_2__8083_, data_stage_2__8082_, data_stage_2__8081_, data_stage_2__8080_, data_stage_2__8079_, data_stage_2__8078_, data_stage_2__8077_, data_stage_2__8076_, data_stage_2__8075_, data_stage_2__8074_, data_stage_2__8073_, data_stage_2__8072_, data_stage_2__8071_, data_stage_2__8070_, data_stage_2__8069_, data_stage_2__8068_, data_stage_2__8067_, data_stage_2__8066_, data_stage_2__8065_, data_stage_2__8064_, data_stage_2__8063_, data_stage_2__8062_, data_stage_2__8061_, data_stage_2__8060_, data_stage_2__8059_, data_stage_2__8058_, data_stage_2__8057_, data_stage_2__8056_, data_stage_2__8055_, data_stage_2__8054_, data_stage_2__8053_, data_stage_2__8052_, data_stage_2__8051_, data_stage_2__8050_, data_stage_2__8049_, data_stage_2__8048_, data_stage_2__8047_, data_stage_2__8046_, data_stage_2__8045_, data_stage_2__8044_, data_stage_2__8043_, data_stage_2__8042_, data_stage_2__8041_, data_stage_2__8040_, data_stage_2__8039_, data_stage_2__8038_, data_stage_2__8037_, data_stage_2__8036_, data_stage_2__8035_, data_stage_2__8034_, data_stage_2__8033_, data_stage_2__8032_, data_stage_2__8031_, data_stage_2__8030_, data_stage_2__8029_, data_stage_2__8028_, data_stage_2__8027_, data_stage_2__8026_, data_stage_2__8025_, data_stage_2__8024_, data_stage_2__8023_, data_stage_2__8022_, data_stage_2__8021_, data_stage_2__8020_, data_stage_2__8019_, data_stage_2__8018_, data_stage_2__8017_, data_stage_2__8016_, data_stage_2__8015_, data_stage_2__8014_, data_stage_2__8013_, data_stage_2__8012_, data_stage_2__8011_, data_stage_2__8010_, data_stage_2__8009_, data_stage_2__8008_, data_stage_2__8007_, data_stage_2__8006_, data_stage_2__8005_, data_stage_2__8004_, data_stage_2__8003_, data_stage_2__8002_, data_stage_2__8001_, data_stage_2__8000_, data_stage_2__7999_, data_stage_2__7998_, data_stage_2__7997_, data_stage_2__7996_, data_stage_2__7995_, data_stage_2__7994_, data_stage_2__7993_, data_stage_2__7992_, data_stage_2__7991_, data_stage_2__7990_, data_stage_2__7989_, data_stage_2__7988_, data_stage_2__7987_, data_stage_2__7986_, data_stage_2__7985_, data_stage_2__7984_, data_stage_2__7983_, data_stage_2__7982_, data_stage_2__7981_, data_stage_2__7980_, data_stage_2__7979_, data_stage_2__7978_, data_stage_2__7977_, data_stage_2__7976_, data_stage_2__7975_, data_stage_2__7974_, data_stage_2__7973_, data_stage_2__7972_, data_stage_2__7971_, data_stage_2__7970_, data_stage_2__7969_, data_stage_2__7968_, data_stage_2__7967_, data_stage_2__7966_, data_stage_2__7965_, data_stage_2__7964_, data_stage_2__7963_, data_stage_2__7962_, data_stage_2__7961_, data_stage_2__7960_, data_stage_2__7959_, data_stage_2__7958_, data_stage_2__7957_, data_stage_2__7956_, data_stage_2__7955_, data_stage_2__7954_, data_stage_2__7953_, data_stage_2__7952_, data_stage_2__7951_, data_stage_2__7950_, data_stage_2__7949_, data_stage_2__7948_, data_stage_2__7947_, data_stage_2__7946_, data_stage_2__7945_, data_stage_2__7944_, data_stage_2__7943_, data_stage_2__7942_, data_stage_2__7941_, data_stage_2__7940_, data_stage_2__7939_, data_stage_2__7938_, data_stage_2__7937_, data_stage_2__7936_, data_stage_2__7935_, data_stage_2__7934_, data_stage_2__7933_, data_stage_2__7932_, data_stage_2__7931_, data_stage_2__7930_, data_stage_2__7929_, data_stage_2__7928_, data_stage_2__7927_, data_stage_2__7926_, data_stage_2__7925_, data_stage_2__7924_, data_stage_2__7923_, data_stage_2__7922_, data_stage_2__7921_, data_stage_2__7920_, data_stage_2__7919_, data_stage_2__7918_, data_stage_2__7917_, data_stage_2__7916_, data_stage_2__7915_, data_stage_2__7914_, data_stage_2__7913_, data_stage_2__7912_, data_stage_2__7911_, data_stage_2__7910_, data_stage_2__7909_, data_stage_2__7908_, data_stage_2__7907_, data_stage_2__7906_, data_stage_2__7905_, data_stage_2__7904_, data_stage_2__7903_, data_stage_2__7902_, data_stage_2__7901_, data_stage_2__7900_, data_stage_2__7899_, data_stage_2__7898_, data_stage_2__7897_, data_stage_2__7896_, data_stage_2__7895_, data_stage_2__7894_, data_stage_2__7893_, data_stage_2__7892_, data_stage_2__7891_, data_stage_2__7890_, data_stage_2__7889_, data_stage_2__7888_, data_stage_2__7887_, data_stage_2__7886_, data_stage_2__7885_, data_stage_2__7884_, data_stage_2__7883_, data_stage_2__7882_, data_stage_2__7881_, data_stage_2__7880_, data_stage_2__7879_, data_stage_2__7878_, data_stage_2__7877_, data_stage_2__7876_, data_stage_2__7875_, data_stage_2__7874_, data_stage_2__7873_, data_stage_2__7872_, data_stage_2__7871_, data_stage_2__7870_, data_stage_2__7869_, data_stage_2__7868_, data_stage_2__7867_, data_stage_2__7866_, data_stage_2__7865_, data_stage_2__7864_, data_stage_2__7863_, data_stage_2__7862_, data_stage_2__7861_, data_stage_2__7860_, data_stage_2__7859_, data_stage_2__7858_, data_stage_2__7857_, data_stage_2__7856_, data_stage_2__7855_, data_stage_2__7854_, data_stage_2__7853_, data_stage_2__7852_, data_stage_2__7851_, data_stage_2__7850_, data_stage_2__7849_, data_stage_2__7848_, data_stage_2__7847_, data_stage_2__7846_, data_stage_2__7845_, data_stage_2__7844_, data_stage_2__7843_, data_stage_2__7842_, data_stage_2__7841_, data_stage_2__7840_, data_stage_2__7839_, data_stage_2__7838_, data_stage_2__7837_, data_stage_2__7836_, data_stage_2__7835_, data_stage_2__7834_, data_stage_2__7833_, data_stage_2__7832_, data_stage_2__7831_, data_stage_2__7830_, data_stage_2__7829_, data_stage_2__7828_, data_stage_2__7827_, data_stage_2__7826_, data_stage_2__7825_, data_stage_2__7824_, data_stage_2__7823_, data_stage_2__7822_, data_stage_2__7821_, data_stage_2__7820_, data_stage_2__7819_, data_stage_2__7818_, data_stage_2__7817_, data_stage_2__7816_, data_stage_2__7815_, data_stage_2__7814_, data_stage_2__7813_, data_stage_2__7812_, data_stage_2__7811_, data_stage_2__7810_, data_stage_2__7809_, data_stage_2__7808_, data_stage_2__7807_, data_stage_2__7806_, data_stage_2__7805_, data_stage_2__7804_, data_stage_2__7803_, data_stage_2__7802_, data_stage_2__7801_, data_stage_2__7800_, data_stage_2__7799_, data_stage_2__7798_, data_stage_2__7797_, data_stage_2__7796_, data_stage_2__7795_, data_stage_2__7794_, data_stage_2__7793_, data_stage_2__7792_, data_stage_2__7791_, data_stage_2__7790_, data_stage_2__7789_, data_stage_2__7788_, data_stage_2__7787_, data_stage_2__7786_, data_stage_2__7785_, data_stage_2__7784_, data_stage_2__7783_, data_stage_2__7782_, data_stage_2__7781_, data_stage_2__7780_, data_stage_2__7779_, data_stage_2__7778_, data_stage_2__7777_, data_stage_2__7776_, data_stage_2__7775_, data_stage_2__7774_, data_stage_2__7773_, data_stage_2__7772_, data_stage_2__7771_, data_stage_2__7770_, data_stage_2__7769_, data_stage_2__7768_, data_stage_2__7767_, data_stage_2__7766_, data_stage_2__7765_, data_stage_2__7764_, data_stage_2__7763_, data_stage_2__7762_, data_stage_2__7761_, data_stage_2__7760_, data_stage_2__7759_, data_stage_2__7758_, data_stage_2__7757_, data_stage_2__7756_, data_stage_2__7755_, data_stage_2__7754_, data_stage_2__7753_, data_stage_2__7752_, data_stage_2__7751_, data_stage_2__7750_, data_stage_2__7749_, data_stage_2__7748_, data_stage_2__7747_, data_stage_2__7746_, data_stage_2__7745_, data_stage_2__7744_, data_stage_2__7743_, data_stage_2__7742_, data_stage_2__7741_, data_stage_2__7740_, data_stage_2__7739_, data_stage_2__7738_, data_stage_2__7737_, data_stage_2__7736_, data_stage_2__7735_, data_stage_2__7734_, data_stage_2__7733_, data_stage_2__7732_, data_stage_2__7731_, data_stage_2__7730_, data_stage_2__7729_, data_stage_2__7728_, data_stage_2__7727_, data_stage_2__7726_, data_stage_2__7725_, data_stage_2__7724_, data_stage_2__7723_, data_stage_2__7722_, data_stage_2__7721_, data_stage_2__7720_, data_stage_2__7719_, data_stage_2__7718_, data_stage_2__7717_, data_stage_2__7716_, data_stage_2__7715_, data_stage_2__7714_, data_stage_2__7713_, data_stage_2__7712_, data_stage_2__7711_, data_stage_2__7710_, data_stage_2__7709_, data_stage_2__7708_, data_stage_2__7707_, data_stage_2__7706_, data_stage_2__7705_, data_stage_2__7704_, data_stage_2__7703_, data_stage_2__7702_, data_stage_2__7701_, data_stage_2__7700_, data_stage_2__7699_, data_stage_2__7698_, data_stage_2__7697_, data_stage_2__7696_, data_stage_2__7695_, data_stage_2__7694_, data_stage_2__7693_, data_stage_2__7692_, data_stage_2__7691_, data_stage_2__7690_, data_stage_2__7689_, data_stage_2__7688_, data_stage_2__7687_, data_stage_2__7686_, data_stage_2__7685_, data_stage_2__7684_, data_stage_2__7683_, data_stage_2__7682_, data_stage_2__7681_, data_stage_2__7680_, data_stage_2__7679_, data_stage_2__7678_, data_stage_2__7677_, data_stage_2__7676_, data_stage_2__7675_, data_stage_2__7674_, data_stage_2__7673_, data_stage_2__7672_, data_stage_2__7671_, data_stage_2__7670_, data_stage_2__7669_, data_stage_2__7668_, data_stage_2__7667_, data_stage_2__7666_, data_stage_2__7665_, data_stage_2__7664_, data_stage_2__7663_, data_stage_2__7662_, data_stage_2__7661_, data_stage_2__7660_, data_stage_2__7659_, data_stage_2__7658_, data_stage_2__7657_, data_stage_2__7656_, data_stage_2__7655_, data_stage_2__7654_, data_stage_2__7653_, data_stage_2__7652_, data_stage_2__7651_, data_stage_2__7650_, data_stage_2__7649_, data_stage_2__7648_, data_stage_2__7647_, data_stage_2__7646_, data_stage_2__7645_, data_stage_2__7644_, data_stage_2__7643_, data_stage_2__7642_, data_stage_2__7641_, data_stage_2__7640_, data_stage_2__7639_, data_stage_2__7638_, data_stage_2__7637_, data_stage_2__7636_, data_stage_2__7635_, data_stage_2__7634_, data_stage_2__7633_, data_stage_2__7632_, data_stage_2__7631_, data_stage_2__7630_, data_stage_2__7629_, data_stage_2__7628_, data_stage_2__7627_, data_stage_2__7626_, data_stage_2__7625_, data_stage_2__7624_, data_stage_2__7623_, data_stage_2__7622_, data_stage_2__7621_, data_stage_2__7620_, data_stage_2__7619_, data_stage_2__7618_, data_stage_2__7617_, data_stage_2__7616_, data_stage_2__7615_, data_stage_2__7614_, data_stage_2__7613_, data_stage_2__7612_, data_stage_2__7611_, data_stage_2__7610_, data_stage_2__7609_, data_stage_2__7608_, data_stage_2__7607_, data_stage_2__7606_, data_stage_2__7605_, data_stage_2__7604_, data_stage_2__7603_, data_stage_2__7602_, data_stage_2__7601_, data_stage_2__7600_, data_stage_2__7599_, data_stage_2__7598_, data_stage_2__7597_, data_stage_2__7596_, data_stage_2__7595_, data_stage_2__7594_, data_stage_2__7593_, data_stage_2__7592_, data_stage_2__7591_, data_stage_2__7590_, data_stage_2__7589_, data_stage_2__7588_, data_stage_2__7587_, data_stage_2__7586_, data_stage_2__7585_, data_stage_2__7584_, data_stage_2__7583_, data_stage_2__7582_, data_stage_2__7581_, data_stage_2__7580_, data_stage_2__7579_, data_stage_2__7578_, data_stage_2__7577_, data_stage_2__7576_, data_stage_2__7575_, data_stage_2__7574_, data_stage_2__7573_, data_stage_2__7572_, data_stage_2__7571_, data_stage_2__7570_, data_stage_2__7569_, data_stage_2__7568_, data_stage_2__7567_, data_stage_2__7566_, data_stage_2__7565_, data_stage_2__7564_, data_stage_2__7563_, data_stage_2__7562_, data_stage_2__7561_, data_stage_2__7560_, data_stage_2__7559_, data_stage_2__7558_, data_stage_2__7557_, data_stage_2__7556_, data_stage_2__7555_, data_stage_2__7554_, data_stage_2__7553_, data_stage_2__7552_, data_stage_2__7551_, data_stage_2__7550_, data_stage_2__7549_, data_stage_2__7548_, data_stage_2__7547_, data_stage_2__7546_, data_stage_2__7545_, data_stage_2__7544_, data_stage_2__7543_, data_stage_2__7542_, data_stage_2__7541_, data_stage_2__7540_, data_stage_2__7539_, data_stage_2__7538_, data_stage_2__7537_, data_stage_2__7536_, data_stage_2__7535_, data_stage_2__7534_, data_stage_2__7533_, data_stage_2__7532_, data_stage_2__7531_, data_stage_2__7530_, data_stage_2__7529_, data_stage_2__7528_, data_stage_2__7527_, data_stage_2__7526_, data_stage_2__7525_, data_stage_2__7524_, data_stage_2__7523_, data_stage_2__7522_, data_stage_2__7521_, data_stage_2__7520_, data_stage_2__7519_, data_stage_2__7518_, data_stage_2__7517_, data_stage_2__7516_, data_stage_2__7515_, data_stage_2__7514_, data_stage_2__7513_, data_stage_2__7512_, data_stage_2__7511_, data_stage_2__7510_, data_stage_2__7509_, data_stage_2__7508_, data_stage_2__7507_, data_stage_2__7506_, data_stage_2__7505_, data_stage_2__7504_, data_stage_2__7503_, data_stage_2__7502_, data_stage_2__7501_, data_stage_2__7500_, data_stage_2__7499_, data_stage_2__7498_, data_stage_2__7497_, data_stage_2__7496_, data_stage_2__7495_, data_stage_2__7494_, data_stage_2__7493_, data_stage_2__7492_, data_stage_2__7491_, data_stage_2__7490_, data_stage_2__7489_, data_stage_2__7488_, data_stage_2__7487_, data_stage_2__7486_, data_stage_2__7485_, data_stage_2__7484_, data_stage_2__7483_, data_stage_2__7482_, data_stage_2__7481_, data_stage_2__7480_, data_stage_2__7479_, data_stage_2__7478_, data_stage_2__7477_, data_stage_2__7476_, data_stage_2__7475_, data_stage_2__7474_, data_stage_2__7473_, data_stage_2__7472_, data_stage_2__7471_, data_stage_2__7470_, data_stage_2__7469_, data_stage_2__7468_, data_stage_2__7467_, data_stage_2__7466_, data_stage_2__7465_, data_stage_2__7464_, data_stage_2__7463_, data_stage_2__7462_, data_stage_2__7461_, data_stage_2__7460_, data_stage_2__7459_, data_stage_2__7458_, data_stage_2__7457_, data_stage_2__7456_, data_stage_2__7455_, data_stage_2__7454_, data_stage_2__7453_, data_stage_2__7452_, data_stage_2__7451_, data_stage_2__7450_, data_stage_2__7449_, data_stage_2__7448_, data_stage_2__7447_, data_stage_2__7446_, data_stage_2__7445_, data_stage_2__7444_, data_stage_2__7443_, data_stage_2__7442_, data_stage_2__7441_, data_stage_2__7440_, data_stage_2__7439_, data_stage_2__7438_, data_stage_2__7437_, data_stage_2__7436_, data_stage_2__7435_, data_stage_2__7434_, data_stage_2__7433_, data_stage_2__7432_, data_stage_2__7431_, data_stage_2__7430_, data_stage_2__7429_, data_stage_2__7428_, data_stage_2__7427_, data_stage_2__7426_, data_stage_2__7425_, data_stage_2__7424_, data_stage_2__7423_, data_stage_2__7422_, data_stage_2__7421_, data_stage_2__7420_, data_stage_2__7419_, data_stage_2__7418_, data_stage_2__7417_, data_stage_2__7416_, data_stage_2__7415_, data_stage_2__7414_, data_stage_2__7413_, data_stage_2__7412_, data_stage_2__7411_, data_stage_2__7410_, data_stage_2__7409_, data_stage_2__7408_, data_stage_2__7407_, data_stage_2__7406_, data_stage_2__7405_, data_stage_2__7404_, data_stage_2__7403_, data_stage_2__7402_, data_stage_2__7401_, data_stage_2__7400_, data_stage_2__7399_, data_stage_2__7398_, data_stage_2__7397_, data_stage_2__7396_, data_stage_2__7395_, data_stage_2__7394_, data_stage_2__7393_, data_stage_2__7392_, data_stage_2__7391_, data_stage_2__7390_, data_stage_2__7389_, data_stage_2__7388_, data_stage_2__7387_, data_stage_2__7386_, data_stage_2__7385_, data_stage_2__7384_, data_stage_2__7383_, data_stage_2__7382_, data_stage_2__7381_, data_stage_2__7380_, data_stage_2__7379_, data_stage_2__7378_, data_stage_2__7377_, data_stage_2__7376_, data_stage_2__7375_, data_stage_2__7374_, data_stage_2__7373_, data_stage_2__7372_, data_stage_2__7371_, data_stage_2__7370_, data_stage_2__7369_, data_stage_2__7368_, data_stage_2__7367_, data_stage_2__7366_, data_stage_2__7365_, data_stage_2__7364_, data_stage_2__7363_, data_stage_2__7362_, data_stage_2__7361_, data_stage_2__7360_, data_stage_2__7359_, data_stage_2__7358_, data_stage_2__7357_, data_stage_2__7356_, data_stage_2__7355_, data_stage_2__7354_, data_stage_2__7353_, data_stage_2__7352_, data_stage_2__7351_, data_stage_2__7350_, data_stage_2__7349_, data_stage_2__7348_, data_stage_2__7347_, data_stage_2__7346_, data_stage_2__7345_, data_stage_2__7344_, data_stage_2__7343_, data_stage_2__7342_, data_stage_2__7341_, data_stage_2__7340_, data_stage_2__7339_, data_stage_2__7338_, data_stage_2__7337_, data_stage_2__7336_, data_stage_2__7335_, data_stage_2__7334_, data_stage_2__7333_, data_stage_2__7332_, data_stage_2__7331_, data_stage_2__7330_, data_stage_2__7329_, data_stage_2__7328_, data_stage_2__7327_, data_stage_2__7326_, data_stage_2__7325_, data_stage_2__7324_, data_stage_2__7323_, data_stage_2__7322_, data_stage_2__7321_, data_stage_2__7320_, data_stage_2__7319_, data_stage_2__7318_, data_stage_2__7317_, data_stage_2__7316_, data_stage_2__7315_, data_stage_2__7314_, data_stage_2__7313_, data_stage_2__7312_, data_stage_2__7311_, data_stage_2__7310_, data_stage_2__7309_, data_stage_2__7308_, data_stage_2__7307_, data_stage_2__7306_, data_stage_2__7305_, data_stage_2__7304_, data_stage_2__7303_, data_stage_2__7302_, data_stage_2__7301_, data_stage_2__7300_, data_stage_2__7299_, data_stage_2__7298_, data_stage_2__7297_, data_stage_2__7296_, data_stage_2__7295_, data_stage_2__7294_, data_stage_2__7293_, data_stage_2__7292_, data_stage_2__7291_, data_stage_2__7290_, data_stage_2__7289_, data_stage_2__7288_, data_stage_2__7287_, data_stage_2__7286_, data_stage_2__7285_, data_stage_2__7284_, data_stage_2__7283_, data_stage_2__7282_, data_stage_2__7281_, data_stage_2__7280_, data_stage_2__7279_, data_stage_2__7278_, data_stage_2__7277_, data_stage_2__7276_, data_stage_2__7275_, data_stage_2__7274_, data_stage_2__7273_, data_stage_2__7272_, data_stage_2__7271_, data_stage_2__7270_, data_stage_2__7269_, data_stage_2__7268_, data_stage_2__7267_, data_stage_2__7266_, data_stage_2__7265_, data_stage_2__7264_, data_stage_2__7263_, data_stage_2__7262_, data_stage_2__7261_, data_stage_2__7260_, data_stage_2__7259_, data_stage_2__7258_, data_stage_2__7257_, data_stage_2__7256_, data_stage_2__7255_, data_stage_2__7254_, data_stage_2__7253_, data_stage_2__7252_, data_stage_2__7251_, data_stage_2__7250_, data_stage_2__7249_, data_stage_2__7248_, data_stage_2__7247_, data_stage_2__7246_, data_stage_2__7245_, data_stage_2__7244_, data_stage_2__7243_, data_stage_2__7242_, data_stage_2__7241_, data_stage_2__7240_, data_stage_2__7239_, data_stage_2__7238_, data_stage_2__7237_, data_stage_2__7236_, data_stage_2__7235_, data_stage_2__7234_, data_stage_2__7233_, data_stage_2__7232_, data_stage_2__7231_, data_stage_2__7230_, data_stage_2__7229_, data_stage_2__7228_, data_stage_2__7227_, data_stage_2__7226_, data_stage_2__7225_, data_stage_2__7224_, data_stage_2__7223_, data_stage_2__7222_, data_stage_2__7221_, data_stage_2__7220_, data_stage_2__7219_, data_stage_2__7218_, data_stage_2__7217_, data_stage_2__7216_, data_stage_2__7215_, data_stage_2__7214_, data_stage_2__7213_, data_stage_2__7212_, data_stage_2__7211_, data_stage_2__7210_, data_stage_2__7209_, data_stage_2__7208_, data_stage_2__7207_, data_stage_2__7206_, data_stage_2__7205_, data_stage_2__7204_, data_stage_2__7203_, data_stage_2__7202_, data_stage_2__7201_, data_stage_2__7200_, data_stage_2__7199_, data_stage_2__7198_, data_stage_2__7197_, data_stage_2__7196_, data_stage_2__7195_, data_stage_2__7194_, data_stage_2__7193_, data_stage_2__7192_, data_stage_2__7191_, data_stage_2__7190_, data_stage_2__7189_, data_stage_2__7188_, data_stage_2__7187_, data_stage_2__7186_, data_stage_2__7185_, data_stage_2__7184_, data_stage_2__7183_, data_stage_2__7182_, data_stage_2__7181_, data_stage_2__7180_, data_stage_2__7179_, data_stage_2__7178_, data_stage_2__7177_, data_stage_2__7176_, data_stage_2__7175_, data_stage_2__7174_, data_stage_2__7173_, data_stage_2__7172_, data_stage_2__7171_, data_stage_2__7170_, data_stage_2__7169_, data_stage_2__7168_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__8191_, data_stage_3__8190_, data_stage_3__8189_, data_stage_3__8188_, data_stage_3__8187_, data_stage_3__8186_, data_stage_3__8185_, data_stage_3__8184_, data_stage_3__8183_, data_stage_3__8182_, data_stage_3__8181_, data_stage_3__8180_, data_stage_3__8179_, data_stage_3__8178_, data_stage_3__8177_, data_stage_3__8176_, data_stage_3__8175_, data_stage_3__8174_, data_stage_3__8173_, data_stage_3__8172_, data_stage_3__8171_, data_stage_3__8170_, data_stage_3__8169_, data_stage_3__8168_, data_stage_3__8167_, data_stage_3__8166_, data_stage_3__8165_, data_stage_3__8164_, data_stage_3__8163_, data_stage_3__8162_, data_stage_3__8161_, data_stage_3__8160_, data_stage_3__8159_, data_stage_3__8158_, data_stage_3__8157_, data_stage_3__8156_, data_stage_3__8155_, data_stage_3__8154_, data_stage_3__8153_, data_stage_3__8152_, data_stage_3__8151_, data_stage_3__8150_, data_stage_3__8149_, data_stage_3__8148_, data_stage_3__8147_, data_stage_3__8146_, data_stage_3__8145_, data_stage_3__8144_, data_stage_3__8143_, data_stage_3__8142_, data_stage_3__8141_, data_stage_3__8140_, data_stage_3__8139_, data_stage_3__8138_, data_stage_3__8137_, data_stage_3__8136_, data_stage_3__8135_, data_stage_3__8134_, data_stage_3__8133_, data_stage_3__8132_, data_stage_3__8131_, data_stage_3__8130_, data_stage_3__8129_, data_stage_3__8128_, data_stage_3__8127_, data_stage_3__8126_, data_stage_3__8125_, data_stage_3__8124_, data_stage_3__8123_, data_stage_3__8122_, data_stage_3__8121_, data_stage_3__8120_, data_stage_3__8119_, data_stage_3__8118_, data_stage_3__8117_, data_stage_3__8116_, data_stage_3__8115_, data_stage_3__8114_, data_stage_3__8113_, data_stage_3__8112_, data_stage_3__8111_, data_stage_3__8110_, data_stage_3__8109_, data_stage_3__8108_, data_stage_3__8107_, data_stage_3__8106_, data_stage_3__8105_, data_stage_3__8104_, data_stage_3__8103_, data_stage_3__8102_, data_stage_3__8101_, data_stage_3__8100_, data_stage_3__8099_, data_stage_3__8098_, data_stage_3__8097_, data_stage_3__8096_, data_stage_3__8095_, data_stage_3__8094_, data_stage_3__8093_, data_stage_3__8092_, data_stage_3__8091_, data_stage_3__8090_, data_stage_3__8089_, data_stage_3__8088_, data_stage_3__8087_, data_stage_3__8086_, data_stage_3__8085_, data_stage_3__8084_, data_stage_3__8083_, data_stage_3__8082_, data_stage_3__8081_, data_stage_3__8080_, data_stage_3__8079_, data_stage_3__8078_, data_stage_3__8077_, data_stage_3__8076_, data_stage_3__8075_, data_stage_3__8074_, data_stage_3__8073_, data_stage_3__8072_, data_stage_3__8071_, data_stage_3__8070_, data_stage_3__8069_, data_stage_3__8068_, data_stage_3__8067_, data_stage_3__8066_, data_stage_3__8065_, data_stage_3__8064_, data_stage_3__8063_, data_stage_3__8062_, data_stage_3__8061_, data_stage_3__8060_, data_stage_3__8059_, data_stage_3__8058_, data_stage_3__8057_, data_stage_3__8056_, data_stage_3__8055_, data_stage_3__8054_, data_stage_3__8053_, data_stage_3__8052_, data_stage_3__8051_, data_stage_3__8050_, data_stage_3__8049_, data_stage_3__8048_, data_stage_3__8047_, data_stage_3__8046_, data_stage_3__8045_, data_stage_3__8044_, data_stage_3__8043_, data_stage_3__8042_, data_stage_3__8041_, data_stage_3__8040_, data_stage_3__8039_, data_stage_3__8038_, data_stage_3__8037_, data_stage_3__8036_, data_stage_3__8035_, data_stage_3__8034_, data_stage_3__8033_, data_stage_3__8032_, data_stage_3__8031_, data_stage_3__8030_, data_stage_3__8029_, data_stage_3__8028_, data_stage_3__8027_, data_stage_3__8026_, data_stage_3__8025_, data_stage_3__8024_, data_stage_3__8023_, data_stage_3__8022_, data_stage_3__8021_, data_stage_3__8020_, data_stage_3__8019_, data_stage_3__8018_, data_stage_3__8017_, data_stage_3__8016_, data_stage_3__8015_, data_stage_3__8014_, data_stage_3__8013_, data_stage_3__8012_, data_stage_3__8011_, data_stage_3__8010_, data_stage_3__8009_, data_stage_3__8008_, data_stage_3__8007_, data_stage_3__8006_, data_stage_3__8005_, data_stage_3__8004_, data_stage_3__8003_, data_stage_3__8002_, data_stage_3__8001_, data_stage_3__8000_, data_stage_3__7999_, data_stage_3__7998_, data_stage_3__7997_, data_stage_3__7996_, data_stage_3__7995_, data_stage_3__7994_, data_stage_3__7993_, data_stage_3__7992_, data_stage_3__7991_, data_stage_3__7990_, data_stage_3__7989_, data_stage_3__7988_, data_stage_3__7987_, data_stage_3__7986_, data_stage_3__7985_, data_stage_3__7984_, data_stage_3__7983_, data_stage_3__7982_, data_stage_3__7981_, data_stage_3__7980_, data_stage_3__7979_, data_stage_3__7978_, data_stage_3__7977_, data_stage_3__7976_, data_stage_3__7975_, data_stage_3__7974_, data_stage_3__7973_, data_stage_3__7972_, data_stage_3__7971_, data_stage_3__7970_, data_stage_3__7969_, data_stage_3__7968_, data_stage_3__7967_, data_stage_3__7966_, data_stage_3__7965_, data_stage_3__7964_, data_stage_3__7963_, data_stage_3__7962_, data_stage_3__7961_, data_stage_3__7960_, data_stage_3__7959_, data_stage_3__7958_, data_stage_3__7957_, data_stage_3__7956_, data_stage_3__7955_, data_stage_3__7954_, data_stage_3__7953_, data_stage_3__7952_, data_stage_3__7951_, data_stage_3__7950_, data_stage_3__7949_, data_stage_3__7948_, data_stage_3__7947_, data_stage_3__7946_, data_stage_3__7945_, data_stage_3__7944_, data_stage_3__7943_, data_stage_3__7942_, data_stage_3__7941_, data_stage_3__7940_, data_stage_3__7939_, data_stage_3__7938_, data_stage_3__7937_, data_stage_3__7936_, data_stage_3__7935_, data_stage_3__7934_, data_stage_3__7933_, data_stage_3__7932_, data_stage_3__7931_, data_stage_3__7930_, data_stage_3__7929_, data_stage_3__7928_, data_stage_3__7927_, data_stage_3__7926_, data_stage_3__7925_, data_stage_3__7924_, data_stage_3__7923_, data_stage_3__7922_, data_stage_3__7921_, data_stage_3__7920_, data_stage_3__7919_, data_stage_3__7918_, data_stage_3__7917_, data_stage_3__7916_, data_stage_3__7915_, data_stage_3__7914_, data_stage_3__7913_, data_stage_3__7912_, data_stage_3__7911_, data_stage_3__7910_, data_stage_3__7909_, data_stage_3__7908_, data_stage_3__7907_, data_stage_3__7906_, data_stage_3__7905_, data_stage_3__7904_, data_stage_3__7903_, data_stage_3__7902_, data_stage_3__7901_, data_stage_3__7900_, data_stage_3__7899_, data_stage_3__7898_, data_stage_3__7897_, data_stage_3__7896_, data_stage_3__7895_, data_stage_3__7894_, data_stage_3__7893_, data_stage_3__7892_, data_stage_3__7891_, data_stage_3__7890_, data_stage_3__7889_, data_stage_3__7888_, data_stage_3__7887_, data_stage_3__7886_, data_stage_3__7885_, data_stage_3__7884_, data_stage_3__7883_, data_stage_3__7882_, data_stage_3__7881_, data_stage_3__7880_, data_stage_3__7879_, data_stage_3__7878_, data_stage_3__7877_, data_stage_3__7876_, data_stage_3__7875_, data_stage_3__7874_, data_stage_3__7873_, data_stage_3__7872_, data_stage_3__7871_, data_stage_3__7870_, data_stage_3__7869_, data_stage_3__7868_, data_stage_3__7867_, data_stage_3__7866_, data_stage_3__7865_, data_stage_3__7864_, data_stage_3__7863_, data_stage_3__7862_, data_stage_3__7861_, data_stage_3__7860_, data_stage_3__7859_, data_stage_3__7858_, data_stage_3__7857_, data_stage_3__7856_, data_stage_3__7855_, data_stage_3__7854_, data_stage_3__7853_, data_stage_3__7852_, data_stage_3__7851_, data_stage_3__7850_, data_stage_3__7849_, data_stage_3__7848_, data_stage_3__7847_, data_stage_3__7846_, data_stage_3__7845_, data_stage_3__7844_, data_stage_3__7843_, data_stage_3__7842_, data_stage_3__7841_, data_stage_3__7840_, data_stage_3__7839_, data_stage_3__7838_, data_stage_3__7837_, data_stage_3__7836_, data_stage_3__7835_, data_stage_3__7834_, data_stage_3__7833_, data_stage_3__7832_, data_stage_3__7831_, data_stage_3__7830_, data_stage_3__7829_, data_stage_3__7828_, data_stage_3__7827_, data_stage_3__7826_, data_stage_3__7825_, data_stage_3__7824_, data_stage_3__7823_, data_stage_3__7822_, data_stage_3__7821_, data_stage_3__7820_, data_stage_3__7819_, data_stage_3__7818_, data_stage_3__7817_, data_stage_3__7816_, data_stage_3__7815_, data_stage_3__7814_, data_stage_3__7813_, data_stage_3__7812_, data_stage_3__7811_, data_stage_3__7810_, data_stage_3__7809_, data_stage_3__7808_, data_stage_3__7807_, data_stage_3__7806_, data_stage_3__7805_, data_stage_3__7804_, data_stage_3__7803_, data_stage_3__7802_, data_stage_3__7801_, data_stage_3__7800_, data_stage_3__7799_, data_stage_3__7798_, data_stage_3__7797_, data_stage_3__7796_, data_stage_3__7795_, data_stage_3__7794_, data_stage_3__7793_, data_stage_3__7792_, data_stage_3__7791_, data_stage_3__7790_, data_stage_3__7789_, data_stage_3__7788_, data_stage_3__7787_, data_stage_3__7786_, data_stage_3__7785_, data_stage_3__7784_, data_stage_3__7783_, data_stage_3__7782_, data_stage_3__7781_, data_stage_3__7780_, data_stage_3__7779_, data_stage_3__7778_, data_stage_3__7777_, data_stage_3__7776_, data_stage_3__7775_, data_stage_3__7774_, data_stage_3__7773_, data_stage_3__7772_, data_stage_3__7771_, data_stage_3__7770_, data_stage_3__7769_, data_stage_3__7768_, data_stage_3__7767_, data_stage_3__7766_, data_stage_3__7765_, data_stage_3__7764_, data_stage_3__7763_, data_stage_3__7762_, data_stage_3__7761_, data_stage_3__7760_, data_stage_3__7759_, data_stage_3__7758_, data_stage_3__7757_, data_stage_3__7756_, data_stage_3__7755_, data_stage_3__7754_, data_stage_3__7753_, data_stage_3__7752_, data_stage_3__7751_, data_stage_3__7750_, data_stage_3__7749_, data_stage_3__7748_, data_stage_3__7747_, data_stage_3__7746_, data_stage_3__7745_, data_stage_3__7744_, data_stage_3__7743_, data_stage_3__7742_, data_stage_3__7741_, data_stage_3__7740_, data_stage_3__7739_, data_stage_3__7738_, data_stage_3__7737_, data_stage_3__7736_, data_stage_3__7735_, data_stage_3__7734_, data_stage_3__7733_, data_stage_3__7732_, data_stage_3__7731_, data_stage_3__7730_, data_stage_3__7729_, data_stage_3__7728_, data_stage_3__7727_, data_stage_3__7726_, data_stage_3__7725_, data_stage_3__7724_, data_stage_3__7723_, data_stage_3__7722_, data_stage_3__7721_, data_stage_3__7720_, data_stage_3__7719_, data_stage_3__7718_, data_stage_3__7717_, data_stage_3__7716_, data_stage_3__7715_, data_stage_3__7714_, data_stage_3__7713_, data_stage_3__7712_, data_stage_3__7711_, data_stage_3__7710_, data_stage_3__7709_, data_stage_3__7708_, data_stage_3__7707_, data_stage_3__7706_, data_stage_3__7705_, data_stage_3__7704_, data_stage_3__7703_, data_stage_3__7702_, data_stage_3__7701_, data_stage_3__7700_, data_stage_3__7699_, data_stage_3__7698_, data_stage_3__7697_, data_stage_3__7696_, data_stage_3__7695_, data_stage_3__7694_, data_stage_3__7693_, data_stage_3__7692_, data_stage_3__7691_, data_stage_3__7690_, data_stage_3__7689_, data_stage_3__7688_, data_stage_3__7687_, data_stage_3__7686_, data_stage_3__7685_, data_stage_3__7684_, data_stage_3__7683_, data_stage_3__7682_, data_stage_3__7681_, data_stage_3__7680_, data_stage_3__7679_, data_stage_3__7678_, data_stage_3__7677_, data_stage_3__7676_, data_stage_3__7675_, data_stage_3__7674_, data_stage_3__7673_, data_stage_3__7672_, data_stage_3__7671_, data_stage_3__7670_, data_stage_3__7669_, data_stage_3__7668_, data_stage_3__7667_, data_stage_3__7666_, data_stage_3__7665_, data_stage_3__7664_, data_stage_3__7663_, data_stage_3__7662_, data_stage_3__7661_, data_stage_3__7660_, data_stage_3__7659_, data_stage_3__7658_, data_stage_3__7657_, data_stage_3__7656_, data_stage_3__7655_, data_stage_3__7654_, data_stage_3__7653_, data_stage_3__7652_, data_stage_3__7651_, data_stage_3__7650_, data_stage_3__7649_, data_stage_3__7648_, data_stage_3__7647_, data_stage_3__7646_, data_stage_3__7645_, data_stage_3__7644_, data_stage_3__7643_, data_stage_3__7642_, data_stage_3__7641_, data_stage_3__7640_, data_stage_3__7639_, data_stage_3__7638_, data_stage_3__7637_, data_stage_3__7636_, data_stage_3__7635_, data_stage_3__7634_, data_stage_3__7633_, data_stage_3__7632_, data_stage_3__7631_, data_stage_3__7630_, data_stage_3__7629_, data_stage_3__7628_, data_stage_3__7627_, data_stage_3__7626_, data_stage_3__7625_, data_stage_3__7624_, data_stage_3__7623_, data_stage_3__7622_, data_stage_3__7621_, data_stage_3__7620_, data_stage_3__7619_, data_stage_3__7618_, data_stage_3__7617_, data_stage_3__7616_, data_stage_3__7615_, data_stage_3__7614_, data_stage_3__7613_, data_stage_3__7612_, data_stage_3__7611_, data_stage_3__7610_, data_stage_3__7609_, data_stage_3__7608_, data_stage_3__7607_, data_stage_3__7606_, data_stage_3__7605_, data_stage_3__7604_, data_stage_3__7603_, data_stage_3__7602_, data_stage_3__7601_, data_stage_3__7600_, data_stage_3__7599_, data_stage_3__7598_, data_stage_3__7597_, data_stage_3__7596_, data_stage_3__7595_, data_stage_3__7594_, data_stage_3__7593_, data_stage_3__7592_, data_stage_3__7591_, data_stage_3__7590_, data_stage_3__7589_, data_stage_3__7588_, data_stage_3__7587_, data_stage_3__7586_, data_stage_3__7585_, data_stage_3__7584_, data_stage_3__7583_, data_stage_3__7582_, data_stage_3__7581_, data_stage_3__7580_, data_stage_3__7579_, data_stage_3__7578_, data_stage_3__7577_, data_stage_3__7576_, data_stage_3__7575_, data_stage_3__7574_, data_stage_3__7573_, data_stage_3__7572_, data_stage_3__7571_, data_stage_3__7570_, data_stage_3__7569_, data_stage_3__7568_, data_stage_3__7567_, data_stage_3__7566_, data_stage_3__7565_, data_stage_3__7564_, data_stage_3__7563_, data_stage_3__7562_, data_stage_3__7561_, data_stage_3__7560_, data_stage_3__7559_, data_stage_3__7558_, data_stage_3__7557_, data_stage_3__7556_, data_stage_3__7555_, data_stage_3__7554_, data_stage_3__7553_, data_stage_3__7552_, data_stage_3__7551_, data_stage_3__7550_, data_stage_3__7549_, data_stage_3__7548_, data_stage_3__7547_, data_stage_3__7546_, data_stage_3__7545_, data_stage_3__7544_, data_stage_3__7543_, data_stage_3__7542_, data_stage_3__7541_, data_stage_3__7540_, data_stage_3__7539_, data_stage_3__7538_, data_stage_3__7537_, data_stage_3__7536_, data_stage_3__7535_, data_stage_3__7534_, data_stage_3__7533_, data_stage_3__7532_, data_stage_3__7531_, data_stage_3__7530_, data_stage_3__7529_, data_stage_3__7528_, data_stage_3__7527_, data_stage_3__7526_, data_stage_3__7525_, data_stage_3__7524_, data_stage_3__7523_, data_stage_3__7522_, data_stage_3__7521_, data_stage_3__7520_, data_stage_3__7519_, data_stage_3__7518_, data_stage_3__7517_, data_stage_3__7516_, data_stage_3__7515_, data_stage_3__7514_, data_stage_3__7513_, data_stage_3__7512_, data_stage_3__7511_, data_stage_3__7510_, data_stage_3__7509_, data_stage_3__7508_, data_stage_3__7507_, data_stage_3__7506_, data_stage_3__7505_, data_stage_3__7504_, data_stage_3__7503_, data_stage_3__7502_, data_stage_3__7501_, data_stage_3__7500_, data_stage_3__7499_, data_stage_3__7498_, data_stage_3__7497_, data_stage_3__7496_, data_stage_3__7495_, data_stage_3__7494_, data_stage_3__7493_, data_stage_3__7492_, data_stage_3__7491_, data_stage_3__7490_, data_stage_3__7489_, data_stage_3__7488_, data_stage_3__7487_, data_stage_3__7486_, data_stage_3__7485_, data_stage_3__7484_, data_stage_3__7483_, data_stage_3__7482_, data_stage_3__7481_, data_stage_3__7480_, data_stage_3__7479_, data_stage_3__7478_, data_stage_3__7477_, data_stage_3__7476_, data_stage_3__7475_, data_stage_3__7474_, data_stage_3__7473_, data_stage_3__7472_, data_stage_3__7471_, data_stage_3__7470_, data_stage_3__7469_, data_stage_3__7468_, data_stage_3__7467_, data_stage_3__7466_, data_stage_3__7465_, data_stage_3__7464_, data_stage_3__7463_, data_stage_3__7462_, data_stage_3__7461_, data_stage_3__7460_, data_stage_3__7459_, data_stage_3__7458_, data_stage_3__7457_, data_stage_3__7456_, data_stage_3__7455_, data_stage_3__7454_, data_stage_3__7453_, data_stage_3__7452_, data_stage_3__7451_, data_stage_3__7450_, data_stage_3__7449_, data_stage_3__7448_, data_stage_3__7447_, data_stage_3__7446_, data_stage_3__7445_, data_stage_3__7444_, data_stage_3__7443_, data_stage_3__7442_, data_stage_3__7441_, data_stage_3__7440_, data_stage_3__7439_, data_stage_3__7438_, data_stage_3__7437_, data_stage_3__7436_, data_stage_3__7435_, data_stage_3__7434_, data_stage_3__7433_, data_stage_3__7432_, data_stage_3__7431_, data_stage_3__7430_, data_stage_3__7429_, data_stage_3__7428_, data_stage_3__7427_, data_stage_3__7426_, data_stage_3__7425_, data_stage_3__7424_, data_stage_3__7423_, data_stage_3__7422_, data_stage_3__7421_, data_stage_3__7420_, data_stage_3__7419_, data_stage_3__7418_, data_stage_3__7417_, data_stage_3__7416_, data_stage_3__7415_, data_stage_3__7414_, data_stage_3__7413_, data_stage_3__7412_, data_stage_3__7411_, data_stage_3__7410_, data_stage_3__7409_, data_stage_3__7408_, data_stage_3__7407_, data_stage_3__7406_, data_stage_3__7405_, data_stage_3__7404_, data_stage_3__7403_, data_stage_3__7402_, data_stage_3__7401_, data_stage_3__7400_, data_stage_3__7399_, data_stage_3__7398_, data_stage_3__7397_, data_stage_3__7396_, data_stage_3__7395_, data_stage_3__7394_, data_stage_3__7393_, data_stage_3__7392_, data_stage_3__7391_, data_stage_3__7390_, data_stage_3__7389_, data_stage_3__7388_, data_stage_3__7387_, data_stage_3__7386_, data_stage_3__7385_, data_stage_3__7384_, data_stage_3__7383_, data_stage_3__7382_, data_stage_3__7381_, data_stage_3__7380_, data_stage_3__7379_, data_stage_3__7378_, data_stage_3__7377_, data_stage_3__7376_, data_stage_3__7375_, data_stage_3__7374_, data_stage_3__7373_, data_stage_3__7372_, data_stage_3__7371_, data_stage_3__7370_, data_stage_3__7369_, data_stage_3__7368_, data_stage_3__7367_, data_stage_3__7366_, data_stage_3__7365_, data_stage_3__7364_, data_stage_3__7363_, data_stage_3__7362_, data_stage_3__7361_, data_stage_3__7360_, data_stage_3__7359_, data_stage_3__7358_, data_stage_3__7357_, data_stage_3__7356_, data_stage_3__7355_, data_stage_3__7354_, data_stage_3__7353_, data_stage_3__7352_, data_stage_3__7351_, data_stage_3__7350_, data_stage_3__7349_, data_stage_3__7348_, data_stage_3__7347_, data_stage_3__7346_, data_stage_3__7345_, data_stage_3__7344_, data_stage_3__7343_, data_stage_3__7342_, data_stage_3__7341_, data_stage_3__7340_, data_stage_3__7339_, data_stage_3__7338_, data_stage_3__7337_, data_stage_3__7336_, data_stage_3__7335_, data_stage_3__7334_, data_stage_3__7333_, data_stage_3__7332_, data_stage_3__7331_, data_stage_3__7330_, data_stage_3__7329_, data_stage_3__7328_, data_stage_3__7327_, data_stage_3__7326_, data_stage_3__7325_, data_stage_3__7324_, data_stage_3__7323_, data_stage_3__7322_, data_stage_3__7321_, data_stage_3__7320_, data_stage_3__7319_, data_stage_3__7318_, data_stage_3__7317_, data_stage_3__7316_, data_stage_3__7315_, data_stage_3__7314_, data_stage_3__7313_, data_stage_3__7312_, data_stage_3__7311_, data_stage_3__7310_, data_stage_3__7309_, data_stage_3__7308_, data_stage_3__7307_, data_stage_3__7306_, data_stage_3__7305_, data_stage_3__7304_, data_stage_3__7303_, data_stage_3__7302_, data_stage_3__7301_, data_stage_3__7300_, data_stage_3__7299_, data_stage_3__7298_, data_stage_3__7297_, data_stage_3__7296_, data_stage_3__7295_, data_stage_3__7294_, data_stage_3__7293_, data_stage_3__7292_, data_stage_3__7291_, data_stage_3__7290_, data_stage_3__7289_, data_stage_3__7288_, data_stage_3__7287_, data_stage_3__7286_, data_stage_3__7285_, data_stage_3__7284_, data_stage_3__7283_, data_stage_3__7282_, data_stage_3__7281_, data_stage_3__7280_, data_stage_3__7279_, data_stage_3__7278_, data_stage_3__7277_, data_stage_3__7276_, data_stage_3__7275_, data_stage_3__7274_, data_stage_3__7273_, data_stage_3__7272_, data_stage_3__7271_, data_stage_3__7270_, data_stage_3__7269_, data_stage_3__7268_, data_stage_3__7267_, data_stage_3__7266_, data_stage_3__7265_, data_stage_3__7264_, data_stage_3__7263_, data_stage_3__7262_, data_stage_3__7261_, data_stage_3__7260_, data_stage_3__7259_, data_stage_3__7258_, data_stage_3__7257_, data_stage_3__7256_, data_stage_3__7255_, data_stage_3__7254_, data_stage_3__7253_, data_stage_3__7252_, data_stage_3__7251_, data_stage_3__7250_, data_stage_3__7249_, data_stage_3__7248_, data_stage_3__7247_, data_stage_3__7246_, data_stage_3__7245_, data_stage_3__7244_, data_stage_3__7243_, data_stage_3__7242_, data_stage_3__7241_, data_stage_3__7240_, data_stage_3__7239_, data_stage_3__7238_, data_stage_3__7237_, data_stage_3__7236_, data_stage_3__7235_, data_stage_3__7234_, data_stage_3__7233_, data_stage_3__7232_, data_stage_3__7231_, data_stage_3__7230_, data_stage_3__7229_, data_stage_3__7228_, data_stage_3__7227_, data_stage_3__7226_, data_stage_3__7225_, data_stage_3__7224_, data_stage_3__7223_, data_stage_3__7222_, data_stage_3__7221_, data_stage_3__7220_, data_stage_3__7219_, data_stage_3__7218_, data_stage_3__7217_, data_stage_3__7216_, data_stage_3__7215_, data_stage_3__7214_, data_stage_3__7213_, data_stage_3__7212_, data_stage_3__7211_, data_stage_3__7210_, data_stage_3__7209_, data_stage_3__7208_, data_stage_3__7207_, data_stage_3__7206_, data_stage_3__7205_, data_stage_3__7204_, data_stage_3__7203_, data_stage_3__7202_, data_stage_3__7201_, data_stage_3__7200_, data_stage_3__7199_, data_stage_3__7198_, data_stage_3__7197_, data_stage_3__7196_, data_stage_3__7195_, data_stage_3__7194_, data_stage_3__7193_, data_stage_3__7192_, data_stage_3__7191_, data_stage_3__7190_, data_stage_3__7189_, data_stage_3__7188_, data_stage_3__7187_, data_stage_3__7186_, data_stage_3__7185_, data_stage_3__7184_, data_stage_3__7183_, data_stage_3__7182_, data_stage_3__7181_, data_stage_3__7180_, data_stage_3__7179_, data_stage_3__7178_, data_stage_3__7177_, data_stage_3__7176_, data_stage_3__7175_, data_stage_3__7174_, data_stage_3__7173_, data_stage_3__7172_, data_stage_3__7171_, data_stage_3__7170_, data_stage_3__7169_, data_stage_3__7168_ })
  );


  bsg_swap_width_p1024
  mux_stage_3__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_3__2047_, data_stage_3__2046_, data_stage_3__2045_, data_stage_3__2044_, data_stage_3__2043_, data_stage_3__2042_, data_stage_3__2041_, data_stage_3__2040_, data_stage_3__2039_, data_stage_3__2038_, data_stage_3__2037_, data_stage_3__2036_, data_stage_3__2035_, data_stage_3__2034_, data_stage_3__2033_, data_stage_3__2032_, data_stage_3__2031_, data_stage_3__2030_, data_stage_3__2029_, data_stage_3__2028_, data_stage_3__2027_, data_stage_3__2026_, data_stage_3__2025_, data_stage_3__2024_, data_stage_3__2023_, data_stage_3__2022_, data_stage_3__2021_, data_stage_3__2020_, data_stage_3__2019_, data_stage_3__2018_, data_stage_3__2017_, data_stage_3__2016_, data_stage_3__2015_, data_stage_3__2014_, data_stage_3__2013_, data_stage_3__2012_, data_stage_3__2011_, data_stage_3__2010_, data_stage_3__2009_, data_stage_3__2008_, data_stage_3__2007_, data_stage_3__2006_, data_stage_3__2005_, data_stage_3__2004_, data_stage_3__2003_, data_stage_3__2002_, data_stage_3__2001_, data_stage_3__2000_, data_stage_3__1999_, data_stage_3__1998_, data_stage_3__1997_, data_stage_3__1996_, data_stage_3__1995_, data_stage_3__1994_, data_stage_3__1993_, data_stage_3__1992_, data_stage_3__1991_, data_stage_3__1990_, data_stage_3__1989_, data_stage_3__1988_, data_stage_3__1987_, data_stage_3__1986_, data_stage_3__1985_, data_stage_3__1984_, data_stage_3__1983_, data_stage_3__1982_, data_stage_3__1981_, data_stage_3__1980_, data_stage_3__1979_, data_stage_3__1978_, data_stage_3__1977_, data_stage_3__1976_, data_stage_3__1975_, data_stage_3__1974_, data_stage_3__1973_, data_stage_3__1972_, data_stage_3__1971_, data_stage_3__1970_, data_stage_3__1969_, data_stage_3__1968_, data_stage_3__1967_, data_stage_3__1966_, data_stage_3__1965_, data_stage_3__1964_, data_stage_3__1963_, data_stage_3__1962_, data_stage_3__1961_, data_stage_3__1960_, data_stage_3__1959_, data_stage_3__1958_, data_stage_3__1957_, data_stage_3__1956_, data_stage_3__1955_, data_stage_3__1954_, data_stage_3__1953_, data_stage_3__1952_, data_stage_3__1951_, data_stage_3__1950_, data_stage_3__1949_, data_stage_3__1948_, data_stage_3__1947_, data_stage_3__1946_, data_stage_3__1945_, data_stage_3__1944_, data_stage_3__1943_, data_stage_3__1942_, data_stage_3__1941_, data_stage_3__1940_, data_stage_3__1939_, data_stage_3__1938_, data_stage_3__1937_, data_stage_3__1936_, data_stage_3__1935_, data_stage_3__1934_, data_stage_3__1933_, data_stage_3__1932_, data_stage_3__1931_, data_stage_3__1930_, data_stage_3__1929_, data_stage_3__1928_, data_stage_3__1927_, data_stage_3__1926_, data_stage_3__1925_, data_stage_3__1924_, data_stage_3__1923_, data_stage_3__1922_, data_stage_3__1921_, data_stage_3__1920_, data_stage_3__1919_, data_stage_3__1918_, data_stage_3__1917_, data_stage_3__1916_, data_stage_3__1915_, data_stage_3__1914_, data_stage_3__1913_, data_stage_3__1912_, data_stage_3__1911_, data_stage_3__1910_, data_stage_3__1909_, data_stage_3__1908_, data_stage_3__1907_, data_stage_3__1906_, data_stage_3__1905_, data_stage_3__1904_, data_stage_3__1903_, data_stage_3__1902_, data_stage_3__1901_, data_stage_3__1900_, data_stage_3__1899_, data_stage_3__1898_, data_stage_3__1897_, data_stage_3__1896_, data_stage_3__1895_, data_stage_3__1894_, data_stage_3__1893_, data_stage_3__1892_, data_stage_3__1891_, data_stage_3__1890_, data_stage_3__1889_, data_stage_3__1888_, data_stage_3__1887_, data_stage_3__1886_, data_stage_3__1885_, data_stage_3__1884_, data_stage_3__1883_, data_stage_3__1882_, data_stage_3__1881_, data_stage_3__1880_, data_stage_3__1879_, data_stage_3__1878_, data_stage_3__1877_, data_stage_3__1876_, data_stage_3__1875_, data_stage_3__1874_, data_stage_3__1873_, data_stage_3__1872_, data_stage_3__1871_, data_stage_3__1870_, data_stage_3__1869_, data_stage_3__1868_, data_stage_3__1867_, data_stage_3__1866_, data_stage_3__1865_, data_stage_3__1864_, data_stage_3__1863_, data_stage_3__1862_, data_stage_3__1861_, data_stage_3__1860_, data_stage_3__1859_, data_stage_3__1858_, data_stage_3__1857_, data_stage_3__1856_, data_stage_3__1855_, data_stage_3__1854_, data_stage_3__1853_, data_stage_3__1852_, data_stage_3__1851_, data_stage_3__1850_, data_stage_3__1849_, data_stage_3__1848_, data_stage_3__1847_, data_stage_3__1846_, data_stage_3__1845_, data_stage_3__1844_, data_stage_3__1843_, data_stage_3__1842_, data_stage_3__1841_, data_stage_3__1840_, data_stage_3__1839_, data_stage_3__1838_, data_stage_3__1837_, data_stage_3__1836_, data_stage_3__1835_, data_stage_3__1834_, data_stage_3__1833_, data_stage_3__1832_, data_stage_3__1831_, data_stage_3__1830_, data_stage_3__1829_, data_stage_3__1828_, data_stage_3__1827_, data_stage_3__1826_, data_stage_3__1825_, data_stage_3__1824_, data_stage_3__1823_, data_stage_3__1822_, data_stage_3__1821_, data_stage_3__1820_, data_stage_3__1819_, data_stage_3__1818_, data_stage_3__1817_, data_stage_3__1816_, data_stage_3__1815_, data_stage_3__1814_, data_stage_3__1813_, data_stage_3__1812_, data_stage_3__1811_, data_stage_3__1810_, data_stage_3__1809_, data_stage_3__1808_, data_stage_3__1807_, data_stage_3__1806_, data_stage_3__1805_, data_stage_3__1804_, data_stage_3__1803_, data_stage_3__1802_, data_stage_3__1801_, data_stage_3__1800_, data_stage_3__1799_, data_stage_3__1798_, data_stage_3__1797_, data_stage_3__1796_, data_stage_3__1795_, data_stage_3__1794_, data_stage_3__1793_, data_stage_3__1792_, data_stage_3__1791_, data_stage_3__1790_, data_stage_3__1789_, data_stage_3__1788_, data_stage_3__1787_, data_stage_3__1786_, data_stage_3__1785_, data_stage_3__1784_, data_stage_3__1783_, data_stage_3__1782_, data_stage_3__1781_, data_stage_3__1780_, data_stage_3__1779_, data_stage_3__1778_, data_stage_3__1777_, data_stage_3__1776_, data_stage_3__1775_, data_stage_3__1774_, data_stage_3__1773_, data_stage_3__1772_, data_stage_3__1771_, data_stage_3__1770_, data_stage_3__1769_, data_stage_3__1768_, data_stage_3__1767_, data_stage_3__1766_, data_stage_3__1765_, data_stage_3__1764_, data_stage_3__1763_, data_stage_3__1762_, data_stage_3__1761_, data_stage_3__1760_, data_stage_3__1759_, data_stage_3__1758_, data_stage_3__1757_, data_stage_3__1756_, data_stage_3__1755_, data_stage_3__1754_, data_stage_3__1753_, data_stage_3__1752_, data_stage_3__1751_, data_stage_3__1750_, data_stage_3__1749_, data_stage_3__1748_, data_stage_3__1747_, data_stage_3__1746_, data_stage_3__1745_, data_stage_3__1744_, data_stage_3__1743_, data_stage_3__1742_, data_stage_3__1741_, data_stage_3__1740_, data_stage_3__1739_, data_stage_3__1738_, data_stage_3__1737_, data_stage_3__1736_, data_stage_3__1735_, data_stage_3__1734_, data_stage_3__1733_, data_stage_3__1732_, data_stage_3__1731_, data_stage_3__1730_, data_stage_3__1729_, data_stage_3__1728_, data_stage_3__1727_, data_stage_3__1726_, data_stage_3__1725_, data_stage_3__1724_, data_stage_3__1723_, data_stage_3__1722_, data_stage_3__1721_, data_stage_3__1720_, data_stage_3__1719_, data_stage_3__1718_, data_stage_3__1717_, data_stage_3__1716_, data_stage_3__1715_, data_stage_3__1714_, data_stage_3__1713_, data_stage_3__1712_, data_stage_3__1711_, data_stage_3__1710_, data_stage_3__1709_, data_stage_3__1708_, data_stage_3__1707_, data_stage_3__1706_, data_stage_3__1705_, data_stage_3__1704_, data_stage_3__1703_, data_stage_3__1702_, data_stage_3__1701_, data_stage_3__1700_, data_stage_3__1699_, data_stage_3__1698_, data_stage_3__1697_, data_stage_3__1696_, data_stage_3__1695_, data_stage_3__1694_, data_stage_3__1693_, data_stage_3__1692_, data_stage_3__1691_, data_stage_3__1690_, data_stage_3__1689_, data_stage_3__1688_, data_stage_3__1687_, data_stage_3__1686_, data_stage_3__1685_, data_stage_3__1684_, data_stage_3__1683_, data_stage_3__1682_, data_stage_3__1681_, data_stage_3__1680_, data_stage_3__1679_, data_stage_3__1678_, data_stage_3__1677_, data_stage_3__1676_, data_stage_3__1675_, data_stage_3__1674_, data_stage_3__1673_, data_stage_3__1672_, data_stage_3__1671_, data_stage_3__1670_, data_stage_3__1669_, data_stage_3__1668_, data_stage_3__1667_, data_stage_3__1666_, data_stage_3__1665_, data_stage_3__1664_, data_stage_3__1663_, data_stage_3__1662_, data_stage_3__1661_, data_stage_3__1660_, data_stage_3__1659_, data_stage_3__1658_, data_stage_3__1657_, data_stage_3__1656_, data_stage_3__1655_, data_stage_3__1654_, data_stage_3__1653_, data_stage_3__1652_, data_stage_3__1651_, data_stage_3__1650_, data_stage_3__1649_, data_stage_3__1648_, data_stage_3__1647_, data_stage_3__1646_, data_stage_3__1645_, data_stage_3__1644_, data_stage_3__1643_, data_stage_3__1642_, data_stage_3__1641_, data_stage_3__1640_, data_stage_3__1639_, data_stage_3__1638_, data_stage_3__1637_, data_stage_3__1636_, data_stage_3__1635_, data_stage_3__1634_, data_stage_3__1633_, data_stage_3__1632_, data_stage_3__1631_, data_stage_3__1630_, data_stage_3__1629_, data_stage_3__1628_, data_stage_3__1627_, data_stage_3__1626_, data_stage_3__1625_, data_stage_3__1624_, data_stage_3__1623_, data_stage_3__1622_, data_stage_3__1621_, data_stage_3__1620_, data_stage_3__1619_, data_stage_3__1618_, data_stage_3__1617_, data_stage_3__1616_, data_stage_3__1615_, data_stage_3__1614_, data_stage_3__1613_, data_stage_3__1612_, data_stage_3__1611_, data_stage_3__1610_, data_stage_3__1609_, data_stage_3__1608_, data_stage_3__1607_, data_stage_3__1606_, data_stage_3__1605_, data_stage_3__1604_, data_stage_3__1603_, data_stage_3__1602_, data_stage_3__1601_, data_stage_3__1600_, data_stage_3__1599_, data_stage_3__1598_, data_stage_3__1597_, data_stage_3__1596_, data_stage_3__1595_, data_stage_3__1594_, data_stage_3__1593_, data_stage_3__1592_, data_stage_3__1591_, data_stage_3__1590_, data_stage_3__1589_, data_stage_3__1588_, data_stage_3__1587_, data_stage_3__1586_, data_stage_3__1585_, data_stage_3__1584_, data_stage_3__1583_, data_stage_3__1582_, data_stage_3__1581_, data_stage_3__1580_, data_stage_3__1579_, data_stage_3__1578_, data_stage_3__1577_, data_stage_3__1576_, data_stage_3__1575_, data_stage_3__1574_, data_stage_3__1573_, data_stage_3__1572_, data_stage_3__1571_, data_stage_3__1570_, data_stage_3__1569_, data_stage_3__1568_, data_stage_3__1567_, data_stage_3__1566_, data_stage_3__1565_, data_stage_3__1564_, data_stage_3__1563_, data_stage_3__1562_, data_stage_3__1561_, data_stage_3__1560_, data_stage_3__1559_, data_stage_3__1558_, data_stage_3__1557_, data_stage_3__1556_, data_stage_3__1555_, data_stage_3__1554_, data_stage_3__1553_, data_stage_3__1552_, data_stage_3__1551_, data_stage_3__1550_, data_stage_3__1549_, data_stage_3__1548_, data_stage_3__1547_, data_stage_3__1546_, data_stage_3__1545_, data_stage_3__1544_, data_stage_3__1543_, data_stage_3__1542_, data_stage_3__1541_, data_stage_3__1540_, data_stage_3__1539_, data_stage_3__1538_, data_stage_3__1537_, data_stage_3__1536_, data_stage_3__1535_, data_stage_3__1534_, data_stage_3__1533_, data_stage_3__1532_, data_stage_3__1531_, data_stage_3__1530_, data_stage_3__1529_, data_stage_3__1528_, data_stage_3__1527_, data_stage_3__1526_, data_stage_3__1525_, data_stage_3__1524_, data_stage_3__1523_, data_stage_3__1522_, data_stage_3__1521_, data_stage_3__1520_, data_stage_3__1519_, data_stage_3__1518_, data_stage_3__1517_, data_stage_3__1516_, data_stage_3__1515_, data_stage_3__1514_, data_stage_3__1513_, data_stage_3__1512_, data_stage_3__1511_, data_stage_3__1510_, data_stage_3__1509_, data_stage_3__1508_, data_stage_3__1507_, data_stage_3__1506_, data_stage_3__1505_, data_stage_3__1504_, data_stage_3__1503_, data_stage_3__1502_, data_stage_3__1501_, data_stage_3__1500_, data_stage_3__1499_, data_stage_3__1498_, data_stage_3__1497_, data_stage_3__1496_, data_stage_3__1495_, data_stage_3__1494_, data_stage_3__1493_, data_stage_3__1492_, data_stage_3__1491_, data_stage_3__1490_, data_stage_3__1489_, data_stage_3__1488_, data_stage_3__1487_, data_stage_3__1486_, data_stage_3__1485_, data_stage_3__1484_, data_stage_3__1483_, data_stage_3__1482_, data_stage_3__1481_, data_stage_3__1480_, data_stage_3__1479_, data_stage_3__1478_, data_stage_3__1477_, data_stage_3__1476_, data_stage_3__1475_, data_stage_3__1474_, data_stage_3__1473_, data_stage_3__1472_, data_stage_3__1471_, data_stage_3__1470_, data_stage_3__1469_, data_stage_3__1468_, data_stage_3__1467_, data_stage_3__1466_, data_stage_3__1465_, data_stage_3__1464_, data_stage_3__1463_, data_stage_3__1462_, data_stage_3__1461_, data_stage_3__1460_, data_stage_3__1459_, data_stage_3__1458_, data_stage_3__1457_, data_stage_3__1456_, data_stage_3__1455_, data_stage_3__1454_, data_stage_3__1453_, data_stage_3__1452_, data_stage_3__1451_, data_stage_3__1450_, data_stage_3__1449_, data_stage_3__1448_, data_stage_3__1447_, data_stage_3__1446_, data_stage_3__1445_, data_stage_3__1444_, data_stage_3__1443_, data_stage_3__1442_, data_stage_3__1441_, data_stage_3__1440_, data_stage_3__1439_, data_stage_3__1438_, data_stage_3__1437_, data_stage_3__1436_, data_stage_3__1435_, data_stage_3__1434_, data_stage_3__1433_, data_stage_3__1432_, data_stage_3__1431_, data_stage_3__1430_, data_stage_3__1429_, data_stage_3__1428_, data_stage_3__1427_, data_stage_3__1426_, data_stage_3__1425_, data_stage_3__1424_, data_stage_3__1423_, data_stage_3__1422_, data_stage_3__1421_, data_stage_3__1420_, data_stage_3__1419_, data_stage_3__1418_, data_stage_3__1417_, data_stage_3__1416_, data_stage_3__1415_, data_stage_3__1414_, data_stage_3__1413_, data_stage_3__1412_, data_stage_3__1411_, data_stage_3__1410_, data_stage_3__1409_, data_stage_3__1408_, data_stage_3__1407_, data_stage_3__1406_, data_stage_3__1405_, data_stage_3__1404_, data_stage_3__1403_, data_stage_3__1402_, data_stage_3__1401_, data_stage_3__1400_, data_stage_3__1399_, data_stage_3__1398_, data_stage_3__1397_, data_stage_3__1396_, data_stage_3__1395_, data_stage_3__1394_, data_stage_3__1393_, data_stage_3__1392_, data_stage_3__1391_, data_stage_3__1390_, data_stage_3__1389_, data_stage_3__1388_, data_stage_3__1387_, data_stage_3__1386_, data_stage_3__1385_, data_stage_3__1384_, data_stage_3__1383_, data_stage_3__1382_, data_stage_3__1381_, data_stage_3__1380_, data_stage_3__1379_, data_stage_3__1378_, data_stage_3__1377_, data_stage_3__1376_, data_stage_3__1375_, data_stage_3__1374_, data_stage_3__1373_, data_stage_3__1372_, data_stage_3__1371_, data_stage_3__1370_, data_stage_3__1369_, data_stage_3__1368_, data_stage_3__1367_, data_stage_3__1366_, data_stage_3__1365_, data_stage_3__1364_, data_stage_3__1363_, data_stage_3__1362_, data_stage_3__1361_, data_stage_3__1360_, data_stage_3__1359_, data_stage_3__1358_, data_stage_3__1357_, data_stage_3__1356_, data_stage_3__1355_, data_stage_3__1354_, data_stage_3__1353_, data_stage_3__1352_, data_stage_3__1351_, data_stage_3__1350_, data_stage_3__1349_, data_stage_3__1348_, data_stage_3__1347_, data_stage_3__1346_, data_stage_3__1345_, data_stage_3__1344_, data_stage_3__1343_, data_stage_3__1342_, data_stage_3__1341_, data_stage_3__1340_, data_stage_3__1339_, data_stage_3__1338_, data_stage_3__1337_, data_stage_3__1336_, data_stage_3__1335_, data_stage_3__1334_, data_stage_3__1333_, data_stage_3__1332_, data_stage_3__1331_, data_stage_3__1330_, data_stage_3__1329_, data_stage_3__1328_, data_stage_3__1327_, data_stage_3__1326_, data_stage_3__1325_, data_stage_3__1324_, data_stage_3__1323_, data_stage_3__1322_, data_stage_3__1321_, data_stage_3__1320_, data_stage_3__1319_, data_stage_3__1318_, data_stage_3__1317_, data_stage_3__1316_, data_stage_3__1315_, data_stage_3__1314_, data_stage_3__1313_, data_stage_3__1312_, data_stage_3__1311_, data_stage_3__1310_, data_stage_3__1309_, data_stage_3__1308_, data_stage_3__1307_, data_stage_3__1306_, data_stage_3__1305_, data_stage_3__1304_, data_stage_3__1303_, data_stage_3__1302_, data_stage_3__1301_, data_stage_3__1300_, data_stage_3__1299_, data_stage_3__1298_, data_stage_3__1297_, data_stage_3__1296_, data_stage_3__1295_, data_stage_3__1294_, data_stage_3__1293_, data_stage_3__1292_, data_stage_3__1291_, data_stage_3__1290_, data_stage_3__1289_, data_stage_3__1288_, data_stage_3__1287_, data_stage_3__1286_, data_stage_3__1285_, data_stage_3__1284_, data_stage_3__1283_, data_stage_3__1282_, data_stage_3__1281_, data_stage_3__1280_, data_stage_3__1279_, data_stage_3__1278_, data_stage_3__1277_, data_stage_3__1276_, data_stage_3__1275_, data_stage_3__1274_, data_stage_3__1273_, data_stage_3__1272_, data_stage_3__1271_, data_stage_3__1270_, data_stage_3__1269_, data_stage_3__1268_, data_stage_3__1267_, data_stage_3__1266_, data_stage_3__1265_, data_stage_3__1264_, data_stage_3__1263_, data_stage_3__1262_, data_stage_3__1261_, data_stage_3__1260_, data_stage_3__1259_, data_stage_3__1258_, data_stage_3__1257_, data_stage_3__1256_, data_stage_3__1255_, data_stage_3__1254_, data_stage_3__1253_, data_stage_3__1252_, data_stage_3__1251_, data_stage_3__1250_, data_stage_3__1249_, data_stage_3__1248_, data_stage_3__1247_, data_stage_3__1246_, data_stage_3__1245_, data_stage_3__1244_, data_stage_3__1243_, data_stage_3__1242_, data_stage_3__1241_, data_stage_3__1240_, data_stage_3__1239_, data_stage_3__1238_, data_stage_3__1237_, data_stage_3__1236_, data_stage_3__1235_, data_stage_3__1234_, data_stage_3__1233_, data_stage_3__1232_, data_stage_3__1231_, data_stage_3__1230_, data_stage_3__1229_, data_stage_3__1228_, data_stage_3__1227_, data_stage_3__1226_, data_stage_3__1225_, data_stage_3__1224_, data_stage_3__1223_, data_stage_3__1222_, data_stage_3__1221_, data_stage_3__1220_, data_stage_3__1219_, data_stage_3__1218_, data_stage_3__1217_, data_stage_3__1216_, data_stage_3__1215_, data_stage_3__1214_, data_stage_3__1213_, data_stage_3__1212_, data_stage_3__1211_, data_stage_3__1210_, data_stage_3__1209_, data_stage_3__1208_, data_stage_3__1207_, data_stage_3__1206_, data_stage_3__1205_, data_stage_3__1204_, data_stage_3__1203_, data_stage_3__1202_, data_stage_3__1201_, data_stage_3__1200_, data_stage_3__1199_, data_stage_3__1198_, data_stage_3__1197_, data_stage_3__1196_, data_stage_3__1195_, data_stage_3__1194_, data_stage_3__1193_, data_stage_3__1192_, data_stage_3__1191_, data_stage_3__1190_, data_stage_3__1189_, data_stage_3__1188_, data_stage_3__1187_, data_stage_3__1186_, data_stage_3__1185_, data_stage_3__1184_, data_stage_3__1183_, data_stage_3__1182_, data_stage_3__1181_, data_stage_3__1180_, data_stage_3__1179_, data_stage_3__1178_, data_stage_3__1177_, data_stage_3__1176_, data_stage_3__1175_, data_stage_3__1174_, data_stage_3__1173_, data_stage_3__1172_, data_stage_3__1171_, data_stage_3__1170_, data_stage_3__1169_, data_stage_3__1168_, data_stage_3__1167_, data_stage_3__1166_, data_stage_3__1165_, data_stage_3__1164_, data_stage_3__1163_, data_stage_3__1162_, data_stage_3__1161_, data_stage_3__1160_, data_stage_3__1159_, data_stage_3__1158_, data_stage_3__1157_, data_stage_3__1156_, data_stage_3__1155_, data_stage_3__1154_, data_stage_3__1153_, data_stage_3__1152_, data_stage_3__1151_, data_stage_3__1150_, data_stage_3__1149_, data_stage_3__1148_, data_stage_3__1147_, data_stage_3__1146_, data_stage_3__1145_, data_stage_3__1144_, data_stage_3__1143_, data_stage_3__1142_, data_stage_3__1141_, data_stage_3__1140_, data_stage_3__1139_, data_stage_3__1138_, data_stage_3__1137_, data_stage_3__1136_, data_stage_3__1135_, data_stage_3__1134_, data_stage_3__1133_, data_stage_3__1132_, data_stage_3__1131_, data_stage_3__1130_, data_stage_3__1129_, data_stage_3__1128_, data_stage_3__1127_, data_stage_3__1126_, data_stage_3__1125_, data_stage_3__1124_, data_stage_3__1123_, data_stage_3__1122_, data_stage_3__1121_, data_stage_3__1120_, data_stage_3__1119_, data_stage_3__1118_, data_stage_3__1117_, data_stage_3__1116_, data_stage_3__1115_, data_stage_3__1114_, data_stage_3__1113_, data_stage_3__1112_, data_stage_3__1111_, data_stage_3__1110_, data_stage_3__1109_, data_stage_3__1108_, data_stage_3__1107_, data_stage_3__1106_, data_stage_3__1105_, data_stage_3__1104_, data_stage_3__1103_, data_stage_3__1102_, data_stage_3__1101_, data_stage_3__1100_, data_stage_3__1099_, data_stage_3__1098_, data_stage_3__1097_, data_stage_3__1096_, data_stage_3__1095_, data_stage_3__1094_, data_stage_3__1093_, data_stage_3__1092_, data_stage_3__1091_, data_stage_3__1090_, data_stage_3__1089_, data_stage_3__1088_, data_stage_3__1087_, data_stage_3__1086_, data_stage_3__1085_, data_stage_3__1084_, data_stage_3__1083_, data_stage_3__1082_, data_stage_3__1081_, data_stage_3__1080_, data_stage_3__1079_, data_stage_3__1078_, data_stage_3__1077_, data_stage_3__1076_, data_stage_3__1075_, data_stage_3__1074_, data_stage_3__1073_, data_stage_3__1072_, data_stage_3__1071_, data_stage_3__1070_, data_stage_3__1069_, data_stage_3__1068_, data_stage_3__1067_, data_stage_3__1066_, data_stage_3__1065_, data_stage_3__1064_, data_stage_3__1063_, data_stage_3__1062_, data_stage_3__1061_, data_stage_3__1060_, data_stage_3__1059_, data_stage_3__1058_, data_stage_3__1057_, data_stage_3__1056_, data_stage_3__1055_, data_stage_3__1054_, data_stage_3__1053_, data_stage_3__1052_, data_stage_3__1051_, data_stage_3__1050_, data_stage_3__1049_, data_stage_3__1048_, data_stage_3__1047_, data_stage_3__1046_, data_stage_3__1045_, data_stage_3__1044_, data_stage_3__1043_, data_stage_3__1042_, data_stage_3__1041_, data_stage_3__1040_, data_stage_3__1039_, data_stage_3__1038_, data_stage_3__1037_, data_stage_3__1036_, data_stage_3__1035_, data_stage_3__1034_, data_stage_3__1033_, data_stage_3__1032_, data_stage_3__1031_, data_stage_3__1030_, data_stage_3__1029_, data_stage_3__1028_, data_stage_3__1027_, data_stage_3__1026_, data_stage_3__1025_, data_stage_3__1024_, data_stage_3__1023_, data_stage_3__1022_, data_stage_3__1021_, data_stage_3__1020_, data_stage_3__1019_, data_stage_3__1018_, data_stage_3__1017_, data_stage_3__1016_, data_stage_3__1015_, data_stage_3__1014_, data_stage_3__1013_, data_stage_3__1012_, data_stage_3__1011_, data_stage_3__1010_, data_stage_3__1009_, data_stage_3__1008_, data_stage_3__1007_, data_stage_3__1006_, data_stage_3__1005_, data_stage_3__1004_, data_stage_3__1003_, data_stage_3__1002_, data_stage_3__1001_, data_stage_3__1000_, data_stage_3__999_, data_stage_3__998_, data_stage_3__997_, data_stage_3__996_, data_stage_3__995_, data_stage_3__994_, data_stage_3__993_, data_stage_3__992_, data_stage_3__991_, data_stage_3__990_, data_stage_3__989_, data_stage_3__988_, data_stage_3__987_, data_stage_3__986_, data_stage_3__985_, data_stage_3__984_, data_stage_3__983_, data_stage_3__982_, data_stage_3__981_, data_stage_3__980_, data_stage_3__979_, data_stage_3__978_, data_stage_3__977_, data_stage_3__976_, data_stage_3__975_, data_stage_3__974_, data_stage_3__973_, data_stage_3__972_, data_stage_3__971_, data_stage_3__970_, data_stage_3__969_, data_stage_3__968_, data_stage_3__967_, data_stage_3__966_, data_stage_3__965_, data_stage_3__964_, data_stage_3__963_, data_stage_3__962_, data_stage_3__961_, data_stage_3__960_, data_stage_3__959_, data_stage_3__958_, data_stage_3__957_, data_stage_3__956_, data_stage_3__955_, data_stage_3__954_, data_stage_3__953_, data_stage_3__952_, data_stage_3__951_, data_stage_3__950_, data_stage_3__949_, data_stage_3__948_, data_stage_3__947_, data_stage_3__946_, data_stage_3__945_, data_stage_3__944_, data_stage_3__943_, data_stage_3__942_, data_stage_3__941_, data_stage_3__940_, data_stage_3__939_, data_stage_3__938_, data_stage_3__937_, data_stage_3__936_, data_stage_3__935_, data_stage_3__934_, data_stage_3__933_, data_stage_3__932_, data_stage_3__931_, data_stage_3__930_, data_stage_3__929_, data_stage_3__928_, data_stage_3__927_, data_stage_3__926_, data_stage_3__925_, data_stage_3__924_, data_stage_3__923_, data_stage_3__922_, data_stage_3__921_, data_stage_3__920_, data_stage_3__919_, data_stage_3__918_, data_stage_3__917_, data_stage_3__916_, data_stage_3__915_, data_stage_3__914_, data_stage_3__913_, data_stage_3__912_, data_stage_3__911_, data_stage_3__910_, data_stage_3__909_, data_stage_3__908_, data_stage_3__907_, data_stage_3__906_, data_stage_3__905_, data_stage_3__904_, data_stage_3__903_, data_stage_3__902_, data_stage_3__901_, data_stage_3__900_, data_stage_3__899_, data_stage_3__898_, data_stage_3__897_, data_stage_3__896_, data_stage_3__895_, data_stage_3__894_, data_stage_3__893_, data_stage_3__892_, data_stage_3__891_, data_stage_3__890_, data_stage_3__889_, data_stage_3__888_, data_stage_3__887_, data_stage_3__886_, data_stage_3__885_, data_stage_3__884_, data_stage_3__883_, data_stage_3__882_, data_stage_3__881_, data_stage_3__880_, data_stage_3__879_, data_stage_3__878_, data_stage_3__877_, data_stage_3__876_, data_stage_3__875_, data_stage_3__874_, data_stage_3__873_, data_stage_3__872_, data_stage_3__871_, data_stage_3__870_, data_stage_3__869_, data_stage_3__868_, data_stage_3__867_, data_stage_3__866_, data_stage_3__865_, data_stage_3__864_, data_stage_3__863_, data_stage_3__862_, data_stage_3__861_, data_stage_3__860_, data_stage_3__859_, data_stage_3__858_, data_stage_3__857_, data_stage_3__856_, data_stage_3__855_, data_stage_3__854_, data_stage_3__853_, data_stage_3__852_, data_stage_3__851_, data_stage_3__850_, data_stage_3__849_, data_stage_3__848_, data_stage_3__847_, data_stage_3__846_, data_stage_3__845_, data_stage_3__844_, data_stage_3__843_, data_stage_3__842_, data_stage_3__841_, data_stage_3__840_, data_stage_3__839_, data_stage_3__838_, data_stage_3__837_, data_stage_3__836_, data_stage_3__835_, data_stage_3__834_, data_stage_3__833_, data_stage_3__832_, data_stage_3__831_, data_stage_3__830_, data_stage_3__829_, data_stage_3__828_, data_stage_3__827_, data_stage_3__826_, data_stage_3__825_, data_stage_3__824_, data_stage_3__823_, data_stage_3__822_, data_stage_3__821_, data_stage_3__820_, data_stage_3__819_, data_stage_3__818_, data_stage_3__817_, data_stage_3__816_, data_stage_3__815_, data_stage_3__814_, data_stage_3__813_, data_stage_3__812_, data_stage_3__811_, data_stage_3__810_, data_stage_3__809_, data_stage_3__808_, data_stage_3__807_, data_stage_3__806_, data_stage_3__805_, data_stage_3__804_, data_stage_3__803_, data_stage_3__802_, data_stage_3__801_, data_stage_3__800_, data_stage_3__799_, data_stage_3__798_, data_stage_3__797_, data_stage_3__796_, data_stage_3__795_, data_stage_3__794_, data_stage_3__793_, data_stage_3__792_, data_stage_3__791_, data_stage_3__790_, data_stage_3__789_, data_stage_3__788_, data_stage_3__787_, data_stage_3__786_, data_stage_3__785_, data_stage_3__784_, data_stage_3__783_, data_stage_3__782_, data_stage_3__781_, data_stage_3__780_, data_stage_3__779_, data_stage_3__778_, data_stage_3__777_, data_stage_3__776_, data_stage_3__775_, data_stage_3__774_, data_stage_3__773_, data_stage_3__772_, data_stage_3__771_, data_stage_3__770_, data_stage_3__769_, data_stage_3__768_, data_stage_3__767_, data_stage_3__766_, data_stage_3__765_, data_stage_3__764_, data_stage_3__763_, data_stage_3__762_, data_stage_3__761_, data_stage_3__760_, data_stage_3__759_, data_stage_3__758_, data_stage_3__757_, data_stage_3__756_, data_stage_3__755_, data_stage_3__754_, data_stage_3__753_, data_stage_3__752_, data_stage_3__751_, data_stage_3__750_, data_stage_3__749_, data_stage_3__748_, data_stage_3__747_, data_stage_3__746_, data_stage_3__745_, data_stage_3__744_, data_stage_3__743_, data_stage_3__742_, data_stage_3__741_, data_stage_3__740_, data_stage_3__739_, data_stage_3__738_, data_stage_3__737_, data_stage_3__736_, data_stage_3__735_, data_stage_3__734_, data_stage_3__733_, data_stage_3__732_, data_stage_3__731_, data_stage_3__730_, data_stage_3__729_, data_stage_3__728_, data_stage_3__727_, data_stage_3__726_, data_stage_3__725_, data_stage_3__724_, data_stage_3__723_, data_stage_3__722_, data_stage_3__721_, data_stage_3__720_, data_stage_3__719_, data_stage_3__718_, data_stage_3__717_, data_stage_3__716_, data_stage_3__715_, data_stage_3__714_, data_stage_3__713_, data_stage_3__712_, data_stage_3__711_, data_stage_3__710_, data_stage_3__709_, data_stage_3__708_, data_stage_3__707_, data_stage_3__706_, data_stage_3__705_, data_stage_3__704_, data_stage_3__703_, data_stage_3__702_, data_stage_3__701_, data_stage_3__700_, data_stage_3__699_, data_stage_3__698_, data_stage_3__697_, data_stage_3__696_, data_stage_3__695_, data_stage_3__694_, data_stage_3__693_, data_stage_3__692_, data_stage_3__691_, data_stage_3__690_, data_stage_3__689_, data_stage_3__688_, data_stage_3__687_, data_stage_3__686_, data_stage_3__685_, data_stage_3__684_, data_stage_3__683_, data_stage_3__682_, data_stage_3__681_, data_stage_3__680_, data_stage_3__679_, data_stage_3__678_, data_stage_3__677_, data_stage_3__676_, data_stage_3__675_, data_stage_3__674_, data_stage_3__673_, data_stage_3__672_, data_stage_3__671_, data_stage_3__670_, data_stage_3__669_, data_stage_3__668_, data_stage_3__667_, data_stage_3__666_, data_stage_3__665_, data_stage_3__664_, data_stage_3__663_, data_stage_3__662_, data_stage_3__661_, data_stage_3__660_, data_stage_3__659_, data_stage_3__658_, data_stage_3__657_, data_stage_3__656_, data_stage_3__655_, data_stage_3__654_, data_stage_3__653_, data_stage_3__652_, data_stage_3__651_, data_stage_3__650_, data_stage_3__649_, data_stage_3__648_, data_stage_3__647_, data_stage_3__646_, data_stage_3__645_, data_stage_3__644_, data_stage_3__643_, data_stage_3__642_, data_stage_3__641_, data_stage_3__640_, data_stage_3__639_, data_stage_3__638_, data_stage_3__637_, data_stage_3__636_, data_stage_3__635_, data_stage_3__634_, data_stage_3__633_, data_stage_3__632_, data_stage_3__631_, data_stage_3__630_, data_stage_3__629_, data_stage_3__628_, data_stage_3__627_, data_stage_3__626_, data_stage_3__625_, data_stage_3__624_, data_stage_3__623_, data_stage_3__622_, data_stage_3__621_, data_stage_3__620_, data_stage_3__619_, data_stage_3__618_, data_stage_3__617_, data_stage_3__616_, data_stage_3__615_, data_stage_3__614_, data_stage_3__613_, data_stage_3__612_, data_stage_3__611_, data_stage_3__610_, data_stage_3__609_, data_stage_3__608_, data_stage_3__607_, data_stage_3__606_, data_stage_3__605_, data_stage_3__604_, data_stage_3__603_, data_stage_3__602_, data_stage_3__601_, data_stage_3__600_, data_stage_3__599_, data_stage_3__598_, data_stage_3__597_, data_stage_3__596_, data_stage_3__595_, data_stage_3__594_, data_stage_3__593_, data_stage_3__592_, data_stage_3__591_, data_stage_3__590_, data_stage_3__589_, data_stage_3__588_, data_stage_3__587_, data_stage_3__586_, data_stage_3__585_, data_stage_3__584_, data_stage_3__583_, data_stage_3__582_, data_stage_3__581_, data_stage_3__580_, data_stage_3__579_, data_stage_3__578_, data_stage_3__577_, data_stage_3__576_, data_stage_3__575_, data_stage_3__574_, data_stage_3__573_, data_stage_3__572_, data_stage_3__571_, data_stage_3__570_, data_stage_3__569_, data_stage_3__568_, data_stage_3__567_, data_stage_3__566_, data_stage_3__565_, data_stage_3__564_, data_stage_3__563_, data_stage_3__562_, data_stage_3__561_, data_stage_3__560_, data_stage_3__559_, data_stage_3__558_, data_stage_3__557_, data_stage_3__556_, data_stage_3__555_, data_stage_3__554_, data_stage_3__553_, data_stage_3__552_, data_stage_3__551_, data_stage_3__550_, data_stage_3__549_, data_stage_3__548_, data_stage_3__547_, data_stage_3__546_, data_stage_3__545_, data_stage_3__544_, data_stage_3__543_, data_stage_3__542_, data_stage_3__541_, data_stage_3__540_, data_stage_3__539_, data_stage_3__538_, data_stage_3__537_, data_stage_3__536_, data_stage_3__535_, data_stage_3__534_, data_stage_3__533_, data_stage_3__532_, data_stage_3__531_, data_stage_3__530_, data_stage_3__529_, data_stage_3__528_, data_stage_3__527_, data_stage_3__526_, data_stage_3__525_, data_stage_3__524_, data_stage_3__523_, data_stage_3__522_, data_stage_3__521_, data_stage_3__520_, data_stage_3__519_, data_stage_3__518_, data_stage_3__517_, data_stage_3__516_, data_stage_3__515_, data_stage_3__514_, data_stage_3__513_, data_stage_3__512_, data_stage_3__511_, data_stage_3__510_, data_stage_3__509_, data_stage_3__508_, data_stage_3__507_, data_stage_3__506_, data_stage_3__505_, data_stage_3__504_, data_stage_3__503_, data_stage_3__502_, data_stage_3__501_, data_stage_3__500_, data_stage_3__499_, data_stage_3__498_, data_stage_3__497_, data_stage_3__496_, data_stage_3__495_, data_stage_3__494_, data_stage_3__493_, data_stage_3__492_, data_stage_3__491_, data_stage_3__490_, data_stage_3__489_, data_stage_3__488_, data_stage_3__487_, data_stage_3__486_, data_stage_3__485_, data_stage_3__484_, data_stage_3__483_, data_stage_3__482_, data_stage_3__481_, data_stage_3__480_, data_stage_3__479_, data_stage_3__478_, data_stage_3__477_, data_stage_3__476_, data_stage_3__475_, data_stage_3__474_, data_stage_3__473_, data_stage_3__472_, data_stage_3__471_, data_stage_3__470_, data_stage_3__469_, data_stage_3__468_, data_stage_3__467_, data_stage_3__466_, data_stage_3__465_, data_stage_3__464_, data_stage_3__463_, data_stage_3__462_, data_stage_3__461_, data_stage_3__460_, data_stage_3__459_, data_stage_3__458_, data_stage_3__457_, data_stage_3__456_, data_stage_3__455_, data_stage_3__454_, data_stage_3__453_, data_stage_3__452_, data_stage_3__451_, data_stage_3__450_, data_stage_3__449_, data_stage_3__448_, data_stage_3__447_, data_stage_3__446_, data_stage_3__445_, data_stage_3__444_, data_stage_3__443_, data_stage_3__442_, data_stage_3__441_, data_stage_3__440_, data_stage_3__439_, data_stage_3__438_, data_stage_3__437_, data_stage_3__436_, data_stage_3__435_, data_stage_3__434_, data_stage_3__433_, data_stage_3__432_, data_stage_3__431_, data_stage_3__430_, data_stage_3__429_, data_stage_3__428_, data_stage_3__427_, data_stage_3__426_, data_stage_3__425_, data_stage_3__424_, data_stage_3__423_, data_stage_3__422_, data_stage_3__421_, data_stage_3__420_, data_stage_3__419_, data_stage_3__418_, data_stage_3__417_, data_stage_3__416_, data_stage_3__415_, data_stage_3__414_, data_stage_3__413_, data_stage_3__412_, data_stage_3__411_, data_stage_3__410_, data_stage_3__409_, data_stage_3__408_, data_stage_3__407_, data_stage_3__406_, data_stage_3__405_, data_stage_3__404_, data_stage_3__403_, data_stage_3__402_, data_stage_3__401_, data_stage_3__400_, data_stage_3__399_, data_stage_3__398_, data_stage_3__397_, data_stage_3__396_, data_stage_3__395_, data_stage_3__394_, data_stage_3__393_, data_stage_3__392_, data_stage_3__391_, data_stage_3__390_, data_stage_3__389_, data_stage_3__388_, data_stage_3__387_, data_stage_3__386_, data_stage_3__385_, data_stage_3__384_, data_stage_3__383_, data_stage_3__382_, data_stage_3__381_, data_stage_3__380_, data_stage_3__379_, data_stage_3__378_, data_stage_3__377_, data_stage_3__376_, data_stage_3__375_, data_stage_3__374_, data_stage_3__373_, data_stage_3__372_, data_stage_3__371_, data_stage_3__370_, data_stage_3__369_, data_stage_3__368_, data_stage_3__367_, data_stage_3__366_, data_stage_3__365_, data_stage_3__364_, data_stage_3__363_, data_stage_3__362_, data_stage_3__361_, data_stage_3__360_, data_stage_3__359_, data_stage_3__358_, data_stage_3__357_, data_stage_3__356_, data_stage_3__355_, data_stage_3__354_, data_stage_3__353_, data_stage_3__352_, data_stage_3__351_, data_stage_3__350_, data_stage_3__349_, data_stage_3__348_, data_stage_3__347_, data_stage_3__346_, data_stage_3__345_, data_stage_3__344_, data_stage_3__343_, data_stage_3__342_, data_stage_3__341_, data_stage_3__340_, data_stage_3__339_, data_stage_3__338_, data_stage_3__337_, data_stage_3__336_, data_stage_3__335_, data_stage_3__334_, data_stage_3__333_, data_stage_3__332_, data_stage_3__331_, data_stage_3__330_, data_stage_3__329_, data_stage_3__328_, data_stage_3__327_, data_stage_3__326_, data_stage_3__325_, data_stage_3__324_, data_stage_3__323_, data_stage_3__322_, data_stage_3__321_, data_stage_3__320_, data_stage_3__319_, data_stage_3__318_, data_stage_3__317_, data_stage_3__316_, data_stage_3__315_, data_stage_3__314_, data_stage_3__313_, data_stage_3__312_, data_stage_3__311_, data_stage_3__310_, data_stage_3__309_, data_stage_3__308_, data_stage_3__307_, data_stage_3__306_, data_stage_3__305_, data_stage_3__304_, data_stage_3__303_, data_stage_3__302_, data_stage_3__301_, data_stage_3__300_, data_stage_3__299_, data_stage_3__298_, data_stage_3__297_, data_stage_3__296_, data_stage_3__295_, data_stage_3__294_, data_stage_3__293_, data_stage_3__292_, data_stage_3__291_, data_stage_3__290_, data_stage_3__289_, data_stage_3__288_, data_stage_3__287_, data_stage_3__286_, data_stage_3__285_, data_stage_3__284_, data_stage_3__283_, data_stage_3__282_, data_stage_3__281_, data_stage_3__280_, data_stage_3__279_, data_stage_3__278_, data_stage_3__277_, data_stage_3__276_, data_stage_3__275_, data_stage_3__274_, data_stage_3__273_, data_stage_3__272_, data_stage_3__271_, data_stage_3__270_, data_stage_3__269_, data_stage_3__268_, data_stage_3__267_, data_stage_3__266_, data_stage_3__265_, data_stage_3__264_, data_stage_3__263_, data_stage_3__262_, data_stage_3__261_, data_stage_3__260_, data_stage_3__259_, data_stage_3__258_, data_stage_3__257_, data_stage_3__256_, data_stage_3__255_, data_stage_3__254_, data_stage_3__253_, data_stage_3__252_, data_stage_3__251_, data_stage_3__250_, data_stage_3__249_, data_stage_3__248_, data_stage_3__247_, data_stage_3__246_, data_stage_3__245_, data_stage_3__244_, data_stage_3__243_, data_stage_3__242_, data_stage_3__241_, data_stage_3__240_, data_stage_3__239_, data_stage_3__238_, data_stage_3__237_, data_stage_3__236_, data_stage_3__235_, data_stage_3__234_, data_stage_3__233_, data_stage_3__232_, data_stage_3__231_, data_stage_3__230_, data_stage_3__229_, data_stage_3__228_, data_stage_3__227_, data_stage_3__226_, data_stage_3__225_, data_stage_3__224_, data_stage_3__223_, data_stage_3__222_, data_stage_3__221_, data_stage_3__220_, data_stage_3__219_, data_stage_3__218_, data_stage_3__217_, data_stage_3__216_, data_stage_3__215_, data_stage_3__214_, data_stage_3__213_, data_stage_3__212_, data_stage_3__211_, data_stage_3__210_, data_stage_3__209_, data_stage_3__208_, data_stage_3__207_, data_stage_3__206_, data_stage_3__205_, data_stage_3__204_, data_stage_3__203_, data_stage_3__202_, data_stage_3__201_, data_stage_3__200_, data_stage_3__199_, data_stage_3__198_, data_stage_3__197_, data_stage_3__196_, data_stage_3__195_, data_stage_3__194_, data_stage_3__193_, data_stage_3__192_, data_stage_3__191_, data_stage_3__190_, data_stage_3__189_, data_stage_3__188_, data_stage_3__187_, data_stage_3__186_, data_stage_3__185_, data_stage_3__184_, data_stage_3__183_, data_stage_3__182_, data_stage_3__181_, data_stage_3__180_, data_stage_3__179_, data_stage_3__178_, data_stage_3__177_, data_stage_3__176_, data_stage_3__175_, data_stage_3__174_, data_stage_3__173_, data_stage_3__172_, data_stage_3__171_, data_stage_3__170_, data_stage_3__169_, data_stage_3__168_, data_stage_3__167_, data_stage_3__166_, data_stage_3__165_, data_stage_3__164_, data_stage_3__163_, data_stage_3__162_, data_stage_3__161_, data_stage_3__160_, data_stage_3__159_, data_stage_3__158_, data_stage_3__157_, data_stage_3__156_, data_stage_3__155_, data_stage_3__154_, data_stage_3__153_, data_stage_3__152_, data_stage_3__151_, data_stage_3__150_, data_stage_3__149_, data_stage_3__148_, data_stage_3__147_, data_stage_3__146_, data_stage_3__145_, data_stage_3__144_, data_stage_3__143_, data_stage_3__142_, data_stage_3__141_, data_stage_3__140_, data_stage_3__139_, data_stage_3__138_, data_stage_3__137_, data_stage_3__136_, data_stage_3__135_, data_stage_3__134_, data_stage_3__133_, data_stage_3__132_, data_stage_3__131_, data_stage_3__130_, data_stage_3__129_, data_stage_3__128_, data_stage_3__127_, data_stage_3__126_, data_stage_3__125_, data_stage_3__124_, data_stage_3__123_, data_stage_3__122_, data_stage_3__121_, data_stage_3__120_, data_stage_3__119_, data_stage_3__118_, data_stage_3__117_, data_stage_3__116_, data_stage_3__115_, data_stage_3__114_, data_stage_3__113_, data_stage_3__112_, data_stage_3__111_, data_stage_3__110_, data_stage_3__109_, data_stage_3__108_, data_stage_3__107_, data_stage_3__106_, data_stage_3__105_, data_stage_3__104_, data_stage_3__103_, data_stage_3__102_, data_stage_3__101_, data_stage_3__100_, data_stage_3__99_, data_stage_3__98_, data_stage_3__97_, data_stage_3__96_, data_stage_3__95_, data_stage_3__94_, data_stage_3__93_, data_stage_3__92_, data_stage_3__91_, data_stage_3__90_, data_stage_3__89_, data_stage_3__88_, data_stage_3__87_, data_stage_3__86_, data_stage_3__85_, data_stage_3__84_, data_stage_3__83_, data_stage_3__82_, data_stage_3__81_, data_stage_3__80_, data_stage_3__79_, data_stage_3__78_, data_stage_3__77_, data_stage_3__76_, data_stage_3__75_, data_stage_3__74_, data_stage_3__73_, data_stage_3__72_, data_stage_3__71_, data_stage_3__70_, data_stage_3__69_, data_stage_3__68_, data_stage_3__67_, data_stage_3__66_, data_stage_3__65_, data_stage_3__64_, data_stage_3__63_, data_stage_3__62_, data_stage_3__61_, data_stage_3__60_, data_stage_3__59_, data_stage_3__58_, data_stage_3__57_, data_stage_3__56_, data_stage_3__55_, data_stage_3__54_, data_stage_3__53_, data_stage_3__52_, data_stage_3__51_, data_stage_3__50_, data_stage_3__49_, data_stage_3__48_, data_stage_3__47_, data_stage_3__46_, data_stage_3__45_, data_stage_3__44_, data_stage_3__43_, data_stage_3__42_, data_stage_3__41_, data_stage_3__40_, data_stage_3__39_, data_stage_3__38_, data_stage_3__37_, data_stage_3__36_, data_stage_3__35_, data_stage_3__34_, data_stage_3__33_, data_stage_3__32_, data_stage_3__31_, data_stage_3__30_, data_stage_3__29_, data_stage_3__28_, data_stage_3__27_, data_stage_3__26_, data_stage_3__25_, data_stage_3__24_, data_stage_3__23_, data_stage_3__22_, data_stage_3__21_, data_stage_3__20_, data_stage_3__19_, data_stage_3__18_, data_stage_3__17_, data_stage_3__16_, data_stage_3__15_, data_stage_3__14_, data_stage_3__13_, data_stage_3__12_, data_stage_3__11_, data_stage_3__10_, data_stage_3__9_, data_stage_3__8_, data_stage_3__7_, data_stage_3__6_, data_stage_3__5_, data_stage_3__4_, data_stage_3__3_, data_stage_3__2_, data_stage_3__1_, data_stage_3__0_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__2047_, data_stage_4__2046_, data_stage_4__2045_, data_stage_4__2044_, data_stage_4__2043_, data_stage_4__2042_, data_stage_4__2041_, data_stage_4__2040_, data_stage_4__2039_, data_stage_4__2038_, data_stage_4__2037_, data_stage_4__2036_, data_stage_4__2035_, data_stage_4__2034_, data_stage_4__2033_, data_stage_4__2032_, data_stage_4__2031_, data_stage_4__2030_, data_stage_4__2029_, data_stage_4__2028_, data_stage_4__2027_, data_stage_4__2026_, data_stage_4__2025_, data_stage_4__2024_, data_stage_4__2023_, data_stage_4__2022_, data_stage_4__2021_, data_stage_4__2020_, data_stage_4__2019_, data_stage_4__2018_, data_stage_4__2017_, data_stage_4__2016_, data_stage_4__2015_, data_stage_4__2014_, data_stage_4__2013_, data_stage_4__2012_, data_stage_4__2011_, data_stage_4__2010_, data_stage_4__2009_, data_stage_4__2008_, data_stage_4__2007_, data_stage_4__2006_, data_stage_4__2005_, data_stage_4__2004_, data_stage_4__2003_, data_stage_4__2002_, data_stage_4__2001_, data_stage_4__2000_, data_stage_4__1999_, data_stage_4__1998_, data_stage_4__1997_, data_stage_4__1996_, data_stage_4__1995_, data_stage_4__1994_, data_stage_4__1993_, data_stage_4__1992_, data_stage_4__1991_, data_stage_4__1990_, data_stage_4__1989_, data_stage_4__1988_, data_stage_4__1987_, data_stage_4__1986_, data_stage_4__1985_, data_stage_4__1984_, data_stage_4__1983_, data_stage_4__1982_, data_stage_4__1981_, data_stage_4__1980_, data_stage_4__1979_, data_stage_4__1978_, data_stage_4__1977_, data_stage_4__1976_, data_stage_4__1975_, data_stage_4__1974_, data_stage_4__1973_, data_stage_4__1972_, data_stage_4__1971_, data_stage_4__1970_, data_stage_4__1969_, data_stage_4__1968_, data_stage_4__1967_, data_stage_4__1966_, data_stage_4__1965_, data_stage_4__1964_, data_stage_4__1963_, data_stage_4__1962_, data_stage_4__1961_, data_stage_4__1960_, data_stage_4__1959_, data_stage_4__1958_, data_stage_4__1957_, data_stage_4__1956_, data_stage_4__1955_, data_stage_4__1954_, data_stage_4__1953_, data_stage_4__1952_, data_stage_4__1951_, data_stage_4__1950_, data_stage_4__1949_, data_stage_4__1948_, data_stage_4__1947_, data_stage_4__1946_, data_stage_4__1945_, data_stage_4__1944_, data_stage_4__1943_, data_stage_4__1942_, data_stage_4__1941_, data_stage_4__1940_, data_stage_4__1939_, data_stage_4__1938_, data_stage_4__1937_, data_stage_4__1936_, data_stage_4__1935_, data_stage_4__1934_, data_stage_4__1933_, data_stage_4__1932_, data_stage_4__1931_, data_stage_4__1930_, data_stage_4__1929_, data_stage_4__1928_, data_stage_4__1927_, data_stage_4__1926_, data_stage_4__1925_, data_stage_4__1924_, data_stage_4__1923_, data_stage_4__1922_, data_stage_4__1921_, data_stage_4__1920_, data_stage_4__1919_, data_stage_4__1918_, data_stage_4__1917_, data_stage_4__1916_, data_stage_4__1915_, data_stage_4__1914_, data_stage_4__1913_, data_stage_4__1912_, data_stage_4__1911_, data_stage_4__1910_, data_stage_4__1909_, data_stage_4__1908_, data_stage_4__1907_, data_stage_4__1906_, data_stage_4__1905_, data_stage_4__1904_, data_stage_4__1903_, data_stage_4__1902_, data_stage_4__1901_, data_stage_4__1900_, data_stage_4__1899_, data_stage_4__1898_, data_stage_4__1897_, data_stage_4__1896_, data_stage_4__1895_, data_stage_4__1894_, data_stage_4__1893_, data_stage_4__1892_, data_stage_4__1891_, data_stage_4__1890_, data_stage_4__1889_, data_stage_4__1888_, data_stage_4__1887_, data_stage_4__1886_, data_stage_4__1885_, data_stage_4__1884_, data_stage_4__1883_, data_stage_4__1882_, data_stage_4__1881_, data_stage_4__1880_, data_stage_4__1879_, data_stage_4__1878_, data_stage_4__1877_, data_stage_4__1876_, data_stage_4__1875_, data_stage_4__1874_, data_stage_4__1873_, data_stage_4__1872_, data_stage_4__1871_, data_stage_4__1870_, data_stage_4__1869_, data_stage_4__1868_, data_stage_4__1867_, data_stage_4__1866_, data_stage_4__1865_, data_stage_4__1864_, data_stage_4__1863_, data_stage_4__1862_, data_stage_4__1861_, data_stage_4__1860_, data_stage_4__1859_, data_stage_4__1858_, data_stage_4__1857_, data_stage_4__1856_, data_stage_4__1855_, data_stage_4__1854_, data_stage_4__1853_, data_stage_4__1852_, data_stage_4__1851_, data_stage_4__1850_, data_stage_4__1849_, data_stage_4__1848_, data_stage_4__1847_, data_stage_4__1846_, data_stage_4__1845_, data_stage_4__1844_, data_stage_4__1843_, data_stage_4__1842_, data_stage_4__1841_, data_stage_4__1840_, data_stage_4__1839_, data_stage_4__1838_, data_stage_4__1837_, data_stage_4__1836_, data_stage_4__1835_, data_stage_4__1834_, data_stage_4__1833_, data_stage_4__1832_, data_stage_4__1831_, data_stage_4__1830_, data_stage_4__1829_, data_stage_4__1828_, data_stage_4__1827_, data_stage_4__1826_, data_stage_4__1825_, data_stage_4__1824_, data_stage_4__1823_, data_stage_4__1822_, data_stage_4__1821_, data_stage_4__1820_, data_stage_4__1819_, data_stage_4__1818_, data_stage_4__1817_, data_stage_4__1816_, data_stage_4__1815_, data_stage_4__1814_, data_stage_4__1813_, data_stage_4__1812_, data_stage_4__1811_, data_stage_4__1810_, data_stage_4__1809_, data_stage_4__1808_, data_stage_4__1807_, data_stage_4__1806_, data_stage_4__1805_, data_stage_4__1804_, data_stage_4__1803_, data_stage_4__1802_, data_stage_4__1801_, data_stage_4__1800_, data_stage_4__1799_, data_stage_4__1798_, data_stage_4__1797_, data_stage_4__1796_, data_stage_4__1795_, data_stage_4__1794_, data_stage_4__1793_, data_stage_4__1792_, data_stage_4__1791_, data_stage_4__1790_, data_stage_4__1789_, data_stage_4__1788_, data_stage_4__1787_, data_stage_4__1786_, data_stage_4__1785_, data_stage_4__1784_, data_stage_4__1783_, data_stage_4__1782_, data_stage_4__1781_, data_stage_4__1780_, data_stage_4__1779_, data_stage_4__1778_, data_stage_4__1777_, data_stage_4__1776_, data_stage_4__1775_, data_stage_4__1774_, data_stage_4__1773_, data_stage_4__1772_, data_stage_4__1771_, data_stage_4__1770_, data_stage_4__1769_, data_stage_4__1768_, data_stage_4__1767_, data_stage_4__1766_, data_stage_4__1765_, data_stage_4__1764_, data_stage_4__1763_, data_stage_4__1762_, data_stage_4__1761_, data_stage_4__1760_, data_stage_4__1759_, data_stage_4__1758_, data_stage_4__1757_, data_stage_4__1756_, data_stage_4__1755_, data_stage_4__1754_, data_stage_4__1753_, data_stage_4__1752_, data_stage_4__1751_, data_stage_4__1750_, data_stage_4__1749_, data_stage_4__1748_, data_stage_4__1747_, data_stage_4__1746_, data_stage_4__1745_, data_stage_4__1744_, data_stage_4__1743_, data_stage_4__1742_, data_stage_4__1741_, data_stage_4__1740_, data_stage_4__1739_, data_stage_4__1738_, data_stage_4__1737_, data_stage_4__1736_, data_stage_4__1735_, data_stage_4__1734_, data_stage_4__1733_, data_stage_4__1732_, data_stage_4__1731_, data_stage_4__1730_, data_stage_4__1729_, data_stage_4__1728_, data_stage_4__1727_, data_stage_4__1726_, data_stage_4__1725_, data_stage_4__1724_, data_stage_4__1723_, data_stage_4__1722_, data_stage_4__1721_, data_stage_4__1720_, data_stage_4__1719_, data_stage_4__1718_, data_stage_4__1717_, data_stage_4__1716_, data_stage_4__1715_, data_stage_4__1714_, data_stage_4__1713_, data_stage_4__1712_, data_stage_4__1711_, data_stage_4__1710_, data_stage_4__1709_, data_stage_4__1708_, data_stage_4__1707_, data_stage_4__1706_, data_stage_4__1705_, data_stage_4__1704_, data_stage_4__1703_, data_stage_4__1702_, data_stage_4__1701_, data_stage_4__1700_, data_stage_4__1699_, data_stage_4__1698_, data_stage_4__1697_, data_stage_4__1696_, data_stage_4__1695_, data_stage_4__1694_, data_stage_4__1693_, data_stage_4__1692_, data_stage_4__1691_, data_stage_4__1690_, data_stage_4__1689_, data_stage_4__1688_, data_stage_4__1687_, data_stage_4__1686_, data_stage_4__1685_, data_stage_4__1684_, data_stage_4__1683_, data_stage_4__1682_, data_stage_4__1681_, data_stage_4__1680_, data_stage_4__1679_, data_stage_4__1678_, data_stage_4__1677_, data_stage_4__1676_, data_stage_4__1675_, data_stage_4__1674_, data_stage_4__1673_, data_stage_4__1672_, data_stage_4__1671_, data_stage_4__1670_, data_stage_4__1669_, data_stage_4__1668_, data_stage_4__1667_, data_stage_4__1666_, data_stage_4__1665_, data_stage_4__1664_, data_stage_4__1663_, data_stage_4__1662_, data_stage_4__1661_, data_stage_4__1660_, data_stage_4__1659_, data_stage_4__1658_, data_stage_4__1657_, data_stage_4__1656_, data_stage_4__1655_, data_stage_4__1654_, data_stage_4__1653_, data_stage_4__1652_, data_stage_4__1651_, data_stage_4__1650_, data_stage_4__1649_, data_stage_4__1648_, data_stage_4__1647_, data_stage_4__1646_, data_stage_4__1645_, data_stage_4__1644_, data_stage_4__1643_, data_stage_4__1642_, data_stage_4__1641_, data_stage_4__1640_, data_stage_4__1639_, data_stage_4__1638_, data_stage_4__1637_, data_stage_4__1636_, data_stage_4__1635_, data_stage_4__1634_, data_stage_4__1633_, data_stage_4__1632_, data_stage_4__1631_, data_stage_4__1630_, data_stage_4__1629_, data_stage_4__1628_, data_stage_4__1627_, data_stage_4__1626_, data_stage_4__1625_, data_stage_4__1624_, data_stage_4__1623_, data_stage_4__1622_, data_stage_4__1621_, data_stage_4__1620_, data_stage_4__1619_, data_stage_4__1618_, data_stage_4__1617_, data_stage_4__1616_, data_stage_4__1615_, data_stage_4__1614_, data_stage_4__1613_, data_stage_4__1612_, data_stage_4__1611_, data_stage_4__1610_, data_stage_4__1609_, data_stage_4__1608_, data_stage_4__1607_, data_stage_4__1606_, data_stage_4__1605_, data_stage_4__1604_, data_stage_4__1603_, data_stage_4__1602_, data_stage_4__1601_, data_stage_4__1600_, data_stage_4__1599_, data_stage_4__1598_, data_stage_4__1597_, data_stage_4__1596_, data_stage_4__1595_, data_stage_4__1594_, data_stage_4__1593_, data_stage_4__1592_, data_stage_4__1591_, data_stage_4__1590_, data_stage_4__1589_, data_stage_4__1588_, data_stage_4__1587_, data_stage_4__1586_, data_stage_4__1585_, data_stage_4__1584_, data_stage_4__1583_, data_stage_4__1582_, data_stage_4__1581_, data_stage_4__1580_, data_stage_4__1579_, data_stage_4__1578_, data_stage_4__1577_, data_stage_4__1576_, data_stage_4__1575_, data_stage_4__1574_, data_stage_4__1573_, data_stage_4__1572_, data_stage_4__1571_, data_stage_4__1570_, data_stage_4__1569_, data_stage_4__1568_, data_stage_4__1567_, data_stage_4__1566_, data_stage_4__1565_, data_stage_4__1564_, data_stage_4__1563_, data_stage_4__1562_, data_stage_4__1561_, data_stage_4__1560_, data_stage_4__1559_, data_stage_4__1558_, data_stage_4__1557_, data_stage_4__1556_, data_stage_4__1555_, data_stage_4__1554_, data_stage_4__1553_, data_stage_4__1552_, data_stage_4__1551_, data_stage_4__1550_, data_stage_4__1549_, data_stage_4__1548_, data_stage_4__1547_, data_stage_4__1546_, data_stage_4__1545_, data_stage_4__1544_, data_stage_4__1543_, data_stage_4__1542_, data_stage_4__1541_, data_stage_4__1540_, data_stage_4__1539_, data_stage_4__1538_, data_stage_4__1537_, data_stage_4__1536_, data_stage_4__1535_, data_stage_4__1534_, data_stage_4__1533_, data_stage_4__1532_, data_stage_4__1531_, data_stage_4__1530_, data_stage_4__1529_, data_stage_4__1528_, data_stage_4__1527_, data_stage_4__1526_, data_stage_4__1525_, data_stage_4__1524_, data_stage_4__1523_, data_stage_4__1522_, data_stage_4__1521_, data_stage_4__1520_, data_stage_4__1519_, data_stage_4__1518_, data_stage_4__1517_, data_stage_4__1516_, data_stage_4__1515_, data_stage_4__1514_, data_stage_4__1513_, data_stage_4__1512_, data_stage_4__1511_, data_stage_4__1510_, data_stage_4__1509_, data_stage_4__1508_, data_stage_4__1507_, data_stage_4__1506_, data_stage_4__1505_, data_stage_4__1504_, data_stage_4__1503_, data_stage_4__1502_, data_stage_4__1501_, data_stage_4__1500_, data_stage_4__1499_, data_stage_4__1498_, data_stage_4__1497_, data_stage_4__1496_, data_stage_4__1495_, data_stage_4__1494_, data_stage_4__1493_, data_stage_4__1492_, data_stage_4__1491_, data_stage_4__1490_, data_stage_4__1489_, data_stage_4__1488_, data_stage_4__1487_, data_stage_4__1486_, data_stage_4__1485_, data_stage_4__1484_, data_stage_4__1483_, data_stage_4__1482_, data_stage_4__1481_, data_stage_4__1480_, data_stage_4__1479_, data_stage_4__1478_, data_stage_4__1477_, data_stage_4__1476_, data_stage_4__1475_, data_stage_4__1474_, data_stage_4__1473_, data_stage_4__1472_, data_stage_4__1471_, data_stage_4__1470_, data_stage_4__1469_, data_stage_4__1468_, data_stage_4__1467_, data_stage_4__1466_, data_stage_4__1465_, data_stage_4__1464_, data_stage_4__1463_, data_stage_4__1462_, data_stage_4__1461_, data_stage_4__1460_, data_stage_4__1459_, data_stage_4__1458_, data_stage_4__1457_, data_stage_4__1456_, data_stage_4__1455_, data_stage_4__1454_, data_stage_4__1453_, data_stage_4__1452_, data_stage_4__1451_, data_stage_4__1450_, data_stage_4__1449_, data_stage_4__1448_, data_stage_4__1447_, data_stage_4__1446_, data_stage_4__1445_, data_stage_4__1444_, data_stage_4__1443_, data_stage_4__1442_, data_stage_4__1441_, data_stage_4__1440_, data_stage_4__1439_, data_stage_4__1438_, data_stage_4__1437_, data_stage_4__1436_, data_stage_4__1435_, data_stage_4__1434_, data_stage_4__1433_, data_stage_4__1432_, data_stage_4__1431_, data_stage_4__1430_, data_stage_4__1429_, data_stage_4__1428_, data_stage_4__1427_, data_stage_4__1426_, data_stage_4__1425_, data_stage_4__1424_, data_stage_4__1423_, data_stage_4__1422_, data_stage_4__1421_, data_stage_4__1420_, data_stage_4__1419_, data_stage_4__1418_, data_stage_4__1417_, data_stage_4__1416_, data_stage_4__1415_, data_stage_4__1414_, data_stage_4__1413_, data_stage_4__1412_, data_stage_4__1411_, data_stage_4__1410_, data_stage_4__1409_, data_stage_4__1408_, data_stage_4__1407_, data_stage_4__1406_, data_stage_4__1405_, data_stage_4__1404_, data_stage_4__1403_, data_stage_4__1402_, data_stage_4__1401_, data_stage_4__1400_, data_stage_4__1399_, data_stage_4__1398_, data_stage_4__1397_, data_stage_4__1396_, data_stage_4__1395_, data_stage_4__1394_, data_stage_4__1393_, data_stage_4__1392_, data_stage_4__1391_, data_stage_4__1390_, data_stage_4__1389_, data_stage_4__1388_, data_stage_4__1387_, data_stage_4__1386_, data_stage_4__1385_, data_stage_4__1384_, data_stage_4__1383_, data_stage_4__1382_, data_stage_4__1381_, data_stage_4__1380_, data_stage_4__1379_, data_stage_4__1378_, data_stage_4__1377_, data_stage_4__1376_, data_stage_4__1375_, data_stage_4__1374_, data_stage_4__1373_, data_stage_4__1372_, data_stage_4__1371_, data_stage_4__1370_, data_stage_4__1369_, data_stage_4__1368_, data_stage_4__1367_, data_stage_4__1366_, data_stage_4__1365_, data_stage_4__1364_, data_stage_4__1363_, data_stage_4__1362_, data_stage_4__1361_, data_stage_4__1360_, data_stage_4__1359_, data_stage_4__1358_, data_stage_4__1357_, data_stage_4__1356_, data_stage_4__1355_, data_stage_4__1354_, data_stage_4__1353_, data_stage_4__1352_, data_stage_4__1351_, data_stage_4__1350_, data_stage_4__1349_, data_stage_4__1348_, data_stage_4__1347_, data_stage_4__1346_, data_stage_4__1345_, data_stage_4__1344_, data_stage_4__1343_, data_stage_4__1342_, data_stage_4__1341_, data_stage_4__1340_, data_stage_4__1339_, data_stage_4__1338_, data_stage_4__1337_, data_stage_4__1336_, data_stage_4__1335_, data_stage_4__1334_, data_stage_4__1333_, data_stage_4__1332_, data_stage_4__1331_, data_stage_4__1330_, data_stage_4__1329_, data_stage_4__1328_, data_stage_4__1327_, data_stage_4__1326_, data_stage_4__1325_, data_stage_4__1324_, data_stage_4__1323_, data_stage_4__1322_, data_stage_4__1321_, data_stage_4__1320_, data_stage_4__1319_, data_stage_4__1318_, data_stage_4__1317_, data_stage_4__1316_, data_stage_4__1315_, data_stage_4__1314_, data_stage_4__1313_, data_stage_4__1312_, data_stage_4__1311_, data_stage_4__1310_, data_stage_4__1309_, data_stage_4__1308_, data_stage_4__1307_, data_stage_4__1306_, data_stage_4__1305_, data_stage_4__1304_, data_stage_4__1303_, data_stage_4__1302_, data_stage_4__1301_, data_stage_4__1300_, data_stage_4__1299_, data_stage_4__1298_, data_stage_4__1297_, data_stage_4__1296_, data_stage_4__1295_, data_stage_4__1294_, data_stage_4__1293_, data_stage_4__1292_, data_stage_4__1291_, data_stage_4__1290_, data_stage_4__1289_, data_stage_4__1288_, data_stage_4__1287_, data_stage_4__1286_, data_stage_4__1285_, data_stage_4__1284_, data_stage_4__1283_, data_stage_4__1282_, data_stage_4__1281_, data_stage_4__1280_, data_stage_4__1279_, data_stage_4__1278_, data_stage_4__1277_, data_stage_4__1276_, data_stage_4__1275_, data_stage_4__1274_, data_stage_4__1273_, data_stage_4__1272_, data_stage_4__1271_, data_stage_4__1270_, data_stage_4__1269_, data_stage_4__1268_, data_stage_4__1267_, data_stage_4__1266_, data_stage_4__1265_, data_stage_4__1264_, data_stage_4__1263_, data_stage_4__1262_, data_stage_4__1261_, data_stage_4__1260_, data_stage_4__1259_, data_stage_4__1258_, data_stage_4__1257_, data_stage_4__1256_, data_stage_4__1255_, data_stage_4__1254_, data_stage_4__1253_, data_stage_4__1252_, data_stage_4__1251_, data_stage_4__1250_, data_stage_4__1249_, data_stage_4__1248_, data_stage_4__1247_, data_stage_4__1246_, data_stage_4__1245_, data_stage_4__1244_, data_stage_4__1243_, data_stage_4__1242_, data_stage_4__1241_, data_stage_4__1240_, data_stage_4__1239_, data_stage_4__1238_, data_stage_4__1237_, data_stage_4__1236_, data_stage_4__1235_, data_stage_4__1234_, data_stage_4__1233_, data_stage_4__1232_, data_stage_4__1231_, data_stage_4__1230_, data_stage_4__1229_, data_stage_4__1228_, data_stage_4__1227_, data_stage_4__1226_, data_stage_4__1225_, data_stage_4__1224_, data_stage_4__1223_, data_stage_4__1222_, data_stage_4__1221_, data_stage_4__1220_, data_stage_4__1219_, data_stage_4__1218_, data_stage_4__1217_, data_stage_4__1216_, data_stage_4__1215_, data_stage_4__1214_, data_stage_4__1213_, data_stage_4__1212_, data_stage_4__1211_, data_stage_4__1210_, data_stage_4__1209_, data_stage_4__1208_, data_stage_4__1207_, data_stage_4__1206_, data_stage_4__1205_, data_stage_4__1204_, data_stage_4__1203_, data_stage_4__1202_, data_stage_4__1201_, data_stage_4__1200_, data_stage_4__1199_, data_stage_4__1198_, data_stage_4__1197_, data_stage_4__1196_, data_stage_4__1195_, data_stage_4__1194_, data_stage_4__1193_, data_stage_4__1192_, data_stage_4__1191_, data_stage_4__1190_, data_stage_4__1189_, data_stage_4__1188_, data_stage_4__1187_, data_stage_4__1186_, data_stage_4__1185_, data_stage_4__1184_, data_stage_4__1183_, data_stage_4__1182_, data_stage_4__1181_, data_stage_4__1180_, data_stage_4__1179_, data_stage_4__1178_, data_stage_4__1177_, data_stage_4__1176_, data_stage_4__1175_, data_stage_4__1174_, data_stage_4__1173_, data_stage_4__1172_, data_stage_4__1171_, data_stage_4__1170_, data_stage_4__1169_, data_stage_4__1168_, data_stage_4__1167_, data_stage_4__1166_, data_stage_4__1165_, data_stage_4__1164_, data_stage_4__1163_, data_stage_4__1162_, data_stage_4__1161_, data_stage_4__1160_, data_stage_4__1159_, data_stage_4__1158_, data_stage_4__1157_, data_stage_4__1156_, data_stage_4__1155_, data_stage_4__1154_, data_stage_4__1153_, data_stage_4__1152_, data_stage_4__1151_, data_stage_4__1150_, data_stage_4__1149_, data_stage_4__1148_, data_stage_4__1147_, data_stage_4__1146_, data_stage_4__1145_, data_stage_4__1144_, data_stage_4__1143_, data_stage_4__1142_, data_stage_4__1141_, data_stage_4__1140_, data_stage_4__1139_, data_stage_4__1138_, data_stage_4__1137_, data_stage_4__1136_, data_stage_4__1135_, data_stage_4__1134_, data_stage_4__1133_, data_stage_4__1132_, data_stage_4__1131_, data_stage_4__1130_, data_stage_4__1129_, data_stage_4__1128_, data_stage_4__1127_, data_stage_4__1126_, data_stage_4__1125_, data_stage_4__1124_, data_stage_4__1123_, data_stage_4__1122_, data_stage_4__1121_, data_stage_4__1120_, data_stage_4__1119_, data_stage_4__1118_, data_stage_4__1117_, data_stage_4__1116_, data_stage_4__1115_, data_stage_4__1114_, data_stage_4__1113_, data_stage_4__1112_, data_stage_4__1111_, data_stage_4__1110_, data_stage_4__1109_, data_stage_4__1108_, data_stage_4__1107_, data_stage_4__1106_, data_stage_4__1105_, data_stage_4__1104_, data_stage_4__1103_, data_stage_4__1102_, data_stage_4__1101_, data_stage_4__1100_, data_stage_4__1099_, data_stage_4__1098_, data_stage_4__1097_, data_stage_4__1096_, data_stage_4__1095_, data_stage_4__1094_, data_stage_4__1093_, data_stage_4__1092_, data_stage_4__1091_, data_stage_4__1090_, data_stage_4__1089_, data_stage_4__1088_, data_stage_4__1087_, data_stage_4__1086_, data_stage_4__1085_, data_stage_4__1084_, data_stage_4__1083_, data_stage_4__1082_, data_stage_4__1081_, data_stage_4__1080_, data_stage_4__1079_, data_stage_4__1078_, data_stage_4__1077_, data_stage_4__1076_, data_stage_4__1075_, data_stage_4__1074_, data_stage_4__1073_, data_stage_4__1072_, data_stage_4__1071_, data_stage_4__1070_, data_stage_4__1069_, data_stage_4__1068_, data_stage_4__1067_, data_stage_4__1066_, data_stage_4__1065_, data_stage_4__1064_, data_stage_4__1063_, data_stage_4__1062_, data_stage_4__1061_, data_stage_4__1060_, data_stage_4__1059_, data_stage_4__1058_, data_stage_4__1057_, data_stage_4__1056_, data_stage_4__1055_, data_stage_4__1054_, data_stage_4__1053_, data_stage_4__1052_, data_stage_4__1051_, data_stage_4__1050_, data_stage_4__1049_, data_stage_4__1048_, data_stage_4__1047_, data_stage_4__1046_, data_stage_4__1045_, data_stage_4__1044_, data_stage_4__1043_, data_stage_4__1042_, data_stage_4__1041_, data_stage_4__1040_, data_stage_4__1039_, data_stage_4__1038_, data_stage_4__1037_, data_stage_4__1036_, data_stage_4__1035_, data_stage_4__1034_, data_stage_4__1033_, data_stage_4__1032_, data_stage_4__1031_, data_stage_4__1030_, data_stage_4__1029_, data_stage_4__1028_, data_stage_4__1027_, data_stage_4__1026_, data_stage_4__1025_, data_stage_4__1024_, data_stage_4__1023_, data_stage_4__1022_, data_stage_4__1021_, data_stage_4__1020_, data_stage_4__1019_, data_stage_4__1018_, data_stage_4__1017_, data_stage_4__1016_, data_stage_4__1015_, data_stage_4__1014_, data_stage_4__1013_, data_stage_4__1012_, data_stage_4__1011_, data_stage_4__1010_, data_stage_4__1009_, data_stage_4__1008_, data_stage_4__1007_, data_stage_4__1006_, data_stage_4__1005_, data_stage_4__1004_, data_stage_4__1003_, data_stage_4__1002_, data_stage_4__1001_, data_stage_4__1000_, data_stage_4__999_, data_stage_4__998_, data_stage_4__997_, data_stage_4__996_, data_stage_4__995_, data_stage_4__994_, data_stage_4__993_, data_stage_4__992_, data_stage_4__991_, data_stage_4__990_, data_stage_4__989_, data_stage_4__988_, data_stage_4__987_, data_stage_4__986_, data_stage_4__985_, data_stage_4__984_, data_stage_4__983_, data_stage_4__982_, data_stage_4__981_, data_stage_4__980_, data_stage_4__979_, data_stage_4__978_, data_stage_4__977_, data_stage_4__976_, data_stage_4__975_, data_stage_4__974_, data_stage_4__973_, data_stage_4__972_, data_stage_4__971_, data_stage_4__970_, data_stage_4__969_, data_stage_4__968_, data_stage_4__967_, data_stage_4__966_, data_stage_4__965_, data_stage_4__964_, data_stage_4__963_, data_stage_4__962_, data_stage_4__961_, data_stage_4__960_, data_stage_4__959_, data_stage_4__958_, data_stage_4__957_, data_stage_4__956_, data_stage_4__955_, data_stage_4__954_, data_stage_4__953_, data_stage_4__952_, data_stage_4__951_, data_stage_4__950_, data_stage_4__949_, data_stage_4__948_, data_stage_4__947_, data_stage_4__946_, data_stage_4__945_, data_stage_4__944_, data_stage_4__943_, data_stage_4__942_, data_stage_4__941_, data_stage_4__940_, data_stage_4__939_, data_stage_4__938_, data_stage_4__937_, data_stage_4__936_, data_stage_4__935_, data_stage_4__934_, data_stage_4__933_, data_stage_4__932_, data_stage_4__931_, data_stage_4__930_, data_stage_4__929_, data_stage_4__928_, data_stage_4__927_, data_stage_4__926_, data_stage_4__925_, data_stage_4__924_, data_stage_4__923_, data_stage_4__922_, data_stage_4__921_, data_stage_4__920_, data_stage_4__919_, data_stage_4__918_, data_stage_4__917_, data_stage_4__916_, data_stage_4__915_, data_stage_4__914_, data_stage_4__913_, data_stage_4__912_, data_stage_4__911_, data_stage_4__910_, data_stage_4__909_, data_stage_4__908_, data_stage_4__907_, data_stage_4__906_, data_stage_4__905_, data_stage_4__904_, data_stage_4__903_, data_stage_4__902_, data_stage_4__901_, data_stage_4__900_, data_stage_4__899_, data_stage_4__898_, data_stage_4__897_, data_stage_4__896_, data_stage_4__895_, data_stage_4__894_, data_stage_4__893_, data_stage_4__892_, data_stage_4__891_, data_stage_4__890_, data_stage_4__889_, data_stage_4__888_, data_stage_4__887_, data_stage_4__886_, data_stage_4__885_, data_stage_4__884_, data_stage_4__883_, data_stage_4__882_, data_stage_4__881_, data_stage_4__880_, data_stage_4__879_, data_stage_4__878_, data_stage_4__877_, data_stage_4__876_, data_stage_4__875_, data_stage_4__874_, data_stage_4__873_, data_stage_4__872_, data_stage_4__871_, data_stage_4__870_, data_stage_4__869_, data_stage_4__868_, data_stage_4__867_, data_stage_4__866_, data_stage_4__865_, data_stage_4__864_, data_stage_4__863_, data_stage_4__862_, data_stage_4__861_, data_stage_4__860_, data_stage_4__859_, data_stage_4__858_, data_stage_4__857_, data_stage_4__856_, data_stage_4__855_, data_stage_4__854_, data_stage_4__853_, data_stage_4__852_, data_stage_4__851_, data_stage_4__850_, data_stage_4__849_, data_stage_4__848_, data_stage_4__847_, data_stage_4__846_, data_stage_4__845_, data_stage_4__844_, data_stage_4__843_, data_stage_4__842_, data_stage_4__841_, data_stage_4__840_, data_stage_4__839_, data_stage_4__838_, data_stage_4__837_, data_stage_4__836_, data_stage_4__835_, data_stage_4__834_, data_stage_4__833_, data_stage_4__832_, data_stage_4__831_, data_stage_4__830_, data_stage_4__829_, data_stage_4__828_, data_stage_4__827_, data_stage_4__826_, data_stage_4__825_, data_stage_4__824_, data_stage_4__823_, data_stage_4__822_, data_stage_4__821_, data_stage_4__820_, data_stage_4__819_, data_stage_4__818_, data_stage_4__817_, data_stage_4__816_, data_stage_4__815_, data_stage_4__814_, data_stage_4__813_, data_stage_4__812_, data_stage_4__811_, data_stage_4__810_, data_stage_4__809_, data_stage_4__808_, data_stage_4__807_, data_stage_4__806_, data_stage_4__805_, data_stage_4__804_, data_stage_4__803_, data_stage_4__802_, data_stage_4__801_, data_stage_4__800_, data_stage_4__799_, data_stage_4__798_, data_stage_4__797_, data_stage_4__796_, data_stage_4__795_, data_stage_4__794_, data_stage_4__793_, data_stage_4__792_, data_stage_4__791_, data_stage_4__790_, data_stage_4__789_, data_stage_4__788_, data_stage_4__787_, data_stage_4__786_, data_stage_4__785_, data_stage_4__784_, data_stage_4__783_, data_stage_4__782_, data_stage_4__781_, data_stage_4__780_, data_stage_4__779_, data_stage_4__778_, data_stage_4__777_, data_stage_4__776_, data_stage_4__775_, data_stage_4__774_, data_stage_4__773_, data_stage_4__772_, data_stage_4__771_, data_stage_4__770_, data_stage_4__769_, data_stage_4__768_, data_stage_4__767_, data_stage_4__766_, data_stage_4__765_, data_stage_4__764_, data_stage_4__763_, data_stage_4__762_, data_stage_4__761_, data_stage_4__760_, data_stage_4__759_, data_stage_4__758_, data_stage_4__757_, data_stage_4__756_, data_stage_4__755_, data_stage_4__754_, data_stage_4__753_, data_stage_4__752_, data_stage_4__751_, data_stage_4__750_, data_stage_4__749_, data_stage_4__748_, data_stage_4__747_, data_stage_4__746_, data_stage_4__745_, data_stage_4__744_, data_stage_4__743_, data_stage_4__742_, data_stage_4__741_, data_stage_4__740_, data_stage_4__739_, data_stage_4__738_, data_stage_4__737_, data_stage_4__736_, data_stage_4__735_, data_stage_4__734_, data_stage_4__733_, data_stage_4__732_, data_stage_4__731_, data_stage_4__730_, data_stage_4__729_, data_stage_4__728_, data_stage_4__727_, data_stage_4__726_, data_stage_4__725_, data_stage_4__724_, data_stage_4__723_, data_stage_4__722_, data_stage_4__721_, data_stage_4__720_, data_stage_4__719_, data_stage_4__718_, data_stage_4__717_, data_stage_4__716_, data_stage_4__715_, data_stage_4__714_, data_stage_4__713_, data_stage_4__712_, data_stage_4__711_, data_stage_4__710_, data_stage_4__709_, data_stage_4__708_, data_stage_4__707_, data_stage_4__706_, data_stage_4__705_, data_stage_4__704_, data_stage_4__703_, data_stage_4__702_, data_stage_4__701_, data_stage_4__700_, data_stage_4__699_, data_stage_4__698_, data_stage_4__697_, data_stage_4__696_, data_stage_4__695_, data_stage_4__694_, data_stage_4__693_, data_stage_4__692_, data_stage_4__691_, data_stage_4__690_, data_stage_4__689_, data_stage_4__688_, data_stage_4__687_, data_stage_4__686_, data_stage_4__685_, data_stage_4__684_, data_stage_4__683_, data_stage_4__682_, data_stage_4__681_, data_stage_4__680_, data_stage_4__679_, data_stage_4__678_, data_stage_4__677_, data_stage_4__676_, data_stage_4__675_, data_stage_4__674_, data_stage_4__673_, data_stage_4__672_, data_stage_4__671_, data_stage_4__670_, data_stage_4__669_, data_stage_4__668_, data_stage_4__667_, data_stage_4__666_, data_stage_4__665_, data_stage_4__664_, data_stage_4__663_, data_stage_4__662_, data_stage_4__661_, data_stage_4__660_, data_stage_4__659_, data_stage_4__658_, data_stage_4__657_, data_stage_4__656_, data_stage_4__655_, data_stage_4__654_, data_stage_4__653_, data_stage_4__652_, data_stage_4__651_, data_stage_4__650_, data_stage_4__649_, data_stage_4__648_, data_stage_4__647_, data_stage_4__646_, data_stage_4__645_, data_stage_4__644_, data_stage_4__643_, data_stage_4__642_, data_stage_4__641_, data_stage_4__640_, data_stage_4__639_, data_stage_4__638_, data_stage_4__637_, data_stage_4__636_, data_stage_4__635_, data_stage_4__634_, data_stage_4__633_, data_stage_4__632_, data_stage_4__631_, data_stage_4__630_, data_stage_4__629_, data_stage_4__628_, data_stage_4__627_, data_stage_4__626_, data_stage_4__625_, data_stage_4__624_, data_stage_4__623_, data_stage_4__622_, data_stage_4__621_, data_stage_4__620_, data_stage_4__619_, data_stage_4__618_, data_stage_4__617_, data_stage_4__616_, data_stage_4__615_, data_stage_4__614_, data_stage_4__613_, data_stage_4__612_, data_stage_4__611_, data_stage_4__610_, data_stage_4__609_, data_stage_4__608_, data_stage_4__607_, data_stage_4__606_, data_stage_4__605_, data_stage_4__604_, data_stage_4__603_, data_stage_4__602_, data_stage_4__601_, data_stage_4__600_, data_stage_4__599_, data_stage_4__598_, data_stage_4__597_, data_stage_4__596_, data_stage_4__595_, data_stage_4__594_, data_stage_4__593_, data_stage_4__592_, data_stage_4__591_, data_stage_4__590_, data_stage_4__589_, data_stage_4__588_, data_stage_4__587_, data_stage_4__586_, data_stage_4__585_, data_stage_4__584_, data_stage_4__583_, data_stage_4__582_, data_stage_4__581_, data_stage_4__580_, data_stage_4__579_, data_stage_4__578_, data_stage_4__577_, data_stage_4__576_, data_stage_4__575_, data_stage_4__574_, data_stage_4__573_, data_stage_4__572_, data_stage_4__571_, data_stage_4__570_, data_stage_4__569_, data_stage_4__568_, data_stage_4__567_, data_stage_4__566_, data_stage_4__565_, data_stage_4__564_, data_stage_4__563_, data_stage_4__562_, data_stage_4__561_, data_stage_4__560_, data_stage_4__559_, data_stage_4__558_, data_stage_4__557_, data_stage_4__556_, data_stage_4__555_, data_stage_4__554_, data_stage_4__553_, data_stage_4__552_, data_stage_4__551_, data_stage_4__550_, data_stage_4__549_, data_stage_4__548_, data_stage_4__547_, data_stage_4__546_, data_stage_4__545_, data_stage_4__544_, data_stage_4__543_, data_stage_4__542_, data_stage_4__541_, data_stage_4__540_, data_stage_4__539_, data_stage_4__538_, data_stage_4__537_, data_stage_4__536_, data_stage_4__535_, data_stage_4__534_, data_stage_4__533_, data_stage_4__532_, data_stage_4__531_, data_stage_4__530_, data_stage_4__529_, data_stage_4__528_, data_stage_4__527_, data_stage_4__526_, data_stage_4__525_, data_stage_4__524_, data_stage_4__523_, data_stage_4__522_, data_stage_4__521_, data_stage_4__520_, data_stage_4__519_, data_stage_4__518_, data_stage_4__517_, data_stage_4__516_, data_stage_4__515_, data_stage_4__514_, data_stage_4__513_, data_stage_4__512_, data_stage_4__511_, data_stage_4__510_, data_stage_4__509_, data_stage_4__508_, data_stage_4__507_, data_stage_4__506_, data_stage_4__505_, data_stage_4__504_, data_stage_4__503_, data_stage_4__502_, data_stage_4__501_, data_stage_4__500_, data_stage_4__499_, data_stage_4__498_, data_stage_4__497_, data_stage_4__496_, data_stage_4__495_, data_stage_4__494_, data_stage_4__493_, data_stage_4__492_, data_stage_4__491_, data_stage_4__490_, data_stage_4__489_, data_stage_4__488_, data_stage_4__487_, data_stage_4__486_, data_stage_4__485_, data_stage_4__484_, data_stage_4__483_, data_stage_4__482_, data_stage_4__481_, data_stage_4__480_, data_stage_4__479_, data_stage_4__478_, data_stage_4__477_, data_stage_4__476_, data_stage_4__475_, data_stage_4__474_, data_stage_4__473_, data_stage_4__472_, data_stage_4__471_, data_stage_4__470_, data_stage_4__469_, data_stage_4__468_, data_stage_4__467_, data_stage_4__466_, data_stage_4__465_, data_stage_4__464_, data_stage_4__463_, data_stage_4__462_, data_stage_4__461_, data_stage_4__460_, data_stage_4__459_, data_stage_4__458_, data_stage_4__457_, data_stage_4__456_, data_stage_4__455_, data_stage_4__454_, data_stage_4__453_, data_stage_4__452_, data_stage_4__451_, data_stage_4__450_, data_stage_4__449_, data_stage_4__448_, data_stage_4__447_, data_stage_4__446_, data_stage_4__445_, data_stage_4__444_, data_stage_4__443_, data_stage_4__442_, data_stage_4__441_, data_stage_4__440_, data_stage_4__439_, data_stage_4__438_, data_stage_4__437_, data_stage_4__436_, data_stage_4__435_, data_stage_4__434_, data_stage_4__433_, data_stage_4__432_, data_stage_4__431_, data_stage_4__430_, data_stage_4__429_, data_stage_4__428_, data_stage_4__427_, data_stage_4__426_, data_stage_4__425_, data_stage_4__424_, data_stage_4__423_, data_stage_4__422_, data_stage_4__421_, data_stage_4__420_, data_stage_4__419_, data_stage_4__418_, data_stage_4__417_, data_stage_4__416_, data_stage_4__415_, data_stage_4__414_, data_stage_4__413_, data_stage_4__412_, data_stage_4__411_, data_stage_4__410_, data_stage_4__409_, data_stage_4__408_, data_stage_4__407_, data_stage_4__406_, data_stage_4__405_, data_stage_4__404_, data_stage_4__403_, data_stage_4__402_, data_stage_4__401_, data_stage_4__400_, data_stage_4__399_, data_stage_4__398_, data_stage_4__397_, data_stage_4__396_, data_stage_4__395_, data_stage_4__394_, data_stage_4__393_, data_stage_4__392_, data_stage_4__391_, data_stage_4__390_, data_stage_4__389_, data_stage_4__388_, data_stage_4__387_, data_stage_4__386_, data_stage_4__385_, data_stage_4__384_, data_stage_4__383_, data_stage_4__382_, data_stage_4__381_, data_stage_4__380_, data_stage_4__379_, data_stage_4__378_, data_stage_4__377_, data_stage_4__376_, data_stage_4__375_, data_stage_4__374_, data_stage_4__373_, data_stage_4__372_, data_stage_4__371_, data_stage_4__370_, data_stage_4__369_, data_stage_4__368_, data_stage_4__367_, data_stage_4__366_, data_stage_4__365_, data_stage_4__364_, data_stage_4__363_, data_stage_4__362_, data_stage_4__361_, data_stage_4__360_, data_stage_4__359_, data_stage_4__358_, data_stage_4__357_, data_stage_4__356_, data_stage_4__355_, data_stage_4__354_, data_stage_4__353_, data_stage_4__352_, data_stage_4__351_, data_stage_4__350_, data_stage_4__349_, data_stage_4__348_, data_stage_4__347_, data_stage_4__346_, data_stage_4__345_, data_stage_4__344_, data_stage_4__343_, data_stage_4__342_, data_stage_4__341_, data_stage_4__340_, data_stage_4__339_, data_stage_4__338_, data_stage_4__337_, data_stage_4__336_, data_stage_4__335_, data_stage_4__334_, data_stage_4__333_, data_stage_4__332_, data_stage_4__331_, data_stage_4__330_, data_stage_4__329_, data_stage_4__328_, data_stage_4__327_, data_stage_4__326_, data_stage_4__325_, data_stage_4__324_, data_stage_4__323_, data_stage_4__322_, data_stage_4__321_, data_stage_4__320_, data_stage_4__319_, data_stage_4__318_, data_stage_4__317_, data_stage_4__316_, data_stage_4__315_, data_stage_4__314_, data_stage_4__313_, data_stage_4__312_, data_stage_4__311_, data_stage_4__310_, data_stage_4__309_, data_stage_4__308_, data_stage_4__307_, data_stage_4__306_, data_stage_4__305_, data_stage_4__304_, data_stage_4__303_, data_stage_4__302_, data_stage_4__301_, data_stage_4__300_, data_stage_4__299_, data_stage_4__298_, data_stage_4__297_, data_stage_4__296_, data_stage_4__295_, data_stage_4__294_, data_stage_4__293_, data_stage_4__292_, data_stage_4__291_, data_stage_4__290_, data_stage_4__289_, data_stage_4__288_, data_stage_4__287_, data_stage_4__286_, data_stage_4__285_, data_stage_4__284_, data_stage_4__283_, data_stage_4__282_, data_stage_4__281_, data_stage_4__280_, data_stage_4__279_, data_stage_4__278_, data_stage_4__277_, data_stage_4__276_, data_stage_4__275_, data_stage_4__274_, data_stage_4__273_, data_stage_4__272_, data_stage_4__271_, data_stage_4__270_, data_stage_4__269_, data_stage_4__268_, data_stage_4__267_, data_stage_4__266_, data_stage_4__265_, data_stage_4__264_, data_stage_4__263_, data_stage_4__262_, data_stage_4__261_, data_stage_4__260_, data_stage_4__259_, data_stage_4__258_, data_stage_4__257_, data_stage_4__256_, data_stage_4__255_, data_stage_4__254_, data_stage_4__253_, data_stage_4__252_, data_stage_4__251_, data_stage_4__250_, data_stage_4__249_, data_stage_4__248_, data_stage_4__247_, data_stage_4__246_, data_stage_4__245_, data_stage_4__244_, data_stage_4__243_, data_stage_4__242_, data_stage_4__241_, data_stage_4__240_, data_stage_4__239_, data_stage_4__238_, data_stage_4__237_, data_stage_4__236_, data_stage_4__235_, data_stage_4__234_, data_stage_4__233_, data_stage_4__232_, data_stage_4__231_, data_stage_4__230_, data_stage_4__229_, data_stage_4__228_, data_stage_4__227_, data_stage_4__226_, data_stage_4__225_, data_stage_4__224_, data_stage_4__223_, data_stage_4__222_, data_stage_4__221_, data_stage_4__220_, data_stage_4__219_, data_stage_4__218_, data_stage_4__217_, data_stage_4__216_, data_stage_4__215_, data_stage_4__214_, data_stage_4__213_, data_stage_4__212_, data_stage_4__211_, data_stage_4__210_, data_stage_4__209_, data_stage_4__208_, data_stage_4__207_, data_stage_4__206_, data_stage_4__205_, data_stage_4__204_, data_stage_4__203_, data_stage_4__202_, data_stage_4__201_, data_stage_4__200_, data_stage_4__199_, data_stage_4__198_, data_stage_4__197_, data_stage_4__196_, data_stage_4__195_, data_stage_4__194_, data_stage_4__193_, data_stage_4__192_, data_stage_4__191_, data_stage_4__190_, data_stage_4__189_, data_stage_4__188_, data_stage_4__187_, data_stage_4__186_, data_stage_4__185_, data_stage_4__184_, data_stage_4__183_, data_stage_4__182_, data_stage_4__181_, data_stage_4__180_, data_stage_4__179_, data_stage_4__178_, data_stage_4__177_, data_stage_4__176_, data_stage_4__175_, data_stage_4__174_, data_stage_4__173_, data_stage_4__172_, data_stage_4__171_, data_stage_4__170_, data_stage_4__169_, data_stage_4__168_, data_stage_4__167_, data_stage_4__166_, data_stage_4__165_, data_stage_4__164_, data_stage_4__163_, data_stage_4__162_, data_stage_4__161_, data_stage_4__160_, data_stage_4__159_, data_stage_4__158_, data_stage_4__157_, data_stage_4__156_, data_stage_4__155_, data_stage_4__154_, data_stage_4__153_, data_stage_4__152_, data_stage_4__151_, data_stage_4__150_, data_stage_4__149_, data_stage_4__148_, data_stage_4__147_, data_stage_4__146_, data_stage_4__145_, data_stage_4__144_, data_stage_4__143_, data_stage_4__142_, data_stage_4__141_, data_stage_4__140_, data_stage_4__139_, data_stage_4__138_, data_stage_4__137_, data_stage_4__136_, data_stage_4__135_, data_stage_4__134_, data_stage_4__133_, data_stage_4__132_, data_stage_4__131_, data_stage_4__130_, data_stage_4__129_, data_stage_4__128_, data_stage_4__127_, data_stage_4__126_, data_stage_4__125_, data_stage_4__124_, data_stage_4__123_, data_stage_4__122_, data_stage_4__121_, data_stage_4__120_, data_stage_4__119_, data_stage_4__118_, data_stage_4__117_, data_stage_4__116_, data_stage_4__115_, data_stage_4__114_, data_stage_4__113_, data_stage_4__112_, data_stage_4__111_, data_stage_4__110_, data_stage_4__109_, data_stage_4__108_, data_stage_4__107_, data_stage_4__106_, data_stage_4__105_, data_stage_4__104_, data_stage_4__103_, data_stage_4__102_, data_stage_4__101_, data_stage_4__100_, data_stage_4__99_, data_stage_4__98_, data_stage_4__97_, data_stage_4__96_, data_stage_4__95_, data_stage_4__94_, data_stage_4__93_, data_stage_4__92_, data_stage_4__91_, data_stage_4__90_, data_stage_4__89_, data_stage_4__88_, data_stage_4__87_, data_stage_4__86_, data_stage_4__85_, data_stage_4__84_, data_stage_4__83_, data_stage_4__82_, data_stage_4__81_, data_stage_4__80_, data_stage_4__79_, data_stage_4__78_, data_stage_4__77_, data_stage_4__76_, data_stage_4__75_, data_stage_4__74_, data_stage_4__73_, data_stage_4__72_, data_stage_4__71_, data_stage_4__70_, data_stage_4__69_, data_stage_4__68_, data_stage_4__67_, data_stage_4__66_, data_stage_4__65_, data_stage_4__64_, data_stage_4__63_, data_stage_4__62_, data_stage_4__61_, data_stage_4__60_, data_stage_4__59_, data_stage_4__58_, data_stage_4__57_, data_stage_4__56_, data_stage_4__55_, data_stage_4__54_, data_stage_4__53_, data_stage_4__52_, data_stage_4__51_, data_stage_4__50_, data_stage_4__49_, data_stage_4__48_, data_stage_4__47_, data_stage_4__46_, data_stage_4__45_, data_stage_4__44_, data_stage_4__43_, data_stage_4__42_, data_stage_4__41_, data_stage_4__40_, data_stage_4__39_, data_stage_4__38_, data_stage_4__37_, data_stage_4__36_, data_stage_4__35_, data_stage_4__34_, data_stage_4__33_, data_stage_4__32_, data_stage_4__31_, data_stage_4__30_, data_stage_4__29_, data_stage_4__28_, data_stage_4__27_, data_stage_4__26_, data_stage_4__25_, data_stage_4__24_, data_stage_4__23_, data_stage_4__22_, data_stage_4__21_, data_stage_4__20_, data_stage_4__19_, data_stage_4__18_, data_stage_4__17_, data_stage_4__16_, data_stage_4__15_, data_stage_4__14_, data_stage_4__13_, data_stage_4__12_, data_stage_4__11_, data_stage_4__10_, data_stage_4__9_, data_stage_4__8_, data_stage_4__7_, data_stage_4__6_, data_stage_4__5_, data_stage_4__4_, data_stage_4__3_, data_stage_4__2_, data_stage_4__1_, data_stage_4__0_ })
  );


  bsg_swap_width_p1024
  mux_stage_3__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_3__4095_, data_stage_3__4094_, data_stage_3__4093_, data_stage_3__4092_, data_stage_3__4091_, data_stage_3__4090_, data_stage_3__4089_, data_stage_3__4088_, data_stage_3__4087_, data_stage_3__4086_, data_stage_3__4085_, data_stage_3__4084_, data_stage_3__4083_, data_stage_3__4082_, data_stage_3__4081_, data_stage_3__4080_, data_stage_3__4079_, data_stage_3__4078_, data_stage_3__4077_, data_stage_3__4076_, data_stage_3__4075_, data_stage_3__4074_, data_stage_3__4073_, data_stage_3__4072_, data_stage_3__4071_, data_stage_3__4070_, data_stage_3__4069_, data_stage_3__4068_, data_stage_3__4067_, data_stage_3__4066_, data_stage_3__4065_, data_stage_3__4064_, data_stage_3__4063_, data_stage_3__4062_, data_stage_3__4061_, data_stage_3__4060_, data_stage_3__4059_, data_stage_3__4058_, data_stage_3__4057_, data_stage_3__4056_, data_stage_3__4055_, data_stage_3__4054_, data_stage_3__4053_, data_stage_3__4052_, data_stage_3__4051_, data_stage_3__4050_, data_stage_3__4049_, data_stage_3__4048_, data_stage_3__4047_, data_stage_3__4046_, data_stage_3__4045_, data_stage_3__4044_, data_stage_3__4043_, data_stage_3__4042_, data_stage_3__4041_, data_stage_3__4040_, data_stage_3__4039_, data_stage_3__4038_, data_stage_3__4037_, data_stage_3__4036_, data_stage_3__4035_, data_stage_3__4034_, data_stage_3__4033_, data_stage_3__4032_, data_stage_3__4031_, data_stage_3__4030_, data_stage_3__4029_, data_stage_3__4028_, data_stage_3__4027_, data_stage_3__4026_, data_stage_3__4025_, data_stage_3__4024_, data_stage_3__4023_, data_stage_3__4022_, data_stage_3__4021_, data_stage_3__4020_, data_stage_3__4019_, data_stage_3__4018_, data_stage_3__4017_, data_stage_3__4016_, data_stage_3__4015_, data_stage_3__4014_, data_stage_3__4013_, data_stage_3__4012_, data_stage_3__4011_, data_stage_3__4010_, data_stage_3__4009_, data_stage_3__4008_, data_stage_3__4007_, data_stage_3__4006_, data_stage_3__4005_, data_stage_3__4004_, data_stage_3__4003_, data_stage_3__4002_, data_stage_3__4001_, data_stage_3__4000_, data_stage_3__3999_, data_stage_3__3998_, data_stage_3__3997_, data_stage_3__3996_, data_stage_3__3995_, data_stage_3__3994_, data_stage_3__3993_, data_stage_3__3992_, data_stage_3__3991_, data_stage_3__3990_, data_stage_3__3989_, data_stage_3__3988_, data_stage_3__3987_, data_stage_3__3986_, data_stage_3__3985_, data_stage_3__3984_, data_stage_3__3983_, data_stage_3__3982_, data_stage_3__3981_, data_stage_3__3980_, data_stage_3__3979_, data_stage_3__3978_, data_stage_3__3977_, data_stage_3__3976_, data_stage_3__3975_, data_stage_3__3974_, data_stage_3__3973_, data_stage_3__3972_, data_stage_3__3971_, data_stage_3__3970_, data_stage_3__3969_, data_stage_3__3968_, data_stage_3__3967_, data_stage_3__3966_, data_stage_3__3965_, data_stage_3__3964_, data_stage_3__3963_, data_stage_3__3962_, data_stage_3__3961_, data_stage_3__3960_, data_stage_3__3959_, data_stage_3__3958_, data_stage_3__3957_, data_stage_3__3956_, data_stage_3__3955_, data_stage_3__3954_, data_stage_3__3953_, data_stage_3__3952_, data_stage_3__3951_, data_stage_3__3950_, data_stage_3__3949_, data_stage_3__3948_, data_stage_3__3947_, data_stage_3__3946_, data_stage_3__3945_, data_stage_3__3944_, data_stage_3__3943_, data_stage_3__3942_, data_stage_3__3941_, data_stage_3__3940_, data_stage_3__3939_, data_stage_3__3938_, data_stage_3__3937_, data_stage_3__3936_, data_stage_3__3935_, data_stage_3__3934_, data_stage_3__3933_, data_stage_3__3932_, data_stage_3__3931_, data_stage_3__3930_, data_stage_3__3929_, data_stage_3__3928_, data_stage_3__3927_, data_stage_3__3926_, data_stage_3__3925_, data_stage_3__3924_, data_stage_3__3923_, data_stage_3__3922_, data_stage_3__3921_, data_stage_3__3920_, data_stage_3__3919_, data_stage_3__3918_, data_stage_3__3917_, data_stage_3__3916_, data_stage_3__3915_, data_stage_3__3914_, data_stage_3__3913_, data_stage_3__3912_, data_stage_3__3911_, data_stage_3__3910_, data_stage_3__3909_, data_stage_3__3908_, data_stage_3__3907_, data_stage_3__3906_, data_stage_3__3905_, data_stage_3__3904_, data_stage_3__3903_, data_stage_3__3902_, data_stage_3__3901_, data_stage_3__3900_, data_stage_3__3899_, data_stage_3__3898_, data_stage_3__3897_, data_stage_3__3896_, data_stage_3__3895_, data_stage_3__3894_, data_stage_3__3893_, data_stage_3__3892_, data_stage_3__3891_, data_stage_3__3890_, data_stage_3__3889_, data_stage_3__3888_, data_stage_3__3887_, data_stage_3__3886_, data_stage_3__3885_, data_stage_3__3884_, data_stage_3__3883_, data_stage_3__3882_, data_stage_3__3881_, data_stage_3__3880_, data_stage_3__3879_, data_stage_3__3878_, data_stage_3__3877_, data_stage_3__3876_, data_stage_3__3875_, data_stage_3__3874_, data_stage_3__3873_, data_stage_3__3872_, data_stage_3__3871_, data_stage_3__3870_, data_stage_3__3869_, data_stage_3__3868_, data_stage_3__3867_, data_stage_3__3866_, data_stage_3__3865_, data_stage_3__3864_, data_stage_3__3863_, data_stage_3__3862_, data_stage_3__3861_, data_stage_3__3860_, data_stage_3__3859_, data_stage_3__3858_, data_stage_3__3857_, data_stage_3__3856_, data_stage_3__3855_, data_stage_3__3854_, data_stage_3__3853_, data_stage_3__3852_, data_stage_3__3851_, data_stage_3__3850_, data_stage_3__3849_, data_stage_3__3848_, data_stage_3__3847_, data_stage_3__3846_, data_stage_3__3845_, data_stage_3__3844_, data_stage_3__3843_, data_stage_3__3842_, data_stage_3__3841_, data_stage_3__3840_, data_stage_3__3839_, data_stage_3__3838_, data_stage_3__3837_, data_stage_3__3836_, data_stage_3__3835_, data_stage_3__3834_, data_stage_3__3833_, data_stage_3__3832_, data_stage_3__3831_, data_stage_3__3830_, data_stage_3__3829_, data_stage_3__3828_, data_stage_3__3827_, data_stage_3__3826_, data_stage_3__3825_, data_stage_3__3824_, data_stage_3__3823_, data_stage_3__3822_, data_stage_3__3821_, data_stage_3__3820_, data_stage_3__3819_, data_stage_3__3818_, data_stage_3__3817_, data_stage_3__3816_, data_stage_3__3815_, data_stage_3__3814_, data_stage_3__3813_, data_stage_3__3812_, data_stage_3__3811_, data_stage_3__3810_, data_stage_3__3809_, data_stage_3__3808_, data_stage_3__3807_, data_stage_3__3806_, data_stage_3__3805_, data_stage_3__3804_, data_stage_3__3803_, data_stage_3__3802_, data_stage_3__3801_, data_stage_3__3800_, data_stage_3__3799_, data_stage_3__3798_, data_stage_3__3797_, data_stage_3__3796_, data_stage_3__3795_, data_stage_3__3794_, data_stage_3__3793_, data_stage_3__3792_, data_stage_3__3791_, data_stage_3__3790_, data_stage_3__3789_, data_stage_3__3788_, data_stage_3__3787_, data_stage_3__3786_, data_stage_3__3785_, data_stage_3__3784_, data_stage_3__3783_, data_stage_3__3782_, data_stage_3__3781_, data_stage_3__3780_, data_stage_3__3779_, data_stage_3__3778_, data_stage_3__3777_, data_stage_3__3776_, data_stage_3__3775_, data_stage_3__3774_, data_stage_3__3773_, data_stage_3__3772_, data_stage_3__3771_, data_stage_3__3770_, data_stage_3__3769_, data_stage_3__3768_, data_stage_3__3767_, data_stage_3__3766_, data_stage_3__3765_, data_stage_3__3764_, data_stage_3__3763_, data_stage_3__3762_, data_stage_3__3761_, data_stage_3__3760_, data_stage_3__3759_, data_stage_3__3758_, data_stage_3__3757_, data_stage_3__3756_, data_stage_3__3755_, data_stage_3__3754_, data_stage_3__3753_, data_stage_3__3752_, data_stage_3__3751_, data_stage_3__3750_, data_stage_3__3749_, data_stage_3__3748_, data_stage_3__3747_, data_stage_3__3746_, data_stage_3__3745_, data_stage_3__3744_, data_stage_3__3743_, data_stage_3__3742_, data_stage_3__3741_, data_stage_3__3740_, data_stage_3__3739_, data_stage_3__3738_, data_stage_3__3737_, data_stage_3__3736_, data_stage_3__3735_, data_stage_3__3734_, data_stage_3__3733_, data_stage_3__3732_, data_stage_3__3731_, data_stage_3__3730_, data_stage_3__3729_, data_stage_3__3728_, data_stage_3__3727_, data_stage_3__3726_, data_stage_3__3725_, data_stage_3__3724_, data_stage_3__3723_, data_stage_3__3722_, data_stage_3__3721_, data_stage_3__3720_, data_stage_3__3719_, data_stage_3__3718_, data_stage_3__3717_, data_stage_3__3716_, data_stage_3__3715_, data_stage_3__3714_, data_stage_3__3713_, data_stage_3__3712_, data_stage_3__3711_, data_stage_3__3710_, data_stage_3__3709_, data_stage_3__3708_, data_stage_3__3707_, data_stage_3__3706_, data_stage_3__3705_, data_stage_3__3704_, data_stage_3__3703_, data_stage_3__3702_, data_stage_3__3701_, data_stage_3__3700_, data_stage_3__3699_, data_stage_3__3698_, data_stage_3__3697_, data_stage_3__3696_, data_stage_3__3695_, data_stage_3__3694_, data_stage_3__3693_, data_stage_3__3692_, data_stage_3__3691_, data_stage_3__3690_, data_stage_3__3689_, data_stage_3__3688_, data_stage_3__3687_, data_stage_3__3686_, data_stage_3__3685_, data_stage_3__3684_, data_stage_3__3683_, data_stage_3__3682_, data_stage_3__3681_, data_stage_3__3680_, data_stage_3__3679_, data_stage_3__3678_, data_stage_3__3677_, data_stage_3__3676_, data_stage_3__3675_, data_stage_3__3674_, data_stage_3__3673_, data_stage_3__3672_, data_stage_3__3671_, data_stage_3__3670_, data_stage_3__3669_, data_stage_3__3668_, data_stage_3__3667_, data_stage_3__3666_, data_stage_3__3665_, data_stage_3__3664_, data_stage_3__3663_, data_stage_3__3662_, data_stage_3__3661_, data_stage_3__3660_, data_stage_3__3659_, data_stage_3__3658_, data_stage_3__3657_, data_stage_3__3656_, data_stage_3__3655_, data_stage_3__3654_, data_stage_3__3653_, data_stage_3__3652_, data_stage_3__3651_, data_stage_3__3650_, data_stage_3__3649_, data_stage_3__3648_, data_stage_3__3647_, data_stage_3__3646_, data_stage_3__3645_, data_stage_3__3644_, data_stage_3__3643_, data_stage_3__3642_, data_stage_3__3641_, data_stage_3__3640_, data_stage_3__3639_, data_stage_3__3638_, data_stage_3__3637_, data_stage_3__3636_, data_stage_3__3635_, data_stage_3__3634_, data_stage_3__3633_, data_stage_3__3632_, data_stage_3__3631_, data_stage_3__3630_, data_stage_3__3629_, data_stage_3__3628_, data_stage_3__3627_, data_stage_3__3626_, data_stage_3__3625_, data_stage_3__3624_, data_stage_3__3623_, data_stage_3__3622_, data_stage_3__3621_, data_stage_3__3620_, data_stage_3__3619_, data_stage_3__3618_, data_stage_3__3617_, data_stage_3__3616_, data_stage_3__3615_, data_stage_3__3614_, data_stage_3__3613_, data_stage_3__3612_, data_stage_3__3611_, data_stage_3__3610_, data_stage_3__3609_, data_stage_3__3608_, data_stage_3__3607_, data_stage_3__3606_, data_stage_3__3605_, data_stage_3__3604_, data_stage_3__3603_, data_stage_3__3602_, data_stage_3__3601_, data_stage_3__3600_, data_stage_3__3599_, data_stage_3__3598_, data_stage_3__3597_, data_stage_3__3596_, data_stage_3__3595_, data_stage_3__3594_, data_stage_3__3593_, data_stage_3__3592_, data_stage_3__3591_, data_stage_3__3590_, data_stage_3__3589_, data_stage_3__3588_, data_stage_3__3587_, data_stage_3__3586_, data_stage_3__3585_, data_stage_3__3584_, data_stage_3__3583_, data_stage_3__3582_, data_stage_3__3581_, data_stage_3__3580_, data_stage_3__3579_, data_stage_3__3578_, data_stage_3__3577_, data_stage_3__3576_, data_stage_3__3575_, data_stage_3__3574_, data_stage_3__3573_, data_stage_3__3572_, data_stage_3__3571_, data_stage_3__3570_, data_stage_3__3569_, data_stage_3__3568_, data_stage_3__3567_, data_stage_3__3566_, data_stage_3__3565_, data_stage_3__3564_, data_stage_3__3563_, data_stage_3__3562_, data_stage_3__3561_, data_stage_3__3560_, data_stage_3__3559_, data_stage_3__3558_, data_stage_3__3557_, data_stage_3__3556_, data_stage_3__3555_, data_stage_3__3554_, data_stage_3__3553_, data_stage_3__3552_, data_stage_3__3551_, data_stage_3__3550_, data_stage_3__3549_, data_stage_3__3548_, data_stage_3__3547_, data_stage_3__3546_, data_stage_3__3545_, data_stage_3__3544_, data_stage_3__3543_, data_stage_3__3542_, data_stage_3__3541_, data_stage_3__3540_, data_stage_3__3539_, data_stage_3__3538_, data_stage_3__3537_, data_stage_3__3536_, data_stage_3__3535_, data_stage_3__3534_, data_stage_3__3533_, data_stage_3__3532_, data_stage_3__3531_, data_stage_3__3530_, data_stage_3__3529_, data_stage_3__3528_, data_stage_3__3527_, data_stage_3__3526_, data_stage_3__3525_, data_stage_3__3524_, data_stage_3__3523_, data_stage_3__3522_, data_stage_3__3521_, data_stage_3__3520_, data_stage_3__3519_, data_stage_3__3518_, data_stage_3__3517_, data_stage_3__3516_, data_stage_3__3515_, data_stage_3__3514_, data_stage_3__3513_, data_stage_3__3512_, data_stage_3__3511_, data_stage_3__3510_, data_stage_3__3509_, data_stage_3__3508_, data_stage_3__3507_, data_stage_3__3506_, data_stage_3__3505_, data_stage_3__3504_, data_stage_3__3503_, data_stage_3__3502_, data_stage_3__3501_, data_stage_3__3500_, data_stage_3__3499_, data_stage_3__3498_, data_stage_3__3497_, data_stage_3__3496_, data_stage_3__3495_, data_stage_3__3494_, data_stage_3__3493_, data_stage_3__3492_, data_stage_3__3491_, data_stage_3__3490_, data_stage_3__3489_, data_stage_3__3488_, data_stage_3__3487_, data_stage_3__3486_, data_stage_3__3485_, data_stage_3__3484_, data_stage_3__3483_, data_stage_3__3482_, data_stage_3__3481_, data_stage_3__3480_, data_stage_3__3479_, data_stage_3__3478_, data_stage_3__3477_, data_stage_3__3476_, data_stage_3__3475_, data_stage_3__3474_, data_stage_3__3473_, data_stage_3__3472_, data_stage_3__3471_, data_stage_3__3470_, data_stage_3__3469_, data_stage_3__3468_, data_stage_3__3467_, data_stage_3__3466_, data_stage_3__3465_, data_stage_3__3464_, data_stage_3__3463_, data_stage_3__3462_, data_stage_3__3461_, data_stage_3__3460_, data_stage_3__3459_, data_stage_3__3458_, data_stage_3__3457_, data_stage_3__3456_, data_stage_3__3455_, data_stage_3__3454_, data_stage_3__3453_, data_stage_3__3452_, data_stage_3__3451_, data_stage_3__3450_, data_stage_3__3449_, data_stage_3__3448_, data_stage_3__3447_, data_stage_3__3446_, data_stage_3__3445_, data_stage_3__3444_, data_stage_3__3443_, data_stage_3__3442_, data_stage_3__3441_, data_stage_3__3440_, data_stage_3__3439_, data_stage_3__3438_, data_stage_3__3437_, data_stage_3__3436_, data_stage_3__3435_, data_stage_3__3434_, data_stage_3__3433_, data_stage_3__3432_, data_stage_3__3431_, data_stage_3__3430_, data_stage_3__3429_, data_stage_3__3428_, data_stage_3__3427_, data_stage_3__3426_, data_stage_3__3425_, data_stage_3__3424_, data_stage_3__3423_, data_stage_3__3422_, data_stage_3__3421_, data_stage_3__3420_, data_stage_3__3419_, data_stage_3__3418_, data_stage_3__3417_, data_stage_3__3416_, data_stage_3__3415_, data_stage_3__3414_, data_stage_3__3413_, data_stage_3__3412_, data_stage_3__3411_, data_stage_3__3410_, data_stage_3__3409_, data_stage_3__3408_, data_stage_3__3407_, data_stage_3__3406_, data_stage_3__3405_, data_stage_3__3404_, data_stage_3__3403_, data_stage_3__3402_, data_stage_3__3401_, data_stage_3__3400_, data_stage_3__3399_, data_stage_3__3398_, data_stage_3__3397_, data_stage_3__3396_, data_stage_3__3395_, data_stage_3__3394_, data_stage_3__3393_, data_stage_3__3392_, data_stage_3__3391_, data_stage_3__3390_, data_stage_3__3389_, data_stage_3__3388_, data_stage_3__3387_, data_stage_3__3386_, data_stage_3__3385_, data_stage_3__3384_, data_stage_3__3383_, data_stage_3__3382_, data_stage_3__3381_, data_stage_3__3380_, data_stage_3__3379_, data_stage_3__3378_, data_stage_3__3377_, data_stage_3__3376_, data_stage_3__3375_, data_stage_3__3374_, data_stage_3__3373_, data_stage_3__3372_, data_stage_3__3371_, data_stage_3__3370_, data_stage_3__3369_, data_stage_3__3368_, data_stage_3__3367_, data_stage_3__3366_, data_stage_3__3365_, data_stage_3__3364_, data_stage_3__3363_, data_stage_3__3362_, data_stage_3__3361_, data_stage_3__3360_, data_stage_3__3359_, data_stage_3__3358_, data_stage_3__3357_, data_stage_3__3356_, data_stage_3__3355_, data_stage_3__3354_, data_stage_3__3353_, data_stage_3__3352_, data_stage_3__3351_, data_stage_3__3350_, data_stage_3__3349_, data_stage_3__3348_, data_stage_3__3347_, data_stage_3__3346_, data_stage_3__3345_, data_stage_3__3344_, data_stage_3__3343_, data_stage_3__3342_, data_stage_3__3341_, data_stage_3__3340_, data_stage_3__3339_, data_stage_3__3338_, data_stage_3__3337_, data_stage_3__3336_, data_stage_3__3335_, data_stage_3__3334_, data_stage_3__3333_, data_stage_3__3332_, data_stage_3__3331_, data_stage_3__3330_, data_stage_3__3329_, data_stage_3__3328_, data_stage_3__3327_, data_stage_3__3326_, data_stage_3__3325_, data_stage_3__3324_, data_stage_3__3323_, data_stage_3__3322_, data_stage_3__3321_, data_stage_3__3320_, data_stage_3__3319_, data_stage_3__3318_, data_stage_3__3317_, data_stage_3__3316_, data_stage_3__3315_, data_stage_3__3314_, data_stage_3__3313_, data_stage_3__3312_, data_stage_3__3311_, data_stage_3__3310_, data_stage_3__3309_, data_stage_3__3308_, data_stage_3__3307_, data_stage_3__3306_, data_stage_3__3305_, data_stage_3__3304_, data_stage_3__3303_, data_stage_3__3302_, data_stage_3__3301_, data_stage_3__3300_, data_stage_3__3299_, data_stage_3__3298_, data_stage_3__3297_, data_stage_3__3296_, data_stage_3__3295_, data_stage_3__3294_, data_stage_3__3293_, data_stage_3__3292_, data_stage_3__3291_, data_stage_3__3290_, data_stage_3__3289_, data_stage_3__3288_, data_stage_3__3287_, data_stage_3__3286_, data_stage_3__3285_, data_stage_3__3284_, data_stage_3__3283_, data_stage_3__3282_, data_stage_3__3281_, data_stage_3__3280_, data_stage_3__3279_, data_stage_3__3278_, data_stage_3__3277_, data_stage_3__3276_, data_stage_3__3275_, data_stage_3__3274_, data_stage_3__3273_, data_stage_3__3272_, data_stage_3__3271_, data_stage_3__3270_, data_stage_3__3269_, data_stage_3__3268_, data_stage_3__3267_, data_stage_3__3266_, data_stage_3__3265_, data_stage_3__3264_, data_stage_3__3263_, data_stage_3__3262_, data_stage_3__3261_, data_stage_3__3260_, data_stage_3__3259_, data_stage_3__3258_, data_stage_3__3257_, data_stage_3__3256_, data_stage_3__3255_, data_stage_3__3254_, data_stage_3__3253_, data_stage_3__3252_, data_stage_3__3251_, data_stage_3__3250_, data_stage_3__3249_, data_stage_3__3248_, data_stage_3__3247_, data_stage_3__3246_, data_stage_3__3245_, data_stage_3__3244_, data_stage_3__3243_, data_stage_3__3242_, data_stage_3__3241_, data_stage_3__3240_, data_stage_3__3239_, data_stage_3__3238_, data_stage_3__3237_, data_stage_3__3236_, data_stage_3__3235_, data_stage_3__3234_, data_stage_3__3233_, data_stage_3__3232_, data_stage_3__3231_, data_stage_3__3230_, data_stage_3__3229_, data_stage_3__3228_, data_stage_3__3227_, data_stage_3__3226_, data_stage_3__3225_, data_stage_3__3224_, data_stage_3__3223_, data_stage_3__3222_, data_stage_3__3221_, data_stage_3__3220_, data_stage_3__3219_, data_stage_3__3218_, data_stage_3__3217_, data_stage_3__3216_, data_stage_3__3215_, data_stage_3__3214_, data_stage_3__3213_, data_stage_3__3212_, data_stage_3__3211_, data_stage_3__3210_, data_stage_3__3209_, data_stage_3__3208_, data_stage_3__3207_, data_stage_3__3206_, data_stage_3__3205_, data_stage_3__3204_, data_stage_3__3203_, data_stage_3__3202_, data_stage_3__3201_, data_stage_3__3200_, data_stage_3__3199_, data_stage_3__3198_, data_stage_3__3197_, data_stage_3__3196_, data_stage_3__3195_, data_stage_3__3194_, data_stage_3__3193_, data_stage_3__3192_, data_stage_3__3191_, data_stage_3__3190_, data_stage_3__3189_, data_stage_3__3188_, data_stage_3__3187_, data_stage_3__3186_, data_stage_3__3185_, data_stage_3__3184_, data_stage_3__3183_, data_stage_3__3182_, data_stage_3__3181_, data_stage_3__3180_, data_stage_3__3179_, data_stage_3__3178_, data_stage_3__3177_, data_stage_3__3176_, data_stage_3__3175_, data_stage_3__3174_, data_stage_3__3173_, data_stage_3__3172_, data_stage_3__3171_, data_stage_3__3170_, data_stage_3__3169_, data_stage_3__3168_, data_stage_3__3167_, data_stage_3__3166_, data_stage_3__3165_, data_stage_3__3164_, data_stage_3__3163_, data_stage_3__3162_, data_stage_3__3161_, data_stage_3__3160_, data_stage_3__3159_, data_stage_3__3158_, data_stage_3__3157_, data_stage_3__3156_, data_stage_3__3155_, data_stage_3__3154_, data_stage_3__3153_, data_stage_3__3152_, data_stage_3__3151_, data_stage_3__3150_, data_stage_3__3149_, data_stage_3__3148_, data_stage_3__3147_, data_stage_3__3146_, data_stage_3__3145_, data_stage_3__3144_, data_stage_3__3143_, data_stage_3__3142_, data_stage_3__3141_, data_stage_3__3140_, data_stage_3__3139_, data_stage_3__3138_, data_stage_3__3137_, data_stage_3__3136_, data_stage_3__3135_, data_stage_3__3134_, data_stage_3__3133_, data_stage_3__3132_, data_stage_3__3131_, data_stage_3__3130_, data_stage_3__3129_, data_stage_3__3128_, data_stage_3__3127_, data_stage_3__3126_, data_stage_3__3125_, data_stage_3__3124_, data_stage_3__3123_, data_stage_3__3122_, data_stage_3__3121_, data_stage_3__3120_, data_stage_3__3119_, data_stage_3__3118_, data_stage_3__3117_, data_stage_3__3116_, data_stage_3__3115_, data_stage_3__3114_, data_stage_3__3113_, data_stage_3__3112_, data_stage_3__3111_, data_stage_3__3110_, data_stage_3__3109_, data_stage_3__3108_, data_stage_3__3107_, data_stage_3__3106_, data_stage_3__3105_, data_stage_3__3104_, data_stage_3__3103_, data_stage_3__3102_, data_stage_3__3101_, data_stage_3__3100_, data_stage_3__3099_, data_stage_3__3098_, data_stage_3__3097_, data_stage_3__3096_, data_stage_3__3095_, data_stage_3__3094_, data_stage_3__3093_, data_stage_3__3092_, data_stage_3__3091_, data_stage_3__3090_, data_stage_3__3089_, data_stage_3__3088_, data_stage_3__3087_, data_stage_3__3086_, data_stage_3__3085_, data_stage_3__3084_, data_stage_3__3083_, data_stage_3__3082_, data_stage_3__3081_, data_stage_3__3080_, data_stage_3__3079_, data_stage_3__3078_, data_stage_3__3077_, data_stage_3__3076_, data_stage_3__3075_, data_stage_3__3074_, data_stage_3__3073_, data_stage_3__3072_, data_stage_3__3071_, data_stage_3__3070_, data_stage_3__3069_, data_stage_3__3068_, data_stage_3__3067_, data_stage_3__3066_, data_stage_3__3065_, data_stage_3__3064_, data_stage_3__3063_, data_stage_3__3062_, data_stage_3__3061_, data_stage_3__3060_, data_stage_3__3059_, data_stage_3__3058_, data_stage_3__3057_, data_stage_3__3056_, data_stage_3__3055_, data_stage_3__3054_, data_stage_3__3053_, data_stage_3__3052_, data_stage_3__3051_, data_stage_3__3050_, data_stage_3__3049_, data_stage_3__3048_, data_stage_3__3047_, data_stage_3__3046_, data_stage_3__3045_, data_stage_3__3044_, data_stage_3__3043_, data_stage_3__3042_, data_stage_3__3041_, data_stage_3__3040_, data_stage_3__3039_, data_stage_3__3038_, data_stage_3__3037_, data_stage_3__3036_, data_stage_3__3035_, data_stage_3__3034_, data_stage_3__3033_, data_stage_3__3032_, data_stage_3__3031_, data_stage_3__3030_, data_stage_3__3029_, data_stage_3__3028_, data_stage_3__3027_, data_stage_3__3026_, data_stage_3__3025_, data_stage_3__3024_, data_stage_3__3023_, data_stage_3__3022_, data_stage_3__3021_, data_stage_3__3020_, data_stage_3__3019_, data_stage_3__3018_, data_stage_3__3017_, data_stage_3__3016_, data_stage_3__3015_, data_stage_3__3014_, data_stage_3__3013_, data_stage_3__3012_, data_stage_3__3011_, data_stage_3__3010_, data_stage_3__3009_, data_stage_3__3008_, data_stage_3__3007_, data_stage_3__3006_, data_stage_3__3005_, data_stage_3__3004_, data_stage_3__3003_, data_stage_3__3002_, data_stage_3__3001_, data_stage_3__3000_, data_stage_3__2999_, data_stage_3__2998_, data_stage_3__2997_, data_stage_3__2996_, data_stage_3__2995_, data_stage_3__2994_, data_stage_3__2993_, data_stage_3__2992_, data_stage_3__2991_, data_stage_3__2990_, data_stage_3__2989_, data_stage_3__2988_, data_stage_3__2987_, data_stage_3__2986_, data_stage_3__2985_, data_stage_3__2984_, data_stage_3__2983_, data_stage_3__2982_, data_stage_3__2981_, data_stage_3__2980_, data_stage_3__2979_, data_stage_3__2978_, data_stage_3__2977_, data_stage_3__2976_, data_stage_3__2975_, data_stage_3__2974_, data_stage_3__2973_, data_stage_3__2972_, data_stage_3__2971_, data_stage_3__2970_, data_stage_3__2969_, data_stage_3__2968_, data_stage_3__2967_, data_stage_3__2966_, data_stage_3__2965_, data_stage_3__2964_, data_stage_3__2963_, data_stage_3__2962_, data_stage_3__2961_, data_stage_3__2960_, data_stage_3__2959_, data_stage_3__2958_, data_stage_3__2957_, data_stage_3__2956_, data_stage_3__2955_, data_stage_3__2954_, data_stage_3__2953_, data_stage_3__2952_, data_stage_3__2951_, data_stage_3__2950_, data_stage_3__2949_, data_stage_3__2948_, data_stage_3__2947_, data_stage_3__2946_, data_stage_3__2945_, data_stage_3__2944_, data_stage_3__2943_, data_stage_3__2942_, data_stage_3__2941_, data_stage_3__2940_, data_stage_3__2939_, data_stage_3__2938_, data_stage_3__2937_, data_stage_3__2936_, data_stage_3__2935_, data_stage_3__2934_, data_stage_3__2933_, data_stage_3__2932_, data_stage_3__2931_, data_stage_3__2930_, data_stage_3__2929_, data_stage_3__2928_, data_stage_3__2927_, data_stage_3__2926_, data_stage_3__2925_, data_stage_3__2924_, data_stage_3__2923_, data_stage_3__2922_, data_stage_3__2921_, data_stage_3__2920_, data_stage_3__2919_, data_stage_3__2918_, data_stage_3__2917_, data_stage_3__2916_, data_stage_3__2915_, data_stage_3__2914_, data_stage_3__2913_, data_stage_3__2912_, data_stage_3__2911_, data_stage_3__2910_, data_stage_3__2909_, data_stage_3__2908_, data_stage_3__2907_, data_stage_3__2906_, data_stage_3__2905_, data_stage_3__2904_, data_stage_3__2903_, data_stage_3__2902_, data_stage_3__2901_, data_stage_3__2900_, data_stage_3__2899_, data_stage_3__2898_, data_stage_3__2897_, data_stage_3__2896_, data_stage_3__2895_, data_stage_3__2894_, data_stage_3__2893_, data_stage_3__2892_, data_stage_3__2891_, data_stage_3__2890_, data_stage_3__2889_, data_stage_3__2888_, data_stage_3__2887_, data_stage_3__2886_, data_stage_3__2885_, data_stage_3__2884_, data_stage_3__2883_, data_stage_3__2882_, data_stage_3__2881_, data_stage_3__2880_, data_stage_3__2879_, data_stage_3__2878_, data_stage_3__2877_, data_stage_3__2876_, data_stage_3__2875_, data_stage_3__2874_, data_stage_3__2873_, data_stage_3__2872_, data_stage_3__2871_, data_stage_3__2870_, data_stage_3__2869_, data_stage_3__2868_, data_stage_3__2867_, data_stage_3__2866_, data_stage_3__2865_, data_stage_3__2864_, data_stage_3__2863_, data_stage_3__2862_, data_stage_3__2861_, data_stage_3__2860_, data_stage_3__2859_, data_stage_3__2858_, data_stage_3__2857_, data_stage_3__2856_, data_stage_3__2855_, data_stage_3__2854_, data_stage_3__2853_, data_stage_3__2852_, data_stage_3__2851_, data_stage_3__2850_, data_stage_3__2849_, data_stage_3__2848_, data_stage_3__2847_, data_stage_3__2846_, data_stage_3__2845_, data_stage_3__2844_, data_stage_3__2843_, data_stage_3__2842_, data_stage_3__2841_, data_stage_3__2840_, data_stage_3__2839_, data_stage_3__2838_, data_stage_3__2837_, data_stage_3__2836_, data_stage_3__2835_, data_stage_3__2834_, data_stage_3__2833_, data_stage_3__2832_, data_stage_3__2831_, data_stage_3__2830_, data_stage_3__2829_, data_stage_3__2828_, data_stage_3__2827_, data_stage_3__2826_, data_stage_3__2825_, data_stage_3__2824_, data_stage_3__2823_, data_stage_3__2822_, data_stage_3__2821_, data_stage_3__2820_, data_stage_3__2819_, data_stage_3__2818_, data_stage_3__2817_, data_stage_3__2816_, data_stage_3__2815_, data_stage_3__2814_, data_stage_3__2813_, data_stage_3__2812_, data_stage_3__2811_, data_stage_3__2810_, data_stage_3__2809_, data_stage_3__2808_, data_stage_3__2807_, data_stage_3__2806_, data_stage_3__2805_, data_stage_3__2804_, data_stage_3__2803_, data_stage_3__2802_, data_stage_3__2801_, data_stage_3__2800_, data_stage_3__2799_, data_stage_3__2798_, data_stage_3__2797_, data_stage_3__2796_, data_stage_3__2795_, data_stage_3__2794_, data_stage_3__2793_, data_stage_3__2792_, data_stage_3__2791_, data_stage_3__2790_, data_stage_3__2789_, data_stage_3__2788_, data_stage_3__2787_, data_stage_3__2786_, data_stage_3__2785_, data_stage_3__2784_, data_stage_3__2783_, data_stage_3__2782_, data_stage_3__2781_, data_stage_3__2780_, data_stage_3__2779_, data_stage_3__2778_, data_stage_3__2777_, data_stage_3__2776_, data_stage_3__2775_, data_stage_3__2774_, data_stage_3__2773_, data_stage_3__2772_, data_stage_3__2771_, data_stage_3__2770_, data_stage_3__2769_, data_stage_3__2768_, data_stage_3__2767_, data_stage_3__2766_, data_stage_3__2765_, data_stage_3__2764_, data_stage_3__2763_, data_stage_3__2762_, data_stage_3__2761_, data_stage_3__2760_, data_stage_3__2759_, data_stage_3__2758_, data_stage_3__2757_, data_stage_3__2756_, data_stage_3__2755_, data_stage_3__2754_, data_stage_3__2753_, data_stage_3__2752_, data_stage_3__2751_, data_stage_3__2750_, data_stage_3__2749_, data_stage_3__2748_, data_stage_3__2747_, data_stage_3__2746_, data_stage_3__2745_, data_stage_3__2744_, data_stage_3__2743_, data_stage_3__2742_, data_stage_3__2741_, data_stage_3__2740_, data_stage_3__2739_, data_stage_3__2738_, data_stage_3__2737_, data_stage_3__2736_, data_stage_3__2735_, data_stage_3__2734_, data_stage_3__2733_, data_stage_3__2732_, data_stage_3__2731_, data_stage_3__2730_, data_stage_3__2729_, data_stage_3__2728_, data_stage_3__2727_, data_stage_3__2726_, data_stage_3__2725_, data_stage_3__2724_, data_stage_3__2723_, data_stage_3__2722_, data_stage_3__2721_, data_stage_3__2720_, data_stage_3__2719_, data_stage_3__2718_, data_stage_3__2717_, data_stage_3__2716_, data_stage_3__2715_, data_stage_3__2714_, data_stage_3__2713_, data_stage_3__2712_, data_stage_3__2711_, data_stage_3__2710_, data_stage_3__2709_, data_stage_3__2708_, data_stage_3__2707_, data_stage_3__2706_, data_stage_3__2705_, data_stage_3__2704_, data_stage_3__2703_, data_stage_3__2702_, data_stage_3__2701_, data_stage_3__2700_, data_stage_3__2699_, data_stage_3__2698_, data_stage_3__2697_, data_stage_3__2696_, data_stage_3__2695_, data_stage_3__2694_, data_stage_3__2693_, data_stage_3__2692_, data_stage_3__2691_, data_stage_3__2690_, data_stage_3__2689_, data_stage_3__2688_, data_stage_3__2687_, data_stage_3__2686_, data_stage_3__2685_, data_stage_3__2684_, data_stage_3__2683_, data_stage_3__2682_, data_stage_3__2681_, data_stage_3__2680_, data_stage_3__2679_, data_stage_3__2678_, data_stage_3__2677_, data_stage_3__2676_, data_stage_3__2675_, data_stage_3__2674_, data_stage_3__2673_, data_stage_3__2672_, data_stage_3__2671_, data_stage_3__2670_, data_stage_3__2669_, data_stage_3__2668_, data_stage_3__2667_, data_stage_3__2666_, data_stage_3__2665_, data_stage_3__2664_, data_stage_3__2663_, data_stage_3__2662_, data_stage_3__2661_, data_stage_3__2660_, data_stage_3__2659_, data_stage_3__2658_, data_stage_3__2657_, data_stage_3__2656_, data_stage_3__2655_, data_stage_3__2654_, data_stage_3__2653_, data_stage_3__2652_, data_stage_3__2651_, data_stage_3__2650_, data_stage_3__2649_, data_stage_3__2648_, data_stage_3__2647_, data_stage_3__2646_, data_stage_3__2645_, data_stage_3__2644_, data_stage_3__2643_, data_stage_3__2642_, data_stage_3__2641_, data_stage_3__2640_, data_stage_3__2639_, data_stage_3__2638_, data_stage_3__2637_, data_stage_3__2636_, data_stage_3__2635_, data_stage_3__2634_, data_stage_3__2633_, data_stage_3__2632_, data_stage_3__2631_, data_stage_3__2630_, data_stage_3__2629_, data_stage_3__2628_, data_stage_3__2627_, data_stage_3__2626_, data_stage_3__2625_, data_stage_3__2624_, data_stage_3__2623_, data_stage_3__2622_, data_stage_3__2621_, data_stage_3__2620_, data_stage_3__2619_, data_stage_3__2618_, data_stage_3__2617_, data_stage_3__2616_, data_stage_3__2615_, data_stage_3__2614_, data_stage_3__2613_, data_stage_3__2612_, data_stage_3__2611_, data_stage_3__2610_, data_stage_3__2609_, data_stage_3__2608_, data_stage_3__2607_, data_stage_3__2606_, data_stage_3__2605_, data_stage_3__2604_, data_stage_3__2603_, data_stage_3__2602_, data_stage_3__2601_, data_stage_3__2600_, data_stage_3__2599_, data_stage_3__2598_, data_stage_3__2597_, data_stage_3__2596_, data_stage_3__2595_, data_stage_3__2594_, data_stage_3__2593_, data_stage_3__2592_, data_stage_3__2591_, data_stage_3__2590_, data_stage_3__2589_, data_stage_3__2588_, data_stage_3__2587_, data_stage_3__2586_, data_stage_3__2585_, data_stage_3__2584_, data_stage_3__2583_, data_stage_3__2582_, data_stage_3__2581_, data_stage_3__2580_, data_stage_3__2579_, data_stage_3__2578_, data_stage_3__2577_, data_stage_3__2576_, data_stage_3__2575_, data_stage_3__2574_, data_stage_3__2573_, data_stage_3__2572_, data_stage_3__2571_, data_stage_3__2570_, data_stage_3__2569_, data_stage_3__2568_, data_stage_3__2567_, data_stage_3__2566_, data_stage_3__2565_, data_stage_3__2564_, data_stage_3__2563_, data_stage_3__2562_, data_stage_3__2561_, data_stage_3__2560_, data_stage_3__2559_, data_stage_3__2558_, data_stage_3__2557_, data_stage_3__2556_, data_stage_3__2555_, data_stage_3__2554_, data_stage_3__2553_, data_stage_3__2552_, data_stage_3__2551_, data_stage_3__2550_, data_stage_3__2549_, data_stage_3__2548_, data_stage_3__2547_, data_stage_3__2546_, data_stage_3__2545_, data_stage_3__2544_, data_stage_3__2543_, data_stage_3__2542_, data_stage_3__2541_, data_stage_3__2540_, data_stage_3__2539_, data_stage_3__2538_, data_stage_3__2537_, data_stage_3__2536_, data_stage_3__2535_, data_stage_3__2534_, data_stage_3__2533_, data_stage_3__2532_, data_stage_3__2531_, data_stage_3__2530_, data_stage_3__2529_, data_stage_3__2528_, data_stage_3__2527_, data_stage_3__2526_, data_stage_3__2525_, data_stage_3__2524_, data_stage_3__2523_, data_stage_3__2522_, data_stage_3__2521_, data_stage_3__2520_, data_stage_3__2519_, data_stage_3__2518_, data_stage_3__2517_, data_stage_3__2516_, data_stage_3__2515_, data_stage_3__2514_, data_stage_3__2513_, data_stage_3__2512_, data_stage_3__2511_, data_stage_3__2510_, data_stage_3__2509_, data_stage_3__2508_, data_stage_3__2507_, data_stage_3__2506_, data_stage_3__2505_, data_stage_3__2504_, data_stage_3__2503_, data_stage_3__2502_, data_stage_3__2501_, data_stage_3__2500_, data_stage_3__2499_, data_stage_3__2498_, data_stage_3__2497_, data_stage_3__2496_, data_stage_3__2495_, data_stage_3__2494_, data_stage_3__2493_, data_stage_3__2492_, data_stage_3__2491_, data_stage_3__2490_, data_stage_3__2489_, data_stage_3__2488_, data_stage_3__2487_, data_stage_3__2486_, data_stage_3__2485_, data_stage_3__2484_, data_stage_3__2483_, data_stage_3__2482_, data_stage_3__2481_, data_stage_3__2480_, data_stage_3__2479_, data_stage_3__2478_, data_stage_3__2477_, data_stage_3__2476_, data_stage_3__2475_, data_stage_3__2474_, data_stage_3__2473_, data_stage_3__2472_, data_stage_3__2471_, data_stage_3__2470_, data_stage_3__2469_, data_stage_3__2468_, data_stage_3__2467_, data_stage_3__2466_, data_stage_3__2465_, data_stage_3__2464_, data_stage_3__2463_, data_stage_3__2462_, data_stage_3__2461_, data_stage_3__2460_, data_stage_3__2459_, data_stage_3__2458_, data_stage_3__2457_, data_stage_3__2456_, data_stage_3__2455_, data_stage_3__2454_, data_stage_3__2453_, data_stage_3__2452_, data_stage_3__2451_, data_stage_3__2450_, data_stage_3__2449_, data_stage_3__2448_, data_stage_3__2447_, data_stage_3__2446_, data_stage_3__2445_, data_stage_3__2444_, data_stage_3__2443_, data_stage_3__2442_, data_stage_3__2441_, data_stage_3__2440_, data_stage_3__2439_, data_stage_3__2438_, data_stage_3__2437_, data_stage_3__2436_, data_stage_3__2435_, data_stage_3__2434_, data_stage_3__2433_, data_stage_3__2432_, data_stage_3__2431_, data_stage_3__2430_, data_stage_3__2429_, data_stage_3__2428_, data_stage_3__2427_, data_stage_3__2426_, data_stage_3__2425_, data_stage_3__2424_, data_stage_3__2423_, data_stage_3__2422_, data_stage_3__2421_, data_stage_3__2420_, data_stage_3__2419_, data_stage_3__2418_, data_stage_3__2417_, data_stage_3__2416_, data_stage_3__2415_, data_stage_3__2414_, data_stage_3__2413_, data_stage_3__2412_, data_stage_3__2411_, data_stage_3__2410_, data_stage_3__2409_, data_stage_3__2408_, data_stage_3__2407_, data_stage_3__2406_, data_stage_3__2405_, data_stage_3__2404_, data_stage_3__2403_, data_stage_3__2402_, data_stage_3__2401_, data_stage_3__2400_, data_stage_3__2399_, data_stage_3__2398_, data_stage_3__2397_, data_stage_3__2396_, data_stage_3__2395_, data_stage_3__2394_, data_stage_3__2393_, data_stage_3__2392_, data_stage_3__2391_, data_stage_3__2390_, data_stage_3__2389_, data_stage_3__2388_, data_stage_3__2387_, data_stage_3__2386_, data_stage_3__2385_, data_stage_3__2384_, data_stage_3__2383_, data_stage_3__2382_, data_stage_3__2381_, data_stage_3__2380_, data_stage_3__2379_, data_stage_3__2378_, data_stage_3__2377_, data_stage_3__2376_, data_stage_3__2375_, data_stage_3__2374_, data_stage_3__2373_, data_stage_3__2372_, data_stage_3__2371_, data_stage_3__2370_, data_stage_3__2369_, data_stage_3__2368_, data_stage_3__2367_, data_stage_3__2366_, data_stage_3__2365_, data_stage_3__2364_, data_stage_3__2363_, data_stage_3__2362_, data_stage_3__2361_, data_stage_3__2360_, data_stage_3__2359_, data_stage_3__2358_, data_stage_3__2357_, data_stage_3__2356_, data_stage_3__2355_, data_stage_3__2354_, data_stage_3__2353_, data_stage_3__2352_, data_stage_3__2351_, data_stage_3__2350_, data_stage_3__2349_, data_stage_3__2348_, data_stage_3__2347_, data_stage_3__2346_, data_stage_3__2345_, data_stage_3__2344_, data_stage_3__2343_, data_stage_3__2342_, data_stage_3__2341_, data_stage_3__2340_, data_stage_3__2339_, data_stage_3__2338_, data_stage_3__2337_, data_stage_3__2336_, data_stage_3__2335_, data_stage_3__2334_, data_stage_3__2333_, data_stage_3__2332_, data_stage_3__2331_, data_stage_3__2330_, data_stage_3__2329_, data_stage_3__2328_, data_stage_3__2327_, data_stage_3__2326_, data_stage_3__2325_, data_stage_3__2324_, data_stage_3__2323_, data_stage_3__2322_, data_stage_3__2321_, data_stage_3__2320_, data_stage_3__2319_, data_stage_3__2318_, data_stage_3__2317_, data_stage_3__2316_, data_stage_3__2315_, data_stage_3__2314_, data_stage_3__2313_, data_stage_3__2312_, data_stage_3__2311_, data_stage_3__2310_, data_stage_3__2309_, data_stage_3__2308_, data_stage_3__2307_, data_stage_3__2306_, data_stage_3__2305_, data_stage_3__2304_, data_stage_3__2303_, data_stage_3__2302_, data_stage_3__2301_, data_stage_3__2300_, data_stage_3__2299_, data_stage_3__2298_, data_stage_3__2297_, data_stage_3__2296_, data_stage_3__2295_, data_stage_3__2294_, data_stage_3__2293_, data_stage_3__2292_, data_stage_3__2291_, data_stage_3__2290_, data_stage_3__2289_, data_stage_3__2288_, data_stage_3__2287_, data_stage_3__2286_, data_stage_3__2285_, data_stage_3__2284_, data_stage_3__2283_, data_stage_3__2282_, data_stage_3__2281_, data_stage_3__2280_, data_stage_3__2279_, data_stage_3__2278_, data_stage_3__2277_, data_stage_3__2276_, data_stage_3__2275_, data_stage_3__2274_, data_stage_3__2273_, data_stage_3__2272_, data_stage_3__2271_, data_stage_3__2270_, data_stage_3__2269_, data_stage_3__2268_, data_stage_3__2267_, data_stage_3__2266_, data_stage_3__2265_, data_stage_3__2264_, data_stage_3__2263_, data_stage_3__2262_, data_stage_3__2261_, data_stage_3__2260_, data_stage_3__2259_, data_stage_3__2258_, data_stage_3__2257_, data_stage_3__2256_, data_stage_3__2255_, data_stage_3__2254_, data_stage_3__2253_, data_stage_3__2252_, data_stage_3__2251_, data_stage_3__2250_, data_stage_3__2249_, data_stage_3__2248_, data_stage_3__2247_, data_stage_3__2246_, data_stage_3__2245_, data_stage_3__2244_, data_stage_3__2243_, data_stage_3__2242_, data_stage_3__2241_, data_stage_3__2240_, data_stage_3__2239_, data_stage_3__2238_, data_stage_3__2237_, data_stage_3__2236_, data_stage_3__2235_, data_stage_3__2234_, data_stage_3__2233_, data_stage_3__2232_, data_stage_3__2231_, data_stage_3__2230_, data_stage_3__2229_, data_stage_3__2228_, data_stage_3__2227_, data_stage_3__2226_, data_stage_3__2225_, data_stage_3__2224_, data_stage_3__2223_, data_stage_3__2222_, data_stage_3__2221_, data_stage_3__2220_, data_stage_3__2219_, data_stage_3__2218_, data_stage_3__2217_, data_stage_3__2216_, data_stage_3__2215_, data_stage_3__2214_, data_stage_3__2213_, data_stage_3__2212_, data_stage_3__2211_, data_stage_3__2210_, data_stage_3__2209_, data_stage_3__2208_, data_stage_3__2207_, data_stage_3__2206_, data_stage_3__2205_, data_stage_3__2204_, data_stage_3__2203_, data_stage_3__2202_, data_stage_3__2201_, data_stage_3__2200_, data_stage_3__2199_, data_stage_3__2198_, data_stage_3__2197_, data_stage_3__2196_, data_stage_3__2195_, data_stage_3__2194_, data_stage_3__2193_, data_stage_3__2192_, data_stage_3__2191_, data_stage_3__2190_, data_stage_3__2189_, data_stage_3__2188_, data_stage_3__2187_, data_stage_3__2186_, data_stage_3__2185_, data_stage_3__2184_, data_stage_3__2183_, data_stage_3__2182_, data_stage_3__2181_, data_stage_3__2180_, data_stage_3__2179_, data_stage_3__2178_, data_stage_3__2177_, data_stage_3__2176_, data_stage_3__2175_, data_stage_3__2174_, data_stage_3__2173_, data_stage_3__2172_, data_stage_3__2171_, data_stage_3__2170_, data_stage_3__2169_, data_stage_3__2168_, data_stage_3__2167_, data_stage_3__2166_, data_stage_3__2165_, data_stage_3__2164_, data_stage_3__2163_, data_stage_3__2162_, data_stage_3__2161_, data_stage_3__2160_, data_stage_3__2159_, data_stage_3__2158_, data_stage_3__2157_, data_stage_3__2156_, data_stage_3__2155_, data_stage_3__2154_, data_stage_3__2153_, data_stage_3__2152_, data_stage_3__2151_, data_stage_3__2150_, data_stage_3__2149_, data_stage_3__2148_, data_stage_3__2147_, data_stage_3__2146_, data_stage_3__2145_, data_stage_3__2144_, data_stage_3__2143_, data_stage_3__2142_, data_stage_3__2141_, data_stage_3__2140_, data_stage_3__2139_, data_stage_3__2138_, data_stage_3__2137_, data_stage_3__2136_, data_stage_3__2135_, data_stage_3__2134_, data_stage_3__2133_, data_stage_3__2132_, data_stage_3__2131_, data_stage_3__2130_, data_stage_3__2129_, data_stage_3__2128_, data_stage_3__2127_, data_stage_3__2126_, data_stage_3__2125_, data_stage_3__2124_, data_stage_3__2123_, data_stage_3__2122_, data_stage_3__2121_, data_stage_3__2120_, data_stage_3__2119_, data_stage_3__2118_, data_stage_3__2117_, data_stage_3__2116_, data_stage_3__2115_, data_stage_3__2114_, data_stage_3__2113_, data_stage_3__2112_, data_stage_3__2111_, data_stage_3__2110_, data_stage_3__2109_, data_stage_3__2108_, data_stage_3__2107_, data_stage_3__2106_, data_stage_3__2105_, data_stage_3__2104_, data_stage_3__2103_, data_stage_3__2102_, data_stage_3__2101_, data_stage_3__2100_, data_stage_3__2099_, data_stage_3__2098_, data_stage_3__2097_, data_stage_3__2096_, data_stage_3__2095_, data_stage_3__2094_, data_stage_3__2093_, data_stage_3__2092_, data_stage_3__2091_, data_stage_3__2090_, data_stage_3__2089_, data_stage_3__2088_, data_stage_3__2087_, data_stage_3__2086_, data_stage_3__2085_, data_stage_3__2084_, data_stage_3__2083_, data_stage_3__2082_, data_stage_3__2081_, data_stage_3__2080_, data_stage_3__2079_, data_stage_3__2078_, data_stage_3__2077_, data_stage_3__2076_, data_stage_3__2075_, data_stage_3__2074_, data_stage_3__2073_, data_stage_3__2072_, data_stage_3__2071_, data_stage_3__2070_, data_stage_3__2069_, data_stage_3__2068_, data_stage_3__2067_, data_stage_3__2066_, data_stage_3__2065_, data_stage_3__2064_, data_stage_3__2063_, data_stage_3__2062_, data_stage_3__2061_, data_stage_3__2060_, data_stage_3__2059_, data_stage_3__2058_, data_stage_3__2057_, data_stage_3__2056_, data_stage_3__2055_, data_stage_3__2054_, data_stage_3__2053_, data_stage_3__2052_, data_stage_3__2051_, data_stage_3__2050_, data_stage_3__2049_, data_stage_3__2048_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__4095_, data_stage_4__4094_, data_stage_4__4093_, data_stage_4__4092_, data_stage_4__4091_, data_stage_4__4090_, data_stage_4__4089_, data_stage_4__4088_, data_stage_4__4087_, data_stage_4__4086_, data_stage_4__4085_, data_stage_4__4084_, data_stage_4__4083_, data_stage_4__4082_, data_stage_4__4081_, data_stage_4__4080_, data_stage_4__4079_, data_stage_4__4078_, data_stage_4__4077_, data_stage_4__4076_, data_stage_4__4075_, data_stage_4__4074_, data_stage_4__4073_, data_stage_4__4072_, data_stage_4__4071_, data_stage_4__4070_, data_stage_4__4069_, data_stage_4__4068_, data_stage_4__4067_, data_stage_4__4066_, data_stage_4__4065_, data_stage_4__4064_, data_stage_4__4063_, data_stage_4__4062_, data_stage_4__4061_, data_stage_4__4060_, data_stage_4__4059_, data_stage_4__4058_, data_stage_4__4057_, data_stage_4__4056_, data_stage_4__4055_, data_stage_4__4054_, data_stage_4__4053_, data_stage_4__4052_, data_stage_4__4051_, data_stage_4__4050_, data_stage_4__4049_, data_stage_4__4048_, data_stage_4__4047_, data_stage_4__4046_, data_stage_4__4045_, data_stage_4__4044_, data_stage_4__4043_, data_stage_4__4042_, data_stage_4__4041_, data_stage_4__4040_, data_stage_4__4039_, data_stage_4__4038_, data_stage_4__4037_, data_stage_4__4036_, data_stage_4__4035_, data_stage_4__4034_, data_stage_4__4033_, data_stage_4__4032_, data_stage_4__4031_, data_stage_4__4030_, data_stage_4__4029_, data_stage_4__4028_, data_stage_4__4027_, data_stage_4__4026_, data_stage_4__4025_, data_stage_4__4024_, data_stage_4__4023_, data_stage_4__4022_, data_stage_4__4021_, data_stage_4__4020_, data_stage_4__4019_, data_stage_4__4018_, data_stage_4__4017_, data_stage_4__4016_, data_stage_4__4015_, data_stage_4__4014_, data_stage_4__4013_, data_stage_4__4012_, data_stage_4__4011_, data_stage_4__4010_, data_stage_4__4009_, data_stage_4__4008_, data_stage_4__4007_, data_stage_4__4006_, data_stage_4__4005_, data_stage_4__4004_, data_stage_4__4003_, data_stage_4__4002_, data_stage_4__4001_, data_stage_4__4000_, data_stage_4__3999_, data_stage_4__3998_, data_stage_4__3997_, data_stage_4__3996_, data_stage_4__3995_, data_stage_4__3994_, data_stage_4__3993_, data_stage_4__3992_, data_stage_4__3991_, data_stage_4__3990_, data_stage_4__3989_, data_stage_4__3988_, data_stage_4__3987_, data_stage_4__3986_, data_stage_4__3985_, data_stage_4__3984_, data_stage_4__3983_, data_stage_4__3982_, data_stage_4__3981_, data_stage_4__3980_, data_stage_4__3979_, data_stage_4__3978_, data_stage_4__3977_, data_stage_4__3976_, data_stage_4__3975_, data_stage_4__3974_, data_stage_4__3973_, data_stage_4__3972_, data_stage_4__3971_, data_stage_4__3970_, data_stage_4__3969_, data_stage_4__3968_, data_stage_4__3967_, data_stage_4__3966_, data_stage_4__3965_, data_stage_4__3964_, data_stage_4__3963_, data_stage_4__3962_, data_stage_4__3961_, data_stage_4__3960_, data_stage_4__3959_, data_stage_4__3958_, data_stage_4__3957_, data_stage_4__3956_, data_stage_4__3955_, data_stage_4__3954_, data_stage_4__3953_, data_stage_4__3952_, data_stage_4__3951_, data_stage_4__3950_, data_stage_4__3949_, data_stage_4__3948_, data_stage_4__3947_, data_stage_4__3946_, data_stage_4__3945_, data_stage_4__3944_, data_stage_4__3943_, data_stage_4__3942_, data_stage_4__3941_, data_stage_4__3940_, data_stage_4__3939_, data_stage_4__3938_, data_stage_4__3937_, data_stage_4__3936_, data_stage_4__3935_, data_stage_4__3934_, data_stage_4__3933_, data_stage_4__3932_, data_stage_4__3931_, data_stage_4__3930_, data_stage_4__3929_, data_stage_4__3928_, data_stage_4__3927_, data_stage_4__3926_, data_stage_4__3925_, data_stage_4__3924_, data_stage_4__3923_, data_stage_4__3922_, data_stage_4__3921_, data_stage_4__3920_, data_stage_4__3919_, data_stage_4__3918_, data_stage_4__3917_, data_stage_4__3916_, data_stage_4__3915_, data_stage_4__3914_, data_stage_4__3913_, data_stage_4__3912_, data_stage_4__3911_, data_stage_4__3910_, data_stage_4__3909_, data_stage_4__3908_, data_stage_4__3907_, data_stage_4__3906_, data_stage_4__3905_, data_stage_4__3904_, data_stage_4__3903_, data_stage_4__3902_, data_stage_4__3901_, data_stage_4__3900_, data_stage_4__3899_, data_stage_4__3898_, data_stage_4__3897_, data_stage_4__3896_, data_stage_4__3895_, data_stage_4__3894_, data_stage_4__3893_, data_stage_4__3892_, data_stage_4__3891_, data_stage_4__3890_, data_stage_4__3889_, data_stage_4__3888_, data_stage_4__3887_, data_stage_4__3886_, data_stage_4__3885_, data_stage_4__3884_, data_stage_4__3883_, data_stage_4__3882_, data_stage_4__3881_, data_stage_4__3880_, data_stage_4__3879_, data_stage_4__3878_, data_stage_4__3877_, data_stage_4__3876_, data_stage_4__3875_, data_stage_4__3874_, data_stage_4__3873_, data_stage_4__3872_, data_stage_4__3871_, data_stage_4__3870_, data_stage_4__3869_, data_stage_4__3868_, data_stage_4__3867_, data_stage_4__3866_, data_stage_4__3865_, data_stage_4__3864_, data_stage_4__3863_, data_stage_4__3862_, data_stage_4__3861_, data_stage_4__3860_, data_stage_4__3859_, data_stage_4__3858_, data_stage_4__3857_, data_stage_4__3856_, data_stage_4__3855_, data_stage_4__3854_, data_stage_4__3853_, data_stage_4__3852_, data_stage_4__3851_, data_stage_4__3850_, data_stage_4__3849_, data_stage_4__3848_, data_stage_4__3847_, data_stage_4__3846_, data_stage_4__3845_, data_stage_4__3844_, data_stage_4__3843_, data_stage_4__3842_, data_stage_4__3841_, data_stage_4__3840_, data_stage_4__3839_, data_stage_4__3838_, data_stage_4__3837_, data_stage_4__3836_, data_stage_4__3835_, data_stage_4__3834_, data_stage_4__3833_, data_stage_4__3832_, data_stage_4__3831_, data_stage_4__3830_, data_stage_4__3829_, data_stage_4__3828_, data_stage_4__3827_, data_stage_4__3826_, data_stage_4__3825_, data_stage_4__3824_, data_stage_4__3823_, data_stage_4__3822_, data_stage_4__3821_, data_stage_4__3820_, data_stage_4__3819_, data_stage_4__3818_, data_stage_4__3817_, data_stage_4__3816_, data_stage_4__3815_, data_stage_4__3814_, data_stage_4__3813_, data_stage_4__3812_, data_stage_4__3811_, data_stage_4__3810_, data_stage_4__3809_, data_stage_4__3808_, data_stage_4__3807_, data_stage_4__3806_, data_stage_4__3805_, data_stage_4__3804_, data_stage_4__3803_, data_stage_4__3802_, data_stage_4__3801_, data_stage_4__3800_, data_stage_4__3799_, data_stage_4__3798_, data_stage_4__3797_, data_stage_4__3796_, data_stage_4__3795_, data_stage_4__3794_, data_stage_4__3793_, data_stage_4__3792_, data_stage_4__3791_, data_stage_4__3790_, data_stage_4__3789_, data_stage_4__3788_, data_stage_4__3787_, data_stage_4__3786_, data_stage_4__3785_, data_stage_4__3784_, data_stage_4__3783_, data_stage_4__3782_, data_stage_4__3781_, data_stage_4__3780_, data_stage_4__3779_, data_stage_4__3778_, data_stage_4__3777_, data_stage_4__3776_, data_stage_4__3775_, data_stage_4__3774_, data_stage_4__3773_, data_stage_4__3772_, data_stage_4__3771_, data_stage_4__3770_, data_stage_4__3769_, data_stage_4__3768_, data_stage_4__3767_, data_stage_4__3766_, data_stage_4__3765_, data_stage_4__3764_, data_stage_4__3763_, data_stage_4__3762_, data_stage_4__3761_, data_stage_4__3760_, data_stage_4__3759_, data_stage_4__3758_, data_stage_4__3757_, data_stage_4__3756_, data_stage_4__3755_, data_stage_4__3754_, data_stage_4__3753_, data_stage_4__3752_, data_stage_4__3751_, data_stage_4__3750_, data_stage_4__3749_, data_stage_4__3748_, data_stage_4__3747_, data_stage_4__3746_, data_stage_4__3745_, data_stage_4__3744_, data_stage_4__3743_, data_stage_4__3742_, data_stage_4__3741_, data_stage_4__3740_, data_stage_4__3739_, data_stage_4__3738_, data_stage_4__3737_, data_stage_4__3736_, data_stage_4__3735_, data_stage_4__3734_, data_stage_4__3733_, data_stage_4__3732_, data_stage_4__3731_, data_stage_4__3730_, data_stage_4__3729_, data_stage_4__3728_, data_stage_4__3727_, data_stage_4__3726_, data_stage_4__3725_, data_stage_4__3724_, data_stage_4__3723_, data_stage_4__3722_, data_stage_4__3721_, data_stage_4__3720_, data_stage_4__3719_, data_stage_4__3718_, data_stage_4__3717_, data_stage_4__3716_, data_stage_4__3715_, data_stage_4__3714_, data_stage_4__3713_, data_stage_4__3712_, data_stage_4__3711_, data_stage_4__3710_, data_stage_4__3709_, data_stage_4__3708_, data_stage_4__3707_, data_stage_4__3706_, data_stage_4__3705_, data_stage_4__3704_, data_stage_4__3703_, data_stage_4__3702_, data_stage_4__3701_, data_stage_4__3700_, data_stage_4__3699_, data_stage_4__3698_, data_stage_4__3697_, data_stage_4__3696_, data_stage_4__3695_, data_stage_4__3694_, data_stage_4__3693_, data_stage_4__3692_, data_stage_4__3691_, data_stage_4__3690_, data_stage_4__3689_, data_stage_4__3688_, data_stage_4__3687_, data_stage_4__3686_, data_stage_4__3685_, data_stage_4__3684_, data_stage_4__3683_, data_stage_4__3682_, data_stage_4__3681_, data_stage_4__3680_, data_stage_4__3679_, data_stage_4__3678_, data_stage_4__3677_, data_stage_4__3676_, data_stage_4__3675_, data_stage_4__3674_, data_stage_4__3673_, data_stage_4__3672_, data_stage_4__3671_, data_stage_4__3670_, data_stage_4__3669_, data_stage_4__3668_, data_stage_4__3667_, data_stage_4__3666_, data_stage_4__3665_, data_stage_4__3664_, data_stage_4__3663_, data_stage_4__3662_, data_stage_4__3661_, data_stage_4__3660_, data_stage_4__3659_, data_stage_4__3658_, data_stage_4__3657_, data_stage_4__3656_, data_stage_4__3655_, data_stage_4__3654_, data_stage_4__3653_, data_stage_4__3652_, data_stage_4__3651_, data_stage_4__3650_, data_stage_4__3649_, data_stage_4__3648_, data_stage_4__3647_, data_stage_4__3646_, data_stage_4__3645_, data_stage_4__3644_, data_stage_4__3643_, data_stage_4__3642_, data_stage_4__3641_, data_stage_4__3640_, data_stage_4__3639_, data_stage_4__3638_, data_stage_4__3637_, data_stage_4__3636_, data_stage_4__3635_, data_stage_4__3634_, data_stage_4__3633_, data_stage_4__3632_, data_stage_4__3631_, data_stage_4__3630_, data_stage_4__3629_, data_stage_4__3628_, data_stage_4__3627_, data_stage_4__3626_, data_stage_4__3625_, data_stage_4__3624_, data_stage_4__3623_, data_stage_4__3622_, data_stage_4__3621_, data_stage_4__3620_, data_stage_4__3619_, data_stage_4__3618_, data_stage_4__3617_, data_stage_4__3616_, data_stage_4__3615_, data_stage_4__3614_, data_stage_4__3613_, data_stage_4__3612_, data_stage_4__3611_, data_stage_4__3610_, data_stage_4__3609_, data_stage_4__3608_, data_stage_4__3607_, data_stage_4__3606_, data_stage_4__3605_, data_stage_4__3604_, data_stage_4__3603_, data_stage_4__3602_, data_stage_4__3601_, data_stage_4__3600_, data_stage_4__3599_, data_stage_4__3598_, data_stage_4__3597_, data_stage_4__3596_, data_stage_4__3595_, data_stage_4__3594_, data_stage_4__3593_, data_stage_4__3592_, data_stage_4__3591_, data_stage_4__3590_, data_stage_4__3589_, data_stage_4__3588_, data_stage_4__3587_, data_stage_4__3586_, data_stage_4__3585_, data_stage_4__3584_, data_stage_4__3583_, data_stage_4__3582_, data_stage_4__3581_, data_stage_4__3580_, data_stage_4__3579_, data_stage_4__3578_, data_stage_4__3577_, data_stage_4__3576_, data_stage_4__3575_, data_stage_4__3574_, data_stage_4__3573_, data_stage_4__3572_, data_stage_4__3571_, data_stage_4__3570_, data_stage_4__3569_, data_stage_4__3568_, data_stage_4__3567_, data_stage_4__3566_, data_stage_4__3565_, data_stage_4__3564_, data_stage_4__3563_, data_stage_4__3562_, data_stage_4__3561_, data_stage_4__3560_, data_stage_4__3559_, data_stage_4__3558_, data_stage_4__3557_, data_stage_4__3556_, data_stage_4__3555_, data_stage_4__3554_, data_stage_4__3553_, data_stage_4__3552_, data_stage_4__3551_, data_stage_4__3550_, data_stage_4__3549_, data_stage_4__3548_, data_stage_4__3547_, data_stage_4__3546_, data_stage_4__3545_, data_stage_4__3544_, data_stage_4__3543_, data_stage_4__3542_, data_stage_4__3541_, data_stage_4__3540_, data_stage_4__3539_, data_stage_4__3538_, data_stage_4__3537_, data_stage_4__3536_, data_stage_4__3535_, data_stage_4__3534_, data_stage_4__3533_, data_stage_4__3532_, data_stage_4__3531_, data_stage_4__3530_, data_stage_4__3529_, data_stage_4__3528_, data_stage_4__3527_, data_stage_4__3526_, data_stage_4__3525_, data_stage_4__3524_, data_stage_4__3523_, data_stage_4__3522_, data_stage_4__3521_, data_stage_4__3520_, data_stage_4__3519_, data_stage_4__3518_, data_stage_4__3517_, data_stage_4__3516_, data_stage_4__3515_, data_stage_4__3514_, data_stage_4__3513_, data_stage_4__3512_, data_stage_4__3511_, data_stage_4__3510_, data_stage_4__3509_, data_stage_4__3508_, data_stage_4__3507_, data_stage_4__3506_, data_stage_4__3505_, data_stage_4__3504_, data_stage_4__3503_, data_stage_4__3502_, data_stage_4__3501_, data_stage_4__3500_, data_stage_4__3499_, data_stage_4__3498_, data_stage_4__3497_, data_stage_4__3496_, data_stage_4__3495_, data_stage_4__3494_, data_stage_4__3493_, data_stage_4__3492_, data_stage_4__3491_, data_stage_4__3490_, data_stage_4__3489_, data_stage_4__3488_, data_stage_4__3487_, data_stage_4__3486_, data_stage_4__3485_, data_stage_4__3484_, data_stage_4__3483_, data_stage_4__3482_, data_stage_4__3481_, data_stage_4__3480_, data_stage_4__3479_, data_stage_4__3478_, data_stage_4__3477_, data_stage_4__3476_, data_stage_4__3475_, data_stage_4__3474_, data_stage_4__3473_, data_stage_4__3472_, data_stage_4__3471_, data_stage_4__3470_, data_stage_4__3469_, data_stage_4__3468_, data_stage_4__3467_, data_stage_4__3466_, data_stage_4__3465_, data_stage_4__3464_, data_stage_4__3463_, data_stage_4__3462_, data_stage_4__3461_, data_stage_4__3460_, data_stage_4__3459_, data_stage_4__3458_, data_stage_4__3457_, data_stage_4__3456_, data_stage_4__3455_, data_stage_4__3454_, data_stage_4__3453_, data_stage_4__3452_, data_stage_4__3451_, data_stage_4__3450_, data_stage_4__3449_, data_stage_4__3448_, data_stage_4__3447_, data_stage_4__3446_, data_stage_4__3445_, data_stage_4__3444_, data_stage_4__3443_, data_stage_4__3442_, data_stage_4__3441_, data_stage_4__3440_, data_stage_4__3439_, data_stage_4__3438_, data_stage_4__3437_, data_stage_4__3436_, data_stage_4__3435_, data_stage_4__3434_, data_stage_4__3433_, data_stage_4__3432_, data_stage_4__3431_, data_stage_4__3430_, data_stage_4__3429_, data_stage_4__3428_, data_stage_4__3427_, data_stage_4__3426_, data_stage_4__3425_, data_stage_4__3424_, data_stage_4__3423_, data_stage_4__3422_, data_stage_4__3421_, data_stage_4__3420_, data_stage_4__3419_, data_stage_4__3418_, data_stage_4__3417_, data_stage_4__3416_, data_stage_4__3415_, data_stage_4__3414_, data_stage_4__3413_, data_stage_4__3412_, data_stage_4__3411_, data_stage_4__3410_, data_stage_4__3409_, data_stage_4__3408_, data_stage_4__3407_, data_stage_4__3406_, data_stage_4__3405_, data_stage_4__3404_, data_stage_4__3403_, data_stage_4__3402_, data_stage_4__3401_, data_stage_4__3400_, data_stage_4__3399_, data_stage_4__3398_, data_stage_4__3397_, data_stage_4__3396_, data_stage_4__3395_, data_stage_4__3394_, data_stage_4__3393_, data_stage_4__3392_, data_stage_4__3391_, data_stage_4__3390_, data_stage_4__3389_, data_stage_4__3388_, data_stage_4__3387_, data_stage_4__3386_, data_stage_4__3385_, data_stage_4__3384_, data_stage_4__3383_, data_stage_4__3382_, data_stage_4__3381_, data_stage_4__3380_, data_stage_4__3379_, data_stage_4__3378_, data_stage_4__3377_, data_stage_4__3376_, data_stage_4__3375_, data_stage_4__3374_, data_stage_4__3373_, data_stage_4__3372_, data_stage_4__3371_, data_stage_4__3370_, data_stage_4__3369_, data_stage_4__3368_, data_stage_4__3367_, data_stage_4__3366_, data_stage_4__3365_, data_stage_4__3364_, data_stage_4__3363_, data_stage_4__3362_, data_stage_4__3361_, data_stage_4__3360_, data_stage_4__3359_, data_stage_4__3358_, data_stage_4__3357_, data_stage_4__3356_, data_stage_4__3355_, data_stage_4__3354_, data_stage_4__3353_, data_stage_4__3352_, data_stage_4__3351_, data_stage_4__3350_, data_stage_4__3349_, data_stage_4__3348_, data_stage_4__3347_, data_stage_4__3346_, data_stage_4__3345_, data_stage_4__3344_, data_stage_4__3343_, data_stage_4__3342_, data_stage_4__3341_, data_stage_4__3340_, data_stage_4__3339_, data_stage_4__3338_, data_stage_4__3337_, data_stage_4__3336_, data_stage_4__3335_, data_stage_4__3334_, data_stage_4__3333_, data_stage_4__3332_, data_stage_4__3331_, data_stage_4__3330_, data_stage_4__3329_, data_stage_4__3328_, data_stage_4__3327_, data_stage_4__3326_, data_stage_4__3325_, data_stage_4__3324_, data_stage_4__3323_, data_stage_4__3322_, data_stage_4__3321_, data_stage_4__3320_, data_stage_4__3319_, data_stage_4__3318_, data_stage_4__3317_, data_stage_4__3316_, data_stage_4__3315_, data_stage_4__3314_, data_stage_4__3313_, data_stage_4__3312_, data_stage_4__3311_, data_stage_4__3310_, data_stage_4__3309_, data_stage_4__3308_, data_stage_4__3307_, data_stage_4__3306_, data_stage_4__3305_, data_stage_4__3304_, data_stage_4__3303_, data_stage_4__3302_, data_stage_4__3301_, data_stage_4__3300_, data_stage_4__3299_, data_stage_4__3298_, data_stage_4__3297_, data_stage_4__3296_, data_stage_4__3295_, data_stage_4__3294_, data_stage_4__3293_, data_stage_4__3292_, data_stage_4__3291_, data_stage_4__3290_, data_stage_4__3289_, data_stage_4__3288_, data_stage_4__3287_, data_stage_4__3286_, data_stage_4__3285_, data_stage_4__3284_, data_stage_4__3283_, data_stage_4__3282_, data_stage_4__3281_, data_stage_4__3280_, data_stage_4__3279_, data_stage_4__3278_, data_stage_4__3277_, data_stage_4__3276_, data_stage_4__3275_, data_stage_4__3274_, data_stage_4__3273_, data_stage_4__3272_, data_stage_4__3271_, data_stage_4__3270_, data_stage_4__3269_, data_stage_4__3268_, data_stage_4__3267_, data_stage_4__3266_, data_stage_4__3265_, data_stage_4__3264_, data_stage_4__3263_, data_stage_4__3262_, data_stage_4__3261_, data_stage_4__3260_, data_stage_4__3259_, data_stage_4__3258_, data_stage_4__3257_, data_stage_4__3256_, data_stage_4__3255_, data_stage_4__3254_, data_stage_4__3253_, data_stage_4__3252_, data_stage_4__3251_, data_stage_4__3250_, data_stage_4__3249_, data_stage_4__3248_, data_stage_4__3247_, data_stage_4__3246_, data_stage_4__3245_, data_stage_4__3244_, data_stage_4__3243_, data_stage_4__3242_, data_stage_4__3241_, data_stage_4__3240_, data_stage_4__3239_, data_stage_4__3238_, data_stage_4__3237_, data_stage_4__3236_, data_stage_4__3235_, data_stage_4__3234_, data_stage_4__3233_, data_stage_4__3232_, data_stage_4__3231_, data_stage_4__3230_, data_stage_4__3229_, data_stage_4__3228_, data_stage_4__3227_, data_stage_4__3226_, data_stage_4__3225_, data_stage_4__3224_, data_stage_4__3223_, data_stage_4__3222_, data_stage_4__3221_, data_stage_4__3220_, data_stage_4__3219_, data_stage_4__3218_, data_stage_4__3217_, data_stage_4__3216_, data_stage_4__3215_, data_stage_4__3214_, data_stage_4__3213_, data_stage_4__3212_, data_stage_4__3211_, data_stage_4__3210_, data_stage_4__3209_, data_stage_4__3208_, data_stage_4__3207_, data_stage_4__3206_, data_stage_4__3205_, data_stage_4__3204_, data_stage_4__3203_, data_stage_4__3202_, data_stage_4__3201_, data_stage_4__3200_, data_stage_4__3199_, data_stage_4__3198_, data_stage_4__3197_, data_stage_4__3196_, data_stage_4__3195_, data_stage_4__3194_, data_stage_4__3193_, data_stage_4__3192_, data_stage_4__3191_, data_stage_4__3190_, data_stage_4__3189_, data_stage_4__3188_, data_stage_4__3187_, data_stage_4__3186_, data_stage_4__3185_, data_stage_4__3184_, data_stage_4__3183_, data_stage_4__3182_, data_stage_4__3181_, data_stage_4__3180_, data_stage_4__3179_, data_stage_4__3178_, data_stage_4__3177_, data_stage_4__3176_, data_stage_4__3175_, data_stage_4__3174_, data_stage_4__3173_, data_stage_4__3172_, data_stage_4__3171_, data_stage_4__3170_, data_stage_4__3169_, data_stage_4__3168_, data_stage_4__3167_, data_stage_4__3166_, data_stage_4__3165_, data_stage_4__3164_, data_stage_4__3163_, data_stage_4__3162_, data_stage_4__3161_, data_stage_4__3160_, data_stage_4__3159_, data_stage_4__3158_, data_stage_4__3157_, data_stage_4__3156_, data_stage_4__3155_, data_stage_4__3154_, data_stage_4__3153_, data_stage_4__3152_, data_stage_4__3151_, data_stage_4__3150_, data_stage_4__3149_, data_stage_4__3148_, data_stage_4__3147_, data_stage_4__3146_, data_stage_4__3145_, data_stage_4__3144_, data_stage_4__3143_, data_stage_4__3142_, data_stage_4__3141_, data_stage_4__3140_, data_stage_4__3139_, data_stage_4__3138_, data_stage_4__3137_, data_stage_4__3136_, data_stage_4__3135_, data_stage_4__3134_, data_stage_4__3133_, data_stage_4__3132_, data_stage_4__3131_, data_stage_4__3130_, data_stage_4__3129_, data_stage_4__3128_, data_stage_4__3127_, data_stage_4__3126_, data_stage_4__3125_, data_stage_4__3124_, data_stage_4__3123_, data_stage_4__3122_, data_stage_4__3121_, data_stage_4__3120_, data_stage_4__3119_, data_stage_4__3118_, data_stage_4__3117_, data_stage_4__3116_, data_stage_4__3115_, data_stage_4__3114_, data_stage_4__3113_, data_stage_4__3112_, data_stage_4__3111_, data_stage_4__3110_, data_stage_4__3109_, data_stage_4__3108_, data_stage_4__3107_, data_stage_4__3106_, data_stage_4__3105_, data_stage_4__3104_, data_stage_4__3103_, data_stage_4__3102_, data_stage_4__3101_, data_stage_4__3100_, data_stage_4__3099_, data_stage_4__3098_, data_stage_4__3097_, data_stage_4__3096_, data_stage_4__3095_, data_stage_4__3094_, data_stage_4__3093_, data_stage_4__3092_, data_stage_4__3091_, data_stage_4__3090_, data_stage_4__3089_, data_stage_4__3088_, data_stage_4__3087_, data_stage_4__3086_, data_stage_4__3085_, data_stage_4__3084_, data_stage_4__3083_, data_stage_4__3082_, data_stage_4__3081_, data_stage_4__3080_, data_stage_4__3079_, data_stage_4__3078_, data_stage_4__3077_, data_stage_4__3076_, data_stage_4__3075_, data_stage_4__3074_, data_stage_4__3073_, data_stage_4__3072_, data_stage_4__3071_, data_stage_4__3070_, data_stage_4__3069_, data_stage_4__3068_, data_stage_4__3067_, data_stage_4__3066_, data_stage_4__3065_, data_stage_4__3064_, data_stage_4__3063_, data_stage_4__3062_, data_stage_4__3061_, data_stage_4__3060_, data_stage_4__3059_, data_stage_4__3058_, data_stage_4__3057_, data_stage_4__3056_, data_stage_4__3055_, data_stage_4__3054_, data_stage_4__3053_, data_stage_4__3052_, data_stage_4__3051_, data_stage_4__3050_, data_stage_4__3049_, data_stage_4__3048_, data_stage_4__3047_, data_stage_4__3046_, data_stage_4__3045_, data_stage_4__3044_, data_stage_4__3043_, data_stage_4__3042_, data_stage_4__3041_, data_stage_4__3040_, data_stage_4__3039_, data_stage_4__3038_, data_stage_4__3037_, data_stage_4__3036_, data_stage_4__3035_, data_stage_4__3034_, data_stage_4__3033_, data_stage_4__3032_, data_stage_4__3031_, data_stage_4__3030_, data_stage_4__3029_, data_stage_4__3028_, data_stage_4__3027_, data_stage_4__3026_, data_stage_4__3025_, data_stage_4__3024_, data_stage_4__3023_, data_stage_4__3022_, data_stage_4__3021_, data_stage_4__3020_, data_stage_4__3019_, data_stage_4__3018_, data_stage_4__3017_, data_stage_4__3016_, data_stage_4__3015_, data_stage_4__3014_, data_stage_4__3013_, data_stage_4__3012_, data_stage_4__3011_, data_stage_4__3010_, data_stage_4__3009_, data_stage_4__3008_, data_stage_4__3007_, data_stage_4__3006_, data_stage_4__3005_, data_stage_4__3004_, data_stage_4__3003_, data_stage_4__3002_, data_stage_4__3001_, data_stage_4__3000_, data_stage_4__2999_, data_stage_4__2998_, data_stage_4__2997_, data_stage_4__2996_, data_stage_4__2995_, data_stage_4__2994_, data_stage_4__2993_, data_stage_4__2992_, data_stage_4__2991_, data_stage_4__2990_, data_stage_4__2989_, data_stage_4__2988_, data_stage_4__2987_, data_stage_4__2986_, data_stage_4__2985_, data_stage_4__2984_, data_stage_4__2983_, data_stage_4__2982_, data_stage_4__2981_, data_stage_4__2980_, data_stage_4__2979_, data_stage_4__2978_, data_stage_4__2977_, data_stage_4__2976_, data_stage_4__2975_, data_stage_4__2974_, data_stage_4__2973_, data_stage_4__2972_, data_stage_4__2971_, data_stage_4__2970_, data_stage_4__2969_, data_stage_4__2968_, data_stage_4__2967_, data_stage_4__2966_, data_stage_4__2965_, data_stage_4__2964_, data_stage_4__2963_, data_stage_4__2962_, data_stage_4__2961_, data_stage_4__2960_, data_stage_4__2959_, data_stage_4__2958_, data_stage_4__2957_, data_stage_4__2956_, data_stage_4__2955_, data_stage_4__2954_, data_stage_4__2953_, data_stage_4__2952_, data_stage_4__2951_, data_stage_4__2950_, data_stage_4__2949_, data_stage_4__2948_, data_stage_4__2947_, data_stage_4__2946_, data_stage_4__2945_, data_stage_4__2944_, data_stage_4__2943_, data_stage_4__2942_, data_stage_4__2941_, data_stage_4__2940_, data_stage_4__2939_, data_stage_4__2938_, data_stage_4__2937_, data_stage_4__2936_, data_stage_4__2935_, data_stage_4__2934_, data_stage_4__2933_, data_stage_4__2932_, data_stage_4__2931_, data_stage_4__2930_, data_stage_4__2929_, data_stage_4__2928_, data_stage_4__2927_, data_stage_4__2926_, data_stage_4__2925_, data_stage_4__2924_, data_stage_4__2923_, data_stage_4__2922_, data_stage_4__2921_, data_stage_4__2920_, data_stage_4__2919_, data_stage_4__2918_, data_stage_4__2917_, data_stage_4__2916_, data_stage_4__2915_, data_stage_4__2914_, data_stage_4__2913_, data_stage_4__2912_, data_stage_4__2911_, data_stage_4__2910_, data_stage_4__2909_, data_stage_4__2908_, data_stage_4__2907_, data_stage_4__2906_, data_stage_4__2905_, data_stage_4__2904_, data_stage_4__2903_, data_stage_4__2902_, data_stage_4__2901_, data_stage_4__2900_, data_stage_4__2899_, data_stage_4__2898_, data_stage_4__2897_, data_stage_4__2896_, data_stage_4__2895_, data_stage_4__2894_, data_stage_4__2893_, data_stage_4__2892_, data_stage_4__2891_, data_stage_4__2890_, data_stage_4__2889_, data_stage_4__2888_, data_stage_4__2887_, data_stage_4__2886_, data_stage_4__2885_, data_stage_4__2884_, data_stage_4__2883_, data_stage_4__2882_, data_stage_4__2881_, data_stage_4__2880_, data_stage_4__2879_, data_stage_4__2878_, data_stage_4__2877_, data_stage_4__2876_, data_stage_4__2875_, data_stage_4__2874_, data_stage_4__2873_, data_stage_4__2872_, data_stage_4__2871_, data_stage_4__2870_, data_stage_4__2869_, data_stage_4__2868_, data_stage_4__2867_, data_stage_4__2866_, data_stage_4__2865_, data_stage_4__2864_, data_stage_4__2863_, data_stage_4__2862_, data_stage_4__2861_, data_stage_4__2860_, data_stage_4__2859_, data_stage_4__2858_, data_stage_4__2857_, data_stage_4__2856_, data_stage_4__2855_, data_stage_4__2854_, data_stage_4__2853_, data_stage_4__2852_, data_stage_4__2851_, data_stage_4__2850_, data_stage_4__2849_, data_stage_4__2848_, data_stage_4__2847_, data_stage_4__2846_, data_stage_4__2845_, data_stage_4__2844_, data_stage_4__2843_, data_stage_4__2842_, data_stage_4__2841_, data_stage_4__2840_, data_stage_4__2839_, data_stage_4__2838_, data_stage_4__2837_, data_stage_4__2836_, data_stage_4__2835_, data_stage_4__2834_, data_stage_4__2833_, data_stage_4__2832_, data_stage_4__2831_, data_stage_4__2830_, data_stage_4__2829_, data_stage_4__2828_, data_stage_4__2827_, data_stage_4__2826_, data_stage_4__2825_, data_stage_4__2824_, data_stage_4__2823_, data_stage_4__2822_, data_stage_4__2821_, data_stage_4__2820_, data_stage_4__2819_, data_stage_4__2818_, data_stage_4__2817_, data_stage_4__2816_, data_stage_4__2815_, data_stage_4__2814_, data_stage_4__2813_, data_stage_4__2812_, data_stage_4__2811_, data_stage_4__2810_, data_stage_4__2809_, data_stage_4__2808_, data_stage_4__2807_, data_stage_4__2806_, data_stage_4__2805_, data_stage_4__2804_, data_stage_4__2803_, data_stage_4__2802_, data_stage_4__2801_, data_stage_4__2800_, data_stage_4__2799_, data_stage_4__2798_, data_stage_4__2797_, data_stage_4__2796_, data_stage_4__2795_, data_stage_4__2794_, data_stage_4__2793_, data_stage_4__2792_, data_stage_4__2791_, data_stage_4__2790_, data_stage_4__2789_, data_stage_4__2788_, data_stage_4__2787_, data_stage_4__2786_, data_stage_4__2785_, data_stage_4__2784_, data_stage_4__2783_, data_stage_4__2782_, data_stage_4__2781_, data_stage_4__2780_, data_stage_4__2779_, data_stage_4__2778_, data_stage_4__2777_, data_stage_4__2776_, data_stage_4__2775_, data_stage_4__2774_, data_stage_4__2773_, data_stage_4__2772_, data_stage_4__2771_, data_stage_4__2770_, data_stage_4__2769_, data_stage_4__2768_, data_stage_4__2767_, data_stage_4__2766_, data_stage_4__2765_, data_stage_4__2764_, data_stage_4__2763_, data_stage_4__2762_, data_stage_4__2761_, data_stage_4__2760_, data_stage_4__2759_, data_stage_4__2758_, data_stage_4__2757_, data_stage_4__2756_, data_stage_4__2755_, data_stage_4__2754_, data_stage_4__2753_, data_stage_4__2752_, data_stage_4__2751_, data_stage_4__2750_, data_stage_4__2749_, data_stage_4__2748_, data_stage_4__2747_, data_stage_4__2746_, data_stage_4__2745_, data_stage_4__2744_, data_stage_4__2743_, data_stage_4__2742_, data_stage_4__2741_, data_stage_4__2740_, data_stage_4__2739_, data_stage_4__2738_, data_stage_4__2737_, data_stage_4__2736_, data_stage_4__2735_, data_stage_4__2734_, data_stage_4__2733_, data_stage_4__2732_, data_stage_4__2731_, data_stage_4__2730_, data_stage_4__2729_, data_stage_4__2728_, data_stage_4__2727_, data_stage_4__2726_, data_stage_4__2725_, data_stage_4__2724_, data_stage_4__2723_, data_stage_4__2722_, data_stage_4__2721_, data_stage_4__2720_, data_stage_4__2719_, data_stage_4__2718_, data_stage_4__2717_, data_stage_4__2716_, data_stage_4__2715_, data_stage_4__2714_, data_stage_4__2713_, data_stage_4__2712_, data_stage_4__2711_, data_stage_4__2710_, data_stage_4__2709_, data_stage_4__2708_, data_stage_4__2707_, data_stage_4__2706_, data_stage_4__2705_, data_stage_4__2704_, data_stage_4__2703_, data_stage_4__2702_, data_stage_4__2701_, data_stage_4__2700_, data_stage_4__2699_, data_stage_4__2698_, data_stage_4__2697_, data_stage_4__2696_, data_stage_4__2695_, data_stage_4__2694_, data_stage_4__2693_, data_stage_4__2692_, data_stage_4__2691_, data_stage_4__2690_, data_stage_4__2689_, data_stage_4__2688_, data_stage_4__2687_, data_stage_4__2686_, data_stage_4__2685_, data_stage_4__2684_, data_stage_4__2683_, data_stage_4__2682_, data_stage_4__2681_, data_stage_4__2680_, data_stage_4__2679_, data_stage_4__2678_, data_stage_4__2677_, data_stage_4__2676_, data_stage_4__2675_, data_stage_4__2674_, data_stage_4__2673_, data_stage_4__2672_, data_stage_4__2671_, data_stage_4__2670_, data_stage_4__2669_, data_stage_4__2668_, data_stage_4__2667_, data_stage_4__2666_, data_stage_4__2665_, data_stage_4__2664_, data_stage_4__2663_, data_stage_4__2662_, data_stage_4__2661_, data_stage_4__2660_, data_stage_4__2659_, data_stage_4__2658_, data_stage_4__2657_, data_stage_4__2656_, data_stage_4__2655_, data_stage_4__2654_, data_stage_4__2653_, data_stage_4__2652_, data_stage_4__2651_, data_stage_4__2650_, data_stage_4__2649_, data_stage_4__2648_, data_stage_4__2647_, data_stage_4__2646_, data_stage_4__2645_, data_stage_4__2644_, data_stage_4__2643_, data_stage_4__2642_, data_stage_4__2641_, data_stage_4__2640_, data_stage_4__2639_, data_stage_4__2638_, data_stage_4__2637_, data_stage_4__2636_, data_stage_4__2635_, data_stage_4__2634_, data_stage_4__2633_, data_stage_4__2632_, data_stage_4__2631_, data_stage_4__2630_, data_stage_4__2629_, data_stage_4__2628_, data_stage_4__2627_, data_stage_4__2626_, data_stage_4__2625_, data_stage_4__2624_, data_stage_4__2623_, data_stage_4__2622_, data_stage_4__2621_, data_stage_4__2620_, data_stage_4__2619_, data_stage_4__2618_, data_stage_4__2617_, data_stage_4__2616_, data_stage_4__2615_, data_stage_4__2614_, data_stage_4__2613_, data_stage_4__2612_, data_stage_4__2611_, data_stage_4__2610_, data_stage_4__2609_, data_stage_4__2608_, data_stage_4__2607_, data_stage_4__2606_, data_stage_4__2605_, data_stage_4__2604_, data_stage_4__2603_, data_stage_4__2602_, data_stage_4__2601_, data_stage_4__2600_, data_stage_4__2599_, data_stage_4__2598_, data_stage_4__2597_, data_stage_4__2596_, data_stage_4__2595_, data_stage_4__2594_, data_stage_4__2593_, data_stage_4__2592_, data_stage_4__2591_, data_stage_4__2590_, data_stage_4__2589_, data_stage_4__2588_, data_stage_4__2587_, data_stage_4__2586_, data_stage_4__2585_, data_stage_4__2584_, data_stage_4__2583_, data_stage_4__2582_, data_stage_4__2581_, data_stage_4__2580_, data_stage_4__2579_, data_stage_4__2578_, data_stage_4__2577_, data_stage_4__2576_, data_stage_4__2575_, data_stage_4__2574_, data_stage_4__2573_, data_stage_4__2572_, data_stage_4__2571_, data_stage_4__2570_, data_stage_4__2569_, data_stage_4__2568_, data_stage_4__2567_, data_stage_4__2566_, data_stage_4__2565_, data_stage_4__2564_, data_stage_4__2563_, data_stage_4__2562_, data_stage_4__2561_, data_stage_4__2560_, data_stage_4__2559_, data_stage_4__2558_, data_stage_4__2557_, data_stage_4__2556_, data_stage_4__2555_, data_stage_4__2554_, data_stage_4__2553_, data_stage_4__2552_, data_stage_4__2551_, data_stage_4__2550_, data_stage_4__2549_, data_stage_4__2548_, data_stage_4__2547_, data_stage_4__2546_, data_stage_4__2545_, data_stage_4__2544_, data_stage_4__2543_, data_stage_4__2542_, data_stage_4__2541_, data_stage_4__2540_, data_stage_4__2539_, data_stage_4__2538_, data_stage_4__2537_, data_stage_4__2536_, data_stage_4__2535_, data_stage_4__2534_, data_stage_4__2533_, data_stage_4__2532_, data_stage_4__2531_, data_stage_4__2530_, data_stage_4__2529_, data_stage_4__2528_, data_stage_4__2527_, data_stage_4__2526_, data_stage_4__2525_, data_stage_4__2524_, data_stage_4__2523_, data_stage_4__2522_, data_stage_4__2521_, data_stage_4__2520_, data_stage_4__2519_, data_stage_4__2518_, data_stage_4__2517_, data_stage_4__2516_, data_stage_4__2515_, data_stage_4__2514_, data_stage_4__2513_, data_stage_4__2512_, data_stage_4__2511_, data_stage_4__2510_, data_stage_4__2509_, data_stage_4__2508_, data_stage_4__2507_, data_stage_4__2506_, data_stage_4__2505_, data_stage_4__2504_, data_stage_4__2503_, data_stage_4__2502_, data_stage_4__2501_, data_stage_4__2500_, data_stage_4__2499_, data_stage_4__2498_, data_stage_4__2497_, data_stage_4__2496_, data_stage_4__2495_, data_stage_4__2494_, data_stage_4__2493_, data_stage_4__2492_, data_stage_4__2491_, data_stage_4__2490_, data_stage_4__2489_, data_stage_4__2488_, data_stage_4__2487_, data_stage_4__2486_, data_stage_4__2485_, data_stage_4__2484_, data_stage_4__2483_, data_stage_4__2482_, data_stage_4__2481_, data_stage_4__2480_, data_stage_4__2479_, data_stage_4__2478_, data_stage_4__2477_, data_stage_4__2476_, data_stage_4__2475_, data_stage_4__2474_, data_stage_4__2473_, data_stage_4__2472_, data_stage_4__2471_, data_stage_4__2470_, data_stage_4__2469_, data_stage_4__2468_, data_stage_4__2467_, data_stage_4__2466_, data_stage_4__2465_, data_stage_4__2464_, data_stage_4__2463_, data_stage_4__2462_, data_stage_4__2461_, data_stage_4__2460_, data_stage_4__2459_, data_stage_4__2458_, data_stage_4__2457_, data_stage_4__2456_, data_stage_4__2455_, data_stage_4__2454_, data_stage_4__2453_, data_stage_4__2452_, data_stage_4__2451_, data_stage_4__2450_, data_stage_4__2449_, data_stage_4__2448_, data_stage_4__2447_, data_stage_4__2446_, data_stage_4__2445_, data_stage_4__2444_, data_stage_4__2443_, data_stage_4__2442_, data_stage_4__2441_, data_stage_4__2440_, data_stage_4__2439_, data_stage_4__2438_, data_stage_4__2437_, data_stage_4__2436_, data_stage_4__2435_, data_stage_4__2434_, data_stage_4__2433_, data_stage_4__2432_, data_stage_4__2431_, data_stage_4__2430_, data_stage_4__2429_, data_stage_4__2428_, data_stage_4__2427_, data_stage_4__2426_, data_stage_4__2425_, data_stage_4__2424_, data_stage_4__2423_, data_stage_4__2422_, data_stage_4__2421_, data_stage_4__2420_, data_stage_4__2419_, data_stage_4__2418_, data_stage_4__2417_, data_stage_4__2416_, data_stage_4__2415_, data_stage_4__2414_, data_stage_4__2413_, data_stage_4__2412_, data_stage_4__2411_, data_stage_4__2410_, data_stage_4__2409_, data_stage_4__2408_, data_stage_4__2407_, data_stage_4__2406_, data_stage_4__2405_, data_stage_4__2404_, data_stage_4__2403_, data_stage_4__2402_, data_stage_4__2401_, data_stage_4__2400_, data_stage_4__2399_, data_stage_4__2398_, data_stage_4__2397_, data_stage_4__2396_, data_stage_4__2395_, data_stage_4__2394_, data_stage_4__2393_, data_stage_4__2392_, data_stage_4__2391_, data_stage_4__2390_, data_stage_4__2389_, data_stage_4__2388_, data_stage_4__2387_, data_stage_4__2386_, data_stage_4__2385_, data_stage_4__2384_, data_stage_4__2383_, data_stage_4__2382_, data_stage_4__2381_, data_stage_4__2380_, data_stage_4__2379_, data_stage_4__2378_, data_stage_4__2377_, data_stage_4__2376_, data_stage_4__2375_, data_stage_4__2374_, data_stage_4__2373_, data_stage_4__2372_, data_stage_4__2371_, data_stage_4__2370_, data_stage_4__2369_, data_stage_4__2368_, data_stage_4__2367_, data_stage_4__2366_, data_stage_4__2365_, data_stage_4__2364_, data_stage_4__2363_, data_stage_4__2362_, data_stage_4__2361_, data_stage_4__2360_, data_stage_4__2359_, data_stage_4__2358_, data_stage_4__2357_, data_stage_4__2356_, data_stage_4__2355_, data_stage_4__2354_, data_stage_4__2353_, data_stage_4__2352_, data_stage_4__2351_, data_stage_4__2350_, data_stage_4__2349_, data_stage_4__2348_, data_stage_4__2347_, data_stage_4__2346_, data_stage_4__2345_, data_stage_4__2344_, data_stage_4__2343_, data_stage_4__2342_, data_stage_4__2341_, data_stage_4__2340_, data_stage_4__2339_, data_stage_4__2338_, data_stage_4__2337_, data_stage_4__2336_, data_stage_4__2335_, data_stage_4__2334_, data_stage_4__2333_, data_stage_4__2332_, data_stage_4__2331_, data_stage_4__2330_, data_stage_4__2329_, data_stage_4__2328_, data_stage_4__2327_, data_stage_4__2326_, data_stage_4__2325_, data_stage_4__2324_, data_stage_4__2323_, data_stage_4__2322_, data_stage_4__2321_, data_stage_4__2320_, data_stage_4__2319_, data_stage_4__2318_, data_stage_4__2317_, data_stage_4__2316_, data_stage_4__2315_, data_stage_4__2314_, data_stage_4__2313_, data_stage_4__2312_, data_stage_4__2311_, data_stage_4__2310_, data_stage_4__2309_, data_stage_4__2308_, data_stage_4__2307_, data_stage_4__2306_, data_stage_4__2305_, data_stage_4__2304_, data_stage_4__2303_, data_stage_4__2302_, data_stage_4__2301_, data_stage_4__2300_, data_stage_4__2299_, data_stage_4__2298_, data_stage_4__2297_, data_stage_4__2296_, data_stage_4__2295_, data_stage_4__2294_, data_stage_4__2293_, data_stage_4__2292_, data_stage_4__2291_, data_stage_4__2290_, data_stage_4__2289_, data_stage_4__2288_, data_stage_4__2287_, data_stage_4__2286_, data_stage_4__2285_, data_stage_4__2284_, data_stage_4__2283_, data_stage_4__2282_, data_stage_4__2281_, data_stage_4__2280_, data_stage_4__2279_, data_stage_4__2278_, data_stage_4__2277_, data_stage_4__2276_, data_stage_4__2275_, data_stage_4__2274_, data_stage_4__2273_, data_stage_4__2272_, data_stage_4__2271_, data_stage_4__2270_, data_stage_4__2269_, data_stage_4__2268_, data_stage_4__2267_, data_stage_4__2266_, data_stage_4__2265_, data_stage_4__2264_, data_stage_4__2263_, data_stage_4__2262_, data_stage_4__2261_, data_stage_4__2260_, data_stage_4__2259_, data_stage_4__2258_, data_stage_4__2257_, data_stage_4__2256_, data_stage_4__2255_, data_stage_4__2254_, data_stage_4__2253_, data_stage_4__2252_, data_stage_4__2251_, data_stage_4__2250_, data_stage_4__2249_, data_stage_4__2248_, data_stage_4__2247_, data_stage_4__2246_, data_stage_4__2245_, data_stage_4__2244_, data_stage_4__2243_, data_stage_4__2242_, data_stage_4__2241_, data_stage_4__2240_, data_stage_4__2239_, data_stage_4__2238_, data_stage_4__2237_, data_stage_4__2236_, data_stage_4__2235_, data_stage_4__2234_, data_stage_4__2233_, data_stage_4__2232_, data_stage_4__2231_, data_stage_4__2230_, data_stage_4__2229_, data_stage_4__2228_, data_stage_4__2227_, data_stage_4__2226_, data_stage_4__2225_, data_stage_4__2224_, data_stage_4__2223_, data_stage_4__2222_, data_stage_4__2221_, data_stage_4__2220_, data_stage_4__2219_, data_stage_4__2218_, data_stage_4__2217_, data_stage_4__2216_, data_stage_4__2215_, data_stage_4__2214_, data_stage_4__2213_, data_stage_4__2212_, data_stage_4__2211_, data_stage_4__2210_, data_stage_4__2209_, data_stage_4__2208_, data_stage_4__2207_, data_stage_4__2206_, data_stage_4__2205_, data_stage_4__2204_, data_stage_4__2203_, data_stage_4__2202_, data_stage_4__2201_, data_stage_4__2200_, data_stage_4__2199_, data_stage_4__2198_, data_stage_4__2197_, data_stage_4__2196_, data_stage_4__2195_, data_stage_4__2194_, data_stage_4__2193_, data_stage_4__2192_, data_stage_4__2191_, data_stage_4__2190_, data_stage_4__2189_, data_stage_4__2188_, data_stage_4__2187_, data_stage_4__2186_, data_stage_4__2185_, data_stage_4__2184_, data_stage_4__2183_, data_stage_4__2182_, data_stage_4__2181_, data_stage_4__2180_, data_stage_4__2179_, data_stage_4__2178_, data_stage_4__2177_, data_stage_4__2176_, data_stage_4__2175_, data_stage_4__2174_, data_stage_4__2173_, data_stage_4__2172_, data_stage_4__2171_, data_stage_4__2170_, data_stage_4__2169_, data_stage_4__2168_, data_stage_4__2167_, data_stage_4__2166_, data_stage_4__2165_, data_stage_4__2164_, data_stage_4__2163_, data_stage_4__2162_, data_stage_4__2161_, data_stage_4__2160_, data_stage_4__2159_, data_stage_4__2158_, data_stage_4__2157_, data_stage_4__2156_, data_stage_4__2155_, data_stage_4__2154_, data_stage_4__2153_, data_stage_4__2152_, data_stage_4__2151_, data_stage_4__2150_, data_stage_4__2149_, data_stage_4__2148_, data_stage_4__2147_, data_stage_4__2146_, data_stage_4__2145_, data_stage_4__2144_, data_stage_4__2143_, data_stage_4__2142_, data_stage_4__2141_, data_stage_4__2140_, data_stage_4__2139_, data_stage_4__2138_, data_stage_4__2137_, data_stage_4__2136_, data_stage_4__2135_, data_stage_4__2134_, data_stage_4__2133_, data_stage_4__2132_, data_stage_4__2131_, data_stage_4__2130_, data_stage_4__2129_, data_stage_4__2128_, data_stage_4__2127_, data_stage_4__2126_, data_stage_4__2125_, data_stage_4__2124_, data_stage_4__2123_, data_stage_4__2122_, data_stage_4__2121_, data_stage_4__2120_, data_stage_4__2119_, data_stage_4__2118_, data_stage_4__2117_, data_stage_4__2116_, data_stage_4__2115_, data_stage_4__2114_, data_stage_4__2113_, data_stage_4__2112_, data_stage_4__2111_, data_stage_4__2110_, data_stage_4__2109_, data_stage_4__2108_, data_stage_4__2107_, data_stage_4__2106_, data_stage_4__2105_, data_stage_4__2104_, data_stage_4__2103_, data_stage_4__2102_, data_stage_4__2101_, data_stage_4__2100_, data_stage_4__2099_, data_stage_4__2098_, data_stage_4__2097_, data_stage_4__2096_, data_stage_4__2095_, data_stage_4__2094_, data_stage_4__2093_, data_stage_4__2092_, data_stage_4__2091_, data_stage_4__2090_, data_stage_4__2089_, data_stage_4__2088_, data_stage_4__2087_, data_stage_4__2086_, data_stage_4__2085_, data_stage_4__2084_, data_stage_4__2083_, data_stage_4__2082_, data_stage_4__2081_, data_stage_4__2080_, data_stage_4__2079_, data_stage_4__2078_, data_stage_4__2077_, data_stage_4__2076_, data_stage_4__2075_, data_stage_4__2074_, data_stage_4__2073_, data_stage_4__2072_, data_stage_4__2071_, data_stage_4__2070_, data_stage_4__2069_, data_stage_4__2068_, data_stage_4__2067_, data_stage_4__2066_, data_stage_4__2065_, data_stage_4__2064_, data_stage_4__2063_, data_stage_4__2062_, data_stage_4__2061_, data_stage_4__2060_, data_stage_4__2059_, data_stage_4__2058_, data_stage_4__2057_, data_stage_4__2056_, data_stage_4__2055_, data_stage_4__2054_, data_stage_4__2053_, data_stage_4__2052_, data_stage_4__2051_, data_stage_4__2050_, data_stage_4__2049_, data_stage_4__2048_ })
  );


  bsg_swap_width_p1024
  mux_stage_3__mux_swap_2__swap_inst
  (
    .data_i({ data_stage_3__6143_, data_stage_3__6142_, data_stage_3__6141_, data_stage_3__6140_, data_stage_3__6139_, data_stage_3__6138_, data_stage_3__6137_, data_stage_3__6136_, data_stage_3__6135_, data_stage_3__6134_, data_stage_3__6133_, data_stage_3__6132_, data_stage_3__6131_, data_stage_3__6130_, data_stage_3__6129_, data_stage_3__6128_, data_stage_3__6127_, data_stage_3__6126_, data_stage_3__6125_, data_stage_3__6124_, data_stage_3__6123_, data_stage_3__6122_, data_stage_3__6121_, data_stage_3__6120_, data_stage_3__6119_, data_stage_3__6118_, data_stage_3__6117_, data_stage_3__6116_, data_stage_3__6115_, data_stage_3__6114_, data_stage_3__6113_, data_stage_3__6112_, data_stage_3__6111_, data_stage_3__6110_, data_stage_3__6109_, data_stage_3__6108_, data_stage_3__6107_, data_stage_3__6106_, data_stage_3__6105_, data_stage_3__6104_, data_stage_3__6103_, data_stage_3__6102_, data_stage_3__6101_, data_stage_3__6100_, data_stage_3__6099_, data_stage_3__6098_, data_stage_3__6097_, data_stage_3__6096_, data_stage_3__6095_, data_stage_3__6094_, data_stage_3__6093_, data_stage_3__6092_, data_stage_3__6091_, data_stage_3__6090_, data_stage_3__6089_, data_stage_3__6088_, data_stage_3__6087_, data_stage_3__6086_, data_stage_3__6085_, data_stage_3__6084_, data_stage_3__6083_, data_stage_3__6082_, data_stage_3__6081_, data_stage_3__6080_, data_stage_3__6079_, data_stage_3__6078_, data_stage_3__6077_, data_stage_3__6076_, data_stage_3__6075_, data_stage_3__6074_, data_stage_3__6073_, data_stage_3__6072_, data_stage_3__6071_, data_stage_3__6070_, data_stage_3__6069_, data_stage_3__6068_, data_stage_3__6067_, data_stage_3__6066_, data_stage_3__6065_, data_stage_3__6064_, data_stage_3__6063_, data_stage_3__6062_, data_stage_3__6061_, data_stage_3__6060_, data_stage_3__6059_, data_stage_3__6058_, data_stage_3__6057_, data_stage_3__6056_, data_stage_3__6055_, data_stage_3__6054_, data_stage_3__6053_, data_stage_3__6052_, data_stage_3__6051_, data_stage_3__6050_, data_stage_3__6049_, data_stage_3__6048_, data_stage_3__6047_, data_stage_3__6046_, data_stage_3__6045_, data_stage_3__6044_, data_stage_3__6043_, data_stage_3__6042_, data_stage_3__6041_, data_stage_3__6040_, data_stage_3__6039_, data_stage_3__6038_, data_stage_3__6037_, data_stage_3__6036_, data_stage_3__6035_, data_stage_3__6034_, data_stage_3__6033_, data_stage_3__6032_, data_stage_3__6031_, data_stage_3__6030_, data_stage_3__6029_, data_stage_3__6028_, data_stage_3__6027_, data_stage_3__6026_, data_stage_3__6025_, data_stage_3__6024_, data_stage_3__6023_, data_stage_3__6022_, data_stage_3__6021_, data_stage_3__6020_, data_stage_3__6019_, data_stage_3__6018_, data_stage_3__6017_, data_stage_3__6016_, data_stage_3__6015_, data_stage_3__6014_, data_stage_3__6013_, data_stage_3__6012_, data_stage_3__6011_, data_stage_3__6010_, data_stage_3__6009_, data_stage_3__6008_, data_stage_3__6007_, data_stage_3__6006_, data_stage_3__6005_, data_stage_3__6004_, data_stage_3__6003_, data_stage_3__6002_, data_stage_3__6001_, data_stage_3__6000_, data_stage_3__5999_, data_stage_3__5998_, data_stage_3__5997_, data_stage_3__5996_, data_stage_3__5995_, data_stage_3__5994_, data_stage_3__5993_, data_stage_3__5992_, data_stage_3__5991_, data_stage_3__5990_, data_stage_3__5989_, data_stage_3__5988_, data_stage_3__5987_, data_stage_3__5986_, data_stage_3__5985_, data_stage_3__5984_, data_stage_3__5983_, data_stage_3__5982_, data_stage_3__5981_, data_stage_3__5980_, data_stage_3__5979_, data_stage_3__5978_, data_stage_3__5977_, data_stage_3__5976_, data_stage_3__5975_, data_stage_3__5974_, data_stage_3__5973_, data_stage_3__5972_, data_stage_3__5971_, data_stage_3__5970_, data_stage_3__5969_, data_stage_3__5968_, data_stage_3__5967_, data_stage_3__5966_, data_stage_3__5965_, data_stage_3__5964_, data_stage_3__5963_, data_stage_3__5962_, data_stage_3__5961_, data_stage_3__5960_, data_stage_3__5959_, data_stage_3__5958_, data_stage_3__5957_, data_stage_3__5956_, data_stage_3__5955_, data_stage_3__5954_, data_stage_3__5953_, data_stage_3__5952_, data_stage_3__5951_, data_stage_3__5950_, data_stage_3__5949_, data_stage_3__5948_, data_stage_3__5947_, data_stage_3__5946_, data_stage_3__5945_, data_stage_3__5944_, data_stage_3__5943_, data_stage_3__5942_, data_stage_3__5941_, data_stage_3__5940_, data_stage_3__5939_, data_stage_3__5938_, data_stage_3__5937_, data_stage_3__5936_, data_stage_3__5935_, data_stage_3__5934_, data_stage_3__5933_, data_stage_3__5932_, data_stage_3__5931_, data_stage_3__5930_, data_stage_3__5929_, data_stage_3__5928_, data_stage_3__5927_, data_stage_3__5926_, data_stage_3__5925_, data_stage_3__5924_, data_stage_3__5923_, data_stage_3__5922_, data_stage_3__5921_, data_stage_3__5920_, data_stage_3__5919_, data_stage_3__5918_, data_stage_3__5917_, data_stage_3__5916_, data_stage_3__5915_, data_stage_3__5914_, data_stage_3__5913_, data_stage_3__5912_, data_stage_3__5911_, data_stage_3__5910_, data_stage_3__5909_, data_stage_3__5908_, data_stage_3__5907_, data_stage_3__5906_, data_stage_3__5905_, data_stage_3__5904_, data_stage_3__5903_, data_stage_3__5902_, data_stage_3__5901_, data_stage_3__5900_, data_stage_3__5899_, data_stage_3__5898_, data_stage_3__5897_, data_stage_3__5896_, data_stage_3__5895_, data_stage_3__5894_, data_stage_3__5893_, data_stage_3__5892_, data_stage_3__5891_, data_stage_3__5890_, data_stage_3__5889_, data_stage_3__5888_, data_stage_3__5887_, data_stage_3__5886_, data_stage_3__5885_, data_stage_3__5884_, data_stage_3__5883_, data_stage_3__5882_, data_stage_3__5881_, data_stage_3__5880_, data_stage_3__5879_, data_stage_3__5878_, data_stage_3__5877_, data_stage_3__5876_, data_stage_3__5875_, data_stage_3__5874_, data_stage_3__5873_, data_stage_3__5872_, data_stage_3__5871_, data_stage_3__5870_, data_stage_3__5869_, data_stage_3__5868_, data_stage_3__5867_, data_stage_3__5866_, data_stage_3__5865_, data_stage_3__5864_, data_stage_3__5863_, data_stage_3__5862_, data_stage_3__5861_, data_stage_3__5860_, data_stage_3__5859_, data_stage_3__5858_, data_stage_3__5857_, data_stage_3__5856_, data_stage_3__5855_, data_stage_3__5854_, data_stage_3__5853_, data_stage_3__5852_, data_stage_3__5851_, data_stage_3__5850_, data_stage_3__5849_, data_stage_3__5848_, data_stage_3__5847_, data_stage_3__5846_, data_stage_3__5845_, data_stage_3__5844_, data_stage_3__5843_, data_stage_3__5842_, data_stage_3__5841_, data_stage_3__5840_, data_stage_3__5839_, data_stage_3__5838_, data_stage_3__5837_, data_stage_3__5836_, data_stage_3__5835_, data_stage_3__5834_, data_stage_3__5833_, data_stage_3__5832_, data_stage_3__5831_, data_stage_3__5830_, data_stage_3__5829_, data_stage_3__5828_, data_stage_3__5827_, data_stage_3__5826_, data_stage_3__5825_, data_stage_3__5824_, data_stage_3__5823_, data_stage_3__5822_, data_stage_3__5821_, data_stage_3__5820_, data_stage_3__5819_, data_stage_3__5818_, data_stage_3__5817_, data_stage_3__5816_, data_stage_3__5815_, data_stage_3__5814_, data_stage_3__5813_, data_stage_3__5812_, data_stage_3__5811_, data_stage_3__5810_, data_stage_3__5809_, data_stage_3__5808_, data_stage_3__5807_, data_stage_3__5806_, data_stage_3__5805_, data_stage_3__5804_, data_stage_3__5803_, data_stage_3__5802_, data_stage_3__5801_, data_stage_3__5800_, data_stage_3__5799_, data_stage_3__5798_, data_stage_3__5797_, data_stage_3__5796_, data_stage_3__5795_, data_stage_3__5794_, data_stage_3__5793_, data_stage_3__5792_, data_stage_3__5791_, data_stage_3__5790_, data_stage_3__5789_, data_stage_3__5788_, data_stage_3__5787_, data_stage_3__5786_, data_stage_3__5785_, data_stage_3__5784_, data_stage_3__5783_, data_stage_3__5782_, data_stage_3__5781_, data_stage_3__5780_, data_stage_3__5779_, data_stage_3__5778_, data_stage_3__5777_, data_stage_3__5776_, data_stage_3__5775_, data_stage_3__5774_, data_stage_3__5773_, data_stage_3__5772_, data_stage_3__5771_, data_stage_3__5770_, data_stage_3__5769_, data_stage_3__5768_, data_stage_3__5767_, data_stage_3__5766_, data_stage_3__5765_, data_stage_3__5764_, data_stage_3__5763_, data_stage_3__5762_, data_stage_3__5761_, data_stage_3__5760_, data_stage_3__5759_, data_stage_3__5758_, data_stage_3__5757_, data_stage_3__5756_, data_stage_3__5755_, data_stage_3__5754_, data_stage_3__5753_, data_stage_3__5752_, data_stage_3__5751_, data_stage_3__5750_, data_stage_3__5749_, data_stage_3__5748_, data_stage_3__5747_, data_stage_3__5746_, data_stage_3__5745_, data_stage_3__5744_, data_stage_3__5743_, data_stage_3__5742_, data_stage_3__5741_, data_stage_3__5740_, data_stage_3__5739_, data_stage_3__5738_, data_stage_3__5737_, data_stage_3__5736_, data_stage_3__5735_, data_stage_3__5734_, data_stage_3__5733_, data_stage_3__5732_, data_stage_3__5731_, data_stage_3__5730_, data_stage_3__5729_, data_stage_3__5728_, data_stage_3__5727_, data_stage_3__5726_, data_stage_3__5725_, data_stage_3__5724_, data_stage_3__5723_, data_stage_3__5722_, data_stage_3__5721_, data_stage_3__5720_, data_stage_3__5719_, data_stage_3__5718_, data_stage_3__5717_, data_stage_3__5716_, data_stage_3__5715_, data_stage_3__5714_, data_stage_3__5713_, data_stage_3__5712_, data_stage_3__5711_, data_stage_3__5710_, data_stage_3__5709_, data_stage_3__5708_, data_stage_3__5707_, data_stage_3__5706_, data_stage_3__5705_, data_stage_3__5704_, data_stage_3__5703_, data_stage_3__5702_, data_stage_3__5701_, data_stage_3__5700_, data_stage_3__5699_, data_stage_3__5698_, data_stage_3__5697_, data_stage_3__5696_, data_stage_3__5695_, data_stage_3__5694_, data_stage_3__5693_, data_stage_3__5692_, data_stage_3__5691_, data_stage_3__5690_, data_stage_3__5689_, data_stage_3__5688_, data_stage_3__5687_, data_stage_3__5686_, data_stage_3__5685_, data_stage_3__5684_, data_stage_3__5683_, data_stage_3__5682_, data_stage_3__5681_, data_stage_3__5680_, data_stage_3__5679_, data_stage_3__5678_, data_stage_3__5677_, data_stage_3__5676_, data_stage_3__5675_, data_stage_3__5674_, data_stage_3__5673_, data_stage_3__5672_, data_stage_3__5671_, data_stage_3__5670_, data_stage_3__5669_, data_stage_3__5668_, data_stage_3__5667_, data_stage_3__5666_, data_stage_3__5665_, data_stage_3__5664_, data_stage_3__5663_, data_stage_3__5662_, data_stage_3__5661_, data_stage_3__5660_, data_stage_3__5659_, data_stage_3__5658_, data_stage_3__5657_, data_stage_3__5656_, data_stage_3__5655_, data_stage_3__5654_, data_stage_3__5653_, data_stage_3__5652_, data_stage_3__5651_, data_stage_3__5650_, data_stage_3__5649_, data_stage_3__5648_, data_stage_3__5647_, data_stage_3__5646_, data_stage_3__5645_, data_stage_3__5644_, data_stage_3__5643_, data_stage_3__5642_, data_stage_3__5641_, data_stage_3__5640_, data_stage_3__5639_, data_stage_3__5638_, data_stage_3__5637_, data_stage_3__5636_, data_stage_3__5635_, data_stage_3__5634_, data_stage_3__5633_, data_stage_3__5632_, data_stage_3__5631_, data_stage_3__5630_, data_stage_3__5629_, data_stage_3__5628_, data_stage_3__5627_, data_stage_3__5626_, data_stage_3__5625_, data_stage_3__5624_, data_stage_3__5623_, data_stage_3__5622_, data_stage_3__5621_, data_stage_3__5620_, data_stage_3__5619_, data_stage_3__5618_, data_stage_3__5617_, data_stage_3__5616_, data_stage_3__5615_, data_stage_3__5614_, data_stage_3__5613_, data_stage_3__5612_, data_stage_3__5611_, data_stage_3__5610_, data_stage_3__5609_, data_stage_3__5608_, data_stage_3__5607_, data_stage_3__5606_, data_stage_3__5605_, data_stage_3__5604_, data_stage_3__5603_, data_stage_3__5602_, data_stage_3__5601_, data_stage_3__5600_, data_stage_3__5599_, data_stage_3__5598_, data_stage_3__5597_, data_stage_3__5596_, data_stage_3__5595_, data_stage_3__5594_, data_stage_3__5593_, data_stage_3__5592_, data_stage_3__5591_, data_stage_3__5590_, data_stage_3__5589_, data_stage_3__5588_, data_stage_3__5587_, data_stage_3__5586_, data_stage_3__5585_, data_stage_3__5584_, data_stage_3__5583_, data_stage_3__5582_, data_stage_3__5581_, data_stage_3__5580_, data_stage_3__5579_, data_stage_3__5578_, data_stage_3__5577_, data_stage_3__5576_, data_stage_3__5575_, data_stage_3__5574_, data_stage_3__5573_, data_stage_3__5572_, data_stage_3__5571_, data_stage_3__5570_, data_stage_3__5569_, data_stage_3__5568_, data_stage_3__5567_, data_stage_3__5566_, data_stage_3__5565_, data_stage_3__5564_, data_stage_3__5563_, data_stage_3__5562_, data_stage_3__5561_, data_stage_3__5560_, data_stage_3__5559_, data_stage_3__5558_, data_stage_3__5557_, data_stage_3__5556_, data_stage_3__5555_, data_stage_3__5554_, data_stage_3__5553_, data_stage_3__5552_, data_stage_3__5551_, data_stage_3__5550_, data_stage_3__5549_, data_stage_3__5548_, data_stage_3__5547_, data_stage_3__5546_, data_stage_3__5545_, data_stage_3__5544_, data_stage_3__5543_, data_stage_3__5542_, data_stage_3__5541_, data_stage_3__5540_, data_stage_3__5539_, data_stage_3__5538_, data_stage_3__5537_, data_stage_3__5536_, data_stage_3__5535_, data_stage_3__5534_, data_stage_3__5533_, data_stage_3__5532_, data_stage_3__5531_, data_stage_3__5530_, data_stage_3__5529_, data_stage_3__5528_, data_stage_3__5527_, data_stage_3__5526_, data_stage_3__5525_, data_stage_3__5524_, data_stage_3__5523_, data_stage_3__5522_, data_stage_3__5521_, data_stage_3__5520_, data_stage_3__5519_, data_stage_3__5518_, data_stage_3__5517_, data_stage_3__5516_, data_stage_3__5515_, data_stage_3__5514_, data_stage_3__5513_, data_stage_3__5512_, data_stage_3__5511_, data_stage_3__5510_, data_stage_3__5509_, data_stage_3__5508_, data_stage_3__5507_, data_stage_3__5506_, data_stage_3__5505_, data_stage_3__5504_, data_stage_3__5503_, data_stage_3__5502_, data_stage_3__5501_, data_stage_3__5500_, data_stage_3__5499_, data_stage_3__5498_, data_stage_3__5497_, data_stage_3__5496_, data_stage_3__5495_, data_stage_3__5494_, data_stage_3__5493_, data_stage_3__5492_, data_stage_3__5491_, data_stage_3__5490_, data_stage_3__5489_, data_stage_3__5488_, data_stage_3__5487_, data_stage_3__5486_, data_stage_3__5485_, data_stage_3__5484_, data_stage_3__5483_, data_stage_3__5482_, data_stage_3__5481_, data_stage_3__5480_, data_stage_3__5479_, data_stage_3__5478_, data_stage_3__5477_, data_stage_3__5476_, data_stage_3__5475_, data_stage_3__5474_, data_stage_3__5473_, data_stage_3__5472_, data_stage_3__5471_, data_stage_3__5470_, data_stage_3__5469_, data_stage_3__5468_, data_stage_3__5467_, data_stage_3__5466_, data_stage_3__5465_, data_stage_3__5464_, data_stage_3__5463_, data_stage_3__5462_, data_stage_3__5461_, data_stage_3__5460_, data_stage_3__5459_, data_stage_3__5458_, data_stage_3__5457_, data_stage_3__5456_, data_stage_3__5455_, data_stage_3__5454_, data_stage_3__5453_, data_stage_3__5452_, data_stage_3__5451_, data_stage_3__5450_, data_stage_3__5449_, data_stage_3__5448_, data_stage_3__5447_, data_stage_3__5446_, data_stage_3__5445_, data_stage_3__5444_, data_stage_3__5443_, data_stage_3__5442_, data_stage_3__5441_, data_stage_3__5440_, data_stage_3__5439_, data_stage_3__5438_, data_stage_3__5437_, data_stage_3__5436_, data_stage_3__5435_, data_stage_3__5434_, data_stage_3__5433_, data_stage_3__5432_, data_stage_3__5431_, data_stage_3__5430_, data_stage_3__5429_, data_stage_3__5428_, data_stage_3__5427_, data_stage_3__5426_, data_stage_3__5425_, data_stage_3__5424_, data_stage_3__5423_, data_stage_3__5422_, data_stage_3__5421_, data_stage_3__5420_, data_stage_3__5419_, data_stage_3__5418_, data_stage_3__5417_, data_stage_3__5416_, data_stage_3__5415_, data_stage_3__5414_, data_stage_3__5413_, data_stage_3__5412_, data_stage_3__5411_, data_stage_3__5410_, data_stage_3__5409_, data_stage_3__5408_, data_stage_3__5407_, data_stage_3__5406_, data_stage_3__5405_, data_stage_3__5404_, data_stage_3__5403_, data_stage_3__5402_, data_stage_3__5401_, data_stage_3__5400_, data_stage_3__5399_, data_stage_3__5398_, data_stage_3__5397_, data_stage_3__5396_, data_stage_3__5395_, data_stage_3__5394_, data_stage_3__5393_, data_stage_3__5392_, data_stage_3__5391_, data_stage_3__5390_, data_stage_3__5389_, data_stage_3__5388_, data_stage_3__5387_, data_stage_3__5386_, data_stage_3__5385_, data_stage_3__5384_, data_stage_3__5383_, data_stage_3__5382_, data_stage_3__5381_, data_stage_3__5380_, data_stage_3__5379_, data_stage_3__5378_, data_stage_3__5377_, data_stage_3__5376_, data_stage_3__5375_, data_stage_3__5374_, data_stage_3__5373_, data_stage_3__5372_, data_stage_3__5371_, data_stage_3__5370_, data_stage_3__5369_, data_stage_3__5368_, data_stage_3__5367_, data_stage_3__5366_, data_stage_3__5365_, data_stage_3__5364_, data_stage_3__5363_, data_stage_3__5362_, data_stage_3__5361_, data_stage_3__5360_, data_stage_3__5359_, data_stage_3__5358_, data_stage_3__5357_, data_stage_3__5356_, data_stage_3__5355_, data_stage_3__5354_, data_stage_3__5353_, data_stage_3__5352_, data_stage_3__5351_, data_stage_3__5350_, data_stage_3__5349_, data_stage_3__5348_, data_stage_3__5347_, data_stage_3__5346_, data_stage_3__5345_, data_stage_3__5344_, data_stage_3__5343_, data_stage_3__5342_, data_stage_3__5341_, data_stage_3__5340_, data_stage_3__5339_, data_stage_3__5338_, data_stage_3__5337_, data_stage_3__5336_, data_stage_3__5335_, data_stage_3__5334_, data_stage_3__5333_, data_stage_3__5332_, data_stage_3__5331_, data_stage_3__5330_, data_stage_3__5329_, data_stage_3__5328_, data_stage_3__5327_, data_stage_3__5326_, data_stage_3__5325_, data_stage_3__5324_, data_stage_3__5323_, data_stage_3__5322_, data_stage_3__5321_, data_stage_3__5320_, data_stage_3__5319_, data_stage_3__5318_, data_stage_3__5317_, data_stage_3__5316_, data_stage_3__5315_, data_stage_3__5314_, data_stage_3__5313_, data_stage_3__5312_, data_stage_3__5311_, data_stage_3__5310_, data_stage_3__5309_, data_stage_3__5308_, data_stage_3__5307_, data_stage_3__5306_, data_stage_3__5305_, data_stage_3__5304_, data_stage_3__5303_, data_stage_3__5302_, data_stage_3__5301_, data_stage_3__5300_, data_stage_3__5299_, data_stage_3__5298_, data_stage_3__5297_, data_stage_3__5296_, data_stage_3__5295_, data_stage_3__5294_, data_stage_3__5293_, data_stage_3__5292_, data_stage_3__5291_, data_stage_3__5290_, data_stage_3__5289_, data_stage_3__5288_, data_stage_3__5287_, data_stage_3__5286_, data_stage_3__5285_, data_stage_3__5284_, data_stage_3__5283_, data_stage_3__5282_, data_stage_3__5281_, data_stage_3__5280_, data_stage_3__5279_, data_stage_3__5278_, data_stage_3__5277_, data_stage_3__5276_, data_stage_3__5275_, data_stage_3__5274_, data_stage_3__5273_, data_stage_3__5272_, data_stage_3__5271_, data_stage_3__5270_, data_stage_3__5269_, data_stage_3__5268_, data_stage_3__5267_, data_stage_3__5266_, data_stage_3__5265_, data_stage_3__5264_, data_stage_3__5263_, data_stage_3__5262_, data_stage_3__5261_, data_stage_3__5260_, data_stage_3__5259_, data_stage_3__5258_, data_stage_3__5257_, data_stage_3__5256_, data_stage_3__5255_, data_stage_3__5254_, data_stage_3__5253_, data_stage_3__5252_, data_stage_3__5251_, data_stage_3__5250_, data_stage_3__5249_, data_stage_3__5248_, data_stage_3__5247_, data_stage_3__5246_, data_stage_3__5245_, data_stage_3__5244_, data_stage_3__5243_, data_stage_3__5242_, data_stage_3__5241_, data_stage_3__5240_, data_stage_3__5239_, data_stage_3__5238_, data_stage_3__5237_, data_stage_3__5236_, data_stage_3__5235_, data_stage_3__5234_, data_stage_3__5233_, data_stage_3__5232_, data_stage_3__5231_, data_stage_3__5230_, data_stage_3__5229_, data_stage_3__5228_, data_stage_3__5227_, data_stage_3__5226_, data_stage_3__5225_, data_stage_3__5224_, data_stage_3__5223_, data_stage_3__5222_, data_stage_3__5221_, data_stage_3__5220_, data_stage_3__5219_, data_stage_3__5218_, data_stage_3__5217_, data_stage_3__5216_, data_stage_3__5215_, data_stage_3__5214_, data_stage_3__5213_, data_stage_3__5212_, data_stage_3__5211_, data_stage_3__5210_, data_stage_3__5209_, data_stage_3__5208_, data_stage_3__5207_, data_stage_3__5206_, data_stage_3__5205_, data_stage_3__5204_, data_stage_3__5203_, data_stage_3__5202_, data_stage_3__5201_, data_stage_3__5200_, data_stage_3__5199_, data_stage_3__5198_, data_stage_3__5197_, data_stage_3__5196_, data_stage_3__5195_, data_stage_3__5194_, data_stage_3__5193_, data_stage_3__5192_, data_stage_3__5191_, data_stage_3__5190_, data_stage_3__5189_, data_stage_3__5188_, data_stage_3__5187_, data_stage_3__5186_, data_stage_3__5185_, data_stage_3__5184_, data_stage_3__5183_, data_stage_3__5182_, data_stage_3__5181_, data_stage_3__5180_, data_stage_3__5179_, data_stage_3__5178_, data_stage_3__5177_, data_stage_3__5176_, data_stage_3__5175_, data_stage_3__5174_, data_stage_3__5173_, data_stage_3__5172_, data_stage_3__5171_, data_stage_3__5170_, data_stage_3__5169_, data_stage_3__5168_, data_stage_3__5167_, data_stage_3__5166_, data_stage_3__5165_, data_stage_3__5164_, data_stage_3__5163_, data_stage_3__5162_, data_stage_3__5161_, data_stage_3__5160_, data_stage_3__5159_, data_stage_3__5158_, data_stage_3__5157_, data_stage_3__5156_, data_stage_3__5155_, data_stage_3__5154_, data_stage_3__5153_, data_stage_3__5152_, data_stage_3__5151_, data_stage_3__5150_, data_stage_3__5149_, data_stage_3__5148_, data_stage_3__5147_, data_stage_3__5146_, data_stage_3__5145_, data_stage_3__5144_, data_stage_3__5143_, data_stage_3__5142_, data_stage_3__5141_, data_stage_3__5140_, data_stage_3__5139_, data_stage_3__5138_, data_stage_3__5137_, data_stage_3__5136_, data_stage_3__5135_, data_stage_3__5134_, data_stage_3__5133_, data_stage_3__5132_, data_stage_3__5131_, data_stage_3__5130_, data_stage_3__5129_, data_stage_3__5128_, data_stage_3__5127_, data_stage_3__5126_, data_stage_3__5125_, data_stage_3__5124_, data_stage_3__5123_, data_stage_3__5122_, data_stage_3__5121_, data_stage_3__5120_, data_stage_3__5119_, data_stage_3__5118_, data_stage_3__5117_, data_stage_3__5116_, data_stage_3__5115_, data_stage_3__5114_, data_stage_3__5113_, data_stage_3__5112_, data_stage_3__5111_, data_stage_3__5110_, data_stage_3__5109_, data_stage_3__5108_, data_stage_3__5107_, data_stage_3__5106_, data_stage_3__5105_, data_stage_3__5104_, data_stage_3__5103_, data_stage_3__5102_, data_stage_3__5101_, data_stage_3__5100_, data_stage_3__5099_, data_stage_3__5098_, data_stage_3__5097_, data_stage_3__5096_, data_stage_3__5095_, data_stage_3__5094_, data_stage_3__5093_, data_stage_3__5092_, data_stage_3__5091_, data_stage_3__5090_, data_stage_3__5089_, data_stage_3__5088_, data_stage_3__5087_, data_stage_3__5086_, data_stage_3__5085_, data_stage_3__5084_, data_stage_3__5083_, data_stage_3__5082_, data_stage_3__5081_, data_stage_3__5080_, data_stage_3__5079_, data_stage_3__5078_, data_stage_3__5077_, data_stage_3__5076_, data_stage_3__5075_, data_stage_3__5074_, data_stage_3__5073_, data_stage_3__5072_, data_stage_3__5071_, data_stage_3__5070_, data_stage_3__5069_, data_stage_3__5068_, data_stage_3__5067_, data_stage_3__5066_, data_stage_3__5065_, data_stage_3__5064_, data_stage_3__5063_, data_stage_3__5062_, data_stage_3__5061_, data_stage_3__5060_, data_stage_3__5059_, data_stage_3__5058_, data_stage_3__5057_, data_stage_3__5056_, data_stage_3__5055_, data_stage_3__5054_, data_stage_3__5053_, data_stage_3__5052_, data_stage_3__5051_, data_stage_3__5050_, data_stage_3__5049_, data_stage_3__5048_, data_stage_3__5047_, data_stage_3__5046_, data_stage_3__5045_, data_stage_3__5044_, data_stage_3__5043_, data_stage_3__5042_, data_stage_3__5041_, data_stage_3__5040_, data_stage_3__5039_, data_stage_3__5038_, data_stage_3__5037_, data_stage_3__5036_, data_stage_3__5035_, data_stage_3__5034_, data_stage_3__5033_, data_stage_3__5032_, data_stage_3__5031_, data_stage_3__5030_, data_stage_3__5029_, data_stage_3__5028_, data_stage_3__5027_, data_stage_3__5026_, data_stage_3__5025_, data_stage_3__5024_, data_stage_3__5023_, data_stage_3__5022_, data_stage_3__5021_, data_stage_3__5020_, data_stage_3__5019_, data_stage_3__5018_, data_stage_3__5017_, data_stage_3__5016_, data_stage_3__5015_, data_stage_3__5014_, data_stage_3__5013_, data_stage_3__5012_, data_stage_3__5011_, data_stage_3__5010_, data_stage_3__5009_, data_stage_3__5008_, data_stage_3__5007_, data_stage_3__5006_, data_stage_3__5005_, data_stage_3__5004_, data_stage_3__5003_, data_stage_3__5002_, data_stage_3__5001_, data_stage_3__5000_, data_stage_3__4999_, data_stage_3__4998_, data_stage_3__4997_, data_stage_3__4996_, data_stage_3__4995_, data_stage_3__4994_, data_stage_3__4993_, data_stage_3__4992_, data_stage_3__4991_, data_stage_3__4990_, data_stage_3__4989_, data_stage_3__4988_, data_stage_3__4987_, data_stage_3__4986_, data_stage_3__4985_, data_stage_3__4984_, data_stage_3__4983_, data_stage_3__4982_, data_stage_3__4981_, data_stage_3__4980_, data_stage_3__4979_, data_stage_3__4978_, data_stage_3__4977_, data_stage_3__4976_, data_stage_3__4975_, data_stage_3__4974_, data_stage_3__4973_, data_stage_3__4972_, data_stage_3__4971_, data_stage_3__4970_, data_stage_3__4969_, data_stage_3__4968_, data_stage_3__4967_, data_stage_3__4966_, data_stage_3__4965_, data_stage_3__4964_, data_stage_3__4963_, data_stage_3__4962_, data_stage_3__4961_, data_stage_3__4960_, data_stage_3__4959_, data_stage_3__4958_, data_stage_3__4957_, data_stage_3__4956_, data_stage_3__4955_, data_stage_3__4954_, data_stage_3__4953_, data_stage_3__4952_, data_stage_3__4951_, data_stage_3__4950_, data_stage_3__4949_, data_stage_3__4948_, data_stage_3__4947_, data_stage_3__4946_, data_stage_3__4945_, data_stage_3__4944_, data_stage_3__4943_, data_stage_3__4942_, data_stage_3__4941_, data_stage_3__4940_, data_stage_3__4939_, data_stage_3__4938_, data_stage_3__4937_, data_stage_3__4936_, data_stage_3__4935_, data_stage_3__4934_, data_stage_3__4933_, data_stage_3__4932_, data_stage_3__4931_, data_stage_3__4930_, data_stage_3__4929_, data_stage_3__4928_, data_stage_3__4927_, data_stage_3__4926_, data_stage_3__4925_, data_stage_3__4924_, data_stage_3__4923_, data_stage_3__4922_, data_stage_3__4921_, data_stage_3__4920_, data_stage_3__4919_, data_stage_3__4918_, data_stage_3__4917_, data_stage_3__4916_, data_stage_3__4915_, data_stage_3__4914_, data_stage_3__4913_, data_stage_3__4912_, data_stage_3__4911_, data_stage_3__4910_, data_stage_3__4909_, data_stage_3__4908_, data_stage_3__4907_, data_stage_3__4906_, data_stage_3__4905_, data_stage_3__4904_, data_stage_3__4903_, data_stage_3__4902_, data_stage_3__4901_, data_stage_3__4900_, data_stage_3__4899_, data_stage_3__4898_, data_stage_3__4897_, data_stage_3__4896_, data_stage_3__4895_, data_stage_3__4894_, data_stage_3__4893_, data_stage_3__4892_, data_stage_3__4891_, data_stage_3__4890_, data_stage_3__4889_, data_stage_3__4888_, data_stage_3__4887_, data_stage_3__4886_, data_stage_3__4885_, data_stage_3__4884_, data_stage_3__4883_, data_stage_3__4882_, data_stage_3__4881_, data_stage_3__4880_, data_stage_3__4879_, data_stage_3__4878_, data_stage_3__4877_, data_stage_3__4876_, data_stage_3__4875_, data_stage_3__4874_, data_stage_3__4873_, data_stage_3__4872_, data_stage_3__4871_, data_stage_3__4870_, data_stage_3__4869_, data_stage_3__4868_, data_stage_3__4867_, data_stage_3__4866_, data_stage_3__4865_, data_stage_3__4864_, data_stage_3__4863_, data_stage_3__4862_, data_stage_3__4861_, data_stage_3__4860_, data_stage_3__4859_, data_stage_3__4858_, data_stage_3__4857_, data_stage_3__4856_, data_stage_3__4855_, data_stage_3__4854_, data_stage_3__4853_, data_stage_3__4852_, data_stage_3__4851_, data_stage_3__4850_, data_stage_3__4849_, data_stage_3__4848_, data_stage_3__4847_, data_stage_3__4846_, data_stage_3__4845_, data_stage_3__4844_, data_stage_3__4843_, data_stage_3__4842_, data_stage_3__4841_, data_stage_3__4840_, data_stage_3__4839_, data_stage_3__4838_, data_stage_3__4837_, data_stage_3__4836_, data_stage_3__4835_, data_stage_3__4834_, data_stage_3__4833_, data_stage_3__4832_, data_stage_3__4831_, data_stage_3__4830_, data_stage_3__4829_, data_stage_3__4828_, data_stage_3__4827_, data_stage_3__4826_, data_stage_3__4825_, data_stage_3__4824_, data_stage_3__4823_, data_stage_3__4822_, data_stage_3__4821_, data_stage_3__4820_, data_stage_3__4819_, data_stage_3__4818_, data_stage_3__4817_, data_stage_3__4816_, data_stage_3__4815_, data_stage_3__4814_, data_stage_3__4813_, data_stage_3__4812_, data_stage_3__4811_, data_stage_3__4810_, data_stage_3__4809_, data_stage_3__4808_, data_stage_3__4807_, data_stage_3__4806_, data_stage_3__4805_, data_stage_3__4804_, data_stage_3__4803_, data_stage_3__4802_, data_stage_3__4801_, data_stage_3__4800_, data_stage_3__4799_, data_stage_3__4798_, data_stage_3__4797_, data_stage_3__4796_, data_stage_3__4795_, data_stage_3__4794_, data_stage_3__4793_, data_stage_3__4792_, data_stage_3__4791_, data_stage_3__4790_, data_stage_3__4789_, data_stage_3__4788_, data_stage_3__4787_, data_stage_3__4786_, data_stage_3__4785_, data_stage_3__4784_, data_stage_3__4783_, data_stage_3__4782_, data_stage_3__4781_, data_stage_3__4780_, data_stage_3__4779_, data_stage_3__4778_, data_stage_3__4777_, data_stage_3__4776_, data_stage_3__4775_, data_stage_3__4774_, data_stage_3__4773_, data_stage_3__4772_, data_stage_3__4771_, data_stage_3__4770_, data_stage_3__4769_, data_stage_3__4768_, data_stage_3__4767_, data_stage_3__4766_, data_stage_3__4765_, data_stage_3__4764_, data_stage_3__4763_, data_stage_3__4762_, data_stage_3__4761_, data_stage_3__4760_, data_stage_3__4759_, data_stage_3__4758_, data_stage_3__4757_, data_stage_3__4756_, data_stage_3__4755_, data_stage_3__4754_, data_stage_3__4753_, data_stage_3__4752_, data_stage_3__4751_, data_stage_3__4750_, data_stage_3__4749_, data_stage_3__4748_, data_stage_3__4747_, data_stage_3__4746_, data_stage_3__4745_, data_stage_3__4744_, data_stage_3__4743_, data_stage_3__4742_, data_stage_3__4741_, data_stage_3__4740_, data_stage_3__4739_, data_stage_3__4738_, data_stage_3__4737_, data_stage_3__4736_, data_stage_3__4735_, data_stage_3__4734_, data_stage_3__4733_, data_stage_3__4732_, data_stage_3__4731_, data_stage_3__4730_, data_stage_3__4729_, data_stage_3__4728_, data_stage_3__4727_, data_stage_3__4726_, data_stage_3__4725_, data_stage_3__4724_, data_stage_3__4723_, data_stage_3__4722_, data_stage_3__4721_, data_stage_3__4720_, data_stage_3__4719_, data_stage_3__4718_, data_stage_3__4717_, data_stage_3__4716_, data_stage_3__4715_, data_stage_3__4714_, data_stage_3__4713_, data_stage_3__4712_, data_stage_3__4711_, data_stage_3__4710_, data_stage_3__4709_, data_stage_3__4708_, data_stage_3__4707_, data_stage_3__4706_, data_stage_3__4705_, data_stage_3__4704_, data_stage_3__4703_, data_stage_3__4702_, data_stage_3__4701_, data_stage_3__4700_, data_stage_3__4699_, data_stage_3__4698_, data_stage_3__4697_, data_stage_3__4696_, data_stage_3__4695_, data_stage_3__4694_, data_stage_3__4693_, data_stage_3__4692_, data_stage_3__4691_, data_stage_3__4690_, data_stage_3__4689_, data_stage_3__4688_, data_stage_3__4687_, data_stage_3__4686_, data_stage_3__4685_, data_stage_3__4684_, data_stage_3__4683_, data_stage_3__4682_, data_stage_3__4681_, data_stage_3__4680_, data_stage_3__4679_, data_stage_3__4678_, data_stage_3__4677_, data_stage_3__4676_, data_stage_3__4675_, data_stage_3__4674_, data_stage_3__4673_, data_stage_3__4672_, data_stage_3__4671_, data_stage_3__4670_, data_stage_3__4669_, data_stage_3__4668_, data_stage_3__4667_, data_stage_3__4666_, data_stage_3__4665_, data_stage_3__4664_, data_stage_3__4663_, data_stage_3__4662_, data_stage_3__4661_, data_stage_3__4660_, data_stage_3__4659_, data_stage_3__4658_, data_stage_3__4657_, data_stage_3__4656_, data_stage_3__4655_, data_stage_3__4654_, data_stage_3__4653_, data_stage_3__4652_, data_stage_3__4651_, data_stage_3__4650_, data_stage_3__4649_, data_stage_3__4648_, data_stage_3__4647_, data_stage_3__4646_, data_stage_3__4645_, data_stage_3__4644_, data_stage_3__4643_, data_stage_3__4642_, data_stage_3__4641_, data_stage_3__4640_, data_stage_3__4639_, data_stage_3__4638_, data_stage_3__4637_, data_stage_3__4636_, data_stage_3__4635_, data_stage_3__4634_, data_stage_3__4633_, data_stage_3__4632_, data_stage_3__4631_, data_stage_3__4630_, data_stage_3__4629_, data_stage_3__4628_, data_stage_3__4627_, data_stage_3__4626_, data_stage_3__4625_, data_stage_3__4624_, data_stage_3__4623_, data_stage_3__4622_, data_stage_3__4621_, data_stage_3__4620_, data_stage_3__4619_, data_stage_3__4618_, data_stage_3__4617_, data_stage_3__4616_, data_stage_3__4615_, data_stage_3__4614_, data_stage_3__4613_, data_stage_3__4612_, data_stage_3__4611_, data_stage_3__4610_, data_stage_3__4609_, data_stage_3__4608_, data_stage_3__4607_, data_stage_3__4606_, data_stage_3__4605_, data_stage_3__4604_, data_stage_3__4603_, data_stage_3__4602_, data_stage_3__4601_, data_stage_3__4600_, data_stage_3__4599_, data_stage_3__4598_, data_stage_3__4597_, data_stage_3__4596_, data_stage_3__4595_, data_stage_3__4594_, data_stage_3__4593_, data_stage_3__4592_, data_stage_3__4591_, data_stage_3__4590_, data_stage_3__4589_, data_stage_3__4588_, data_stage_3__4587_, data_stage_3__4586_, data_stage_3__4585_, data_stage_3__4584_, data_stage_3__4583_, data_stage_3__4582_, data_stage_3__4581_, data_stage_3__4580_, data_stage_3__4579_, data_stage_3__4578_, data_stage_3__4577_, data_stage_3__4576_, data_stage_3__4575_, data_stage_3__4574_, data_stage_3__4573_, data_stage_3__4572_, data_stage_3__4571_, data_stage_3__4570_, data_stage_3__4569_, data_stage_3__4568_, data_stage_3__4567_, data_stage_3__4566_, data_stage_3__4565_, data_stage_3__4564_, data_stage_3__4563_, data_stage_3__4562_, data_stage_3__4561_, data_stage_3__4560_, data_stage_3__4559_, data_stage_3__4558_, data_stage_3__4557_, data_stage_3__4556_, data_stage_3__4555_, data_stage_3__4554_, data_stage_3__4553_, data_stage_3__4552_, data_stage_3__4551_, data_stage_3__4550_, data_stage_3__4549_, data_stage_3__4548_, data_stage_3__4547_, data_stage_3__4546_, data_stage_3__4545_, data_stage_3__4544_, data_stage_3__4543_, data_stage_3__4542_, data_stage_3__4541_, data_stage_3__4540_, data_stage_3__4539_, data_stage_3__4538_, data_stage_3__4537_, data_stage_3__4536_, data_stage_3__4535_, data_stage_3__4534_, data_stage_3__4533_, data_stage_3__4532_, data_stage_3__4531_, data_stage_3__4530_, data_stage_3__4529_, data_stage_3__4528_, data_stage_3__4527_, data_stage_3__4526_, data_stage_3__4525_, data_stage_3__4524_, data_stage_3__4523_, data_stage_3__4522_, data_stage_3__4521_, data_stage_3__4520_, data_stage_3__4519_, data_stage_3__4518_, data_stage_3__4517_, data_stage_3__4516_, data_stage_3__4515_, data_stage_3__4514_, data_stage_3__4513_, data_stage_3__4512_, data_stage_3__4511_, data_stage_3__4510_, data_stage_3__4509_, data_stage_3__4508_, data_stage_3__4507_, data_stage_3__4506_, data_stage_3__4505_, data_stage_3__4504_, data_stage_3__4503_, data_stage_3__4502_, data_stage_3__4501_, data_stage_3__4500_, data_stage_3__4499_, data_stage_3__4498_, data_stage_3__4497_, data_stage_3__4496_, data_stage_3__4495_, data_stage_3__4494_, data_stage_3__4493_, data_stage_3__4492_, data_stage_3__4491_, data_stage_3__4490_, data_stage_3__4489_, data_stage_3__4488_, data_stage_3__4487_, data_stage_3__4486_, data_stage_3__4485_, data_stage_3__4484_, data_stage_3__4483_, data_stage_3__4482_, data_stage_3__4481_, data_stage_3__4480_, data_stage_3__4479_, data_stage_3__4478_, data_stage_3__4477_, data_stage_3__4476_, data_stage_3__4475_, data_stage_3__4474_, data_stage_3__4473_, data_stage_3__4472_, data_stage_3__4471_, data_stage_3__4470_, data_stage_3__4469_, data_stage_3__4468_, data_stage_3__4467_, data_stage_3__4466_, data_stage_3__4465_, data_stage_3__4464_, data_stage_3__4463_, data_stage_3__4462_, data_stage_3__4461_, data_stage_3__4460_, data_stage_3__4459_, data_stage_3__4458_, data_stage_3__4457_, data_stage_3__4456_, data_stage_3__4455_, data_stage_3__4454_, data_stage_3__4453_, data_stage_3__4452_, data_stage_3__4451_, data_stage_3__4450_, data_stage_3__4449_, data_stage_3__4448_, data_stage_3__4447_, data_stage_3__4446_, data_stage_3__4445_, data_stage_3__4444_, data_stage_3__4443_, data_stage_3__4442_, data_stage_3__4441_, data_stage_3__4440_, data_stage_3__4439_, data_stage_3__4438_, data_stage_3__4437_, data_stage_3__4436_, data_stage_3__4435_, data_stage_3__4434_, data_stage_3__4433_, data_stage_3__4432_, data_stage_3__4431_, data_stage_3__4430_, data_stage_3__4429_, data_stage_3__4428_, data_stage_3__4427_, data_stage_3__4426_, data_stage_3__4425_, data_stage_3__4424_, data_stage_3__4423_, data_stage_3__4422_, data_stage_3__4421_, data_stage_3__4420_, data_stage_3__4419_, data_stage_3__4418_, data_stage_3__4417_, data_stage_3__4416_, data_stage_3__4415_, data_stage_3__4414_, data_stage_3__4413_, data_stage_3__4412_, data_stage_3__4411_, data_stage_3__4410_, data_stage_3__4409_, data_stage_3__4408_, data_stage_3__4407_, data_stage_3__4406_, data_stage_3__4405_, data_stage_3__4404_, data_stage_3__4403_, data_stage_3__4402_, data_stage_3__4401_, data_stage_3__4400_, data_stage_3__4399_, data_stage_3__4398_, data_stage_3__4397_, data_stage_3__4396_, data_stage_3__4395_, data_stage_3__4394_, data_stage_3__4393_, data_stage_3__4392_, data_stage_3__4391_, data_stage_3__4390_, data_stage_3__4389_, data_stage_3__4388_, data_stage_3__4387_, data_stage_3__4386_, data_stage_3__4385_, data_stage_3__4384_, data_stage_3__4383_, data_stage_3__4382_, data_stage_3__4381_, data_stage_3__4380_, data_stage_3__4379_, data_stage_3__4378_, data_stage_3__4377_, data_stage_3__4376_, data_stage_3__4375_, data_stage_3__4374_, data_stage_3__4373_, data_stage_3__4372_, data_stage_3__4371_, data_stage_3__4370_, data_stage_3__4369_, data_stage_3__4368_, data_stage_3__4367_, data_stage_3__4366_, data_stage_3__4365_, data_stage_3__4364_, data_stage_3__4363_, data_stage_3__4362_, data_stage_3__4361_, data_stage_3__4360_, data_stage_3__4359_, data_stage_3__4358_, data_stage_3__4357_, data_stage_3__4356_, data_stage_3__4355_, data_stage_3__4354_, data_stage_3__4353_, data_stage_3__4352_, data_stage_3__4351_, data_stage_3__4350_, data_stage_3__4349_, data_stage_3__4348_, data_stage_3__4347_, data_stage_3__4346_, data_stage_3__4345_, data_stage_3__4344_, data_stage_3__4343_, data_stage_3__4342_, data_stage_3__4341_, data_stage_3__4340_, data_stage_3__4339_, data_stage_3__4338_, data_stage_3__4337_, data_stage_3__4336_, data_stage_3__4335_, data_stage_3__4334_, data_stage_3__4333_, data_stage_3__4332_, data_stage_3__4331_, data_stage_3__4330_, data_stage_3__4329_, data_stage_3__4328_, data_stage_3__4327_, data_stage_3__4326_, data_stage_3__4325_, data_stage_3__4324_, data_stage_3__4323_, data_stage_3__4322_, data_stage_3__4321_, data_stage_3__4320_, data_stage_3__4319_, data_stage_3__4318_, data_stage_3__4317_, data_stage_3__4316_, data_stage_3__4315_, data_stage_3__4314_, data_stage_3__4313_, data_stage_3__4312_, data_stage_3__4311_, data_stage_3__4310_, data_stage_3__4309_, data_stage_3__4308_, data_stage_3__4307_, data_stage_3__4306_, data_stage_3__4305_, data_stage_3__4304_, data_stage_3__4303_, data_stage_3__4302_, data_stage_3__4301_, data_stage_3__4300_, data_stage_3__4299_, data_stage_3__4298_, data_stage_3__4297_, data_stage_3__4296_, data_stage_3__4295_, data_stage_3__4294_, data_stage_3__4293_, data_stage_3__4292_, data_stage_3__4291_, data_stage_3__4290_, data_stage_3__4289_, data_stage_3__4288_, data_stage_3__4287_, data_stage_3__4286_, data_stage_3__4285_, data_stage_3__4284_, data_stage_3__4283_, data_stage_3__4282_, data_stage_3__4281_, data_stage_3__4280_, data_stage_3__4279_, data_stage_3__4278_, data_stage_3__4277_, data_stage_3__4276_, data_stage_3__4275_, data_stage_3__4274_, data_stage_3__4273_, data_stage_3__4272_, data_stage_3__4271_, data_stage_3__4270_, data_stage_3__4269_, data_stage_3__4268_, data_stage_3__4267_, data_stage_3__4266_, data_stage_3__4265_, data_stage_3__4264_, data_stage_3__4263_, data_stage_3__4262_, data_stage_3__4261_, data_stage_3__4260_, data_stage_3__4259_, data_stage_3__4258_, data_stage_3__4257_, data_stage_3__4256_, data_stage_3__4255_, data_stage_3__4254_, data_stage_3__4253_, data_stage_3__4252_, data_stage_3__4251_, data_stage_3__4250_, data_stage_3__4249_, data_stage_3__4248_, data_stage_3__4247_, data_stage_3__4246_, data_stage_3__4245_, data_stage_3__4244_, data_stage_3__4243_, data_stage_3__4242_, data_stage_3__4241_, data_stage_3__4240_, data_stage_3__4239_, data_stage_3__4238_, data_stage_3__4237_, data_stage_3__4236_, data_stage_3__4235_, data_stage_3__4234_, data_stage_3__4233_, data_stage_3__4232_, data_stage_3__4231_, data_stage_3__4230_, data_stage_3__4229_, data_stage_3__4228_, data_stage_3__4227_, data_stage_3__4226_, data_stage_3__4225_, data_stage_3__4224_, data_stage_3__4223_, data_stage_3__4222_, data_stage_3__4221_, data_stage_3__4220_, data_stage_3__4219_, data_stage_3__4218_, data_stage_3__4217_, data_stage_3__4216_, data_stage_3__4215_, data_stage_3__4214_, data_stage_3__4213_, data_stage_3__4212_, data_stage_3__4211_, data_stage_3__4210_, data_stage_3__4209_, data_stage_3__4208_, data_stage_3__4207_, data_stage_3__4206_, data_stage_3__4205_, data_stage_3__4204_, data_stage_3__4203_, data_stage_3__4202_, data_stage_3__4201_, data_stage_3__4200_, data_stage_3__4199_, data_stage_3__4198_, data_stage_3__4197_, data_stage_3__4196_, data_stage_3__4195_, data_stage_3__4194_, data_stage_3__4193_, data_stage_3__4192_, data_stage_3__4191_, data_stage_3__4190_, data_stage_3__4189_, data_stage_3__4188_, data_stage_3__4187_, data_stage_3__4186_, data_stage_3__4185_, data_stage_3__4184_, data_stage_3__4183_, data_stage_3__4182_, data_stage_3__4181_, data_stage_3__4180_, data_stage_3__4179_, data_stage_3__4178_, data_stage_3__4177_, data_stage_3__4176_, data_stage_3__4175_, data_stage_3__4174_, data_stage_3__4173_, data_stage_3__4172_, data_stage_3__4171_, data_stage_3__4170_, data_stage_3__4169_, data_stage_3__4168_, data_stage_3__4167_, data_stage_3__4166_, data_stage_3__4165_, data_stage_3__4164_, data_stage_3__4163_, data_stage_3__4162_, data_stage_3__4161_, data_stage_3__4160_, data_stage_3__4159_, data_stage_3__4158_, data_stage_3__4157_, data_stage_3__4156_, data_stage_3__4155_, data_stage_3__4154_, data_stage_3__4153_, data_stage_3__4152_, data_stage_3__4151_, data_stage_3__4150_, data_stage_3__4149_, data_stage_3__4148_, data_stage_3__4147_, data_stage_3__4146_, data_stage_3__4145_, data_stage_3__4144_, data_stage_3__4143_, data_stage_3__4142_, data_stage_3__4141_, data_stage_3__4140_, data_stage_3__4139_, data_stage_3__4138_, data_stage_3__4137_, data_stage_3__4136_, data_stage_3__4135_, data_stage_3__4134_, data_stage_3__4133_, data_stage_3__4132_, data_stage_3__4131_, data_stage_3__4130_, data_stage_3__4129_, data_stage_3__4128_, data_stage_3__4127_, data_stage_3__4126_, data_stage_3__4125_, data_stage_3__4124_, data_stage_3__4123_, data_stage_3__4122_, data_stage_3__4121_, data_stage_3__4120_, data_stage_3__4119_, data_stage_3__4118_, data_stage_3__4117_, data_stage_3__4116_, data_stage_3__4115_, data_stage_3__4114_, data_stage_3__4113_, data_stage_3__4112_, data_stage_3__4111_, data_stage_3__4110_, data_stage_3__4109_, data_stage_3__4108_, data_stage_3__4107_, data_stage_3__4106_, data_stage_3__4105_, data_stage_3__4104_, data_stage_3__4103_, data_stage_3__4102_, data_stage_3__4101_, data_stage_3__4100_, data_stage_3__4099_, data_stage_3__4098_, data_stage_3__4097_, data_stage_3__4096_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__6143_, data_stage_4__6142_, data_stage_4__6141_, data_stage_4__6140_, data_stage_4__6139_, data_stage_4__6138_, data_stage_4__6137_, data_stage_4__6136_, data_stage_4__6135_, data_stage_4__6134_, data_stage_4__6133_, data_stage_4__6132_, data_stage_4__6131_, data_stage_4__6130_, data_stage_4__6129_, data_stage_4__6128_, data_stage_4__6127_, data_stage_4__6126_, data_stage_4__6125_, data_stage_4__6124_, data_stage_4__6123_, data_stage_4__6122_, data_stage_4__6121_, data_stage_4__6120_, data_stage_4__6119_, data_stage_4__6118_, data_stage_4__6117_, data_stage_4__6116_, data_stage_4__6115_, data_stage_4__6114_, data_stage_4__6113_, data_stage_4__6112_, data_stage_4__6111_, data_stage_4__6110_, data_stage_4__6109_, data_stage_4__6108_, data_stage_4__6107_, data_stage_4__6106_, data_stage_4__6105_, data_stage_4__6104_, data_stage_4__6103_, data_stage_4__6102_, data_stage_4__6101_, data_stage_4__6100_, data_stage_4__6099_, data_stage_4__6098_, data_stage_4__6097_, data_stage_4__6096_, data_stage_4__6095_, data_stage_4__6094_, data_stage_4__6093_, data_stage_4__6092_, data_stage_4__6091_, data_stage_4__6090_, data_stage_4__6089_, data_stage_4__6088_, data_stage_4__6087_, data_stage_4__6086_, data_stage_4__6085_, data_stage_4__6084_, data_stage_4__6083_, data_stage_4__6082_, data_stage_4__6081_, data_stage_4__6080_, data_stage_4__6079_, data_stage_4__6078_, data_stage_4__6077_, data_stage_4__6076_, data_stage_4__6075_, data_stage_4__6074_, data_stage_4__6073_, data_stage_4__6072_, data_stage_4__6071_, data_stage_4__6070_, data_stage_4__6069_, data_stage_4__6068_, data_stage_4__6067_, data_stage_4__6066_, data_stage_4__6065_, data_stage_4__6064_, data_stage_4__6063_, data_stage_4__6062_, data_stage_4__6061_, data_stage_4__6060_, data_stage_4__6059_, data_stage_4__6058_, data_stage_4__6057_, data_stage_4__6056_, data_stage_4__6055_, data_stage_4__6054_, data_stage_4__6053_, data_stage_4__6052_, data_stage_4__6051_, data_stage_4__6050_, data_stage_4__6049_, data_stage_4__6048_, data_stage_4__6047_, data_stage_4__6046_, data_stage_4__6045_, data_stage_4__6044_, data_stage_4__6043_, data_stage_4__6042_, data_stage_4__6041_, data_stage_4__6040_, data_stage_4__6039_, data_stage_4__6038_, data_stage_4__6037_, data_stage_4__6036_, data_stage_4__6035_, data_stage_4__6034_, data_stage_4__6033_, data_stage_4__6032_, data_stage_4__6031_, data_stage_4__6030_, data_stage_4__6029_, data_stage_4__6028_, data_stage_4__6027_, data_stage_4__6026_, data_stage_4__6025_, data_stage_4__6024_, data_stage_4__6023_, data_stage_4__6022_, data_stage_4__6021_, data_stage_4__6020_, data_stage_4__6019_, data_stage_4__6018_, data_stage_4__6017_, data_stage_4__6016_, data_stage_4__6015_, data_stage_4__6014_, data_stage_4__6013_, data_stage_4__6012_, data_stage_4__6011_, data_stage_4__6010_, data_stage_4__6009_, data_stage_4__6008_, data_stage_4__6007_, data_stage_4__6006_, data_stage_4__6005_, data_stage_4__6004_, data_stage_4__6003_, data_stage_4__6002_, data_stage_4__6001_, data_stage_4__6000_, data_stage_4__5999_, data_stage_4__5998_, data_stage_4__5997_, data_stage_4__5996_, data_stage_4__5995_, data_stage_4__5994_, data_stage_4__5993_, data_stage_4__5992_, data_stage_4__5991_, data_stage_4__5990_, data_stage_4__5989_, data_stage_4__5988_, data_stage_4__5987_, data_stage_4__5986_, data_stage_4__5985_, data_stage_4__5984_, data_stage_4__5983_, data_stage_4__5982_, data_stage_4__5981_, data_stage_4__5980_, data_stage_4__5979_, data_stage_4__5978_, data_stage_4__5977_, data_stage_4__5976_, data_stage_4__5975_, data_stage_4__5974_, data_stage_4__5973_, data_stage_4__5972_, data_stage_4__5971_, data_stage_4__5970_, data_stage_4__5969_, data_stage_4__5968_, data_stage_4__5967_, data_stage_4__5966_, data_stage_4__5965_, data_stage_4__5964_, data_stage_4__5963_, data_stage_4__5962_, data_stage_4__5961_, data_stage_4__5960_, data_stage_4__5959_, data_stage_4__5958_, data_stage_4__5957_, data_stage_4__5956_, data_stage_4__5955_, data_stage_4__5954_, data_stage_4__5953_, data_stage_4__5952_, data_stage_4__5951_, data_stage_4__5950_, data_stage_4__5949_, data_stage_4__5948_, data_stage_4__5947_, data_stage_4__5946_, data_stage_4__5945_, data_stage_4__5944_, data_stage_4__5943_, data_stage_4__5942_, data_stage_4__5941_, data_stage_4__5940_, data_stage_4__5939_, data_stage_4__5938_, data_stage_4__5937_, data_stage_4__5936_, data_stage_4__5935_, data_stage_4__5934_, data_stage_4__5933_, data_stage_4__5932_, data_stage_4__5931_, data_stage_4__5930_, data_stage_4__5929_, data_stage_4__5928_, data_stage_4__5927_, data_stage_4__5926_, data_stage_4__5925_, data_stage_4__5924_, data_stage_4__5923_, data_stage_4__5922_, data_stage_4__5921_, data_stage_4__5920_, data_stage_4__5919_, data_stage_4__5918_, data_stage_4__5917_, data_stage_4__5916_, data_stage_4__5915_, data_stage_4__5914_, data_stage_4__5913_, data_stage_4__5912_, data_stage_4__5911_, data_stage_4__5910_, data_stage_4__5909_, data_stage_4__5908_, data_stage_4__5907_, data_stage_4__5906_, data_stage_4__5905_, data_stage_4__5904_, data_stage_4__5903_, data_stage_4__5902_, data_stage_4__5901_, data_stage_4__5900_, data_stage_4__5899_, data_stage_4__5898_, data_stage_4__5897_, data_stage_4__5896_, data_stage_4__5895_, data_stage_4__5894_, data_stage_4__5893_, data_stage_4__5892_, data_stage_4__5891_, data_stage_4__5890_, data_stage_4__5889_, data_stage_4__5888_, data_stage_4__5887_, data_stage_4__5886_, data_stage_4__5885_, data_stage_4__5884_, data_stage_4__5883_, data_stage_4__5882_, data_stage_4__5881_, data_stage_4__5880_, data_stage_4__5879_, data_stage_4__5878_, data_stage_4__5877_, data_stage_4__5876_, data_stage_4__5875_, data_stage_4__5874_, data_stage_4__5873_, data_stage_4__5872_, data_stage_4__5871_, data_stage_4__5870_, data_stage_4__5869_, data_stage_4__5868_, data_stage_4__5867_, data_stage_4__5866_, data_stage_4__5865_, data_stage_4__5864_, data_stage_4__5863_, data_stage_4__5862_, data_stage_4__5861_, data_stage_4__5860_, data_stage_4__5859_, data_stage_4__5858_, data_stage_4__5857_, data_stage_4__5856_, data_stage_4__5855_, data_stage_4__5854_, data_stage_4__5853_, data_stage_4__5852_, data_stage_4__5851_, data_stage_4__5850_, data_stage_4__5849_, data_stage_4__5848_, data_stage_4__5847_, data_stage_4__5846_, data_stage_4__5845_, data_stage_4__5844_, data_stage_4__5843_, data_stage_4__5842_, data_stage_4__5841_, data_stage_4__5840_, data_stage_4__5839_, data_stage_4__5838_, data_stage_4__5837_, data_stage_4__5836_, data_stage_4__5835_, data_stage_4__5834_, data_stage_4__5833_, data_stage_4__5832_, data_stage_4__5831_, data_stage_4__5830_, data_stage_4__5829_, data_stage_4__5828_, data_stage_4__5827_, data_stage_4__5826_, data_stage_4__5825_, data_stage_4__5824_, data_stage_4__5823_, data_stage_4__5822_, data_stage_4__5821_, data_stage_4__5820_, data_stage_4__5819_, data_stage_4__5818_, data_stage_4__5817_, data_stage_4__5816_, data_stage_4__5815_, data_stage_4__5814_, data_stage_4__5813_, data_stage_4__5812_, data_stage_4__5811_, data_stage_4__5810_, data_stage_4__5809_, data_stage_4__5808_, data_stage_4__5807_, data_stage_4__5806_, data_stage_4__5805_, data_stage_4__5804_, data_stage_4__5803_, data_stage_4__5802_, data_stage_4__5801_, data_stage_4__5800_, data_stage_4__5799_, data_stage_4__5798_, data_stage_4__5797_, data_stage_4__5796_, data_stage_4__5795_, data_stage_4__5794_, data_stage_4__5793_, data_stage_4__5792_, data_stage_4__5791_, data_stage_4__5790_, data_stage_4__5789_, data_stage_4__5788_, data_stage_4__5787_, data_stage_4__5786_, data_stage_4__5785_, data_stage_4__5784_, data_stage_4__5783_, data_stage_4__5782_, data_stage_4__5781_, data_stage_4__5780_, data_stage_4__5779_, data_stage_4__5778_, data_stage_4__5777_, data_stage_4__5776_, data_stage_4__5775_, data_stage_4__5774_, data_stage_4__5773_, data_stage_4__5772_, data_stage_4__5771_, data_stage_4__5770_, data_stage_4__5769_, data_stage_4__5768_, data_stage_4__5767_, data_stage_4__5766_, data_stage_4__5765_, data_stage_4__5764_, data_stage_4__5763_, data_stage_4__5762_, data_stage_4__5761_, data_stage_4__5760_, data_stage_4__5759_, data_stage_4__5758_, data_stage_4__5757_, data_stage_4__5756_, data_stage_4__5755_, data_stage_4__5754_, data_stage_4__5753_, data_stage_4__5752_, data_stage_4__5751_, data_stage_4__5750_, data_stage_4__5749_, data_stage_4__5748_, data_stage_4__5747_, data_stage_4__5746_, data_stage_4__5745_, data_stage_4__5744_, data_stage_4__5743_, data_stage_4__5742_, data_stage_4__5741_, data_stage_4__5740_, data_stage_4__5739_, data_stage_4__5738_, data_stage_4__5737_, data_stage_4__5736_, data_stage_4__5735_, data_stage_4__5734_, data_stage_4__5733_, data_stage_4__5732_, data_stage_4__5731_, data_stage_4__5730_, data_stage_4__5729_, data_stage_4__5728_, data_stage_4__5727_, data_stage_4__5726_, data_stage_4__5725_, data_stage_4__5724_, data_stage_4__5723_, data_stage_4__5722_, data_stage_4__5721_, data_stage_4__5720_, data_stage_4__5719_, data_stage_4__5718_, data_stage_4__5717_, data_stage_4__5716_, data_stage_4__5715_, data_stage_4__5714_, data_stage_4__5713_, data_stage_4__5712_, data_stage_4__5711_, data_stage_4__5710_, data_stage_4__5709_, data_stage_4__5708_, data_stage_4__5707_, data_stage_4__5706_, data_stage_4__5705_, data_stage_4__5704_, data_stage_4__5703_, data_stage_4__5702_, data_stage_4__5701_, data_stage_4__5700_, data_stage_4__5699_, data_stage_4__5698_, data_stage_4__5697_, data_stage_4__5696_, data_stage_4__5695_, data_stage_4__5694_, data_stage_4__5693_, data_stage_4__5692_, data_stage_4__5691_, data_stage_4__5690_, data_stage_4__5689_, data_stage_4__5688_, data_stage_4__5687_, data_stage_4__5686_, data_stage_4__5685_, data_stage_4__5684_, data_stage_4__5683_, data_stage_4__5682_, data_stage_4__5681_, data_stage_4__5680_, data_stage_4__5679_, data_stage_4__5678_, data_stage_4__5677_, data_stage_4__5676_, data_stage_4__5675_, data_stage_4__5674_, data_stage_4__5673_, data_stage_4__5672_, data_stage_4__5671_, data_stage_4__5670_, data_stage_4__5669_, data_stage_4__5668_, data_stage_4__5667_, data_stage_4__5666_, data_stage_4__5665_, data_stage_4__5664_, data_stage_4__5663_, data_stage_4__5662_, data_stage_4__5661_, data_stage_4__5660_, data_stage_4__5659_, data_stage_4__5658_, data_stage_4__5657_, data_stage_4__5656_, data_stage_4__5655_, data_stage_4__5654_, data_stage_4__5653_, data_stage_4__5652_, data_stage_4__5651_, data_stage_4__5650_, data_stage_4__5649_, data_stage_4__5648_, data_stage_4__5647_, data_stage_4__5646_, data_stage_4__5645_, data_stage_4__5644_, data_stage_4__5643_, data_stage_4__5642_, data_stage_4__5641_, data_stage_4__5640_, data_stage_4__5639_, data_stage_4__5638_, data_stage_4__5637_, data_stage_4__5636_, data_stage_4__5635_, data_stage_4__5634_, data_stage_4__5633_, data_stage_4__5632_, data_stage_4__5631_, data_stage_4__5630_, data_stage_4__5629_, data_stage_4__5628_, data_stage_4__5627_, data_stage_4__5626_, data_stage_4__5625_, data_stage_4__5624_, data_stage_4__5623_, data_stage_4__5622_, data_stage_4__5621_, data_stage_4__5620_, data_stage_4__5619_, data_stage_4__5618_, data_stage_4__5617_, data_stage_4__5616_, data_stage_4__5615_, data_stage_4__5614_, data_stage_4__5613_, data_stage_4__5612_, data_stage_4__5611_, data_stage_4__5610_, data_stage_4__5609_, data_stage_4__5608_, data_stage_4__5607_, data_stage_4__5606_, data_stage_4__5605_, data_stage_4__5604_, data_stage_4__5603_, data_stage_4__5602_, data_stage_4__5601_, data_stage_4__5600_, data_stage_4__5599_, data_stage_4__5598_, data_stage_4__5597_, data_stage_4__5596_, data_stage_4__5595_, data_stage_4__5594_, data_stage_4__5593_, data_stage_4__5592_, data_stage_4__5591_, data_stage_4__5590_, data_stage_4__5589_, data_stage_4__5588_, data_stage_4__5587_, data_stage_4__5586_, data_stage_4__5585_, data_stage_4__5584_, data_stage_4__5583_, data_stage_4__5582_, data_stage_4__5581_, data_stage_4__5580_, data_stage_4__5579_, data_stage_4__5578_, data_stage_4__5577_, data_stage_4__5576_, data_stage_4__5575_, data_stage_4__5574_, data_stage_4__5573_, data_stage_4__5572_, data_stage_4__5571_, data_stage_4__5570_, data_stage_4__5569_, data_stage_4__5568_, data_stage_4__5567_, data_stage_4__5566_, data_stage_4__5565_, data_stage_4__5564_, data_stage_4__5563_, data_stage_4__5562_, data_stage_4__5561_, data_stage_4__5560_, data_stage_4__5559_, data_stage_4__5558_, data_stage_4__5557_, data_stage_4__5556_, data_stage_4__5555_, data_stage_4__5554_, data_stage_4__5553_, data_stage_4__5552_, data_stage_4__5551_, data_stage_4__5550_, data_stage_4__5549_, data_stage_4__5548_, data_stage_4__5547_, data_stage_4__5546_, data_stage_4__5545_, data_stage_4__5544_, data_stage_4__5543_, data_stage_4__5542_, data_stage_4__5541_, data_stage_4__5540_, data_stage_4__5539_, data_stage_4__5538_, data_stage_4__5537_, data_stage_4__5536_, data_stage_4__5535_, data_stage_4__5534_, data_stage_4__5533_, data_stage_4__5532_, data_stage_4__5531_, data_stage_4__5530_, data_stage_4__5529_, data_stage_4__5528_, data_stage_4__5527_, data_stage_4__5526_, data_stage_4__5525_, data_stage_4__5524_, data_stage_4__5523_, data_stage_4__5522_, data_stage_4__5521_, data_stage_4__5520_, data_stage_4__5519_, data_stage_4__5518_, data_stage_4__5517_, data_stage_4__5516_, data_stage_4__5515_, data_stage_4__5514_, data_stage_4__5513_, data_stage_4__5512_, data_stage_4__5511_, data_stage_4__5510_, data_stage_4__5509_, data_stage_4__5508_, data_stage_4__5507_, data_stage_4__5506_, data_stage_4__5505_, data_stage_4__5504_, data_stage_4__5503_, data_stage_4__5502_, data_stage_4__5501_, data_stage_4__5500_, data_stage_4__5499_, data_stage_4__5498_, data_stage_4__5497_, data_stage_4__5496_, data_stage_4__5495_, data_stage_4__5494_, data_stage_4__5493_, data_stage_4__5492_, data_stage_4__5491_, data_stage_4__5490_, data_stage_4__5489_, data_stage_4__5488_, data_stage_4__5487_, data_stage_4__5486_, data_stage_4__5485_, data_stage_4__5484_, data_stage_4__5483_, data_stage_4__5482_, data_stage_4__5481_, data_stage_4__5480_, data_stage_4__5479_, data_stage_4__5478_, data_stage_4__5477_, data_stage_4__5476_, data_stage_4__5475_, data_stage_4__5474_, data_stage_4__5473_, data_stage_4__5472_, data_stage_4__5471_, data_stage_4__5470_, data_stage_4__5469_, data_stage_4__5468_, data_stage_4__5467_, data_stage_4__5466_, data_stage_4__5465_, data_stage_4__5464_, data_stage_4__5463_, data_stage_4__5462_, data_stage_4__5461_, data_stage_4__5460_, data_stage_4__5459_, data_stage_4__5458_, data_stage_4__5457_, data_stage_4__5456_, data_stage_4__5455_, data_stage_4__5454_, data_stage_4__5453_, data_stage_4__5452_, data_stage_4__5451_, data_stage_4__5450_, data_stage_4__5449_, data_stage_4__5448_, data_stage_4__5447_, data_stage_4__5446_, data_stage_4__5445_, data_stage_4__5444_, data_stage_4__5443_, data_stage_4__5442_, data_stage_4__5441_, data_stage_4__5440_, data_stage_4__5439_, data_stage_4__5438_, data_stage_4__5437_, data_stage_4__5436_, data_stage_4__5435_, data_stage_4__5434_, data_stage_4__5433_, data_stage_4__5432_, data_stage_4__5431_, data_stage_4__5430_, data_stage_4__5429_, data_stage_4__5428_, data_stage_4__5427_, data_stage_4__5426_, data_stage_4__5425_, data_stage_4__5424_, data_stage_4__5423_, data_stage_4__5422_, data_stage_4__5421_, data_stage_4__5420_, data_stage_4__5419_, data_stage_4__5418_, data_stage_4__5417_, data_stage_4__5416_, data_stage_4__5415_, data_stage_4__5414_, data_stage_4__5413_, data_stage_4__5412_, data_stage_4__5411_, data_stage_4__5410_, data_stage_4__5409_, data_stage_4__5408_, data_stage_4__5407_, data_stage_4__5406_, data_stage_4__5405_, data_stage_4__5404_, data_stage_4__5403_, data_stage_4__5402_, data_stage_4__5401_, data_stage_4__5400_, data_stage_4__5399_, data_stage_4__5398_, data_stage_4__5397_, data_stage_4__5396_, data_stage_4__5395_, data_stage_4__5394_, data_stage_4__5393_, data_stage_4__5392_, data_stage_4__5391_, data_stage_4__5390_, data_stage_4__5389_, data_stage_4__5388_, data_stage_4__5387_, data_stage_4__5386_, data_stage_4__5385_, data_stage_4__5384_, data_stage_4__5383_, data_stage_4__5382_, data_stage_4__5381_, data_stage_4__5380_, data_stage_4__5379_, data_stage_4__5378_, data_stage_4__5377_, data_stage_4__5376_, data_stage_4__5375_, data_stage_4__5374_, data_stage_4__5373_, data_stage_4__5372_, data_stage_4__5371_, data_stage_4__5370_, data_stage_4__5369_, data_stage_4__5368_, data_stage_4__5367_, data_stage_4__5366_, data_stage_4__5365_, data_stage_4__5364_, data_stage_4__5363_, data_stage_4__5362_, data_stage_4__5361_, data_stage_4__5360_, data_stage_4__5359_, data_stage_4__5358_, data_stage_4__5357_, data_stage_4__5356_, data_stage_4__5355_, data_stage_4__5354_, data_stage_4__5353_, data_stage_4__5352_, data_stage_4__5351_, data_stage_4__5350_, data_stage_4__5349_, data_stage_4__5348_, data_stage_4__5347_, data_stage_4__5346_, data_stage_4__5345_, data_stage_4__5344_, data_stage_4__5343_, data_stage_4__5342_, data_stage_4__5341_, data_stage_4__5340_, data_stage_4__5339_, data_stage_4__5338_, data_stage_4__5337_, data_stage_4__5336_, data_stage_4__5335_, data_stage_4__5334_, data_stage_4__5333_, data_stage_4__5332_, data_stage_4__5331_, data_stage_4__5330_, data_stage_4__5329_, data_stage_4__5328_, data_stage_4__5327_, data_stage_4__5326_, data_stage_4__5325_, data_stage_4__5324_, data_stage_4__5323_, data_stage_4__5322_, data_stage_4__5321_, data_stage_4__5320_, data_stage_4__5319_, data_stage_4__5318_, data_stage_4__5317_, data_stage_4__5316_, data_stage_4__5315_, data_stage_4__5314_, data_stage_4__5313_, data_stage_4__5312_, data_stage_4__5311_, data_stage_4__5310_, data_stage_4__5309_, data_stage_4__5308_, data_stage_4__5307_, data_stage_4__5306_, data_stage_4__5305_, data_stage_4__5304_, data_stage_4__5303_, data_stage_4__5302_, data_stage_4__5301_, data_stage_4__5300_, data_stage_4__5299_, data_stage_4__5298_, data_stage_4__5297_, data_stage_4__5296_, data_stage_4__5295_, data_stage_4__5294_, data_stage_4__5293_, data_stage_4__5292_, data_stage_4__5291_, data_stage_4__5290_, data_stage_4__5289_, data_stage_4__5288_, data_stage_4__5287_, data_stage_4__5286_, data_stage_4__5285_, data_stage_4__5284_, data_stage_4__5283_, data_stage_4__5282_, data_stage_4__5281_, data_stage_4__5280_, data_stage_4__5279_, data_stage_4__5278_, data_stage_4__5277_, data_stage_4__5276_, data_stage_4__5275_, data_stage_4__5274_, data_stage_4__5273_, data_stage_4__5272_, data_stage_4__5271_, data_stage_4__5270_, data_stage_4__5269_, data_stage_4__5268_, data_stage_4__5267_, data_stage_4__5266_, data_stage_4__5265_, data_stage_4__5264_, data_stage_4__5263_, data_stage_4__5262_, data_stage_4__5261_, data_stage_4__5260_, data_stage_4__5259_, data_stage_4__5258_, data_stage_4__5257_, data_stage_4__5256_, data_stage_4__5255_, data_stage_4__5254_, data_stage_4__5253_, data_stage_4__5252_, data_stage_4__5251_, data_stage_4__5250_, data_stage_4__5249_, data_stage_4__5248_, data_stage_4__5247_, data_stage_4__5246_, data_stage_4__5245_, data_stage_4__5244_, data_stage_4__5243_, data_stage_4__5242_, data_stage_4__5241_, data_stage_4__5240_, data_stage_4__5239_, data_stage_4__5238_, data_stage_4__5237_, data_stage_4__5236_, data_stage_4__5235_, data_stage_4__5234_, data_stage_4__5233_, data_stage_4__5232_, data_stage_4__5231_, data_stage_4__5230_, data_stage_4__5229_, data_stage_4__5228_, data_stage_4__5227_, data_stage_4__5226_, data_stage_4__5225_, data_stage_4__5224_, data_stage_4__5223_, data_stage_4__5222_, data_stage_4__5221_, data_stage_4__5220_, data_stage_4__5219_, data_stage_4__5218_, data_stage_4__5217_, data_stage_4__5216_, data_stage_4__5215_, data_stage_4__5214_, data_stage_4__5213_, data_stage_4__5212_, data_stage_4__5211_, data_stage_4__5210_, data_stage_4__5209_, data_stage_4__5208_, data_stage_4__5207_, data_stage_4__5206_, data_stage_4__5205_, data_stage_4__5204_, data_stage_4__5203_, data_stage_4__5202_, data_stage_4__5201_, data_stage_4__5200_, data_stage_4__5199_, data_stage_4__5198_, data_stage_4__5197_, data_stage_4__5196_, data_stage_4__5195_, data_stage_4__5194_, data_stage_4__5193_, data_stage_4__5192_, data_stage_4__5191_, data_stage_4__5190_, data_stage_4__5189_, data_stage_4__5188_, data_stage_4__5187_, data_stage_4__5186_, data_stage_4__5185_, data_stage_4__5184_, data_stage_4__5183_, data_stage_4__5182_, data_stage_4__5181_, data_stage_4__5180_, data_stage_4__5179_, data_stage_4__5178_, data_stage_4__5177_, data_stage_4__5176_, data_stage_4__5175_, data_stage_4__5174_, data_stage_4__5173_, data_stage_4__5172_, data_stage_4__5171_, data_stage_4__5170_, data_stage_4__5169_, data_stage_4__5168_, data_stage_4__5167_, data_stage_4__5166_, data_stage_4__5165_, data_stage_4__5164_, data_stage_4__5163_, data_stage_4__5162_, data_stage_4__5161_, data_stage_4__5160_, data_stage_4__5159_, data_stage_4__5158_, data_stage_4__5157_, data_stage_4__5156_, data_stage_4__5155_, data_stage_4__5154_, data_stage_4__5153_, data_stage_4__5152_, data_stage_4__5151_, data_stage_4__5150_, data_stage_4__5149_, data_stage_4__5148_, data_stage_4__5147_, data_stage_4__5146_, data_stage_4__5145_, data_stage_4__5144_, data_stage_4__5143_, data_stage_4__5142_, data_stage_4__5141_, data_stage_4__5140_, data_stage_4__5139_, data_stage_4__5138_, data_stage_4__5137_, data_stage_4__5136_, data_stage_4__5135_, data_stage_4__5134_, data_stage_4__5133_, data_stage_4__5132_, data_stage_4__5131_, data_stage_4__5130_, data_stage_4__5129_, data_stage_4__5128_, data_stage_4__5127_, data_stage_4__5126_, data_stage_4__5125_, data_stage_4__5124_, data_stage_4__5123_, data_stage_4__5122_, data_stage_4__5121_, data_stage_4__5120_, data_stage_4__5119_, data_stage_4__5118_, data_stage_4__5117_, data_stage_4__5116_, data_stage_4__5115_, data_stage_4__5114_, data_stage_4__5113_, data_stage_4__5112_, data_stage_4__5111_, data_stage_4__5110_, data_stage_4__5109_, data_stage_4__5108_, data_stage_4__5107_, data_stage_4__5106_, data_stage_4__5105_, data_stage_4__5104_, data_stage_4__5103_, data_stage_4__5102_, data_stage_4__5101_, data_stage_4__5100_, data_stage_4__5099_, data_stage_4__5098_, data_stage_4__5097_, data_stage_4__5096_, data_stage_4__5095_, data_stage_4__5094_, data_stage_4__5093_, data_stage_4__5092_, data_stage_4__5091_, data_stage_4__5090_, data_stage_4__5089_, data_stage_4__5088_, data_stage_4__5087_, data_stage_4__5086_, data_stage_4__5085_, data_stage_4__5084_, data_stage_4__5083_, data_stage_4__5082_, data_stage_4__5081_, data_stage_4__5080_, data_stage_4__5079_, data_stage_4__5078_, data_stage_4__5077_, data_stage_4__5076_, data_stage_4__5075_, data_stage_4__5074_, data_stage_4__5073_, data_stage_4__5072_, data_stage_4__5071_, data_stage_4__5070_, data_stage_4__5069_, data_stage_4__5068_, data_stage_4__5067_, data_stage_4__5066_, data_stage_4__5065_, data_stage_4__5064_, data_stage_4__5063_, data_stage_4__5062_, data_stage_4__5061_, data_stage_4__5060_, data_stage_4__5059_, data_stage_4__5058_, data_stage_4__5057_, data_stage_4__5056_, data_stage_4__5055_, data_stage_4__5054_, data_stage_4__5053_, data_stage_4__5052_, data_stage_4__5051_, data_stage_4__5050_, data_stage_4__5049_, data_stage_4__5048_, data_stage_4__5047_, data_stage_4__5046_, data_stage_4__5045_, data_stage_4__5044_, data_stage_4__5043_, data_stage_4__5042_, data_stage_4__5041_, data_stage_4__5040_, data_stage_4__5039_, data_stage_4__5038_, data_stage_4__5037_, data_stage_4__5036_, data_stage_4__5035_, data_stage_4__5034_, data_stage_4__5033_, data_stage_4__5032_, data_stage_4__5031_, data_stage_4__5030_, data_stage_4__5029_, data_stage_4__5028_, data_stage_4__5027_, data_stage_4__5026_, data_stage_4__5025_, data_stage_4__5024_, data_stage_4__5023_, data_stage_4__5022_, data_stage_4__5021_, data_stage_4__5020_, data_stage_4__5019_, data_stage_4__5018_, data_stage_4__5017_, data_stage_4__5016_, data_stage_4__5015_, data_stage_4__5014_, data_stage_4__5013_, data_stage_4__5012_, data_stage_4__5011_, data_stage_4__5010_, data_stage_4__5009_, data_stage_4__5008_, data_stage_4__5007_, data_stage_4__5006_, data_stage_4__5005_, data_stage_4__5004_, data_stage_4__5003_, data_stage_4__5002_, data_stage_4__5001_, data_stage_4__5000_, data_stage_4__4999_, data_stage_4__4998_, data_stage_4__4997_, data_stage_4__4996_, data_stage_4__4995_, data_stage_4__4994_, data_stage_4__4993_, data_stage_4__4992_, data_stage_4__4991_, data_stage_4__4990_, data_stage_4__4989_, data_stage_4__4988_, data_stage_4__4987_, data_stage_4__4986_, data_stage_4__4985_, data_stage_4__4984_, data_stage_4__4983_, data_stage_4__4982_, data_stage_4__4981_, data_stage_4__4980_, data_stage_4__4979_, data_stage_4__4978_, data_stage_4__4977_, data_stage_4__4976_, data_stage_4__4975_, data_stage_4__4974_, data_stage_4__4973_, data_stage_4__4972_, data_stage_4__4971_, data_stage_4__4970_, data_stage_4__4969_, data_stage_4__4968_, data_stage_4__4967_, data_stage_4__4966_, data_stage_4__4965_, data_stage_4__4964_, data_stage_4__4963_, data_stage_4__4962_, data_stage_4__4961_, data_stage_4__4960_, data_stage_4__4959_, data_stage_4__4958_, data_stage_4__4957_, data_stage_4__4956_, data_stage_4__4955_, data_stage_4__4954_, data_stage_4__4953_, data_stage_4__4952_, data_stage_4__4951_, data_stage_4__4950_, data_stage_4__4949_, data_stage_4__4948_, data_stage_4__4947_, data_stage_4__4946_, data_stage_4__4945_, data_stage_4__4944_, data_stage_4__4943_, data_stage_4__4942_, data_stage_4__4941_, data_stage_4__4940_, data_stage_4__4939_, data_stage_4__4938_, data_stage_4__4937_, data_stage_4__4936_, data_stage_4__4935_, data_stage_4__4934_, data_stage_4__4933_, data_stage_4__4932_, data_stage_4__4931_, data_stage_4__4930_, data_stage_4__4929_, data_stage_4__4928_, data_stage_4__4927_, data_stage_4__4926_, data_stage_4__4925_, data_stage_4__4924_, data_stage_4__4923_, data_stage_4__4922_, data_stage_4__4921_, data_stage_4__4920_, data_stage_4__4919_, data_stage_4__4918_, data_stage_4__4917_, data_stage_4__4916_, data_stage_4__4915_, data_stage_4__4914_, data_stage_4__4913_, data_stage_4__4912_, data_stage_4__4911_, data_stage_4__4910_, data_stage_4__4909_, data_stage_4__4908_, data_stage_4__4907_, data_stage_4__4906_, data_stage_4__4905_, data_stage_4__4904_, data_stage_4__4903_, data_stage_4__4902_, data_stage_4__4901_, data_stage_4__4900_, data_stage_4__4899_, data_stage_4__4898_, data_stage_4__4897_, data_stage_4__4896_, data_stage_4__4895_, data_stage_4__4894_, data_stage_4__4893_, data_stage_4__4892_, data_stage_4__4891_, data_stage_4__4890_, data_stage_4__4889_, data_stage_4__4888_, data_stage_4__4887_, data_stage_4__4886_, data_stage_4__4885_, data_stage_4__4884_, data_stage_4__4883_, data_stage_4__4882_, data_stage_4__4881_, data_stage_4__4880_, data_stage_4__4879_, data_stage_4__4878_, data_stage_4__4877_, data_stage_4__4876_, data_stage_4__4875_, data_stage_4__4874_, data_stage_4__4873_, data_stage_4__4872_, data_stage_4__4871_, data_stage_4__4870_, data_stage_4__4869_, data_stage_4__4868_, data_stage_4__4867_, data_stage_4__4866_, data_stage_4__4865_, data_stage_4__4864_, data_stage_4__4863_, data_stage_4__4862_, data_stage_4__4861_, data_stage_4__4860_, data_stage_4__4859_, data_stage_4__4858_, data_stage_4__4857_, data_stage_4__4856_, data_stage_4__4855_, data_stage_4__4854_, data_stage_4__4853_, data_stage_4__4852_, data_stage_4__4851_, data_stage_4__4850_, data_stage_4__4849_, data_stage_4__4848_, data_stage_4__4847_, data_stage_4__4846_, data_stage_4__4845_, data_stage_4__4844_, data_stage_4__4843_, data_stage_4__4842_, data_stage_4__4841_, data_stage_4__4840_, data_stage_4__4839_, data_stage_4__4838_, data_stage_4__4837_, data_stage_4__4836_, data_stage_4__4835_, data_stage_4__4834_, data_stage_4__4833_, data_stage_4__4832_, data_stage_4__4831_, data_stage_4__4830_, data_stage_4__4829_, data_stage_4__4828_, data_stage_4__4827_, data_stage_4__4826_, data_stage_4__4825_, data_stage_4__4824_, data_stage_4__4823_, data_stage_4__4822_, data_stage_4__4821_, data_stage_4__4820_, data_stage_4__4819_, data_stage_4__4818_, data_stage_4__4817_, data_stage_4__4816_, data_stage_4__4815_, data_stage_4__4814_, data_stage_4__4813_, data_stage_4__4812_, data_stage_4__4811_, data_stage_4__4810_, data_stage_4__4809_, data_stage_4__4808_, data_stage_4__4807_, data_stage_4__4806_, data_stage_4__4805_, data_stage_4__4804_, data_stage_4__4803_, data_stage_4__4802_, data_stage_4__4801_, data_stage_4__4800_, data_stage_4__4799_, data_stage_4__4798_, data_stage_4__4797_, data_stage_4__4796_, data_stage_4__4795_, data_stage_4__4794_, data_stage_4__4793_, data_stage_4__4792_, data_stage_4__4791_, data_stage_4__4790_, data_stage_4__4789_, data_stage_4__4788_, data_stage_4__4787_, data_stage_4__4786_, data_stage_4__4785_, data_stage_4__4784_, data_stage_4__4783_, data_stage_4__4782_, data_stage_4__4781_, data_stage_4__4780_, data_stage_4__4779_, data_stage_4__4778_, data_stage_4__4777_, data_stage_4__4776_, data_stage_4__4775_, data_stage_4__4774_, data_stage_4__4773_, data_stage_4__4772_, data_stage_4__4771_, data_stage_4__4770_, data_stage_4__4769_, data_stage_4__4768_, data_stage_4__4767_, data_stage_4__4766_, data_stage_4__4765_, data_stage_4__4764_, data_stage_4__4763_, data_stage_4__4762_, data_stage_4__4761_, data_stage_4__4760_, data_stage_4__4759_, data_stage_4__4758_, data_stage_4__4757_, data_stage_4__4756_, data_stage_4__4755_, data_stage_4__4754_, data_stage_4__4753_, data_stage_4__4752_, data_stage_4__4751_, data_stage_4__4750_, data_stage_4__4749_, data_stage_4__4748_, data_stage_4__4747_, data_stage_4__4746_, data_stage_4__4745_, data_stage_4__4744_, data_stage_4__4743_, data_stage_4__4742_, data_stage_4__4741_, data_stage_4__4740_, data_stage_4__4739_, data_stage_4__4738_, data_stage_4__4737_, data_stage_4__4736_, data_stage_4__4735_, data_stage_4__4734_, data_stage_4__4733_, data_stage_4__4732_, data_stage_4__4731_, data_stage_4__4730_, data_stage_4__4729_, data_stage_4__4728_, data_stage_4__4727_, data_stage_4__4726_, data_stage_4__4725_, data_stage_4__4724_, data_stage_4__4723_, data_stage_4__4722_, data_stage_4__4721_, data_stage_4__4720_, data_stage_4__4719_, data_stage_4__4718_, data_stage_4__4717_, data_stage_4__4716_, data_stage_4__4715_, data_stage_4__4714_, data_stage_4__4713_, data_stage_4__4712_, data_stage_4__4711_, data_stage_4__4710_, data_stage_4__4709_, data_stage_4__4708_, data_stage_4__4707_, data_stage_4__4706_, data_stage_4__4705_, data_stage_4__4704_, data_stage_4__4703_, data_stage_4__4702_, data_stage_4__4701_, data_stage_4__4700_, data_stage_4__4699_, data_stage_4__4698_, data_stage_4__4697_, data_stage_4__4696_, data_stage_4__4695_, data_stage_4__4694_, data_stage_4__4693_, data_stage_4__4692_, data_stage_4__4691_, data_stage_4__4690_, data_stage_4__4689_, data_stage_4__4688_, data_stage_4__4687_, data_stage_4__4686_, data_stage_4__4685_, data_stage_4__4684_, data_stage_4__4683_, data_stage_4__4682_, data_stage_4__4681_, data_stage_4__4680_, data_stage_4__4679_, data_stage_4__4678_, data_stage_4__4677_, data_stage_4__4676_, data_stage_4__4675_, data_stage_4__4674_, data_stage_4__4673_, data_stage_4__4672_, data_stage_4__4671_, data_stage_4__4670_, data_stage_4__4669_, data_stage_4__4668_, data_stage_4__4667_, data_stage_4__4666_, data_stage_4__4665_, data_stage_4__4664_, data_stage_4__4663_, data_stage_4__4662_, data_stage_4__4661_, data_stage_4__4660_, data_stage_4__4659_, data_stage_4__4658_, data_stage_4__4657_, data_stage_4__4656_, data_stage_4__4655_, data_stage_4__4654_, data_stage_4__4653_, data_stage_4__4652_, data_stage_4__4651_, data_stage_4__4650_, data_stage_4__4649_, data_stage_4__4648_, data_stage_4__4647_, data_stage_4__4646_, data_stage_4__4645_, data_stage_4__4644_, data_stage_4__4643_, data_stage_4__4642_, data_stage_4__4641_, data_stage_4__4640_, data_stage_4__4639_, data_stage_4__4638_, data_stage_4__4637_, data_stage_4__4636_, data_stage_4__4635_, data_stage_4__4634_, data_stage_4__4633_, data_stage_4__4632_, data_stage_4__4631_, data_stage_4__4630_, data_stage_4__4629_, data_stage_4__4628_, data_stage_4__4627_, data_stage_4__4626_, data_stage_4__4625_, data_stage_4__4624_, data_stage_4__4623_, data_stage_4__4622_, data_stage_4__4621_, data_stage_4__4620_, data_stage_4__4619_, data_stage_4__4618_, data_stage_4__4617_, data_stage_4__4616_, data_stage_4__4615_, data_stage_4__4614_, data_stage_4__4613_, data_stage_4__4612_, data_stage_4__4611_, data_stage_4__4610_, data_stage_4__4609_, data_stage_4__4608_, data_stage_4__4607_, data_stage_4__4606_, data_stage_4__4605_, data_stage_4__4604_, data_stage_4__4603_, data_stage_4__4602_, data_stage_4__4601_, data_stage_4__4600_, data_stage_4__4599_, data_stage_4__4598_, data_stage_4__4597_, data_stage_4__4596_, data_stage_4__4595_, data_stage_4__4594_, data_stage_4__4593_, data_stage_4__4592_, data_stage_4__4591_, data_stage_4__4590_, data_stage_4__4589_, data_stage_4__4588_, data_stage_4__4587_, data_stage_4__4586_, data_stage_4__4585_, data_stage_4__4584_, data_stage_4__4583_, data_stage_4__4582_, data_stage_4__4581_, data_stage_4__4580_, data_stage_4__4579_, data_stage_4__4578_, data_stage_4__4577_, data_stage_4__4576_, data_stage_4__4575_, data_stage_4__4574_, data_stage_4__4573_, data_stage_4__4572_, data_stage_4__4571_, data_stage_4__4570_, data_stage_4__4569_, data_stage_4__4568_, data_stage_4__4567_, data_stage_4__4566_, data_stage_4__4565_, data_stage_4__4564_, data_stage_4__4563_, data_stage_4__4562_, data_stage_4__4561_, data_stage_4__4560_, data_stage_4__4559_, data_stage_4__4558_, data_stage_4__4557_, data_stage_4__4556_, data_stage_4__4555_, data_stage_4__4554_, data_stage_4__4553_, data_stage_4__4552_, data_stage_4__4551_, data_stage_4__4550_, data_stage_4__4549_, data_stage_4__4548_, data_stage_4__4547_, data_stage_4__4546_, data_stage_4__4545_, data_stage_4__4544_, data_stage_4__4543_, data_stage_4__4542_, data_stage_4__4541_, data_stage_4__4540_, data_stage_4__4539_, data_stage_4__4538_, data_stage_4__4537_, data_stage_4__4536_, data_stage_4__4535_, data_stage_4__4534_, data_stage_4__4533_, data_stage_4__4532_, data_stage_4__4531_, data_stage_4__4530_, data_stage_4__4529_, data_stage_4__4528_, data_stage_4__4527_, data_stage_4__4526_, data_stage_4__4525_, data_stage_4__4524_, data_stage_4__4523_, data_stage_4__4522_, data_stage_4__4521_, data_stage_4__4520_, data_stage_4__4519_, data_stage_4__4518_, data_stage_4__4517_, data_stage_4__4516_, data_stage_4__4515_, data_stage_4__4514_, data_stage_4__4513_, data_stage_4__4512_, data_stage_4__4511_, data_stage_4__4510_, data_stage_4__4509_, data_stage_4__4508_, data_stage_4__4507_, data_stage_4__4506_, data_stage_4__4505_, data_stage_4__4504_, data_stage_4__4503_, data_stage_4__4502_, data_stage_4__4501_, data_stage_4__4500_, data_stage_4__4499_, data_stage_4__4498_, data_stage_4__4497_, data_stage_4__4496_, data_stage_4__4495_, data_stage_4__4494_, data_stage_4__4493_, data_stage_4__4492_, data_stage_4__4491_, data_stage_4__4490_, data_stage_4__4489_, data_stage_4__4488_, data_stage_4__4487_, data_stage_4__4486_, data_stage_4__4485_, data_stage_4__4484_, data_stage_4__4483_, data_stage_4__4482_, data_stage_4__4481_, data_stage_4__4480_, data_stage_4__4479_, data_stage_4__4478_, data_stage_4__4477_, data_stage_4__4476_, data_stage_4__4475_, data_stage_4__4474_, data_stage_4__4473_, data_stage_4__4472_, data_stage_4__4471_, data_stage_4__4470_, data_stage_4__4469_, data_stage_4__4468_, data_stage_4__4467_, data_stage_4__4466_, data_stage_4__4465_, data_stage_4__4464_, data_stage_4__4463_, data_stage_4__4462_, data_stage_4__4461_, data_stage_4__4460_, data_stage_4__4459_, data_stage_4__4458_, data_stage_4__4457_, data_stage_4__4456_, data_stage_4__4455_, data_stage_4__4454_, data_stage_4__4453_, data_stage_4__4452_, data_stage_4__4451_, data_stage_4__4450_, data_stage_4__4449_, data_stage_4__4448_, data_stage_4__4447_, data_stage_4__4446_, data_stage_4__4445_, data_stage_4__4444_, data_stage_4__4443_, data_stage_4__4442_, data_stage_4__4441_, data_stage_4__4440_, data_stage_4__4439_, data_stage_4__4438_, data_stage_4__4437_, data_stage_4__4436_, data_stage_4__4435_, data_stage_4__4434_, data_stage_4__4433_, data_stage_4__4432_, data_stage_4__4431_, data_stage_4__4430_, data_stage_4__4429_, data_stage_4__4428_, data_stage_4__4427_, data_stage_4__4426_, data_stage_4__4425_, data_stage_4__4424_, data_stage_4__4423_, data_stage_4__4422_, data_stage_4__4421_, data_stage_4__4420_, data_stage_4__4419_, data_stage_4__4418_, data_stage_4__4417_, data_stage_4__4416_, data_stage_4__4415_, data_stage_4__4414_, data_stage_4__4413_, data_stage_4__4412_, data_stage_4__4411_, data_stage_4__4410_, data_stage_4__4409_, data_stage_4__4408_, data_stage_4__4407_, data_stage_4__4406_, data_stage_4__4405_, data_stage_4__4404_, data_stage_4__4403_, data_stage_4__4402_, data_stage_4__4401_, data_stage_4__4400_, data_stage_4__4399_, data_stage_4__4398_, data_stage_4__4397_, data_stage_4__4396_, data_stage_4__4395_, data_stage_4__4394_, data_stage_4__4393_, data_stage_4__4392_, data_stage_4__4391_, data_stage_4__4390_, data_stage_4__4389_, data_stage_4__4388_, data_stage_4__4387_, data_stage_4__4386_, data_stage_4__4385_, data_stage_4__4384_, data_stage_4__4383_, data_stage_4__4382_, data_stage_4__4381_, data_stage_4__4380_, data_stage_4__4379_, data_stage_4__4378_, data_stage_4__4377_, data_stage_4__4376_, data_stage_4__4375_, data_stage_4__4374_, data_stage_4__4373_, data_stage_4__4372_, data_stage_4__4371_, data_stage_4__4370_, data_stage_4__4369_, data_stage_4__4368_, data_stage_4__4367_, data_stage_4__4366_, data_stage_4__4365_, data_stage_4__4364_, data_stage_4__4363_, data_stage_4__4362_, data_stage_4__4361_, data_stage_4__4360_, data_stage_4__4359_, data_stage_4__4358_, data_stage_4__4357_, data_stage_4__4356_, data_stage_4__4355_, data_stage_4__4354_, data_stage_4__4353_, data_stage_4__4352_, data_stage_4__4351_, data_stage_4__4350_, data_stage_4__4349_, data_stage_4__4348_, data_stage_4__4347_, data_stage_4__4346_, data_stage_4__4345_, data_stage_4__4344_, data_stage_4__4343_, data_stage_4__4342_, data_stage_4__4341_, data_stage_4__4340_, data_stage_4__4339_, data_stage_4__4338_, data_stage_4__4337_, data_stage_4__4336_, data_stage_4__4335_, data_stage_4__4334_, data_stage_4__4333_, data_stage_4__4332_, data_stage_4__4331_, data_stage_4__4330_, data_stage_4__4329_, data_stage_4__4328_, data_stage_4__4327_, data_stage_4__4326_, data_stage_4__4325_, data_stage_4__4324_, data_stage_4__4323_, data_stage_4__4322_, data_stage_4__4321_, data_stage_4__4320_, data_stage_4__4319_, data_stage_4__4318_, data_stage_4__4317_, data_stage_4__4316_, data_stage_4__4315_, data_stage_4__4314_, data_stage_4__4313_, data_stage_4__4312_, data_stage_4__4311_, data_stage_4__4310_, data_stage_4__4309_, data_stage_4__4308_, data_stage_4__4307_, data_stage_4__4306_, data_stage_4__4305_, data_stage_4__4304_, data_stage_4__4303_, data_stage_4__4302_, data_stage_4__4301_, data_stage_4__4300_, data_stage_4__4299_, data_stage_4__4298_, data_stage_4__4297_, data_stage_4__4296_, data_stage_4__4295_, data_stage_4__4294_, data_stage_4__4293_, data_stage_4__4292_, data_stage_4__4291_, data_stage_4__4290_, data_stage_4__4289_, data_stage_4__4288_, data_stage_4__4287_, data_stage_4__4286_, data_stage_4__4285_, data_stage_4__4284_, data_stage_4__4283_, data_stage_4__4282_, data_stage_4__4281_, data_stage_4__4280_, data_stage_4__4279_, data_stage_4__4278_, data_stage_4__4277_, data_stage_4__4276_, data_stage_4__4275_, data_stage_4__4274_, data_stage_4__4273_, data_stage_4__4272_, data_stage_4__4271_, data_stage_4__4270_, data_stage_4__4269_, data_stage_4__4268_, data_stage_4__4267_, data_stage_4__4266_, data_stage_4__4265_, data_stage_4__4264_, data_stage_4__4263_, data_stage_4__4262_, data_stage_4__4261_, data_stage_4__4260_, data_stage_4__4259_, data_stage_4__4258_, data_stage_4__4257_, data_stage_4__4256_, data_stage_4__4255_, data_stage_4__4254_, data_stage_4__4253_, data_stage_4__4252_, data_stage_4__4251_, data_stage_4__4250_, data_stage_4__4249_, data_stage_4__4248_, data_stage_4__4247_, data_stage_4__4246_, data_stage_4__4245_, data_stage_4__4244_, data_stage_4__4243_, data_stage_4__4242_, data_stage_4__4241_, data_stage_4__4240_, data_stage_4__4239_, data_stage_4__4238_, data_stage_4__4237_, data_stage_4__4236_, data_stage_4__4235_, data_stage_4__4234_, data_stage_4__4233_, data_stage_4__4232_, data_stage_4__4231_, data_stage_4__4230_, data_stage_4__4229_, data_stage_4__4228_, data_stage_4__4227_, data_stage_4__4226_, data_stage_4__4225_, data_stage_4__4224_, data_stage_4__4223_, data_stage_4__4222_, data_stage_4__4221_, data_stage_4__4220_, data_stage_4__4219_, data_stage_4__4218_, data_stage_4__4217_, data_stage_4__4216_, data_stage_4__4215_, data_stage_4__4214_, data_stage_4__4213_, data_stage_4__4212_, data_stage_4__4211_, data_stage_4__4210_, data_stage_4__4209_, data_stage_4__4208_, data_stage_4__4207_, data_stage_4__4206_, data_stage_4__4205_, data_stage_4__4204_, data_stage_4__4203_, data_stage_4__4202_, data_stage_4__4201_, data_stage_4__4200_, data_stage_4__4199_, data_stage_4__4198_, data_stage_4__4197_, data_stage_4__4196_, data_stage_4__4195_, data_stage_4__4194_, data_stage_4__4193_, data_stage_4__4192_, data_stage_4__4191_, data_stage_4__4190_, data_stage_4__4189_, data_stage_4__4188_, data_stage_4__4187_, data_stage_4__4186_, data_stage_4__4185_, data_stage_4__4184_, data_stage_4__4183_, data_stage_4__4182_, data_stage_4__4181_, data_stage_4__4180_, data_stage_4__4179_, data_stage_4__4178_, data_stage_4__4177_, data_stage_4__4176_, data_stage_4__4175_, data_stage_4__4174_, data_stage_4__4173_, data_stage_4__4172_, data_stage_4__4171_, data_stage_4__4170_, data_stage_4__4169_, data_stage_4__4168_, data_stage_4__4167_, data_stage_4__4166_, data_stage_4__4165_, data_stage_4__4164_, data_stage_4__4163_, data_stage_4__4162_, data_stage_4__4161_, data_stage_4__4160_, data_stage_4__4159_, data_stage_4__4158_, data_stage_4__4157_, data_stage_4__4156_, data_stage_4__4155_, data_stage_4__4154_, data_stage_4__4153_, data_stage_4__4152_, data_stage_4__4151_, data_stage_4__4150_, data_stage_4__4149_, data_stage_4__4148_, data_stage_4__4147_, data_stage_4__4146_, data_stage_4__4145_, data_stage_4__4144_, data_stage_4__4143_, data_stage_4__4142_, data_stage_4__4141_, data_stage_4__4140_, data_stage_4__4139_, data_stage_4__4138_, data_stage_4__4137_, data_stage_4__4136_, data_stage_4__4135_, data_stage_4__4134_, data_stage_4__4133_, data_stage_4__4132_, data_stage_4__4131_, data_stage_4__4130_, data_stage_4__4129_, data_stage_4__4128_, data_stage_4__4127_, data_stage_4__4126_, data_stage_4__4125_, data_stage_4__4124_, data_stage_4__4123_, data_stage_4__4122_, data_stage_4__4121_, data_stage_4__4120_, data_stage_4__4119_, data_stage_4__4118_, data_stage_4__4117_, data_stage_4__4116_, data_stage_4__4115_, data_stage_4__4114_, data_stage_4__4113_, data_stage_4__4112_, data_stage_4__4111_, data_stage_4__4110_, data_stage_4__4109_, data_stage_4__4108_, data_stage_4__4107_, data_stage_4__4106_, data_stage_4__4105_, data_stage_4__4104_, data_stage_4__4103_, data_stage_4__4102_, data_stage_4__4101_, data_stage_4__4100_, data_stage_4__4099_, data_stage_4__4098_, data_stage_4__4097_, data_stage_4__4096_ })
  );


  bsg_swap_width_p1024
  mux_stage_3__mux_swap_3__swap_inst
  (
    .data_i({ data_stage_3__8191_, data_stage_3__8190_, data_stage_3__8189_, data_stage_3__8188_, data_stage_3__8187_, data_stage_3__8186_, data_stage_3__8185_, data_stage_3__8184_, data_stage_3__8183_, data_stage_3__8182_, data_stage_3__8181_, data_stage_3__8180_, data_stage_3__8179_, data_stage_3__8178_, data_stage_3__8177_, data_stage_3__8176_, data_stage_3__8175_, data_stage_3__8174_, data_stage_3__8173_, data_stage_3__8172_, data_stage_3__8171_, data_stage_3__8170_, data_stage_3__8169_, data_stage_3__8168_, data_stage_3__8167_, data_stage_3__8166_, data_stage_3__8165_, data_stage_3__8164_, data_stage_3__8163_, data_stage_3__8162_, data_stage_3__8161_, data_stage_3__8160_, data_stage_3__8159_, data_stage_3__8158_, data_stage_3__8157_, data_stage_3__8156_, data_stage_3__8155_, data_stage_3__8154_, data_stage_3__8153_, data_stage_3__8152_, data_stage_3__8151_, data_stage_3__8150_, data_stage_3__8149_, data_stage_3__8148_, data_stage_3__8147_, data_stage_3__8146_, data_stage_3__8145_, data_stage_3__8144_, data_stage_3__8143_, data_stage_3__8142_, data_stage_3__8141_, data_stage_3__8140_, data_stage_3__8139_, data_stage_3__8138_, data_stage_3__8137_, data_stage_3__8136_, data_stage_3__8135_, data_stage_3__8134_, data_stage_3__8133_, data_stage_3__8132_, data_stage_3__8131_, data_stage_3__8130_, data_stage_3__8129_, data_stage_3__8128_, data_stage_3__8127_, data_stage_3__8126_, data_stage_3__8125_, data_stage_3__8124_, data_stage_3__8123_, data_stage_3__8122_, data_stage_3__8121_, data_stage_3__8120_, data_stage_3__8119_, data_stage_3__8118_, data_stage_3__8117_, data_stage_3__8116_, data_stage_3__8115_, data_stage_3__8114_, data_stage_3__8113_, data_stage_3__8112_, data_stage_3__8111_, data_stage_3__8110_, data_stage_3__8109_, data_stage_3__8108_, data_stage_3__8107_, data_stage_3__8106_, data_stage_3__8105_, data_stage_3__8104_, data_stage_3__8103_, data_stage_3__8102_, data_stage_3__8101_, data_stage_3__8100_, data_stage_3__8099_, data_stage_3__8098_, data_stage_3__8097_, data_stage_3__8096_, data_stage_3__8095_, data_stage_3__8094_, data_stage_3__8093_, data_stage_3__8092_, data_stage_3__8091_, data_stage_3__8090_, data_stage_3__8089_, data_stage_3__8088_, data_stage_3__8087_, data_stage_3__8086_, data_stage_3__8085_, data_stage_3__8084_, data_stage_3__8083_, data_stage_3__8082_, data_stage_3__8081_, data_stage_3__8080_, data_stage_3__8079_, data_stage_3__8078_, data_stage_3__8077_, data_stage_3__8076_, data_stage_3__8075_, data_stage_3__8074_, data_stage_3__8073_, data_stage_3__8072_, data_stage_3__8071_, data_stage_3__8070_, data_stage_3__8069_, data_stage_3__8068_, data_stage_3__8067_, data_stage_3__8066_, data_stage_3__8065_, data_stage_3__8064_, data_stage_3__8063_, data_stage_3__8062_, data_stage_3__8061_, data_stage_3__8060_, data_stage_3__8059_, data_stage_3__8058_, data_stage_3__8057_, data_stage_3__8056_, data_stage_3__8055_, data_stage_3__8054_, data_stage_3__8053_, data_stage_3__8052_, data_stage_3__8051_, data_stage_3__8050_, data_stage_3__8049_, data_stage_3__8048_, data_stage_3__8047_, data_stage_3__8046_, data_stage_3__8045_, data_stage_3__8044_, data_stage_3__8043_, data_stage_3__8042_, data_stage_3__8041_, data_stage_3__8040_, data_stage_3__8039_, data_stage_3__8038_, data_stage_3__8037_, data_stage_3__8036_, data_stage_3__8035_, data_stage_3__8034_, data_stage_3__8033_, data_stage_3__8032_, data_stage_3__8031_, data_stage_3__8030_, data_stage_3__8029_, data_stage_3__8028_, data_stage_3__8027_, data_stage_3__8026_, data_stage_3__8025_, data_stage_3__8024_, data_stage_3__8023_, data_stage_3__8022_, data_stage_3__8021_, data_stage_3__8020_, data_stage_3__8019_, data_stage_3__8018_, data_stage_3__8017_, data_stage_3__8016_, data_stage_3__8015_, data_stage_3__8014_, data_stage_3__8013_, data_stage_3__8012_, data_stage_3__8011_, data_stage_3__8010_, data_stage_3__8009_, data_stage_3__8008_, data_stage_3__8007_, data_stage_3__8006_, data_stage_3__8005_, data_stage_3__8004_, data_stage_3__8003_, data_stage_3__8002_, data_stage_3__8001_, data_stage_3__8000_, data_stage_3__7999_, data_stage_3__7998_, data_stage_3__7997_, data_stage_3__7996_, data_stage_3__7995_, data_stage_3__7994_, data_stage_3__7993_, data_stage_3__7992_, data_stage_3__7991_, data_stage_3__7990_, data_stage_3__7989_, data_stage_3__7988_, data_stage_3__7987_, data_stage_3__7986_, data_stage_3__7985_, data_stage_3__7984_, data_stage_3__7983_, data_stage_3__7982_, data_stage_3__7981_, data_stage_3__7980_, data_stage_3__7979_, data_stage_3__7978_, data_stage_3__7977_, data_stage_3__7976_, data_stage_3__7975_, data_stage_3__7974_, data_stage_3__7973_, data_stage_3__7972_, data_stage_3__7971_, data_stage_3__7970_, data_stage_3__7969_, data_stage_3__7968_, data_stage_3__7967_, data_stage_3__7966_, data_stage_3__7965_, data_stage_3__7964_, data_stage_3__7963_, data_stage_3__7962_, data_stage_3__7961_, data_stage_3__7960_, data_stage_3__7959_, data_stage_3__7958_, data_stage_3__7957_, data_stage_3__7956_, data_stage_3__7955_, data_stage_3__7954_, data_stage_3__7953_, data_stage_3__7952_, data_stage_3__7951_, data_stage_3__7950_, data_stage_3__7949_, data_stage_3__7948_, data_stage_3__7947_, data_stage_3__7946_, data_stage_3__7945_, data_stage_3__7944_, data_stage_3__7943_, data_stage_3__7942_, data_stage_3__7941_, data_stage_3__7940_, data_stage_3__7939_, data_stage_3__7938_, data_stage_3__7937_, data_stage_3__7936_, data_stage_3__7935_, data_stage_3__7934_, data_stage_3__7933_, data_stage_3__7932_, data_stage_3__7931_, data_stage_3__7930_, data_stage_3__7929_, data_stage_3__7928_, data_stage_3__7927_, data_stage_3__7926_, data_stage_3__7925_, data_stage_3__7924_, data_stage_3__7923_, data_stage_3__7922_, data_stage_3__7921_, data_stage_3__7920_, data_stage_3__7919_, data_stage_3__7918_, data_stage_3__7917_, data_stage_3__7916_, data_stage_3__7915_, data_stage_3__7914_, data_stage_3__7913_, data_stage_3__7912_, data_stage_3__7911_, data_stage_3__7910_, data_stage_3__7909_, data_stage_3__7908_, data_stage_3__7907_, data_stage_3__7906_, data_stage_3__7905_, data_stage_3__7904_, data_stage_3__7903_, data_stage_3__7902_, data_stage_3__7901_, data_stage_3__7900_, data_stage_3__7899_, data_stage_3__7898_, data_stage_3__7897_, data_stage_3__7896_, data_stage_3__7895_, data_stage_3__7894_, data_stage_3__7893_, data_stage_3__7892_, data_stage_3__7891_, data_stage_3__7890_, data_stage_3__7889_, data_stage_3__7888_, data_stage_3__7887_, data_stage_3__7886_, data_stage_3__7885_, data_stage_3__7884_, data_stage_3__7883_, data_stage_3__7882_, data_stage_3__7881_, data_stage_3__7880_, data_stage_3__7879_, data_stage_3__7878_, data_stage_3__7877_, data_stage_3__7876_, data_stage_3__7875_, data_stage_3__7874_, data_stage_3__7873_, data_stage_3__7872_, data_stage_3__7871_, data_stage_3__7870_, data_stage_3__7869_, data_stage_3__7868_, data_stage_3__7867_, data_stage_3__7866_, data_stage_3__7865_, data_stage_3__7864_, data_stage_3__7863_, data_stage_3__7862_, data_stage_3__7861_, data_stage_3__7860_, data_stage_3__7859_, data_stage_3__7858_, data_stage_3__7857_, data_stage_3__7856_, data_stage_3__7855_, data_stage_3__7854_, data_stage_3__7853_, data_stage_3__7852_, data_stage_3__7851_, data_stage_3__7850_, data_stage_3__7849_, data_stage_3__7848_, data_stage_3__7847_, data_stage_3__7846_, data_stage_3__7845_, data_stage_3__7844_, data_stage_3__7843_, data_stage_3__7842_, data_stage_3__7841_, data_stage_3__7840_, data_stage_3__7839_, data_stage_3__7838_, data_stage_3__7837_, data_stage_3__7836_, data_stage_3__7835_, data_stage_3__7834_, data_stage_3__7833_, data_stage_3__7832_, data_stage_3__7831_, data_stage_3__7830_, data_stage_3__7829_, data_stage_3__7828_, data_stage_3__7827_, data_stage_3__7826_, data_stage_3__7825_, data_stage_3__7824_, data_stage_3__7823_, data_stage_3__7822_, data_stage_3__7821_, data_stage_3__7820_, data_stage_3__7819_, data_stage_3__7818_, data_stage_3__7817_, data_stage_3__7816_, data_stage_3__7815_, data_stage_3__7814_, data_stage_3__7813_, data_stage_3__7812_, data_stage_3__7811_, data_stage_3__7810_, data_stage_3__7809_, data_stage_3__7808_, data_stage_3__7807_, data_stage_3__7806_, data_stage_3__7805_, data_stage_3__7804_, data_stage_3__7803_, data_stage_3__7802_, data_stage_3__7801_, data_stage_3__7800_, data_stage_3__7799_, data_stage_3__7798_, data_stage_3__7797_, data_stage_3__7796_, data_stage_3__7795_, data_stage_3__7794_, data_stage_3__7793_, data_stage_3__7792_, data_stage_3__7791_, data_stage_3__7790_, data_stage_3__7789_, data_stage_3__7788_, data_stage_3__7787_, data_stage_3__7786_, data_stage_3__7785_, data_stage_3__7784_, data_stage_3__7783_, data_stage_3__7782_, data_stage_3__7781_, data_stage_3__7780_, data_stage_3__7779_, data_stage_3__7778_, data_stage_3__7777_, data_stage_3__7776_, data_stage_3__7775_, data_stage_3__7774_, data_stage_3__7773_, data_stage_3__7772_, data_stage_3__7771_, data_stage_3__7770_, data_stage_3__7769_, data_stage_3__7768_, data_stage_3__7767_, data_stage_3__7766_, data_stage_3__7765_, data_stage_3__7764_, data_stage_3__7763_, data_stage_3__7762_, data_stage_3__7761_, data_stage_3__7760_, data_stage_3__7759_, data_stage_3__7758_, data_stage_3__7757_, data_stage_3__7756_, data_stage_3__7755_, data_stage_3__7754_, data_stage_3__7753_, data_stage_3__7752_, data_stage_3__7751_, data_stage_3__7750_, data_stage_3__7749_, data_stage_3__7748_, data_stage_3__7747_, data_stage_3__7746_, data_stage_3__7745_, data_stage_3__7744_, data_stage_3__7743_, data_stage_3__7742_, data_stage_3__7741_, data_stage_3__7740_, data_stage_3__7739_, data_stage_3__7738_, data_stage_3__7737_, data_stage_3__7736_, data_stage_3__7735_, data_stage_3__7734_, data_stage_3__7733_, data_stage_3__7732_, data_stage_3__7731_, data_stage_3__7730_, data_stage_3__7729_, data_stage_3__7728_, data_stage_3__7727_, data_stage_3__7726_, data_stage_3__7725_, data_stage_3__7724_, data_stage_3__7723_, data_stage_3__7722_, data_stage_3__7721_, data_stage_3__7720_, data_stage_3__7719_, data_stage_3__7718_, data_stage_3__7717_, data_stage_3__7716_, data_stage_3__7715_, data_stage_3__7714_, data_stage_3__7713_, data_stage_3__7712_, data_stage_3__7711_, data_stage_3__7710_, data_stage_3__7709_, data_stage_3__7708_, data_stage_3__7707_, data_stage_3__7706_, data_stage_3__7705_, data_stage_3__7704_, data_stage_3__7703_, data_stage_3__7702_, data_stage_3__7701_, data_stage_3__7700_, data_stage_3__7699_, data_stage_3__7698_, data_stage_3__7697_, data_stage_3__7696_, data_stage_3__7695_, data_stage_3__7694_, data_stage_3__7693_, data_stage_3__7692_, data_stage_3__7691_, data_stage_3__7690_, data_stage_3__7689_, data_stage_3__7688_, data_stage_3__7687_, data_stage_3__7686_, data_stage_3__7685_, data_stage_3__7684_, data_stage_3__7683_, data_stage_3__7682_, data_stage_3__7681_, data_stage_3__7680_, data_stage_3__7679_, data_stage_3__7678_, data_stage_3__7677_, data_stage_3__7676_, data_stage_3__7675_, data_stage_3__7674_, data_stage_3__7673_, data_stage_3__7672_, data_stage_3__7671_, data_stage_3__7670_, data_stage_3__7669_, data_stage_3__7668_, data_stage_3__7667_, data_stage_3__7666_, data_stage_3__7665_, data_stage_3__7664_, data_stage_3__7663_, data_stage_3__7662_, data_stage_3__7661_, data_stage_3__7660_, data_stage_3__7659_, data_stage_3__7658_, data_stage_3__7657_, data_stage_3__7656_, data_stage_3__7655_, data_stage_3__7654_, data_stage_3__7653_, data_stage_3__7652_, data_stage_3__7651_, data_stage_3__7650_, data_stage_3__7649_, data_stage_3__7648_, data_stage_3__7647_, data_stage_3__7646_, data_stage_3__7645_, data_stage_3__7644_, data_stage_3__7643_, data_stage_3__7642_, data_stage_3__7641_, data_stage_3__7640_, data_stage_3__7639_, data_stage_3__7638_, data_stage_3__7637_, data_stage_3__7636_, data_stage_3__7635_, data_stage_3__7634_, data_stage_3__7633_, data_stage_3__7632_, data_stage_3__7631_, data_stage_3__7630_, data_stage_3__7629_, data_stage_3__7628_, data_stage_3__7627_, data_stage_3__7626_, data_stage_3__7625_, data_stage_3__7624_, data_stage_3__7623_, data_stage_3__7622_, data_stage_3__7621_, data_stage_3__7620_, data_stage_3__7619_, data_stage_3__7618_, data_stage_3__7617_, data_stage_3__7616_, data_stage_3__7615_, data_stage_3__7614_, data_stage_3__7613_, data_stage_3__7612_, data_stage_3__7611_, data_stage_3__7610_, data_stage_3__7609_, data_stage_3__7608_, data_stage_3__7607_, data_stage_3__7606_, data_stage_3__7605_, data_stage_3__7604_, data_stage_3__7603_, data_stage_3__7602_, data_stage_3__7601_, data_stage_3__7600_, data_stage_3__7599_, data_stage_3__7598_, data_stage_3__7597_, data_stage_3__7596_, data_stage_3__7595_, data_stage_3__7594_, data_stage_3__7593_, data_stage_3__7592_, data_stage_3__7591_, data_stage_3__7590_, data_stage_3__7589_, data_stage_3__7588_, data_stage_3__7587_, data_stage_3__7586_, data_stage_3__7585_, data_stage_3__7584_, data_stage_3__7583_, data_stage_3__7582_, data_stage_3__7581_, data_stage_3__7580_, data_stage_3__7579_, data_stage_3__7578_, data_stage_3__7577_, data_stage_3__7576_, data_stage_3__7575_, data_stage_3__7574_, data_stage_3__7573_, data_stage_3__7572_, data_stage_3__7571_, data_stage_3__7570_, data_stage_3__7569_, data_stage_3__7568_, data_stage_3__7567_, data_stage_3__7566_, data_stage_3__7565_, data_stage_3__7564_, data_stage_3__7563_, data_stage_3__7562_, data_stage_3__7561_, data_stage_3__7560_, data_stage_3__7559_, data_stage_3__7558_, data_stage_3__7557_, data_stage_3__7556_, data_stage_3__7555_, data_stage_3__7554_, data_stage_3__7553_, data_stage_3__7552_, data_stage_3__7551_, data_stage_3__7550_, data_stage_3__7549_, data_stage_3__7548_, data_stage_3__7547_, data_stage_3__7546_, data_stage_3__7545_, data_stage_3__7544_, data_stage_3__7543_, data_stage_3__7542_, data_stage_3__7541_, data_stage_3__7540_, data_stage_3__7539_, data_stage_3__7538_, data_stage_3__7537_, data_stage_3__7536_, data_stage_3__7535_, data_stage_3__7534_, data_stage_3__7533_, data_stage_3__7532_, data_stage_3__7531_, data_stage_3__7530_, data_stage_3__7529_, data_stage_3__7528_, data_stage_3__7527_, data_stage_3__7526_, data_stage_3__7525_, data_stage_3__7524_, data_stage_3__7523_, data_stage_3__7522_, data_stage_3__7521_, data_stage_3__7520_, data_stage_3__7519_, data_stage_3__7518_, data_stage_3__7517_, data_stage_3__7516_, data_stage_3__7515_, data_stage_3__7514_, data_stage_3__7513_, data_stage_3__7512_, data_stage_3__7511_, data_stage_3__7510_, data_stage_3__7509_, data_stage_3__7508_, data_stage_3__7507_, data_stage_3__7506_, data_stage_3__7505_, data_stage_3__7504_, data_stage_3__7503_, data_stage_3__7502_, data_stage_3__7501_, data_stage_3__7500_, data_stage_3__7499_, data_stage_3__7498_, data_stage_3__7497_, data_stage_3__7496_, data_stage_3__7495_, data_stage_3__7494_, data_stage_3__7493_, data_stage_3__7492_, data_stage_3__7491_, data_stage_3__7490_, data_stage_3__7489_, data_stage_3__7488_, data_stage_3__7487_, data_stage_3__7486_, data_stage_3__7485_, data_stage_3__7484_, data_stage_3__7483_, data_stage_3__7482_, data_stage_3__7481_, data_stage_3__7480_, data_stage_3__7479_, data_stage_3__7478_, data_stage_3__7477_, data_stage_3__7476_, data_stage_3__7475_, data_stage_3__7474_, data_stage_3__7473_, data_stage_3__7472_, data_stage_3__7471_, data_stage_3__7470_, data_stage_3__7469_, data_stage_3__7468_, data_stage_3__7467_, data_stage_3__7466_, data_stage_3__7465_, data_stage_3__7464_, data_stage_3__7463_, data_stage_3__7462_, data_stage_3__7461_, data_stage_3__7460_, data_stage_3__7459_, data_stage_3__7458_, data_stage_3__7457_, data_stage_3__7456_, data_stage_3__7455_, data_stage_3__7454_, data_stage_3__7453_, data_stage_3__7452_, data_stage_3__7451_, data_stage_3__7450_, data_stage_3__7449_, data_stage_3__7448_, data_stage_3__7447_, data_stage_3__7446_, data_stage_3__7445_, data_stage_3__7444_, data_stage_3__7443_, data_stage_3__7442_, data_stage_3__7441_, data_stage_3__7440_, data_stage_3__7439_, data_stage_3__7438_, data_stage_3__7437_, data_stage_3__7436_, data_stage_3__7435_, data_stage_3__7434_, data_stage_3__7433_, data_stage_3__7432_, data_stage_3__7431_, data_stage_3__7430_, data_stage_3__7429_, data_stage_3__7428_, data_stage_3__7427_, data_stage_3__7426_, data_stage_3__7425_, data_stage_3__7424_, data_stage_3__7423_, data_stage_3__7422_, data_stage_3__7421_, data_stage_3__7420_, data_stage_3__7419_, data_stage_3__7418_, data_stage_3__7417_, data_stage_3__7416_, data_stage_3__7415_, data_stage_3__7414_, data_stage_3__7413_, data_stage_3__7412_, data_stage_3__7411_, data_stage_3__7410_, data_stage_3__7409_, data_stage_3__7408_, data_stage_3__7407_, data_stage_3__7406_, data_stage_3__7405_, data_stage_3__7404_, data_stage_3__7403_, data_stage_3__7402_, data_stage_3__7401_, data_stage_3__7400_, data_stage_3__7399_, data_stage_3__7398_, data_stage_3__7397_, data_stage_3__7396_, data_stage_3__7395_, data_stage_3__7394_, data_stage_3__7393_, data_stage_3__7392_, data_stage_3__7391_, data_stage_3__7390_, data_stage_3__7389_, data_stage_3__7388_, data_stage_3__7387_, data_stage_3__7386_, data_stage_3__7385_, data_stage_3__7384_, data_stage_3__7383_, data_stage_3__7382_, data_stage_3__7381_, data_stage_3__7380_, data_stage_3__7379_, data_stage_3__7378_, data_stage_3__7377_, data_stage_3__7376_, data_stage_3__7375_, data_stage_3__7374_, data_stage_3__7373_, data_stage_3__7372_, data_stage_3__7371_, data_stage_3__7370_, data_stage_3__7369_, data_stage_3__7368_, data_stage_3__7367_, data_stage_3__7366_, data_stage_3__7365_, data_stage_3__7364_, data_stage_3__7363_, data_stage_3__7362_, data_stage_3__7361_, data_stage_3__7360_, data_stage_3__7359_, data_stage_3__7358_, data_stage_3__7357_, data_stage_3__7356_, data_stage_3__7355_, data_stage_3__7354_, data_stage_3__7353_, data_stage_3__7352_, data_stage_3__7351_, data_stage_3__7350_, data_stage_3__7349_, data_stage_3__7348_, data_stage_3__7347_, data_stage_3__7346_, data_stage_3__7345_, data_stage_3__7344_, data_stage_3__7343_, data_stage_3__7342_, data_stage_3__7341_, data_stage_3__7340_, data_stage_3__7339_, data_stage_3__7338_, data_stage_3__7337_, data_stage_3__7336_, data_stage_3__7335_, data_stage_3__7334_, data_stage_3__7333_, data_stage_3__7332_, data_stage_3__7331_, data_stage_3__7330_, data_stage_3__7329_, data_stage_3__7328_, data_stage_3__7327_, data_stage_3__7326_, data_stage_3__7325_, data_stage_3__7324_, data_stage_3__7323_, data_stage_3__7322_, data_stage_3__7321_, data_stage_3__7320_, data_stage_3__7319_, data_stage_3__7318_, data_stage_3__7317_, data_stage_3__7316_, data_stage_3__7315_, data_stage_3__7314_, data_stage_3__7313_, data_stage_3__7312_, data_stage_3__7311_, data_stage_3__7310_, data_stage_3__7309_, data_stage_3__7308_, data_stage_3__7307_, data_stage_3__7306_, data_stage_3__7305_, data_stage_3__7304_, data_stage_3__7303_, data_stage_3__7302_, data_stage_3__7301_, data_stage_3__7300_, data_stage_3__7299_, data_stage_3__7298_, data_stage_3__7297_, data_stage_3__7296_, data_stage_3__7295_, data_stage_3__7294_, data_stage_3__7293_, data_stage_3__7292_, data_stage_3__7291_, data_stage_3__7290_, data_stage_3__7289_, data_stage_3__7288_, data_stage_3__7287_, data_stage_3__7286_, data_stage_3__7285_, data_stage_3__7284_, data_stage_3__7283_, data_stage_3__7282_, data_stage_3__7281_, data_stage_3__7280_, data_stage_3__7279_, data_stage_3__7278_, data_stage_3__7277_, data_stage_3__7276_, data_stage_3__7275_, data_stage_3__7274_, data_stage_3__7273_, data_stage_3__7272_, data_stage_3__7271_, data_stage_3__7270_, data_stage_3__7269_, data_stage_3__7268_, data_stage_3__7267_, data_stage_3__7266_, data_stage_3__7265_, data_stage_3__7264_, data_stage_3__7263_, data_stage_3__7262_, data_stage_3__7261_, data_stage_3__7260_, data_stage_3__7259_, data_stage_3__7258_, data_stage_3__7257_, data_stage_3__7256_, data_stage_3__7255_, data_stage_3__7254_, data_stage_3__7253_, data_stage_3__7252_, data_stage_3__7251_, data_stage_3__7250_, data_stage_3__7249_, data_stage_3__7248_, data_stage_3__7247_, data_stage_3__7246_, data_stage_3__7245_, data_stage_3__7244_, data_stage_3__7243_, data_stage_3__7242_, data_stage_3__7241_, data_stage_3__7240_, data_stage_3__7239_, data_stage_3__7238_, data_stage_3__7237_, data_stage_3__7236_, data_stage_3__7235_, data_stage_3__7234_, data_stage_3__7233_, data_stage_3__7232_, data_stage_3__7231_, data_stage_3__7230_, data_stage_3__7229_, data_stage_3__7228_, data_stage_3__7227_, data_stage_3__7226_, data_stage_3__7225_, data_stage_3__7224_, data_stage_3__7223_, data_stage_3__7222_, data_stage_3__7221_, data_stage_3__7220_, data_stage_3__7219_, data_stage_3__7218_, data_stage_3__7217_, data_stage_3__7216_, data_stage_3__7215_, data_stage_3__7214_, data_stage_3__7213_, data_stage_3__7212_, data_stage_3__7211_, data_stage_3__7210_, data_stage_3__7209_, data_stage_3__7208_, data_stage_3__7207_, data_stage_3__7206_, data_stage_3__7205_, data_stage_3__7204_, data_stage_3__7203_, data_stage_3__7202_, data_stage_3__7201_, data_stage_3__7200_, data_stage_3__7199_, data_stage_3__7198_, data_stage_3__7197_, data_stage_3__7196_, data_stage_3__7195_, data_stage_3__7194_, data_stage_3__7193_, data_stage_3__7192_, data_stage_3__7191_, data_stage_3__7190_, data_stage_3__7189_, data_stage_3__7188_, data_stage_3__7187_, data_stage_3__7186_, data_stage_3__7185_, data_stage_3__7184_, data_stage_3__7183_, data_stage_3__7182_, data_stage_3__7181_, data_stage_3__7180_, data_stage_3__7179_, data_stage_3__7178_, data_stage_3__7177_, data_stage_3__7176_, data_stage_3__7175_, data_stage_3__7174_, data_stage_3__7173_, data_stage_3__7172_, data_stage_3__7171_, data_stage_3__7170_, data_stage_3__7169_, data_stage_3__7168_, data_stage_3__7167_, data_stage_3__7166_, data_stage_3__7165_, data_stage_3__7164_, data_stage_3__7163_, data_stage_3__7162_, data_stage_3__7161_, data_stage_3__7160_, data_stage_3__7159_, data_stage_3__7158_, data_stage_3__7157_, data_stage_3__7156_, data_stage_3__7155_, data_stage_3__7154_, data_stage_3__7153_, data_stage_3__7152_, data_stage_3__7151_, data_stage_3__7150_, data_stage_3__7149_, data_stage_3__7148_, data_stage_3__7147_, data_stage_3__7146_, data_stage_3__7145_, data_stage_3__7144_, data_stage_3__7143_, data_stage_3__7142_, data_stage_3__7141_, data_stage_3__7140_, data_stage_3__7139_, data_stage_3__7138_, data_stage_3__7137_, data_stage_3__7136_, data_stage_3__7135_, data_stage_3__7134_, data_stage_3__7133_, data_stage_3__7132_, data_stage_3__7131_, data_stage_3__7130_, data_stage_3__7129_, data_stage_3__7128_, data_stage_3__7127_, data_stage_3__7126_, data_stage_3__7125_, data_stage_3__7124_, data_stage_3__7123_, data_stage_3__7122_, data_stage_3__7121_, data_stage_3__7120_, data_stage_3__7119_, data_stage_3__7118_, data_stage_3__7117_, data_stage_3__7116_, data_stage_3__7115_, data_stage_3__7114_, data_stage_3__7113_, data_stage_3__7112_, data_stage_3__7111_, data_stage_3__7110_, data_stage_3__7109_, data_stage_3__7108_, data_stage_3__7107_, data_stage_3__7106_, data_stage_3__7105_, data_stage_3__7104_, data_stage_3__7103_, data_stage_3__7102_, data_stage_3__7101_, data_stage_3__7100_, data_stage_3__7099_, data_stage_3__7098_, data_stage_3__7097_, data_stage_3__7096_, data_stage_3__7095_, data_stage_3__7094_, data_stage_3__7093_, data_stage_3__7092_, data_stage_3__7091_, data_stage_3__7090_, data_stage_3__7089_, data_stage_3__7088_, data_stage_3__7087_, data_stage_3__7086_, data_stage_3__7085_, data_stage_3__7084_, data_stage_3__7083_, data_stage_3__7082_, data_stage_3__7081_, data_stage_3__7080_, data_stage_3__7079_, data_stage_3__7078_, data_stage_3__7077_, data_stage_3__7076_, data_stage_3__7075_, data_stage_3__7074_, data_stage_3__7073_, data_stage_3__7072_, data_stage_3__7071_, data_stage_3__7070_, data_stage_3__7069_, data_stage_3__7068_, data_stage_3__7067_, data_stage_3__7066_, data_stage_3__7065_, data_stage_3__7064_, data_stage_3__7063_, data_stage_3__7062_, data_stage_3__7061_, data_stage_3__7060_, data_stage_3__7059_, data_stage_3__7058_, data_stage_3__7057_, data_stage_3__7056_, data_stage_3__7055_, data_stage_3__7054_, data_stage_3__7053_, data_stage_3__7052_, data_stage_3__7051_, data_stage_3__7050_, data_stage_3__7049_, data_stage_3__7048_, data_stage_3__7047_, data_stage_3__7046_, data_stage_3__7045_, data_stage_3__7044_, data_stage_3__7043_, data_stage_3__7042_, data_stage_3__7041_, data_stage_3__7040_, data_stage_3__7039_, data_stage_3__7038_, data_stage_3__7037_, data_stage_3__7036_, data_stage_3__7035_, data_stage_3__7034_, data_stage_3__7033_, data_stage_3__7032_, data_stage_3__7031_, data_stage_3__7030_, data_stage_3__7029_, data_stage_3__7028_, data_stage_3__7027_, data_stage_3__7026_, data_stage_3__7025_, data_stage_3__7024_, data_stage_3__7023_, data_stage_3__7022_, data_stage_3__7021_, data_stage_3__7020_, data_stage_3__7019_, data_stage_3__7018_, data_stage_3__7017_, data_stage_3__7016_, data_stage_3__7015_, data_stage_3__7014_, data_stage_3__7013_, data_stage_3__7012_, data_stage_3__7011_, data_stage_3__7010_, data_stage_3__7009_, data_stage_3__7008_, data_stage_3__7007_, data_stage_3__7006_, data_stage_3__7005_, data_stage_3__7004_, data_stage_3__7003_, data_stage_3__7002_, data_stage_3__7001_, data_stage_3__7000_, data_stage_3__6999_, data_stage_3__6998_, data_stage_3__6997_, data_stage_3__6996_, data_stage_3__6995_, data_stage_3__6994_, data_stage_3__6993_, data_stage_3__6992_, data_stage_3__6991_, data_stage_3__6990_, data_stage_3__6989_, data_stage_3__6988_, data_stage_3__6987_, data_stage_3__6986_, data_stage_3__6985_, data_stage_3__6984_, data_stage_3__6983_, data_stage_3__6982_, data_stage_3__6981_, data_stage_3__6980_, data_stage_3__6979_, data_stage_3__6978_, data_stage_3__6977_, data_stage_3__6976_, data_stage_3__6975_, data_stage_3__6974_, data_stage_3__6973_, data_stage_3__6972_, data_stage_3__6971_, data_stage_3__6970_, data_stage_3__6969_, data_stage_3__6968_, data_stage_3__6967_, data_stage_3__6966_, data_stage_3__6965_, data_stage_3__6964_, data_stage_3__6963_, data_stage_3__6962_, data_stage_3__6961_, data_stage_3__6960_, data_stage_3__6959_, data_stage_3__6958_, data_stage_3__6957_, data_stage_3__6956_, data_stage_3__6955_, data_stage_3__6954_, data_stage_3__6953_, data_stage_3__6952_, data_stage_3__6951_, data_stage_3__6950_, data_stage_3__6949_, data_stage_3__6948_, data_stage_3__6947_, data_stage_3__6946_, data_stage_3__6945_, data_stage_3__6944_, data_stage_3__6943_, data_stage_3__6942_, data_stage_3__6941_, data_stage_3__6940_, data_stage_3__6939_, data_stage_3__6938_, data_stage_3__6937_, data_stage_3__6936_, data_stage_3__6935_, data_stage_3__6934_, data_stage_3__6933_, data_stage_3__6932_, data_stage_3__6931_, data_stage_3__6930_, data_stage_3__6929_, data_stage_3__6928_, data_stage_3__6927_, data_stage_3__6926_, data_stage_3__6925_, data_stage_3__6924_, data_stage_3__6923_, data_stage_3__6922_, data_stage_3__6921_, data_stage_3__6920_, data_stage_3__6919_, data_stage_3__6918_, data_stage_3__6917_, data_stage_3__6916_, data_stage_3__6915_, data_stage_3__6914_, data_stage_3__6913_, data_stage_3__6912_, data_stage_3__6911_, data_stage_3__6910_, data_stage_3__6909_, data_stage_3__6908_, data_stage_3__6907_, data_stage_3__6906_, data_stage_3__6905_, data_stage_3__6904_, data_stage_3__6903_, data_stage_3__6902_, data_stage_3__6901_, data_stage_3__6900_, data_stage_3__6899_, data_stage_3__6898_, data_stage_3__6897_, data_stage_3__6896_, data_stage_3__6895_, data_stage_3__6894_, data_stage_3__6893_, data_stage_3__6892_, data_stage_3__6891_, data_stage_3__6890_, data_stage_3__6889_, data_stage_3__6888_, data_stage_3__6887_, data_stage_3__6886_, data_stage_3__6885_, data_stage_3__6884_, data_stage_3__6883_, data_stage_3__6882_, data_stage_3__6881_, data_stage_3__6880_, data_stage_3__6879_, data_stage_3__6878_, data_stage_3__6877_, data_stage_3__6876_, data_stage_3__6875_, data_stage_3__6874_, data_stage_3__6873_, data_stage_3__6872_, data_stage_3__6871_, data_stage_3__6870_, data_stage_3__6869_, data_stage_3__6868_, data_stage_3__6867_, data_stage_3__6866_, data_stage_3__6865_, data_stage_3__6864_, data_stage_3__6863_, data_stage_3__6862_, data_stage_3__6861_, data_stage_3__6860_, data_stage_3__6859_, data_stage_3__6858_, data_stage_3__6857_, data_stage_3__6856_, data_stage_3__6855_, data_stage_3__6854_, data_stage_3__6853_, data_stage_3__6852_, data_stage_3__6851_, data_stage_3__6850_, data_stage_3__6849_, data_stage_3__6848_, data_stage_3__6847_, data_stage_3__6846_, data_stage_3__6845_, data_stage_3__6844_, data_stage_3__6843_, data_stage_3__6842_, data_stage_3__6841_, data_stage_3__6840_, data_stage_3__6839_, data_stage_3__6838_, data_stage_3__6837_, data_stage_3__6836_, data_stage_3__6835_, data_stage_3__6834_, data_stage_3__6833_, data_stage_3__6832_, data_stage_3__6831_, data_stage_3__6830_, data_stage_3__6829_, data_stage_3__6828_, data_stage_3__6827_, data_stage_3__6826_, data_stage_3__6825_, data_stage_3__6824_, data_stage_3__6823_, data_stage_3__6822_, data_stage_3__6821_, data_stage_3__6820_, data_stage_3__6819_, data_stage_3__6818_, data_stage_3__6817_, data_stage_3__6816_, data_stage_3__6815_, data_stage_3__6814_, data_stage_3__6813_, data_stage_3__6812_, data_stage_3__6811_, data_stage_3__6810_, data_stage_3__6809_, data_stage_3__6808_, data_stage_3__6807_, data_stage_3__6806_, data_stage_3__6805_, data_stage_3__6804_, data_stage_3__6803_, data_stage_3__6802_, data_stage_3__6801_, data_stage_3__6800_, data_stage_3__6799_, data_stage_3__6798_, data_stage_3__6797_, data_stage_3__6796_, data_stage_3__6795_, data_stage_3__6794_, data_stage_3__6793_, data_stage_3__6792_, data_stage_3__6791_, data_stage_3__6790_, data_stage_3__6789_, data_stage_3__6788_, data_stage_3__6787_, data_stage_3__6786_, data_stage_3__6785_, data_stage_3__6784_, data_stage_3__6783_, data_stage_3__6782_, data_stage_3__6781_, data_stage_3__6780_, data_stage_3__6779_, data_stage_3__6778_, data_stage_3__6777_, data_stage_3__6776_, data_stage_3__6775_, data_stage_3__6774_, data_stage_3__6773_, data_stage_3__6772_, data_stage_3__6771_, data_stage_3__6770_, data_stage_3__6769_, data_stage_3__6768_, data_stage_3__6767_, data_stage_3__6766_, data_stage_3__6765_, data_stage_3__6764_, data_stage_3__6763_, data_stage_3__6762_, data_stage_3__6761_, data_stage_3__6760_, data_stage_3__6759_, data_stage_3__6758_, data_stage_3__6757_, data_stage_3__6756_, data_stage_3__6755_, data_stage_3__6754_, data_stage_3__6753_, data_stage_3__6752_, data_stage_3__6751_, data_stage_3__6750_, data_stage_3__6749_, data_stage_3__6748_, data_stage_3__6747_, data_stage_3__6746_, data_stage_3__6745_, data_stage_3__6744_, data_stage_3__6743_, data_stage_3__6742_, data_stage_3__6741_, data_stage_3__6740_, data_stage_3__6739_, data_stage_3__6738_, data_stage_3__6737_, data_stage_3__6736_, data_stage_3__6735_, data_stage_3__6734_, data_stage_3__6733_, data_stage_3__6732_, data_stage_3__6731_, data_stage_3__6730_, data_stage_3__6729_, data_stage_3__6728_, data_stage_3__6727_, data_stage_3__6726_, data_stage_3__6725_, data_stage_3__6724_, data_stage_3__6723_, data_stage_3__6722_, data_stage_3__6721_, data_stage_3__6720_, data_stage_3__6719_, data_stage_3__6718_, data_stage_3__6717_, data_stage_3__6716_, data_stage_3__6715_, data_stage_3__6714_, data_stage_3__6713_, data_stage_3__6712_, data_stage_3__6711_, data_stage_3__6710_, data_stage_3__6709_, data_stage_3__6708_, data_stage_3__6707_, data_stage_3__6706_, data_stage_3__6705_, data_stage_3__6704_, data_stage_3__6703_, data_stage_3__6702_, data_stage_3__6701_, data_stage_3__6700_, data_stage_3__6699_, data_stage_3__6698_, data_stage_3__6697_, data_stage_3__6696_, data_stage_3__6695_, data_stage_3__6694_, data_stage_3__6693_, data_stage_3__6692_, data_stage_3__6691_, data_stage_3__6690_, data_stage_3__6689_, data_stage_3__6688_, data_stage_3__6687_, data_stage_3__6686_, data_stage_3__6685_, data_stage_3__6684_, data_stage_3__6683_, data_stage_3__6682_, data_stage_3__6681_, data_stage_3__6680_, data_stage_3__6679_, data_stage_3__6678_, data_stage_3__6677_, data_stage_3__6676_, data_stage_3__6675_, data_stage_3__6674_, data_stage_3__6673_, data_stage_3__6672_, data_stage_3__6671_, data_stage_3__6670_, data_stage_3__6669_, data_stage_3__6668_, data_stage_3__6667_, data_stage_3__6666_, data_stage_3__6665_, data_stage_3__6664_, data_stage_3__6663_, data_stage_3__6662_, data_stage_3__6661_, data_stage_3__6660_, data_stage_3__6659_, data_stage_3__6658_, data_stage_3__6657_, data_stage_3__6656_, data_stage_3__6655_, data_stage_3__6654_, data_stage_3__6653_, data_stage_3__6652_, data_stage_3__6651_, data_stage_3__6650_, data_stage_3__6649_, data_stage_3__6648_, data_stage_3__6647_, data_stage_3__6646_, data_stage_3__6645_, data_stage_3__6644_, data_stage_3__6643_, data_stage_3__6642_, data_stage_3__6641_, data_stage_3__6640_, data_stage_3__6639_, data_stage_3__6638_, data_stage_3__6637_, data_stage_3__6636_, data_stage_3__6635_, data_stage_3__6634_, data_stage_3__6633_, data_stage_3__6632_, data_stage_3__6631_, data_stage_3__6630_, data_stage_3__6629_, data_stage_3__6628_, data_stage_3__6627_, data_stage_3__6626_, data_stage_3__6625_, data_stage_3__6624_, data_stage_3__6623_, data_stage_3__6622_, data_stage_3__6621_, data_stage_3__6620_, data_stage_3__6619_, data_stage_3__6618_, data_stage_3__6617_, data_stage_3__6616_, data_stage_3__6615_, data_stage_3__6614_, data_stage_3__6613_, data_stage_3__6612_, data_stage_3__6611_, data_stage_3__6610_, data_stage_3__6609_, data_stage_3__6608_, data_stage_3__6607_, data_stage_3__6606_, data_stage_3__6605_, data_stage_3__6604_, data_stage_3__6603_, data_stage_3__6602_, data_stage_3__6601_, data_stage_3__6600_, data_stage_3__6599_, data_stage_3__6598_, data_stage_3__6597_, data_stage_3__6596_, data_stage_3__6595_, data_stage_3__6594_, data_stage_3__6593_, data_stage_3__6592_, data_stage_3__6591_, data_stage_3__6590_, data_stage_3__6589_, data_stage_3__6588_, data_stage_3__6587_, data_stage_3__6586_, data_stage_3__6585_, data_stage_3__6584_, data_stage_3__6583_, data_stage_3__6582_, data_stage_3__6581_, data_stage_3__6580_, data_stage_3__6579_, data_stage_3__6578_, data_stage_3__6577_, data_stage_3__6576_, data_stage_3__6575_, data_stage_3__6574_, data_stage_3__6573_, data_stage_3__6572_, data_stage_3__6571_, data_stage_3__6570_, data_stage_3__6569_, data_stage_3__6568_, data_stage_3__6567_, data_stage_3__6566_, data_stage_3__6565_, data_stage_3__6564_, data_stage_3__6563_, data_stage_3__6562_, data_stage_3__6561_, data_stage_3__6560_, data_stage_3__6559_, data_stage_3__6558_, data_stage_3__6557_, data_stage_3__6556_, data_stage_3__6555_, data_stage_3__6554_, data_stage_3__6553_, data_stage_3__6552_, data_stage_3__6551_, data_stage_3__6550_, data_stage_3__6549_, data_stage_3__6548_, data_stage_3__6547_, data_stage_3__6546_, data_stage_3__6545_, data_stage_3__6544_, data_stage_3__6543_, data_stage_3__6542_, data_stage_3__6541_, data_stage_3__6540_, data_stage_3__6539_, data_stage_3__6538_, data_stage_3__6537_, data_stage_3__6536_, data_stage_3__6535_, data_stage_3__6534_, data_stage_3__6533_, data_stage_3__6532_, data_stage_3__6531_, data_stage_3__6530_, data_stage_3__6529_, data_stage_3__6528_, data_stage_3__6527_, data_stage_3__6526_, data_stage_3__6525_, data_stage_3__6524_, data_stage_3__6523_, data_stage_3__6522_, data_stage_3__6521_, data_stage_3__6520_, data_stage_3__6519_, data_stage_3__6518_, data_stage_3__6517_, data_stage_3__6516_, data_stage_3__6515_, data_stage_3__6514_, data_stage_3__6513_, data_stage_3__6512_, data_stage_3__6511_, data_stage_3__6510_, data_stage_3__6509_, data_stage_3__6508_, data_stage_3__6507_, data_stage_3__6506_, data_stage_3__6505_, data_stage_3__6504_, data_stage_3__6503_, data_stage_3__6502_, data_stage_3__6501_, data_stage_3__6500_, data_stage_3__6499_, data_stage_3__6498_, data_stage_3__6497_, data_stage_3__6496_, data_stage_3__6495_, data_stage_3__6494_, data_stage_3__6493_, data_stage_3__6492_, data_stage_3__6491_, data_stage_3__6490_, data_stage_3__6489_, data_stage_3__6488_, data_stage_3__6487_, data_stage_3__6486_, data_stage_3__6485_, data_stage_3__6484_, data_stage_3__6483_, data_stage_3__6482_, data_stage_3__6481_, data_stage_3__6480_, data_stage_3__6479_, data_stage_3__6478_, data_stage_3__6477_, data_stage_3__6476_, data_stage_3__6475_, data_stage_3__6474_, data_stage_3__6473_, data_stage_3__6472_, data_stage_3__6471_, data_stage_3__6470_, data_stage_3__6469_, data_stage_3__6468_, data_stage_3__6467_, data_stage_3__6466_, data_stage_3__6465_, data_stage_3__6464_, data_stage_3__6463_, data_stage_3__6462_, data_stage_3__6461_, data_stage_3__6460_, data_stage_3__6459_, data_stage_3__6458_, data_stage_3__6457_, data_stage_3__6456_, data_stage_3__6455_, data_stage_3__6454_, data_stage_3__6453_, data_stage_3__6452_, data_stage_3__6451_, data_stage_3__6450_, data_stage_3__6449_, data_stage_3__6448_, data_stage_3__6447_, data_stage_3__6446_, data_stage_3__6445_, data_stage_3__6444_, data_stage_3__6443_, data_stage_3__6442_, data_stage_3__6441_, data_stage_3__6440_, data_stage_3__6439_, data_stage_3__6438_, data_stage_3__6437_, data_stage_3__6436_, data_stage_3__6435_, data_stage_3__6434_, data_stage_3__6433_, data_stage_3__6432_, data_stage_3__6431_, data_stage_3__6430_, data_stage_3__6429_, data_stage_3__6428_, data_stage_3__6427_, data_stage_3__6426_, data_stage_3__6425_, data_stage_3__6424_, data_stage_3__6423_, data_stage_3__6422_, data_stage_3__6421_, data_stage_3__6420_, data_stage_3__6419_, data_stage_3__6418_, data_stage_3__6417_, data_stage_3__6416_, data_stage_3__6415_, data_stage_3__6414_, data_stage_3__6413_, data_stage_3__6412_, data_stage_3__6411_, data_stage_3__6410_, data_stage_3__6409_, data_stage_3__6408_, data_stage_3__6407_, data_stage_3__6406_, data_stage_3__6405_, data_stage_3__6404_, data_stage_3__6403_, data_stage_3__6402_, data_stage_3__6401_, data_stage_3__6400_, data_stage_3__6399_, data_stage_3__6398_, data_stage_3__6397_, data_stage_3__6396_, data_stage_3__6395_, data_stage_3__6394_, data_stage_3__6393_, data_stage_3__6392_, data_stage_3__6391_, data_stage_3__6390_, data_stage_3__6389_, data_stage_3__6388_, data_stage_3__6387_, data_stage_3__6386_, data_stage_3__6385_, data_stage_3__6384_, data_stage_3__6383_, data_stage_3__6382_, data_stage_3__6381_, data_stage_3__6380_, data_stage_3__6379_, data_stage_3__6378_, data_stage_3__6377_, data_stage_3__6376_, data_stage_3__6375_, data_stage_3__6374_, data_stage_3__6373_, data_stage_3__6372_, data_stage_3__6371_, data_stage_3__6370_, data_stage_3__6369_, data_stage_3__6368_, data_stage_3__6367_, data_stage_3__6366_, data_stage_3__6365_, data_stage_3__6364_, data_stage_3__6363_, data_stage_3__6362_, data_stage_3__6361_, data_stage_3__6360_, data_stage_3__6359_, data_stage_3__6358_, data_stage_3__6357_, data_stage_3__6356_, data_stage_3__6355_, data_stage_3__6354_, data_stage_3__6353_, data_stage_3__6352_, data_stage_3__6351_, data_stage_3__6350_, data_stage_3__6349_, data_stage_3__6348_, data_stage_3__6347_, data_stage_3__6346_, data_stage_3__6345_, data_stage_3__6344_, data_stage_3__6343_, data_stage_3__6342_, data_stage_3__6341_, data_stage_3__6340_, data_stage_3__6339_, data_stage_3__6338_, data_stage_3__6337_, data_stage_3__6336_, data_stage_3__6335_, data_stage_3__6334_, data_stage_3__6333_, data_stage_3__6332_, data_stage_3__6331_, data_stage_3__6330_, data_stage_3__6329_, data_stage_3__6328_, data_stage_3__6327_, data_stage_3__6326_, data_stage_3__6325_, data_stage_3__6324_, data_stage_3__6323_, data_stage_3__6322_, data_stage_3__6321_, data_stage_3__6320_, data_stage_3__6319_, data_stage_3__6318_, data_stage_3__6317_, data_stage_3__6316_, data_stage_3__6315_, data_stage_3__6314_, data_stage_3__6313_, data_stage_3__6312_, data_stage_3__6311_, data_stage_3__6310_, data_stage_3__6309_, data_stage_3__6308_, data_stage_3__6307_, data_stage_3__6306_, data_stage_3__6305_, data_stage_3__6304_, data_stage_3__6303_, data_stage_3__6302_, data_stage_3__6301_, data_stage_3__6300_, data_stage_3__6299_, data_stage_3__6298_, data_stage_3__6297_, data_stage_3__6296_, data_stage_3__6295_, data_stage_3__6294_, data_stage_3__6293_, data_stage_3__6292_, data_stage_3__6291_, data_stage_3__6290_, data_stage_3__6289_, data_stage_3__6288_, data_stage_3__6287_, data_stage_3__6286_, data_stage_3__6285_, data_stage_3__6284_, data_stage_3__6283_, data_stage_3__6282_, data_stage_3__6281_, data_stage_3__6280_, data_stage_3__6279_, data_stage_3__6278_, data_stage_3__6277_, data_stage_3__6276_, data_stage_3__6275_, data_stage_3__6274_, data_stage_3__6273_, data_stage_3__6272_, data_stage_3__6271_, data_stage_3__6270_, data_stage_3__6269_, data_stage_3__6268_, data_stage_3__6267_, data_stage_3__6266_, data_stage_3__6265_, data_stage_3__6264_, data_stage_3__6263_, data_stage_3__6262_, data_stage_3__6261_, data_stage_3__6260_, data_stage_3__6259_, data_stage_3__6258_, data_stage_3__6257_, data_stage_3__6256_, data_stage_3__6255_, data_stage_3__6254_, data_stage_3__6253_, data_stage_3__6252_, data_stage_3__6251_, data_stage_3__6250_, data_stage_3__6249_, data_stage_3__6248_, data_stage_3__6247_, data_stage_3__6246_, data_stage_3__6245_, data_stage_3__6244_, data_stage_3__6243_, data_stage_3__6242_, data_stage_3__6241_, data_stage_3__6240_, data_stage_3__6239_, data_stage_3__6238_, data_stage_3__6237_, data_stage_3__6236_, data_stage_3__6235_, data_stage_3__6234_, data_stage_3__6233_, data_stage_3__6232_, data_stage_3__6231_, data_stage_3__6230_, data_stage_3__6229_, data_stage_3__6228_, data_stage_3__6227_, data_stage_3__6226_, data_stage_3__6225_, data_stage_3__6224_, data_stage_3__6223_, data_stage_3__6222_, data_stage_3__6221_, data_stage_3__6220_, data_stage_3__6219_, data_stage_3__6218_, data_stage_3__6217_, data_stage_3__6216_, data_stage_3__6215_, data_stage_3__6214_, data_stage_3__6213_, data_stage_3__6212_, data_stage_3__6211_, data_stage_3__6210_, data_stage_3__6209_, data_stage_3__6208_, data_stage_3__6207_, data_stage_3__6206_, data_stage_3__6205_, data_stage_3__6204_, data_stage_3__6203_, data_stage_3__6202_, data_stage_3__6201_, data_stage_3__6200_, data_stage_3__6199_, data_stage_3__6198_, data_stage_3__6197_, data_stage_3__6196_, data_stage_3__6195_, data_stage_3__6194_, data_stage_3__6193_, data_stage_3__6192_, data_stage_3__6191_, data_stage_3__6190_, data_stage_3__6189_, data_stage_3__6188_, data_stage_3__6187_, data_stage_3__6186_, data_stage_3__6185_, data_stage_3__6184_, data_stage_3__6183_, data_stage_3__6182_, data_stage_3__6181_, data_stage_3__6180_, data_stage_3__6179_, data_stage_3__6178_, data_stage_3__6177_, data_stage_3__6176_, data_stage_3__6175_, data_stage_3__6174_, data_stage_3__6173_, data_stage_3__6172_, data_stage_3__6171_, data_stage_3__6170_, data_stage_3__6169_, data_stage_3__6168_, data_stage_3__6167_, data_stage_3__6166_, data_stage_3__6165_, data_stage_3__6164_, data_stage_3__6163_, data_stage_3__6162_, data_stage_3__6161_, data_stage_3__6160_, data_stage_3__6159_, data_stage_3__6158_, data_stage_3__6157_, data_stage_3__6156_, data_stage_3__6155_, data_stage_3__6154_, data_stage_3__6153_, data_stage_3__6152_, data_stage_3__6151_, data_stage_3__6150_, data_stage_3__6149_, data_stage_3__6148_, data_stage_3__6147_, data_stage_3__6146_, data_stage_3__6145_, data_stage_3__6144_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__8191_, data_stage_4__8190_, data_stage_4__8189_, data_stage_4__8188_, data_stage_4__8187_, data_stage_4__8186_, data_stage_4__8185_, data_stage_4__8184_, data_stage_4__8183_, data_stage_4__8182_, data_stage_4__8181_, data_stage_4__8180_, data_stage_4__8179_, data_stage_4__8178_, data_stage_4__8177_, data_stage_4__8176_, data_stage_4__8175_, data_stage_4__8174_, data_stage_4__8173_, data_stage_4__8172_, data_stage_4__8171_, data_stage_4__8170_, data_stage_4__8169_, data_stage_4__8168_, data_stage_4__8167_, data_stage_4__8166_, data_stage_4__8165_, data_stage_4__8164_, data_stage_4__8163_, data_stage_4__8162_, data_stage_4__8161_, data_stage_4__8160_, data_stage_4__8159_, data_stage_4__8158_, data_stage_4__8157_, data_stage_4__8156_, data_stage_4__8155_, data_stage_4__8154_, data_stage_4__8153_, data_stage_4__8152_, data_stage_4__8151_, data_stage_4__8150_, data_stage_4__8149_, data_stage_4__8148_, data_stage_4__8147_, data_stage_4__8146_, data_stage_4__8145_, data_stage_4__8144_, data_stage_4__8143_, data_stage_4__8142_, data_stage_4__8141_, data_stage_4__8140_, data_stage_4__8139_, data_stage_4__8138_, data_stage_4__8137_, data_stage_4__8136_, data_stage_4__8135_, data_stage_4__8134_, data_stage_4__8133_, data_stage_4__8132_, data_stage_4__8131_, data_stage_4__8130_, data_stage_4__8129_, data_stage_4__8128_, data_stage_4__8127_, data_stage_4__8126_, data_stage_4__8125_, data_stage_4__8124_, data_stage_4__8123_, data_stage_4__8122_, data_stage_4__8121_, data_stage_4__8120_, data_stage_4__8119_, data_stage_4__8118_, data_stage_4__8117_, data_stage_4__8116_, data_stage_4__8115_, data_stage_4__8114_, data_stage_4__8113_, data_stage_4__8112_, data_stage_4__8111_, data_stage_4__8110_, data_stage_4__8109_, data_stage_4__8108_, data_stage_4__8107_, data_stage_4__8106_, data_stage_4__8105_, data_stage_4__8104_, data_stage_4__8103_, data_stage_4__8102_, data_stage_4__8101_, data_stage_4__8100_, data_stage_4__8099_, data_stage_4__8098_, data_stage_4__8097_, data_stage_4__8096_, data_stage_4__8095_, data_stage_4__8094_, data_stage_4__8093_, data_stage_4__8092_, data_stage_4__8091_, data_stage_4__8090_, data_stage_4__8089_, data_stage_4__8088_, data_stage_4__8087_, data_stage_4__8086_, data_stage_4__8085_, data_stage_4__8084_, data_stage_4__8083_, data_stage_4__8082_, data_stage_4__8081_, data_stage_4__8080_, data_stage_4__8079_, data_stage_4__8078_, data_stage_4__8077_, data_stage_4__8076_, data_stage_4__8075_, data_stage_4__8074_, data_stage_4__8073_, data_stage_4__8072_, data_stage_4__8071_, data_stage_4__8070_, data_stage_4__8069_, data_stage_4__8068_, data_stage_4__8067_, data_stage_4__8066_, data_stage_4__8065_, data_stage_4__8064_, data_stage_4__8063_, data_stage_4__8062_, data_stage_4__8061_, data_stage_4__8060_, data_stage_4__8059_, data_stage_4__8058_, data_stage_4__8057_, data_stage_4__8056_, data_stage_4__8055_, data_stage_4__8054_, data_stage_4__8053_, data_stage_4__8052_, data_stage_4__8051_, data_stage_4__8050_, data_stage_4__8049_, data_stage_4__8048_, data_stage_4__8047_, data_stage_4__8046_, data_stage_4__8045_, data_stage_4__8044_, data_stage_4__8043_, data_stage_4__8042_, data_stage_4__8041_, data_stage_4__8040_, data_stage_4__8039_, data_stage_4__8038_, data_stage_4__8037_, data_stage_4__8036_, data_stage_4__8035_, data_stage_4__8034_, data_stage_4__8033_, data_stage_4__8032_, data_stage_4__8031_, data_stage_4__8030_, data_stage_4__8029_, data_stage_4__8028_, data_stage_4__8027_, data_stage_4__8026_, data_stage_4__8025_, data_stage_4__8024_, data_stage_4__8023_, data_stage_4__8022_, data_stage_4__8021_, data_stage_4__8020_, data_stage_4__8019_, data_stage_4__8018_, data_stage_4__8017_, data_stage_4__8016_, data_stage_4__8015_, data_stage_4__8014_, data_stage_4__8013_, data_stage_4__8012_, data_stage_4__8011_, data_stage_4__8010_, data_stage_4__8009_, data_stage_4__8008_, data_stage_4__8007_, data_stage_4__8006_, data_stage_4__8005_, data_stage_4__8004_, data_stage_4__8003_, data_stage_4__8002_, data_stage_4__8001_, data_stage_4__8000_, data_stage_4__7999_, data_stage_4__7998_, data_stage_4__7997_, data_stage_4__7996_, data_stage_4__7995_, data_stage_4__7994_, data_stage_4__7993_, data_stage_4__7992_, data_stage_4__7991_, data_stage_4__7990_, data_stage_4__7989_, data_stage_4__7988_, data_stage_4__7987_, data_stage_4__7986_, data_stage_4__7985_, data_stage_4__7984_, data_stage_4__7983_, data_stage_4__7982_, data_stage_4__7981_, data_stage_4__7980_, data_stage_4__7979_, data_stage_4__7978_, data_stage_4__7977_, data_stage_4__7976_, data_stage_4__7975_, data_stage_4__7974_, data_stage_4__7973_, data_stage_4__7972_, data_stage_4__7971_, data_stage_4__7970_, data_stage_4__7969_, data_stage_4__7968_, data_stage_4__7967_, data_stage_4__7966_, data_stage_4__7965_, data_stage_4__7964_, data_stage_4__7963_, data_stage_4__7962_, data_stage_4__7961_, data_stage_4__7960_, data_stage_4__7959_, data_stage_4__7958_, data_stage_4__7957_, data_stage_4__7956_, data_stage_4__7955_, data_stage_4__7954_, data_stage_4__7953_, data_stage_4__7952_, data_stage_4__7951_, data_stage_4__7950_, data_stage_4__7949_, data_stage_4__7948_, data_stage_4__7947_, data_stage_4__7946_, data_stage_4__7945_, data_stage_4__7944_, data_stage_4__7943_, data_stage_4__7942_, data_stage_4__7941_, data_stage_4__7940_, data_stage_4__7939_, data_stage_4__7938_, data_stage_4__7937_, data_stage_4__7936_, data_stage_4__7935_, data_stage_4__7934_, data_stage_4__7933_, data_stage_4__7932_, data_stage_4__7931_, data_stage_4__7930_, data_stage_4__7929_, data_stage_4__7928_, data_stage_4__7927_, data_stage_4__7926_, data_stage_4__7925_, data_stage_4__7924_, data_stage_4__7923_, data_stage_4__7922_, data_stage_4__7921_, data_stage_4__7920_, data_stage_4__7919_, data_stage_4__7918_, data_stage_4__7917_, data_stage_4__7916_, data_stage_4__7915_, data_stage_4__7914_, data_stage_4__7913_, data_stage_4__7912_, data_stage_4__7911_, data_stage_4__7910_, data_stage_4__7909_, data_stage_4__7908_, data_stage_4__7907_, data_stage_4__7906_, data_stage_4__7905_, data_stage_4__7904_, data_stage_4__7903_, data_stage_4__7902_, data_stage_4__7901_, data_stage_4__7900_, data_stage_4__7899_, data_stage_4__7898_, data_stage_4__7897_, data_stage_4__7896_, data_stage_4__7895_, data_stage_4__7894_, data_stage_4__7893_, data_stage_4__7892_, data_stage_4__7891_, data_stage_4__7890_, data_stage_4__7889_, data_stage_4__7888_, data_stage_4__7887_, data_stage_4__7886_, data_stage_4__7885_, data_stage_4__7884_, data_stage_4__7883_, data_stage_4__7882_, data_stage_4__7881_, data_stage_4__7880_, data_stage_4__7879_, data_stage_4__7878_, data_stage_4__7877_, data_stage_4__7876_, data_stage_4__7875_, data_stage_4__7874_, data_stage_4__7873_, data_stage_4__7872_, data_stage_4__7871_, data_stage_4__7870_, data_stage_4__7869_, data_stage_4__7868_, data_stage_4__7867_, data_stage_4__7866_, data_stage_4__7865_, data_stage_4__7864_, data_stage_4__7863_, data_stage_4__7862_, data_stage_4__7861_, data_stage_4__7860_, data_stage_4__7859_, data_stage_4__7858_, data_stage_4__7857_, data_stage_4__7856_, data_stage_4__7855_, data_stage_4__7854_, data_stage_4__7853_, data_stage_4__7852_, data_stage_4__7851_, data_stage_4__7850_, data_stage_4__7849_, data_stage_4__7848_, data_stage_4__7847_, data_stage_4__7846_, data_stage_4__7845_, data_stage_4__7844_, data_stage_4__7843_, data_stage_4__7842_, data_stage_4__7841_, data_stage_4__7840_, data_stage_4__7839_, data_stage_4__7838_, data_stage_4__7837_, data_stage_4__7836_, data_stage_4__7835_, data_stage_4__7834_, data_stage_4__7833_, data_stage_4__7832_, data_stage_4__7831_, data_stage_4__7830_, data_stage_4__7829_, data_stage_4__7828_, data_stage_4__7827_, data_stage_4__7826_, data_stage_4__7825_, data_stage_4__7824_, data_stage_4__7823_, data_stage_4__7822_, data_stage_4__7821_, data_stage_4__7820_, data_stage_4__7819_, data_stage_4__7818_, data_stage_4__7817_, data_stage_4__7816_, data_stage_4__7815_, data_stage_4__7814_, data_stage_4__7813_, data_stage_4__7812_, data_stage_4__7811_, data_stage_4__7810_, data_stage_4__7809_, data_stage_4__7808_, data_stage_4__7807_, data_stage_4__7806_, data_stage_4__7805_, data_stage_4__7804_, data_stage_4__7803_, data_stage_4__7802_, data_stage_4__7801_, data_stage_4__7800_, data_stage_4__7799_, data_stage_4__7798_, data_stage_4__7797_, data_stage_4__7796_, data_stage_4__7795_, data_stage_4__7794_, data_stage_4__7793_, data_stage_4__7792_, data_stage_4__7791_, data_stage_4__7790_, data_stage_4__7789_, data_stage_4__7788_, data_stage_4__7787_, data_stage_4__7786_, data_stage_4__7785_, data_stage_4__7784_, data_stage_4__7783_, data_stage_4__7782_, data_stage_4__7781_, data_stage_4__7780_, data_stage_4__7779_, data_stage_4__7778_, data_stage_4__7777_, data_stage_4__7776_, data_stage_4__7775_, data_stage_4__7774_, data_stage_4__7773_, data_stage_4__7772_, data_stage_4__7771_, data_stage_4__7770_, data_stage_4__7769_, data_stage_4__7768_, data_stage_4__7767_, data_stage_4__7766_, data_stage_4__7765_, data_stage_4__7764_, data_stage_4__7763_, data_stage_4__7762_, data_stage_4__7761_, data_stage_4__7760_, data_stage_4__7759_, data_stage_4__7758_, data_stage_4__7757_, data_stage_4__7756_, data_stage_4__7755_, data_stage_4__7754_, data_stage_4__7753_, data_stage_4__7752_, data_stage_4__7751_, data_stage_4__7750_, data_stage_4__7749_, data_stage_4__7748_, data_stage_4__7747_, data_stage_4__7746_, data_stage_4__7745_, data_stage_4__7744_, data_stage_4__7743_, data_stage_4__7742_, data_stage_4__7741_, data_stage_4__7740_, data_stage_4__7739_, data_stage_4__7738_, data_stage_4__7737_, data_stage_4__7736_, data_stage_4__7735_, data_stage_4__7734_, data_stage_4__7733_, data_stage_4__7732_, data_stage_4__7731_, data_stage_4__7730_, data_stage_4__7729_, data_stage_4__7728_, data_stage_4__7727_, data_stage_4__7726_, data_stage_4__7725_, data_stage_4__7724_, data_stage_4__7723_, data_stage_4__7722_, data_stage_4__7721_, data_stage_4__7720_, data_stage_4__7719_, data_stage_4__7718_, data_stage_4__7717_, data_stage_4__7716_, data_stage_4__7715_, data_stage_4__7714_, data_stage_4__7713_, data_stage_4__7712_, data_stage_4__7711_, data_stage_4__7710_, data_stage_4__7709_, data_stage_4__7708_, data_stage_4__7707_, data_stage_4__7706_, data_stage_4__7705_, data_stage_4__7704_, data_stage_4__7703_, data_stage_4__7702_, data_stage_4__7701_, data_stage_4__7700_, data_stage_4__7699_, data_stage_4__7698_, data_stage_4__7697_, data_stage_4__7696_, data_stage_4__7695_, data_stage_4__7694_, data_stage_4__7693_, data_stage_4__7692_, data_stage_4__7691_, data_stage_4__7690_, data_stage_4__7689_, data_stage_4__7688_, data_stage_4__7687_, data_stage_4__7686_, data_stage_4__7685_, data_stage_4__7684_, data_stage_4__7683_, data_stage_4__7682_, data_stage_4__7681_, data_stage_4__7680_, data_stage_4__7679_, data_stage_4__7678_, data_stage_4__7677_, data_stage_4__7676_, data_stage_4__7675_, data_stage_4__7674_, data_stage_4__7673_, data_stage_4__7672_, data_stage_4__7671_, data_stage_4__7670_, data_stage_4__7669_, data_stage_4__7668_, data_stage_4__7667_, data_stage_4__7666_, data_stage_4__7665_, data_stage_4__7664_, data_stage_4__7663_, data_stage_4__7662_, data_stage_4__7661_, data_stage_4__7660_, data_stage_4__7659_, data_stage_4__7658_, data_stage_4__7657_, data_stage_4__7656_, data_stage_4__7655_, data_stage_4__7654_, data_stage_4__7653_, data_stage_4__7652_, data_stage_4__7651_, data_stage_4__7650_, data_stage_4__7649_, data_stage_4__7648_, data_stage_4__7647_, data_stage_4__7646_, data_stage_4__7645_, data_stage_4__7644_, data_stage_4__7643_, data_stage_4__7642_, data_stage_4__7641_, data_stage_4__7640_, data_stage_4__7639_, data_stage_4__7638_, data_stage_4__7637_, data_stage_4__7636_, data_stage_4__7635_, data_stage_4__7634_, data_stage_4__7633_, data_stage_4__7632_, data_stage_4__7631_, data_stage_4__7630_, data_stage_4__7629_, data_stage_4__7628_, data_stage_4__7627_, data_stage_4__7626_, data_stage_4__7625_, data_stage_4__7624_, data_stage_4__7623_, data_stage_4__7622_, data_stage_4__7621_, data_stage_4__7620_, data_stage_4__7619_, data_stage_4__7618_, data_stage_4__7617_, data_stage_4__7616_, data_stage_4__7615_, data_stage_4__7614_, data_stage_4__7613_, data_stage_4__7612_, data_stage_4__7611_, data_stage_4__7610_, data_stage_4__7609_, data_stage_4__7608_, data_stage_4__7607_, data_stage_4__7606_, data_stage_4__7605_, data_stage_4__7604_, data_stage_4__7603_, data_stage_4__7602_, data_stage_4__7601_, data_stage_4__7600_, data_stage_4__7599_, data_stage_4__7598_, data_stage_4__7597_, data_stage_4__7596_, data_stage_4__7595_, data_stage_4__7594_, data_stage_4__7593_, data_stage_4__7592_, data_stage_4__7591_, data_stage_4__7590_, data_stage_4__7589_, data_stage_4__7588_, data_stage_4__7587_, data_stage_4__7586_, data_stage_4__7585_, data_stage_4__7584_, data_stage_4__7583_, data_stage_4__7582_, data_stage_4__7581_, data_stage_4__7580_, data_stage_4__7579_, data_stage_4__7578_, data_stage_4__7577_, data_stage_4__7576_, data_stage_4__7575_, data_stage_4__7574_, data_stage_4__7573_, data_stage_4__7572_, data_stage_4__7571_, data_stage_4__7570_, data_stage_4__7569_, data_stage_4__7568_, data_stage_4__7567_, data_stage_4__7566_, data_stage_4__7565_, data_stage_4__7564_, data_stage_4__7563_, data_stage_4__7562_, data_stage_4__7561_, data_stage_4__7560_, data_stage_4__7559_, data_stage_4__7558_, data_stage_4__7557_, data_stage_4__7556_, data_stage_4__7555_, data_stage_4__7554_, data_stage_4__7553_, data_stage_4__7552_, data_stage_4__7551_, data_stage_4__7550_, data_stage_4__7549_, data_stage_4__7548_, data_stage_4__7547_, data_stage_4__7546_, data_stage_4__7545_, data_stage_4__7544_, data_stage_4__7543_, data_stage_4__7542_, data_stage_4__7541_, data_stage_4__7540_, data_stage_4__7539_, data_stage_4__7538_, data_stage_4__7537_, data_stage_4__7536_, data_stage_4__7535_, data_stage_4__7534_, data_stage_4__7533_, data_stage_4__7532_, data_stage_4__7531_, data_stage_4__7530_, data_stage_4__7529_, data_stage_4__7528_, data_stage_4__7527_, data_stage_4__7526_, data_stage_4__7525_, data_stage_4__7524_, data_stage_4__7523_, data_stage_4__7522_, data_stage_4__7521_, data_stage_4__7520_, data_stage_4__7519_, data_stage_4__7518_, data_stage_4__7517_, data_stage_4__7516_, data_stage_4__7515_, data_stage_4__7514_, data_stage_4__7513_, data_stage_4__7512_, data_stage_4__7511_, data_stage_4__7510_, data_stage_4__7509_, data_stage_4__7508_, data_stage_4__7507_, data_stage_4__7506_, data_stage_4__7505_, data_stage_4__7504_, data_stage_4__7503_, data_stage_4__7502_, data_stage_4__7501_, data_stage_4__7500_, data_stage_4__7499_, data_stage_4__7498_, data_stage_4__7497_, data_stage_4__7496_, data_stage_4__7495_, data_stage_4__7494_, data_stage_4__7493_, data_stage_4__7492_, data_stage_4__7491_, data_stage_4__7490_, data_stage_4__7489_, data_stage_4__7488_, data_stage_4__7487_, data_stage_4__7486_, data_stage_4__7485_, data_stage_4__7484_, data_stage_4__7483_, data_stage_4__7482_, data_stage_4__7481_, data_stage_4__7480_, data_stage_4__7479_, data_stage_4__7478_, data_stage_4__7477_, data_stage_4__7476_, data_stage_4__7475_, data_stage_4__7474_, data_stage_4__7473_, data_stage_4__7472_, data_stage_4__7471_, data_stage_4__7470_, data_stage_4__7469_, data_stage_4__7468_, data_stage_4__7467_, data_stage_4__7466_, data_stage_4__7465_, data_stage_4__7464_, data_stage_4__7463_, data_stage_4__7462_, data_stage_4__7461_, data_stage_4__7460_, data_stage_4__7459_, data_stage_4__7458_, data_stage_4__7457_, data_stage_4__7456_, data_stage_4__7455_, data_stage_4__7454_, data_stage_4__7453_, data_stage_4__7452_, data_stage_4__7451_, data_stage_4__7450_, data_stage_4__7449_, data_stage_4__7448_, data_stage_4__7447_, data_stage_4__7446_, data_stage_4__7445_, data_stage_4__7444_, data_stage_4__7443_, data_stage_4__7442_, data_stage_4__7441_, data_stage_4__7440_, data_stage_4__7439_, data_stage_4__7438_, data_stage_4__7437_, data_stage_4__7436_, data_stage_4__7435_, data_stage_4__7434_, data_stage_4__7433_, data_stage_4__7432_, data_stage_4__7431_, data_stage_4__7430_, data_stage_4__7429_, data_stage_4__7428_, data_stage_4__7427_, data_stage_4__7426_, data_stage_4__7425_, data_stage_4__7424_, data_stage_4__7423_, data_stage_4__7422_, data_stage_4__7421_, data_stage_4__7420_, data_stage_4__7419_, data_stage_4__7418_, data_stage_4__7417_, data_stage_4__7416_, data_stage_4__7415_, data_stage_4__7414_, data_stage_4__7413_, data_stage_4__7412_, data_stage_4__7411_, data_stage_4__7410_, data_stage_4__7409_, data_stage_4__7408_, data_stage_4__7407_, data_stage_4__7406_, data_stage_4__7405_, data_stage_4__7404_, data_stage_4__7403_, data_stage_4__7402_, data_stage_4__7401_, data_stage_4__7400_, data_stage_4__7399_, data_stage_4__7398_, data_stage_4__7397_, data_stage_4__7396_, data_stage_4__7395_, data_stage_4__7394_, data_stage_4__7393_, data_stage_4__7392_, data_stage_4__7391_, data_stage_4__7390_, data_stage_4__7389_, data_stage_4__7388_, data_stage_4__7387_, data_stage_4__7386_, data_stage_4__7385_, data_stage_4__7384_, data_stage_4__7383_, data_stage_4__7382_, data_stage_4__7381_, data_stage_4__7380_, data_stage_4__7379_, data_stage_4__7378_, data_stage_4__7377_, data_stage_4__7376_, data_stage_4__7375_, data_stage_4__7374_, data_stage_4__7373_, data_stage_4__7372_, data_stage_4__7371_, data_stage_4__7370_, data_stage_4__7369_, data_stage_4__7368_, data_stage_4__7367_, data_stage_4__7366_, data_stage_4__7365_, data_stage_4__7364_, data_stage_4__7363_, data_stage_4__7362_, data_stage_4__7361_, data_stage_4__7360_, data_stage_4__7359_, data_stage_4__7358_, data_stage_4__7357_, data_stage_4__7356_, data_stage_4__7355_, data_stage_4__7354_, data_stage_4__7353_, data_stage_4__7352_, data_stage_4__7351_, data_stage_4__7350_, data_stage_4__7349_, data_stage_4__7348_, data_stage_4__7347_, data_stage_4__7346_, data_stage_4__7345_, data_stage_4__7344_, data_stage_4__7343_, data_stage_4__7342_, data_stage_4__7341_, data_stage_4__7340_, data_stage_4__7339_, data_stage_4__7338_, data_stage_4__7337_, data_stage_4__7336_, data_stage_4__7335_, data_stage_4__7334_, data_stage_4__7333_, data_stage_4__7332_, data_stage_4__7331_, data_stage_4__7330_, data_stage_4__7329_, data_stage_4__7328_, data_stage_4__7327_, data_stage_4__7326_, data_stage_4__7325_, data_stage_4__7324_, data_stage_4__7323_, data_stage_4__7322_, data_stage_4__7321_, data_stage_4__7320_, data_stage_4__7319_, data_stage_4__7318_, data_stage_4__7317_, data_stage_4__7316_, data_stage_4__7315_, data_stage_4__7314_, data_stage_4__7313_, data_stage_4__7312_, data_stage_4__7311_, data_stage_4__7310_, data_stage_4__7309_, data_stage_4__7308_, data_stage_4__7307_, data_stage_4__7306_, data_stage_4__7305_, data_stage_4__7304_, data_stage_4__7303_, data_stage_4__7302_, data_stage_4__7301_, data_stage_4__7300_, data_stage_4__7299_, data_stage_4__7298_, data_stage_4__7297_, data_stage_4__7296_, data_stage_4__7295_, data_stage_4__7294_, data_stage_4__7293_, data_stage_4__7292_, data_stage_4__7291_, data_stage_4__7290_, data_stage_4__7289_, data_stage_4__7288_, data_stage_4__7287_, data_stage_4__7286_, data_stage_4__7285_, data_stage_4__7284_, data_stage_4__7283_, data_stage_4__7282_, data_stage_4__7281_, data_stage_4__7280_, data_stage_4__7279_, data_stage_4__7278_, data_stage_4__7277_, data_stage_4__7276_, data_stage_4__7275_, data_stage_4__7274_, data_stage_4__7273_, data_stage_4__7272_, data_stage_4__7271_, data_stage_4__7270_, data_stage_4__7269_, data_stage_4__7268_, data_stage_4__7267_, data_stage_4__7266_, data_stage_4__7265_, data_stage_4__7264_, data_stage_4__7263_, data_stage_4__7262_, data_stage_4__7261_, data_stage_4__7260_, data_stage_4__7259_, data_stage_4__7258_, data_stage_4__7257_, data_stage_4__7256_, data_stage_4__7255_, data_stage_4__7254_, data_stage_4__7253_, data_stage_4__7252_, data_stage_4__7251_, data_stage_4__7250_, data_stage_4__7249_, data_stage_4__7248_, data_stage_4__7247_, data_stage_4__7246_, data_stage_4__7245_, data_stage_4__7244_, data_stage_4__7243_, data_stage_4__7242_, data_stage_4__7241_, data_stage_4__7240_, data_stage_4__7239_, data_stage_4__7238_, data_stage_4__7237_, data_stage_4__7236_, data_stage_4__7235_, data_stage_4__7234_, data_stage_4__7233_, data_stage_4__7232_, data_stage_4__7231_, data_stage_4__7230_, data_stage_4__7229_, data_stage_4__7228_, data_stage_4__7227_, data_stage_4__7226_, data_stage_4__7225_, data_stage_4__7224_, data_stage_4__7223_, data_stage_4__7222_, data_stage_4__7221_, data_stage_4__7220_, data_stage_4__7219_, data_stage_4__7218_, data_stage_4__7217_, data_stage_4__7216_, data_stage_4__7215_, data_stage_4__7214_, data_stage_4__7213_, data_stage_4__7212_, data_stage_4__7211_, data_stage_4__7210_, data_stage_4__7209_, data_stage_4__7208_, data_stage_4__7207_, data_stage_4__7206_, data_stage_4__7205_, data_stage_4__7204_, data_stage_4__7203_, data_stage_4__7202_, data_stage_4__7201_, data_stage_4__7200_, data_stage_4__7199_, data_stage_4__7198_, data_stage_4__7197_, data_stage_4__7196_, data_stage_4__7195_, data_stage_4__7194_, data_stage_4__7193_, data_stage_4__7192_, data_stage_4__7191_, data_stage_4__7190_, data_stage_4__7189_, data_stage_4__7188_, data_stage_4__7187_, data_stage_4__7186_, data_stage_4__7185_, data_stage_4__7184_, data_stage_4__7183_, data_stage_4__7182_, data_stage_4__7181_, data_stage_4__7180_, data_stage_4__7179_, data_stage_4__7178_, data_stage_4__7177_, data_stage_4__7176_, data_stage_4__7175_, data_stage_4__7174_, data_stage_4__7173_, data_stage_4__7172_, data_stage_4__7171_, data_stage_4__7170_, data_stage_4__7169_, data_stage_4__7168_, data_stage_4__7167_, data_stage_4__7166_, data_stage_4__7165_, data_stage_4__7164_, data_stage_4__7163_, data_stage_4__7162_, data_stage_4__7161_, data_stage_4__7160_, data_stage_4__7159_, data_stage_4__7158_, data_stage_4__7157_, data_stage_4__7156_, data_stage_4__7155_, data_stage_4__7154_, data_stage_4__7153_, data_stage_4__7152_, data_stage_4__7151_, data_stage_4__7150_, data_stage_4__7149_, data_stage_4__7148_, data_stage_4__7147_, data_stage_4__7146_, data_stage_4__7145_, data_stage_4__7144_, data_stage_4__7143_, data_stage_4__7142_, data_stage_4__7141_, data_stage_4__7140_, data_stage_4__7139_, data_stage_4__7138_, data_stage_4__7137_, data_stage_4__7136_, data_stage_4__7135_, data_stage_4__7134_, data_stage_4__7133_, data_stage_4__7132_, data_stage_4__7131_, data_stage_4__7130_, data_stage_4__7129_, data_stage_4__7128_, data_stage_4__7127_, data_stage_4__7126_, data_stage_4__7125_, data_stage_4__7124_, data_stage_4__7123_, data_stage_4__7122_, data_stage_4__7121_, data_stage_4__7120_, data_stage_4__7119_, data_stage_4__7118_, data_stage_4__7117_, data_stage_4__7116_, data_stage_4__7115_, data_stage_4__7114_, data_stage_4__7113_, data_stage_4__7112_, data_stage_4__7111_, data_stage_4__7110_, data_stage_4__7109_, data_stage_4__7108_, data_stage_4__7107_, data_stage_4__7106_, data_stage_4__7105_, data_stage_4__7104_, data_stage_4__7103_, data_stage_4__7102_, data_stage_4__7101_, data_stage_4__7100_, data_stage_4__7099_, data_stage_4__7098_, data_stage_4__7097_, data_stage_4__7096_, data_stage_4__7095_, data_stage_4__7094_, data_stage_4__7093_, data_stage_4__7092_, data_stage_4__7091_, data_stage_4__7090_, data_stage_4__7089_, data_stage_4__7088_, data_stage_4__7087_, data_stage_4__7086_, data_stage_4__7085_, data_stage_4__7084_, data_stage_4__7083_, data_stage_4__7082_, data_stage_4__7081_, data_stage_4__7080_, data_stage_4__7079_, data_stage_4__7078_, data_stage_4__7077_, data_stage_4__7076_, data_stage_4__7075_, data_stage_4__7074_, data_stage_4__7073_, data_stage_4__7072_, data_stage_4__7071_, data_stage_4__7070_, data_stage_4__7069_, data_stage_4__7068_, data_stage_4__7067_, data_stage_4__7066_, data_stage_4__7065_, data_stage_4__7064_, data_stage_4__7063_, data_stage_4__7062_, data_stage_4__7061_, data_stage_4__7060_, data_stage_4__7059_, data_stage_4__7058_, data_stage_4__7057_, data_stage_4__7056_, data_stage_4__7055_, data_stage_4__7054_, data_stage_4__7053_, data_stage_4__7052_, data_stage_4__7051_, data_stage_4__7050_, data_stage_4__7049_, data_stage_4__7048_, data_stage_4__7047_, data_stage_4__7046_, data_stage_4__7045_, data_stage_4__7044_, data_stage_4__7043_, data_stage_4__7042_, data_stage_4__7041_, data_stage_4__7040_, data_stage_4__7039_, data_stage_4__7038_, data_stage_4__7037_, data_stage_4__7036_, data_stage_4__7035_, data_stage_4__7034_, data_stage_4__7033_, data_stage_4__7032_, data_stage_4__7031_, data_stage_4__7030_, data_stage_4__7029_, data_stage_4__7028_, data_stage_4__7027_, data_stage_4__7026_, data_stage_4__7025_, data_stage_4__7024_, data_stage_4__7023_, data_stage_4__7022_, data_stage_4__7021_, data_stage_4__7020_, data_stage_4__7019_, data_stage_4__7018_, data_stage_4__7017_, data_stage_4__7016_, data_stage_4__7015_, data_stage_4__7014_, data_stage_4__7013_, data_stage_4__7012_, data_stage_4__7011_, data_stage_4__7010_, data_stage_4__7009_, data_stage_4__7008_, data_stage_4__7007_, data_stage_4__7006_, data_stage_4__7005_, data_stage_4__7004_, data_stage_4__7003_, data_stage_4__7002_, data_stage_4__7001_, data_stage_4__7000_, data_stage_4__6999_, data_stage_4__6998_, data_stage_4__6997_, data_stage_4__6996_, data_stage_4__6995_, data_stage_4__6994_, data_stage_4__6993_, data_stage_4__6992_, data_stage_4__6991_, data_stage_4__6990_, data_stage_4__6989_, data_stage_4__6988_, data_stage_4__6987_, data_stage_4__6986_, data_stage_4__6985_, data_stage_4__6984_, data_stage_4__6983_, data_stage_4__6982_, data_stage_4__6981_, data_stage_4__6980_, data_stage_4__6979_, data_stage_4__6978_, data_stage_4__6977_, data_stage_4__6976_, data_stage_4__6975_, data_stage_4__6974_, data_stage_4__6973_, data_stage_4__6972_, data_stage_4__6971_, data_stage_4__6970_, data_stage_4__6969_, data_stage_4__6968_, data_stage_4__6967_, data_stage_4__6966_, data_stage_4__6965_, data_stage_4__6964_, data_stage_4__6963_, data_stage_4__6962_, data_stage_4__6961_, data_stage_4__6960_, data_stage_4__6959_, data_stage_4__6958_, data_stage_4__6957_, data_stage_4__6956_, data_stage_4__6955_, data_stage_4__6954_, data_stage_4__6953_, data_stage_4__6952_, data_stage_4__6951_, data_stage_4__6950_, data_stage_4__6949_, data_stage_4__6948_, data_stage_4__6947_, data_stage_4__6946_, data_stage_4__6945_, data_stage_4__6944_, data_stage_4__6943_, data_stage_4__6942_, data_stage_4__6941_, data_stage_4__6940_, data_stage_4__6939_, data_stage_4__6938_, data_stage_4__6937_, data_stage_4__6936_, data_stage_4__6935_, data_stage_4__6934_, data_stage_4__6933_, data_stage_4__6932_, data_stage_4__6931_, data_stage_4__6930_, data_stage_4__6929_, data_stage_4__6928_, data_stage_4__6927_, data_stage_4__6926_, data_stage_4__6925_, data_stage_4__6924_, data_stage_4__6923_, data_stage_4__6922_, data_stage_4__6921_, data_stage_4__6920_, data_stage_4__6919_, data_stage_4__6918_, data_stage_4__6917_, data_stage_4__6916_, data_stage_4__6915_, data_stage_4__6914_, data_stage_4__6913_, data_stage_4__6912_, data_stage_4__6911_, data_stage_4__6910_, data_stage_4__6909_, data_stage_4__6908_, data_stage_4__6907_, data_stage_4__6906_, data_stage_4__6905_, data_stage_4__6904_, data_stage_4__6903_, data_stage_4__6902_, data_stage_4__6901_, data_stage_4__6900_, data_stage_4__6899_, data_stage_4__6898_, data_stage_4__6897_, data_stage_4__6896_, data_stage_4__6895_, data_stage_4__6894_, data_stage_4__6893_, data_stage_4__6892_, data_stage_4__6891_, data_stage_4__6890_, data_stage_4__6889_, data_stage_4__6888_, data_stage_4__6887_, data_stage_4__6886_, data_stage_4__6885_, data_stage_4__6884_, data_stage_4__6883_, data_stage_4__6882_, data_stage_4__6881_, data_stage_4__6880_, data_stage_4__6879_, data_stage_4__6878_, data_stage_4__6877_, data_stage_4__6876_, data_stage_4__6875_, data_stage_4__6874_, data_stage_4__6873_, data_stage_4__6872_, data_stage_4__6871_, data_stage_4__6870_, data_stage_4__6869_, data_stage_4__6868_, data_stage_4__6867_, data_stage_4__6866_, data_stage_4__6865_, data_stage_4__6864_, data_stage_4__6863_, data_stage_4__6862_, data_stage_4__6861_, data_stage_4__6860_, data_stage_4__6859_, data_stage_4__6858_, data_stage_4__6857_, data_stage_4__6856_, data_stage_4__6855_, data_stage_4__6854_, data_stage_4__6853_, data_stage_4__6852_, data_stage_4__6851_, data_stage_4__6850_, data_stage_4__6849_, data_stage_4__6848_, data_stage_4__6847_, data_stage_4__6846_, data_stage_4__6845_, data_stage_4__6844_, data_stage_4__6843_, data_stage_4__6842_, data_stage_4__6841_, data_stage_4__6840_, data_stage_4__6839_, data_stage_4__6838_, data_stage_4__6837_, data_stage_4__6836_, data_stage_4__6835_, data_stage_4__6834_, data_stage_4__6833_, data_stage_4__6832_, data_stage_4__6831_, data_stage_4__6830_, data_stage_4__6829_, data_stage_4__6828_, data_stage_4__6827_, data_stage_4__6826_, data_stage_4__6825_, data_stage_4__6824_, data_stage_4__6823_, data_stage_4__6822_, data_stage_4__6821_, data_stage_4__6820_, data_stage_4__6819_, data_stage_4__6818_, data_stage_4__6817_, data_stage_4__6816_, data_stage_4__6815_, data_stage_4__6814_, data_stage_4__6813_, data_stage_4__6812_, data_stage_4__6811_, data_stage_4__6810_, data_stage_4__6809_, data_stage_4__6808_, data_stage_4__6807_, data_stage_4__6806_, data_stage_4__6805_, data_stage_4__6804_, data_stage_4__6803_, data_stage_4__6802_, data_stage_4__6801_, data_stage_4__6800_, data_stage_4__6799_, data_stage_4__6798_, data_stage_4__6797_, data_stage_4__6796_, data_stage_4__6795_, data_stage_4__6794_, data_stage_4__6793_, data_stage_4__6792_, data_stage_4__6791_, data_stage_4__6790_, data_stage_4__6789_, data_stage_4__6788_, data_stage_4__6787_, data_stage_4__6786_, data_stage_4__6785_, data_stage_4__6784_, data_stage_4__6783_, data_stage_4__6782_, data_stage_4__6781_, data_stage_4__6780_, data_stage_4__6779_, data_stage_4__6778_, data_stage_4__6777_, data_stage_4__6776_, data_stage_4__6775_, data_stage_4__6774_, data_stage_4__6773_, data_stage_4__6772_, data_stage_4__6771_, data_stage_4__6770_, data_stage_4__6769_, data_stage_4__6768_, data_stage_4__6767_, data_stage_4__6766_, data_stage_4__6765_, data_stage_4__6764_, data_stage_4__6763_, data_stage_4__6762_, data_stage_4__6761_, data_stage_4__6760_, data_stage_4__6759_, data_stage_4__6758_, data_stage_4__6757_, data_stage_4__6756_, data_stage_4__6755_, data_stage_4__6754_, data_stage_4__6753_, data_stage_4__6752_, data_stage_4__6751_, data_stage_4__6750_, data_stage_4__6749_, data_stage_4__6748_, data_stage_4__6747_, data_stage_4__6746_, data_stage_4__6745_, data_stage_4__6744_, data_stage_4__6743_, data_stage_4__6742_, data_stage_4__6741_, data_stage_4__6740_, data_stage_4__6739_, data_stage_4__6738_, data_stage_4__6737_, data_stage_4__6736_, data_stage_4__6735_, data_stage_4__6734_, data_stage_4__6733_, data_stage_4__6732_, data_stage_4__6731_, data_stage_4__6730_, data_stage_4__6729_, data_stage_4__6728_, data_stage_4__6727_, data_stage_4__6726_, data_stage_4__6725_, data_stage_4__6724_, data_stage_4__6723_, data_stage_4__6722_, data_stage_4__6721_, data_stage_4__6720_, data_stage_4__6719_, data_stage_4__6718_, data_stage_4__6717_, data_stage_4__6716_, data_stage_4__6715_, data_stage_4__6714_, data_stage_4__6713_, data_stage_4__6712_, data_stage_4__6711_, data_stage_4__6710_, data_stage_4__6709_, data_stage_4__6708_, data_stage_4__6707_, data_stage_4__6706_, data_stage_4__6705_, data_stage_4__6704_, data_stage_4__6703_, data_stage_4__6702_, data_stage_4__6701_, data_stage_4__6700_, data_stage_4__6699_, data_stage_4__6698_, data_stage_4__6697_, data_stage_4__6696_, data_stage_4__6695_, data_stage_4__6694_, data_stage_4__6693_, data_stage_4__6692_, data_stage_4__6691_, data_stage_4__6690_, data_stage_4__6689_, data_stage_4__6688_, data_stage_4__6687_, data_stage_4__6686_, data_stage_4__6685_, data_stage_4__6684_, data_stage_4__6683_, data_stage_4__6682_, data_stage_4__6681_, data_stage_4__6680_, data_stage_4__6679_, data_stage_4__6678_, data_stage_4__6677_, data_stage_4__6676_, data_stage_4__6675_, data_stage_4__6674_, data_stage_4__6673_, data_stage_4__6672_, data_stage_4__6671_, data_stage_4__6670_, data_stage_4__6669_, data_stage_4__6668_, data_stage_4__6667_, data_stage_4__6666_, data_stage_4__6665_, data_stage_4__6664_, data_stage_4__6663_, data_stage_4__6662_, data_stage_4__6661_, data_stage_4__6660_, data_stage_4__6659_, data_stage_4__6658_, data_stage_4__6657_, data_stage_4__6656_, data_stage_4__6655_, data_stage_4__6654_, data_stage_4__6653_, data_stage_4__6652_, data_stage_4__6651_, data_stage_4__6650_, data_stage_4__6649_, data_stage_4__6648_, data_stage_4__6647_, data_stage_4__6646_, data_stage_4__6645_, data_stage_4__6644_, data_stage_4__6643_, data_stage_4__6642_, data_stage_4__6641_, data_stage_4__6640_, data_stage_4__6639_, data_stage_4__6638_, data_stage_4__6637_, data_stage_4__6636_, data_stage_4__6635_, data_stage_4__6634_, data_stage_4__6633_, data_stage_4__6632_, data_stage_4__6631_, data_stage_4__6630_, data_stage_4__6629_, data_stage_4__6628_, data_stage_4__6627_, data_stage_4__6626_, data_stage_4__6625_, data_stage_4__6624_, data_stage_4__6623_, data_stage_4__6622_, data_stage_4__6621_, data_stage_4__6620_, data_stage_4__6619_, data_stage_4__6618_, data_stage_4__6617_, data_stage_4__6616_, data_stage_4__6615_, data_stage_4__6614_, data_stage_4__6613_, data_stage_4__6612_, data_stage_4__6611_, data_stage_4__6610_, data_stage_4__6609_, data_stage_4__6608_, data_stage_4__6607_, data_stage_4__6606_, data_stage_4__6605_, data_stage_4__6604_, data_stage_4__6603_, data_stage_4__6602_, data_stage_4__6601_, data_stage_4__6600_, data_stage_4__6599_, data_stage_4__6598_, data_stage_4__6597_, data_stage_4__6596_, data_stage_4__6595_, data_stage_4__6594_, data_stage_4__6593_, data_stage_4__6592_, data_stage_4__6591_, data_stage_4__6590_, data_stage_4__6589_, data_stage_4__6588_, data_stage_4__6587_, data_stage_4__6586_, data_stage_4__6585_, data_stage_4__6584_, data_stage_4__6583_, data_stage_4__6582_, data_stage_4__6581_, data_stage_4__6580_, data_stage_4__6579_, data_stage_4__6578_, data_stage_4__6577_, data_stage_4__6576_, data_stage_4__6575_, data_stage_4__6574_, data_stage_4__6573_, data_stage_4__6572_, data_stage_4__6571_, data_stage_4__6570_, data_stage_4__6569_, data_stage_4__6568_, data_stage_4__6567_, data_stage_4__6566_, data_stage_4__6565_, data_stage_4__6564_, data_stage_4__6563_, data_stage_4__6562_, data_stage_4__6561_, data_stage_4__6560_, data_stage_4__6559_, data_stage_4__6558_, data_stage_4__6557_, data_stage_4__6556_, data_stage_4__6555_, data_stage_4__6554_, data_stage_4__6553_, data_stage_4__6552_, data_stage_4__6551_, data_stage_4__6550_, data_stage_4__6549_, data_stage_4__6548_, data_stage_4__6547_, data_stage_4__6546_, data_stage_4__6545_, data_stage_4__6544_, data_stage_4__6543_, data_stage_4__6542_, data_stage_4__6541_, data_stage_4__6540_, data_stage_4__6539_, data_stage_4__6538_, data_stage_4__6537_, data_stage_4__6536_, data_stage_4__6535_, data_stage_4__6534_, data_stage_4__6533_, data_stage_4__6532_, data_stage_4__6531_, data_stage_4__6530_, data_stage_4__6529_, data_stage_4__6528_, data_stage_4__6527_, data_stage_4__6526_, data_stage_4__6525_, data_stage_4__6524_, data_stage_4__6523_, data_stage_4__6522_, data_stage_4__6521_, data_stage_4__6520_, data_stage_4__6519_, data_stage_4__6518_, data_stage_4__6517_, data_stage_4__6516_, data_stage_4__6515_, data_stage_4__6514_, data_stage_4__6513_, data_stage_4__6512_, data_stage_4__6511_, data_stage_4__6510_, data_stage_4__6509_, data_stage_4__6508_, data_stage_4__6507_, data_stage_4__6506_, data_stage_4__6505_, data_stage_4__6504_, data_stage_4__6503_, data_stage_4__6502_, data_stage_4__6501_, data_stage_4__6500_, data_stage_4__6499_, data_stage_4__6498_, data_stage_4__6497_, data_stage_4__6496_, data_stage_4__6495_, data_stage_4__6494_, data_stage_4__6493_, data_stage_4__6492_, data_stage_4__6491_, data_stage_4__6490_, data_stage_4__6489_, data_stage_4__6488_, data_stage_4__6487_, data_stage_4__6486_, data_stage_4__6485_, data_stage_4__6484_, data_stage_4__6483_, data_stage_4__6482_, data_stage_4__6481_, data_stage_4__6480_, data_stage_4__6479_, data_stage_4__6478_, data_stage_4__6477_, data_stage_4__6476_, data_stage_4__6475_, data_stage_4__6474_, data_stage_4__6473_, data_stage_4__6472_, data_stage_4__6471_, data_stage_4__6470_, data_stage_4__6469_, data_stage_4__6468_, data_stage_4__6467_, data_stage_4__6466_, data_stage_4__6465_, data_stage_4__6464_, data_stage_4__6463_, data_stage_4__6462_, data_stage_4__6461_, data_stage_4__6460_, data_stage_4__6459_, data_stage_4__6458_, data_stage_4__6457_, data_stage_4__6456_, data_stage_4__6455_, data_stage_4__6454_, data_stage_4__6453_, data_stage_4__6452_, data_stage_4__6451_, data_stage_4__6450_, data_stage_4__6449_, data_stage_4__6448_, data_stage_4__6447_, data_stage_4__6446_, data_stage_4__6445_, data_stage_4__6444_, data_stage_4__6443_, data_stage_4__6442_, data_stage_4__6441_, data_stage_4__6440_, data_stage_4__6439_, data_stage_4__6438_, data_stage_4__6437_, data_stage_4__6436_, data_stage_4__6435_, data_stage_4__6434_, data_stage_4__6433_, data_stage_4__6432_, data_stage_4__6431_, data_stage_4__6430_, data_stage_4__6429_, data_stage_4__6428_, data_stage_4__6427_, data_stage_4__6426_, data_stage_4__6425_, data_stage_4__6424_, data_stage_4__6423_, data_stage_4__6422_, data_stage_4__6421_, data_stage_4__6420_, data_stage_4__6419_, data_stage_4__6418_, data_stage_4__6417_, data_stage_4__6416_, data_stage_4__6415_, data_stage_4__6414_, data_stage_4__6413_, data_stage_4__6412_, data_stage_4__6411_, data_stage_4__6410_, data_stage_4__6409_, data_stage_4__6408_, data_stage_4__6407_, data_stage_4__6406_, data_stage_4__6405_, data_stage_4__6404_, data_stage_4__6403_, data_stage_4__6402_, data_stage_4__6401_, data_stage_4__6400_, data_stage_4__6399_, data_stage_4__6398_, data_stage_4__6397_, data_stage_4__6396_, data_stage_4__6395_, data_stage_4__6394_, data_stage_4__6393_, data_stage_4__6392_, data_stage_4__6391_, data_stage_4__6390_, data_stage_4__6389_, data_stage_4__6388_, data_stage_4__6387_, data_stage_4__6386_, data_stage_4__6385_, data_stage_4__6384_, data_stage_4__6383_, data_stage_4__6382_, data_stage_4__6381_, data_stage_4__6380_, data_stage_4__6379_, data_stage_4__6378_, data_stage_4__6377_, data_stage_4__6376_, data_stage_4__6375_, data_stage_4__6374_, data_stage_4__6373_, data_stage_4__6372_, data_stage_4__6371_, data_stage_4__6370_, data_stage_4__6369_, data_stage_4__6368_, data_stage_4__6367_, data_stage_4__6366_, data_stage_4__6365_, data_stage_4__6364_, data_stage_4__6363_, data_stage_4__6362_, data_stage_4__6361_, data_stage_4__6360_, data_stage_4__6359_, data_stage_4__6358_, data_stage_4__6357_, data_stage_4__6356_, data_stage_4__6355_, data_stage_4__6354_, data_stage_4__6353_, data_stage_4__6352_, data_stage_4__6351_, data_stage_4__6350_, data_stage_4__6349_, data_stage_4__6348_, data_stage_4__6347_, data_stage_4__6346_, data_stage_4__6345_, data_stage_4__6344_, data_stage_4__6343_, data_stage_4__6342_, data_stage_4__6341_, data_stage_4__6340_, data_stage_4__6339_, data_stage_4__6338_, data_stage_4__6337_, data_stage_4__6336_, data_stage_4__6335_, data_stage_4__6334_, data_stage_4__6333_, data_stage_4__6332_, data_stage_4__6331_, data_stage_4__6330_, data_stage_4__6329_, data_stage_4__6328_, data_stage_4__6327_, data_stage_4__6326_, data_stage_4__6325_, data_stage_4__6324_, data_stage_4__6323_, data_stage_4__6322_, data_stage_4__6321_, data_stage_4__6320_, data_stage_4__6319_, data_stage_4__6318_, data_stage_4__6317_, data_stage_4__6316_, data_stage_4__6315_, data_stage_4__6314_, data_stage_4__6313_, data_stage_4__6312_, data_stage_4__6311_, data_stage_4__6310_, data_stage_4__6309_, data_stage_4__6308_, data_stage_4__6307_, data_stage_4__6306_, data_stage_4__6305_, data_stage_4__6304_, data_stage_4__6303_, data_stage_4__6302_, data_stage_4__6301_, data_stage_4__6300_, data_stage_4__6299_, data_stage_4__6298_, data_stage_4__6297_, data_stage_4__6296_, data_stage_4__6295_, data_stage_4__6294_, data_stage_4__6293_, data_stage_4__6292_, data_stage_4__6291_, data_stage_4__6290_, data_stage_4__6289_, data_stage_4__6288_, data_stage_4__6287_, data_stage_4__6286_, data_stage_4__6285_, data_stage_4__6284_, data_stage_4__6283_, data_stage_4__6282_, data_stage_4__6281_, data_stage_4__6280_, data_stage_4__6279_, data_stage_4__6278_, data_stage_4__6277_, data_stage_4__6276_, data_stage_4__6275_, data_stage_4__6274_, data_stage_4__6273_, data_stage_4__6272_, data_stage_4__6271_, data_stage_4__6270_, data_stage_4__6269_, data_stage_4__6268_, data_stage_4__6267_, data_stage_4__6266_, data_stage_4__6265_, data_stage_4__6264_, data_stage_4__6263_, data_stage_4__6262_, data_stage_4__6261_, data_stage_4__6260_, data_stage_4__6259_, data_stage_4__6258_, data_stage_4__6257_, data_stage_4__6256_, data_stage_4__6255_, data_stage_4__6254_, data_stage_4__6253_, data_stage_4__6252_, data_stage_4__6251_, data_stage_4__6250_, data_stage_4__6249_, data_stage_4__6248_, data_stage_4__6247_, data_stage_4__6246_, data_stage_4__6245_, data_stage_4__6244_, data_stage_4__6243_, data_stage_4__6242_, data_stage_4__6241_, data_stage_4__6240_, data_stage_4__6239_, data_stage_4__6238_, data_stage_4__6237_, data_stage_4__6236_, data_stage_4__6235_, data_stage_4__6234_, data_stage_4__6233_, data_stage_4__6232_, data_stage_4__6231_, data_stage_4__6230_, data_stage_4__6229_, data_stage_4__6228_, data_stage_4__6227_, data_stage_4__6226_, data_stage_4__6225_, data_stage_4__6224_, data_stage_4__6223_, data_stage_4__6222_, data_stage_4__6221_, data_stage_4__6220_, data_stage_4__6219_, data_stage_4__6218_, data_stage_4__6217_, data_stage_4__6216_, data_stage_4__6215_, data_stage_4__6214_, data_stage_4__6213_, data_stage_4__6212_, data_stage_4__6211_, data_stage_4__6210_, data_stage_4__6209_, data_stage_4__6208_, data_stage_4__6207_, data_stage_4__6206_, data_stage_4__6205_, data_stage_4__6204_, data_stage_4__6203_, data_stage_4__6202_, data_stage_4__6201_, data_stage_4__6200_, data_stage_4__6199_, data_stage_4__6198_, data_stage_4__6197_, data_stage_4__6196_, data_stage_4__6195_, data_stage_4__6194_, data_stage_4__6193_, data_stage_4__6192_, data_stage_4__6191_, data_stage_4__6190_, data_stage_4__6189_, data_stage_4__6188_, data_stage_4__6187_, data_stage_4__6186_, data_stage_4__6185_, data_stage_4__6184_, data_stage_4__6183_, data_stage_4__6182_, data_stage_4__6181_, data_stage_4__6180_, data_stage_4__6179_, data_stage_4__6178_, data_stage_4__6177_, data_stage_4__6176_, data_stage_4__6175_, data_stage_4__6174_, data_stage_4__6173_, data_stage_4__6172_, data_stage_4__6171_, data_stage_4__6170_, data_stage_4__6169_, data_stage_4__6168_, data_stage_4__6167_, data_stage_4__6166_, data_stage_4__6165_, data_stage_4__6164_, data_stage_4__6163_, data_stage_4__6162_, data_stage_4__6161_, data_stage_4__6160_, data_stage_4__6159_, data_stage_4__6158_, data_stage_4__6157_, data_stage_4__6156_, data_stage_4__6155_, data_stage_4__6154_, data_stage_4__6153_, data_stage_4__6152_, data_stage_4__6151_, data_stage_4__6150_, data_stage_4__6149_, data_stage_4__6148_, data_stage_4__6147_, data_stage_4__6146_, data_stage_4__6145_, data_stage_4__6144_ })
  );


  bsg_swap_width_p2048
  mux_stage_4__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_4__4095_, data_stage_4__4094_, data_stage_4__4093_, data_stage_4__4092_, data_stage_4__4091_, data_stage_4__4090_, data_stage_4__4089_, data_stage_4__4088_, data_stage_4__4087_, data_stage_4__4086_, data_stage_4__4085_, data_stage_4__4084_, data_stage_4__4083_, data_stage_4__4082_, data_stage_4__4081_, data_stage_4__4080_, data_stage_4__4079_, data_stage_4__4078_, data_stage_4__4077_, data_stage_4__4076_, data_stage_4__4075_, data_stage_4__4074_, data_stage_4__4073_, data_stage_4__4072_, data_stage_4__4071_, data_stage_4__4070_, data_stage_4__4069_, data_stage_4__4068_, data_stage_4__4067_, data_stage_4__4066_, data_stage_4__4065_, data_stage_4__4064_, data_stage_4__4063_, data_stage_4__4062_, data_stage_4__4061_, data_stage_4__4060_, data_stage_4__4059_, data_stage_4__4058_, data_stage_4__4057_, data_stage_4__4056_, data_stage_4__4055_, data_stage_4__4054_, data_stage_4__4053_, data_stage_4__4052_, data_stage_4__4051_, data_stage_4__4050_, data_stage_4__4049_, data_stage_4__4048_, data_stage_4__4047_, data_stage_4__4046_, data_stage_4__4045_, data_stage_4__4044_, data_stage_4__4043_, data_stage_4__4042_, data_stage_4__4041_, data_stage_4__4040_, data_stage_4__4039_, data_stage_4__4038_, data_stage_4__4037_, data_stage_4__4036_, data_stage_4__4035_, data_stage_4__4034_, data_stage_4__4033_, data_stage_4__4032_, data_stage_4__4031_, data_stage_4__4030_, data_stage_4__4029_, data_stage_4__4028_, data_stage_4__4027_, data_stage_4__4026_, data_stage_4__4025_, data_stage_4__4024_, data_stage_4__4023_, data_stage_4__4022_, data_stage_4__4021_, data_stage_4__4020_, data_stage_4__4019_, data_stage_4__4018_, data_stage_4__4017_, data_stage_4__4016_, data_stage_4__4015_, data_stage_4__4014_, data_stage_4__4013_, data_stage_4__4012_, data_stage_4__4011_, data_stage_4__4010_, data_stage_4__4009_, data_stage_4__4008_, data_stage_4__4007_, data_stage_4__4006_, data_stage_4__4005_, data_stage_4__4004_, data_stage_4__4003_, data_stage_4__4002_, data_stage_4__4001_, data_stage_4__4000_, data_stage_4__3999_, data_stage_4__3998_, data_stage_4__3997_, data_stage_4__3996_, data_stage_4__3995_, data_stage_4__3994_, data_stage_4__3993_, data_stage_4__3992_, data_stage_4__3991_, data_stage_4__3990_, data_stage_4__3989_, data_stage_4__3988_, data_stage_4__3987_, data_stage_4__3986_, data_stage_4__3985_, data_stage_4__3984_, data_stage_4__3983_, data_stage_4__3982_, data_stage_4__3981_, data_stage_4__3980_, data_stage_4__3979_, data_stage_4__3978_, data_stage_4__3977_, data_stage_4__3976_, data_stage_4__3975_, data_stage_4__3974_, data_stage_4__3973_, data_stage_4__3972_, data_stage_4__3971_, data_stage_4__3970_, data_stage_4__3969_, data_stage_4__3968_, data_stage_4__3967_, data_stage_4__3966_, data_stage_4__3965_, data_stage_4__3964_, data_stage_4__3963_, data_stage_4__3962_, data_stage_4__3961_, data_stage_4__3960_, data_stage_4__3959_, data_stage_4__3958_, data_stage_4__3957_, data_stage_4__3956_, data_stage_4__3955_, data_stage_4__3954_, data_stage_4__3953_, data_stage_4__3952_, data_stage_4__3951_, data_stage_4__3950_, data_stage_4__3949_, data_stage_4__3948_, data_stage_4__3947_, data_stage_4__3946_, data_stage_4__3945_, data_stage_4__3944_, data_stage_4__3943_, data_stage_4__3942_, data_stage_4__3941_, data_stage_4__3940_, data_stage_4__3939_, data_stage_4__3938_, data_stage_4__3937_, data_stage_4__3936_, data_stage_4__3935_, data_stage_4__3934_, data_stage_4__3933_, data_stage_4__3932_, data_stage_4__3931_, data_stage_4__3930_, data_stage_4__3929_, data_stage_4__3928_, data_stage_4__3927_, data_stage_4__3926_, data_stage_4__3925_, data_stage_4__3924_, data_stage_4__3923_, data_stage_4__3922_, data_stage_4__3921_, data_stage_4__3920_, data_stage_4__3919_, data_stage_4__3918_, data_stage_4__3917_, data_stage_4__3916_, data_stage_4__3915_, data_stage_4__3914_, data_stage_4__3913_, data_stage_4__3912_, data_stage_4__3911_, data_stage_4__3910_, data_stage_4__3909_, data_stage_4__3908_, data_stage_4__3907_, data_stage_4__3906_, data_stage_4__3905_, data_stage_4__3904_, data_stage_4__3903_, data_stage_4__3902_, data_stage_4__3901_, data_stage_4__3900_, data_stage_4__3899_, data_stage_4__3898_, data_stage_4__3897_, data_stage_4__3896_, data_stage_4__3895_, data_stage_4__3894_, data_stage_4__3893_, data_stage_4__3892_, data_stage_4__3891_, data_stage_4__3890_, data_stage_4__3889_, data_stage_4__3888_, data_stage_4__3887_, data_stage_4__3886_, data_stage_4__3885_, data_stage_4__3884_, data_stage_4__3883_, data_stage_4__3882_, data_stage_4__3881_, data_stage_4__3880_, data_stage_4__3879_, data_stage_4__3878_, data_stage_4__3877_, data_stage_4__3876_, data_stage_4__3875_, data_stage_4__3874_, data_stage_4__3873_, data_stage_4__3872_, data_stage_4__3871_, data_stage_4__3870_, data_stage_4__3869_, data_stage_4__3868_, data_stage_4__3867_, data_stage_4__3866_, data_stage_4__3865_, data_stage_4__3864_, data_stage_4__3863_, data_stage_4__3862_, data_stage_4__3861_, data_stage_4__3860_, data_stage_4__3859_, data_stage_4__3858_, data_stage_4__3857_, data_stage_4__3856_, data_stage_4__3855_, data_stage_4__3854_, data_stage_4__3853_, data_stage_4__3852_, data_stage_4__3851_, data_stage_4__3850_, data_stage_4__3849_, data_stage_4__3848_, data_stage_4__3847_, data_stage_4__3846_, data_stage_4__3845_, data_stage_4__3844_, data_stage_4__3843_, data_stage_4__3842_, data_stage_4__3841_, data_stage_4__3840_, data_stage_4__3839_, data_stage_4__3838_, data_stage_4__3837_, data_stage_4__3836_, data_stage_4__3835_, data_stage_4__3834_, data_stage_4__3833_, data_stage_4__3832_, data_stage_4__3831_, data_stage_4__3830_, data_stage_4__3829_, data_stage_4__3828_, data_stage_4__3827_, data_stage_4__3826_, data_stage_4__3825_, data_stage_4__3824_, data_stage_4__3823_, data_stage_4__3822_, data_stage_4__3821_, data_stage_4__3820_, data_stage_4__3819_, data_stage_4__3818_, data_stage_4__3817_, data_stage_4__3816_, data_stage_4__3815_, data_stage_4__3814_, data_stage_4__3813_, data_stage_4__3812_, data_stage_4__3811_, data_stage_4__3810_, data_stage_4__3809_, data_stage_4__3808_, data_stage_4__3807_, data_stage_4__3806_, data_stage_4__3805_, data_stage_4__3804_, data_stage_4__3803_, data_stage_4__3802_, data_stage_4__3801_, data_stage_4__3800_, data_stage_4__3799_, data_stage_4__3798_, data_stage_4__3797_, data_stage_4__3796_, data_stage_4__3795_, data_stage_4__3794_, data_stage_4__3793_, data_stage_4__3792_, data_stage_4__3791_, data_stage_4__3790_, data_stage_4__3789_, data_stage_4__3788_, data_stage_4__3787_, data_stage_4__3786_, data_stage_4__3785_, data_stage_4__3784_, data_stage_4__3783_, data_stage_4__3782_, data_stage_4__3781_, data_stage_4__3780_, data_stage_4__3779_, data_stage_4__3778_, data_stage_4__3777_, data_stage_4__3776_, data_stage_4__3775_, data_stage_4__3774_, data_stage_4__3773_, data_stage_4__3772_, data_stage_4__3771_, data_stage_4__3770_, data_stage_4__3769_, data_stage_4__3768_, data_stage_4__3767_, data_stage_4__3766_, data_stage_4__3765_, data_stage_4__3764_, data_stage_4__3763_, data_stage_4__3762_, data_stage_4__3761_, data_stage_4__3760_, data_stage_4__3759_, data_stage_4__3758_, data_stage_4__3757_, data_stage_4__3756_, data_stage_4__3755_, data_stage_4__3754_, data_stage_4__3753_, data_stage_4__3752_, data_stage_4__3751_, data_stage_4__3750_, data_stage_4__3749_, data_stage_4__3748_, data_stage_4__3747_, data_stage_4__3746_, data_stage_4__3745_, data_stage_4__3744_, data_stage_4__3743_, data_stage_4__3742_, data_stage_4__3741_, data_stage_4__3740_, data_stage_4__3739_, data_stage_4__3738_, data_stage_4__3737_, data_stage_4__3736_, data_stage_4__3735_, data_stage_4__3734_, data_stage_4__3733_, data_stage_4__3732_, data_stage_4__3731_, data_stage_4__3730_, data_stage_4__3729_, data_stage_4__3728_, data_stage_4__3727_, data_stage_4__3726_, data_stage_4__3725_, data_stage_4__3724_, data_stage_4__3723_, data_stage_4__3722_, data_stage_4__3721_, data_stage_4__3720_, data_stage_4__3719_, data_stage_4__3718_, data_stage_4__3717_, data_stage_4__3716_, data_stage_4__3715_, data_stage_4__3714_, data_stage_4__3713_, data_stage_4__3712_, data_stage_4__3711_, data_stage_4__3710_, data_stage_4__3709_, data_stage_4__3708_, data_stage_4__3707_, data_stage_4__3706_, data_stage_4__3705_, data_stage_4__3704_, data_stage_4__3703_, data_stage_4__3702_, data_stage_4__3701_, data_stage_4__3700_, data_stage_4__3699_, data_stage_4__3698_, data_stage_4__3697_, data_stage_4__3696_, data_stage_4__3695_, data_stage_4__3694_, data_stage_4__3693_, data_stage_4__3692_, data_stage_4__3691_, data_stage_4__3690_, data_stage_4__3689_, data_stage_4__3688_, data_stage_4__3687_, data_stage_4__3686_, data_stage_4__3685_, data_stage_4__3684_, data_stage_4__3683_, data_stage_4__3682_, data_stage_4__3681_, data_stage_4__3680_, data_stage_4__3679_, data_stage_4__3678_, data_stage_4__3677_, data_stage_4__3676_, data_stage_4__3675_, data_stage_4__3674_, data_stage_4__3673_, data_stage_4__3672_, data_stage_4__3671_, data_stage_4__3670_, data_stage_4__3669_, data_stage_4__3668_, data_stage_4__3667_, data_stage_4__3666_, data_stage_4__3665_, data_stage_4__3664_, data_stage_4__3663_, data_stage_4__3662_, data_stage_4__3661_, data_stage_4__3660_, data_stage_4__3659_, data_stage_4__3658_, data_stage_4__3657_, data_stage_4__3656_, data_stage_4__3655_, data_stage_4__3654_, data_stage_4__3653_, data_stage_4__3652_, data_stage_4__3651_, data_stage_4__3650_, data_stage_4__3649_, data_stage_4__3648_, data_stage_4__3647_, data_stage_4__3646_, data_stage_4__3645_, data_stage_4__3644_, data_stage_4__3643_, data_stage_4__3642_, data_stage_4__3641_, data_stage_4__3640_, data_stage_4__3639_, data_stage_4__3638_, data_stage_4__3637_, data_stage_4__3636_, data_stage_4__3635_, data_stage_4__3634_, data_stage_4__3633_, data_stage_4__3632_, data_stage_4__3631_, data_stage_4__3630_, data_stage_4__3629_, data_stage_4__3628_, data_stage_4__3627_, data_stage_4__3626_, data_stage_4__3625_, data_stage_4__3624_, data_stage_4__3623_, data_stage_4__3622_, data_stage_4__3621_, data_stage_4__3620_, data_stage_4__3619_, data_stage_4__3618_, data_stage_4__3617_, data_stage_4__3616_, data_stage_4__3615_, data_stage_4__3614_, data_stage_4__3613_, data_stage_4__3612_, data_stage_4__3611_, data_stage_4__3610_, data_stage_4__3609_, data_stage_4__3608_, data_stage_4__3607_, data_stage_4__3606_, data_stage_4__3605_, data_stage_4__3604_, data_stage_4__3603_, data_stage_4__3602_, data_stage_4__3601_, data_stage_4__3600_, data_stage_4__3599_, data_stage_4__3598_, data_stage_4__3597_, data_stage_4__3596_, data_stage_4__3595_, data_stage_4__3594_, data_stage_4__3593_, data_stage_4__3592_, data_stage_4__3591_, data_stage_4__3590_, data_stage_4__3589_, data_stage_4__3588_, data_stage_4__3587_, data_stage_4__3586_, data_stage_4__3585_, data_stage_4__3584_, data_stage_4__3583_, data_stage_4__3582_, data_stage_4__3581_, data_stage_4__3580_, data_stage_4__3579_, data_stage_4__3578_, data_stage_4__3577_, data_stage_4__3576_, data_stage_4__3575_, data_stage_4__3574_, data_stage_4__3573_, data_stage_4__3572_, data_stage_4__3571_, data_stage_4__3570_, data_stage_4__3569_, data_stage_4__3568_, data_stage_4__3567_, data_stage_4__3566_, data_stage_4__3565_, data_stage_4__3564_, data_stage_4__3563_, data_stage_4__3562_, data_stage_4__3561_, data_stage_4__3560_, data_stage_4__3559_, data_stage_4__3558_, data_stage_4__3557_, data_stage_4__3556_, data_stage_4__3555_, data_stage_4__3554_, data_stage_4__3553_, data_stage_4__3552_, data_stage_4__3551_, data_stage_4__3550_, data_stage_4__3549_, data_stage_4__3548_, data_stage_4__3547_, data_stage_4__3546_, data_stage_4__3545_, data_stage_4__3544_, data_stage_4__3543_, data_stage_4__3542_, data_stage_4__3541_, data_stage_4__3540_, data_stage_4__3539_, data_stage_4__3538_, data_stage_4__3537_, data_stage_4__3536_, data_stage_4__3535_, data_stage_4__3534_, data_stage_4__3533_, data_stage_4__3532_, data_stage_4__3531_, data_stage_4__3530_, data_stage_4__3529_, data_stage_4__3528_, data_stage_4__3527_, data_stage_4__3526_, data_stage_4__3525_, data_stage_4__3524_, data_stage_4__3523_, data_stage_4__3522_, data_stage_4__3521_, data_stage_4__3520_, data_stage_4__3519_, data_stage_4__3518_, data_stage_4__3517_, data_stage_4__3516_, data_stage_4__3515_, data_stage_4__3514_, data_stage_4__3513_, data_stage_4__3512_, data_stage_4__3511_, data_stage_4__3510_, data_stage_4__3509_, data_stage_4__3508_, data_stage_4__3507_, data_stage_4__3506_, data_stage_4__3505_, data_stage_4__3504_, data_stage_4__3503_, data_stage_4__3502_, data_stage_4__3501_, data_stage_4__3500_, data_stage_4__3499_, data_stage_4__3498_, data_stage_4__3497_, data_stage_4__3496_, data_stage_4__3495_, data_stage_4__3494_, data_stage_4__3493_, data_stage_4__3492_, data_stage_4__3491_, data_stage_4__3490_, data_stage_4__3489_, data_stage_4__3488_, data_stage_4__3487_, data_stage_4__3486_, data_stage_4__3485_, data_stage_4__3484_, data_stage_4__3483_, data_stage_4__3482_, data_stage_4__3481_, data_stage_4__3480_, data_stage_4__3479_, data_stage_4__3478_, data_stage_4__3477_, data_stage_4__3476_, data_stage_4__3475_, data_stage_4__3474_, data_stage_4__3473_, data_stage_4__3472_, data_stage_4__3471_, data_stage_4__3470_, data_stage_4__3469_, data_stage_4__3468_, data_stage_4__3467_, data_stage_4__3466_, data_stage_4__3465_, data_stage_4__3464_, data_stage_4__3463_, data_stage_4__3462_, data_stage_4__3461_, data_stage_4__3460_, data_stage_4__3459_, data_stage_4__3458_, data_stage_4__3457_, data_stage_4__3456_, data_stage_4__3455_, data_stage_4__3454_, data_stage_4__3453_, data_stage_4__3452_, data_stage_4__3451_, data_stage_4__3450_, data_stage_4__3449_, data_stage_4__3448_, data_stage_4__3447_, data_stage_4__3446_, data_stage_4__3445_, data_stage_4__3444_, data_stage_4__3443_, data_stage_4__3442_, data_stage_4__3441_, data_stage_4__3440_, data_stage_4__3439_, data_stage_4__3438_, data_stage_4__3437_, data_stage_4__3436_, data_stage_4__3435_, data_stage_4__3434_, data_stage_4__3433_, data_stage_4__3432_, data_stage_4__3431_, data_stage_4__3430_, data_stage_4__3429_, data_stage_4__3428_, data_stage_4__3427_, data_stage_4__3426_, data_stage_4__3425_, data_stage_4__3424_, data_stage_4__3423_, data_stage_4__3422_, data_stage_4__3421_, data_stage_4__3420_, data_stage_4__3419_, data_stage_4__3418_, data_stage_4__3417_, data_stage_4__3416_, data_stage_4__3415_, data_stage_4__3414_, data_stage_4__3413_, data_stage_4__3412_, data_stage_4__3411_, data_stage_4__3410_, data_stage_4__3409_, data_stage_4__3408_, data_stage_4__3407_, data_stage_4__3406_, data_stage_4__3405_, data_stage_4__3404_, data_stage_4__3403_, data_stage_4__3402_, data_stage_4__3401_, data_stage_4__3400_, data_stage_4__3399_, data_stage_4__3398_, data_stage_4__3397_, data_stage_4__3396_, data_stage_4__3395_, data_stage_4__3394_, data_stage_4__3393_, data_stage_4__3392_, data_stage_4__3391_, data_stage_4__3390_, data_stage_4__3389_, data_stage_4__3388_, data_stage_4__3387_, data_stage_4__3386_, data_stage_4__3385_, data_stage_4__3384_, data_stage_4__3383_, data_stage_4__3382_, data_stage_4__3381_, data_stage_4__3380_, data_stage_4__3379_, data_stage_4__3378_, data_stage_4__3377_, data_stage_4__3376_, data_stage_4__3375_, data_stage_4__3374_, data_stage_4__3373_, data_stage_4__3372_, data_stage_4__3371_, data_stage_4__3370_, data_stage_4__3369_, data_stage_4__3368_, data_stage_4__3367_, data_stage_4__3366_, data_stage_4__3365_, data_stage_4__3364_, data_stage_4__3363_, data_stage_4__3362_, data_stage_4__3361_, data_stage_4__3360_, data_stage_4__3359_, data_stage_4__3358_, data_stage_4__3357_, data_stage_4__3356_, data_stage_4__3355_, data_stage_4__3354_, data_stage_4__3353_, data_stage_4__3352_, data_stage_4__3351_, data_stage_4__3350_, data_stage_4__3349_, data_stage_4__3348_, data_stage_4__3347_, data_stage_4__3346_, data_stage_4__3345_, data_stage_4__3344_, data_stage_4__3343_, data_stage_4__3342_, data_stage_4__3341_, data_stage_4__3340_, data_stage_4__3339_, data_stage_4__3338_, data_stage_4__3337_, data_stage_4__3336_, data_stage_4__3335_, data_stage_4__3334_, data_stage_4__3333_, data_stage_4__3332_, data_stage_4__3331_, data_stage_4__3330_, data_stage_4__3329_, data_stage_4__3328_, data_stage_4__3327_, data_stage_4__3326_, data_stage_4__3325_, data_stage_4__3324_, data_stage_4__3323_, data_stage_4__3322_, data_stage_4__3321_, data_stage_4__3320_, data_stage_4__3319_, data_stage_4__3318_, data_stage_4__3317_, data_stage_4__3316_, data_stage_4__3315_, data_stage_4__3314_, data_stage_4__3313_, data_stage_4__3312_, data_stage_4__3311_, data_stage_4__3310_, data_stage_4__3309_, data_stage_4__3308_, data_stage_4__3307_, data_stage_4__3306_, data_stage_4__3305_, data_stage_4__3304_, data_stage_4__3303_, data_stage_4__3302_, data_stage_4__3301_, data_stage_4__3300_, data_stage_4__3299_, data_stage_4__3298_, data_stage_4__3297_, data_stage_4__3296_, data_stage_4__3295_, data_stage_4__3294_, data_stage_4__3293_, data_stage_4__3292_, data_stage_4__3291_, data_stage_4__3290_, data_stage_4__3289_, data_stage_4__3288_, data_stage_4__3287_, data_stage_4__3286_, data_stage_4__3285_, data_stage_4__3284_, data_stage_4__3283_, data_stage_4__3282_, data_stage_4__3281_, data_stage_4__3280_, data_stage_4__3279_, data_stage_4__3278_, data_stage_4__3277_, data_stage_4__3276_, data_stage_4__3275_, data_stage_4__3274_, data_stage_4__3273_, data_stage_4__3272_, data_stage_4__3271_, data_stage_4__3270_, data_stage_4__3269_, data_stage_4__3268_, data_stage_4__3267_, data_stage_4__3266_, data_stage_4__3265_, data_stage_4__3264_, data_stage_4__3263_, data_stage_4__3262_, data_stage_4__3261_, data_stage_4__3260_, data_stage_4__3259_, data_stage_4__3258_, data_stage_4__3257_, data_stage_4__3256_, data_stage_4__3255_, data_stage_4__3254_, data_stage_4__3253_, data_stage_4__3252_, data_stage_4__3251_, data_stage_4__3250_, data_stage_4__3249_, data_stage_4__3248_, data_stage_4__3247_, data_stage_4__3246_, data_stage_4__3245_, data_stage_4__3244_, data_stage_4__3243_, data_stage_4__3242_, data_stage_4__3241_, data_stage_4__3240_, data_stage_4__3239_, data_stage_4__3238_, data_stage_4__3237_, data_stage_4__3236_, data_stage_4__3235_, data_stage_4__3234_, data_stage_4__3233_, data_stage_4__3232_, data_stage_4__3231_, data_stage_4__3230_, data_stage_4__3229_, data_stage_4__3228_, data_stage_4__3227_, data_stage_4__3226_, data_stage_4__3225_, data_stage_4__3224_, data_stage_4__3223_, data_stage_4__3222_, data_stage_4__3221_, data_stage_4__3220_, data_stage_4__3219_, data_stage_4__3218_, data_stage_4__3217_, data_stage_4__3216_, data_stage_4__3215_, data_stage_4__3214_, data_stage_4__3213_, data_stage_4__3212_, data_stage_4__3211_, data_stage_4__3210_, data_stage_4__3209_, data_stage_4__3208_, data_stage_4__3207_, data_stage_4__3206_, data_stage_4__3205_, data_stage_4__3204_, data_stage_4__3203_, data_stage_4__3202_, data_stage_4__3201_, data_stage_4__3200_, data_stage_4__3199_, data_stage_4__3198_, data_stage_4__3197_, data_stage_4__3196_, data_stage_4__3195_, data_stage_4__3194_, data_stage_4__3193_, data_stage_4__3192_, data_stage_4__3191_, data_stage_4__3190_, data_stage_4__3189_, data_stage_4__3188_, data_stage_4__3187_, data_stage_4__3186_, data_stage_4__3185_, data_stage_4__3184_, data_stage_4__3183_, data_stage_4__3182_, data_stage_4__3181_, data_stage_4__3180_, data_stage_4__3179_, data_stage_4__3178_, data_stage_4__3177_, data_stage_4__3176_, data_stage_4__3175_, data_stage_4__3174_, data_stage_4__3173_, data_stage_4__3172_, data_stage_4__3171_, data_stage_4__3170_, data_stage_4__3169_, data_stage_4__3168_, data_stage_4__3167_, data_stage_4__3166_, data_stage_4__3165_, data_stage_4__3164_, data_stage_4__3163_, data_stage_4__3162_, data_stage_4__3161_, data_stage_4__3160_, data_stage_4__3159_, data_stage_4__3158_, data_stage_4__3157_, data_stage_4__3156_, data_stage_4__3155_, data_stage_4__3154_, data_stage_4__3153_, data_stage_4__3152_, data_stage_4__3151_, data_stage_4__3150_, data_stage_4__3149_, data_stage_4__3148_, data_stage_4__3147_, data_stage_4__3146_, data_stage_4__3145_, data_stage_4__3144_, data_stage_4__3143_, data_stage_4__3142_, data_stage_4__3141_, data_stage_4__3140_, data_stage_4__3139_, data_stage_4__3138_, data_stage_4__3137_, data_stage_4__3136_, data_stage_4__3135_, data_stage_4__3134_, data_stage_4__3133_, data_stage_4__3132_, data_stage_4__3131_, data_stage_4__3130_, data_stage_4__3129_, data_stage_4__3128_, data_stage_4__3127_, data_stage_4__3126_, data_stage_4__3125_, data_stage_4__3124_, data_stage_4__3123_, data_stage_4__3122_, data_stage_4__3121_, data_stage_4__3120_, data_stage_4__3119_, data_stage_4__3118_, data_stage_4__3117_, data_stage_4__3116_, data_stage_4__3115_, data_stage_4__3114_, data_stage_4__3113_, data_stage_4__3112_, data_stage_4__3111_, data_stage_4__3110_, data_stage_4__3109_, data_stage_4__3108_, data_stage_4__3107_, data_stage_4__3106_, data_stage_4__3105_, data_stage_4__3104_, data_stage_4__3103_, data_stage_4__3102_, data_stage_4__3101_, data_stage_4__3100_, data_stage_4__3099_, data_stage_4__3098_, data_stage_4__3097_, data_stage_4__3096_, data_stage_4__3095_, data_stage_4__3094_, data_stage_4__3093_, data_stage_4__3092_, data_stage_4__3091_, data_stage_4__3090_, data_stage_4__3089_, data_stage_4__3088_, data_stage_4__3087_, data_stage_4__3086_, data_stage_4__3085_, data_stage_4__3084_, data_stage_4__3083_, data_stage_4__3082_, data_stage_4__3081_, data_stage_4__3080_, data_stage_4__3079_, data_stage_4__3078_, data_stage_4__3077_, data_stage_4__3076_, data_stage_4__3075_, data_stage_4__3074_, data_stage_4__3073_, data_stage_4__3072_, data_stage_4__3071_, data_stage_4__3070_, data_stage_4__3069_, data_stage_4__3068_, data_stage_4__3067_, data_stage_4__3066_, data_stage_4__3065_, data_stage_4__3064_, data_stage_4__3063_, data_stage_4__3062_, data_stage_4__3061_, data_stage_4__3060_, data_stage_4__3059_, data_stage_4__3058_, data_stage_4__3057_, data_stage_4__3056_, data_stage_4__3055_, data_stage_4__3054_, data_stage_4__3053_, data_stage_4__3052_, data_stage_4__3051_, data_stage_4__3050_, data_stage_4__3049_, data_stage_4__3048_, data_stage_4__3047_, data_stage_4__3046_, data_stage_4__3045_, data_stage_4__3044_, data_stage_4__3043_, data_stage_4__3042_, data_stage_4__3041_, data_stage_4__3040_, data_stage_4__3039_, data_stage_4__3038_, data_stage_4__3037_, data_stage_4__3036_, data_stage_4__3035_, data_stage_4__3034_, data_stage_4__3033_, data_stage_4__3032_, data_stage_4__3031_, data_stage_4__3030_, data_stage_4__3029_, data_stage_4__3028_, data_stage_4__3027_, data_stage_4__3026_, data_stage_4__3025_, data_stage_4__3024_, data_stage_4__3023_, data_stage_4__3022_, data_stage_4__3021_, data_stage_4__3020_, data_stage_4__3019_, data_stage_4__3018_, data_stage_4__3017_, data_stage_4__3016_, data_stage_4__3015_, data_stage_4__3014_, data_stage_4__3013_, data_stage_4__3012_, data_stage_4__3011_, data_stage_4__3010_, data_stage_4__3009_, data_stage_4__3008_, data_stage_4__3007_, data_stage_4__3006_, data_stage_4__3005_, data_stage_4__3004_, data_stage_4__3003_, data_stage_4__3002_, data_stage_4__3001_, data_stage_4__3000_, data_stage_4__2999_, data_stage_4__2998_, data_stage_4__2997_, data_stage_4__2996_, data_stage_4__2995_, data_stage_4__2994_, data_stage_4__2993_, data_stage_4__2992_, data_stage_4__2991_, data_stage_4__2990_, data_stage_4__2989_, data_stage_4__2988_, data_stage_4__2987_, data_stage_4__2986_, data_stage_4__2985_, data_stage_4__2984_, data_stage_4__2983_, data_stage_4__2982_, data_stage_4__2981_, data_stage_4__2980_, data_stage_4__2979_, data_stage_4__2978_, data_stage_4__2977_, data_stage_4__2976_, data_stage_4__2975_, data_stage_4__2974_, data_stage_4__2973_, data_stage_4__2972_, data_stage_4__2971_, data_stage_4__2970_, data_stage_4__2969_, data_stage_4__2968_, data_stage_4__2967_, data_stage_4__2966_, data_stage_4__2965_, data_stage_4__2964_, data_stage_4__2963_, data_stage_4__2962_, data_stage_4__2961_, data_stage_4__2960_, data_stage_4__2959_, data_stage_4__2958_, data_stage_4__2957_, data_stage_4__2956_, data_stage_4__2955_, data_stage_4__2954_, data_stage_4__2953_, data_stage_4__2952_, data_stage_4__2951_, data_stage_4__2950_, data_stage_4__2949_, data_stage_4__2948_, data_stage_4__2947_, data_stage_4__2946_, data_stage_4__2945_, data_stage_4__2944_, data_stage_4__2943_, data_stage_4__2942_, data_stage_4__2941_, data_stage_4__2940_, data_stage_4__2939_, data_stage_4__2938_, data_stage_4__2937_, data_stage_4__2936_, data_stage_4__2935_, data_stage_4__2934_, data_stage_4__2933_, data_stage_4__2932_, data_stage_4__2931_, data_stage_4__2930_, data_stage_4__2929_, data_stage_4__2928_, data_stage_4__2927_, data_stage_4__2926_, data_stage_4__2925_, data_stage_4__2924_, data_stage_4__2923_, data_stage_4__2922_, data_stage_4__2921_, data_stage_4__2920_, data_stage_4__2919_, data_stage_4__2918_, data_stage_4__2917_, data_stage_4__2916_, data_stage_4__2915_, data_stage_4__2914_, data_stage_4__2913_, data_stage_4__2912_, data_stage_4__2911_, data_stage_4__2910_, data_stage_4__2909_, data_stage_4__2908_, data_stage_4__2907_, data_stage_4__2906_, data_stage_4__2905_, data_stage_4__2904_, data_stage_4__2903_, data_stage_4__2902_, data_stage_4__2901_, data_stage_4__2900_, data_stage_4__2899_, data_stage_4__2898_, data_stage_4__2897_, data_stage_4__2896_, data_stage_4__2895_, data_stage_4__2894_, data_stage_4__2893_, data_stage_4__2892_, data_stage_4__2891_, data_stage_4__2890_, data_stage_4__2889_, data_stage_4__2888_, data_stage_4__2887_, data_stage_4__2886_, data_stage_4__2885_, data_stage_4__2884_, data_stage_4__2883_, data_stage_4__2882_, data_stage_4__2881_, data_stage_4__2880_, data_stage_4__2879_, data_stage_4__2878_, data_stage_4__2877_, data_stage_4__2876_, data_stage_4__2875_, data_stage_4__2874_, data_stage_4__2873_, data_stage_4__2872_, data_stage_4__2871_, data_stage_4__2870_, data_stage_4__2869_, data_stage_4__2868_, data_stage_4__2867_, data_stage_4__2866_, data_stage_4__2865_, data_stage_4__2864_, data_stage_4__2863_, data_stage_4__2862_, data_stage_4__2861_, data_stage_4__2860_, data_stage_4__2859_, data_stage_4__2858_, data_stage_4__2857_, data_stage_4__2856_, data_stage_4__2855_, data_stage_4__2854_, data_stage_4__2853_, data_stage_4__2852_, data_stage_4__2851_, data_stage_4__2850_, data_stage_4__2849_, data_stage_4__2848_, data_stage_4__2847_, data_stage_4__2846_, data_stage_4__2845_, data_stage_4__2844_, data_stage_4__2843_, data_stage_4__2842_, data_stage_4__2841_, data_stage_4__2840_, data_stage_4__2839_, data_stage_4__2838_, data_stage_4__2837_, data_stage_4__2836_, data_stage_4__2835_, data_stage_4__2834_, data_stage_4__2833_, data_stage_4__2832_, data_stage_4__2831_, data_stage_4__2830_, data_stage_4__2829_, data_stage_4__2828_, data_stage_4__2827_, data_stage_4__2826_, data_stage_4__2825_, data_stage_4__2824_, data_stage_4__2823_, data_stage_4__2822_, data_stage_4__2821_, data_stage_4__2820_, data_stage_4__2819_, data_stage_4__2818_, data_stage_4__2817_, data_stage_4__2816_, data_stage_4__2815_, data_stage_4__2814_, data_stage_4__2813_, data_stage_4__2812_, data_stage_4__2811_, data_stage_4__2810_, data_stage_4__2809_, data_stage_4__2808_, data_stage_4__2807_, data_stage_4__2806_, data_stage_4__2805_, data_stage_4__2804_, data_stage_4__2803_, data_stage_4__2802_, data_stage_4__2801_, data_stage_4__2800_, data_stage_4__2799_, data_stage_4__2798_, data_stage_4__2797_, data_stage_4__2796_, data_stage_4__2795_, data_stage_4__2794_, data_stage_4__2793_, data_stage_4__2792_, data_stage_4__2791_, data_stage_4__2790_, data_stage_4__2789_, data_stage_4__2788_, data_stage_4__2787_, data_stage_4__2786_, data_stage_4__2785_, data_stage_4__2784_, data_stage_4__2783_, data_stage_4__2782_, data_stage_4__2781_, data_stage_4__2780_, data_stage_4__2779_, data_stage_4__2778_, data_stage_4__2777_, data_stage_4__2776_, data_stage_4__2775_, data_stage_4__2774_, data_stage_4__2773_, data_stage_4__2772_, data_stage_4__2771_, data_stage_4__2770_, data_stage_4__2769_, data_stage_4__2768_, data_stage_4__2767_, data_stage_4__2766_, data_stage_4__2765_, data_stage_4__2764_, data_stage_4__2763_, data_stage_4__2762_, data_stage_4__2761_, data_stage_4__2760_, data_stage_4__2759_, data_stage_4__2758_, data_stage_4__2757_, data_stage_4__2756_, data_stage_4__2755_, data_stage_4__2754_, data_stage_4__2753_, data_stage_4__2752_, data_stage_4__2751_, data_stage_4__2750_, data_stage_4__2749_, data_stage_4__2748_, data_stage_4__2747_, data_stage_4__2746_, data_stage_4__2745_, data_stage_4__2744_, data_stage_4__2743_, data_stage_4__2742_, data_stage_4__2741_, data_stage_4__2740_, data_stage_4__2739_, data_stage_4__2738_, data_stage_4__2737_, data_stage_4__2736_, data_stage_4__2735_, data_stage_4__2734_, data_stage_4__2733_, data_stage_4__2732_, data_stage_4__2731_, data_stage_4__2730_, data_stage_4__2729_, data_stage_4__2728_, data_stage_4__2727_, data_stage_4__2726_, data_stage_4__2725_, data_stage_4__2724_, data_stage_4__2723_, data_stage_4__2722_, data_stage_4__2721_, data_stage_4__2720_, data_stage_4__2719_, data_stage_4__2718_, data_stage_4__2717_, data_stage_4__2716_, data_stage_4__2715_, data_stage_4__2714_, data_stage_4__2713_, data_stage_4__2712_, data_stage_4__2711_, data_stage_4__2710_, data_stage_4__2709_, data_stage_4__2708_, data_stage_4__2707_, data_stage_4__2706_, data_stage_4__2705_, data_stage_4__2704_, data_stage_4__2703_, data_stage_4__2702_, data_stage_4__2701_, data_stage_4__2700_, data_stage_4__2699_, data_stage_4__2698_, data_stage_4__2697_, data_stage_4__2696_, data_stage_4__2695_, data_stage_4__2694_, data_stage_4__2693_, data_stage_4__2692_, data_stage_4__2691_, data_stage_4__2690_, data_stage_4__2689_, data_stage_4__2688_, data_stage_4__2687_, data_stage_4__2686_, data_stage_4__2685_, data_stage_4__2684_, data_stage_4__2683_, data_stage_4__2682_, data_stage_4__2681_, data_stage_4__2680_, data_stage_4__2679_, data_stage_4__2678_, data_stage_4__2677_, data_stage_4__2676_, data_stage_4__2675_, data_stage_4__2674_, data_stage_4__2673_, data_stage_4__2672_, data_stage_4__2671_, data_stage_4__2670_, data_stage_4__2669_, data_stage_4__2668_, data_stage_4__2667_, data_stage_4__2666_, data_stage_4__2665_, data_stage_4__2664_, data_stage_4__2663_, data_stage_4__2662_, data_stage_4__2661_, data_stage_4__2660_, data_stage_4__2659_, data_stage_4__2658_, data_stage_4__2657_, data_stage_4__2656_, data_stage_4__2655_, data_stage_4__2654_, data_stage_4__2653_, data_stage_4__2652_, data_stage_4__2651_, data_stage_4__2650_, data_stage_4__2649_, data_stage_4__2648_, data_stage_4__2647_, data_stage_4__2646_, data_stage_4__2645_, data_stage_4__2644_, data_stage_4__2643_, data_stage_4__2642_, data_stage_4__2641_, data_stage_4__2640_, data_stage_4__2639_, data_stage_4__2638_, data_stage_4__2637_, data_stage_4__2636_, data_stage_4__2635_, data_stage_4__2634_, data_stage_4__2633_, data_stage_4__2632_, data_stage_4__2631_, data_stage_4__2630_, data_stage_4__2629_, data_stage_4__2628_, data_stage_4__2627_, data_stage_4__2626_, data_stage_4__2625_, data_stage_4__2624_, data_stage_4__2623_, data_stage_4__2622_, data_stage_4__2621_, data_stage_4__2620_, data_stage_4__2619_, data_stage_4__2618_, data_stage_4__2617_, data_stage_4__2616_, data_stage_4__2615_, data_stage_4__2614_, data_stage_4__2613_, data_stage_4__2612_, data_stage_4__2611_, data_stage_4__2610_, data_stage_4__2609_, data_stage_4__2608_, data_stage_4__2607_, data_stage_4__2606_, data_stage_4__2605_, data_stage_4__2604_, data_stage_4__2603_, data_stage_4__2602_, data_stage_4__2601_, data_stage_4__2600_, data_stage_4__2599_, data_stage_4__2598_, data_stage_4__2597_, data_stage_4__2596_, data_stage_4__2595_, data_stage_4__2594_, data_stage_4__2593_, data_stage_4__2592_, data_stage_4__2591_, data_stage_4__2590_, data_stage_4__2589_, data_stage_4__2588_, data_stage_4__2587_, data_stage_4__2586_, data_stage_4__2585_, data_stage_4__2584_, data_stage_4__2583_, data_stage_4__2582_, data_stage_4__2581_, data_stage_4__2580_, data_stage_4__2579_, data_stage_4__2578_, data_stage_4__2577_, data_stage_4__2576_, data_stage_4__2575_, data_stage_4__2574_, data_stage_4__2573_, data_stage_4__2572_, data_stage_4__2571_, data_stage_4__2570_, data_stage_4__2569_, data_stage_4__2568_, data_stage_4__2567_, data_stage_4__2566_, data_stage_4__2565_, data_stage_4__2564_, data_stage_4__2563_, data_stage_4__2562_, data_stage_4__2561_, data_stage_4__2560_, data_stage_4__2559_, data_stage_4__2558_, data_stage_4__2557_, data_stage_4__2556_, data_stage_4__2555_, data_stage_4__2554_, data_stage_4__2553_, data_stage_4__2552_, data_stage_4__2551_, data_stage_4__2550_, data_stage_4__2549_, data_stage_4__2548_, data_stage_4__2547_, data_stage_4__2546_, data_stage_4__2545_, data_stage_4__2544_, data_stage_4__2543_, data_stage_4__2542_, data_stage_4__2541_, data_stage_4__2540_, data_stage_4__2539_, data_stage_4__2538_, data_stage_4__2537_, data_stage_4__2536_, data_stage_4__2535_, data_stage_4__2534_, data_stage_4__2533_, data_stage_4__2532_, data_stage_4__2531_, data_stage_4__2530_, data_stage_4__2529_, data_stage_4__2528_, data_stage_4__2527_, data_stage_4__2526_, data_stage_4__2525_, data_stage_4__2524_, data_stage_4__2523_, data_stage_4__2522_, data_stage_4__2521_, data_stage_4__2520_, data_stage_4__2519_, data_stage_4__2518_, data_stage_4__2517_, data_stage_4__2516_, data_stage_4__2515_, data_stage_4__2514_, data_stage_4__2513_, data_stage_4__2512_, data_stage_4__2511_, data_stage_4__2510_, data_stage_4__2509_, data_stage_4__2508_, data_stage_4__2507_, data_stage_4__2506_, data_stage_4__2505_, data_stage_4__2504_, data_stage_4__2503_, data_stage_4__2502_, data_stage_4__2501_, data_stage_4__2500_, data_stage_4__2499_, data_stage_4__2498_, data_stage_4__2497_, data_stage_4__2496_, data_stage_4__2495_, data_stage_4__2494_, data_stage_4__2493_, data_stage_4__2492_, data_stage_4__2491_, data_stage_4__2490_, data_stage_4__2489_, data_stage_4__2488_, data_stage_4__2487_, data_stage_4__2486_, data_stage_4__2485_, data_stage_4__2484_, data_stage_4__2483_, data_stage_4__2482_, data_stage_4__2481_, data_stage_4__2480_, data_stage_4__2479_, data_stage_4__2478_, data_stage_4__2477_, data_stage_4__2476_, data_stage_4__2475_, data_stage_4__2474_, data_stage_4__2473_, data_stage_4__2472_, data_stage_4__2471_, data_stage_4__2470_, data_stage_4__2469_, data_stage_4__2468_, data_stage_4__2467_, data_stage_4__2466_, data_stage_4__2465_, data_stage_4__2464_, data_stage_4__2463_, data_stage_4__2462_, data_stage_4__2461_, data_stage_4__2460_, data_stage_4__2459_, data_stage_4__2458_, data_stage_4__2457_, data_stage_4__2456_, data_stage_4__2455_, data_stage_4__2454_, data_stage_4__2453_, data_stage_4__2452_, data_stage_4__2451_, data_stage_4__2450_, data_stage_4__2449_, data_stage_4__2448_, data_stage_4__2447_, data_stage_4__2446_, data_stage_4__2445_, data_stage_4__2444_, data_stage_4__2443_, data_stage_4__2442_, data_stage_4__2441_, data_stage_4__2440_, data_stage_4__2439_, data_stage_4__2438_, data_stage_4__2437_, data_stage_4__2436_, data_stage_4__2435_, data_stage_4__2434_, data_stage_4__2433_, data_stage_4__2432_, data_stage_4__2431_, data_stage_4__2430_, data_stage_4__2429_, data_stage_4__2428_, data_stage_4__2427_, data_stage_4__2426_, data_stage_4__2425_, data_stage_4__2424_, data_stage_4__2423_, data_stage_4__2422_, data_stage_4__2421_, data_stage_4__2420_, data_stage_4__2419_, data_stage_4__2418_, data_stage_4__2417_, data_stage_4__2416_, data_stage_4__2415_, data_stage_4__2414_, data_stage_4__2413_, data_stage_4__2412_, data_stage_4__2411_, data_stage_4__2410_, data_stage_4__2409_, data_stage_4__2408_, data_stage_4__2407_, data_stage_4__2406_, data_stage_4__2405_, data_stage_4__2404_, data_stage_4__2403_, data_stage_4__2402_, data_stage_4__2401_, data_stage_4__2400_, data_stage_4__2399_, data_stage_4__2398_, data_stage_4__2397_, data_stage_4__2396_, data_stage_4__2395_, data_stage_4__2394_, data_stage_4__2393_, data_stage_4__2392_, data_stage_4__2391_, data_stage_4__2390_, data_stage_4__2389_, data_stage_4__2388_, data_stage_4__2387_, data_stage_4__2386_, data_stage_4__2385_, data_stage_4__2384_, data_stage_4__2383_, data_stage_4__2382_, data_stage_4__2381_, data_stage_4__2380_, data_stage_4__2379_, data_stage_4__2378_, data_stage_4__2377_, data_stage_4__2376_, data_stage_4__2375_, data_stage_4__2374_, data_stage_4__2373_, data_stage_4__2372_, data_stage_4__2371_, data_stage_4__2370_, data_stage_4__2369_, data_stage_4__2368_, data_stage_4__2367_, data_stage_4__2366_, data_stage_4__2365_, data_stage_4__2364_, data_stage_4__2363_, data_stage_4__2362_, data_stage_4__2361_, data_stage_4__2360_, data_stage_4__2359_, data_stage_4__2358_, data_stage_4__2357_, data_stage_4__2356_, data_stage_4__2355_, data_stage_4__2354_, data_stage_4__2353_, data_stage_4__2352_, data_stage_4__2351_, data_stage_4__2350_, data_stage_4__2349_, data_stage_4__2348_, data_stage_4__2347_, data_stage_4__2346_, data_stage_4__2345_, data_stage_4__2344_, data_stage_4__2343_, data_stage_4__2342_, data_stage_4__2341_, data_stage_4__2340_, data_stage_4__2339_, data_stage_4__2338_, data_stage_4__2337_, data_stage_4__2336_, data_stage_4__2335_, data_stage_4__2334_, data_stage_4__2333_, data_stage_4__2332_, data_stage_4__2331_, data_stage_4__2330_, data_stage_4__2329_, data_stage_4__2328_, data_stage_4__2327_, data_stage_4__2326_, data_stage_4__2325_, data_stage_4__2324_, data_stage_4__2323_, data_stage_4__2322_, data_stage_4__2321_, data_stage_4__2320_, data_stage_4__2319_, data_stage_4__2318_, data_stage_4__2317_, data_stage_4__2316_, data_stage_4__2315_, data_stage_4__2314_, data_stage_4__2313_, data_stage_4__2312_, data_stage_4__2311_, data_stage_4__2310_, data_stage_4__2309_, data_stage_4__2308_, data_stage_4__2307_, data_stage_4__2306_, data_stage_4__2305_, data_stage_4__2304_, data_stage_4__2303_, data_stage_4__2302_, data_stage_4__2301_, data_stage_4__2300_, data_stage_4__2299_, data_stage_4__2298_, data_stage_4__2297_, data_stage_4__2296_, data_stage_4__2295_, data_stage_4__2294_, data_stage_4__2293_, data_stage_4__2292_, data_stage_4__2291_, data_stage_4__2290_, data_stage_4__2289_, data_stage_4__2288_, data_stage_4__2287_, data_stage_4__2286_, data_stage_4__2285_, data_stage_4__2284_, data_stage_4__2283_, data_stage_4__2282_, data_stage_4__2281_, data_stage_4__2280_, data_stage_4__2279_, data_stage_4__2278_, data_stage_4__2277_, data_stage_4__2276_, data_stage_4__2275_, data_stage_4__2274_, data_stage_4__2273_, data_stage_4__2272_, data_stage_4__2271_, data_stage_4__2270_, data_stage_4__2269_, data_stage_4__2268_, data_stage_4__2267_, data_stage_4__2266_, data_stage_4__2265_, data_stage_4__2264_, data_stage_4__2263_, data_stage_4__2262_, data_stage_4__2261_, data_stage_4__2260_, data_stage_4__2259_, data_stage_4__2258_, data_stage_4__2257_, data_stage_4__2256_, data_stage_4__2255_, data_stage_4__2254_, data_stage_4__2253_, data_stage_4__2252_, data_stage_4__2251_, data_stage_4__2250_, data_stage_4__2249_, data_stage_4__2248_, data_stage_4__2247_, data_stage_4__2246_, data_stage_4__2245_, data_stage_4__2244_, data_stage_4__2243_, data_stage_4__2242_, data_stage_4__2241_, data_stage_4__2240_, data_stage_4__2239_, data_stage_4__2238_, data_stage_4__2237_, data_stage_4__2236_, data_stage_4__2235_, data_stage_4__2234_, data_stage_4__2233_, data_stage_4__2232_, data_stage_4__2231_, data_stage_4__2230_, data_stage_4__2229_, data_stage_4__2228_, data_stage_4__2227_, data_stage_4__2226_, data_stage_4__2225_, data_stage_4__2224_, data_stage_4__2223_, data_stage_4__2222_, data_stage_4__2221_, data_stage_4__2220_, data_stage_4__2219_, data_stage_4__2218_, data_stage_4__2217_, data_stage_4__2216_, data_stage_4__2215_, data_stage_4__2214_, data_stage_4__2213_, data_stage_4__2212_, data_stage_4__2211_, data_stage_4__2210_, data_stage_4__2209_, data_stage_4__2208_, data_stage_4__2207_, data_stage_4__2206_, data_stage_4__2205_, data_stage_4__2204_, data_stage_4__2203_, data_stage_4__2202_, data_stage_4__2201_, data_stage_4__2200_, data_stage_4__2199_, data_stage_4__2198_, data_stage_4__2197_, data_stage_4__2196_, data_stage_4__2195_, data_stage_4__2194_, data_stage_4__2193_, data_stage_4__2192_, data_stage_4__2191_, data_stage_4__2190_, data_stage_4__2189_, data_stage_4__2188_, data_stage_4__2187_, data_stage_4__2186_, data_stage_4__2185_, data_stage_4__2184_, data_stage_4__2183_, data_stage_4__2182_, data_stage_4__2181_, data_stage_4__2180_, data_stage_4__2179_, data_stage_4__2178_, data_stage_4__2177_, data_stage_4__2176_, data_stage_4__2175_, data_stage_4__2174_, data_stage_4__2173_, data_stage_4__2172_, data_stage_4__2171_, data_stage_4__2170_, data_stage_4__2169_, data_stage_4__2168_, data_stage_4__2167_, data_stage_4__2166_, data_stage_4__2165_, data_stage_4__2164_, data_stage_4__2163_, data_stage_4__2162_, data_stage_4__2161_, data_stage_4__2160_, data_stage_4__2159_, data_stage_4__2158_, data_stage_4__2157_, data_stage_4__2156_, data_stage_4__2155_, data_stage_4__2154_, data_stage_4__2153_, data_stage_4__2152_, data_stage_4__2151_, data_stage_4__2150_, data_stage_4__2149_, data_stage_4__2148_, data_stage_4__2147_, data_stage_4__2146_, data_stage_4__2145_, data_stage_4__2144_, data_stage_4__2143_, data_stage_4__2142_, data_stage_4__2141_, data_stage_4__2140_, data_stage_4__2139_, data_stage_4__2138_, data_stage_4__2137_, data_stage_4__2136_, data_stage_4__2135_, data_stage_4__2134_, data_stage_4__2133_, data_stage_4__2132_, data_stage_4__2131_, data_stage_4__2130_, data_stage_4__2129_, data_stage_4__2128_, data_stage_4__2127_, data_stage_4__2126_, data_stage_4__2125_, data_stage_4__2124_, data_stage_4__2123_, data_stage_4__2122_, data_stage_4__2121_, data_stage_4__2120_, data_stage_4__2119_, data_stage_4__2118_, data_stage_4__2117_, data_stage_4__2116_, data_stage_4__2115_, data_stage_4__2114_, data_stage_4__2113_, data_stage_4__2112_, data_stage_4__2111_, data_stage_4__2110_, data_stage_4__2109_, data_stage_4__2108_, data_stage_4__2107_, data_stage_4__2106_, data_stage_4__2105_, data_stage_4__2104_, data_stage_4__2103_, data_stage_4__2102_, data_stage_4__2101_, data_stage_4__2100_, data_stage_4__2099_, data_stage_4__2098_, data_stage_4__2097_, data_stage_4__2096_, data_stage_4__2095_, data_stage_4__2094_, data_stage_4__2093_, data_stage_4__2092_, data_stage_4__2091_, data_stage_4__2090_, data_stage_4__2089_, data_stage_4__2088_, data_stage_4__2087_, data_stage_4__2086_, data_stage_4__2085_, data_stage_4__2084_, data_stage_4__2083_, data_stage_4__2082_, data_stage_4__2081_, data_stage_4__2080_, data_stage_4__2079_, data_stage_4__2078_, data_stage_4__2077_, data_stage_4__2076_, data_stage_4__2075_, data_stage_4__2074_, data_stage_4__2073_, data_stage_4__2072_, data_stage_4__2071_, data_stage_4__2070_, data_stage_4__2069_, data_stage_4__2068_, data_stage_4__2067_, data_stage_4__2066_, data_stage_4__2065_, data_stage_4__2064_, data_stage_4__2063_, data_stage_4__2062_, data_stage_4__2061_, data_stage_4__2060_, data_stage_4__2059_, data_stage_4__2058_, data_stage_4__2057_, data_stage_4__2056_, data_stage_4__2055_, data_stage_4__2054_, data_stage_4__2053_, data_stage_4__2052_, data_stage_4__2051_, data_stage_4__2050_, data_stage_4__2049_, data_stage_4__2048_, data_stage_4__2047_, data_stage_4__2046_, data_stage_4__2045_, data_stage_4__2044_, data_stage_4__2043_, data_stage_4__2042_, data_stage_4__2041_, data_stage_4__2040_, data_stage_4__2039_, data_stage_4__2038_, data_stage_4__2037_, data_stage_4__2036_, data_stage_4__2035_, data_stage_4__2034_, data_stage_4__2033_, data_stage_4__2032_, data_stage_4__2031_, data_stage_4__2030_, data_stage_4__2029_, data_stage_4__2028_, data_stage_4__2027_, data_stage_4__2026_, data_stage_4__2025_, data_stage_4__2024_, data_stage_4__2023_, data_stage_4__2022_, data_stage_4__2021_, data_stage_4__2020_, data_stage_4__2019_, data_stage_4__2018_, data_stage_4__2017_, data_stage_4__2016_, data_stage_4__2015_, data_stage_4__2014_, data_stage_4__2013_, data_stage_4__2012_, data_stage_4__2011_, data_stage_4__2010_, data_stage_4__2009_, data_stage_4__2008_, data_stage_4__2007_, data_stage_4__2006_, data_stage_4__2005_, data_stage_4__2004_, data_stage_4__2003_, data_stage_4__2002_, data_stage_4__2001_, data_stage_4__2000_, data_stage_4__1999_, data_stage_4__1998_, data_stage_4__1997_, data_stage_4__1996_, data_stage_4__1995_, data_stage_4__1994_, data_stage_4__1993_, data_stage_4__1992_, data_stage_4__1991_, data_stage_4__1990_, data_stage_4__1989_, data_stage_4__1988_, data_stage_4__1987_, data_stage_4__1986_, data_stage_4__1985_, data_stage_4__1984_, data_stage_4__1983_, data_stage_4__1982_, data_stage_4__1981_, data_stage_4__1980_, data_stage_4__1979_, data_stage_4__1978_, data_stage_4__1977_, data_stage_4__1976_, data_stage_4__1975_, data_stage_4__1974_, data_stage_4__1973_, data_stage_4__1972_, data_stage_4__1971_, data_stage_4__1970_, data_stage_4__1969_, data_stage_4__1968_, data_stage_4__1967_, data_stage_4__1966_, data_stage_4__1965_, data_stage_4__1964_, data_stage_4__1963_, data_stage_4__1962_, data_stage_4__1961_, data_stage_4__1960_, data_stage_4__1959_, data_stage_4__1958_, data_stage_4__1957_, data_stage_4__1956_, data_stage_4__1955_, data_stage_4__1954_, data_stage_4__1953_, data_stage_4__1952_, data_stage_4__1951_, data_stage_4__1950_, data_stage_4__1949_, data_stage_4__1948_, data_stage_4__1947_, data_stage_4__1946_, data_stage_4__1945_, data_stage_4__1944_, data_stage_4__1943_, data_stage_4__1942_, data_stage_4__1941_, data_stage_4__1940_, data_stage_4__1939_, data_stage_4__1938_, data_stage_4__1937_, data_stage_4__1936_, data_stage_4__1935_, data_stage_4__1934_, data_stage_4__1933_, data_stage_4__1932_, data_stage_4__1931_, data_stage_4__1930_, data_stage_4__1929_, data_stage_4__1928_, data_stage_4__1927_, data_stage_4__1926_, data_stage_4__1925_, data_stage_4__1924_, data_stage_4__1923_, data_stage_4__1922_, data_stage_4__1921_, data_stage_4__1920_, data_stage_4__1919_, data_stage_4__1918_, data_stage_4__1917_, data_stage_4__1916_, data_stage_4__1915_, data_stage_4__1914_, data_stage_4__1913_, data_stage_4__1912_, data_stage_4__1911_, data_stage_4__1910_, data_stage_4__1909_, data_stage_4__1908_, data_stage_4__1907_, data_stage_4__1906_, data_stage_4__1905_, data_stage_4__1904_, data_stage_4__1903_, data_stage_4__1902_, data_stage_4__1901_, data_stage_4__1900_, data_stage_4__1899_, data_stage_4__1898_, data_stage_4__1897_, data_stage_4__1896_, data_stage_4__1895_, data_stage_4__1894_, data_stage_4__1893_, data_stage_4__1892_, data_stage_4__1891_, data_stage_4__1890_, data_stage_4__1889_, data_stage_4__1888_, data_stage_4__1887_, data_stage_4__1886_, data_stage_4__1885_, data_stage_4__1884_, data_stage_4__1883_, data_stage_4__1882_, data_stage_4__1881_, data_stage_4__1880_, data_stage_4__1879_, data_stage_4__1878_, data_stage_4__1877_, data_stage_4__1876_, data_stage_4__1875_, data_stage_4__1874_, data_stage_4__1873_, data_stage_4__1872_, data_stage_4__1871_, data_stage_4__1870_, data_stage_4__1869_, data_stage_4__1868_, data_stage_4__1867_, data_stage_4__1866_, data_stage_4__1865_, data_stage_4__1864_, data_stage_4__1863_, data_stage_4__1862_, data_stage_4__1861_, data_stage_4__1860_, data_stage_4__1859_, data_stage_4__1858_, data_stage_4__1857_, data_stage_4__1856_, data_stage_4__1855_, data_stage_4__1854_, data_stage_4__1853_, data_stage_4__1852_, data_stage_4__1851_, data_stage_4__1850_, data_stage_4__1849_, data_stage_4__1848_, data_stage_4__1847_, data_stage_4__1846_, data_stage_4__1845_, data_stage_4__1844_, data_stage_4__1843_, data_stage_4__1842_, data_stage_4__1841_, data_stage_4__1840_, data_stage_4__1839_, data_stage_4__1838_, data_stage_4__1837_, data_stage_4__1836_, data_stage_4__1835_, data_stage_4__1834_, data_stage_4__1833_, data_stage_4__1832_, data_stage_4__1831_, data_stage_4__1830_, data_stage_4__1829_, data_stage_4__1828_, data_stage_4__1827_, data_stage_4__1826_, data_stage_4__1825_, data_stage_4__1824_, data_stage_4__1823_, data_stage_4__1822_, data_stage_4__1821_, data_stage_4__1820_, data_stage_4__1819_, data_stage_4__1818_, data_stage_4__1817_, data_stage_4__1816_, data_stage_4__1815_, data_stage_4__1814_, data_stage_4__1813_, data_stage_4__1812_, data_stage_4__1811_, data_stage_4__1810_, data_stage_4__1809_, data_stage_4__1808_, data_stage_4__1807_, data_stage_4__1806_, data_stage_4__1805_, data_stage_4__1804_, data_stage_4__1803_, data_stage_4__1802_, data_stage_4__1801_, data_stage_4__1800_, data_stage_4__1799_, data_stage_4__1798_, data_stage_4__1797_, data_stage_4__1796_, data_stage_4__1795_, data_stage_4__1794_, data_stage_4__1793_, data_stage_4__1792_, data_stage_4__1791_, data_stage_4__1790_, data_stage_4__1789_, data_stage_4__1788_, data_stage_4__1787_, data_stage_4__1786_, data_stage_4__1785_, data_stage_4__1784_, data_stage_4__1783_, data_stage_4__1782_, data_stage_4__1781_, data_stage_4__1780_, data_stage_4__1779_, data_stage_4__1778_, data_stage_4__1777_, data_stage_4__1776_, data_stage_4__1775_, data_stage_4__1774_, data_stage_4__1773_, data_stage_4__1772_, data_stage_4__1771_, data_stage_4__1770_, data_stage_4__1769_, data_stage_4__1768_, data_stage_4__1767_, data_stage_4__1766_, data_stage_4__1765_, data_stage_4__1764_, data_stage_4__1763_, data_stage_4__1762_, data_stage_4__1761_, data_stage_4__1760_, data_stage_4__1759_, data_stage_4__1758_, data_stage_4__1757_, data_stage_4__1756_, data_stage_4__1755_, data_stage_4__1754_, data_stage_4__1753_, data_stage_4__1752_, data_stage_4__1751_, data_stage_4__1750_, data_stage_4__1749_, data_stage_4__1748_, data_stage_4__1747_, data_stage_4__1746_, data_stage_4__1745_, data_stage_4__1744_, data_stage_4__1743_, data_stage_4__1742_, data_stage_4__1741_, data_stage_4__1740_, data_stage_4__1739_, data_stage_4__1738_, data_stage_4__1737_, data_stage_4__1736_, data_stage_4__1735_, data_stage_4__1734_, data_stage_4__1733_, data_stage_4__1732_, data_stage_4__1731_, data_stage_4__1730_, data_stage_4__1729_, data_stage_4__1728_, data_stage_4__1727_, data_stage_4__1726_, data_stage_4__1725_, data_stage_4__1724_, data_stage_4__1723_, data_stage_4__1722_, data_stage_4__1721_, data_stage_4__1720_, data_stage_4__1719_, data_stage_4__1718_, data_stage_4__1717_, data_stage_4__1716_, data_stage_4__1715_, data_stage_4__1714_, data_stage_4__1713_, data_stage_4__1712_, data_stage_4__1711_, data_stage_4__1710_, data_stage_4__1709_, data_stage_4__1708_, data_stage_4__1707_, data_stage_4__1706_, data_stage_4__1705_, data_stage_4__1704_, data_stage_4__1703_, data_stage_4__1702_, data_stage_4__1701_, data_stage_4__1700_, data_stage_4__1699_, data_stage_4__1698_, data_stage_4__1697_, data_stage_4__1696_, data_stage_4__1695_, data_stage_4__1694_, data_stage_4__1693_, data_stage_4__1692_, data_stage_4__1691_, data_stage_4__1690_, data_stage_4__1689_, data_stage_4__1688_, data_stage_4__1687_, data_stage_4__1686_, data_stage_4__1685_, data_stage_4__1684_, data_stage_4__1683_, data_stage_4__1682_, data_stage_4__1681_, data_stage_4__1680_, data_stage_4__1679_, data_stage_4__1678_, data_stage_4__1677_, data_stage_4__1676_, data_stage_4__1675_, data_stage_4__1674_, data_stage_4__1673_, data_stage_4__1672_, data_stage_4__1671_, data_stage_4__1670_, data_stage_4__1669_, data_stage_4__1668_, data_stage_4__1667_, data_stage_4__1666_, data_stage_4__1665_, data_stage_4__1664_, data_stage_4__1663_, data_stage_4__1662_, data_stage_4__1661_, data_stage_4__1660_, data_stage_4__1659_, data_stage_4__1658_, data_stage_4__1657_, data_stage_4__1656_, data_stage_4__1655_, data_stage_4__1654_, data_stage_4__1653_, data_stage_4__1652_, data_stage_4__1651_, data_stage_4__1650_, data_stage_4__1649_, data_stage_4__1648_, data_stage_4__1647_, data_stage_4__1646_, data_stage_4__1645_, data_stage_4__1644_, data_stage_4__1643_, data_stage_4__1642_, data_stage_4__1641_, data_stage_4__1640_, data_stage_4__1639_, data_stage_4__1638_, data_stage_4__1637_, data_stage_4__1636_, data_stage_4__1635_, data_stage_4__1634_, data_stage_4__1633_, data_stage_4__1632_, data_stage_4__1631_, data_stage_4__1630_, data_stage_4__1629_, data_stage_4__1628_, data_stage_4__1627_, data_stage_4__1626_, data_stage_4__1625_, data_stage_4__1624_, data_stage_4__1623_, data_stage_4__1622_, data_stage_4__1621_, data_stage_4__1620_, data_stage_4__1619_, data_stage_4__1618_, data_stage_4__1617_, data_stage_4__1616_, data_stage_4__1615_, data_stage_4__1614_, data_stage_4__1613_, data_stage_4__1612_, data_stage_4__1611_, data_stage_4__1610_, data_stage_4__1609_, data_stage_4__1608_, data_stage_4__1607_, data_stage_4__1606_, data_stage_4__1605_, data_stage_4__1604_, data_stage_4__1603_, data_stage_4__1602_, data_stage_4__1601_, data_stage_4__1600_, data_stage_4__1599_, data_stage_4__1598_, data_stage_4__1597_, data_stage_4__1596_, data_stage_4__1595_, data_stage_4__1594_, data_stage_4__1593_, data_stage_4__1592_, data_stage_4__1591_, data_stage_4__1590_, data_stage_4__1589_, data_stage_4__1588_, data_stage_4__1587_, data_stage_4__1586_, data_stage_4__1585_, data_stage_4__1584_, data_stage_4__1583_, data_stage_4__1582_, data_stage_4__1581_, data_stage_4__1580_, data_stage_4__1579_, data_stage_4__1578_, data_stage_4__1577_, data_stage_4__1576_, data_stage_4__1575_, data_stage_4__1574_, data_stage_4__1573_, data_stage_4__1572_, data_stage_4__1571_, data_stage_4__1570_, data_stage_4__1569_, data_stage_4__1568_, data_stage_4__1567_, data_stage_4__1566_, data_stage_4__1565_, data_stage_4__1564_, data_stage_4__1563_, data_stage_4__1562_, data_stage_4__1561_, data_stage_4__1560_, data_stage_4__1559_, data_stage_4__1558_, data_stage_4__1557_, data_stage_4__1556_, data_stage_4__1555_, data_stage_4__1554_, data_stage_4__1553_, data_stage_4__1552_, data_stage_4__1551_, data_stage_4__1550_, data_stage_4__1549_, data_stage_4__1548_, data_stage_4__1547_, data_stage_4__1546_, data_stage_4__1545_, data_stage_4__1544_, data_stage_4__1543_, data_stage_4__1542_, data_stage_4__1541_, data_stage_4__1540_, data_stage_4__1539_, data_stage_4__1538_, data_stage_4__1537_, data_stage_4__1536_, data_stage_4__1535_, data_stage_4__1534_, data_stage_4__1533_, data_stage_4__1532_, data_stage_4__1531_, data_stage_4__1530_, data_stage_4__1529_, data_stage_4__1528_, data_stage_4__1527_, data_stage_4__1526_, data_stage_4__1525_, data_stage_4__1524_, data_stage_4__1523_, data_stage_4__1522_, data_stage_4__1521_, data_stage_4__1520_, data_stage_4__1519_, data_stage_4__1518_, data_stage_4__1517_, data_stage_4__1516_, data_stage_4__1515_, data_stage_4__1514_, data_stage_4__1513_, data_stage_4__1512_, data_stage_4__1511_, data_stage_4__1510_, data_stage_4__1509_, data_stage_4__1508_, data_stage_4__1507_, data_stage_4__1506_, data_stage_4__1505_, data_stage_4__1504_, data_stage_4__1503_, data_stage_4__1502_, data_stage_4__1501_, data_stage_4__1500_, data_stage_4__1499_, data_stage_4__1498_, data_stage_4__1497_, data_stage_4__1496_, data_stage_4__1495_, data_stage_4__1494_, data_stage_4__1493_, data_stage_4__1492_, data_stage_4__1491_, data_stage_4__1490_, data_stage_4__1489_, data_stage_4__1488_, data_stage_4__1487_, data_stage_4__1486_, data_stage_4__1485_, data_stage_4__1484_, data_stage_4__1483_, data_stage_4__1482_, data_stage_4__1481_, data_stage_4__1480_, data_stage_4__1479_, data_stage_4__1478_, data_stage_4__1477_, data_stage_4__1476_, data_stage_4__1475_, data_stage_4__1474_, data_stage_4__1473_, data_stage_4__1472_, data_stage_4__1471_, data_stage_4__1470_, data_stage_4__1469_, data_stage_4__1468_, data_stage_4__1467_, data_stage_4__1466_, data_stage_4__1465_, data_stage_4__1464_, data_stage_4__1463_, data_stage_4__1462_, data_stage_4__1461_, data_stage_4__1460_, data_stage_4__1459_, data_stage_4__1458_, data_stage_4__1457_, data_stage_4__1456_, data_stage_4__1455_, data_stage_4__1454_, data_stage_4__1453_, data_stage_4__1452_, data_stage_4__1451_, data_stage_4__1450_, data_stage_4__1449_, data_stage_4__1448_, data_stage_4__1447_, data_stage_4__1446_, data_stage_4__1445_, data_stage_4__1444_, data_stage_4__1443_, data_stage_4__1442_, data_stage_4__1441_, data_stage_4__1440_, data_stage_4__1439_, data_stage_4__1438_, data_stage_4__1437_, data_stage_4__1436_, data_stage_4__1435_, data_stage_4__1434_, data_stage_4__1433_, data_stage_4__1432_, data_stage_4__1431_, data_stage_4__1430_, data_stage_4__1429_, data_stage_4__1428_, data_stage_4__1427_, data_stage_4__1426_, data_stage_4__1425_, data_stage_4__1424_, data_stage_4__1423_, data_stage_4__1422_, data_stage_4__1421_, data_stage_4__1420_, data_stage_4__1419_, data_stage_4__1418_, data_stage_4__1417_, data_stage_4__1416_, data_stage_4__1415_, data_stage_4__1414_, data_stage_4__1413_, data_stage_4__1412_, data_stage_4__1411_, data_stage_4__1410_, data_stage_4__1409_, data_stage_4__1408_, data_stage_4__1407_, data_stage_4__1406_, data_stage_4__1405_, data_stage_4__1404_, data_stage_4__1403_, data_stage_4__1402_, data_stage_4__1401_, data_stage_4__1400_, data_stage_4__1399_, data_stage_4__1398_, data_stage_4__1397_, data_stage_4__1396_, data_stage_4__1395_, data_stage_4__1394_, data_stage_4__1393_, data_stage_4__1392_, data_stage_4__1391_, data_stage_4__1390_, data_stage_4__1389_, data_stage_4__1388_, data_stage_4__1387_, data_stage_4__1386_, data_stage_4__1385_, data_stage_4__1384_, data_stage_4__1383_, data_stage_4__1382_, data_stage_4__1381_, data_stage_4__1380_, data_stage_4__1379_, data_stage_4__1378_, data_stage_4__1377_, data_stage_4__1376_, data_stage_4__1375_, data_stage_4__1374_, data_stage_4__1373_, data_stage_4__1372_, data_stage_4__1371_, data_stage_4__1370_, data_stage_4__1369_, data_stage_4__1368_, data_stage_4__1367_, data_stage_4__1366_, data_stage_4__1365_, data_stage_4__1364_, data_stage_4__1363_, data_stage_4__1362_, data_stage_4__1361_, data_stage_4__1360_, data_stage_4__1359_, data_stage_4__1358_, data_stage_4__1357_, data_stage_4__1356_, data_stage_4__1355_, data_stage_4__1354_, data_stage_4__1353_, data_stage_4__1352_, data_stage_4__1351_, data_stage_4__1350_, data_stage_4__1349_, data_stage_4__1348_, data_stage_4__1347_, data_stage_4__1346_, data_stage_4__1345_, data_stage_4__1344_, data_stage_4__1343_, data_stage_4__1342_, data_stage_4__1341_, data_stage_4__1340_, data_stage_4__1339_, data_stage_4__1338_, data_stage_4__1337_, data_stage_4__1336_, data_stage_4__1335_, data_stage_4__1334_, data_stage_4__1333_, data_stage_4__1332_, data_stage_4__1331_, data_stage_4__1330_, data_stage_4__1329_, data_stage_4__1328_, data_stage_4__1327_, data_stage_4__1326_, data_stage_4__1325_, data_stage_4__1324_, data_stage_4__1323_, data_stage_4__1322_, data_stage_4__1321_, data_stage_4__1320_, data_stage_4__1319_, data_stage_4__1318_, data_stage_4__1317_, data_stage_4__1316_, data_stage_4__1315_, data_stage_4__1314_, data_stage_4__1313_, data_stage_4__1312_, data_stage_4__1311_, data_stage_4__1310_, data_stage_4__1309_, data_stage_4__1308_, data_stage_4__1307_, data_stage_4__1306_, data_stage_4__1305_, data_stage_4__1304_, data_stage_4__1303_, data_stage_4__1302_, data_stage_4__1301_, data_stage_4__1300_, data_stage_4__1299_, data_stage_4__1298_, data_stage_4__1297_, data_stage_4__1296_, data_stage_4__1295_, data_stage_4__1294_, data_stage_4__1293_, data_stage_4__1292_, data_stage_4__1291_, data_stage_4__1290_, data_stage_4__1289_, data_stage_4__1288_, data_stage_4__1287_, data_stage_4__1286_, data_stage_4__1285_, data_stage_4__1284_, data_stage_4__1283_, data_stage_4__1282_, data_stage_4__1281_, data_stage_4__1280_, data_stage_4__1279_, data_stage_4__1278_, data_stage_4__1277_, data_stage_4__1276_, data_stage_4__1275_, data_stage_4__1274_, data_stage_4__1273_, data_stage_4__1272_, data_stage_4__1271_, data_stage_4__1270_, data_stage_4__1269_, data_stage_4__1268_, data_stage_4__1267_, data_stage_4__1266_, data_stage_4__1265_, data_stage_4__1264_, data_stage_4__1263_, data_stage_4__1262_, data_stage_4__1261_, data_stage_4__1260_, data_stage_4__1259_, data_stage_4__1258_, data_stage_4__1257_, data_stage_4__1256_, data_stage_4__1255_, data_stage_4__1254_, data_stage_4__1253_, data_stage_4__1252_, data_stage_4__1251_, data_stage_4__1250_, data_stage_4__1249_, data_stage_4__1248_, data_stage_4__1247_, data_stage_4__1246_, data_stage_4__1245_, data_stage_4__1244_, data_stage_4__1243_, data_stage_4__1242_, data_stage_4__1241_, data_stage_4__1240_, data_stage_4__1239_, data_stage_4__1238_, data_stage_4__1237_, data_stage_4__1236_, data_stage_4__1235_, data_stage_4__1234_, data_stage_4__1233_, data_stage_4__1232_, data_stage_4__1231_, data_stage_4__1230_, data_stage_4__1229_, data_stage_4__1228_, data_stage_4__1227_, data_stage_4__1226_, data_stage_4__1225_, data_stage_4__1224_, data_stage_4__1223_, data_stage_4__1222_, data_stage_4__1221_, data_stage_4__1220_, data_stage_4__1219_, data_stage_4__1218_, data_stage_4__1217_, data_stage_4__1216_, data_stage_4__1215_, data_stage_4__1214_, data_stage_4__1213_, data_stage_4__1212_, data_stage_4__1211_, data_stage_4__1210_, data_stage_4__1209_, data_stage_4__1208_, data_stage_4__1207_, data_stage_4__1206_, data_stage_4__1205_, data_stage_4__1204_, data_stage_4__1203_, data_stage_4__1202_, data_stage_4__1201_, data_stage_4__1200_, data_stage_4__1199_, data_stage_4__1198_, data_stage_4__1197_, data_stage_4__1196_, data_stage_4__1195_, data_stage_4__1194_, data_stage_4__1193_, data_stage_4__1192_, data_stage_4__1191_, data_stage_4__1190_, data_stage_4__1189_, data_stage_4__1188_, data_stage_4__1187_, data_stage_4__1186_, data_stage_4__1185_, data_stage_4__1184_, data_stage_4__1183_, data_stage_4__1182_, data_stage_4__1181_, data_stage_4__1180_, data_stage_4__1179_, data_stage_4__1178_, data_stage_4__1177_, data_stage_4__1176_, data_stage_4__1175_, data_stage_4__1174_, data_stage_4__1173_, data_stage_4__1172_, data_stage_4__1171_, data_stage_4__1170_, data_stage_4__1169_, data_stage_4__1168_, data_stage_4__1167_, data_stage_4__1166_, data_stage_4__1165_, data_stage_4__1164_, data_stage_4__1163_, data_stage_4__1162_, data_stage_4__1161_, data_stage_4__1160_, data_stage_4__1159_, data_stage_4__1158_, data_stage_4__1157_, data_stage_4__1156_, data_stage_4__1155_, data_stage_4__1154_, data_stage_4__1153_, data_stage_4__1152_, data_stage_4__1151_, data_stage_4__1150_, data_stage_4__1149_, data_stage_4__1148_, data_stage_4__1147_, data_stage_4__1146_, data_stage_4__1145_, data_stage_4__1144_, data_stage_4__1143_, data_stage_4__1142_, data_stage_4__1141_, data_stage_4__1140_, data_stage_4__1139_, data_stage_4__1138_, data_stage_4__1137_, data_stage_4__1136_, data_stage_4__1135_, data_stage_4__1134_, data_stage_4__1133_, data_stage_4__1132_, data_stage_4__1131_, data_stage_4__1130_, data_stage_4__1129_, data_stage_4__1128_, data_stage_4__1127_, data_stage_4__1126_, data_stage_4__1125_, data_stage_4__1124_, data_stage_4__1123_, data_stage_4__1122_, data_stage_4__1121_, data_stage_4__1120_, data_stage_4__1119_, data_stage_4__1118_, data_stage_4__1117_, data_stage_4__1116_, data_stage_4__1115_, data_stage_4__1114_, data_stage_4__1113_, data_stage_4__1112_, data_stage_4__1111_, data_stage_4__1110_, data_stage_4__1109_, data_stage_4__1108_, data_stage_4__1107_, data_stage_4__1106_, data_stage_4__1105_, data_stage_4__1104_, data_stage_4__1103_, data_stage_4__1102_, data_stage_4__1101_, data_stage_4__1100_, data_stage_4__1099_, data_stage_4__1098_, data_stage_4__1097_, data_stage_4__1096_, data_stage_4__1095_, data_stage_4__1094_, data_stage_4__1093_, data_stage_4__1092_, data_stage_4__1091_, data_stage_4__1090_, data_stage_4__1089_, data_stage_4__1088_, data_stage_4__1087_, data_stage_4__1086_, data_stage_4__1085_, data_stage_4__1084_, data_stage_4__1083_, data_stage_4__1082_, data_stage_4__1081_, data_stage_4__1080_, data_stage_4__1079_, data_stage_4__1078_, data_stage_4__1077_, data_stage_4__1076_, data_stage_4__1075_, data_stage_4__1074_, data_stage_4__1073_, data_stage_4__1072_, data_stage_4__1071_, data_stage_4__1070_, data_stage_4__1069_, data_stage_4__1068_, data_stage_4__1067_, data_stage_4__1066_, data_stage_4__1065_, data_stage_4__1064_, data_stage_4__1063_, data_stage_4__1062_, data_stage_4__1061_, data_stage_4__1060_, data_stage_4__1059_, data_stage_4__1058_, data_stage_4__1057_, data_stage_4__1056_, data_stage_4__1055_, data_stage_4__1054_, data_stage_4__1053_, data_stage_4__1052_, data_stage_4__1051_, data_stage_4__1050_, data_stage_4__1049_, data_stage_4__1048_, data_stage_4__1047_, data_stage_4__1046_, data_stage_4__1045_, data_stage_4__1044_, data_stage_4__1043_, data_stage_4__1042_, data_stage_4__1041_, data_stage_4__1040_, data_stage_4__1039_, data_stage_4__1038_, data_stage_4__1037_, data_stage_4__1036_, data_stage_4__1035_, data_stage_4__1034_, data_stage_4__1033_, data_stage_4__1032_, data_stage_4__1031_, data_stage_4__1030_, data_stage_4__1029_, data_stage_4__1028_, data_stage_4__1027_, data_stage_4__1026_, data_stage_4__1025_, data_stage_4__1024_, data_stage_4__1023_, data_stage_4__1022_, data_stage_4__1021_, data_stage_4__1020_, data_stage_4__1019_, data_stage_4__1018_, data_stage_4__1017_, data_stage_4__1016_, data_stage_4__1015_, data_stage_4__1014_, data_stage_4__1013_, data_stage_4__1012_, data_stage_4__1011_, data_stage_4__1010_, data_stage_4__1009_, data_stage_4__1008_, data_stage_4__1007_, data_stage_4__1006_, data_stage_4__1005_, data_stage_4__1004_, data_stage_4__1003_, data_stage_4__1002_, data_stage_4__1001_, data_stage_4__1000_, data_stage_4__999_, data_stage_4__998_, data_stage_4__997_, data_stage_4__996_, data_stage_4__995_, data_stage_4__994_, data_stage_4__993_, data_stage_4__992_, data_stage_4__991_, data_stage_4__990_, data_stage_4__989_, data_stage_4__988_, data_stage_4__987_, data_stage_4__986_, data_stage_4__985_, data_stage_4__984_, data_stage_4__983_, data_stage_4__982_, data_stage_4__981_, data_stage_4__980_, data_stage_4__979_, data_stage_4__978_, data_stage_4__977_, data_stage_4__976_, data_stage_4__975_, data_stage_4__974_, data_stage_4__973_, data_stage_4__972_, data_stage_4__971_, data_stage_4__970_, data_stage_4__969_, data_stage_4__968_, data_stage_4__967_, data_stage_4__966_, data_stage_4__965_, data_stage_4__964_, data_stage_4__963_, data_stage_4__962_, data_stage_4__961_, data_stage_4__960_, data_stage_4__959_, data_stage_4__958_, data_stage_4__957_, data_stage_4__956_, data_stage_4__955_, data_stage_4__954_, data_stage_4__953_, data_stage_4__952_, data_stage_4__951_, data_stage_4__950_, data_stage_4__949_, data_stage_4__948_, data_stage_4__947_, data_stage_4__946_, data_stage_4__945_, data_stage_4__944_, data_stage_4__943_, data_stage_4__942_, data_stage_4__941_, data_stage_4__940_, data_stage_4__939_, data_stage_4__938_, data_stage_4__937_, data_stage_4__936_, data_stage_4__935_, data_stage_4__934_, data_stage_4__933_, data_stage_4__932_, data_stage_4__931_, data_stage_4__930_, data_stage_4__929_, data_stage_4__928_, data_stage_4__927_, data_stage_4__926_, data_stage_4__925_, data_stage_4__924_, data_stage_4__923_, data_stage_4__922_, data_stage_4__921_, data_stage_4__920_, data_stage_4__919_, data_stage_4__918_, data_stage_4__917_, data_stage_4__916_, data_stage_4__915_, data_stage_4__914_, data_stage_4__913_, data_stage_4__912_, data_stage_4__911_, data_stage_4__910_, data_stage_4__909_, data_stage_4__908_, data_stage_4__907_, data_stage_4__906_, data_stage_4__905_, data_stage_4__904_, data_stage_4__903_, data_stage_4__902_, data_stage_4__901_, data_stage_4__900_, data_stage_4__899_, data_stage_4__898_, data_stage_4__897_, data_stage_4__896_, data_stage_4__895_, data_stage_4__894_, data_stage_4__893_, data_stage_4__892_, data_stage_4__891_, data_stage_4__890_, data_stage_4__889_, data_stage_4__888_, data_stage_4__887_, data_stage_4__886_, data_stage_4__885_, data_stage_4__884_, data_stage_4__883_, data_stage_4__882_, data_stage_4__881_, data_stage_4__880_, data_stage_4__879_, data_stage_4__878_, data_stage_4__877_, data_stage_4__876_, data_stage_4__875_, data_stage_4__874_, data_stage_4__873_, data_stage_4__872_, data_stage_4__871_, data_stage_4__870_, data_stage_4__869_, data_stage_4__868_, data_stage_4__867_, data_stage_4__866_, data_stage_4__865_, data_stage_4__864_, data_stage_4__863_, data_stage_4__862_, data_stage_4__861_, data_stage_4__860_, data_stage_4__859_, data_stage_4__858_, data_stage_4__857_, data_stage_4__856_, data_stage_4__855_, data_stage_4__854_, data_stage_4__853_, data_stage_4__852_, data_stage_4__851_, data_stage_4__850_, data_stage_4__849_, data_stage_4__848_, data_stage_4__847_, data_stage_4__846_, data_stage_4__845_, data_stage_4__844_, data_stage_4__843_, data_stage_4__842_, data_stage_4__841_, data_stage_4__840_, data_stage_4__839_, data_stage_4__838_, data_stage_4__837_, data_stage_4__836_, data_stage_4__835_, data_stage_4__834_, data_stage_4__833_, data_stage_4__832_, data_stage_4__831_, data_stage_4__830_, data_stage_4__829_, data_stage_4__828_, data_stage_4__827_, data_stage_4__826_, data_stage_4__825_, data_stage_4__824_, data_stage_4__823_, data_stage_4__822_, data_stage_4__821_, data_stage_4__820_, data_stage_4__819_, data_stage_4__818_, data_stage_4__817_, data_stage_4__816_, data_stage_4__815_, data_stage_4__814_, data_stage_4__813_, data_stage_4__812_, data_stage_4__811_, data_stage_4__810_, data_stage_4__809_, data_stage_4__808_, data_stage_4__807_, data_stage_4__806_, data_stage_4__805_, data_stage_4__804_, data_stage_4__803_, data_stage_4__802_, data_stage_4__801_, data_stage_4__800_, data_stage_4__799_, data_stage_4__798_, data_stage_4__797_, data_stage_4__796_, data_stage_4__795_, data_stage_4__794_, data_stage_4__793_, data_stage_4__792_, data_stage_4__791_, data_stage_4__790_, data_stage_4__789_, data_stage_4__788_, data_stage_4__787_, data_stage_4__786_, data_stage_4__785_, data_stage_4__784_, data_stage_4__783_, data_stage_4__782_, data_stage_4__781_, data_stage_4__780_, data_stage_4__779_, data_stage_4__778_, data_stage_4__777_, data_stage_4__776_, data_stage_4__775_, data_stage_4__774_, data_stage_4__773_, data_stage_4__772_, data_stage_4__771_, data_stage_4__770_, data_stage_4__769_, data_stage_4__768_, data_stage_4__767_, data_stage_4__766_, data_stage_4__765_, data_stage_4__764_, data_stage_4__763_, data_stage_4__762_, data_stage_4__761_, data_stage_4__760_, data_stage_4__759_, data_stage_4__758_, data_stage_4__757_, data_stage_4__756_, data_stage_4__755_, data_stage_4__754_, data_stage_4__753_, data_stage_4__752_, data_stage_4__751_, data_stage_4__750_, data_stage_4__749_, data_stage_4__748_, data_stage_4__747_, data_stage_4__746_, data_stage_4__745_, data_stage_4__744_, data_stage_4__743_, data_stage_4__742_, data_stage_4__741_, data_stage_4__740_, data_stage_4__739_, data_stage_4__738_, data_stage_4__737_, data_stage_4__736_, data_stage_4__735_, data_stage_4__734_, data_stage_4__733_, data_stage_4__732_, data_stage_4__731_, data_stage_4__730_, data_stage_4__729_, data_stage_4__728_, data_stage_4__727_, data_stage_4__726_, data_stage_4__725_, data_stage_4__724_, data_stage_4__723_, data_stage_4__722_, data_stage_4__721_, data_stage_4__720_, data_stage_4__719_, data_stage_4__718_, data_stage_4__717_, data_stage_4__716_, data_stage_4__715_, data_stage_4__714_, data_stage_4__713_, data_stage_4__712_, data_stage_4__711_, data_stage_4__710_, data_stage_4__709_, data_stage_4__708_, data_stage_4__707_, data_stage_4__706_, data_stage_4__705_, data_stage_4__704_, data_stage_4__703_, data_stage_4__702_, data_stage_4__701_, data_stage_4__700_, data_stage_4__699_, data_stage_4__698_, data_stage_4__697_, data_stage_4__696_, data_stage_4__695_, data_stage_4__694_, data_stage_4__693_, data_stage_4__692_, data_stage_4__691_, data_stage_4__690_, data_stage_4__689_, data_stage_4__688_, data_stage_4__687_, data_stage_4__686_, data_stage_4__685_, data_stage_4__684_, data_stage_4__683_, data_stage_4__682_, data_stage_4__681_, data_stage_4__680_, data_stage_4__679_, data_stage_4__678_, data_stage_4__677_, data_stage_4__676_, data_stage_4__675_, data_stage_4__674_, data_stage_4__673_, data_stage_4__672_, data_stage_4__671_, data_stage_4__670_, data_stage_4__669_, data_stage_4__668_, data_stage_4__667_, data_stage_4__666_, data_stage_4__665_, data_stage_4__664_, data_stage_4__663_, data_stage_4__662_, data_stage_4__661_, data_stage_4__660_, data_stage_4__659_, data_stage_4__658_, data_stage_4__657_, data_stage_4__656_, data_stage_4__655_, data_stage_4__654_, data_stage_4__653_, data_stage_4__652_, data_stage_4__651_, data_stage_4__650_, data_stage_4__649_, data_stage_4__648_, data_stage_4__647_, data_stage_4__646_, data_stage_4__645_, data_stage_4__644_, data_stage_4__643_, data_stage_4__642_, data_stage_4__641_, data_stage_4__640_, data_stage_4__639_, data_stage_4__638_, data_stage_4__637_, data_stage_4__636_, data_stage_4__635_, data_stage_4__634_, data_stage_4__633_, data_stage_4__632_, data_stage_4__631_, data_stage_4__630_, data_stage_4__629_, data_stage_4__628_, data_stage_4__627_, data_stage_4__626_, data_stage_4__625_, data_stage_4__624_, data_stage_4__623_, data_stage_4__622_, data_stage_4__621_, data_stage_4__620_, data_stage_4__619_, data_stage_4__618_, data_stage_4__617_, data_stage_4__616_, data_stage_4__615_, data_stage_4__614_, data_stage_4__613_, data_stage_4__612_, data_stage_4__611_, data_stage_4__610_, data_stage_4__609_, data_stage_4__608_, data_stage_4__607_, data_stage_4__606_, data_stage_4__605_, data_stage_4__604_, data_stage_4__603_, data_stage_4__602_, data_stage_4__601_, data_stage_4__600_, data_stage_4__599_, data_stage_4__598_, data_stage_4__597_, data_stage_4__596_, data_stage_4__595_, data_stage_4__594_, data_stage_4__593_, data_stage_4__592_, data_stage_4__591_, data_stage_4__590_, data_stage_4__589_, data_stage_4__588_, data_stage_4__587_, data_stage_4__586_, data_stage_4__585_, data_stage_4__584_, data_stage_4__583_, data_stage_4__582_, data_stage_4__581_, data_stage_4__580_, data_stage_4__579_, data_stage_4__578_, data_stage_4__577_, data_stage_4__576_, data_stage_4__575_, data_stage_4__574_, data_stage_4__573_, data_stage_4__572_, data_stage_4__571_, data_stage_4__570_, data_stage_4__569_, data_stage_4__568_, data_stage_4__567_, data_stage_4__566_, data_stage_4__565_, data_stage_4__564_, data_stage_4__563_, data_stage_4__562_, data_stage_4__561_, data_stage_4__560_, data_stage_4__559_, data_stage_4__558_, data_stage_4__557_, data_stage_4__556_, data_stage_4__555_, data_stage_4__554_, data_stage_4__553_, data_stage_4__552_, data_stage_4__551_, data_stage_4__550_, data_stage_4__549_, data_stage_4__548_, data_stage_4__547_, data_stage_4__546_, data_stage_4__545_, data_stage_4__544_, data_stage_4__543_, data_stage_4__542_, data_stage_4__541_, data_stage_4__540_, data_stage_4__539_, data_stage_4__538_, data_stage_4__537_, data_stage_4__536_, data_stage_4__535_, data_stage_4__534_, data_stage_4__533_, data_stage_4__532_, data_stage_4__531_, data_stage_4__530_, data_stage_4__529_, data_stage_4__528_, data_stage_4__527_, data_stage_4__526_, data_stage_4__525_, data_stage_4__524_, data_stage_4__523_, data_stage_4__522_, data_stage_4__521_, data_stage_4__520_, data_stage_4__519_, data_stage_4__518_, data_stage_4__517_, data_stage_4__516_, data_stage_4__515_, data_stage_4__514_, data_stage_4__513_, data_stage_4__512_, data_stage_4__511_, data_stage_4__510_, data_stage_4__509_, data_stage_4__508_, data_stage_4__507_, data_stage_4__506_, data_stage_4__505_, data_stage_4__504_, data_stage_4__503_, data_stage_4__502_, data_stage_4__501_, data_stage_4__500_, data_stage_4__499_, data_stage_4__498_, data_stage_4__497_, data_stage_4__496_, data_stage_4__495_, data_stage_4__494_, data_stage_4__493_, data_stage_4__492_, data_stage_4__491_, data_stage_4__490_, data_stage_4__489_, data_stage_4__488_, data_stage_4__487_, data_stage_4__486_, data_stage_4__485_, data_stage_4__484_, data_stage_4__483_, data_stage_4__482_, data_stage_4__481_, data_stage_4__480_, data_stage_4__479_, data_stage_4__478_, data_stage_4__477_, data_stage_4__476_, data_stage_4__475_, data_stage_4__474_, data_stage_4__473_, data_stage_4__472_, data_stage_4__471_, data_stage_4__470_, data_stage_4__469_, data_stage_4__468_, data_stage_4__467_, data_stage_4__466_, data_stage_4__465_, data_stage_4__464_, data_stage_4__463_, data_stage_4__462_, data_stage_4__461_, data_stage_4__460_, data_stage_4__459_, data_stage_4__458_, data_stage_4__457_, data_stage_4__456_, data_stage_4__455_, data_stage_4__454_, data_stage_4__453_, data_stage_4__452_, data_stage_4__451_, data_stage_4__450_, data_stage_4__449_, data_stage_4__448_, data_stage_4__447_, data_stage_4__446_, data_stage_4__445_, data_stage_4__444_, data_stage_4__443_, data_stage_4__442_, data_stage_4__441_, data_stage_4__440_, data_stage_4__439_, data_stage_4__438_, data_stage_4__437_, data_stage_4__436_, data_stage_4__435_, data_stage_4__434_, data_stage_4__433_, data_stage_4__432_, data_stage_4__431_, data_stage_4__430_, data_stage_4__429_, data_stage_4__428_, data_stage_4__427_, data_stage_4__426_, data_stage_4__425_, data_stage_4__424_, data_stage_4__423_, data_stage_4__422_, data_stage_4__421_, data_stage_4__420_, data_stage_4__419_, data_stage_4__418_, data_stage_4__417_, data_stage_4__416_, data_stage_4__415_, data_stage_4__414_, data_stage_4__413_, data_stage_4__412_, data_stage_4__411_, data_stage_4__410_, data_stage_4__409_, data_stage_4__408_, data_stage_4__407_, data_stage_4__406_, data_stage_4__405_, data_stage_4__404_, data_stage_4__403_, data_stage_4__402_, data_stage_4__401_, data_stage_4__400_, data_stage_4__399_, data_stage_4__398_, data_stage_4__397_, data_stage_4__396_, data_stage_4__395_, data_stage_4__394_, data_stage_4__393_, data_stage_4__392_, data_stage_4__391_, data_stage_4__390_, data_stage_4__389_, data_stage_4__388_, data_stage_4__387_, data_stage_4__386_, data_stage_4__385_, data_stage_4__384_, data_stage_4__383_, data_stage_4__382_, data_stage_4__381_, data_stage_4__380_, data_stage_4__379_, data_stage_4__378_, data_stage_4__377_, data_stage_4__376_, data_stage_4__375_, data_stage_4__374_, data_stage_4__373_, data_stage_4__372_, data_stage_4__371_, data_stage_4__370_, data_stage_4__369_, data_stage_4__368_, data_stage_4__367_, data_stage_4__366_, data_stage_4__365_, data_stage_4__364_, data_stage_4__363_, data_stage_4__362_, data_stage_4__361_, data_stage_4__360_, data_stage_4__359_, data_stage_4__358_, data_stage_4__357_, data_stage_4__356_, data_stage_4__355_, data_stage_4__354_, data_stage_4__353_, data_stage_4__352_, data_stage_4__351_, data_stage_4__350_, data_stage_4__349_, data_stage_4__348_, data_stage_4__347_, data_stage_4__346_, data_stage_4__345_, data_stage_4__344_, data_stage_4__343_, data_stage_4__342_, data_stage_4__341_, data_stage_4__340_, data_stage_4__339_, data_stage_4__338_, data_stage_4__337_, data_stage_4__336_, data_stage_4__335_, data_stage_4__334_, data_stage_4__333_, data_stage_4__332_, data_stage_4__331_, data_stage_4__330_, data_stage_4__329_, data_stage_4__328_, data_stage_4__327_, data_stage_4__326_, data_stage_4__325_, data_stage_4__324_, data_stage_4__323_, data_stage_4__322_, data_stage_4__321_, data_stage_4__320_, data_stage_4__319_, data_stage_4__318_, data_stage_4__317_, data_stage_4__316_, data_stage_4__315_, data_stage_4__314_, data_stage_4__313_, data_stage_4__312_, data_stage_4__311_, data_stage_4__310_, data_stage_4__309_, data_stage_4__308_, data_stage_4__307_, data_stage_4__306_, data_stage_4__305_, data_stage_4__304_, data_stage_4__303_, data_stage_4__302_, data_stage_4__301_, data_stage_4__300_, data_stage_4__299_, data_stage_4__298_, data_stage_4__297_, data_stage_4__296_, data_stage_4__295_, data_stage_4__294_, data_stage_4__293_, data_stage_4__292_, data_stage_4__291_, data_stage_4__290_, data_stage_4__289_, data_stage_4__288_, data_stage_4__287_, data_stage_4__286_, data_stage_4__285_, data_stage_4__284_, data_stage_4__283_, data_stage_4__282_, data_stage_4__281_, data_stage_4__280_, data_stage_4__279_, data_stage_4__278_, data_stage_4__277_, data_stage_4__276_, data_stage_4__275_, data_stage_4__274_, data_stage_4__273_, data_stage_4__272_, data_stage_4__271_, data_stage_4__270_, data_stage_4__269_, data_stage_4__268_, data_stage_4__267_, data_stage_4__266_, data_stage_4__265_, data_stage_4__264_, data_stage_4__263_, data_stage_4__262_, data_stage_4__261_, data_stage_4__260_, data_stage_4__259_, data_stage_4__258_, data_stage_4__257_, data_stage_4__256_, data_stage_4__255_, data_stage_4__254_, data_stage_4__253_, data_stage_4__252_, data_stage_4__251_, data_stage_4__250_, data_stage_4__249_, data_stage_4__248_, data_stage_4__247_, data_stage_4__246_, data_stage_4__245_, data_stage_4__244_, data_stage_4__243_, data_stage_4__242_, data_stage_4__241_, data_stage_4__240_, data_stage_4__239_, data_stage_4__238_, data_stage_4__237_, data_stage_4__236_, data_stage_4__235_, data_stage_4__234_, data_stage_4__233_, data_stage_4__232_, data_stage_4__231_, data_stage_4__230_, data_stage_4__229_, data_stage_4__228_, data_stage_4__227_, data_stage_4__226_, data_stage_4__225_, data_stage_4__224_, data_stage_4__223_, data_stage_4__222_, data_stage_4__221_, data_stage_4__220_, data_stage_4__219_, data_stage_4__218_, data_stage_4__217_, data_stage_4__216_, data_stage_4__215_, data_stage_4__214_, data_stage_4__213_, data_stage_4__212_, data_stage_4__211_, data_stage_4__210_, data_stage_4__209_, data_stage_4__208_, data_stage_4__207_, data_stage_4__206_, data_stage_4__205_, data_stage_4__204_, data_stage_4__203_, data_stage_4__202_, data_stage_4__201_, data_stage_4__200_, data_stage_4__199_, data_stage_4__198_, data_stage_4__197_, data_stage_4__196_, data_stage_4__195_, data_stage_4__194_, data_stage_4__193_, data_stage_4__192_, data_stage_4__191_, data_stage_4__190_, data_stage_4__189_, data_stage_4__188_, data_stage_4__187_, data_stage_4__186_, data_stage_4__185_, data_stage_4__184_, data_stage_4__183_, data_stage_4__182_, data_stage_4__181_, data_stage_4__180_, data_stage_4__179_, data_stage_4__178_, data_stage_4__177_, data_stage_4__176_, data_stage_4__175_, data_stage_4__174_, data_stage_4__173_, data_stage_4__172_, data_stage_4__171_, data_stage_4__170_, data_stage_4__169_, data_stage_4__168_, data_stage_4__167_, data_stage_4__166_, data_stage_4__165_, data_stage_4__164_, data_stage_4__163_, data_stage_4__162_, data_stage_4__161_, data_stage_4__160_, data_stage_4__159_, data_stage_4__158_, data_stage_4__157_, data_stage_4__156_, data_stage_4__155_, data_stage_4__154_, data_stage_4__153_, data_stage_4__152_, data_stage_4__151_, data_stage_4__150_, data_stage_4__149_, data_stage_4__148_, data_stage_4__147_, data_stage_4__146_, data_stage_4__145_, data_stage_4__144_, data_stage_4__143_, data_stage_4__142_, data_stage_4__141_, data_stage_4__140_, data_stage_4__139_, data_stage_4__138_, data_stage_4__137_, data_stage_4__136_, data_stage_4__135_, data_stage_4__134_, data_stage_4__133_, data_stage_4__132_, data_stage_4__131_, data_stage_4__130_, data_stage_4__129_, data_stage_4__128_, data_stage_4__127_, data_stage_4__126_, data_stage_4__125_, data_stage_4__124_, data_stage_4__123_, data_stage_4__122_, data_stage_4__121_, data_stage_4__120_, data_stage_4__119_, data_stage_4__118_, data_stage_4__117_, data_stage_4__116_, data_stage_4__115_, data_stage_4__114_, data_stage_4__113_, data_stage_4__112_, data_stage_4__111_, data_stage_4__110_, data_stage_4__109_, data_stage_4__108_, data_stage_4__107_, data_stage_4__106_, data_stage_4__105_, data_stage_4__104_, data_stage_4__103_, data_stage_4__102_, data_stage_4__101_, data_stage_4__100_, data_stage_4__99_, data_stage_4__98_, data_stage_4__97_, data_stage_4__96_, data_stage_4__95_, data_stage_4__94_, data_stage_4__93_, data_stage_4__92_, data_stage_4__91_, data_stage_4__90_, data_stage_4__89_, data_stage_4__88_, data_stage_4__87_, data_stage_4__86_, data_stage_4__85_, data_stage_4__84_, data_stage_4__83_, data_stage_4__82_, data_stage_4__81_, data_stage_4__80_, data_stage_4__79_, data_stage_4__78_, data_stage_4__77_, data_stage_4__76_, data_stage_4__75_, data_stage_4__74_, data_stage_4__73_, data_stage_4__72_, data_stage_4__71_, data_stage_4__70_, data_stage_4__69_, data_stage_4__68_, data_stage_4__67_, data_stage_4__66_, data_stage_4__65_, data_stage_4__64_, data_stage_4__63_, data_stage_4__62_, data_stage_4__61_, data_stage_4__60_, data_stage_4__59_, data_stage_4__58_, data_stage_4__57_, data_stage_4__56_, data_stage_4__55_, data_stage_4__54_, data_stage_4__53_, data_stage_4__52_, data_stage_4__51_, data_stage_4__50_, data_stage_4__49_, data_stage_4__48_, data_stage_4__47_, data_stage_4__46_, data_stage_4__45_, data_stage_4__44_, data_stage_4__43_, data_stage_4__42_, data_stage_4__41_, data_stage_4__40_, data_stage_4__39_, data_stage_4__38_, data_stage_4__37_, data_stage_4__36_, data_stage_4__35_, data_stage_4__34_, data_stage_4__33_, data_stage_4__32_, data_stage_4__31_, data_stage_4__30_, data_stage_4__29_, data_stage_4__28_, data_stage_4__27_, data_stage_4__26_, data_stage_4__25_, data_stage_4__24_, data_stage_4__23_, data_stage_4__22_, data_stage_4__21_, data_stage_4__20_, data_stage_4__19_, data_stage_4__18_, data_stage_4__17_, data_stage_4__16_, data_stage_4__15_, data_stage_4__14_, data_stage_4__13_, data_stage_4__12_, data_stage_4__11_, data_stage_4__10_, data_stage_4__9_, data_stage_4__8_, data_stage_4__7_, data_stage_4__6_, data_stage_4__5_, data_stage_4__4_, data_stage_4__3_, data_stage_4__2_, data_stage_4__1_, data_stage_4__0_ }),
    .swap_i(sel_i[4]),
    .data_o({ data_stage_5__4095_, data_stage_5__4094_, data_stage_5__4093_, data_stage_5__4092_, data_stage_5__4091_, data_stage_5__4090_, data_stage_5__4089_, data_stage_5__4088_, data_stage_5__4087_, data_stage_5__4086_, data_stage_5__4085_, data_stage_5__4084_, data_stage_5__4083_, data_stage_5__4082_, data_stage_5__4081_, data_stage_5__4080_, data_stage_5__4079_, data_stage_5__4078_, data_stage_5__4077_, data_stage_5__4076_, data_stage_5__4075_, data_stage_5__4074_, data_stage_5__4073_, data_stage_5__4072_, data_stage_5__4071_, data_stage_5__4070_, data_stage_5__4069_, data_stage_5__4068_, data_stage_5__4067_, data_stage_5__4066_, data_stage_5__4065_, data_stage_5__4064_, data_stage_5__4063_, data_stage_5__4062_, data_stage_5__4061_, data_stage_5__4060_, data_stage_5__4059_, data_stage_5__4058_, data_stage_5__4057_, data_stage_5__4056_, data_stage_5__4055_, data_stage_5__4054_, data_stage_5__4053_, data_stage_5__4052_, data_stage_5__4051_, data_stage_5__4050_, data_stage_5__4049_, data_stage_5__4048_, data_stage_5__4047_, data_stage_5__4046_, data_stage_5__4045_, data_stage_5__4044_, data_stage_5__4043_, data_stage_5__4042_, data_stage_5__4041_, data_stage_5__4040_, data_stage_5__4039_, data_stage_5__4038_, data_stage_5__4037_, data_stage_5__4036_, data_stage_5__4035_, data_stage_5__4034_, data_stage_5__4033_, data_stage_5__4032_, data_stage_5__4031_, data_stage_5__4030_, data_stage_5__4029_, data_stage_5__4028_, data_stage_5__4027_, data_stage_5__4026_, data_stage_5__4025_, data_stage_5__4024_, data_stage_5__4023_, data_stage_5__4022_, data_stage_5__4021_, data_stage_5__4020_, data_stage_5__4019_, data_stage_5__4018_, data_stage_5__4017_, data_stage_5__4016_, data_stage_5__4015_, data_stage_5__4014_, data_stage_5__4013_, data_stage_5__4012_, data_stage_5__4011_, data_stage_5__4010_, data_stage_5__4009_, data_stage_5__4008_, data_stage_5__4007_, data_stage_5__4006_, data_stage_5__4005_, data_stage_5__4004_, data_stage_5__4003_, data_stage_5__4002_, data_stage_5__4001_, data_stage_5__4000_, data_stage_5__3999_, data_stage_5__3998_, data_stage_5__3997_, data_stage_5__3996_, data_stage_5__3995_, data_stage_5__3994_, data_stage_5__3993_, data_stage_5__3992_, data_stage_5__3991_, data_stage_5__3990_, data_stage_5__3989_, data_stage_5__3988_, data_stage_5__3987_, data_stage_5__3986_, data_stage_5__3985_, data_stage_5__3984_, data_stage_5__3983_, data_stage_5__3982_, data_stage_5__3981_, data_stage_5__3980_, data_stage_5__3979_, data_stage_5__3978_, data_stage_5__3977_, data_stage_5__3976_, data_stage_5__3975_, data_stage_5__3974_, data_stage_5__3973_, data_stage_5__3972_, data_stage_5__3971_, data_stage_5__3970_, data_stage_5__3969_, data_stage_5__3968_, data_stage_5__3967_, data_stage_5__3966_, data_stage_5__3965_, data_stage_5__3964_, data_stage_5__3963_, data_stage_5__3962_, data_stage_5__3961_, data_stage_5__3960_, data_stage_5__3959_, data_stage_5__3958_, data_stage_5__3957_, data_stage_5__3956_, data_stage_5__3955_, data_stage_5__3954_, data_stage_5__3953_, data_stage_5__3952_, data_stage_5__3951_, data_stage_5__3950_, data_stage_5__3949_, data_stage_5__3948_, data_stage_5__3947_, data_stage_5__3946_, data_stage_5__3945_, data_stage_5__3944_, data_stage_5__3943_, data_stage_5__3942_, data_stage_5__3941_, data_stage_5__3940_, data_stage_5__3939_, data_stage_5__3938_, data_stage_5__3937_, data_stage_5__3936_, data_stage_5__3935_, data_stage_5__3934_, data_stage_5__3933_, data_stage_5__3932_, data_stage_5__3931_, data_stage_5__3930_, data_stage_5__3929_, data_stage_5__3928_, data_stage_5__3927_, data_stage_5__3926_, data_stage_5__3925_, data_stage_5__3924_, data_stage_5__3923_, data_stage_5__3922_, data_stage_5__3921_, data_stage_5__3920_, data_stage_5__3919_, data_stage_5__3918_, data_stage_5__3917_, data_stage_5__3916_, data_stage_5__3915_, data_stage_5__3914_, data_stage_5__3913_, data_stage_5__3912_, data_stage_5__3911_, data_stage_5__3910_, data_stage_5__3909_, data_stage_5__3908_, data_stage_5__3907_, data_stage_5__3906_, data_stage_5__3905_, data_stage_5__3904_, data_stage_5__3903_, data_stage_5__3902_, data_stage_5__3901_, data_stage_5__3900_, data_stage_5__3899_, data_stage_5__3898_, data_stage_5__3897_, data_stage_5__3896_, data_stage_5__3895_, data_stage_5__3894_, data_stage_5__3893_, data_stage_5__3892_, data_stage_5__3891_, data_stage_5__3890_, data_stage_5__3889_, data_stage_5__3888_, data_stage_5__3887_, data_stage_5__3886_, data_stage_5__3885_, data_stage_5__3884_, data_stage_5__3883_, data_stage_5__3882_, data_stage_5__3881_, data_stage_5__3880_, data_stage_5__3879_, data_stage_5__3878_, data_stage_5__3877_, data_stage_5__3876_, data_stage_5__3875_, data_stage_5__3874_, data_stage_5__3873_, data_stage_5__3872_, data_stage_5__3871_, data_stage_5__3870_, data_stage_5__3869_, data_stage_5__3868_, data_stage_5__3867_, data_stage_5__3866_, data_stage_5__3865_, data_stage_5__3864_, data_stage_5__3863_, data_stage_5__3862_, data_stage_5__3861_, data_stage_5__3860_, data_stage_5__3859_, data_stage_5__3858_, data_stage_5__3857_, data_stage_5__3856_, data_stage_5__3855_, data_stage_5__3854_, data_stage_5__3853_, data_stage_5__3852_, data_stage_5__3851_, data_stage_5__3850_, data_stage_5__3849_, data_stage_5__3848_, data_stage_5__3847_, data_stage_5__3846_, data_stage_5__3845_, data_stage_5__3844_, data_stage_5__3843_, data_stage_5__3842_, data_stage_5__3841_, data_stage_5__3840_, data_stage_5__3839_, data_stage_5__3838_, data_stage_5__3837_, data_stage_5__3836_, data_stage_5__3835_, data_stage_5__3834_, data_stage_5__3833_, data_stage_5__3832_, data_stage_5__3831_, data_stage_5__3830_, data_stage_5__3829_, data_stage_5__3828_, data_stage_5__3827_, data_stage_5__3826_, data_stage_5__3825_, data_stage_5__3824_, data_stage_5__3823_, data_stage_5__3822_, data_stage_5__3821_, data_stage_5__3820_, data_stage_5__3819_, data_stage_5__3818_, data_stage_5__3817_, data_stage_5__3816_, data_stage_5__3815_, data_stage_5__3814_, data_stage_5__3813_, data_stage_5__3812_, data_stage_5__3811_, data_stage_5__3810_, data_stage_5__3809_, data_stage_5__3808_, data_stage_5__3807_, data_stage_5__3806_, data_stage_5__3805_, data_stage_5__3804_, data_stage_5__3803_, data_stage_5__3802_, data_stage_5__3801_, data_stage_5__3800_, data_stage_5__3799_, data_stage_5__3798_, data_stage_5__3797_, data_stage_5__3796_, data_stage_5__3795_, data_stage_5__3794_, data_stage_5__3793_, data_stage_5__3792_, data_stage_5__3791_, data_stage_5__3790_, data_stage_5__3789_, data_stage_5__3788_, data_stage_5__3787_, data_stage_5__3786_, data_stage_5__3785_, data_stage_5__3784_, data_stage_5__3783_, data_stage_5__3782_, data_stage_5__3781_, data_stage_5__3780_, data_stage_5__3779_, data_stage_5__3778_, data_stage_5__3777_, data_stage_5__3776_, data_stage_5__3775_, data_stage_5__3774_, data_stage_5__3773_, data_stage_5__3772_, data_stage_5__3771_, data_stage_5__3770_, data_stage_5__3769_, data_stage_5__3768_, data_stage_5__3767_, data_stage_5__3766_, data_stage_5__3765_, data_stage_5__3764_, data_stage_5__3763_, data_stage_5__3762_, data_stage_5__3761_, data_stage_5__3760_, data_stage_5__3759_, data_stage_5__3758_, data_stage_5__3757_, data_stage_5__3756_, data_stage_5__3755_, data_stage_5__3754_, data_stage_5__3753_, data_stage_5__3752_, data_stage_5__3751_, data_stage_5__3750_, data_stage_5__3749_, data_stage_5__3748_, data_stage_5__3747_, data_stage_5__3746_, data_stage_5__3745_, data_stage_5__3744_, data_stage_5__3743_, data_stage_5__3742_, data_stage_5__3741_, data_stage_5__3740_, data_stage_5__3739_, data_stage_5__3738_, data_stage_5__3737_, data_stage_5__3736_, data_stage_5__3735_, data_stage_5__3734_, data_stage_5__3733_, data_stage_5__3732_, data_stage_5__3731_, data_stage_5__3730_, data_stage_5__3729_, data_stage_5__3728_, data_stage_5__3727_, data_stage_5__3726_, data_stage_5__3725_, data_stage_5__3724_, data_stage_5__3723_, data_stage_5__3722_, data_stage_5__3721_, data_stage_5__3720_, data_stage_5__3719_, data_stage_5__3718_, data_stage_5__3717_, data_stage_5__3716_, data_stage_5__3715_, data_stage_5__3714_, data_stage_5__3713_, data_stage_5__3712_, data_stage_5__3711_, data_stage_5__3710_, data_stage_5__3709_, data_stage_5__3708_, data_stage_5__3707_, data_stage_5__3706_, data_stage_5__3705_, data_stage_5__3704_, data_stage_5__3703_, data_stage_5__3702_, data_stage_5__3701_, data_stage_5__3700_, data_stage_5__3699_, data_stage_5__3698_, data_stage_5__3697_, data_stage_5__3696_, data_stage_5__3695_, data_stage_5__3694_, data_stage_5__3693_, data_stage_5__3692_, data_stage_5__3691_, data_stage_5__3690_, data_stage_5__3689_, data_stage_5__3688_, data_stage_5__3687_, data_stage_5__3686_, data_stage_5__3685_, data_stage_5__3684_, data_stage_5__3683_, data_stage_5__3682_, data_stage_5__3681_, data_stage_5__3680_, data_stage_5__3679_, data_stage_5__3678_, data_stage_5__3677_, data_stage_5__3676_, data_stage_5__3675_, data_stage_5__3674_, data_stage_5__3673_, data_stage_5__3672_, data_stage_5__3671_, data_stage_5__3670_, data_stage_5__3669_, data_stage_5__3668_, data_stage_5__3667_, data_stage_5__3666_, data_stage_5__3665_, data_stage_5__3664_, data_stage_5__3663_, data_stage_5__3662_, data_stage_5__3661_, data_stage_5__3660_, data_stage_5__3659_, data_stage_5__3658_, data_stage_5__3657_, data_stage_5__3656_, data_stage_5__3655_, data_stage_5__3654_, data_stage_5__3653_, data_stage_5__3652_, data_stage_5__3651_, data_stage_5__3650_, data_stage_5__3649_, data_stage_5__3648_, data_stage_5__3647_, data_stage_5__3646_, data_stage_5__3645_, data_stage_5__3644_, data_stage_5__3643_, data_stage_5__3642_, data_stage_5__3641_, data_stage_5__3640_, data_stage_5__3639_, data_stage_5__3638_, data_stage_5__3637_, data_stage_5__3636_, data_stage_5__3635_, data_stage_5__3634_, data_stage_5__3633_, data_stage_5__3632_, data_stage_5__3631_, data_stage_5__3630_, data_stage_5__3629_, data_stage_5__3628_, data_stage_5__3627_, data_stage_5__3626_, data_stage_5__3625_, data_stage_5__3624_, data_stage_5__3623_, data_stage_5__3622_, data_stage_5__3621_, data_stage_5__3620_, data_stage_5__3619_, data_stage_5__3618_, data_stage_5__3617_, data_stage_5__3616_, data_stage_5__3615_, data_stage_5__3614_, data_stage_5__3613_, data_stage_5__3612_, data_stage_5__3611_, data_stage_5__3610_, data_stage_5__3609_, data_stage_5__3608_, data_stage_5__3607_, data_stage_5__3606_, data_stage_5__3605_, data_stage_5__3604_, data_stage_5__3603_, data_stage_5__3602_, data_stage_5__3601_, data_stage_5__3600_, data_stage_5__3599_, data_stage_5__3598_, data_stage_5__3597_, data_stage_5__3596_, data_stage_5__3595_, data_stage_5__3594_, data_stage_5__3593_, data_stage_5__3592_, data_stage_5__3591_, data_stage_5__3590_, data_stage_5__3589_, data_stage_5__3588_, data_stage_5__3587_, data_stage_5__3586_, data_stage_5__3585_, data_stage_5__3584_, data_stage_5__3583_, data_stage_5__3582_, data_stage_5__3581_, data_stage_5__3580_, data_stage_5__3579_, data_stage_5__3578_, data_stage_5__3577_, data_stage_5__3576_, data_stage_5__3575_, data_stage_5__3574_, data_stage_5__3573_, data_stage_5__3572_, data_stage_5__3571_, data_stage_5__3570_, data_stage_5__3569_, data_stage_5__3568_, data_stage_5__3567_, data_stage_5__3566_, data_stage_5__3565_, data_stage_5__3564_, data_stage_5__3563_, data_stage_5__3562_, data_stage_5__3561_, data_stage_5__3560_, data_stage_5__3559_, data_stage_5__3558_, data_stage_5__3557_, data_stage_5__3556_, data_stage_5__3555_, data_stage_5__3554_, data_stage_5__3553_, data_stage_5__3552_, data_stage_5__3551_, data_stage_5__3550_, data_stage_5__3549_, data_stage_5__3548_, data_stage_5__3547_, data_stage_5__3546_, data_stage_5__3545_, data_stage_5__3544_, data_stage_5__3543_, data_stage_5__3542_, data_stage_5__3541_, data_stage_5__3540_, data_stage_5__3539_, data_stage_5__3538_, data_stage_5__3537_, data_stage_5__3536_, data_stage_5__3535_, data_stage_5__3534_, data_stage_5__3533_, data_stage_5__3532_, data_stage_5__3531_, data_stage_5__3530_, data_stage_5__3529_, data_stage_5__3528_, data_stage_5__3527_, data_stage_5__3526_, data_stage_5__3525_, data_stage_5__3524_, data_stage_5__3523_, data_stage_5__3522_, data_stage_5__3521_, data_stage_5__3520_, data_stage_5__3519_, data_stage_5__3518_, data_stage_5__3517_, data_stage_5__3516_, data_stage_5__3515_, data_stage_5__3514_, data_stage_5__3513_, data_stage_5__3512_, data_stage_5__3511_, data_stage_5__3510_, data_stage_5__3509_, data_stage_5__3508_, data_stage_5__3507_, data_stage_5__3506_, data_stage_5__3505_, data_stage_5__3504_, data_stage_5__3503_, data_stage_5__3502_, data_stage_5__3501_, data_stage_5__3500_, data_stage_5__3499_, data_stage_5__3498_, data_stage_5__3497_, data_stage_5__3496_, data_stage_5__3495_, data_stage_5__3494_, data_stage_5__3493_, data_stage_5__3492_, data_stage_5__3491_, data_stage_5__3490_, data_stage_5__3489_, data_stage_5__3488_, data_stage_5__3487_, data_stage_5__3486_, data_stage_5__3485_, data_stage_5__3484_, data_stage_5__3483_, data_stage_5__3482_, data_stage_5__3481_, data_stage_5__3480_, data_stage_5__3479_, data_stage_5__3478_, data_stage_5__3477_, data_stage_5__3476_, data_stage_5__3475_, data_stage_5__3474_, data_stage_5__3473_, data_stage_5__3472_, data_stage_5__3471_, data_stage_5__3470_, data_stage_5__3469_, data_stage_5__3468_, data_stage_5__3467_, data_stage_5__3466_, data_stage_5__3465_, data_stage_5__3464_, data_stage_5__3463_, data_stage_5__3462_, data_stage_5__3461_, data_stage_5__3460_, data_stage_5__3459_, data_stage_5__3458_, data_stage_5__3457_, data_stage_5__3456_, data_stage_5__3455_, data_stage_5__3454_, data_stage_5__3453_, data_stage_5__3452_, data_stage_5__3451_, data_stage_5__3450_, data_stage_5__3449_, data_stage_5__3448_, data_stage_5__3447_, data_stage_5__3446_, data_stage_5__3445_, data_stage_5__3444_, data_stage_5__3443_, data_stage_5__3442_, data_stage_5__3441_, data_stage_5__3440_, data_stage_5__3439_, data_stage_5__3438_, data_stage_5__3437_, data_stage_5__3436_, data_stage_5__3435_, data_stage_5__3434_, data_stage_5__3433_, data_stage_5__3432_, data_stage_5__3431_, data_stage_5__3430_, data_stage_5__3429_, data_stage_5__3428_, data_stage_5__3427_, data_stage_5__3426_, data_stage_5__3425_, data_stage_5__3424_, data_stage_5__3423_, data_stage_5__3422_, data_stage_5__3421_, data_stage_5__3420_, data_stage_5__3419_, data_stage_5__3418_, data_stage_5__3417_, data_stage_5__3416_, data_stage_5__3415_, data_stage_5__3414_, data_stage_5__3413_, data_stage_5__3412_, data_stage_5__3411_, data_stage_5__3410_, data_stage_5__3409_, data_stage_5__3408_, data_stage_5__3407_, data_stage_5__3406_, data_stage_5__3405_, data_stage_5__3404_, data_stage_5__3403_, data_stage_5__3402_, data_stage_5__3401_, data_stage_5__3400_, data_stage_5__3399_, data_stage_5__3398_, data_stage_5__3397_, data_stage_5__3396_, data_stage_5__3395_, data_stage_5__3394_, data_stage_5__3393_, data_stage_5__3392_, data_stage_5__3391_, data_stage_5__3390_, data_stage_5__3389_, data_stage_5__3388_, data_stage_5__3387_, data_stage_5__3386_, data_stage_5__3385_, data_stage_5__3384_, data_stage_5__3383_, data_stage_5__3382_, data_stage_5__3381_, data_stage_5__3380_, data_stage_5__3379_, data_stage_5__3378_, data_stage_5__3377_, data_stage_5__3376_, data_stage_5__3375_, data_stage_5__3374_, data_stage_5__3373_, data_stage_5__3372_, data_stage_5__3371_, data_stage_5__3370_, data_stage_5__3369_, data_stage_5__3368_, data_stage_5__3367_, data_stage_5__3366_, data_stage_5__3365_, data_stage_5__3364_, data_stage_5__3363_, data_stage_5__3362_, data_stage_5__3361_, data_stage_5__3360_, data_stage_5__3359_, data_stage_5__3358_, data_stage_5__3357_, data_stage_5__3356_, data_stage_5__3355_, data_stage_5__3354_, data_stage_5__3353_, data_stage_5__3352_, data_stage_5__3351_, data_stage_5__3350_, data_stage_5__3349_, data_stage_5__3348_, data_stage_5__3347_, data_stage_5__3346_, data_stage_5__3345_, data_stage_5__3344_, data_stage_5__3343_, data_stage_5__3342_, data_stage_5__3341_, data_stage_5__3340_, data_stage_5__3339_, data_stage_5__3338_, data_stage_5__3337_, data_stage_5__3336_, data_stage_5__3335_, data_stage_5__3334_, data_stage_5__3333_, data_stage_5__3332_, data_stage_5__3331_, data_stage_5__3330_, data_stage_5__3329_, data_stage_5__3328_, data_stage_5__3327_, data_stage_5__3326_, data_stage_5__3325_, data_stage_5__3324_, data_stage_5__3323_, data_stage_5__3322_, data_stage_5__3321_, data_stage_5__3320_, data_stage_5__3319_, data_stage_5__3318_, data_stage_5__3317_, data_stage_5__3316_, data_stage_5__3315_, data_stage_5__3314_, data_stage_5__3313_, data_stage_5__3312_, data_stage_5__3311_, data_stage_5__3310_, data_stage_5__3309_, data_stage_5__3308_, data_stage_5__3307_, data_stage_5__3306_, data_stage_5__3305_, data_stage_5__3304_, data_stage_5__3303_, data_stage_5__3302_, data_stage_5__3301_, data_stage_5__3300_, data_stage_5__3299_, data_stage_5__3298_, data_stage_5__3297_, data_stage_5__3296_, data_stage_5__3295_, data_stage_5__3294_, data_stage_5__3293_, data_stage_5__3292_, data_stage_5__3291_, data_stage_5__3290_, data_stage_5__3289_, data_stage_5__3288_, data_stage_5__3287_, data_stage_5__3286_, data_stage_5__3285_, data_stage_5__3284_, data_stage_5__3283_, data_stage_5__3282_, data_stage_5__3281_, data_stage_5__3280_, data_stage_5__3279_, data_stage_5__3278_, data_stage_5__3277_, data_stage_5__3276_, data_stage_5__3275_, data_stage_5__3274_, data_stage_5__3273_, data_stage_5__3272_, data_stage_5__3271_, data_stage_5__3270_, data_stage_5__3269_, data_stage_5__3268_, data_stage_5__3267_, data_stage_5__3266_, data_stage_5__3265_, data_stage_5__3264_, data_stage_5__3263_, data_stage_5__3262_, data_stage_5__3261_, data_stage_5__3260_, data_stage_5__3259_, data_stage_5__3258_, data_stage_5__3257_, data_stage_5__3256_, data_stage_5__3255_, data_stage_5__3254_, data_stage_5__3253_, data_stage_5__3252_, data_stage_5__3251_, data_stage_5__3250_, data_stage_5__3249_, data_stage_5__3248_, data_stage_5__3247_, data_stage_5__3246_, data_stage_5__3245_, data_stage_5__3244_, data_stage_5__3243_, data_stage_5__3242_, data_stage_5__3241_, data_stage_5__3240_, data_stage_5__3239_, data_stage_5__3238_, data_stage_5__3237_, data_stage_5__3236_, data_stage_5__3235_, data_stage_5__3234_, data_stage_5__3233_, data_stage_5__3232_, data_stage_5__3231_, data_stage_5__3230_, data_stage_5__3229_, data_stage_5__3228_, data_stage_5__3227_, data_stage_5__3226_, data_stage_5__3225_, data_stage_5__3224_, data_stage_5__3223_, data_stage_5__3222_, data_stage_5__3221_, data_stage_5__3220_, data_stage_5__3219_, data_stage_5__3218_, data_stage_5__3217_, data_stage_5__3216_, data_stage_5__3215_, data_stage_5__3214_, data_stage_5__3213_, data_stage_5__3212_, data_stage_5__3211_, data_stage_5__3210_, data_stage_5__3209_, data_stage_5__3208_, data_stage_5__3207_, data_stage_5__3206_, data_stage_5__3205_, data_stage_5__3204_, data_stage_5__3203_, data_stage_5__3202_, data_stage_5__3201_, data_stage_5__3200_, data_stage_5__3199_, data_stage_5__3198_, data_stage_5__3197_, data_stage_5__3196_, data_stage_5__3195_, data_stage_5__3194_, data_stage_5__3193_, data_stage_5__3192_, data_stage_5__3191_, data_stage_5__3190_, data_stage_5__3189_, data_stage_5__3188_, data_stage_5__3187_, data_stage_5__3186_, data_stage_5__3185_, data_stage_5__3184_, data_stage_5__3183_, data_stage_5__3182_, data_stage_5__3181_, data_stage_5__3180_, data_stage_5__3179_, data_stage_5__3178_, data_stage_5__3177_, data_stage_5__3176_, data_stage_5__3175_, data_stage_5__3174_, data_stage_5__3173_, data_stage_5__3172_, data_stage_5__3171_, data_stage_5__3170_, data_stage_5__3169_, data_stage_5__3168_, data_stage_5__3167_, data_stage_5__3166_, data_stage_5__3165_, data_stage_5__3164_, data_stage_5__3163_, data_stage_5__3162_, data_stage_5__3161_, data_stage_5__3160_, data_stage_5__3159_, data_stage_5__3158_, data_stage_5__3157_, data_stage_5__3156_, data_stage_5__3155_, data_stage_5__3154_, data_stage_5__3153_, data_stage_5__3152_, data_stage_5__3151_, data_stage_5__3150_, data_stage_5__3149_, data_stage_5__3148_, data_stage_5__3147_, data_stage_5__3146_, data_stage_5__3145_, data_stage_5__3144_, data_stage_5__3143_, data_stage_5__3142_, data_stage_5__3141_, data_stage_5__3140_, data_stage_5__3139_, data_stage_5__3138_, data_stage_5__3137_, data_stage_5__3136_, data_stage_5__3135_, data_stage_5__3134_, data_stage_5__3133_, data_stage_5__3132_, data_stage_5__3131_, data_stage_5__3130_, data_stage_5__3129_, data_stage_5__3128_, data_stage_5__3127_, data_stage_5__3126_, data_stage_5__3125_, data_stage_5__3124_, data_stage_5__3123_, data_stage_5__3122_, data_stage_5__3121_, data_stage_5__3120_, data_stage_5__3119_, data_stage_5__3118_, data_stage_5__3117_, data_stage_5__3116_, data_stage_5__3115_, data_stage_5__3114_, data_stage_5__3113_, data_stage_5__3112_, data_stage_5__3111_, data_stage_5__3110_, data_stage_5__3109_, data_stage_5__3108_, data_stage_5__3107_, data_stage_5__3106_, data_stage_5__3105_, data_stage_5__3104_, data_stage_5__3103_, data_stage_5__3102_, data_stage_5__3101_, data_stage_5__3100_, data_stage_5__3099_, data_stage_5__3098_, data_stage_5__3097_, data_stage_5__3096_, data_stage_5__3095_, data_stage_5__3094_, data_stage_5__3093_, data_stage_5__3092_, data_stage_5__3091_, data_stage_5__3090_, data_stage_5__3089_, data_stage_5__3088_, data_stage_5__3087_, data_stage_5__3086_, data_stage_5__3085_, data_stage_5__3084_, data_stage_5__3083_, data_stage_5__3082_, data_stage_5__3081_, data_stage_5__3080_, data_stage_5__3079_, data_stage_5__3078_, data_stage_5__3077_, data_stage_5__3076_, data_stage_5__3075_, data_stage_5__3074_, data_stage_5__3073_, data_stage_5__3072_, data_stage_5__3071_, data_stage_5__3070_, data_stage_5__3069_, data_stage_5__3068_, data_stage_5__3067_, data_stage_5__3066_, data_stage_5__3065_, data_stage_5__3064_, data_stage_5__3063_, data_stage_5__3062_, data_stage_5__3061_, data_stage_5__3060_, data_stage_5__3059_, data_stage_5__3058_, data_stage_5__3057_, data_stage_5__3056_, data_stage_5__3055_, data_stage_5__3054_, data_stage_5__3053_, data_stage_5__3052_, data_stage_5__3051_, data_stage_5__3050_, data_stage_5__3049_, data_stage_5__3048_, data_stage_5__3047_, data_stage_5__3046_, data_stage_5__3045_, data_stage_5__3044_, data_stage_5__3043_, data_stage_5__3042_, data_stage_5__3041_, data_stage_5__3040_, data_stage_5__3039_, data_stage_5__3038_, data_stage_5__3037_, data_stage_5__3036_, data_stage_5__3035_, data_stage_5__3034_, data_stage_5__3033_, data_stage_5__3032_, data_stage_5__3031_, data_stage_5__3030_, data_stage_5__3029_, data_stage_5__3028_, data_stage_5__3027_, data_stage_5__3026_, data_stage_5__3025_, data_stage_5__3024_, data_stage_5__3023_, data_stage_5__3022_, data_stage_5__3021_, data_stage_5__3020_, data_stage_5__3019_, data_stage_5__3018_, data_stage_5__3017_, data_stage_5__3016_, data_stage_5__3015_, data_stage_5__3014_, data_stage_5__3013_, data_stage_5__3012_, data_stage_5__3011_, data_stage_5__3010_, data_stage_5__3009_, data_stage_5__3008_, data_stage_5__3007_, data_stage_5__3006_, data_stage_5__3005_, data_stage_5__3004_, data_stage_5__3003_, data_stage_5__3002_, data_stage_5__3001_, data_stage_5__3000_, data_stage_5__2999_, data_stage_5__2998_, data_stage_5__2997_, data_stage_5__2996_, data_stage_5__2995_, data_stage_5__2994_, data_stage_5__2993_, data_stage_5__2992_, data_stage_5__2991_, data_stage_5__2990_, data_stage_5__2989_, data_stage_5__2988_, data_stage_5__2987_, data_stage_5__2986_, data_stage_5__2985_, data_stage_5__2984_, data_stage_5__2983_, data_stage_5__2982_, data_stage_5__2981_, data_stage_5__2980_, data_stage_5__2979_, data_stage_5__2978_, data_stage_5__2977_, data_stage_5__2976_, data_stage_5__2975_, data_stage_5__2974_, data_stage_5__2973_, data_stage_5__2972_, data_stage_5__2971_, data_stage_5__2970_, data_stage_5__2969_, data_stage_5__2968_, data_stage_5__2967_, data_stage_5__2966_, data_stage_5__2965_, data_stage_5__2964_, data_stage_5__2963_, data_stage_5__2962_, data_stage_5__2961_, data_stage_5__2960_, data_stage_5__2959_, data_stage_5__2958_, data_stage_5__2957_, data_stage_5__2956_, data_stage_5__2955_, data_stage_5__2954_, data_stage_5__2953_, data_stage_5__2952_, data_stage_5__2951_, data_stage_5__2950_, data_stage_5__2949_, data_stage_5__2948_, data_stage_5__2947_, data_stage_5__2946_, data_stage_5__2945_, data_stage_5__2944_, data_stage_5__2943_, data_stage_5__2942_, data_stage_5__2941_, data_stage_5__2940_, data_stage_5__2939_, data_stage_5__2938_, data_stage_5__2937_, data_stage_5__2936_, data_stage_5__2935_, data_stage_5__2934_, data_stage_5__2933_, data_stage_5__2932_, data_stage_5__2931_, data_stage_5__2930_, data_stage_5__2929_, data_stage_5__2928_, data_stage_5__2927_, data_stage_5__2926_, data_stage_5__2925_, data_stage_5__2924_, data_stage_5__2923_, data_stage_5__2922_, data_stage_5__2921_, data_stage_5__2920_, data_stage_5__2919_, data_stage_5__2918_, data_stage_5__2917_, data_stage_5__2916_, data_stage_5__2915_, data_stage_5__2914_, data_stage_5__2913_, data_stage_5__2912_, data_stage_5__2911_, data_stage_5__2910_, data_stage_5__2909_, data_stage_5__2908_, data_stage_5__2907_, data_stage_5__2906_, data_stage_5__2905_, data_stage_5__2904_, data_stage_5__2903_, data_stage_5__2902_, data_stage_5__2901_, data_stage_5__2900_, data_stage_5__2899_, data_stage_5__2898_, data_stage_5__2897_, data_stage_5__2896_, data_stage_5__2895_, data_stage_5__2894_, data_stage_5__2893_, data_stage_5__2892_, data_stage_5__2891_, data_stage_5__2890_, data_stage_5__2889_, data_stage_5__2888_, data_stage_5__2887_, data_stage_5__2886_, data_stage_5__2885_, data_stage_5__2884_, data_stage_5__2883_, data_stage_5__2882_, data_stage_5__2881_, data_stage_5__2880_, data_stage_5__2879_, data_stage_5__2878_, data_stage_5__2877_, data_stage_5__2876_, data_stage_5__2875_, data_stage_5__2874_, data_stage_5__2873_, data_stage_5__2872_, data_stage_5__2871_, data_stage_5__2870_, data_stage_5__2869_, data_stage_5__2868_, data_stage_5__2867_, data_stage_5__2866_, data_stage_5__2865_, data_stage_5__2864_, data_stage_5__2863_, data_stage_5__2862_, data_stage_5__2861_, data_stage_5__2860_, data_stage_5__2859_, data_stage_5__2858_, data_stage_5__2857_, data_stage_5__2856_, data_stage_5__2855_, data_stage_5__2854_, data_stage_5__2853_, data_stage_5__2852_, data_stage_5__2851_, data_stage_5__2850_, data_stage_5__2849_, data_stage_5__2848_, data_stage_5__2847_, data_stage_5__2846_, data_stage_5__2845_, data_stage_5__2844_, data_stage_5__2843_, data_stage_5__2842_, data_stage_5__2841_, data_stage_5__2840_, data_stage_5__2839_, data_stage_5__2838_, data_stage_5__2837_, data_stage_5__2836_, data_stage_5__2835_, data_stage_5__2834_, data_stage_5__2833_, data_stage_5__2832_, data_stage_5__2831_, data_stage_5__2830_, data_stage_5__2829_, data_stage_5__2828_, data_stage_5__2827_, data_stage_5__2826_, data_stage_5__2825_, data_stage_5__2824_, data_stage_5__2823_, data_stage_5__2822_, data_stage_5__2821_, data_stage_5__2820_, data_stage_5__2819_, data_stage_5__2818_, data_stage_5__2817_, data_stage_5__2816_, data_stage_5__2815_, data_stage_5__2814_, data_stage_5__2813_, data_stage_5__2812_, data_stage_5__2811_, data_stage_5__2810_, data_stage_5__2809_, data_stage_5__2808_, data_stage_5__2807_, data_stage_5__2806_, data_stage_5__2805_, data_stage_5__2804_, data_stage_5__2803_, data_stage_5__2802_, data_stage_5__2801_, data_stage_5__2800_, data_stage_5__2799_, data_stage_5__2798_, data_stage_5__2797_, data_stage_5__2796_, data_stage_5__2795_, data_stage_5__2794_, data_stage_5__2793_, data_stage_5__2792_, data_stage_5__2791_, data_stage_5__2790_, data_stage_5__2789_, data_stage_5__2788_, data_stage_5__2787_, data_stage_5__2786_, data_stage_5__2785_, data_stage_5__2784_, data_stage_5__2783_, data_stage_5__2782_, data_stage_5__2781_, data_stage_5__2780_, data_stage_5__2779_, data_stage_5__2778_, data_stage_5__2777_, data_stage_5__2776_, data_stage_5__2775_, data_stage_5__2774_, data_stage_5__2773_, data_stage_5__2772_, data_stage_5__2771_, data_stage_5__2770_, data_stage_5__2769_, data_stage_5__2768_, data_stage_5__2767_, data_stage_5__2766_, data_stage_5__2765_, data_stage_5__2764_, data_stage_5__2763_, data_stage_5__2762_, data_stage_5__2761_, data_stage_5__2760_, data_stage_5__2759_, data_stage_5__2758_, data_stage_5__2757_, data_stage_5__2756_, data_stage_5__2755_, data_stage_5__2754_, data_stage_5__2753_, data_stage_5__2752_, data_stage_5__2751_, data_stage_5__2750_, data_stage_5__2749_, data_stage_5__2748_, data_stage_5__2747_, data_stage_5__2746_, data_stage_5__2745_, data_stage_5__2744_, data_stage_5__2743_, data_stage_5__2742_, data_stage_5__2741_, data_stage_5__2740_, data_stage_5__2739_, data_stage_5__2738_, data_stage_5__2737_, data_stage_5__2736_, data_stage_5__2735_, data_stage_5__2734_, data_stage_5__2733_, data_stage_5__2732_, data_stage_5__2731_, data_stage_5__2730_, data_stage_5__2729_, data_stage_5__2728_, data_stage_5__2727_, data_stage_5__2726_, data_stage_5__2725_, data_stage_5__2724_, data_stage_5__2723_, data_stage_5__2722_, data_stage_5__2721_, data_stage_5__2720_, data_stage_5__2719_, data_stage_5__2718_, data_stage_5__2717_, data_stage_5__2716_, data_stage_5__2715_, data_stage_5__2714_, data_stage_5__2713_, data_stage_5__2712_, data_stage_5__2711_, data_stage_5__2710_, data_stage_5__2709_, data_stage_5__2708_, data_stage_5__2707_, data_stage_5__2706_, data_stage_5__2705_, data_stage_5__2704_, data_stage_5__2703_, data_stage_5__2702_, data_stage_5__2701_, data_stage_5__2700_, data_stage_5__2699_, data_stage_5__2698_, data_stage_5__2697_, data_stage_5__2696_, data_stage_5__2695_, data_stage_5__2694_, data_stage_5__2693_, data_stage_5__2692_, data_stage_5__2691_, data_stage_5__2690_, data_stage_5__2689_, data_stage_5__2688_, data_stage_5__2687_, data_stage_5__2686_, data_stage_5__2685_, data_stage_5__2684_, data_stage_5__2683_, data_stage_5__2682_, data_stage_5__2681_, data_stage_5__2680_, data_stage_5__2679_, data_stage_5__2678_, data_stage_5__2677_, data_stage_5__2676_, data_stage_5__2675_, data_stage_5__2674_, data_stage_5__2673_, data_stage_5__2672_, data_stage_5__2671_, data_stage_5__2670_, data_stage_5__2669_, data_stage_5__2668_, data_stage_5__2667_, data_stage_5__2666_, data_stage_5__2665_, data_stage_5__2664_, data_stage_5__2663_, data_stage_5__2662_, data_stage_5__2661_, data_stage_5__2660_, data_stage_5__2659_, data_stage_5__2658_, data_stage_5__2657_, data_stage_5__2656_, data_stage_5__2655_, data_stage_5__2654_, data_stage_5__2653_, data_stage_5__2652_, data_stage_5__2651_, data_stage_5__2650_, data_stage_5__2649_, data_stage_5__2648_, data_stage_5__2647_, data_stage_5__2646_, data_stage_5__2645_, data_stage_5__2644_, data_stage_5__2643_, data_stage_5__2642_, data_stage_5__2641_, data_stage_5__2640_, data_stage_5__2639_, data_stage_5__2638_, data_stage_5__2637_, data_stage_5__2636_, data_stage_5__2635_, data_stage_5__2634_, data_stage_5__2633_, data_stage_5__2632_, data_stage_5__2631_, data_stage_5__2630_, data_stage_5__2629_, data_stage_5__2628_, data_stage_5__2627_, data_stage_5__2626_, data_stage_5__2625_, data_stage_5__2624_, data_stage_5__2623_, data_stage_5__2622_, data_stage_5__2621_, data_stage_5__2620_, data_stage_5__2619_, data_stage_5__2618_, data_stage_5__2617_, data_stage_5__2616_, data_stage_5__2615_, data_stage_5__2614_, data_stage_5__2613_, data_stage_5__2612_, data_stage_5__2611_, data_stage_5__2610_, data_stage_5__2609_, data_stage_5__2608_, data_stage_5__2607_, data_stage_5__2606_, data_stage_5__2605_, data_stage_5__2604_, data_stage_5__2603_, data_stage_5__2602_, data_stage_5__2601_, data_stage_5__2600_, data_stage_5__2599_, data_stage_5__2598_, data_stage_5__2597_, data_stage_5__2596_, data_stage_5__2595_, data_stage_5__2594_, data_stage_5__2593_, data_stage_5__2592_, data_stage_5__2591_, data_stage_5__2590_, data_stage_5__2589_, data_stage_5__2588_, data_stage_5__2587_, data_stage_5__2586_, data_stage_5__2585_, data_stage_5__2584_, data_stage_5__2583_, data_stage_5__2582_, data_stage_5__2581_, data_stage_5__2580_, data_stage_5__2579_, data_stage_5__2578_, data_stage_5__2577_, data_stage_5__2576_, data_stage_5__2575_, data_stage_5__2574_, data_stage_5__2573_, data_stage_5__2572_, data_stage_5__2571_, data_stage_5__2570_, data_stage_5__2569_, data_stage_5__2568_, data_stage_5__2567_, data_stage_5__2566_, data_stage_5__2565_, data_stage_5__2564_, data_stage_5__2563_, data_stage_5__2562_, data_stage_5__2561_, data_stage_5__2560_, data_stage_5__2559_, data_stage_5__2558_, data_stage_5__2557_, data_stage_5__2556_, data_stage_5__2555_, data_stage_5__2554_, data_stage_5__2553_, data_stage_5__2552_, data_stage_5__2551_, data_stage_5__2550_, data_stage_5__2549_, data_stage_5__2548_, data_stage_5__2547_, data_stage_5__2546_, data_stage_5__2545_, data_stage_5__2544_, data_stage_5__2543_, data_stage_5__2542_, data_stage_5__2541_, data_stage_5__2540_, data_stage_5__2539_, data_stage_5__2538_, data_stage_5__2537_, data_stage_5__2536_, data_stage_5__2535_, data_stage_5__2534_, data_stage_5__2533_, data_stage_5__2532_, data_stage_5__2531_, data_stage_5__2530_, data_stage_5__2529_, data_stage_5__2528_, data_stage_5__2527_, data_stage_5__2526_, data_stage_5__2525_, data_stage_5__2524_, data_stage_5__2523_, data_stage_5__2522_, data_stage_5__2521_, data_stage_5__2520_, data_stage_5__2519_, data_stage_5__2518_, data_stage_5__2517_, data_stage_5__2516_, data_stage_5__2515_, data_stage_5__2514_, data_stage_5__2513_, data_stage_5__2512_, data_stage_5__2511_, data_stage_5__2510_, data_stage_5__2509_, data_stage_5__2508_, data_stage_5__2507_, data_stage_5__2506_, data_stage_5__2505_, data_stage_5__2504_, data_stage_5__2503_, data_stage_5__2502_, data_stage_5__2501_, data_stage_5__2500_, data_stage_5__2499_, data_stage_5__2498_, data_stage_5__2497_, data_stage_5__2496_, data_stage_5__2495_, data_stage_5__2494_, data_stage_5__2493_, data_stage_5__2492_, data_stage_5__2491_, data_stage_5__2490_, data_stage_5__2489_, data_stage_5__2488_, data_stage_5__2487_, data_stage_5__2486_, data_stage_5__2485_, data_stage_5__2484_, data_stage_5__2483_, data_stage_5__2482_, data_stage_5__2481_, data_stage_5__2480_, data_stage_5__2479_, data_stage_5__2478_, data_stage_5__2477_, data_stage_5__2476_, data_stage_5__2475_, data_stage_5__2474_, data_stage_5__2473_, data_stage_5__2472_, data_stage_5__2471_, data_stage_5__2470_, data_stage_5__2469_, data_stage_5__2468_, data_stage_5__2467_, data_stage_5__2466_, data_stage_5__2465_, data_stage_5__2464_, data_stage_5__2463_, data_stage_5__2462_, data_stage_5__2461_, data_stage_5__2460_, data_stage_5__2459_, data_stage_5__2458_, data_stage_5__2457_, data_stage_5__2456_, data_stage_5__2455_, data_stage_5__2454_, data_stage_5__2453_, data_stage_5__2452_, data_stage_5__2451_, data_stage_5__2450_, data_stage_5__2449_, data_stage_5__2448_, data_stage_5__2447_, data_stage_5__2446_, data_stage_5__2445_, data_stage_5__2444_, data_stage_5__2443_, data_stage_5__2442_, data_stage_5__2441_, data_stage_5__2440_, data_stage_5__2439_, data_stage_5__2438_, data_stage_5__2437_, data_stage_5__2436_, data_stage_5__2435_, data_stage_5__2434_, data_stage_5__2433_, data_stage_5__2432_, data_stage_5__2431_, data_stage_5__2430_, data_stage_5__2429_, data_stage_5__2428_, data_stage_5__2427_, data_stage_5__2426_, data_stage_5__2425_, data_stage_5__2424_, data_stage_5__2423_, data_stage_5__2422_, data_stage_5__2421_, data_stage_5__2420_, data_stage_5__2419_, data_stage_5__2418_, data_stage_5__2417_, data_stage_5__2416_, data_stage_5__2415_, data_stage_5__2414_, data_stage_5__2413_, data_stage_5__2412_, data_stage_5__2411_, data_stage_5__2410_, data_stage_5__2409_, data_stage_5__2408_, data_stage_5__2407_, data_stage_5__2406_, data_stage_5__2405_, data_stage_5__2404_, data_stage_5__2403_, data_stage_5__2402_, data_stage_5__2401_, data_stage_5__2400_, data_stage_5__2399_, data_stage_5__2398_, data_stage_5__2397_, data_stage_5__2396_, data_stage_5__2395_, data_stage_5__2394_, data_stage_5__2393_, data_stage_5__2392_, data_stage_5__2391_, data_stage_5__2390_, data_stage_5__2389_, data_stage_5__2388_, data_stage_5__2387_, data_stage_5__2386_, data_stage_5__2385_, data_stage_5__2384_, data_stage_5__2383_, data_stage_5__2382_, data_stage_5__2381_, data_stage_5__2380_, data_stage_5__2379_, data_stage_5__2378_, data_stage_5__2377_, data_stage_5__2376_, data_stage_5__2375_, data_stage_5__2374_, data_stage_5__2373_, data_stage_5__2372_, data_stage_5__2371_, data_stage_5__2370_, data_stage_5__2369_, data_stage_5__2368_, data_stage_5__2367_, data_stage_5__2366_, data_stage_5__2365_, data_stage_5__2364_, data_stage_5__2363_, data_stage_5__2362_, data_stage_5__2361_, data_stage_5__2360_, data_stage_5__2359_, data_stage_5__2358_, data_stage_5__2357_, data_stage_5__2356_, data_stage_5__2355_, data_stage_5__2354_, data_stage_5__2353_, data_stage_5__2352_, data_stage_5__2351_, data_stage_5__2350_, data_stage_5__2349_, data_stage_5__2348_, data_stage_5__2347_, data_stage_5__2346_, data_stage_5__2345_, data_stage_5__2344_, data_stage_5__2343_, data_stage_5__2342_, data_stage_5__2341_, data_stage_5__2340_, data_stage_5__2339_, data_stage_5__2338_, data_stage_5__2337_, data_stage_5__2336_, data_stage_5__2335_, data_stage_5__2334_, data_stage_5__2333_, data_stage_5__2332_, data_stage_5__2331_, data_stage_5__2330_, data_stage_5__2329_, data_stage_5__2328_, data_stage_5__2327_, data_stage_5__2326_, data_stage_5__2325_, data_stage_5__2324_, data_stage_5__2323_, data_stage_5__2322_, data_stage_5__2321_, data_stage_5__2320_, data_stage_5__2319_, data_stage_5__2318_, data_stage_5__2317_, data_stage_5__2316_, data_stage_5__2315_, data_stage_5__2314_, data_stage_5__2313_, data_stage_5__2312_, data_stage_5__2311_, data_stage_5__2310_, data_stage_5__2309_, data_stage_5__2308_, data_stage_5__2307_, data_stage_5__2306_, data_stage_5__2305_, data_stage_5__2304_, data_stage_5__2303_, data_stage_5__2302_, data_stage_5__2301_, data_stage_5__2300_, data_stage_5__2299_, data_stage_5__2298_, data_stage_5__2297_, data_stage_5__2296_, data_stage_5__2295_, data_stage_5__2294_, data_stage_5__2293_, data_stage_5__2292_, data_stage_5__2291_, data_stage_5__2290_, data_stage_5__2289_, data_stage_5__2288_, data_stage_5__2287_, data_stage_5__2286_, data_stage_5__2285_, data_stage_5__2284_, data_stage_5__2283_, data_stage_5__2282_, data_stage_5__2281_, data_stage_5__2280_, data_stage_5__2279_, data_stage_5__2278_, data_stage_5__2277_, data_stage_5__2276_, data_stage_5__2275_, data_stage_5__2274_, data_stage_5__2273_, data_stage_5__2272_, data_stage_5__2271_, data_stage_5__2270_, data_stage_5__2269_, data_stage_5__2268_, data_stage_5__2267_, data_stage_5__2266_, data_stage_5__2265_, data_stage_5__2264_, data_stage_5__2263_, data_stage_5__2262_, data_stage_5__2261_, data_stage_5__2260_, data_stage_5__2259_, data_stage_5__2258_, data_stage_5__2257_, data_stage_5__2256_, data_stage_5__2255_, data_stage_5__2254_, data_stage_5__2253_, data_stage_5__2252_, data_stage_5__2251_, data_stage_5__2250_, data_stage_5__2249_, data_stage_5__2248_, data_stage_5__2247_, data_stage_5__2246_, data_stage_5__2245_, data_stage_5__2244_, data_stage_5__2243_, data_stage_5__2242_, data_stage_5__2241_, data_stage_5__2240_, data_stage_5__2239_, data_stage_5__2238_, data_stage_5__2237_, data_stage_5__2236_, data_stage_5__2235_, data_stage_5__2234_, data_stage_5__2233_, data_stage_5__2232_, data_stage_5__2231_, data_stage_5__2230_, data_stage_5__2229_, data_stage_5__2228_, data_stage_5__2227_, data_stage_5__2226_, data_stage_5__2225_, data_stage_5__2224_, data_stage_5__2223_, data_stage_5__2222_, data_stage_5__2221_, data_stage_5__2220_, data_stage_5__2219_, data_stage_5__2218_, data_stage_5__2217_, data_stage_5__2216_, data_stage_5__2215_, data_stage_5__2214_, data_stage_5__2213_, data_stage_5__2212_, data_stage_5__2211_, data_stage_5__2210_, data_stage_5__2209_, data_stage_5__2208_, data_stage_5__2207_, data_stage_5__2206_, data_stage_5__2205_, data_stage_5__2204_, data_stage_5__2203_, data_stage_5__2202_, data_stage_5__2201_, data_stage_5__2200_, data_stage_5__2199_, data_stage_5__2198_, data_stage_5__2197_, data_stage_5__2196_, data_stage_5__2195_, data_stage_5__2194_, data_stage_5__2193_, data_stage_5__2192_, data_stage_5__2191_, data_stage_5__2190_, data_stage_5__2189_, data_stage_5__2188_, data_stage_5__2187_, data_stage_5__2186_, data_stage_5__2185_, data_stage_5__2184_, data_stage_5__2183_, data_stage_5__2182_, data_stage_5__2181_, data_stage_5__2180_, data_stage_5__2179_, data_stage_5__2178_, data_stage_5__2177_, data_stage_5__2176_, data_stage_5__2175_, data_stage_5__2174_, data_stage_5__2173_, data_stage_5__2172_, data_stage_5__2171_, data_stage_5__2170_, data_stage_5__2169_, data_stage_5__2168_, data_stage_5__2167_, data_stage_5__2166_, data_stage_5__2165_, data_stage_5__2164_, data_stage_5__2163_, data_stage_5__2162_, data_stage_5__2161_, data_stage_5__2160_, data_stage_5__2159_, data_stage_5__2158_, data_stage_5__2157_, data_stage_5__2156_, data_stage_5__2155_, data_stage_5__2154_, data_stage_5__2153_, data_stage_5__2152_, data_stage_5__2151_, data_stage_5__2150_, data_stage_5__2149_, data_stage_5__2148_, data_stage_5__2147_, data_stage_5__2146_, data_stage_5__2145_, data_stage_5__2144_, data_stage_5__2143_, data_stage_5__2142_, data_stage_5__2141_, data_stage_5__2140_, data_stage_5__2139_, data_stage_5__2138_, data_stage_5__2137_, data_stage_5__2136_, data_stage_5__2135_, data_stage_5__2134_, data_stage_5__2133_, data_stage_5__2132_, data_stage_5__2131_, data_stage_5__2130_, data_stage_5__2129_, data_stage_5__2128_, data_stage_5__2127_, data_stage_5__2126_, data_stage_5__2125_, data_stage_5__2124_, data_stage_5__2123_, data_stage_5__2122_, data_stage_5__2121_, data_stage_5__2120_, data_stage_5__2119_, data_stage_5__2118_, data_stage_5__2117_, data_stage_5__2116_, data_stage_5__2115_, data_stage_5__2114_, data_stage_5__2113_, data_stage_5__2112_, data_stage_5__2111_, data_stage_5__2110_, data_stage_5__2109_, data_stage_5__2108_, data_stage_5__2107_, data_stage_5__2106_, data_stage_5__2105_, data_stage_5__2104_, data_stage_5__2103_, data_stage_5__2102_, data_stage_5__2101_, data_stage_5__2100_, data_stage_5__2099_, data_stage_5__2098_, data_stage_5__2097_, data_stage_5__2096_, data_stage_5__2095_, data_stage_5__2094_, data_stage_5__2093_, data_stage_5__2092_, data_stage_5__2091_, data_stage_5__2090_, data_stage_5__2089_, data_stage_5__2088_, data_stage_5__2087_, data_stage_5__2086_, data_stage_5__2085_, data_stage_5__2084_, data_stage_5__2083_, data_stage_5__2082_, data_stage_5__2081_, data_stage_5__2080_, data_stage_5__2079_, data_stage_5__2078_, data_stage_5__2077_, data_stage_5__2076_, data_stage_5__2075_, data_stage_5__2074_, data_stage_5__2073_, data_stage_5__2072_, data_stage_5__2071_, data_stage_5__2070_, data_stage_5__2069_, data_stage_5__2068_, data_stage_5__2067_, data_stage_5__2066_, data_stage_5__2065_, data_stage_5__2064_, data_stage_5__2063_, data_stage_5__2062_, data_stage_5__2061_, data_stage_5__2060_, data_stage_5__2059_, data_stage_5__2058_, data_stage_5__2057_, data_stage_5__2056_, data_stage_5__2055_, data_stage_5__2054_, data_stage_5__2053_, data_stage_5__2052_, data_stage_5__2051_, data_stage_5__2050_, data_stage_5__2049_, data_stage_5__2048_, data_stage_5__2047_, data_stage_5__2046_, data_stage_5__2045_, data_stage_5__2044_, data_stage_5__2043_, data_stage_5__2042_, data_stage_5__2041_, data_stage_5__2040_, data_stage_5__2039_, data_stage_5__2038_, data_stage_5__2037_, data_stage_5__2036_, data_stage_5__2035_, data_stage_5__2034_, data_stage_5__2033_, data_stage_5__2032_, data_stage_5__2031_, data_stage_5__2030_, data_stage_5__2029_, data_stage_5__2028_, data_stage_5__2027_, data_stage_5__2026_, data_stage_5__2025_, data_stage_5__2024_, data_stage_5__2023_, data_stage_5__2022_, data_stage_5__2021_, data_stage_5__2020_, data_stage_5__2019_, data_stage_5__2018_, data_stage_5__2017_, data_stage_5__2016_, data_stage_5__2015_, data_stage_5__2014_, data_stage_5__2013_, data_stage_5__2012_, data_stage_5__2011_, data_stage_5__2010_, data_stage_5__2009_, data_stage_5__2008_, data_stage_5__2007_, data_stage_5__2006_, data_stage_5__2005_, data_stage_5__2004_, data_stage_5__2003_, data_stage_5__2002_, data_stage_5__2001_, data_stage_5__2000_, data_stage_5__1999_, data_stage_5__1998_, data_stage_5__1997_, data_stage_5__1996_, data_stage_5__1995_, data_stage_5__1994_, data_stage_5__1993_, data_stage_5__1992_, data_stage_5__1991_, data_stage_5__1990_, data_stage_5__1989_, data_stage_5__1988_, data_stage_5__1987_, data_stage_5__1986_, data_stage_5__1985_, data_stage_5__1984_, data_stage_5__1983_, data_stage_5__1982_, data_stage_5__1981_, data_stage_5__1980_, data_stage_5__1979_, data_stage_5__1978_, data_stage_5__1977_, data_stage_5__1976_, data_stage_5__1975_, data_stage_5__1974_, data_stage_5__1973_, data_stage_5__1972_, data_stage_5__1971_, data_stage_5__1970_, data_stage_5__1969_, data_stage_5__1968_, data_stage_5__1967_, data_stage_5__1966_, data_stage_5__1965_, data_stage_5__1964_, data_stage_5__1963_, data_stage_5__1962_, data_stage_5__1961_, data_stage_5__1960_, data_stage_5__1959_, data_stage_5__1958_, data_stage_5__1957_, data_stage_5__1956_, data_stage_5__1955_, data_stage_5__1954_, data_stage_5__1953_, data_stage_5__1952_, data_stage_5__1951_, data_stage_5__1950_, data_stage_5__1949_, data_stage_5__1948_, data_stage_5__1947_, data_stage_5__1946_, data_stage_5__1945_, data_stage_5__1944_, data_stage_5__1943_, data_stage_5__1942_, data_stage_5__1941_, data_stage_5__1940_, data_stage_5__1939_, data_stage_5__1938_, data_stage_5__1937_, data_stage_5__1936_, data_stage_5__1935_, data_stage_5__1934_, data_stage_5__1933_, data_stage_5__1932_, data_stage_5__1931_, data_stage_5__1930_, data_stage_5__1929_, data_stage_5__1928_, data_stage_5__1927_, data_stage_5__1926_, data_stage_5__1925_, data_stage_5__1924_, data_stage_5__1923_, data_stage_5__1922_, data_stage_5__1921_, data_stage_5__1920_, data_stage_5__1919_, data_stage_5__1918_, data_stage_5__1917_, data_stage_5__1916_, data_stage_5__1915_, data_stage_5__1914_, data_stage_5__1913_, data_stage_5__1912_, data_stage_5__1911_, data_stage_5__1910_, data_stage_5__1909_, data_stage_5__1908_, data_stage_5__1907_, data_stage_5__1906_, data_stage_5__1905_, data_stage_5__1904_, data_stage_5__1903_, data_stage_5__1902_, data_stage_5__1901_, data_stage_5__1900_, data_stage_5__1899_, data_stage_5__1898_, data_stage_5__1897_, data_stage_5__1896_, data_stage_5__1895_, data_stage_5__1894_, data_stage_5__1893_, data_stage_5__1892_, data_stage_5__1891_, data_stage_5__1890_, data_stage_5__1889_, data_stage_5__1888_, data_stage_5__1887_, data_stage_5__1886_, data_stage_5__1885_, data_stage_5__1884_, data_stage_5__1883_, data_stage_5__1882_, data_stage_5__1881_, data_stage_5__1880_, data_stage_5__1879_, data_stage_5__1878_, data_stage_5__1877_, data_stage_5__1876_, data_stage_5__1875_, data_stage_5__1874_, data_stage_5__1873_, data_stage_5__1872_, data_stage_5__1871_, data_stage_5__1870_, data_stage_5__1869_, data_stage_5__1868_, data_stage_5__1867_, data_stage_5__1866_, data_stage_5__1865_, data_stage_5__1864_, data_stage_5__1863_, data_stage_5__1862_, data_stage_5__1861_, data_stage_5__1860_, data_stage_5__1859_, data_stage_5__1858_, data_stage_5__1857_, data_stage_5__1856_, data_stage_5__1855_, data_stage_5__1854_, data_stage_5__1853_, data_stage_5__1852_, data_stage_5__1851_, data_stage_5__1850_, data_stage_5__1849_, data_stage_5__1848_, data_stage_5__1847_, data_stage_5__1846_, data_stage_5__1845_, data_stage_5__1844_, data_stage_5__1843_, data_stage_5__1842_, data_stage_5__1841_, data_stage_5__1840_, data_stage_5__1839_, data_stage_5__1838_, data_stage_5__1837_, data_stage_5__1836_, data_stage_5__1835_, data_stage_5__1834_, data_stage_5__1833_, data_stage_5__1832_, data_stage_5__1831_, data_stage_5__1830_, data_stage_5__1829_, data_stage_5__1828_, data_stage_5__1827_, data_stage_5__1826_, data_stage_5__1825_, data_stage_5__1824_, data_stage_5__1823_, data_stage_5__1822_, data_stage_5__1821_, data_stage_5__1820_, data_stage_5__1819_, data_stage_5__1818_, data_stage_5__1817_, data_stage_5__1816_, data_stage_5__1815_, data_stage_5__1814_, data_stage_5__1813_, data_stage_5__1812_, data_stage_5__1811_, data_stage_5__1810_, data_stage_5__1809_, data_stage_5__1808_, data_stage_5__1807_, data_stage_5__1806_, data_stage_5__1805_, data_stage_5__1804_, data_stage_5__1803_, data_stage_5__1802_, data_stage_5__1801_, data_stage_5__1800_, data_stage_5__1799_, data_stage_5__1798_, data_stage_5__1797_, data_stage_5__1796_, data_stage_5__1795_, data_stage_5__1794_, data_stage_5__1793_, data_stage_5__1792_, data_stage_5__1791_, data_stage_5__1790_, data_stage_5__1789_, data_stage_5__1788_, data_stage_5__1787_, data_stage_5__1786_, data_stage_5__1785_, data_stage_5__1784_, data_stage_5__1783_, data_stage_5__1782_, data_stage_5__1781_, data_stage_5__1780_, data_stage_5__1779_, data_stage_5__1778_, data_stage_5__1777_, data_stage_5__1776_, data_stage_5__1775_, data_stage_5__1774_, data_stage_5__1773_, data_stage_5__1772_, data_stage_5__1771_, data_stage_5__1770_, data_stage_5__1769_, data_stage_5__1768_, data_stage_5__1767_, data_stage_5__1766_, data_stage_5__1765_, data_stage_5__1764_, data_stage_5__1763_, data_stage_5__1762_, data_stage_5__1761_, data_stage_5__1760_, data_stage_5__1759_, data_stage_5__1758_, data_stage_5__1757_, data_stage_5__1756_, data_stage_5__1755_, data_stage_5__1754_, data_stage_5__1753_, data_stage_5__1752_, data_stage_5__1751_, data_stage_5__1750_, data_stage_5__1749_, data_stage_5__1748_, data_stage_5__1747_, data_stage_5__1746_, data_stage_5__1745_, data_stage_5__1744_, data_stage_5__1743_, data_stage_5__1742_, data_stage_5__1741_, data_stage_5__1740_, data_stage_5__1739_, data_stage_5__1738_, data_stage_5__1737_, data_stage_5__1736_, data_stage_5__1735_, data_stage_5__1734_, data_stage_5__1733_, data_stage_5__1732_, data_stage_5__1731_, data_stage_5__1730_, data_stage_5__1729_, data_stage_5__1728_, data_stage_5__1727_, data_stage_5__1726_, data_stage_5__1725_, data_stage_5__1724_, data_stage_5__1723_, data_stage_5__1722_, data_stage_5__1721_, data_stage_5__1720_, data_stage_5__1719_, data_stage_5__1718_, data_stage_5__1717_, data_stage_5__1716_, data_stage_5__1715_, data_stage_5__1714_, data_stage_5__1713_, data_stage_5__1712_, data_stage_5__1711_, data_stage_5__1710_, data_stage_5__1709_, data_stage_5__1708_, data_stage_5__1707_, data_stage_5__1706_, data_stage_5__1705_, data_stage_5__1704_, data_stage_5__1703_, data_stage_5__1702_, data_stage_5__1701_, data_stage_5__1700_, data_stage_5__1699_, data_stage_5__1698_, data_stage_5__1697_, data_stage_5__1696_, data_stage_5__1695_, data_stage_5__1694_, data_stage_5__1693_, data_stage_5__1692_, data_stage_5__1691_, data_stage_5__1690_, data_stage_5__1689_, data_stage_5__1688_, data_stage_5__1687_, data_stage_5__1686_, data_stage_5__1685_, data_stage_5__1684_, data_stage_5__1683_, data_stage_5__1682_, data_stage_5__1681_, data_stage_5__1680_, data_stage_5__1679_, data_stage_5__1678_, data_stage_5__1677_, data_stage_5__1676_, data_stage_5__1675_, data_stage_5__1674_, data_stage_5__1673_, data_stage_5__1672_, data_stage_5__1671_, data_stage_5__1670_, data_stage_5__1669_, data_stage_5__1668_, data_stage_5__1667_, data_stage_5__1666_, data_stage_5__1665_, data_stage_5__1664_, data_stage_5__1663_, data_stage_5__1662_, data_stage_5__1661_, data_stage_5__1660_, data_stage_5__1659_, data_stage_5__1658_, data_stage_5__1657_, data_stage_5__1656_, data_stage_5__1655_, data_stage_5__1654_, data_stage_5__1653_, data_stage_5__1652_, data_stage_5__1651_, data_stage_5__1650_, data_stage_5__1649_, data_stage_5__1648_, data_stage_5__1647_, data_stage_5__1646_, data_stage_5__1645_, data_stage_5__1644_, data_stage_5__1643_, data_stage_5__1642_, data_stage_5__1641_, data_stage_5__1640_, data_stage_5__1639_, data_stage_5__1638_, data_stage_5__1637_, data_stage_5__1636_, data_stage_5__1635_, data_stage_5__1634_, data_stage_5__1633_, data_stage_5__1632_, data_stage_5__1631_, data_stage_5__1630_, data_stage_5__1629_, data_stage_5__1628_, data_stage_5__1627_, data_stage_5__1626_, data_stage_5__1625_, data_stage_5__1624_, data_stage_5__1623_, data_stage_5__1622_, data_stage_5__1621_, data_stage_5__1620_, data_stage_5__1619_, data_stage_5__1618_, data_stage_5__1617_, data_stage_5__1616_, data_stage_5__1615_, data_stage_5__1614_, data_stage_5__1613_, data_stage_5__1612_, data_stage_5__1611_, data_stage_5__1610_, data_stage_5__1609_, data_stage_5__1608_, data_stage_5__1607_, data_stage_5__1606_, data_stage_5__1605_, data_stage_5__1604_, data_stage_5__1603_, data_stage_5__1602_, data_stage_5__1601_, data_stage_5__1600_, data_stage_5__1599_, data_stage_5__1598_, data_stage_5__1597_, data_stage_5__1596_, data_stage_5__1595_, data_stage_5__1594_, data_stage_5__1593_, data_stage_5__1592_, data_stage_5__1591_, data_stage_5__1590_, data_stage_5__1589_, data_stage_5__1588_, data_stage_5__1587_, data_stage_5__1586_, data_stage_5__1585_, data_stage_5__1584_, data_stage_5__1583_, data_stage_5__1582_, data_stage_5__1581_, data_stage_5__1580_, data_stage_5__1579_, data_stage_5__1578_, data_stage_5__1577_, data_stage_5__1576_, data_stage_5__1575_, data_stage_5__1574_, data_stage_5__1573_, data_stage_5__1572_, data_stage_5__1571_, data_stage_5__1570_, data_stage_5__1569_, data_stage_5__1568_, data_stage_5__1567_, data_stage_5__1566_, data_stage_5__1565_, data_stage_5__1564_, data_stage_5__1563_, data_stage_5__1562_, data_stage_5__1561_, data_stage_5__1560_, data_stage_5__1559_, data_stage_5__1558_, data_stage_5__1557_, data_stage_5__1556_, data_stage_5__1555_, data_stage_5__1554_, data_stage_5__1553_, data_stage_5__1552_, data_stage_5__1551_, data_stage_5__1550_, data_stage_5__1549_, data_stage_5__1548_, data_stage_5__1547_, data_stage_5__1546_, data_stage_5__1545_, data_stage_5__1544_, data_stage_5__1543_, data_stage_5__1542_, data_stage_5__1541_, data_stage_5__1540_, data_stage_5__1539_, data_stage_5__1538_, data_stage_5__1537_, data_stage_5__1536_, data_stage_5__1535_, data_stage_5__1534_, data_stage_5__1533_, data_stage_5__1532_, data_stage_5__1531_, data_stage_5__1530_, data_stage_5__1529_, data_stage_5__1528_, data_stage_5__1527_, data_stage_5__1526_, data_stage_5__1525_, data_stage_5__1524_, data_stage_5__1523_, data_stage_5__1522_, data_stage_5__1521_, data_stage_5__1520_, data_stage_5__1519_, data_stage_5__1518_, data_stage_5__1517_, data_stage_5__1516_, data_stage_5__1515_, data_stage_5__1514_, data_stage_5__1513_, data_stage_5__1512_, data_stage_5__1511_, data_stage_5__1510_, data_stage_5__1509_, data_stage_5__1508_, data_stage_5__1507_, data_stage_5__1506_, data_stage_5__1505_, data_stage_5__1504_, data_stage_5__1503_, data_stage_5__1502_, data_stage_5__1501_, data_stage_5__1500_, data_stage_5__1499_, data_stage_5__1498_, data_stage_5__1497_, data_stage_5__1496_, data_stage_5__1495_, data_stage_5__1494_, data_stage_5__1493_, data_stage_5__1492_, data_stage_5__1491_, data_stage_5__1490_, data_stage_5__1489_, data_stage_5__1488_, data_stage_5__1487_, data_stage_5__1486_, data_stage_5__1485_, data_stage_5__1484_, data_stage_5__1483_, data_stage_5__1482_, data_stage_5__1481_, data_stage_5__1480_, data_stage_5__1479_, data_stage_5__1478_, data_stage_5__1477_, data_stage_5__1476_, data_stage_5__1475_, data_stage_5__1474_, data_stage_5__1473_, data_stage_5__1472_, data_stage_5__1471_, data_stage_5__1470_, data_stage_5__1469_, data_stage_5__1468_, data_stage_5__1467_, data_stage_5__1466_, data_stage_5__1465_, data_stage_5__1464_, data_stage_5__1463_, data_stage_5__1462_, data_stage_5__1461_, data_stage_5__1460_, data_stage_5__1459_, data_stage_5__1458_, data_stage_5__1457_, data_stage_5__1456_, data_stage_5__1455_, data_stage_5__1454_, data_stage_5__1453_, data_stage_5__1452_, data_stage_5__1451_, data_stage_5__1450_, data_stage_5__1449_, data_stage_5__1448_, data_stage_5__1447_, data_stage_5__1446_, data_stage_5__1445_, data_stage_5__1444_, data_stage_5__1443_, data_stage_5__1442_, data_stage_5__1441_, data_stage_5__1440_, data_stage_5__1439_, data_stage_5__1438_, data_stage_5__1437_, data_stage_5__1436_, data_stage_5__1435_, data_stage_5__1434_, data_stage_5__1433_, data_stage_5__1432_, data_stage_5__1431_, data_stage_5__1430_, data_stage_5__1429_, data_stage_5__1428_, data_stage_5__1427_, data_stage_5__1426_, data_stage_5__1425_, data_stage_5__1424_, data_stage_5__1423_, data_stage_5__1422_, data_stage_5__1421_, data_stage_5__1420_, data_stage_5__1419_, data_stage_5__1418_, data_stage_5__1417_, data_stage_5__1416_, data_stage_5__1415_, data_stage_5__1414_, data_stage_5__1413_, data_stage_5__1412_, data_stage_5__1411_, data_stage_5__1410_, data_stage_5__1409_, data_stage_5__1408_, data_stage_5__1407_, data_stage_5__1406_, data_stage_5__1405_, data_stage_5__1404_, data_stage_5__1403_, data_stage_5__1402_, data_stage_5__1401_, data_stage_5__1400_, data_stage_5__1399_, data_stage_5__1398_, data_stage_5__1397_, data_stage_5__1396_, data_stage_5__1395_, data_stage_5__1394_, data_stage_5__1393_, data_stage_5__1392_, data_stage_5__1391_, data_stage_5__1390_, data_stage_5__1389_, data_stage_5__1388_, data_stage_5__1387_, data_stage_5__1386_, data_stage_5__1385_, data_stage_5__1384_, data_stage_5__1383_, data_stage_5__1382_, data_stage_5__1381_, data_stage_5__1380_, data_stage_5__1379_, data_stage_5__1378_, data_stage_5__1377_, data_stage_5__1376_, data_stage_5__1375_, data_stage_5__1374_, data_stage_5__1373_, data_stage_5__1372_, data_stage_5__1371_, data_stage_5__1370_, data_stage_5__1369_, data_stage_5__1368_, data_stage_5__1367_, data_stage_5__1366_, data_stage_5__1365_, data_stage_5__1364_, data_stage_5__1363_, data_stage_5__1362_, data_stage_5__1361_, data_stage_5__1360_, data_stage_5__1359_, data_stage_5__1358_, data_stage_5__1357_, data_stage_5__1356_, data_stage_5__1355_, data_stage_5__1354_, data_stage_5__1353_, data_stage_5__1352_, data_stage_5__1351_, data_stage_5__1350_, data_stage_5__1349_, data_stage_5__1348_, data_stage_5__1347_, data_stage_5__1346_, data_stage_5__1345_, data_stage_5__1344_, data_stage_5__1343_, data_stage_5__1342_, data_stage_5__1341_, data_stage_5__1340_, data_stage_5__1339_, data_stage_5__1338_, data_stage_5__1337_, data_stage_5__1336_, data_stage_5__1335_, data_stage_5__1334_, data_stage_5__1333_, data_stage_5__1332_, data_stage_5__1331_, data_stage_5__1330_, data_stage_5__1329_, data_stage_5__1328_, data_stage_5__1327_, data_stage_5__1326_, data_stage_5__1325_, data_stage_5__1324_, data_stage_5__1323_, data_stage_5__1322_, data_stage_5__1321_, data_stage_5__1320_, data_stage_5__1319_, data_stage_5__1318_, data_stage_5__1317_, data_stage_5__1316_, data_stage_5__1315_, data_stage_5__1314_, data_stage_5__1313_, data_stage_5__1312_, data_stage_5__1311_, data_stage_5__1310_, data_stage_5__1309_, data_stage_5__1308_, data_stage_5__1307_, data_stage_5__1306_, data_stage_5__1305_, data_stage_5__1304_, data_stage_5__1303_, data_stage_5__1302_, data_stage_5__1301_, data_stage_5__1300_, data_stage_5__1299_, data_stage_5__1298_, data_stage_5__1297_, data_stage_5__1296_, data_stage_5__1295_, data_stage_5__1294_, data_stage_5__1293_, data_stage_5__1292_, data_stage_5__1291_, data_stage_5__1290_, data_stage_5__1289_, data_stage_5__1288_, data_stage_5__1287_, data_stage_5__1286_, data_stage_5__1285_, data_stage_5__1284_, data_stage_5__1283_, data_stage_5__1282_, data_stage_5__1281_, data_stage_5__1280_, data_stage_5__1279_, data_stage_5__1278_, data_stage_5__1277_, data_stage_5__1276_, data_stage_5__1275_, data_stage_5__1274_, data_stage_5__1273_, data_stage_5__1272_, data_stage_5__1271_, data_stage_5__1270_, data_stage_5__1269_, data_stage_5__1268_, data_stage_5__1267_, data_stage_5__1266_, data_stage_5__1265_, data_stage_5__1264_, data_stage_5__1263_, data_stage_5__1262_, data_stage_5__1261_, data_stage_5__1260_, data_stage_5__1259_, data_stage_5__1258_, data_stage_5__1257_, data_stage_5__1256_, data_stage_5__1255_, data_stage_5__1254_, data_stage_5__1253_, data_stage_5__1252_, data_stage_5__1251_, data_stage_5__1250_, data_stage_5__1249_, data_stage_5__1248_, data_stage_5__1247_, data_stage_5__1246_, data_stage_5__1245_, data_stage_5__1244_, data_stage_5__1243_, data_stage_5__1242_, data_stage_5__1241_, data_stage_5__1240_, data_stage_5__1239_, data_stage_5__1238_, data_stage_5__1237_, data_stage_5__1236_, data_stage_5__1235_, data_stage_5__1234_, data_stage_5__1233_, data_stage_5__1232_, data_stage_5__1231_, data_stage_5__1230_, data_stage_5__1229_, data_stage_5__1228_, data_stage_5__1227_, data_stage_5__1226_, data_stage_5__1225_, data_stage_5__1224_, data_stage_5__1223_, data_stage_5__1222_, data_stage_5__1221_, data_stage_5__1220_, data_stage_5__1219_, data_stage_5__1218_, data_stage_5__1217_, data_stage_5__1216_, data_stage_5__1215_, data_stage_5__1214_, data_stage_5__1213_, data_stage_5__1212_, data_stage_5__1211_, data_stage_5__1210_, data_stage_5__1209_, data_stage_5__1208_, data_stage_5__1207_, data_stage_5__1206_, data_stage_5__1205_, data_stage_5__1204_, data_stage_5__1203_, data_stage_5__1202_, data_stage_5__1201_, data_stage_5__1200_, data_stage_5__1199_, data_stage_5__1198_, data_stage_5__1197_, data_stage_5__1196_, data_stage_5__1195_, data_stage_5__1194_, data_stage_5__1193_, data_stage_5__1192_, data_stage_5__1191_, data_stage_5__1190_, data_stage_5__1189_, data_stage_5__1188_, data_stage_5__1187_, data_stage_5__1186_, data_stage_5__1185_, data_stage_5__1184_, data_stage_5__1183_, data_stage_5__1182_, data_stage_5__1181_, data_stage_5__1180_, data_stage_5__1179_, data_stage_5__1178_, data_stage_5__1177_, data_stage_5__1176_, data_stage_5__1175_, data_stage_5__1174_, data_stage_5__1173_, data_stage_5__1172_, data_stage_5__1171_, data_stage_5__1170_, data_stage_5__1169_, data_stage_5__1168_, data_stage_5__1167_, data_stage_5__1166_, data_stage_5__1165_, data_stage_5__1164_, data_stage_5__1163_, data_stage_5__1162_, data_stage_5__1161_, data_stage_5__1160_, data_stage_5__1159_, data_stage_5__1158_, data_stage_5__1157_, data_stage_5__1156_, data_stage_5__1155_, data_stage_5__1154_, data_stage_5__1153_, data_stage_5__1152_, data_stage_5__1151_, data_stage_5__1150_, data_stage_5__1149_, data_stage_5__1148_, data_stage_5__1147_, data_stage_5__1146_, data_stage_5__1145_, data_stage_5__1144_, data_stage_5__1143_, data_stage_5__1142_, data_stage_5__1141_, data_stage_5__1140_, data_stage_5__1139_, data_stage_5__1138_, data_stage_5__1137_, data_stage_5__1136_, data_stage_5__1135_, data_stage_5__1134_, data_stage_5__1133_, data_stage_5__1132_, data_stage_5__1131_, data_stage_5__1130_, data_stage_5__1129_, data_stage_5__1128_, data_stage_5__1127_, data_stage_5__1126_, data_stage_5__1125_, data_stage_5__1124_, data_stage_5__1123_, data_stage_5__1122_, data_stage_5__1121_, data_stage_5__1120_, data_stage_5__1119_, data_stage_5__1118_, data_stage_5__1117_, data_stage_5__1116_, data_stage_5__1115_, data_stage_5__1114_, data_stage_5__1113_, data_stage_5__1112_, data_stage_5__1111_, data_stage_5__1110_, data_stage_5__1109_, data_stage_5__1108_, data_stage_5__1107_, data_stage_5__1106_, data_stage_5__1105_, data_stage_5__1104_, data_stage_5__1103_, data_stage_5__1102_, data_stage_5__1101_, data_stage_5__1100_, data_stage_5__1099_, data_stage_5__1098_, data_stage_5__1097_, data_stage_5__1096_, data_stage_5__1095_, data_stage_5__1094_, data_stage_5__1093_, data_stage_5__1092_, data_stage_5__1091_, data_stage_5__1090_, data_stage_5__1089_, data_stage_5__1088_, data_stage_5__1087_, data_stage_5__1086_, data_stage_5__1085_, data_stage_5__1084_, data_stage_5__1083_, data_stage_5__1082_, data_stage_5__1081_, data_stage_5__1080_, data_stage_5__1079_, data_stage_5__1078_, data_stage_5__1077_, data_stage_5__1076_, data_stage_5__1075_, data_stage_5__1074_, data_stage_5__1073_, data_stage_5__1072_, data_stage_5__1071_, data_stage_5__1070_, data_stage_5__1069_, data_stage_5__1068_, data_stage_5__1067_, data_stage_5__1066_, data_stage_5__1065_, data_stage_5__1064_, data_stage_5__1063_, data_stage_5__1062_, data_stage_5__1061_, data_stage_5__1060_, data_stage_5__1059_, data_stage_5__1058_, data_stage_5__1057_, data_stage_5__1056_, data_stage_5__1055_, data_stage_5__1054_, data_stage_5__1053_, data_stage_5__1052_, data_stage_5__1051_, data_stage_5__1050_, data_stage_5__1049_, data_stage_5__1048_, data_stage_5__1047_, data_stage_5__1046_, data_stage_5__1045_, data_stage_5__1044_, data_stage_5__1043_, data_stage_5__1042_, data_stage_5__1041_, data_stage_5__1040_, data_stage_5__1039_, data_stage_5__1038_, data_stage_5__1037_, data_stage_5__1036_, data_stage_5__1035_, data_stage_5__1034_, data_stage_5__1033_, data_stage_5__1032_, data_stage_5__1031_, data_stage_5__1030_, data_stage_5__1029_, data_stage_5__1028_, data_stage_5__1027_, data_stage_5__1026_, data_stage_5__1025_, data_stage_5__1024_, data_stage_5__1023_, data_stage_5__1022_, data_stage_5__1021_, data_stage_5__1020_, data_stage_5__1019_, data_stage_5__1018_, data_stage_5__1017_, data_stage_5__1016_, data_stage_5__1015_, data_stage_5__1014_, data_stage_5__1013_, data_stage_5__1012_, data_stage_5__1011_, data_stage_5__1010_, data_stage_5__1009_, data_stage_5__1008_, data_stage_5__1007_, data_stage_5__1006_, data_stage_5__1005_, data_stage_5__1004_, data_stage_5__1003_, data_stage_5__1002_, data_stage_5__1001_, data_stage_5__1000_, data_stage_5__999_, data_stage_5__998_, data_stage_5__997_, data_stage_5__996_, data_stage_5__995_, data_stage_5__994_, data_stage_5__993_, data_stage_5__992_, data_stage_5__991_, data_stage_5__990_, data_stage_5__989_, data_stage_5__988_, data_stage_5__987_, data_stage_5__986_, data_stage_5__985_, data_stage_5__984_, data_stage_5__983_, data_stage_5__982_, data_stage_5__981_, data_stage_5__980_, data_stage_5__979_, data_stage_5__978_, data_stage_5__977_, data_stage_5__976_, data_stage_5__975_, data_stage_5__974_, data_stage_5__973_, data_stage_5__972_, data_stage_5__971_, data_stage_5__970_, data_stage_5__969_, data_stage_5__968_, data_stage_5__967_, data_stage_5__966_, data_stage_5__965_, data_stage_5__964_, data_stage_5__963_, data_stage_5__962_, data_stage_5__961_, data_stage_5__960_, data_stage_5__959_, data_stage_5__958_, data_stage_5__957_, data_stage_5__956_, data_stage_5__955_, data_stage_5__954_, data_stage_5__953_, data_stage_5__952_, data_stage_5__951_, data_stage_5__950_, data_stage_5__949_, data_stage_5__948_, data_stage_5__947_, data_stage_5__946_, data_stage_5__945_, data_stage_5__944_, data_stage_5__943_, data_stage_5__942_, data_stage_5__941_, data_stage_5__940_, data_stage_5__939_, data_stage_5__938_, data_stage_5__937_, data_stage_5__936_, data_stage_5__935_, data_stage_5__934_, data_stage_5__933_, data_stage_5__932_, data_stage_5__931_, data_stage_5__930_, data_stage_5__929_, data_stage_5__928_, data_stage_5__927_, data_stage_5__926_, data_stage_5__925_, data_stage_5__924_, data_stage_5__923_, data_stage_5__922_, data_stage_5__921_, data_stage_5__920_, data_stage_5__919_, data_stage_5__918_, data_stage_5__917_, data_stage_5__916_, data_stage_5__915_, data_stage_5__914_, data_stage_5__913_, data_stage_5__912_, data_stage_5__911_, data_stage_5__910_, data_stage_5__909_, data_stage_5__908_, data_stage_5__907_, data_stage_5__906_, data_stage_5__905_, data_stage_5__904_, data_stage_5__903_, data_stage_5__902_, data_stage_5__901_, data_stage_5__900_, data_stage_5__899_, data_stage_5__898_, data_stage_5__897_, data_stage_5__896_, data_stage_5__895_, data_stage_5__894_, data_stage_5__893_, data_stage_5__892_, data_stage_5__891_, data_stage_5__890_, data_stage_5__889_, data_stage_5__888_, data_stage_5__887_, data_stage_5__886_, data_stage_5__885_, data_stage_5__884_, data_stage_5__883_, data_stage_5__882_, data_stage_5__881_, data_stage_5__880_, data_stage_5__879_, data_stage_5__878_, data_stage_5__877_, data_stage_5__876_, data_stage_5__875_, data_stage_5__874_, data_stage_5__873_, data_stage_5__872_, data_stage_5__871_, data_stage_5__870_, data_stage_5__869_, data_stage_5__868_, data_stage_5__867_, data_stage_5__866_, data_stage_5__865_, data_stage_5__864_, data_stage_5__863_, data_stage_5__862_, data_stage_5__861_, data_stage_5__860_, data_stage_5__859_, data_stage_5__858_, data_stage_5__857_, data_stage_5__856_, data_stage_5__855_, data_stage_5__854_, data_stage_5__853_, data_stage_5__852_, data_stage_5__851_, data_stage_5__850_, data_stage_5__849_, data_stage_5__848_, data_stage_5__847_, data_stage_5__846_, data_stage_5__845_, data_stage_5__844_, data_stage_5__843_, data_stage_5__842_, data_stage_5__841_, data_stage_5__840_, data_stage_5__839_, data_stage_5__838_, data_stage_5__837_, data_stage_5__836_, data_stage_5__835_, data_stage_5__834_, data_stage_5__833_, data_stage_5__832_, data_stage_5__831_, data_stage_5__830_, data_stage_5__829_, data_stage_5__828_, data_stage_5__827_, data_stage_5__826_, data_stage_5__825_, data_stage_5__824_, data_stage_5__823_, data_stage_5__822_, data_stage_5__821_, data_stage_5__820_, data_stage_5__819_, data_stage_5__818_, data_stage_5__817_, data_stage_5__816_, data_stage_5__815_, data_stage_5__814_, data_stage_5__813_, data_stage_5__812_, data_stage_5__811_, data_stage_5__810_, data_stage_5__809_, data_stage_5__808_, data_stage_5__807_, data_stage_5__806_, data_stage_5__805_, data_stage_5__804_, data_stage_5__803_, data_stage_5__802_, data_stage_5__801_, data_stage_5__800_, data_stage_5__799_, data_stage_5__798_, data_stage_5__797_, data_stage_5__796_, data_stage_5__795_, data_stage_5__794_, data_stage_5__793_, data_stage_5__792_, data_stage_5__791_, data_stage_5__790_, data_stage_5__789_, data_stage_5__788_, data_stage_5__787_, data_stage_5__786_, data_stage_5__785_, data_stage_5__784_, data_stage_5__783_, data_stage_5__782_, data_stage_5__781_, data_stage_5__780_, data_stage_5__779_, data_stage_5__778_, data_stage_5__777_, data_stage_5__776_, data_stage_5__775_, data_stage_5__774_, data_stage_5__773_, data_stage_5__772_, data_stage_5__771_, data_stage_5__770_, data_stage_5__769_, data_stage_5__768_, data_stage_5__767_, data_stage_5__766_, data_stage_5__765_, data_stage_5__764_, data_stage_5__763_, data_stage_5__762_, data_stage_5__761_, data_stage_5__760_, data_stage_5__759_, data_stage_5__758_, data_stage_5__757_, data_stage_5__756_, data_stage_5__755_, data_stage_5__754_, data_stage_5__753_, data_stage_5__752_, data_stage_5__751_, data_stage_5__750_, data_stage_5__749_, data_stage_5__748_, data_stage_5__747_, data_stage_5__746_, data_stage_5__745_, data_stage_5__744_, data_stage_5__743_, data_stage_5__742_, data_stage_5__741_, data_stage_5__740_, data_stage_5__739_, data_stage_5__738_, data_stage_5__737_, data_stage_5__736_, data_stage_5__735_, data_stage_5__734_, data_stage_5__733_, data_stage_5__732_, data_stage_5__731_, data_stage_5__730_, data_stage_5__729_, data_stage_5__728_, data_stage_5__727_, data_stage_5__726_, data_stage_5__725_, data_stage_5__724_, data_stage_5__723_, data_stage_5__722_, data_stage_5__721_, data_stage_5__720_, data_stage_5__719_, data_stage_5__718_, data_stage_5__717_, data_stage_5__716_, data_stage_5__715_, data_stage_5__714_, data_stage_5__713_, data_stage_5__712_, data_stage_5__711_, data_stage_5__710_, data_stage_5__709_, data_stage_5__708_, data_stage_5__707_, data_stage_5__706_, data_stage_5__705_, data_stage_5__704_, data_stage_5__703_, data_stage_5__702_, data_stage_5__701_, data_stage_5__700_, data_stage_5__699_, data_stage_5__698_, data_stage_5__697_, data_stage_5__696_, data_stage_5__695_, data_stage_5__694_, data_stage_5__693_, data_stage_5__692_, data_stage_5__691_, data_stage_5__690_, data_stage_5__689_, data_stage_5__688_, data_stage_5__687_, data_stage_5__686_, data_stage_5__685_, data_stage_5__684_, data_stage_5__683_, data_stage_5__682_, data_stage_5__681_, data_stage_5__680_, data_stage_5__679_, data_stage_5__678_, data_stage_5__677_, data_stage_5__676_, data_stage_5__675_, data_stage_5__674_, data_stage_5__673_, data_stage_5__672_, data_stage_5__671_, data_stage_5__670_, data_stage_5__669_, data_stage_5__668_, data_stage_5__667_, data_stage_5__666_, data_stage_5__665_, data_stage_5__664_, data_stage_5__663_, data_stage_5__662_, data_stage_5__661_, data_stage_5__660_, data_stage_5__659_, data_stage_5__658_, data_stage_5__657_, data_stage_5__656_, data_stage_5__655_, data_stage_5__654_, data_stage_5__653_, data_stage_5__652_, data_stage_5__651_, data_stage_5__650_, data_stage_5__649_, data_stage_5__648_, data_stage_5__647_, data_stage_5__646_, data_stage_5__645_, data_stage_5__644_, data_stage_5__643_, data_stage_5__642_, data_stage_5__641_, data_stage_5__640_, data_stage_5__639_, data_stage_5__638_, data_stage_5__637_, data_stage_5__636_, data_stage_5__635_, data_stage_5__634_, data_stage_5__633_, data_stage_5__632_, data_stage_5__631_, data_stage_5__630_, data_stage_5__629_, data_stage_5__628_, data_stage_5__627_, data_stage_5__626_, data_stage_5__625_, data_stage_5__624_, data_stage_5__623_, data_stage_5__622_, data_stage_5__621_, data_stage_5__620_, data_stage_5__619_, data_stage_5__618_, data_stage_5__617_, data_stage_5__616_, data_stage_5__615_, data_stage_5__614_, data_stage_5__613_, data_stage_5__612_, data_stage_5__611_, data_stage_5__610_, data_stage_5__609_, data_stage_5__608_, data_stage_5__607_, data_stage_5__606_, data_stage_5__605_, data_stage_5__604_, data_stage_5__603_, data_stage_5__602_, data_stage_5__601_, data_stage_5__600_, data_stage_5__599_, data_stage_5__598_, data_stage_5__597_, data_stage_5__596_, data_stage_5__595_, data_stage_5__594_, data_stage_5__593_, data_stage_5__592_, data_stage_5__591_, data_stage_5__590_, data_stage_5__589_, data_stage_5__588_, data_stage_5__587_, data_stage_5__586_, data_stage_5__585_, data_stage_5__584_, data_stage_5__583_, data_stage_5__582_, data_stage_5__581_, data_stage_5__580_, data_stage_5__579_, data_stage_5__578_, data_stage_5__577_, data_stage_5__576_, data_stage_5__575_, data_stage_5__574_, data_stage_5__573_, data_stage_5__572_, data_stage_5__571_, data_stage_5__570_, data_stage_5__569_, data_stage_5__568_, data_stage_5__567_, data_stage_5__566_, data_stage_5__565_, data_stage_5__564_, data_stage_5__563_, data_stage_5__562_, data_stage_5__561_, data_stage_5__560_, data_stage_5__559_, data_stage_5__558_, data_stage_5__557_, data_stage_5__556_, data_stage_5__555_, data_stage_5__554_, data_stage_5__553_, data_stage_5__552_, data_stage_5__551_, data_stage_5__550_, data_stage_5__549_, data_stage_5__548_, data_stage_5__547_, data_stage_5__546_, data_stage_5__545_, data_stage_5__544_, data_stage_5__543_, data_stage_5__542_, data_stage_5__541_, data_stage_5__540_, data_stage_5__539_, data_stage_5__538_, data_stage_5__537_, data_stage_5__536_, data_stage_5__535_, data_stage_5__534_, data_stage_5__533_, data_stage_5__532_, data_stage_5__531_, data_stage_5__530_, data_stage_5__529_, data_stage_5__528_, data_stage_5__527_, data_stage_5__526_, data_stage_5__525_, data_stage_5__524_, data_stage_5__523_, data_stage_5__522_, data_stage_5__521_, data_stage_5__520_, data_stage_5__519_, data_stage_5__518_, data_stage_5__517_, data_stage_5__516_, data_stage_5__515_, data_stage_5__514_, data_stage_5__513_, data_stage_5__512_, data_stage_5__511_, data_stage_5__510_, data_stage_5__509_, data_stage_5__508_, data_stage_5__507_, data_stage_5__506_, data_stage_5__505_, data_stage_5__504_, data_stage_5__503_, data_stage_5__502_, data_stage_5__501_, data_stage_5__500_, data_stage_5__499_, data_stage_5__498_, data_stage_5__497_, data_stage_5__496_, data_stage_5__495_, data_stage_5__494_, data_stage_5__493_, data_stage_5__492_, data_stage_5__491_, data_stage_5__490_, data_stage_5__489_, data_stage_5__488_, data_stage_5__487_, data_stage_5__486_, data_stage_5__485_, data_stage_5__484_, data_stage_5__483_, data_stage_5__482_, data_stage_5__481_, data_stage_5__480_, data_stage_5__479_, data_stage_5__478_, data_stage_5__477_, data_stage_5__476_, data_stage_5__475_, data_stage_5__474_, data_stage_5__473_, data_stage_5__472_, data_stage_5__471_, data_stage_5__470_, data_stage_5__469_, data_stage_5__468_, data_stage_5__467_, data_stage_5__466_, data_stage_5__465_, data_stage_5__464_, data_stage_5__463_, data_stage_5__462_, data_stage_5__461_, data_stage_5__460_, data_stage_5__459_, data_stage_5__458_, data_stage_5__457_, data_stage_5__456_, data_stage_5__455_, data_stage_5__454_, data_stage_5__453_, data_stage_5__452_, data_stage_5__451_, data_stage_5__450_, data_stage_5__449_, data_stage_5__448_, data_stage_5__447_, data_stage_5__446_, data_stage_5__445_, data_stage_5__444_, data_stage_5__443_, data_stage_5__442_, data_stage_5__441_, data_stage_5__440_, data_stage_5__439_, data_stage_5__438_, data_stage_5__437_, data_stage_5__436_, data_stage_5__435_, data_stage_5__434_, data_stage_5__433_, data_stage_5__432_, data_stage_5__431_, data_stage_5__430_, data_stage_5__429_, data_stage_5__428_, data_stage_5__427_, data_stage_5__426_, data_stage_5__425_, data_stage_5__424_, data_stage_5__423_, data_stage_5__422_, data_stage_5__421_, data_stage_5__420_, data_stage_5__419_, data_stage_5__418_, data_stage_5__417_, data_stage_5__416_, data_stage_5__415_, data_stage_5__414_, data_stage_5__413_, data_stage_5__412_, data_stage_5__411_, data_stage_5__410_, data_stage_5__409_, data_stage_5__408_, data_stage_5__407_, data_stage_5__406_, data_stage_5__405_, data_stage_5__404_, data_stage_5__403_, data_stage_5__402_, data_stage_5__401_, data_stage_5__400_, data_stage_5__399_, data_stage_5__398_, data_stage_5__397_, data_stage_5__396_, data_stage_5__395_, data_stage_5__394_, data_stage_5__393_, data_stage_5__392_, data_stage_5__391_, data_stage_5__390_, data_stage_5__389_, data_stage_5__388_, data_stage_5__387_, data_stage_5__386_, data_stage_5__385_, data_stage_5__384_, data_stage_5__383_, data_stage_5__382_, data_stage_5__381_, data_stage_5__380_, data_stage_5__379_, data_stage_5__378_, data_stage_5__377_, data_stage_5__376_, data_stage_5__375_, data_stage_5__374_, data_stage_5__373_, data_stage_5__372_, data_stage_5__371_, data_stage_5__370_, data_stage_5__369_, data_stage_5__368_, data_stage_5__367_, data_stage_5__366_, data_stage_5__365_, data_stage_5__364_, data_stage_5__363_, data_stage_5__362_, data_stage_5__361_, data_stage_5__360_, data_stage_5__359_, data_stage_5__358_, data_stage_5__357_, data_stage_5__356_, data_stage_5__355_, data_stage_5__354_, data_stage_5__353_, data_stage_5__352_, data_stage_5__351_, data_stage_5__350_, data_stage_5__349_, data_stage_5__348_, data_stage_5__347_, data_stage_5__346_, data_stage_5__345_, data_stage_5__344_, data_stage_5__343_, data_stage_5__342_, data_stage_5__341_, data_stage_5__340_, data_stage_5__339_, data_stage_5__338_, data_stage_5__337_, data_stage_5__336_, data_stage_5__335_, data_stage_5__334_, data_stage_5__333_, data_stage_5__332_, data_stage_5__331_, data_stage_5__330_, data_stage_5__329_, data_stage_5__328_, data_stage_5__327_, data_stage_5__326_, data_stage_5__325_, data_stage_5__324_, data_stage_5__323_, data_stage_5__322_, data_stage_5__321_, data_stage_5__320_, data_stage_5__319_, data_stage_5__318_, data_stage_5__317_, data_stage_5__316_, data_stage_5__315_, data_stage_5__314_, data_stage_5__313_, data_stage_5__312_, data_stage_5__311_, data_stage_5__310_, data_stage_5__309_, data_stage_5__308_, data_stage_5__307_, data_stage_5__306_, data_stage_5__305_, data_stage_5__304_, data_stage_5__303_, data_stage_5__302_, data_stage_5__301_, data_stage_5__300_, data_stage_5__299_, data_stage_5__298_, data_stage_5__297_, data_stage_5__296_, data_stage_5__295_, data_stage_5__294_, data_stage_5__293_, data_stage_5__292_, data_stage_5__291_, data_stage_5__290_, data_stage_5__289_, data_stage_5__288_, data_stage_5__287_, data_stage_5__286_, data_stage_5__285_, data_stage_5__284_, data_stage_5__283_, data_stage_5__282_, data_stage_5__281_, data_stage_5__280_, data_stage_5__279_, data_stage_5__278_, data_stage_5__277_, data_stage_5__276_, data_stage_5__275_, data_stage_5__274_, data_stage_5__273_, data_stage_5__272_, data_stage_5__271_, data_stage_5__270_, data_stage_5__269_, data_stage_5__268_, data_stage_5__267_, data_stage_5__266_, data_stage_5__265_, data_stage_5__264_, data_stage_5__263_, data_stage_5__262_, data_stage_5__261_, data_stage_5__260_, data_stage_5__259_, data_stage_5__258_, data_stage_5__257_, data_stage_5__256_, data_stage_5__255_, data_stage_5__254_, data_stage_5__253_, data_stage_5__252_, data_stage_5__251_, data_stage_5__250_, data_stage_5__249_, data_stage_5__248_, data_stage_5__247_, data_stage_5__246_, data_stage_5__245_, data_stage_5__244_, data_stage_5__243_, data_stage_5__242_, data_stage_5__241_, data_stage_5__240_, data_stage_5__239_, data_stage_5__238_, data_stage_5__237_, data_stage_5__236_, data_stage_5__235_, data_stage_5__234_, data_stage_5__233_, data_stage_5__232_, data_stage_5__231_, data_stage_5__230_, data_stage_5__229_, data_stage_5__228_, data_stage_5__227_, data_stage_5__226_, data_stage_5__225_, data_stage_5__224_, data_stage_5__223_, data_stage_5__222_, data_stage_5__221_, data_stage_5__220_, data_stage_5__219_, data_stage_5__218_, data_stage_5__217_, data_stage_5__216_, data_stage_5__215_, data_stage_5__214_, data_stage_5__213_, data_stage_5__212_, data_stage_5__211_, data_stage_5__210_, data_stage_5__209_, data_stage_5__208_, data_stage_5__207_, data_stage_5__206_, data_stage_5__205_, data_stage_5__204_, data_stage_5__203_, data_stage_5__202_, data_stage_5__201_, data_stage_5__200_, data_stage_5__199_, data_stage_5__198_, data_stage_5__197_, data_stage_5__196_, data_stage_5__195_, data_stage_5__194_, data_stage_5__193_, data_stage_5__192_, data_stage_5__191_, data_stage_5__190_, data_stage_5__189_, data_stage_5__188_, data_stage_5__187_, data_stage_5__186_, data_stage_5__185_, data_stage_5__184_, data_stage_5__183_, data_stage_5__182_, data_stage_5__181_, data_stage_5__180_, data_stage_5__179_, data_stage_5__178_, data_stage_5__177_, data_stage_5__176_, data_stage_5__175_, data_stage_5__174_, data_stage_5__173_, data_stage_5__172_, data_stage_5__171_, data_stage_5__170_, data_stage_5__169_, data_stage_5__168_, data_stage_5__167_, data_stage_5__166_, data_stage_5__165_, data_stage_5__164_, data_stage_5__163_, data_stage_5__162_, data_stage_5__161_, data_stage_5__160_, data_stage_5__159_, data_stage_5__158_, data_stage_5__157_, data_stage_5__156_, data_stage_5__155_, data_stage_5__154_, data_stage_5__153_, data_stage_5__152_, data_stage_5__151_, data_stage_5__150_, data_stage_5__149_, data_stage_5__148_, data_stage_5__147_, data_stage_5__146_, data_stage_5__145_, data_stage_5__144_, data_stage_5__143_, data_stage_5__142_, data_stage_5__141_, data_stage_5__140_, data_stage_5__139_, data_stage_5__138_, data_stage_5__137_, data_stage_5__136_, data_stage_5__135_, data_stage_5__134_, data_stage_5__133_, data_stage_5__132_, data_stage_5__131_, data_stage_5__130_, data_stage_5__129_, data_stage_5__128_, data_stage_5__127_, data_stage_5__126_, data_stage_5__125_, data_stage_5__124_, data_stage_5__123_, data_stage_5__122_, data_stage_5__121_, data_stage_5__120_, data_stage_5__119_, data_stage_5__118_, data_stage_5__117_, data_stage_5__116_, data_stage_5__115_, data_stage_5__114_, data_stage_5__113_, data_stage_5__112_, data_stage_5__111_, data_stage_5__110_, data_stage_5__109_, data_stage_5__108_, data_stage_5__107_, data_stage_5__106_, data_stage_5__105_, data_stage_5__104_, data_stage_5__103_, data_stage_5__102_, data_stage_5__101_, data_stage_5__100_, data_stage_5__99_, data_stage_5__98_, data_stage_5__97_, data_stage_5__96_, data_stage_5__95_, data_stage_5__94_, data_stage_5__93_, data_stage_5__92_, data_stage_5__91_, data_stage_5__90_, data_stage_5__89_, data_stage_5__88_, data_stage_5__87_, data_stage_5__86_, data_stage_5__85_, data_stage_5__84_, data_stage_5__83_, data_stage_5__82_, data_stage_5__81_, data_stage_5__80_, data_stage_5__79_, data_stage_5__78_, data_stage_5__77_, data_stage_5__76_, data_stage_5__75_, data_stage_5__74_, data_stage_5__73_, data_stage_5__72_, data_stage_5__71_, data_stage_5__70_, data_stage_5__69_, data_stage_5__68_, data_stage_5__67_, data_stage_5__66_, data_stage_5__65_, data_stage_5__64_, data_stage_5__63_, data_stage_5__62_, data_stage_5__61_, data_stage_5__60_, data_stage_5__59_, data_stage_5__58_, data_stage_5__57_, data_stage_5__56_, data_stage_5__55_, data_stage_5__54_, data_stage_5__53_, data_stage_5__52_, data_stage_5__51_, data_stage_5__50_, data_stage_5__49_, data_stage_5__48_, data_stage_5__47_, data_stage_5__46_, data_stage_5__45_, data_stage_5__44_, data_stage_5__43_, data_stage_5__42_, data_stage_5__41_, data_stage_5__40_, data_stage_5__39_, data_stage_5__38_, data_stage_5__37_, data_stage_5__36_, data_stage_5__35_, data_stage_5__34_, data_stage_5__33_, data_stage_5__32_, data_stage_5__31_, data_stage_5__30_, data_stage_5__29_, data_stage_5__28_, data_stage_5__27_, data_stage_5__26_, data_stage_5__25_, data_stage_5__24_, data_stage_5__23_, data_stage_5__22_, data_stage_5__21_, data_stage_5__20_, data_stage_5__19_, data_stage_5__18_, data_stage_5__17_, data_stage_5__16_, data_stage_5__15_, data_stage_5__14_, data_stage_5__13_, data_stage_5__12_, data_stage_5__11_, data_stage_5__10_, data_stage_5__9_, data_stage_5__8_, data_stage_5__7_, data_stage_5__6_, data_stage_5__5_, data_stage_5__4_, data_stage_5__3_, data_stage_5__2_, data_stage_5__1_, data_stage_5__0_ })
  );


  bsg_swap_width_p2048
  mux_stage_4__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_4__8191_, data_stage_4__8190_, data_stage_4__8189_, data_stage_4__8188_, data_stage_4__8187_, data_stage_4__8186_, data_stage_4__8185_, data_stage_4__8184_, data_stage_4__8183_, data_stage_4__8182_, data_stage_4__8181_, data_stage_4__8180_, data_stage_4__8179_, data_stage_4__8178_, data_stage_4__8177_, data_stage_4__8176_, data_stage_4__8175_, data_stage_4__8174_, data_stage_4__8173_, data_stage_4__8172_, data_stage_4__8171_, data_stage_4__8170_, data_stage_4__8169_, data_stage_4__8168_, data_stage_4__8167_, data_stage_4__8166_, data_stage_4__8165_, data_stage_4__8164_, data_stage_4__8163_, data_stage_4__8162_, data_stage_4__8161_, data_stage_4__8160_, data_stage_4__8159_, data_stage_4__8158_, data_stage_4__8157_, data_stage_4__8156_, data_stage_4__8155_, data_stage_4__8154_, data_stage_4__8153_, data_stage_4__8152_, data_stage_4__8151_, data_stage_4__8150_, data_stage_4__8149_, data_stage_4__8148_, data_stage_4__8147_, data_stage_4__8146_, data_stage_4__8145_, data_stage_4__8144_, data_stage_4__8143_, data_stage_4__8142_, data_stage_4__8141_, data_stage_4__8140_, data_stage_4__8139_, data_stage_4__8138_, data_stage_4__8137_, data_stage_4__8136_, data_stage_4__8135_, data_stage_4__8134_, data_stage_4__8133_, data_stage_4__8132_, data_stage_4__8131_, data_stage_4__8130_, data_stage_4__8129_, data_stage_4__8128_, data_stage_4__8127_, data_stage_4__8126_, data_stage_4__8125_, data_stage_4__8124_, data_stage_4__8123_, data_stage_4__8122_, data_stage_4__8121_, data_stage_4__8120_, data_stage_4__8119_, data_stage_4__8118_, data_stage_4__8117_, data_stage_4__8116_, data_stage_4__8115_, data_stage_4__8114_, data_stage_4__8113_, data_stage_4__8112_, data_stage_4__8111_, data_stage_4__8110_, data_stage_4__8109_, data_stage_4__8108_, data_stage_4__8107_, data_stage_4__8106_, data_stage_4__8105_, data_stage_4__8104_, data_stage_4__8103_, data_stage_4__8102_, data_stage_4__8101_, data_stage_4__8100_, data_stage_4__8099_, data_stage_4__8098_, data_stage_4__8097_, data_stage_4__8096_, data_stage_4__8095_, data_stage_4__8094_, data_stage_4__8093_, data_stage_4__8092_, data_stage_4__8091_, data_stage_4__8090_, data_stage_4__8089_, data_stage_4__8088_, data_stage_4__8087_, data_stage_4__8086_, data_stage_4__8085_, data_stage_4__8084_, data_stage_4__8083_, data_stage_4__8082_, data_stage_4__8081_, data_stage_4__8080_, data_stage_4__8079_, data_stage_4__8078_, data_stage_4__8077_, data_stage_4__8076_, data_stage_4__8075_, data_stage_4__8074_, data_stage_4__8073_, data_stage_4__8072_, data_stage_4__8071_, data_stage_4__8070_, data_stage_4__8069_, data_stage_4__8068_, data_stage_4__8067_, data_stage_4__8066_, data_stage_4__8065_, data_stage_4__8064_, data_stage_4__8063_, data_stage_4__8062_, data_stage_4__8061_, data_stage_4__8060_, data_stage_4__8059_, data_stage_4__8058_, data_stage_4__8057_, data_stage_4__8056_, data_stage_4__8055_, data_stage_4__8054_, data_stage_4__8053_, data_stage_4__8052_, data_stage_4__8051_, data_stage_4__8050_, data_stage_4__8049_, data_stage_4__8048_, data_stage_4__8047_, data_stage_4__8046_, data_stage_4__8045_, data_stage_4__8044_, data_stage_4__8043_, data_stage_4__8042_, data_stage_4__8041_, data_stage_4__8040_, data_stage_4__8039_, data_stage_4__8038_, data_stage_4__8037_, data_stage_4__8036_, data_stage_4__8035_, data_stage_4__8034_, data_stage_4__8033_, data_stage_4__8032_, data_stage_4__8031_, data_stage_4__8030_, data_stage_4__8029_, data_stage_4__8028_, data_stage_4__8027_, data_stage_4__8026_, data_stage_4__8025_, data_stage_4__8024_, data_stage_4__8023_, data_stage_4__8022_, data_stage_4__8021_, data_stage_4__8020_, data_stage_4__8019_, data_stage_4__8018_, data_stage_4__8017_, data_stage_4__8016_, data_stage_4__8015_, data_stage_4__8014_, data_stage_4__8013_, data_stage_4__8012_, data_stage_4__8011_, data_stage_4__8010_, data_stage_4__8009_, data_stage_4__8008_, data_stage_4__8007_, data_stage_4__8006_, data_stage_4__8005_, data_stage_4__8004_, data_stage_4__8003_, data_stage_4__8002_, data_stage_4__8001_, data_stage_4__8000_, data_stage_4__7999_, data_stage_4__7998_, data_stage_4__7997_, data_stage_4__7996_, data_stage_4__7995_, data_stage_4__7994_, data_stage_4__7993_, data_stage_4__7992_, data_stage_4__7991_, data_stage_4__7990_, data_stage_4__7989_, data_stage_4__7988_, data_stage_4__7987_, data_stage_4__7986_, data_stage_4__7985_, data_stage_4__7984_, data_stage_4__7983_, data_stage_4__7982_, data_stage_4__7981_, data_stage_4__7980_, data_stage_4__7979_, data_stage_4__7978_, data_stage_4__7977_, data_stage_4__7976_, data_stage_4__7975_, data_stage_4__7974_, data_stage_4__7973_, data_stage_4__7972_, data_stage_4__7971_, data_stage_4__7970_, data_stage_4__7969_, data_stage_4__7968_, data_stage_4__7967_, data_stage_4__7966_, data_stage_4__7965_, data_stage_4__7964_, data_stage_4__7963_, data_stage_4__7962_, data_stage_4__7961_, data_stage_4__7960_, data_stage_4__7959_, data_stage_4__7958_, data_stage_4__7957_, data_stage_4__7956_, data_stage_4__7955_, data_stage_4__7954_, data_stage_4__7953_, data_stage_4__7952_, data_stage_4__7951_, data_stage_4__7950_, data_stage_4__7949_, data_stage_4__7948_, data_stage_4__7947_, data_stage_4__7946_, data_stage_4__7945_, data_stage_4__7944_, data_stage_4__7943_, data_stage_4__7942_, data_stage_4__7941_, data_stage_4__7940_, data_stage_4__7939_, data_stage_4__7938_, data_stage_4__7937_, data_stage_4__7936_, data_stage_4__7935_, data_stage_4__7934_, data_stage_4__7933_, data_stage_4__7932_, data_stage_4__7931_, data_stage_4__7930_, data_stage_4__7929_, data_stage_4__7928_, data_stage_4__7927_, data_stage_4__7926_, data_stage_4__7925_, data_stage_4__7924_, data_stage_4__7923_, data_stage_4__7922_, data_stage_4__7921_, data_stage_4__7920_, data_stage_4__7919_, data_stage_4__7918_, data_stage_4__7917_, data_stage_4__7916_, data_stage_4__7915_, data_stage_4__7914_, data_stage_4__7913_, data_stage_4__7912_, data_stage_4__7911_, data_stage_4__7910_, data_stage_4__7909_, data_stage_4__7908_, data_stage_4__7907_, data_stage_4__7906_, data_stage_4__7905_, data_stage_4__7904_, data_stage_4__7903_, data_stage_4__7902_, data_stage_4__7901_, data_stage_4__7900_, data_stage_4__7899_, data_stage_4__7898_, data_stage_4__7897_, data_stage_4__7896_, data_stage_4__7895_, data_stage_4__7894_, data_stage_4__7893_, data_stage_4__7892_, data_stage_4__7891_, data_stage_4__7890_, data_stage_4__7889_, data_stage_4__7888_, data_stage_4__7887_, data_stage_4__7886_, data_stage_4__7885_, data_stage_4__7884_, data_stage_4__7883_, data_stage_4__7882_, data_stage_4__7881_, data_stage_4__7880_, data_stage_4__7879_, data_stage_4__7878_, data_stage_4__7877_, data_stage_4__7876_, data_stage_4__7875_, data_stage_4__7874_, data_stage_4__7873_, data_stage_4__7872_, data_stage_4__7871_, data_stage_4__7870_, data_stage_4__7869_, data_stage_4__7868_, data_stage_4__7867_, data_stage_4__7866_, data_stage_4__7865_, data_stage_4__7864_, data_stage_4__7863_, data_stage_4__7862_, data_stage_4__7861_, data_stage_4__7860_, data_stage_4__7859_, data_stage_4__7858_, data_stage_4__7857_, data_stage_4__7856_, data_stage_4__7855_, data_stage_4__7854_, data_stage_4__7853_, data_stage_4__7852_, data_stage_4__7851_, data_stage_4__7850_, data_stage_4__7849_, data_stage_4__7848_, data_stage_4__7847_, data_stage_4__7846_, data_stage_4__7845_, data_stage_4__7844_, data_stage_4__7843_, data_stage_4__7842_, data_stage_4__7841_, data_stage_4__7840_, data_stage_4__7839_, data_stage_4__7838_, data_stage_4__7837_, data_stage_4__7836_, data_stage_4__7835_, data_stage_4__7834_, data_stage_4__7833_, data_stage_4__7832_, data_stage_4__7831_, data_stage_4__7830_, data_stage_4__7829_, data_stage_4__7828_, data_stage_4__7827_, data_stage_4__7826_, data_stage_4__7825_, data_stage_4__7824_, data_stage_4__7823_, data_stage_4__7822_, data_stage_4__7821_, data_stage_4__7820_, data_stage_4__7819_, data_stage_4__7818_, data_stage_4__7817_, data_stage_4__7816_, data_stage_4__7815_, data_stage_4__7814_, data_stage_4__7813_, data_stage_4__7812_, data_stage_4__7811_, data_stage_4__7810_, data_stage_4__7809_, data_stage_4__7808_, data_stage_4__7807_, data_stage_4__7806_, data_stage_4__7805_, data_stage_4__7804_, data_stage_4__7803_, data_stage_4__7802_, data_stage_4__7801_, data_stage_4__7800_, data_stage_4__7799_, data_stage_4__7798_, data_stage_4__7797_, data_stage_4__7796_, data_stage_4__7795_, data_stage_4__7794_, data_stage_4__7793_, data_stage_4__7792_, data_stage_4__7791_, data_stage_4__7790_, data_stage_4__7789_, data_stage_4__7788_, data_stage_4__7787_, data_stage_4__7786_, data_stage_4__7785_, data_stage_4__7784_, data_stage_4__7783_, data_stage_4__7782_, data_stage_4__7781_, data_stage_4__7780_, data_stage_4__7779_, data_stage_4__7778_, data_stage_4__7777_, data_stage_4__7776_, data_stage_4__7775_, data_stage_4__7774_, data_stage_4__7773_, data_stage_4__7772_, data_stage_4__7771_, data_stage_4__7770_, data_stage_4__7769_, data_stage_4__7768_, data_stage_4__7767_, data_stage_4__7766_, data_stage_4__7765_, data_stage_4__7764_, data_stage_4__7763_, data_stage_4__7762_, data_stage_4__7761_, data_stage_4__7760_, data_stage_4__7759_, data_stage_4__7758_, data_stage_4__7757_, data_stage_4__7756_, data_stage_4__7755_, data_stage_4__7754_, data_stage_4__7753_, data_stage_4__7752_, data_stage_4__7751_, data_stage_4__7750_, data_stage_4__7749_, data_stage_4__7748_, data_stage_4__7747_, data_stage_4__7746_, data_stage_4__7745_, data_stage_4__7744_, data_stage_4__7743_, data_stage_4__7742_, data_stage_4__7741_, data_stage_4__7740_, data_stage_4__7739_, data_stage_4__7738_, data_stage_4__7737_, data_stage_4__7736_, data_stage_4__7735_, data_stage_4__7734_, data_stage_4__7733_, data_stage_4__7732_, data_stage_4__7731_, data_stage_4__7730_, data_stage_4__7729_, data_stage_4__7728_, data_stage_4__7727_, data_stage_4__7726_, data_stage_4__7725_, data_stage_4__7724_, data_stage_4__7723_, data_stage_4__7722_, data_stage_4__7721_, data_stage_4__7720_, data_stage_4__7719_, data_stage_4__7718_, data_stage_4__7717_, data_stage_4__7716_, data_stage_4__7715_, data_stage_4__7714_, data_stage_4__7713_, data_stage_4__7712_, data_stage_4__7711_, data_stage_4__7710_, data_stage_4__7709_, data_stage_4__7708_, data_stage_4__7707_, data_stage_4__7706_, data_stage_4__7705_, data_stage_4__7704_, data_stage_4__7703_, data_stage_4__7702_, data_stage_4__7701_, data_stage_4__7700_, data_stage_4__7699_, data_stage_4__7698_, data_stage_4__7697_, data_stage_4__7696_, data_stage_4__7695_, data_stage_4__7694_, data_stage_4__7693_, data_stage_4__7692_, data_stage_4__7691_, data_stage_4__7690_, data_stage_4__7689_, data_stage_4__7688_, data_stage_4__7687_, data_stage_4__7686_, data_stage_4__7685_, data_stage_4__7684_, data_stage_4__7683_, data_stage_4__7682_, data_stage_4__7681_, data_stage_4__7680_, data_stage_4__7679_, data_stage_4__7678_, data_stage_4__7677_, data_stage_4__7676_, data_stage_4__7675_, data_stage_4__7674_, data_stage_4__7673_, data_stage_4__7672_, data_stage_4__7671_, data_stage_4__7670_, data_stage_4__7669_, data_stage_4__7668_, data_stage_4__7667_, data_stage_4__7666_, data_stage_4__7665_, data_stage_4__7664_, data_stage_4__7663_, data_stage_4__7662_, data_stage_4__7661_, data_stage_4__7660_, data_stage_4__7659_, data_stage_4__7658_, data_stage_4__7657_, data_stage_4__7656_, data_stage_4__7655_, data_stage_4__7654_, data_stage_4__7653_, data_stage_4__7652_, data_stage_4__7651_, data_stage_4__7650_, data_stage_4__7649_, data_stage_4__7648_, data_stage_4__7647_, data_stage_4__7646_, data_stage_4__7645_, data_stage_4__7644_, data_stage_4__7643_, data_stage_4__7642_, data_stage_4__7641_, data_stage_4__7640_, data_stage_4__7639_, data_stage_4__7638_, data_stage_4__7637_, data_stage_4__7636_, data_stage_4__7635_, data_stage_4__7634_, data_stage_4__7633_, data_stage_4__7632_, data_stage_4__7631_, data_stage_4__7630_, data_stage_4__7629_, data_stage_4__7628_, data_stage_4__7627_, data_stage_4__7626_, data_stage_4__7625_, data_stage_4__7624_, data_stage_4__7623_, data_stage_4__7622_, data_stage_4__7621_, data_stage_4__7620_, data_stage_4__7619_, data_stage_4__7618_, data_stage_4__7617_, data_stage_4__7616_, data_stage_4__7615_, data_stage_4__7614_, data_stage_4__7613_, data_stage_4__7612_, data_stage_4__7611_, data_stage_4__7610_, data_stage_4__7609_, data_stage_4__7608_, data_stage_4__7607_, data_stage_4__7606_, data_stage_4__7605_, data_stage_4__7604_, data_stage_4__7603_, data_stage_4__7602_, data_stage_4__7601_, data_stage_4__7600_, data_stage_4__7599_, data_stage_4__7598_, data_stage_4__7597_, data_stage_4__7596_, data_stage_4__7595_, data_stage_4__7594_, data_stage_4__7593_, data_stage_4__7592_, data_stage_4__7591_, data_stage_4__7590_, data_stage_4__7589_, data_stage_4__7588_, data_stage_4__7587_, data_stage_4__7586_, data_stage_4__7585_, data_stage_4__7584_, data_stage_4__7583_, data_stage_4__7582_, data_stage_4__7581_, data_stage_4__7580_, data_stage_4__7579_, data_stage_4__7578_, data_stage_4__7577_, data_stage_4__7576_, data_stage_4__7575_, data_stage_4__7574_, data_stage_4__7573_, data_stage_4__7572_, data_stage_4__7571_, data_stage_4__7570_, data_stage_4__7569_, data_stage_4__7568_, data_stage_4__7567_, data_stage_4__7566_, data_stage_4__7565_, data_stage_4__7564_, data_stage_4__7563_, data_stage_4__7562_, data_stage_4__7561_, data_stage_4__7560_, data_stage_4__7559_, data_stage_4__7558_, data_stage_4__7557_, data_stage_4__7556_, data_stage_4__7555_, data_stage_4__7554_, data_stage_4__7553_, data_stage_4__7552_, data_stage_4__7551_, data_stage_4__7550_, data_stage_4__7549_, data_stage_4__7548_, data_stage_4__7547_, data_stage_4__7546_, data_stage_4__7545_, data_stage_4__7544_, data_stage_4__7543_, data_stage_4__7542_, data_stage_4__7541_, data_stage_4__7540_, data_stage_4__7539_, data_stage_4__7538_, data_stage_4__7537_, data_stage_4__7536_, data_stage_4__7535_, data_stage_4__7534_, data_stage_4__7533_, data_stage_4__7532_, data_stage_4__7531_, data_stage_4__7530_, data_stage_4__7529_, data_stage_4__7528_, data_stage_4__7527_, data_stage_4__7526_, data_stage_4__7525_, data_stage_4__7524_, data_stage_4__7523_, data_stage_4__7522_, data_stage_4__7521_, data_stage_4__7520_, data_stage_4__7519_, data_stage_4__7518_, data_stage_4__7517_, data_stage_4__7516_, data_stage_4__7515_, data_stage_4__7514_, data_stage_4__7513_, data_stage_4__7512_, data_stage_4__7511_, data_stage_4__7510_, data_stage_4__7509_, data_stage_4__7508_, data_stage_4__7507_, data_stage_4__7506_, data_stage_4__7505_, data_stage_4__7504_, data_stage_4__7503_, data_stage_4__7502_, data_stage_4__7501_, data_stage_4__7500_, data_stage_4__7499_, data_stage_4__7498_, data_stage_4__7497_, data_stage_4__7496_, data_stage_4__7495_, data_stage_4__7494_, data_stage_4__7493_, data_stage_4__7492_, data_stage_4__7491_, data_stage_4__7490_, data_stage_4__7489_, data_stage_4__7488_, data_stage_4__7487_, data_stage_4__7486_, data_stage_4__7485_, data_stage_4__7484_, data_stage_4__7483_, data_stage_4__7482_, data_stage_4__7481_, data_stage_4__7480_, data_stage_4__7479_, data_stage_4__7478_, data_stage_4__7477_, data_stage_4__7476_, data_stage_4__7475_, data_stage_4__7474_, data_stage_4__7473_, data_stage_4__7472_, data_stage_4__7471_, data_stage_4__7470_, data_stage_4__7469_, data_stage_4__7468_, data_stage_4__7467_, data_stage_4__7466_, data_stage_4__7465_, data_stage_4__7464_, data_stage_4__7463_, data_stage_4__7462_, data_stage_4__7461_, data_stage_4__7460_, data_stage_4__7459_, data_stage_4__7458_, data_stage_4__7457_, data_stage_4__7456_, data_stage_4__7455_, data_stage_4__7454_, data_stage_4__7453_, data_stage_4__7452_, data_stage_4__7451_, data_stage_4__7450_, data_stage_4__7449_, data_stage_4__7448_, data_stage_4__7447_, data_stage_4__7446_, data_stage_4__7445_, data_stage_4__7444_, data_stage_4__7443_, data_stage_4__7442_, data_stage_4__7441_, data_stage_4__7440_, data_stage_4__7439_, data_stage_4__7438_, data_stage_4__7437_, data_stage_4__7436_, data_stage_4__7435_, data_stage_4__7434_, data_stage_4__7433_, data_stage_4__7432_, data_stage_4__7431_, data_stage_4__7430_, data_stage_4__7429_, data_stage_4__7428_, data_stage_4__7427_, data_stage_4__7426_, data_stage_4__7425_, data_stage_4__7424_, data_stage_4__7423_, data_stage_4__7422_, data_stage_4__7421_, data_stage_4__7420_, data_stage_4__7419_, data_stage_4__7418_, data_stage_4__7417_, data_stage_4__7416_, data_stage_4__7415_, data_stage_4__7414_, data_stage_4__7413_, data_stage_4__7412_, data_stage_4__7411_, data_stage_4__7410_, data_stage_4__7409_, data_stage_4__7408_, data_stage_4__7407_, data_stage_4__7406_, data_stage_4__7405_, data_stage_4__7404_, data_stage_4__7403_, data_stage_4__7402_, data_stage_4__7401_, data_stage_4__7400_, data_stage_4__7399_, data_stage_4__7398_, data_stage_4__7397_, data_stage_4__7396_, data_stage_4__7395_, data_stage_4__7394_, data_stage_4__7393_, data_stage_4__7392_, data_stage_4__7391_, data_stage_4__7390_, data_stage_4__7389_, data_stage_4__7388_, data_stage_4__7387_, data_stage_4__7386_, data_stage_4__7385_, data_stage_4__7384_, data_stage_4__7383_, data_stage_4__7382_, data_stage_4__7381_, data_stage_4__7380_, data_stage_4__7379_, data_stage_4__7378_, data_stage_4__7377_, data_stage_4__7376_, data_stage_4__7375_, data_stage_4__7374_, data_stage_4__7373_, data_stage_4__7372_, data_stage_4__7371_, data_stage_4__7370_, data_stage_4__7369_, data_stage_4__7368_, data_stage_4__7367_, data_stage_4__7366_, data_stage_4__7365_, data_stage_4__7364_, data_stage_4__7363_, data_stage_4__7362_, data_stage_4__7361_, data_stage_4__7360_, data_stage_4__7359_, data_stage_4__7358_, data_stage_4__7357_, data_stage_4__7356_, data_stage_4__7355_, data_stage_4__7354_, data_stage_4__7353_, data_stage_4__7352_, data_stage_4__7351_, data_stage_4__7350_, data_stage_4__7349_, data_stage_4__7348_, data_stage_4__7347_, data_stage_4__7346_, data_stage_4__7345_, data_stage_4__7344_, data_stage_4__7343_, data_stage_4__7342_, data_stage_4__7341_, data_stage_4__7340_, data_stage_4__7339_, data_stage_4__7338_, data_stage_4__7337_, data_stage_4__7336_, data_stage_4__7335_, data_stage_4__7334_, data_stage_4__7333_, data_stage_4__7332_, data_stage_4__7331_, data_stage_4__7330_, data_stage_4__7329_, data_stage_4__7328_, data_stage_4__7327_, data_stage_4__7326_, data_stage_4__7325_, data_stage_4__7324_, data_stage_4__7323_, data_stage_4__7322_, data_stage_4__7321_, data_stage_4__7320_, data_stage_4__7319_, data_stage_4__7318_, data_stage_4__7317_, data_stage_4__7316_, data_stage_4__7315_, data_stage_4__7314_, data_stage_4__7313_, data_stage_4__7312_, data_stage_4__7311_, data_stage_4__7310_, data_stage_4__7309_, data_stage_4__7308_, data_stage_4__7307_, data_stage_4__7306_, data_stage_4__7305_, data_stage_4__7304_, data_stage_4__7303_, data_stage_4__7302_, data_stage_4__7301_, data_stage_4__7300_, data_stage_4__7299_, data_stage_4__7298_, data_stage_4__7297_, data_stage_4__7296_, data_stage_4__7295_, data_stage_4__7294_, data_stage_4__7293_, data_stage_4__7292_, data_stage_4__7291_, data_stage_4__7290_, data_stage_4__7289_, data_stage_4__7288_, data_stage_4__7287_, data_stage_4__7286_, data_stage_4__7285_, data_stage_4__7284_, data_stage_4__7283_, data_stage_4__7282_, data_stage_4__7281_, data_stage_4__7280_, data_stage_4__7279_, data_stage_4__7278_, data_stage_4__7277_, data_stage_4__7276_, data_stage_4__7275_, data_stage_4__7274_, data_stage_4__7273_, data_stage_4__7272_, data_stage_4__7271_, data_stage_4__7270_, data_stage_4__7269_, data_stage_4__7268_, data_stage_4__7267_, data_stage_4__7266_, data_stage_4__7265_, data_stage_4__7264_, data_stage_4__7263_, data_stage_4__7262_, data_stage_4__7261_, data_stage_4__7260_, data_stage_4__7259_, data_stage_4__7258_, data_stage_4__7257_, data_stage_4__7256_, data_stage_4__7255_, data_stage_4__7254_, data_stage_4__7253_, data_stage_4__7252_, data_stage_4__7251_, data_stage_4__7250_, data_stage_4__7249_, data_stage_4__7248_, data_stage_4__7247_, data_stage_4__7246_, data_stage_4__7245_, data_stage_4__7244_, data_stage_4__7243_, data_stage_4__7242_, data_stage_4__7241_, data_stage_4__7240_, data_stage_4__7239_, data_stage_4__7238_, data_stage_4__7237_, data_stage_4__7236_, data_stage_4__7235_, data_stage_4__7234_, data_stage_4__7233_, data_stage_4__7232_, data_stage_4__7231_, data_stage_4__7230_, data_stage_4__7229_, data_stage_4__7228_, data_stage_4__7227_, data_stage_4__7226_, data_stage_4__7225_, data_stage_4__7224_, data_stage_4__7223_, data_stage_4__7222_, data_stage_4__7221_, data_stage_4__7220_, data_stage_4__7219_, data_stage_4__7218_, data_stage_4__7217_, data_stage_4__7216_, data_stage_4__7215_, data_stage_4__7214_, data_stage_4__7213_, data_stage_4__7212_, data_stage_4__7211_, data_stage_4__7210_, data_stage_4__7209_, data_stage_4__7208_, data_stage_4__7207_, data_stage_4__7206_, data_stage_4__7205_, data_stage_4__7204_, data_stage_4__7203_, data_stage_4__7202_, data_stage_4__7201_, data_stage_4__7200_, data_stage_4__7199_, data_stage_4__7198_, data_stage_4__7197_, data_stage_4__7196_, data_stage_4__7195_, data_stage_4__7194_, data_stage_4__7193_, data_stage_4__7192_, data_stage_4__7191_, data_stage_4__7190_, data_stage_4__7189_, data_stage_4__7188_, data_stage_4__7187_, data_stage_4__7186_, data_stage_4__7185_, data_stage_4__7184_, data_stage_4__7183_, data_stage_4__7182_, data_stage_4__7181_, data_stage_4__7180_, data_stage_4__7179_, data_stage_4__7178_, data_stage_4__7177_, data_stage_4__7176_, data_stage_4__7175_, data_stage_4__7174_, data_stage_4__7173_, data_stage_4__7172_, data_stage_4__7171_, data_stage_4__7170_, data_stage_4__7169_, data_stage_4__7168_, data_stage_4__7167_, data_stage_4__7166_, data_stage_4__7165_, data_stage_4__7164_, data_stage_4__7163_, data_stage_4__7162_, data_stage_4__7161_, data_stage_4__7160_, data_stage_4__7159_, data_stage_4__7158_, data_stage_4__7157_, data_stage_4__7156_, data_stage_4__7155_, data_stage_4__7154_, data_stage_4__7153_, data_stage_4__7152_, data_stage_4__7151_, data_stage_4__7150_, data_stage_4__7149_, data_stage_4__7148_, data_stage_4__7147_, data_stage_4__7146_, data_stage_4__7145_, data_stage_4__7144_, data_stage_4__7143_, data_stage_4__7142_, data_stage_4__7141_, data_stage_4__7140_, data_stage_4__7139_, data_stage_4__7138_, data_stage_4__7137_, data_stage_4__7136_, data_stage_4__7135_, data_stage_4__7134_, data_stage_4__7133_, data_stage_4__7132_, data_stage_4__7131_, data_stage_4__7130_, data_stage_4__7129_, data_stage_4__7128_, data_stage_4__7127_, data_stage_4__7126_, data_stage_4__7125_, data_stage_4__7124_, data_stage_4__7123_, data_stage_4__7122_, data_stage_4__7121_, data_stage_4__7120_, data_stage_4__7119_, data_stage_4__7118_, data_stage_4__7117_, data_stage_4__7116_, data_stage_4__7115_, data_stage_4__7114_, data_stage_4__7113_, data_stage_4__7112_, data_stage_4__7111_, data_stage_4__7110_, data_stage_4__7109_, data_stage_4__7108_, data_stage_4__7107_, data_stage_4__7106_, data_stage_4__7105_, data_stage_4__7104_, data_stage_4__7103_, data_stage_4__7102_, data_stage_4__7101_, data_stage_4__7100_, data_stage_4__7099_, data_stage_4__7098_, data_stage_4__7097_, data_stage_4__7096_, data_stage_4__7095_, data_stage_4__7094_, data_stage_4__7093_, data_stage_4__7092_, data_stage_4__7091_, data_stage_4__7090_, data_stage_4__7089_, data_stage_4__7088_, data_stage_4__7087_, data_stage_4__7086_, data_stage_4__7085_, data_stage_4__7084_, data_stage_4__7083_, data_stage_4__7082_, data_stage_4__7081_, data_stage_4__7080_, data_stage_4__7079_, data_stage_4__7078_, data_stage_4__7077_, data_stage_4__7076_, data_stage_4__7075_, data_stage_4__7074_, data_stage_4__7073_, data_stage_4__7072_, data_stage_4__7071_, data_stage_4__7070_, data_stage_4__7069_, data_stage_4__7068_, data_stage_4__7067_, data_stage_4__7066_, data_stage_4__7065_, data_stage_4__7064_, data_stage_4__7063_, data_stage_4__7062_, data_stage_4__7061_, data_stage_4__7060_, data_stage_4__7059_, data_stage_4__7058_, data_stage_4__7057_, data_stage_4__7056_, data_stage_4__7055_, data_stage_4__7054_, data_stage_4__7053_, data_stage_4__7052_, data_stage_4__7051_, data_stage_4__7050_, data_stage_4__7049_, data_stage_4__7048_, data_stage_4__7047_, data_stage_4__7046_, data_stage_4__7045_, data_stage_4__7044_, data_stage_4__7043_, data_stage_4__7042_, data_stage_4__7041_, data_stage_4__7040_, data_stage_4__7039_, data_stage_4__7038_, data_stage_4__7037_, data_stage_4__7036_, data_stage_4__7035_, data_stage_4__7034_, data_stage_4__7033_, data_stage_4__7032_, data_stage_4__7031_, data_stage_4__7030_, data_stage_4__7029_, data_stage_4__7028_, data_stage_4__7027_, data_stage_4__7026_, data_stage_4__7025_, data_stage_4__7024_, data_stage_4__7023_, data_stage_4__7022_, data_stage_4__7021_, data_stage_4__7020_, data_stage_4__7019_, data_stage_4__7018_, data_stage_4__7017_, data_stage_4__7016_, data_stage_4__7015_, data_stage_4__7014_, data_stage_4__7013_, data_stage_4__7012_, data_stage_4__7011_, data_stage_4__7010_, data_stage_4__7009_, data_stage_4__7008_, data_stage_4__7007_, data_stage_4__7006_, data_stage_4__7005_, data_stage_4__7004_, data_stage_4__7003_, data_stage_4__7002_, data_stage_4__7001_, data_stage_4__7000_, data_stage_4__6999_, data_stage_4__6998_, data_stage_4__6997_, data_stage_4__6996_, data_stage_4__6995_, data_stage_4__6994_, data_stage_4__6993_, data_stage_4__6992_, data_stage_4__6991_, data_stage_4__6990_, data_stage_4__6989_, data_stage_4__6988_, data_stage_4__6987_, data_stage_4__6986_, data_stage_4__6985_, data_stage_4__6984_, data_stage_4__6983_, data_stage_4__6982_, data_stage_4__6981_, data_stage_4__6980_, data_stage_4__6979_, data_stage_4__6978_, data_stage_4__6977_, data_stage_4__6976_, data_stage_4__6975_, data_stage_4__6974_, data_stage_4__6973_, data_stage_4__6972_, data_stage_4__6971_, data_stage_4__6970_, data_stage_4__6969_, data_stage_4__6968_, data_stage_4__6967_, data_stage_4__6966_, data_stage_4__6965_, data_stage_4__6964_, data_stage_4__6963_, data_stage_4__6962_, data_stage_4__6961_, data_stage_4__6960_, data_stage_4__6959_, data_stage_4__6958_, data_stage_4__6957_, data_stage_4__6956_, data_stage_4__6955_, data_stage_4__6954_, data_stage_4__6953_, data_stage_4__6952_, data_stage_4__6951_, data_stage_4__6950_, data_stage_4__6949_, data_stage_4__6948_, data_stage_4__6947_, data_stage_4__6946_, data_stage_4__6945_, data_stage_4__6944_, data_stage_4__6943_, data_stage_4__6942_, data_stage_4__6941_, data_stage_4__6940_, data_stage_4__6939_, data_stage_4__6938_, data_stage_4__6937_, data_stage_4__6936_, data_stage_4__6935_, data_stage_4__6934_, data_stage_4__6933_, data_stage_4__6932_, data_stage_4__6931_, data_stage_4__6930_, data_stage_4__6929_, data_stage_4__6928_, data_stage_4__6927_, data_stage_4__6926_, data_stage_4__6925_, data_stage_4__6924_, data_stage_4__6923_, data_stage_4__6922_, data_stage_4__6921_, data_stage_4__6920_, data_stage_4__6919_, data_stage_4__6918_, data_stage_4__6917_, data_stage_4__6916_, data_stage_4__6915_, data_stage_4__6914_, data_stage_4__6913_, data_stage_4__6912_, data_stage_4__6911_, data_stage_4__6910_, data_stage_4__6909_, data_stage_4__6908_, data_stage_4__6907_, data_stage_4__6906_, data_stage_4__6905_, data_stage_4__6904_, data_stage_4__6903_, data_stage_4__6902_, data_stage_4__6901_, data_stage_4__6900_, data_stage_4__6899_, data_stage_4__6898_, data_stage_4__6897_, data_stage_4__6896_, data_stage_4__6895_, data_stage_4__6894_, data_stage_4__6893_, data_stage_4__6892_, data_stage_4__6891_, data_stage_4__6890_, data_stage_4__6889_, data_stage_4__6888_, data_stage_4__6887_, data_stage_4__6886_, data_stage_4__6885_, data_stage_4__6884_, data_stage_4__6883_, data_stage_4__6882_, data_stage_4__6881_, data_stage_4__6880_, data_stage_4__6879_, data_stage_4__6878_, data_stage_4__6877_, data_stage_4__6876_, data_stage_4__6875_, data_stage_4__6874_, data_stage_4__6873_, data_stage_4__6872_, data_stage_4__6871_, data_stage_4__6870_, data_stage_4__6869_, data_stage_4__6868_, data_stage_4__6867_, data_stage_4__6866_, data_stage_4__6865_, data_stage_4__6864_, data_stage_4__6863_, data_stage_4__6862_, data_stage_4__6861_, data_stage_4__6860_, data_stage_4__6859_, data_stage_4__6858_, data_stage_4__6857_, data_stage_4__6856_, data_stage_4__6855_, data_stage_4__6854_, data_stage_4__6853_, data_stage_4__6852_, data_stage_4__6851_, data_stage_4__6850_, data_stage_4__6849_, data_stage_4__6848_, data_stage_4__6847_, data_stage_4__6846_, data_stage_4__6845_, data_stage_4__6844_, data_stage_4__6843_, data_stage_4__6842_, data_stage_4__6841_, data_stage_4__6840_, data_stage_4__6839_, data_stage_4__6838_, data_stage_4__6837_, data_stage_4__6836_, data_stage_4__6835_, data_stage_4__6834_, data_stage_4__6833_, data_stage_4__6832_, data_stage_4__6831_, data_stage_4__6830_, data_stage_4__6829_, data_stage_4__6828_, data_stage_4__6827_, data_stage_4__6826_, data_stage_4__6825_, data_stage_4__6824_, data_stage_4__6823_, data_stage_4__6822_, data_stage_4__6821_, data_stage_4__6820_, data_stage_4__6819_, data_stage_4__6818_, data_stage_4__6817_, data_stage_4__6816_, data_stage_4__6815_, data_stage_4__6814_, data_stage_4__6813_, data_stage_4__6812_, data_stage_4__6811_, data_stage_4__6810_, data_stage_4__6809_, data_stage_4__6808_, data_stage_4__6807_, data_stage_4__6806_, data_stage_4__6805_, data_stage_4__6804_, data_stage_4__6803_, data_stage_4__6802_, data_stage_4__6801_, data_stage_4__6800_, data_stage_4__6799_, data_stage_4__6798_, data_stage_4__6797_, data_stage_4__6796_, data_stage_4__6795_, data_stage_4__6794_, data_stage_4__6793_, data_stage_4__6792_, data_stage_4__6791_, data_stage_4__6790_, data_stage_4__6789_, data_stage_4__6788_, data_stage_4__6787_, data_stage_4__6786_, data_stage_4__6785_, data_stage_4__6784_, data_stage_4__6783_, data_stage_4__6782_, data_stage_4__6781_, data_stage_4__6780_, data_stage_4__6779_, data_stage_4__6778_, data_stage_4__6777_, data_stage_4__6776_, data_stage_4__6775_, data_stage_4__6774_, data_stage_4__6773_, data_stage_4__6772_, data_stage_4__6771_, data_stage_4__6770_, data_stage_4__6769_, data_stage_4__6768_, data_stage_4__6767_, data_stage_4__6766_, data_stage_4__6765_, data_stage_4__6764_, data_stage_4__6763_, data_stage_4__6762_, data_stage_4__6761_, data_stage_4__6760_, data_stage_4__6759_, data_stage_4__6758_, data_stage_4__6757_, data_stage_4__6756_, data_stage_4__6755_, data_stage_4__6754_, data_stage_4__6753_, data_stage_4__6752_, data_stage_4__6751_, data_stage_4__6750_, data_stage_4__6749_, data_stage_4__6748_, data_stage_4__6747_, data_stage_4__6746_, data_stage_4__6745_, data_stage_4__6744_, data_stage_4__6743_, data_stage_4__6742_, data_stage_4__6741_, data_stage_4__6740_, data_stage_4__6739_, data_stage_4__6738_, data_stage_4__6737_, data_stage_4__6736_, data_stage_4__6735_, data_stage_4__6734_, data_stage_4__6733_, data_stage_4__6732_, data_stage_4__6731_, data_stage_4__6730_, data_stage_4__6729_, data_stage_4__6728_, data_stage_4__6727_, data_stage_4__6726_, data_stage_4__6725_, data_stage_4__6724_, data_stage_4__6723_, data_stage_4__6722_, data_stage_4__6721_, data_stage_4__6720_, data_stage_4__6719_, data_stage_4__6718_, data_stage_4__6717_, data_stage_4__6716_, data_stage_4__6715_, data_stage_4__6714_, data_stage_4__6713_, data_stage_4__6712_, data_stage_4__6711_, data_stage_4__6710_, data_stage_4__6709_, data_stage_4__6708_, data_stage_4__6707_, data_stage_4__6706_, data_stage_4__6705_, data_stage_4__6704_, data_stage_4__6703_, data_stage_4__6702_, data_stage_4__6701_, data_stage_4__6700_, data_stage_4__6699_, data_stage_4__6698_, data_stage_4__6697_, data_stage_4__6696_, data_stage_4__6695_, data_stage_4__6694_, data_stage_4__6693_, data_stage_4__6692_, data_stage_4__6691_, data_stage_4__6690_, data_stage_4__6689_, data_stage_4__6688_, data_stage_4__6687_, data_stage_4__6686_, data_stage_4__6685_, data_stage_4__6684_, data_stage_4__6683_, data_stage_4__6682_, data_stage_4__6681_, data_stage_4__6680_, data_stage_4__6679_, data_stage_4__6678_, data_stage_4__6677_, data_stage_4__6676_, data_stage_4__6675_, data_stage_4__6674_, data_stage_4__6673_, data_stage_4__6672_, data_stage_4__6671_, data_stage_4__6670_, data_stage_4__6669_, data_stage_4__6668_, data_stage_4__6667_, data_stage_4__6666_, data_stage_4__6665_, data_stage_4__6664_, data_stage_4__6663_, data_stage_4__6662_, data_stage_4__6661_, data_stage_4__6660_, data_stage_4__6659_, data_stage_4__6658_, data_stage_4__6657_, data_stage_4__6656_, data_stage_4__6655_, data_stage_4__6654_, data_stage_4__6653_, data_stage_4__6652_, data_stage_4__6651_, data_stage_4__6650_, data_stage_4__6649_, data_stage_4__6648_, data_stage_4__6647_, data_stage_4__6646_, data_stage_4__6645_, data_stage_4__6644_, data_stage_4__6643_, data_stage_4__6642_, data_stage_4__6641_, data_stage_4__6640_, data_stage_4__6639_, data_stage_4__6638_, data_stage_4__6637_, data_stage_4__6636_, data_stage_4__6635_, data_stage_4__6634_, data_stage_4__6633_, data_stage_4__6632_, data_stage_4__6631_, data_stage_4__6630_, data_stage_4__6629_, data_stage_4__6628_, data_stage_4__6627_, data_stage_4__6626_, data_stage_4__6625_, data_stage_4__6624_, data_stage_4__6623_, data_stage_4__6622_, data_stage_4__6621_, data_stage_4__6620_, data_stage_4__6619_, data_stage_4__6618_, data_stage_4__6617_, data_stage_4__6616_, data_stage_4__6615_, data_stage_4__6614_, data_stage_4__6613_, data_stage_4__6612_, data_stage_4__6611_, data_stage_4__6610_, data_stage_4__6609_, data_stage_4__6608_, data_stage_4__6607_, data_stage_4__6606_, data_stage_4__6605_, data_stage_4__6604_, data_stage_4__6603_, data_stage_4__6602_, data_stage_4__6601_, data_stage_4__6600_, data_stage_4__6599_, data_stage_4__6598_, data_stage_4__6597_, data_stage_4__6596_, data_stage_4__6595_, data_stage_4__6594_, data_stage_4__6593_, data_stage_4__6592_, data_stage_4__6591_, data_stage_4__6590_, data_stage_4__6589_, data_stage_4__6588_, data_stage_4__6587_, data_stage_4__6586_, data_stage_4__6585_, data_stage_4__6584_, data_stage_4__6583_, data_stage_4__6582_, data_stage_4__6581_, data_stage_4__6580_, data_stage_4__6579_, data_stage_4__6578_, data_stage_4__6577_, data_stage_4__6576_, data_stage_4__6575_, data_stage_4__6574_, data_stage_4__6573_, data_stage_4__6572_, data_stage_4__6571_, data_stage_4__6570_, data_stage_4__6569_, data_stage_4__6568_, data_stage_4__6567_, data_stage_4__6566_, data_stage_4__6565_, data_stage_4__6564_, data_stage_4__6563_, data_stage_4__6562_, data_stage_4__6561_, data_stage_4__6560_, data_stage_4__6559_, data_stage_4__6558_, data_stage_4__6557_, data_stage_4__6556_, data_stage_4__6555_, data_stage_4__6554_, data_stage_4__6553_, data_stage_4__6552_, data_stage_4__6551_, data_stage_4__6550_, data_stage_4__6549_, data_stage_4__6548_, data_stage_4__6547_, data_stage_4__6546_, data_stage_4__6545_, data_stage_4__6544_, data_stage_4__6543_, data_stage_4__6542_, data_stage_4__6541_, data_stage_4__6540_, data_stage_4__6539_, data_stage_4__6538_, data_stage_4__6537_, data_stage_4__6536_, data_stage_4__6535_, data_stage_4__6534_, data_stage_4__6533_, data_stage_4__6532_, data_stage_4__6531_, data_stage_4__6530_, data_stage_4__6529_, data_stage_4__6528_, data_stage_4__6527_, data_stage_4__6526_, data_stage_4__6525_, data_stage_4__6524_, data_stage_4__6523_, data_stage_4__6522_, data_stage_4__6521_, data_stage_4__6520_, data_stage_4__6519_, data_stage_4__6518_, data_stage_4__6517_, data_stage_4__6516_, data_stage_4__6515_, data_stage_4__6514_, data_stage_4__6513_, data_stage_4__6512_, data_stage_4__6511_, data_stage_4__6510_, data_stage_4__6509_, data_stage_4__6508_, data_stage_4__6507_, data_stage_4__6506_, data_stage_4__6505_, data_stage_4__6504_, data_stage_4__6503_, data_stage_4__6502_, data_stage_4__6501_, data_stage_4__6500_, data_stage_4__6499_, data_stage_4__6498_, data_stage_4__6497_, data_stage_4__6496_, data_stage_4__6495_, data_stage_4__6494_, data_stage_4__6493_, data_stage_4__6492_, data_stage_4__6491_, data_stage_4__6490_, data_stage_4__6489_, data_stage_4__6488_, data_stage_4__6487_, data_stage_4__6486_, data_stage_4__6485_, data_stage_4__6484_, data_stage_4__6483_, data_stage_4__6482_, data_stage_4__6481_, data_stage_4__6480_, data_stage_4__6479_, data_stage_4__6478_, data_stage_4__6477_, data_stage_4__6476_, data_stage_4__6475_, data_stage_4__6474_, data_stage_4__6473_, data_stage_4__6472_, data_stage_4__6471_, data_stage_4__6470_, data_stage_4__6469_, data_stage_4__6468_, data_stage_4__6467_, data_stage_4__6466_, data_stage_4__6465_, data_stage_4__6464_, data_stage_4__6463_, data_stage_4__6462_, data_stage_4__6461_, data_stage_4__6460_, data_stage_4__6459_, data_stage_4__6458_, data_stage_4__6457_, data_stage_4__6456_, data_stage_4__6455_, data_stage_4__6454_, data_stage_4__6453_, data_stage_4__6452_, data_stage_4__6451_, data_stage_4__6450_, data_stage_4__6449_, data_stage_4__6448_, data_stage_4__6447_, data_stage_4__6446_, data_stage_4__6445_, data_stage_4__6444_, data_stage_4__6443_, data_stage_4__6442_, data_stage_4__6441_, data_stage_4__6440_, data_stage_4__6439_, data_stage_4__6438_, data_stage_4__6437_, data_stage_4__6436_, data_stage_4__6435_, data_stage_4__6434_, data_stage_4__6433_, data_stage_4__6432_, data_stage_4__6431_, data_stage_4__6430_, data_stage_4__6429_, data_stage_4__6428_, data_stage_4__6427_, data_stage_4__6426_, data_stage_4__6425_, data_stage_4__6424_, data_stage_4__6423_, data_stage_4__6422_, data_stage_4__6421_, data_stage_4__6420_, data_stage_4__6419_, data_stage_4__6418_, data_stage_4__6417_, data_stage_4__6416_, data_stage_4__6415_, data_stage_4__6414_, data_stage_4__6413_, data_stage_4__6412_, data_stage_4__6411_, data_stage_4__6410_, data_stage_4__6409_, data_stage_4__6408_, data_stage_4__6407_, data_stage_4__6406_, data_stage_4__6405_, data_stage_4__6404_, data_stage_4__6403_, data_stage_4__6402_, data_stage_4__6401_, data_stage_4__6400_, data_stage_4__6399_, data_stage_4__6398_, data_stage_4__6397_, data_stage_4__6396_, data_stage_4__6395_, data_stage_4__6394_, data_stage_4__6393_, data_stage_4__6392_, data_stage_4__6391_, data_stage_4__6390_, data_stage_4__6389_, data_stage_4__6388_, data_stage_4__6387_, data_stage_4__6386_, data_stage_4__6385_, data_stage_4__6384_, data_stage_4__6383_, data_stage_4__6382_, data_stage_4__6381_, data_stage_4__6380_, data_stage_4__6379_, data_stage_4__6378_, data_stage_4__6377_, data_stage_4__6376_, data_stage_4__6375_, data_stage_4__6374_, data_stage_4__6373_, data_stage_4__6372_, data_stage_4__6371_, data_stage_4__6370_, data_stage_4__6369_, data_stage_4__6368_, data_stage_4__6367_, data_stage_4__6366_, data_stage_4__6365_, data_stage_4__6364_, data_stage_4__6363_, data_stage_4__6362_, data_stage_4__6361_, data_stage_4__6360_, data_stage_4__6359_, data_stage_4__6358_, data_stage_4__6357_, data_stage_4__6356_, data_stage_4__6355_, data_stage_4__6354_, data_stage_4__6353_, data_stage_4__6352_, data_stage_4__6351_, data_stage_4__6350_, data_stage_4__6349_, data_stage_4__6348_, data_stage_4__6347_, data_stage_4__6346_, data_stage_4__6345_, data_stage_4__6344_, data_stage_4__6343_, data_stage_4__6342_, data_stage_4__6341_, data_stage_4__6340_, data_stage_4__6339_, data_stage_4__6338_, data_stage_4__6337_, data_stage_4__6336_, data_stage_4__6335_, data_stage_4__6334_, data_stage_4__6333_, data_stage_4__6332_, data_stage_4__6331_, data_stage_4__6330_, data_stage_4__6329_, data_stage_4__6328_, data_stage_4__6327_, data_stage_4__6326_, data_stage_4__6325_, data_stage_4__6324_, data_stage_4__6323_, data_stage_4__6322_, data_stage_4__6321_, data_stage_4__6320_, data_stage_4__6319_, data_stage_4__6318_, data_stage_4__6317_, data_stage_4__6316_, data_stage_4__6315_, data_stage_4__6314_, data_stage_4__6313_, data_stage_4__6312_, data_stage_4__6311_, data_stage_4__6310_, data_stage_4__6309_, data_stage_4__6308_, data_stage_4__6307_, data_stage_4__6306_, data_stage_4__6305_, data_stage_4__6304_, data_stage_4__6303_, data_stage_4__6302_, data_stage_4__6301_, data_stage_4__6300_, data_stage_4__6299_, data_stage_4__6298_, data_stage_4__6297_, data_stage_4__6296_, data_stage_4__6295_, data_stage_4__6294_, data_stage_4__6293_, data_stage_4__6292_, data_stage_4__6291_, data_stage_4__6290_, data_stage_4__6289_, data_stage_4__6288_, data_stage_4__6287_, data_stage_4__6286_, data_stage_4__6285_, data_stage_4__6284_, data_stage_4__6283_, data_stage_4__6282_, data_stage_4__6281_, data_stage_4__6280_, data_stage_4__6279_, data_stage_4__6278_, data_stage_4__6277_, data_stage_4__6276_, data_stage_4__6275_, data_stage_4__6274_, data_stage_4__6273_, data_stage_4__6272_, data_stage_4__6271_, data_stage_4__6270_, data_stage_4__6269_, data_stage_4__6268_, data_stage_4__6267_, data_stage_4__6266_, data_stage_4__6265_, data_stage_4__6264_, data_stage_4__6263_, data_stage_4__6262_, data_stage_4__6261_, data_stage_4__6260_, data_stage_4__6259_, data_stage_4__6258_, data_stage_4__6257_, data_stage_4__6256_, data_stage_4__6255_, data_stage_4__6254_, data_stage_4__6253_, data_stage_4__6252_, data_stage_4__6251_, data_stage_4__6250_, data_stage_4__6249_, data_stage_4__6248_, data_stage_4__6247_, data_stage_4__6246_, data_stage_4__6245_, data_stage_4__6244_, data_stage_4__6243_, data_stage_4__6242_, data_stage_4__6241_, data_stage_4__6240_, data_stage_4__6239_, data_stage_4__6238_, data_stage_4__6237_, data_stage_4__6236_, data_stage_4__6235_, data_stage_4__6234_, data_stage_4__6233_, data_stage_4__6232_, data_stage_4__6231_, data_stage_4__6230_, data_stage_4__6229_, data_stage_4__6228_, data_stage_4__6227_, data_stage_4__6226_, data_stage_4__6225_, data_stage_4__6224_, data_stage_4__6223_, data_stage_4__6222_, data_stage_4__6221_, data_stage_4__6220_, data_stage_4__6219_, data_stage_4__6218_, data_stage_4__6217_, data_stage_4__6216_, data_stage_4__6215_, data_stage_4__6214_, data_stage_4__6213_, data_stage_4__6212_, data_stage_4__6211_, data_stage_4__6210_, data_stage_4__6209_, data_stage_4__6208_, data_stage_4__6207_, data_stage_4__6206_, data_stage_4__6205_, data_stage_4__6204_, data_stage_4__6203_, data_stage_4__6202_, data_stage_4__6201_, data_stage_4__6200_, data_stage_4__6199_, data_stage_4__6198_, data_stage_4__6197_, data_stage_4__6196_, data_stage_4__6195_, data_stage_4__6194_, data_stage_4__6193_, data_stage_4__6192_, data_stage_4__6191_, data_stage_4__6190_, data_stage_4__6189_, data_stage_4__6188_, data_stage_4__6187_, data_stage_4__6186_, data_stage_4__6185_, data_stage_4__6184_, data_stage_4__6183_, data_stage_4__6182_, data_stage_4__6181_, data_stage_4__6180_, data_stage_4__6179_, data_stage_4__6178_, data_stage_4__6177_, data_stage_4__6176_, data_stage_4__6175_, data_stage_4__6174_, data_stage_4__6173_, data_stage_4__6172_, data_stage_4__6171_, data_stage_4__6170_, data_stage_4__6169_, data_stage_4__6168_, data_stage_4__6167_, data_stage_4__6166_, data_stage_4__6165_, data_stage_4__6164_, data_stage_4__6163_, data_stage_4__6162_, data_stage_4__6161_, data_stage_4__6160_, data_stage_4__6159_, data_stage_4__6158_, data_stage_4__6157_, data_stage_4__6156_, data_stage_4__6155_, data_stage_4__6154_, data_stage_4__6153_, data_stage_4__6152_, data_stage_4__6151_, data_stage_4__6150_, data_stage_4__6149_, data_stage_4__6148_, data_stage_4__6147_, data_stage_4__6146_, data_stage_4__6145_, data_stage_4__6144_, data_stage_4__6143_, data_stage_4__6142_, data_stage_4__6141_, data_stage_4__6140_, data_stage_4__6139_, data_stage_4__6138_, data_stage_4__6137_, data_stage_4__6136_, data_stage_4__6135_, data_stage_4__6134_, data_stage_4__6133_, data_stage_4__6132_, data_stage_4__6131_, data_stage_4__6130_, data_stage_4__6129_, data_stage_4__6128_, data_stage_4__6127_, data_stage_4__6126_, data_stage_4__6125_, data_stage_4__6124_, data_stage_4__6123_, data_stage_4__6122_, data_stage_4__6121_, data_stage_4__6120_, data_stage_4__6119_, data_stage_4__6118_, data_stage_4__6117_, data_stage_4__6116_, data_stage_4__6115_, data_stage_4__6114_, data_stage_4__6113_, data_stage_4__6112_, data_stage_4__6111_, data_stage_4__6110_, data_stage_4__6109_, data_stage_4__6108_, data_stage_4__6107_, data_stage_4__6106_, data_stage_4__6105_, data_stage_4__6104_, data_stage_4__6103_, data_stage_4__6102_, data_stage_4__6101_, data_stage_4__6100_, data_stage_4__6099_, data_stage_4__6098_, data_stage_4__6097_, data_stage_4__6096_, data_stage_4__6095_, data_stage_4__6094_, data_stage_4__6093_, data_stage_4__6092_, data_stage_4__6091_, data_stage_4__6090_, data_stage_4__6089_, data_stage_4__6088_, data_stage_4__6087_, data_stage_4__6086_, data_stage_4__6085_, data_stage_4__6084_, data_stage_4__6083_, data_stage_4__6082_, data_stage_4__6081_, data_stage_4__6080_, data_stage_4__6079_, data_stage_4__6078_, data_stage_4__6077_, data_stage_4__6076_, data_stage_4__6075_, data_stage_4__6074_, data_stage_4__6073_, data_stage_4__6072_, data_stage_4__6071_, data_stage_4__6070_, data_stage_4__6069_, data_stage_4__6068_, data_stage_4__6067_, data_stage_4__6066_, data_stage_4__6065_, data_stage_4__6064_, data_stage_4__6063_, data_stage_4__6062_, data_stage_4__6061_, data_stage_4__6060_, data_stage_4__6059_, data_stage_4__6058_, data_stage_4__6057_, data_stage_4__6056_, data_stage_4__6055_, data_stage_4__6054_, data_stage_4__6053_, data_stage_4__6052_, data_stage_4__6051_, data_stage_4__6050_, data_stage_4__6049_, data_stage_4__6048_, data_stage_4__6047_, data_stage_4__6046_, data_stage_4__6045_, data_stage_4__6044_, data_stage_4__6043_, data_stage_4__6042_, data_stage_4__6041_, data_stage_4__6040_, data_stage_4__6039_, data_stage_4__6038_, data_stage_4__6037_, data_stage_4__6036_, data_stage_4__6035_, data_stage_4__6034_, data_stage_4__6033_, data_stage_4__6032_, data_stage_4__6031_, data_stage_4__6030_, data_stage_4__6029_, data_stage_4__6028_, data_stage_4__6027_, data_stage_4__6026_, data_stage_4__6025_, data_stage_4__6024_, data_stage_4__6023_, data_stage_4__6022_, data_stage_4__6021_, data_stage_4__6020_, data_stage_4__6019_, data_stage_4__6018_, data_stage_4__6017_, data_stage_4__6016_, data_stage_4__6015_, data_stage_4__6014_, data_stage_4__6013_, data_stage_4__6012_, data_stage_4__6011_, data_stage_4__6010_, data_stage_4__6009_, data_stage_4__6008_, data_stage_4__6007_, data_stage_4__6006_, data_stage_4__6005_, data_stage_4__6004_, data_stage_4__6003_, data_stage_4__6002_, data_stage_4__6001_, data_stage_4__6000_, data_stage_4__5999_, data_stage_4__5998_, data_stage_4__5997_, data_stage_4__5996_, data_stage_4__5995_, data_stage_4__5994_, data_stage_4__5993_, data_stage_4__5992_, data_stage_4__5991_, data_stage_4__5990_, data_stage_4__5989_, data_stage_4__5988_, data_stage_4__5987_, data_stage_4__5986_, data_stage_4__5985_, data_stage_4__5984_, data_stage_4__5983_, data_stage_4__5982_, data_stage_4__5981_, data_stage_4__5980_, data_stage_4__5979_, data_stage_4__5978_, data_stage_4__5977_, data_stage_4__5976_, data_stage_4__5975_, data_stage_4__5974_, data_stage_4__5973_, data_stage_4__5972_, data_stage_4__5971_, data_stage_4__5970_, data_stage_4__5969_, data_stage_4__5968_, data_stage_4__5967_, data_stage_4__5966_, data_stage_4__5965_, data_stage_4__5964_, data_stage_4__5963_, data_stage_4__5962_, data_stage_4__5961_, data_stage_4__5960_, data_stage_4__5959_, data_stage_4__5958_, data_stage_4__5957_, data_stage_4__5956_, data_stage_4__5955_, data_stage_4__5954_, data_stage_4__5953_, data_stage_4__5952_, data_stage_4__5951_, data_stage_4__5950_, data_stage_4__5949_, data_stage_4__5948_, data_stage_4__5947_, data_stage_4__5946_, data_stage_4__5945_, data_stage_4__5944_, data_stage_4__5943_, data_stage_4__5942_, data_stage_4__5941_, data_stage_4__5940_, data_stage_4__5939_, data_stage_4__5938_, data_stage_4__5937_, data_stage_4__5936_, data_stage_4__5935_, data_stage_4__5934_, data_stage_4__5933_, data_stage_4__5932_, data_stage_4__5931_, data_stage_4__5930_, data_stage_4__5929_, data_stage_4__5928_, data_stage_4__5927_, data_stage_4__5926_, data_stage_4__5925_, data_stage_4__5924_, data_stage_4__5923_, data_stage_4__5922_, data_stage_4__5921_, data_stage_4__5920_, data_stage_4__5919_, data_stage_4__5918_, data_stage_4__5917_, data_stage_4__5916_, data_stage_4__5915_, data_stage_4__5914_, data_stage_4__5913_, data_stage_4__5912_, data_stage_4__5911_, data_stage_4__5910_, data_stage_4__5909_, data_stage_4__5908_, data_stage_4__5907_, data_stage_4__5906_, data_stage_4__5905_, data_stage_4__5904_, data_stage_4__5903_, data_stage_4__5902_, data_stage_4__5901_, data_stage_4__5900_, data_stage_4__5899_, data_stage_4__5898_, data_stage_4__5897_, data_stage_4__5896_, data_stage_4__5895_, data_stage_4__5894_, data_stage_4__5893_, data_stage_4__5892_, data_stage_4__5891_, data_stage_4__5890_, data_stage_4__5889_, data_stage_4__5888_, data_stage_4__5887_, data_stage_4__5886_, data_stage_4__5885_, data_stage_4__5884_, data_stage_4__5883_, data_stage_4__5882_, data_stage_4__5881_, data_stage_4__5880_, data_stage_4__5879_, data_stage_4__5878_, data_stage_4__5877_, data_stage_4__5876_, data_stage_4__5875_, data_stage_4__5874_, data_stage_4__5873_, data_stage_4__5872_, data_stage_4__5871_, data_stage_4__5870_, data_stage_4__5869_, data_stage_4__5868_, data_stage_4__5867_, data_stage_4__5866_, data_stage_4__5865_, data_stage_4__5864_, data_stage_4__5863_, data_stage_4__5862_, data_stage_4__5861_, data_stage_4__5860_, data_stage_4__5859_, data_stage_4__5858_, data_stage_4__5857_, data_stage_4__5856_, data_stage_4__5855_, data_stage_4__5854_, data_stage_4__5853_, data_stage_4__5852_, data_stage_4__5851_, data_stage_4__5850_, data_stage_4__5849_, data_stage_4__5848_, data_stage_4__5847_, data_stage_4__5846_, data_stage_4__5845_, data_stage_4__5844_, data_stage_4__5843_, data_stage_4__5842_, data_stage_4__5841_, data_stage_4__5840_, data_stage_4__5839_, data_stage_4__5838_, data_stage_4__5837_, data_stage_4__5836_, data_stage_4__5835_, data_stage_4__5834_, data_stage_4__5833_, data_stage_4__5832_, data_stage_4__5831_, data_stage_4__5830_, data_stage_4__5829_, data_stage_4__5828_, data_stage_4__5827_, data_stage_4__5826_, data_stage_4__5825_, data_stage_4__5824_, data_stage_4__5823_, data_stage_4__5822_, data_stage_4__5821_, data_stage_4__5820_, data_stage_4__5819_, data_stage_4__5818_, data_stage_4__5817_, data_stage_4__5816_, data_stage_4__5815_, data_stage_4__5814_, data_stage_4__5813_, data_stage_4__5812_, data_stage_4__5811_, data_stage_4__5810_, data_stage_4__5809_, data_stage_4__5808_, data_stage_4__5807_, data_stage_4__5806_, data_stage_4__5805_, data_stage_4__5804_, data_stage_4__5803_, data_stage_4__5802_, data_stage_4__5801_, data_stage_4__5800_, data_stage_4__5799_, data_stage_4__5798_, data_stage_4__5797_, data_stage_4__5796_, data_stage_4__5795_, data_stage_4__5794_, data_stage_4__5793_, data_stage_4__5792_, data_stage_4__5791_, data_stage_4__5790_, data_stage_4__5789_, data_stage_4__5788_, data_stage_4__5787_, data_stage_4__5786_, data_stage_4__5785_, data_stage_4__5784_, data_stage_4__5783_, data_stage_4__5782_, data_stage_4__5781_, data_stage_4__5780_, data_stage_4__5779_, data_stage_4__5778_, data_stage_4__5777_, data_stage_4__5776_, data_stage_4__5775_, data_stage_4__5774_, data_stage_4__5773_, data_stage_4__5772_, data_stage_4__5771_, data_stage_4__5770_, data_stage_4__5769_, data_stage_4__5768_, data_stage_4__5767_, data_stage_4__5766_, data_stage_4__5765_, data_stage_4__5764_, data_stage_4__5763_, data_stage_4__5762_, data_stage_4__5761_, data_stage_4__5760_, data_stage_4__5759_, data_stage_4__5758_, data_stage_4__5757_, data_stage_4__5756_, data_stage_4__5755_, data_stage_4__5754_, data_stage_4__5753_, data_stage_4__5752_, data_stage_4__5751_, data_stage_4__5750_, data_stage_4__5749_, data_stage_4__5748_, data_stage_4__5747_, data_stage_4__5746_, data_stage_4__5745_, data_stage_4__5744_, data_stage_4__5743_, data_stage_4__5742_, data_stage_4__5741_, data_stage_4__5740_, data_stage_4__5739_, data_stage_4__5738_, data_stage_4__5737_, data_stage_4__5736_, data_stage_4__5735_, data_stage_4__5734_, data_stage_4__5733_, data_stage_4__5732_, data_stage_4__5731_, data_stage_4__5730_, data_stage_4__5729_, data_stage_4__5728_, data_stage_4__5727_, data_stage_4__5726_, data_stage_4__5725_, data_stage_4__5724_, data_stage_4__5723_, data_stage_4__5722_, data_stage_4__5721_, data_stage_4__5720_, data_stage_4__5719_, data_stage_4__5718_, data_stage_4__5717_, data_stage_4__5716_, data_stage_4__5715_, data_stage_4__5714_, data_stage_4__5713_, data_stage_4__5712_, data_stage_4__5711_, data_stage_4__5710_, data_stage_4__5709_, data_stage_4__5708_, data_stage_4__5707_, data_stage_4__5706_, data_stage_4__5705_, data_stage_4__5704_, data_stage_4__5703_, data_stage_4__5702_, data_stage_4__5701_, data_stage_4__5700_, data_stage_4__5699_, data_stage_4__5698_, data_stage_4__5697_, data_stage_4__5696_, data_stage_4__5695_, data_stage_4__5694_, data_stage_4__5693_, data_stage_4__5692_, data_stage_4__5691_, data_stage_4__5690_, data_stage_4__5689_, data_stage_4__5688_, data_stage_4__5687_, data_stage_4__5686_, data_stage_4__5685_, data_stage_4__5684_, data_stage_4__5683_, data_stage_4__5682_, data_stage_4__5681_, data_stage_4__5680_, data_stage_4__5679_, data_stage_4__5678_, data_stage_4__5677_, data_stage_4__5676_, data_stage_4__5675_, data_stage_4__5674_, data_stage_4__5673_, data_stage_4__5672_, data_stage_4__5671_, data_stage_4__5670_, data_stage_4__5669_, data_stage_4__5668_, data_stage_4__5667_, data_stage_4__5666_, data_stage_4__5665_, data_stage_4__5664_, data_stage_4__5663_, data_stage_4__5662_, data_stage_4__5661_, data_stage_4__5660_, data_stage_4__5659_, data_stage_4__5658_, data_stage_4__5657_, data_stage_4__5656_, data_stage_4__5655_, data_stage_4__5654_, data_stage_4__5653_, data_stage_4__5652_, data_stage_4__5651_, data_stage_4__5650_, data_stage_4__5649_, data_stage_4__5648_, data_stage_4__5647_, data_stage_4__5646_, data_stage_4__5645_, data_stage_4__5644_, data_stage_4__5643_, data_stage_4__5642_, data_stage_4__5641_, data_stage_4__5640_, data_stage_4__5639_, data_stage_4__5638_, data_stage_4__5637_, data_stage_4__5636_, data_stage_4__5635_, data_stage_4__5634_, data_stage_4__5633_, data_stage_4__5632_, data_stage_4__5631_, data_stage_4__5630_, data_stage_4__5629_, data_stage_4__5628_, data_stage_4__5627_, data_stage_4__5626_, data_stage_4__5625_, data_stage_4__5624_, data_stage_4__5623_, data_stage_4__5622_, data_stage_4__5621_, data_stage_4__5620_, data_stage_4__5619_, data_stage_4__5618_, data_stage_4__5617_, data_stage_4__5616_, data_stage_4__5615_, data_stage_4__5614_, data_stage_4__5613_, data_stage_4__5612_, data_stage_4__5611_, data_stage_4__5610_, data_stage_4__5609_, data_stage_4__5608_, data_stage_4__5607_, data_stage_4__5606_, data_stage_4__5605_, data_stage_4__5604_, data_stage_4__5603_, data_stage_4__5602_, data_stage_4__5601_, data_stage_4__5600_, data_stage_4__5599_, data_stage_4__5598_, data_stage_4__5597_, data_stage_4__5596_, data_stage_4__5595_, data_stage_4__5594_, data_stage_4__5593_, data_stage_4__5592_, data_stage_4__5591_, data_stage_4__5590_, data_stage_4__5589_, data_stage_4__5588_, data_stage_4__5587_, data_stage_4__5586_, data_stage_4__5585_, data_stage_4__5584_, data_stage_4__5583_, data_stage_4__5582_, data_stage_4__5581_, data_stage_4__5580_, data_stage_4__5579_, data_stage_4__5578_, data_stage_4__5577_, data_stage_4__5576_, data_stage_4__5575_, data_stage_4__5574_, data_stage_4__5573_, data_stage_4__5572_, data_stage_4__5571_, data_stage_4__5570_, data_stage_4__5569_, data_stage_4__5568_, data_stage_4__5567_, data_stage_4__5566_, data_stage_4__5565_, data_stage_4__5564_, data_stage_4__5563_, data_stage_4__5562_, data_stage_4__5561_, data_stage_4__5560_, data_stage_4__5559_, data_stage_4__5558_, data_stage_4__5557_, data_stage_4__5556_, data_stage_4__5555_, data_stage_4__5554_, data_stage_4__5553_, data_stage_4__5552_, data_stage_4__5551_, data_stage_4__5550_, data_stage_4__5549_, data_stage_4__5548_, data_stage_4__5547_, data_stage_4__5546_, data_stage_4__5545_, data_stage_4__5544_, data_stage_4__5543_, data_stage_4__5542_, data_stage_4__5541_, data_stage_4__5540_, data_stage_4__5539_, data_stage_4__5538_, data_stage_4__5537_, data_stage_4__5536_, data_stage_4__5535_, data_stage_4__5534_, data_stage_4__5533_, data_stage_4__5532_, data_stage_4__5531_, data_stage_4__5530_, data_stage_4__5529_, data_stage_4__5528_, data_stage_4__5527_, data_stage_4__5526_, data_stage_4__5525_, data_stage_4__5524_, data_stage_4__5523_, data_stage_4__5522_, data_stage_4__5521_, data_stage_4__5520_, data_stage_4__5519_, data_stage_4__5518_, data_stage_4__5517_, data_stage_4__5516_, data_stage_4__5515_, data_stage_4__5514_, data_stage_4__5513_, data_stage_4__5512_, data_stage_4__5511_, data_stage_4__5510_, data_stage_4__5509_, data_stage_4__5508_, data_stage_4__5507_, data_stage_4__5506_, data_stage_4__5505_, data_stage_4__5504_, data_stage_4__5503_, data_stage_4__5502_, data_stage_4__5501_, data_stage_4__5500_, data_stage_4__5499_, data_stage_4__5498_, data_stage_4__5497_, data_stage_4__5496_, data_stage_4__5495_, data_stage_4__5494_, data_stage_4__5493_, data_stage_4__5492_, data_stage_4__5491_, data_stage_4__5490_, data_stage_4__5489_, data_stage_4__5488_, data_stage_4__5487_, data_stage_4__5486_, data_stage_4__5485_, data_stage_4__5484_, data_stage_4__5483_, data_stage_4__5482_, data_stage_4__5481_, data_stage_4__5480_, data_stage_4__5479_, data_stage_4__5478_, data_stage_4__5477_, data_stage_4__5476_, data_stage_4__5475_, data_stage_4__5474_, data_stage_4__5473_, data_stage_4__5472_, data_stage_4__5471_, data_stage_4__5470_, data_stage_4__5469_, data_stage_4__5468_, data_stage_4__5467_, data_stage_4__5466_, data_stage_4__5465_, data_stage_4__5464_, data_stage_4__5463_, data_stage_4__5462_, data_stage_4__5461_, data_stage_4__5460_, data_stage_4__5459_, data_stage_4__5458_, data_stage_4__5457_, data_stage_4__5456_, data_stage_4__5455_, data_stage_4__5454_, data_stage_4__5453_, data_stage_4__5452_, data_stage_4__5451_, data_stage_4__5450_, data_stage_4__5449_, data_stage_4__5448_, data_stage_4__5447_, data_stage_4__5446_, data_stage_4__5445_, data_stage_4__5444_, data_stage_4__5443_, data_stage_4__5442_, data_stage_4__5441_, data_stage_4__5440_, data_stage_4__5439_, data_stage_4__5438_, data_stage_4__5437_, data_stage_4__5436_, data_stage_4__5435_, data_stage_4__5434_, data_stage_4__5433_, data_stage_4__5432_, data_stage_4__5431_, data_stage_4__5430_, data_stage_4__5429_, data_stage_4__5428_, data_stage_4__5427_, data_stage_4__5426_, data_stage_4__5425_, data_stage_4__5424_, data_stage_4__5423_, data_stage_4__5422_, data_stage_4__5421_, data_stage_4__5420_, data_stage_4__5419_, data_stage_4__5418_, data_stage_4__5417_, data_stage_4__5416_, data_stage_4__5415_, data_stage_4__5414_, data_stage_4__5413_, data_stage_4__5412_, data_stage_4__5411_, data_stage_4__5410_, data_stage_4__5409_, data_stage_4__5408_, data_stage_4__5407_, data_stage_4__5406_, data_stage_4__5405_, data_stage_4__5404_, data_stage_4__5403_, data_stage_4__5402_, data_stage_4__5401_, data_stage_4__5400_, data_stage_4__5399_, data_stage_4__5398_, data_stage_4__5397_, data_stage_4__5396_, data_stage_4__5395_, data_stage_4__5394_, data_stage_4__5393_, data_stage_4__5392_, data_stage_4__5391_, data_stage_4__5390_, data_stage_4__5389_, data_stage_4__5388_, data_stage_4__5387_, data_stage_4__5386_, data_stage_4__5385_, data_stage_4__5384_, data_stage_4__5383_, data_stage_4__5382_, data_stage_4__5381_, data_stage_4__5380_, data_stage_4__5379_, data_stage_4__5378_, data_stage_4__5377_, data_stage_4__5376_, data_stage_4__5375_, data_stage_4__5374_, data_stage_4__5373_, data_stage_4__5372_, data_stage_4__5371_, data_stage_4__5370_, data_stage_4__5369_, data_stage_4__5368_, data_stage_4__5367_, data_stage_4__5366_, data_stage_4__5365_, data_stage_4__5364_, data_stage_4__5363_, data_stage_4__5362_, data_stage_4__5361_, data_stage_4__5360_, data_stage_4__5359_, data_stage_4__5358_, data_stage_4__5357_, data_stage_4__5356_, data_stage_4__5355_, data_stage_4__5354_, data_stage_4__5353_, data_stage_4__5352_, data_stage_4__5351_, data_stage_4__5350_, data_stage_4__5349_, data_stage_4__5348_, data_stage_4__5347_, data_stage_4__5346_, data_stage_4__5345_, data_stage_4__5344_, data_stage_4__5343_, data_stage_4__5342_, data_stage_4__5341_, data_stage_4__5340_, data_stage_4__5339_, data_stage_4__5338_, data_stage_4__5337_, data_stage_4__5336_, data_stage_4__5335_, data_stage_4__5334_, data_stage_4__5333_, data_stage_4__5332_, data_stage_4__5331_, data_stage_4__5330_, data_stage_4__5329_, data_stage_4__5328_, data_stage_4__5327_, data_stage_4__5326_, data_stage_4__5325_, data_stage_4__5324_, data_stage_4__5323_, data_stage_4__5322_, data_stage_4__5321_, data_stage_4__5320_, data_stage_4__5319_, data_stage_4__5318_, data_stage_4__5317_, data_stage_4__5316_, data_stage_4__5315_, data_stage_4__5314_, data_stage_4__5313_, data_stage_4__5312_, data_stage_4__5311_, data_stage_4__5310_, data_stage_4__5309_, data_stage_4__5308_, data_stage_4__5307_, data_stage_4__5306_, data_stage_4__5305_, data_stage_4__5304_, data_stage_4__5303_, data_stage_4__5302_, data_stage_4__5301_, data_stage_4__5300_, data_stage_4__5299_, data_stage_4__5298_, data_stage_4__5297_, data_stage_4__5296_, data_stage_4__5295_, data_stage_4__5294_, data_stage_4__5293_, data_stage_4__5292_, data_stage_4__5291_, data_stage_4__5290_, data_stage_4__5289_, data_stage_4__5288_, data_stage_4__5287_, data_stage_4__5286_, data_stage_4__5285_, data_stage_4__5284_, data_stage_4__5283_, data_stage_4__5282_, data_stage_4__5281_, data_stage_4__5280_, data_stage_4__5279_, data_stage_4__5278_, data_stage_4__5277_, data_stage_4__5276_, data_stage_4__5275_, data_stage_4__5274_, data_stage_4__5273_, data_stage_4__5272_, data_stage_4__5271_, data_stage_4__5270_, data_stage_4__5269_, data_stage_4__5268_, data_stage_4__5267_, data_stage_4__5266_, data_stage_4__5265_, data_stage_4__5264_, data_stage_4__5263_, data_stage_4__5262_, data_stage_4__5261_, data_stage_4__5260_, data_stage_4__5259_, data_stage_4__5258_, data_stage_4__5257_, data_stage_4__5256_, data_stage_4__5255_, data_stage_4__5254_, data_stage_4__5253_, data_stage_4__5252_, data_stage_4__5251_, data_stage_4__5250_, data_stage_4__5249_, data_stage_4__5248_, data_stage_4__5247_, data_stage_4__5246_, data_stage_4__5245_, data_stage_4__5244_, data_stage_4__5243_, data_stage_4__5242_, data_stage_4__5241_, data_stage_4__5240_, data_stage_4__5239_, data_stage_4__5238_, data_stage_4__5237_, data_stage_4__5236_, data_stage_4__5235_, data_stage_4__5234_, data_stage_4__5233_, data_stage_4__5232_, data_stage_4__5231_, data_stage_4__5230_, data_stage_4__5229_, data_stage_4__5228_, data_stage_4__5227_, data_stage_4__5226_, data_stage_4__5225_, data_stage_4__5224_, data_stage_4__5223_, data_stage_4__5222_, data_stage_4__5221_, data_stage_4__5220_, data_stage_4__5219_, data_stage_4__5218_, data_stage_4__5217_, data_stage_4__5216_, data_stage_4__5215_, data_stage_4__5214_, data_stage_4__5213_, data_stage_4__5212_, data_stage_4__5211_, data_stage_4__5210_, data_stage_4__5209_, data_stage_4__5208_, data_stage_4__5207_, data_stage_4__5206_, data_stage_4__5205_, data_stage_4__5204_, data_stage_4__5203_, data_stage_4__5202_, data_stage_4__5201_, data_stage_4__5200_, data_stage_4__5199_, data_stage_4__5198_, data_stage_4__5197_, data_stage_4__5196_, data_stage_4__5195_, data_stage_4__5194_, data_stage_4__5193_, data_stage_4__5192_, data_stage_4__5191_, data_stage_4__5190_, data_stage_4__5189_, data_stage_4__5188_, data_stage_4__5187_, data_stage_4__5186_, data_stage_4__5185_, data_stage_4__5184_, data_stage_4__5183_, data_stage_4__5182_, data_stage_4__5181_, data_stage_4__5180_, data_stage_4__5179_, data_stage_4__5178_, data_stage_4__5177_, data_stage_4__5176_, data_stage_4__5175_, data_stage_4__5174_, data_stage_4__5173_, data_stage_4__5172_, data_stage_4__5171_, data_stage_4__5170_, data_stage_4__5169_, data_stage_4__5168_, data_stage_4__5167_, data_stage_4__5166_, data_stage_4__5165_, data_stage_4__5164_, data_stage_4__5163_, data_stage_4__5162_, data_stage_4__5161_, data_stage_4__5160_, data_stage_4__5159_, data_stage_4__5158_, data_stage_4__5157_, data_stage_4__5156_, data_stage_4__5155_, data_stage_4__5154_, data_stage_4__5153_, data_stage_4__5152_, data_stage_4__5151_, data_stage_4__5150_, data_stage_4__5149_, data_stage_4__5148_, data_stage_4__5147_, data_stage_4__5146_, data_stage_4__5145_, data_stage_4__5144_, data_stage_4__5143_, data_stage_4__5142_, data_stage_4__5141_, data_stage_4__5140_, data_stage_4__5139_, data_stage_4__5138_, data_stage_4__5137_, data_stage_4__5136_, data_stage_4__5135_, data_stage_4__5134_, data_stage_4__5133_, data_stage_4__5132_, data_stage_4__5131_, data_stage_4__5130_, data_stage_4__5129_, data_stage_4__5128_, data_stage_4__5127_, data_stage_4__5126_, data_stage_4__5125_, data_stage_4__5124_, data_stage_4__5123_, data_stage_4__5122_, data_stage_4__5121_, data_stage_4__5120_, data_stage_4__5119_, data_stage_4__5118_, data_stage_4__5117_, data_stage_4__5116_, data_stage_4__5115_, data_stage_4__5114_, data_stage_4__5113_, data_stage_4__5112_, data_stage_4__5111_, data_stage_4__5110_, data_stage_4__5109_, data_stage_4__5108_, data_stage_4__5107_, data_stage_4__5106_, data_stage_4__5105_, data_stage_4__5104_, data_stage_4__5103_, data_stage_4__5102_, data_stage_4__5101_, data_stage_4__5100_, data_stage_4__5099_, data_stage_4__5098_, data_stage_4__5097_, data_stage_4__5096_, data_stage_4__5095_, data_stage_4__5094_, data_stage_4__5093_, data_stage_4__5092_, data_stage_4__5091_, data_stage_4__5090_, data_stage_4__5089_, data_stage_4__5088_, data_stage_4__5087_, data_stage_4__5086_, data_stage_4__5085_, data_stage_4__5084_, data_stage_4__5083_, data_stage_4__5082_, data_stage_4__5081_, data_stage_4__5080_, data_stage_4__5079_, data_stage_4__5078_, data_stage_4__5077_, data_stage_4__5076_, data_stage_4__5075_, data_stage_4__5074_, data_stage_4__5073_, data_stage_4__5072_, data_stage_4__5071_, data_stage_4__5070_, data_stage_4__5069_, data_stage_4__5068_, data_stage_4__5067_, data_stage_4__5066_, data_stage_4__5065_, data_stage_4__5064_, data_stage_4__5063_, data_stage_4__5062_, data_stage_4__5061_, data_stage_4__5060_, data_stage_4__5059_, data_stage_4__5058_, data_stage_4__5057_, data_stage_4__5056_, data_stage_4__5055_, data_stage_4__5054_, data_stage_4__5053_, data_stage_4__5052_, data_stage_4__5051_, data_stage_4__5050_, data_stage_4__5049_, data_stage_4__5048_, data_stage_4__5047_, data_stage_4__5046_, data_stage_4__5045_, data_stage_4__5044_, data_stage_4__5043_, data_stage_4__5042_, data_stage_4__5041_, data_stage_4__5040_, data_stage_4__5039_, data_stage_4__5038_, data_stage_4__5037_, data_stage_4__5036_, data_stage_4__5035_, data_stage_4__5034_, data_stage_4__5033_, data_stage_4__5032_, data_stage_4__5031_, data_stage_4__5030_, data_stage_4__5029_, data_stage_4__5028_, data_stage_4__5027_, data_stage_4__5026_, data_stage_4__5025_, data_stage_4__5024_, data_stage_4__5023_, data_stage_4__5022_, data_stage_4__5021_, data_stage_4__5020_, data_stage_4__5019_, data_stage_4__5018_, data_stage_4__5017_, data_stage_4__5016_, data_stage_4__5015_, data_stage_4__5014_, data_stage_4__5013_, data_stage_4__5012_, data_stage_4__5011_, data_stage_4__5010_, data_stage_4__5009_, data_stage_4__5008_, data_stage_4__5007_, data_stage_4__5006_, data_stage_4__5005_, data_stage_4__5004_, data_stage_4__5003_, data_stage_4__5002_, data_stage_4__5001_, data_stage_4__5000_, data_stage_4__4999_, data_stage_4__4998_, data_stage_4__4997_, data_stage_4__4996_, data_stage_4__4995_, data_stage_4__4994_, data_stage_4__4993_, data_stage_4__4992_, data_stage_4__4991_, data_stage_4__4990_, data_stage_4__4989_, data_stage_4__4988_, data_stage_4__4987_, data_stage_4__4986_, data_stage_4__4985_, data_stage_4__4984_, data_stage_4__4983_, data_stage_4__4982_, data_stage_4__4981_, data_stage_4__4980_, data_stage_4__4979_, data_stage_4__4978_, data_stage_4__4977_, data_stage_4__4976_, data_stage_4__4975_, data_stage_4__4974_, data_stage_4__4973_, data_stage_4__4972_, data_stage_4__4971_, data_stage_4__4970_, data_stage_4__4969_, data_stage_4__4968_, data_stage_4__4967_, data_stage_4__4966_, data_stage_4__4965_, data_stage_4__4964_, data_stage_4__4963_, data_stage_4__4962_, data_stage_4__4961_, data_stage_4__4960_, data_stage_4__4959_, data_stage_4__4958_, data_stage_4__4957_, data_stage_4__4956_, data_stage_4__4955_, data_stage_4__4954_, data_stage_4__4953_, data_stage_4__4952_, data_stage_4__4951_, data_stage_4__4950_, data_stage_4__4949_, data_stage_4__4948_, data_stage_4__4947_, data_stage_4__4946_, data_stage_4__4945_, data_stage_4__4944_, data_stage_4__4943_, data_stage_4__4942_, data_stage_4__4941_, data_stage_4__4940_, data_stage_4__4939_, data_stage_4__4938_, data_stage_4__4937_, data_stage_4__4936_, data_stage_4__4935_, data_stage_4__4934_, data_stage_4__4933_, data_stage_4__4932_, data_stage_4__4931_, data_stage_4__4930_, data_stage_4__4929_, data_stage_4__4928_, data_stage_4__4927_, data_stage_4__4926_, data_stage_4__4925_, data_stage_4__4924_, data_stage_4__4923_, data_stage_4__4922_, data_stage_4__4921_, data_stage_4__4920_, data_stage_4__4919_, data_stage_4__4918_, data_stage_4__4917_, data_stage_4__4916_, data_stage_4__4915_, data_stage_4__4914_, data_stage_4__4913_, data_stage_4__4912_, data_stage_4__4911_, data_stage_4__4910_, data_stage_4__4909_, data_stage_4__4908_, data_stage_4__4907_, data_stage_4__4906_, data_stage_4__4905_, data_stage_4__4904_, data_stage_4__4903_, data_stage_4__4902_, data_stage_4__4901_, data_stage_4__4900_, data_stage_4__4899_, data_stage_4__4898_, data_stage_4__4897_, data_stage_4__4896_, data_stage_4__4895_, data_stage_4__4894_, data_stage_4__4893_, data_stage_4__4892_, data_stage_4__4891_, data_stage_4__4890_, data_stage_4__4889_, data_stage_4__4888_, data_stage_4__4887_, data_stage_4__4886_, data_stage_4__4885_, data_stage_4__4884_, data_stage_4__4883_, data_stage_4__4882_, data_stage_4__4881_, data_stage_4__4880_, data_stage_4__4879_, data_stage_4__4878_, data_stage_4__4877_, data_stage_4__4876_, data_stage_4__4875_, data_stage_4__4874_, data_stage_4__4873_, data_stage_4__4872_, data_stage_4__4871_, data_stage_4__4870_, data_stage_4__4869_, data_stage_4__4868_, data_stage_4__4867_, data_stage_4__4866_, data_stage_4__4865_, data_stage_4__4864_, data_stage_4__4863_, data_stage_4__4862_, data_stage_4__4861_, data_stage_4__4860_, data_stage_4__4859_, data_stage_4__4858_, data_stage_4__4857_, data_stage_4__4856_, data_stage_4__4855_, data_stage_4__4854_, data_stage_4__4853_, data_stage_4__4852_, data_stage_4__4851_, data_stage_4__4850_, data_stage_4__4849_, data_stage_4__4848_, data_stage_4__4847_, data_stage_4__4846_, data_stage_4__4845_, data_stage_4__4844_, data_stage_4__4843_, data_stage_4__4842_, data_stage_4__4841_, data_stage_4__4840_, data_stage_4__4839_, data_stage_4__4838_, data_stage_4__4837_, data_stage_4__4836_, data_stage_4__4835_, data_stage_4__4834_, data_stage_4__4833_, data_stage_4__4832_, data_stage_4__4831_, data_stage_4__4830_, data_stage_4__4829_, data_stage_4__4828_, data_stage_4__4827_, data_stage_4__4826_, data_stage_4__4825_, data_stage_4__4824_, data_stage_4__4823_, data_stage_4__4822_, data_stage_4__4821_, data_stage_4__4820_, data_stage_4__4819_, data_stage_4__4818_, data_stage_4__4817_, data_stage_4__4816_, data_stage_4__4815_, data_stage_4__4814_, data_stage_4__4813_, data_stage_4__4812_, data_stage_4__4811_, data_stage_4__4810_, data_stage_4__4809_, data_stage_4__4808_, data_stage_4__4807_, data_stage_4__4806_, data_stage_4__4805_, data_stage_4__4804_, data_stage_4__4803_, data_stage_4__4802_, data_stage_4__4801_, data_stage_4__4800_, data_stage_4__4799_, data_stage_4__4798_, data_stage_4__4797_, data_stage_4__4796_, data_stage_4__4795_, data_stage_4__4794_, data_stage_4__4793_, data_stage_4__4792_, data_stage_4__4791_, data_stage_4__4790_, data_stage_4__4789_, data_stage_4__4788_, data_stage_4__4787_, data_stage_4__4786_, data_stage_4__4785_, data_stage_4__4784_, data_stage_4__4783_, data_stage_4__4782_, data_stage_4__4781_, data_stage_4__4780_, data_stage_4__4779_, data_stage_4__4778_, data_stage_4__4777_, data_stage_4__4776_, data_stage_4__4775_, data_stage_4__4774_, data_stage_4__4773_, data_stage_4__4772_, data_stage_4__4771_, data_stage_4__4770_, data_stage_4__4769_, data_stage_4__4768_, data_stage_4__4767_, data_stage_4__4766_, data_stage_4__4765_, data_stage_4__4764_, data_stage_4__4763_, data_stage_4__4762_, data_stage_4__4761_, data_stage_4__4760_, data_stage_4__4759_, data_stage_4__4758_, data_stage_4__4757_, data_stage_4__4756_, data_stage_4__4755_, data_stage_4__4754_, data_stage_4__4753_, data_stage_4__4752_, data_stage_4__4751_, data_stage_4__4750_, data_stage_4__4749_, data_stage_4__4748_, data_stage_4__4747_, data_stage_4__4746_, data_stage_4__4745_, data_stage_4__4744_, data_stage_4__4743_, data_stage_4__4742_, data_stage_4__4741_, data_stage_4__4740_, data_stage_4__4739_, data_stage_4__4738_, data_stage_4__4737_, data_stage_4__4736_, data_stage_4__4735_, data_stage_4__4734_, data_stage_4__4733_, data_stage_4__4732_, data_stage_4__4731_, data_stage_4__4730_, data_stage_4__4729_, data_stage_4__4728_, data_stage_4__4727_, data_stage_4__4726_, data_stage_4__4725_, data_stage_4__4724_, data_stage_4__4723_, data_stage_4__4722_, data_stage_4__4721_, data_stage_4__4720_, data_stage_4__4719_, data_stage_4__4718_, data_stage_4__4717_, data_stage_4__4716_, data_stage_4__4715_, data_stage_4__4714_, data_stage_4__4713_, data_stage_4__4712_, data_stage_4__4711_, data_stage_4__4710_, data_stage_4__4709_, data_stage_4__4708_, data_stage_4__4707_, data_stage_4__4706_, data_stage_4__4705_, data_stage_4__4704_, data_stage_4__4703_, data_stage_4__4702_, data_stage_4__4701_, data_stage_4__4700_, data_stage_4__4699_, data_stage_4__4698_, data_stage_4__4697_, data_stage_4__4696_, data_stage_4__4695_, data_stage_4__4694_, data_stage_4__4693_, data_stage_4__4692_, data_stage_4__4691_, data_stage_4__4690_, data_stage_4__4689_, data_stage_4__4688_, data_stage_4__4687_, data_stage_4__4686_, data_stage_4__4685_, data_stage_4__4684_, data_stage_4__4683_, data_stage_4__4682_, data_stage_4__4681_, data_stage_4__4680_, data_stage_4__4679_, data_stage_4__4678_, data_stage_4__4677_, data_stage_4__4676_, data_stage_4__4675_, data_stage_4__4674_, data_stage_4__4673_, data_stage_4__4672_, data_stage_4__4671_, data_stage_4__4670_, data_stage_4__4669_, data_stage_4__4668_, data_stage_4__4667_, data_stage_4__4666_, data_stage_4__4665_, data_stage_4__4664_, data_stage_4__4663_, data_stage_4__4662_, data_stage_4__4661_, data_stage_4__4660_, data_stage_4__4659_, data_stage_4__4658_, data_stage_4__4657_, data_stage_4__4656_, data_stage_4__4655_, data_stage_4__4654_, data_stage_4__4653_, data_stage_4__4652_, data_stage_4__4651_, data_stage_4__4650_, data_stage_4__4649_, data_stage_4__4648_, data_stage_4__4647_, data_stage_4__4646_, data_stage_4__4645_, data_stage_4__4644_, data_stage_4__4643_, data_stage_4__4642_, data_stage_4__4641_, data_stage_4__4640_, data_stage_4__4639_, data_stage_4__4638_, data_stage_4__4637_, data_stage_4__4636_, data_stage_4__4635_, data_stage_4__4634_, data_stage_4__4633_, data_stage_4__4632_, data_stage_4__4631_, data_stage_4__4630_, data_stage_4__4629_, data_stage_4__4628_, data_stage_4__4627_, data_stage_4__4626_, data_stage_4__4625_, data_stage_4__4624_, data_stage_4__4623_, data_stage_4__4622_, data_stage_4__4621_, data_stage_4__4620_, data_stage_4__4619_, data_stage_4__4618_, data_stage_4__4617_, data_stage_4__4616_, data_stage_4__4615_, data_stage_4__4614_, data_stage_4__4613_, data_stage_4__4612_, data_stage_4__4611_, data_stage_4__4610_, data_stage_4__4609_, data_stage_4__4608_, data_stage_4__4607_, data_stage_4__4606_, data_stage_4__4605_, data_stage_4__4604_, data_stage_4__4603_, data_stage_4__4602_, data_stage_4__4601_, data_stage_4__4600_, data_stage_4__4599_, data_stage_4__4598_, data_stage_4__4597_, data_stage_4__4596_, data_stage_4__4595_, data_stage_4__4594_, data_stage_4__4593_, data_stage_4__4592_, data_stage_4__4591_, data_stage_4__4590_, data_stage_4__4589_, data_stage_4__4588_, data_stage_4__4587_, data_stage_4__4586_, data_stage_4__4585_, data_stage_4__4584_, data_stage_4__4583_, data_stage_4__4582_, data_stage_4__4581_, data_stage_4__4580_, data_stage_4__4579_, data_stage_4__4578_, data_stage_4__4577_, data_stage_4__4576_, data_stage_4__4575_, data_stage_4__4574_, data_stage_4__4573_, data_stage_4__4572_, data_stage_4__4571_, data_stage_4__4570_, data_stage_4__4569_, data_stage_4__4568_, data_stage_4__4567_, data_stage_4__4566_, data_stage_4__4565_, data_stage_4__4564_, data_stage_4__4563_, data_stage_4__4562_, data_stage_4__4561_, data_stage_4__4560_, data_stage_4__4559_, data_stage_4__4558_, data_stage_4__4557_, data_stage_4__4556_, data_stage_4__4555_, data_stage_4__4554_, data_stage_4__4553_, data_stage_4__4552_, data_stage_4__4551_, data_stage_4__4550_, data_stage_4__4549_, data_stage_4__4548_, data_stage_4__4547_, data_stage_4__4546_, data_stage_4__4545_, data_stage_4__4544_, data_stage_4__4543_, data_stage_4__4542_, data_stage_4__4541_, data_stage_4__4540_, data_stage_4__4539_, data_stage_4__4538_, data_stage_4__4537_, data_stage_4__4536_, data_stage_4__4535_, data_stage_4__4534_, data_stage_4__4533_, data_stage_4__4532_, data_stage_4__4531_, data_stage_4__4530_, data_stage_4__4529_, data_stage_4__4528_, data_stage_4__4527_, data_stage_4__4526_, data_stage_4__4525_, data_stage_4__4524_, data_stage_4__4523_, data_stage_4__4522_, data_stage_4__4521_, data_stage_4__4520_, data_stage_4__4519_, data_stage_4__4518_, data_stage_4__4517_, data_stage_4__4516_, data_stage_4__4515_, data_stage_4__4514_, data_stage_4__4513_, data_stage_4__4512_, data_stage_4__4511_, data_stage_4__4510_, data_stage_4__4509_, data_stage_4__4508_, data_stage_4__4507_, data_stage_4__4506_, data_stage_4__4505_, data_stage_4__4504_, data_stage_4__4503_, data_stage_4__4502_, data_stage_4__4501_, data_stage_4__4500_, data_stage_4__4499_, data_stage_4__4498_, data_stage_4__4497_, data_stage_4__4496_, data_stage_4__4495_, data_stage_4__4494_, data_stage_4__4493_, data_stage_4__4492_, data_stage_4__4491_, data_stage_4__4490_, data_stage_4__4489_, data_stage_4__4488_, data_stage_4__4487_, data_stage_4__4486_, data_stage_4__4485_, data_stage_4__4484_, data_stage_4__4483_, data_stage_4__4482_, data_stage_4__4481_, data_stage_4__4480_, data_stage_4__4479_, data_stage_4__4478_, data_stage_4__4477_, data_stage_4__4476_, data_stage_4__4475_, data_stage_4__4474_, data_stage_4__4473_, data_stage_4__4472_, data_stage_4__4471_, data_stage_4__4470_, data_stage_4__4469_, data_stage_4__4468_, data_stage_4__4467_, data_stage_4__4466_, data_stage_4__4465_, data_stage_4__4464_, data_stage_4__4463_, data_stage_4__4462_, data_stage_4__4461_, data_stage_4__4460_, data_stage_4__4459_, data_stage_4__4458_, data_stage_4__4457_, data_stage_4__4456_, data_stage_4__4455_, data_stage_4__4454_, data_stage_4__4453_, data_stage_4__4452_, data_stage_4__4451_, data_stage_4__4450_, data_stage_4__4449_, data_stage_4__4448_, data_stage_4__4447_, data_stage_4__4446_, data_stage_4__4445_, data_stage_4__4444_, data_stage_4__4443_, data_stage_4__4442_, data_stage_4__4441_, data_stage_4__4440_, data_stage_4__4439_, data_stage_4__4438_, data_stage_4__4437_, data_stage_4__4436_, data_stage_4__4435_, data_stage_4__4434_, data_stage_4__4433_, data_stage_4__4432_, data_stage_4__4431_, data_stage_4__4430_, data_stage_4__4429_, data_stage_4__4428_, data_stage_4__4427_, data_stage_4__4426_, data_stage_4__4425_, data_stage_4__4424_, data_stage_4__4423_, data_stage_4__4422_, data_stage_4__4421_, data_stage_4__4420_, data_stage_4__4419_, data_stage_4__4418_, data_stage_4__4417_, data_stage_4__4416_, data_stage_4__4415_, data_stage_4__4414_, data_stage_4__4413_, data_stage_4__4412_, data_stage_4__4411_, data_stage_4__4410_, data_stage_4__4409_, data_stage_4__4408_, data_stage_4__4407_, data_stage_4__4406_, data_stage_4__4405_, data_stage_4__4404_, data_stage_4__4403_, data_stage_4__4402_, data_stage_4__4401_, data_stage_4__4400_, data_stage_4__4399_, data_stage_4__4398_, data_stage_4__4397_, data_stage_4__4396_, data_stage_4__4395_, data_stage_4__4394_, data_stage_4__4393_, data_stage_4__4392_, data_stage_4__4391_, data_stage_4__4390_, data_stage_4__4389_, data_stage_4__4388_, data_stage_4__4387_, data_stage_4__4386_, data_stage_4__4385_, data_stage_4__4384_, data_stage_4__4383_, data_stage_4__4382_, data_stage_4__4381_, data_stage_4__4380_, data_stage_4__4379_, data_stage_4__4378_, data_stage_4__4377_, data_stage_4__4376_, data_stage_4__4375_, data_stage_4__4374_, data_stage_4__4373_, data_stage_4__4372_, data_stage_4__4371_, data_stage_4__4370_, data_stage_4__4369_, data_stage_4__4368_, data_stage_4__4367_, data_stage_4__4366_, data_stage_4__4365_, data_stage_4__4364_, data_stage_4__4363_, data_stage_4__4362_, data_stage_4__4361_, data_stage_4__4360_, data_stage_4__4359_, data_stage_4__4358_, data_stage_4__4357_, data_stage_4__4356_, data_stage_4__4355_, data_stage_4__4354_, data_stage_4__4353_, data_stage_4__4352_, data_stage_4__4351_, data_stage_4__4350_, data_stage_4__4349_, data_stage_4__4348_, data_stage_4__4347_, data_stage_4__4346_, data_stage_4__4345_, data_stage_4__4344_, data_stage_4__4343_, data_stage_4__4342_, data_stage_4__4341_, data_stage_4__4340_, data_stage_4__4339_, data_stage_4__4338_, data_stage_4__4337_, data_stage_4__4336_, data_stage_4__4335_, data_stage_4__4334_, data_stage_4__4333_, data_stage_4__4332_, data_stage_4__4331_, data_stage_4__4330_, data_stage_4__4329_, data_stage_4__4328_, data_stage_4__4327_, data_stage_4__4326_, data_stage_4__4325_, data_stage_4__4324_, data_stage_4__4323_, data_stage_4__4322_, data_stage_4__4321_, data_stage_4__4320_, data_stage_4__4319_, data_stage_4__4318_, data_stage_4__4317_, data_stage_4__4316_, data_stage_4__4315_, data_stage_4__4314_, data_stage_4__4313_, data_stage_4__4312_, data_stage_4__4311_, data_stage_4__4310_, data_stage_4__4309_, data_stage_4__4308_, data_stage_4__4307_, data_stage_4__4306_, data_stage_4__4305_, data_stage_4__4304_, data_stage_4__4303_, data_stage_4__4302_, data_stage_4__4301_, data_stage_4__4300_, data_stage_4__4299_, data_stage_4__4298_, data_stage_4__4297_, data_stage_4__4296_, data_stage_4__4295_, data_stage_4__4294_, data_stage_4__4293_, data_stage_4__4292_, data_stage_4__4291_, data_stage_4__4290_, data_stage_4__4289_, data_stage_4__4288_, data_stage_4__4287_, data_stage_4__4286_, data_stage_4__4285_, data_stage_4__4284_, data_stage_4__4283_, data_stage_4__4282_, data_stage_4__4281_, data_stage_4__4280_, data_stage_4__4279_, data_stage_4__4278_, data_stage_4__4277_, data_stage_4__4276_, data_stage_4__4275_, data_stage_4__4274_, data_stage_4__4273_, data_stage_4__4272_, data_stage_4__4271_, data_stage_4__4270_, data_stage_4__4269_, data_stage_4__4268_, data_stage_4__4267_, data_stage_4__4266_, data_stage_4__4265_, data_stage_4__4264_, data_stage_4__4263_, data_stage_4__4262_, data_stage_4__4261_, data_stage_4__4260_, data_stage_4__4259_, data_stage_4__4258_, data_stage_4__4257_, data_stage_4__4256_, data_stage_4__4255_, data_stage_4__4254_, data_stage_4__4253_, data_stage_4__4252_, data_stage_4__4251_, data_stage_4__4250_, data_stage_4__4249_, data_stage_4__4248_, data_stage_4__4247_, data_stage_4__4246_, data_stage_4__4245_, data_stage_4__4244_, data_stage_4__4243_, data_stage_4__4242_, data_stage_4__4241_, data_stage_4__4240_, data_stage_4__4239_, data_stage_4__4238_, data_stage_4__4237_, data_stage_4__4236_, data_stage_4__4235_, data_stage_4__4234_, data_stage_4__4233_, data_stage_4__4232_, data_stage_4__4231_, data_stage_4__4230_, data_stage_4__4229_, data_stage_4__4228_, data_stage_4__4227_, data_stage_4__4226_, data_stage_4__4225_, data_stage_4__4224_, data_stage_4__4223_, data_stage_4__4222_, data_stage_4__4221_, data_stage_4__4220_, data_stage_4__4219_, data_stage_4__4218_, data_stage_4__4217_, data_stage_4__4216_, data_stage_4__4215_, data_stage_4__4214_, data_stage_4__4213_, data_stage_4__4212_, data_stage_4__4211_, data_stage_4__4210_, data_stage_4__4209_, data_stage_4__4208_, data_stage_4__4207_, data_stage_4__4206_, data_stage_4__4205_, data_stage_4__4204_, data_stage_4__4203_, data_stage_4__4202_, data_stage_4__4201_, data_stage_4__4200_, data_stage_4__4199_, data_stage_4__4198_, data_stage_4__4197_, data_stage_4__4196_, data_stage_4__4195_, data_stage_4__4194_, data_stage_4__4193_, data_stage_4__4192_, data_stage_4__4191_, data_stage_4__4190_, data_stage_4__4189_, data_stage_4__4188_, data_stage_4__4187_, data_stage_4__4186_, data_stage_4__4185_, data_stage_4__4184_, data_stage_4__4183_, data_stage_4__4182_, data_stage_4__4181_, data_stage_4__4180_, data_stage_4__4179_, data_stage_4__4178_, data_stage_4__4177_, data_stage_4__4176_, data_stage_4__4175_, data_stage_4__4174_, data_stage_4__4173_, data_stage_4__4172_, data_stage_4__4171_, data_stage_4__4170_, data_stage_4__4169_, data_stage_4__4168_, data_stage_4__4167_, data_stage_4__4166_, data_stage_4__4165_, data_stage_4__4164_, data_stage_4__4163_, data_stage_4__4162_, data_stage_4__4161_, data_stage_4__4160_, data_stage_4__4159_, data_stage_4__4158_, data_stage_4__4157_, data_stage_4__4156_, data_stage_4__4155_, data_stage_4__4154_, data_stage_4__4153_, data_stage_4__4152_, data_stage_4__4151_, data_stage_4__4150_, data_stage_4__4149_, data_stage_4__4148_, data_stage_4__4147_, data_stage_4__4146_, data_stage_4__4145_, data_stage_4__4144_, data_stage_4__4143_, data_stage_4__4142_, data_stage_4__4141_, data_stage_4__4140_, data_stage_4__4139_, data_stage_4__4138_, data_stage_4__4137_, data_stage_4__4136_, data_stage_4__4135_, data_stage_4__4134_, data_stage_4__4133_, data_stage_4__4132_, data_stage_4__4131_, data_stage_4__4130_, data_stage_4__4129_, data_stage_4__4128_, data_stage_4__4127_, data_stage_4__4126_, data_stage_4__4125_, data_stage_4__4124_, data_stage_4__4123_, data_stage_4__4122_, data_stage_4__4121_, data_stage_4__4120_, data_stage_4__4119_, data_stage_4__4118_, data_stage_4__4117_, data_stage_4__4116_, data_stage_4__4115_, data_stage_4__4114_, data_stage_4__4113_, data_stage_4__4112_, data_stage_4__4111_, data_stage_4__4110_, data_stage_4__4109_, data_stage_4__4108_, data_stage_4__4107_, data_stage_4__4106_, data_stage_4__4105_, data_stage_4__4104_, data_stage_4__4103_, data_stage_4__4102_, data_stage_4__4101_, data_stage_4__4100_, data_stage_4__4099_, data_stage_4__4098_, data_stage_4__4097_, data_stage_4__4096_ }),
    .swap_i(sel_i[4]),
    .data_o({ data_stage_5__8191_, data_stage_5__8190_, data_stage_5__8189_, data_stage_5__8188_, data_stage_5__8187_, data_stage_5__8186_, data_stage_5__8185_, data_stage_5__8184_, data_stage_5__8183_, data_stage_5__8182_, data_stage_5__8181_, data_stage_5__8180_, data_stage_5__8179_, data_stage_5__8178_, data_stage_5__8177_, data_stage_5__8176_, data_stage_5__8175_, data_stage_5__8174_, data_stage_5__8173_, data_stage_5__8172_, data_stage_5__8171_, data_stage_5__8170_, data_stage_5__8169_, data_stage_5__8168_, data_stage_5__8167_, data_stage_5__8166_, data_stage_5__8165_, data_stage_5__8164_, data_stage_5__8163_, data_stage_5__8162_, data_stage_5__8161_, data_stage_5__8160_, data_stage_5__8159_, data_stage_5__8158_, data_stage_5__8157_, data_stage_5__8156_, data_stage_5__8155_, data_stage_5__8154_, data_stage_5__8153_, data_stage_5__8152_, data_stage_5__8151_, data_stage_5__8150_, data_stage_5__8149_, data_stage_5__8148_, data_stage_5__8147_, data_stage_5__8146_, data_stage_5__8145_, data_stage_5__8144_, data_stage_5__8143_, data_stage_5__8142_, data_stage_5__8141_, data_stage_5__8140_, data_stage_5__8139_, data_stage_5__8138_, data_stage_5__8137_, data_stage_5__8136_, data_stage_5__8135_, data_stage_5__8134_, data_stage_5__8133_, data_stage_5__8132_, data_stage_5__8131_, data_stage_5__8130_, data_stage_5__8129_, data_stage_5__8128_, data_stage_5__8127_, data_stage_5__8126_, data_stage_5__8125_, data_stage_5__8124_, data_stage_5__8123_, data_stage_5__8122_, data_stage_5__8121_, data_stage_5__8120_, data_stage_5__8119_, data_stage_5__8118_, data_stage_5__8117_, data_stage_5__8116_, data_stage_5__8115_, data_stage_5__8114_, data_stage_5__8113_, data_stage_5__8112_, data_stage_5__8111_, data_stage_5__8110_, data_stage_5__8109_, data_stage_5__8108_, data_stage_5__8107_, data_stage_5__8106_, data_stage_5__8105_, data_stage_5__8104_, data_stage_5__8103_, data_stage_5__8102_, data_stage_5__8101_, data_stage_5__8100_, data_stage_5__8099_, data_stage_5__8098_, data_stage_5__8097_, data_stage_5__8096_, data_stage_5__8095_, data_stage_5__8094_, data_stage_5__8093_, data_stage_5__8092_, data_stage_5__8091_, data_stage_5__8090_, data_stage_5__8089_, data_stage_5__8088_, data_stage_5__8087_, data_stage_5__8086_, data_stage_5__8085_, data_stage_5__8084_, data_stage_5__8083_, data_stage_5__8082_, data_stage_5__8081_, data_stage_5__8080_, data_stage_5__8079_, data_stage_5__8078_, data_stage_5__8077_, data_stage_5__8076_, data_stage_5__8075_, data_stage_5__8074_, data_stage_5__8073_, data_stage_5__8072_, data_stage_5__8071_, data_stage_5__8070_, data_stage_5__8069_, data_stage_5__8068_, data_stage_5__8067_, data_stage_5__8066_, data_stage_5__8065_, data_stage_5__8064_, data_stage_5__8063_, data_stage_5__8062_, data_stage_5__8061_, data_stage_5__8060_, data_stage_5__8059_, data_stage_5__8058_, data_stage_5__8057_, data_stage_5__8056_, data_stage_5__8055_, data_stage_5__8054_, data_stage_5__8053_, data_stage_5__8052_, data_stage_5__8051_, data_stage_5__8050_, data_stage_5__8049_, data_stage_5__8048_, data_stage_5__8047_, data_stage_5__8046_, data_stage_5__8045_, data_stage_5__8044_, data_stage_5__8043_, data_stage_5__8042_, data_stage_5__8041_, data_stage_5__8040_, data_stage_5__8039_, data_stage_5__8038_, data_stage_5__8037_, data_stage_5__8036_, data_stage_5__8035_, data_stage_5__8034_, data_stage_5__8033_, data_stage_5__8032_, data_stage_5__8031_, data_stage_5__8030_, data_stage_5__8029_, data_stage_5__8028_, data_stage_5__8027_, data_stage_5__8026_, data_stage_5__8025_, data_stage_5__8024_, data_stage_5__8023_, data_stage_5__8022_, data_stage_5__8021_, data_stage_5__8020_, data_stage_5__8019_, data_stage_5__8018_, data_stage_5__8017_, data_stage_5__8016_, data_stage_5__8015_, data_stage_5__8014_, data_stage_5__8013_, data_stage_5__8012_, data_stage_5__8011_, data_stage_5__8010_, data_stage_5__8009_, data_stage_5__8008_, data_stage_5__8007_, data_stage_5__8006_, data_stage_5__8005_, data_stage_5__8004_, data_stage_5__8003_, data_stage_5__8002_, data_stage_5__8001_, data_stage_5__8000_, data_stage_5__7999_, data_stage_5__7998_, data_stage_5__7997_, data_stage_5__7996_, data_stage_5__7995_, data_stage_5__7994_, data_stage_5__7993_, data_stage_5__7992_, data_stage_5__7991_, data_stage_5__7990_, data_stage_5__7989_, data_stage_5__7988_, data_stage_5__7987_, data_stage_5__7986_, data_stage_5__7985_, data_stage_5__7984_, data_stage_5__7983_, data_stage_5__7982_, data_stage_5__7981_, data_stage_5__7980_, data_stage_5__7979_, data_stage_5__7978_, data_stage_5__7977_, data_stage_5__7976_, data_stage_5__7975_, data_stage_5__7974_, data_stage_5__7973_, data_stage_5__7972_, data_stage_5__7971_, data_stage_5__7970_, data_stage_5__7969_, data_stage_5__7968_, data_stage_5__7967_, data_stage_5__7966_, data_stage_5__7965_, data_stage_5__7964_, data_stage_5__7963_, data_stage_5__7962_, data_stage_5__7961_, data_stage_5__7960_, data_stage_5__7959_, data_stage_5__7958_, data_stage_5__7957_, data_stage_5__7956_, data_stage_5__7955_, data_stage_5__7954_, data_stage_5__7953_, data_stage_5__7952_, data_stage_5__7951_, data_stage_5__7950_, data_stage_5__7949_, data_stage_5__7948_, data_stage_5__7947_, data_stage_5__7946_, data_stage_5__7945_, data_stage_5__7944_, data_stage_5__7943_, data_stage_5__7942_, data_stage_5__7941_, data_stage_5__7940_, data_stage_5__7939_, data_stage_5__7938_, data_stage_5__7937_, data_stage_5__7936_, data_stage_5__7935_, data_stage_5__7934_, data_stage_5__7933_, data_stage_5__7932_, data_stage_5__7931_, data_stage_5__7930_, data_stage_5__7929_, data_stage_5__7928_, data_stage_5__7927_, data_stage_5__7926_, data_stage_5__7925_, data_stage_5__7924_, data_stage_5__7923_, data_stage_5__7922_, data_stage_5__7921_, data_stage_5__7920_, data_stage_5__7919_, data_stage_5__7918_, data_stage_5__7917_, data_stage_5__7916_, data_stage_5__7915_, data_stage_5__7914_, data_stage_5__7913_, data_stage_5__7912_, data_stage_5__7911_, data_stage_5__7910_, data_stage_5__7909_, data_stage_5__7908_, data_stage_5__7907_, data_stage_5__7906_, data_stage_5__7905_, data_stage_5__7904_, data_stage_5__7903_, data_stage_5__7902_, data_stage_5__7901_, data_stage_5__7900_, data_stage_5__7899_, data_stage_5__7898_, data_stage_5__7897_, data_stage_5__7896_, data_stage_5__7895_, data_stage_5__7894_, data_stage_5__7893_, data_stage_5__7892_, data_stage_5__7891_, data_stage_5__7890_, data_stage_5__7889_, data_stage_5__7888_, data_stage_5__7887_, data_stage_5__7886_, data_stage_5__7885_, data_stage_5__7884_, data_stage_5__7883_, data_stage_5__7882_, data_stage_5__7881_, data_stage_5__7880_, data_stage_5__7879_, data_stage_5__7878_, data_stage_5__7877_, data_stage_5__7876_, data_stage_5__7875_, data_stage_5__7874_, data_stage_5__7873_, data_stage_5__7872_, data_stage_5__7871_, data_stage_5__7870_, data_stage_5__7869_, data_stage_5__7868_, data_stage_5__7867_, data_stage_5__7866_, data_stage_5__7865_, data_stage_5__7864_, data_stage_5__7863_, data_stage_5__7862_, data_stage_5__7861_, data_stage_5__7860_, data_stage_5__7859_, data_stage_5__7858_, data_stage_5__7857_, data_stage_5__7856_, data_stage_5__7855_, data_stage_5__7854_, data_stage_5__7853_, data_stage_5__7852_, data_stage_5__7851_, data_stage_5__7850_, data_stage_5__7849_, data_stage_5__7848_, data_stage_5__7847_, data_stage_5__7846_, data_stage_5__7845_, data_stage_5__7844_, data_stage_5__7843_, data_stage_5__7842_, data_stage_5__7841_, data_stage_5__7840_, data_stage_5__7839_, data_stage_5__7838_, data_stage_5__7837_, data_stage_5__7836_, data_stage_5__7835_, data_stage_5__7834_, data_stage_5__7833_, data_stage_5__7832_, data_stage_5__7831_, data_stage_5__7830_, data_stage_5__7829_, data_stage_5__7828_, data_stage_5__7827_, data_stage_5__7826_, data_stage_5__7825_, data_stage_5__7824_, data_stage_5__7823_, data_stage_5__7822_, data_stage_5__7821_, data_stage_5__7820_, data_stage_5__7819_, data_stage_5__7818_, data_stage_5__7817_, data_stage_5__7816_, data_stage_5__7815_, data_stage_5__7814_, data_stage_5__7813_, data_stage_5__7812_, data_stage_5__7811_, data_stage_5__7810_, data_stage_5__7809_, data_stage_5__7808_, data_stage_5__7807_, data_stage_5__7806_, data_stage_5__7805_, data_stage_5__7804_, data_stage_5__7803_, data_stage_5__7802_, data_stage_5__7801_, data_stage_5__7800_, data_stage_5__7799_, data_stage_5__7798_, data_stage_5__7797_, data_stage_5__7796_, data_stage_5__7795_, data_stage_5__7794_, data_stage_5__7793_, data_stage_5__7792_, data_stage_5__7791_, data_stage_5__7790_, data_stage_5__7789_, data_stage_5__7788_, data_stage_5__7787_, data_stage_5__7786_, data_stage_5__7785_, data_stage_5__7784_, data_stage_5__7783_, data_stage_5__7782_, data_stage_5__7781_, data_stage_5__7780_, data_stage_5__7779_, data_stage_5__7778_, data_stage_5__7777_, data_stage_5__7776_, data_stage_5__7775_, data_stage_5__7774_, data_stage_5__7773_, data_stage_5__7772_, data_stage_5__7771_, data_stage_5__7770_, data_stage_5__7769_, data_stage_5__7768_, data_stage_5__7767_, data_stage_5__7766_, data_stage_5__7765_, data_stage_5__7764_, data_stage_5__7763_, data_stage_5__7762_, data_stage_5__7761_, data_stage_5__7760_, data_stage_5__7759_, data_stage_5__7758_, data_stage_5__7757_, data_stage_5__7756_, data_stage_5__7755_, data_stage_5__7754_, data_stage_5__7753_, data_stage_5__7752_, data_stage_5__7751_, data_stage_5__7750_, data_stage_5__7749_, data_stage_5__7748_, data_stage_5__7747_, data_stage_5__7746_, data_stage_5__7745_, data_stage_5__7744_, data_stage_5__7743_, data_stage_5__7742_, data_stage_5__7741_, data_stage_5__7740_, data_stage_5__7739_, data_stage_5__7738_, data_stage_5__7737_, data_stage_5__7736_, data_stage_5__7735_, data_stage_5__7734_, data_stage_5__7733_, data_stage_5__7732_, data_stage_5__7731_, data_stage_5__7730_, data_stage_5__7729_, data_stage_5__7728_, data_stage_5__7727_, data_stage_5__7726_, data_stage_5__7725_, data_stage_5__7724_, data_stage_5__7723_, data_stage_5__7722_, data_stage_5__7721_, data_stage_5__7720_, data_stage_5__7719_, data_stage_5__7718_, data_stage_5__7717_, data_stage_5__7716_, data_stage_5__7715_, data_stage_5__7714_, data_stage_5__7713_, data_stage_5__7712_, data_stage_5__7711_, data_stage_5__7710_, data_stage_5__7709_, data_stage_5__7708_, data_stage_5__7707_, data_stage_5__7706_, data_stage_5__7705_, data_stage_5__7704_, data_stage_5__7703_, data_stage_5__7702_, data_stage_5__7701_, data_stage_5__7700_, data_stage_5__7699_, data_stage_5__7698_, data_stage_5__7697_, data_stage_5__7696_, data_stage_5__7695_, data_stage_5__7694_, data_stage_5__7693_, data_stage_5__7692_, data_stage_5__7691_, data_stage_5__7690_, data_stage_5__7689_, data_stage_5__7688_, data_stage_5__7687_, data_stage_5__7686_, data_stage_5__7685_, data_stage_5__7684_, data_stage_5__7683_, data_stage_5__7682_, data_stage_5__7681_, data_stage_5__7680_, data_stage_5__7679_, data_stage_5__7678_, data_stage_5__7677_, data_stage_5__7676_, data_stage_5__7675_, data_stage_5__7674_, data_stage_5__7673_, data_stage_5__7672_, data_stage_5__7671_, data_stage_5__7670_, data_stage_5__7669_, data_stage_5__7668_, data_stage_5__7667_, data_stage_5__7666_, data_stage_5__7665_, data_stage_5__7664_, data_stage_5__7663_, data_stage_5__7662_, data_stage_5__7661_, data_stage_5__7660_, data_stage_5__7659_, data_stage_5__7658_, data_stage_5__7657_, data_stage_5__7656_, data_stage_5__7655_, data_stage_5__7654_, data_stage_5__7653_, data_stage_5__7652_, data_stage_5__7651_, data_stage_5__7650_, data_stage_5__7649_, data_stage_5__7648_, data_stage_5__7647_, data_stage_5__7646_, data_stage_5__7645_, data_stage_5__7644_, data_stage_5__7643_, data_stage_5__7642_, data_stage_5__7641_, data_stage_5__7640_, data_stage_5__7639_, data_stage_5__7638_, data_stage_5__7637_, data_stage_5__7636_, data_stage_5__7635_, data_stage_5__7634_, data_stage_5__7633_, data_stage_5__7632_, data_stage_5__7631_, data_stage_5__7630_, data_stage_5__7629_, data_stage_5__7628_, data_stage_5__7627_, data_stage_5__7626_, data_stage_5__7625_, data_stage_5__7624_, data_stage_5__7623_, data_stage_5__7622_, data_stage_5__7621_, data_stage_5__7620_, data_stage_5__7619_, data_stage_5__7618_, data_stage_5__7617_, data_stage_5__7616_, data_stage_5__7615_, data_stage_5__7614_, data_stage_5__7613_, data_stage_5__7612_, data_stage_5__7611_, data_stage_5__7610_, data_stage_5__7609_, data_stage_5__7608_, data_stage_5__7607_, data_stage_5__7606_, data_stage_5__7605_, data_stage_5__7604_, data_stage_5__7603_, data_stage_5__7602_, data_stage_5__7601_, data_stage_5__7600_, data_stage_5__7599_, data_stage_5__7598_, data_stage_5__7597_, data_stage_5__7596_, data_stage_5__7595_, data_stage_5__7594_, data_stage_5__7593_, data_stage_5__7592_, data_stage_5__7591_, data_stage_5__7590_, data_stage_5__7589_, data_stage_5__7588_, data_stage_5__7587_, data_stage_5__7586_, data_stage_5__7585_, data_stage_5__7584_, data_stage_5__7583_, data_stage_5__7582_, data_stage_5__7581_, data_stage_5__7580_, data_stage_5__7579_, data_stage_5__7578_, data_stage_5__7577_, data_stage_5__7576_, data_stage_5__7575_, data_stage_5__7574_, data_stage_5__7573_, data_stage_5__7572_, data_stage_5__7571_, data_stage_5__7570_, data_stage_5__7569_, data_stage_5__7568_, data_stage_5__7567_, data_stage_5__7566_, data_stage_5__7565_, data_stage_5__7564_, data_stage_5__7563_, data_stage_5__7562_, data_stage_5__7561_, data_stage_5__7560_, data_stage_5__7559_, data_stage_5__7558_, data_stage_5__7557_, data_stage_5__7556_, data_stage_5__7555_, data_stage_5__7554_, data_stage_5__7553_, data_stage_5__7552_, data_stage_5__7551_, data_stage_5__7550_, data_stage_5__7549_, data_stage_5__7548_, data_stage_5__7547_, data_stage_5__7546_, data_stage_5__7545_, data_stage_5__7544_, data_stage_5__7543_, data_stage_5__7542_, data_stage_5__7541_, data_stage_5__7540_, data_stage_5__7539_, data_stage_5__7538_, data_stage_5__7537_, data_stage_5__7536_, data_stage_5__7535_, data_stage_5__7534_, data_stage_5__7533_, data_stage_5__7532_, data_stage_5__7531_, data_stage_5__7530_, data_stage_5__7529_, data_stage_5__7528_, data_stage_5__7527_, data_stage_5__7526_, data_stage_5__7525_, data_stage_5__7524_, data_stage_5__7523_, data_stage_5__7522_, data_stage_5__7521_, data_stage_5__7520_, data_stage_5__7519_, data_stage_5__7518_, data_stage_5__7517_, data_stage_5__7516_, data_stage_5__7515_, data_stage_5__7514_, data_stage_5__7513_, data_stage_5__7512_, data_stage_5__7511_, data_stage_5__7510_, data_stage_5__7509_, data_stage_5__7508_, data_stage_5__7507_, data_stage_5__7506_, data_stage_5__7505_, data_stage_5__7504_, data_stage_5__7503_, data_stage_5__7502_, data_stage_5__7501_, data_stage_5__7500_, data_stage_5__7499_, data_stage_5__7498_, data_stage_5__7497_, data_stage_5__7496_, data_stage_5__7495_, data_stage_5__7494_, data_stage_5__7493_, data_stage_5__7492_, data_stage_5__7491_, data_stage_5__7490_, data_stage_5__7489_, data_stage_5__7488_, data_stage_5__7487_, data_stage_5__7486_, data_stage_5__7485_, data_stage_5__7484_, data_stage_5__7483_, data_stage_5__7482_, data_stage_5__7481_, data_stage_5__7480_, data_stage_5__7479_, data_stage_5__7478_, data_stage_5__7477_, data_stage_5__7476_, data_stage_5__7475_, data_stage_5__7474_, data_stage_5__7473_, data_stage_5__7472_, data_stage_5__7471_, data_stage_5__7470_, data_stage_5__7469_, data_stage_5__7468_, data_stage_5__7467_, data_stage_5__7466_, data_stage_5__7465_, data_stage_5__7464_, data_stage_5__7463_, data_stage_5__7462_, data_stage_5__7461_, data_stage_5__7460_, data_stage_5__7459_, data_stage_5__7458_, data_stage_5__7457_, data_stage_5__7456_, data_stage_5__7455_, data_stage_5__7454_, data_stage_5__7453_, data_stage_5__7452_, data_stage_5__7451_, data_stage_5__7450_, data_stage_5__7449_, data_stage_5__7448_, data_stage_5__7447_, data_stage_5__7446_, data_stage_5__7445_, data_stage_5__7444_, data_stage_5__7443_, data_stage_5__7442_, data_stage_5__7441_, data_stage_5__7440_, data_stage_5__7439_, data_stage_5__7438_, data_stage_5__7437_, data_stage_5__7436_, data_stage_5__7435_, data_stage_5__7434_, data_stage_5__7433_, data_stage_5__7432_, data_stage_5__7431_, data_stage_5__7430_, data_stage_5__7429_, data_stage_5__7428_, data_stage_5__7427_, data_stage_5__7426_, data_stage_5__7425_, data_stage_5__7424_, data_stage_5__7423_, data_stage_5__7422_, data_stage_5__7421_, data_stage_5__7420_, data_stage_5__7419_, data_stage_5__7418_, data_stage_5__7417_, data_stage_5__7416_, data_stage_5__7415_, data_stage_5__7414_, data_stage_5__7413_, data_stage_5__7412_, data_stage_5__7411_, data_stage_5__7410_, data_stage_5__7409_, data_stage_5__7408_, data_stage_5__7407_, data_stage_5__7406_, data_stage_5__7405_, data_stage_5__7404_, data_stage_5__7403_, data_stage_5__7402_, data_stage_5__7401_, data_stage_5__7400_, data_stage_5__7399_, data_stage_5__7398_, data_stage_5__7397_, data_stage_5__7396_, data_stage_5__7395_, data_stage_5__7394_, data_stage_5__7393_, data_stage_5__7392_, data_stage_5__7391_, data_stage_5__7390_, data_stage_5__7389_, data_stage_5__7388_, data_stage_5__7387_, data_stage_5__7386_, data_stage_5__7385_, data_stage_5__7384_, data_stage_5__7383_, data_stage_5__7382_, data_stage_5__7381_, data_stage_5__7380_, data_stage_5__7379_, data_stage_5__7378_, data_stage_5__7377_, data_stage_5__7376_, data_stage_5__7375_, data_stage_5__7374_, data_stage_5__7373_, data_stage_5__7372_, data_stage_5__7371_, data_stage_5__7370_, data_stage_5__7369_, data_stage_5__7368_, data_stage_5__7367_, data_stage_5__7366_, data_stage_5__7365_, data_stage_5__7364_, data_stage_5__7363_, data_stage_5__7362_, data_stage_5__7361_, data_stage_5__7360_, data_stage_5__7359_, data_stage_5__7358_, data_stage_5__7357_, data_stage_5__7356_, data_stage_5__7355_, data_stage_5__7354_, data_stage_5__7353_, data_stage_5__7352_, data_stage_5__7351_, data_stage_5__7350_, data_stage_5__7349_, data_stage_5__7348_, data_stage_5__7347_, data_stage_5__7346_, data_stage_5__7345_, data_stage_5__7344_, data_stage_5__7343_, data_stage_5__7342_, data_stage_5__7341_, data_stage_5__7340_, data_stage_5__7339_, data_stage_5__7338_, data_stage_5__7337_, data_stage_5__7336_, data_stage_5__7335_, data_stage_5__7334_, data_stage_5__7333_, data_stage_5__7332_, data_stage_5__7331_, data_stage_5__7330_, data_stage_5__7329_, data_stage_5__7328_, data_stage_5__7327_, data_stage_5__7326_, data_stage_5__7325_, data_stage_5__7324_, data_stage_5__7323_, data_stage_5__7322_, data_stage_5__7321_, data_stage_5__7320_, data_stage_5__7319_, data_stage_5__7318_, data_stage_5__7317_, data_stage_5__7316_, data_stage_5__7315_, data_stage_5__7314_, data_stage_5__7313_, data_stage_5__7312_, data_stage_5__7311_, data_stage_5__7310_, data_stage_5__7309_, data_stage_5__7308_, data_stage_5__7307_, data_stage_5__7306_, data_stage_5__7305_, data_stage_5__7304_, data_stage_5__7303_, data_stage_5__7302_, data_stage_5__7301_, data_stage_5__7300_, data_stage_5__7299_, data_stage_5__7298_, data_stage_5__7297_, data_stage_5__7296_, data_stage_5__7295_, data_stage_5__7294_, data_stage_5__7293_, data_stage_5__7292_, data_stage_5__7291_, data_stage_5__7290_, data_stage_5__7289_, data_stage_5__7288_, data_stage_5__7287_, data_stage_5__7286_, data_stage_5__7285_, data_stage_5__7284_, data_stage_5__7283_, data_stage_5__7282_, data_stage_5__7281_, data_stage_5__7280_, data_stage_5__7279_, data_stage_5__7278_, data_stage_5__7277_, data_stage_5__7276_, data_stage_5__7275_, data_stage_5__7274_, data_stage_5__7273_, data_stage_5__7272_, data_stage_5__7271_, data_stage_5__7270_, data_stage_5__7269_, data_stage_5__7268_, data_stage_5__7267_, data_stage_5__7266_, data_stage_5__7265_, data_stage_5__7264_, data_stage_5__7263_, data_stage_5__7262_, data_stage_5__7261_, data_stage_5__7260_, data_stage_5__7259_, data_stage_5__7258_, data_stage_5__7257_, data_stage_5__7256_, data_stage_5__7255_, data_stage_5__7254_, data_stage_5__7253_, data_stage_5__7252_, data_stage_5__7251_, data_stage_5__7250_, data_stage_5__7249_, data_stage_5__7248_, data_stage_5__7247_, data_stage_5__7246_, data_stage_5__7245_, data_stage_5__7244_, data_stage_5__7243_, data_stage_5__7242_, data_stage_5__7241_, data_stage_5__7240_, data_stage_5__7239_, data_stage_5__7238_, data_stage_5__7237_, data_stage_5__7236_, data_stage_5__7235_, data_stage_5__7234_, data_stage_5__7233_, data_stage_5__7232_, data_stage_5__7231_, data_stage_5__7230_, data_stage_5__7229_, data_stage_5__7228_, data_stage_5__7227_, data_stage_5__7226_, data_stage_5__7225_, data_stage_5__7224_, data_stage_5__7223_, data_stage_5__7222_, data_stage_5__7221_, data_stage_5__7220_, data_stage_5__7219_, data_stage_5__7218_, data_stage_5__7217_, data_stage_5__7216_, data_stage_5__7215_, data_stage_5__7214_, data_stage_5__7213_, data_stage_5__7212_, data_stage_5__7211_, data_stage_5__7210_, data_stage_5__7209_, data_stage_5__7208_, data_stage_5__7207_, data_stage_5__7206_, data_stage_5__7205_, data_stage_5__7204_, data_stage_5__7203_, data_stage_5__7202_, data_stage_5__7201_, data_stage_5__7200_, data_stage_5__7199_, data_stage_5__7198_, data_stage_5__7197_, data_stage_5__7196_, data_stage_5__7195_, data_stage_5__7194_, data_stage_5__7193_, data_stage_5__7192_, data_stage_5__7191_, data_stage_5__7190_, data_stage_5__7189_, data_stage_5__7188_, data_stage_5__7187_, data_stage_5__7186_, data_stage_5__7185_, data_stage_5__7184_, data_stage_5__7183_, data_stage_5__7182_, data_stage_5__7181_, data_stage_5__7180_, data_stage_5__7179_, data_stage_5__7178_, data_stage_5__7177_, data_stage_5__7176_, data_stage_5__7175_, data_stage_5__7174_, data_stage_5__7173_, data_stage_5__7172_, data_stage_5__7171_, data_stage_5__7170_, data_stage_5__7169_, data_stage_5__7168_, data_stage_5__7167_, data_stage_5__7166_, data_stage_5__7165_, data_stage_5__7164_, data_stage_5__7163_, data_stage_5__7162_, data_stage_5__7161_, data_stage_5__7160_, data_stage_5__7159_, data_stage_5__7158_, data_stage_5__7157_, data_stage_5__7156_, data_stage_5__7155_, data_stage_5__7154_, data_stage_5__7153_, data_stage_5__7152_, data_stage_5__7151_, data_stage_5__7150_, data_stage_5__7149_, data_stage_5__7148_, data_stage_5__7147_, data_stage_5__7146_, data_stage_5__7145_, data_stage_5__7144_, data_stage_5__7143_, data_stage_5__7142_, data_stage_5__7141_, data_stage_5__7140_, data_stage_5__7139_, data_stage_5__7138_, data_stage_5__7137_, data_stage_5__7136_, data_stage_5__7135_, data_stage_5__7134_, data_stage_5__7133_, data_stage_5__7132_, data_stage_5__7131_, data_stage_5__7130_, data_stage_5__7129_, data_stage_5__7128_, data_stage_5__7127_, data_stage_5__7126_, data_stage_5__7125_, data_stage_5__7124_, data_stage_5__7123_, data_stage_5__7122_, data_stage_5__7121_, data_stage_5__7120_, data_stage_5__7119_, data_stage_5__7118_, data_stage_5__7117_, data_stage_5__7116_, data_stage_5__7115_, data_stage_5__7114_, data_stage_5__7113_, data_stage_5__7112_, data_stage_5__7111_, data_stage_5__7110_, data_stage_5__7109_, data_stage_5__7108_, data_stage_5__7107_, data_stage_5__7106_, data_stage_5__7105_, data_stage_5__7104_, data_stage_5__7103_, data_stage_5__7102_, data_stage_5__7101_, data_stage_5__7100_, data_stage_5__7099_, data_stage_5__7098_, data_stage_5__7097_, data_stage_5__7096_, data_stage_5__7095_, data_stage_5__7094_, data_stage_5__7093_, data_stage_5__7092_, data_stage_5__7091_, data_stage_5__7090_, data_stage_5__7089_, data_stage_5__7088_, data_stage_5__7087_, data_stage_5__7086_, data_stage_5__7085_, data_stage_5__7084_, data_stage_5__7083_, data_stage_5__7082_, data_stage_5__7081_, data_stage_5__7080_, data_stage_5__7079_, data_stage_5__7078_, data_stage_5__7077_, data_stage_5__7076_, data_stage_5__7075_, data_stage_5__7074_, data_stage_5__7073_, data_stage_5__7072_, data_stage_5__7071_, data_stage_5__7070_, data_stage_5__7069_, data_stage_5__7068_, data_stage_5__7067_, data_stage_5__7066_, data_stage_5__7065_, data_stage_5__7064_, data_stage_5__7063_, data_stage_5__7062_, data_stage_5__7061_, data_stage_5__7060_, data_stage_5__7059_, data_stage_5__7058_, data_stage_5__7057_, data_stage_5__7056_, data_stage_5__7055_, data_stage_5__7054_, data_stage_5__7053_, data_stage_5__7052_, data_stage_5__7051_, data_stage_5__7050_, data_stage_5__7049_, data_stage_5__7048_, data_stage_5__7047_, data_stage_5__7046_, data_stage_5__7045_, data_stage_5__7044_, data_stage_5__7043_, data_stage_5__7042_, data_stage_5__7041_, data_stage_5__7040_, data_stage_5__7039_, data_stage_5__7038_, data_stage_5__7037_, data_stage_5__7036_, data_stage_5__7035_, data_stage_5__7034_, data_stage_5__7033_, data_stage_5__7032_, data_stage_5__7031_, data_stage_5__7030_, data_stage_5__7029_, data_stage_5__7028_, data_stage_5__7027_, data_stage_5__7026_, data_stage_5__7025_, data_stage_5__7024_, data_stage_5__7023_, data_stage_5__7022_, data_stage_5__7021_, data_stage_5__7020_, data_stage_5__7019_, data_stage_5__7018_, data_stage_5__7017_, data_stage_5__7016_, data_stage_5__7015_, data_stage_5__7014_, data_stage_5__7013_, data_stage_5__7012_, data_stage_5__7011_, data_stage_5__7010_, data_stage_5__7009_, data_stage_5__7008_, data_stage_5__7007_, data_stage_5__7006_, data_stage_5__7005_, data_stage_5__7004_, data_stage_5__7003_, data_stage_5__7002_, data_stage_5__7001_, data_stage_5__7000_, data_stage_5__6999_, data_stage_5__6998_, data_stage_5__6997_, data_stage_5__6996_, data_stage_5__6995_, data_stage_5__6994_, data_stage_5__6993_, data_stage_5__6992_, data_stage_5__6991_, data_stage_5__6990_, data_stage_5__6989_, data_stage_5__6988_, data_stage_5__6987_, data_stage_5__6986_, data_stage_5__6985_, data_stage_5__6984_, data_stage_5__6983_, data_stage_5__6982_, data_stage_5__6981_, data_stage_5__6980_, data_stage_5__6979_, data_stage_5__6978_, data_stage_5__6977_, data_stage_5__6976_, data_stage_5__6975_, data_stage_5__6974_, data_stage_5__6973_, data_stage_5__6972_, data_stage_5__6971_, data_stage_5__6970_, data_stage_5__6969_, data_stage_5__6968_, data_stage_5__6967_, data_stage_5__6966_, data_stage_5__6965_, data_stage_5__6964_, data_stage_5__6963_, data_stage_5__6962_, data_stage_5__6961_, data_stage_5__6960_, data_stage_5__6959_, data_stage_5__6958_, data_stage_5__6957_, data_stage_5__6956_, data_stage_5__6955_, data_stage_5__6954_, data_stage_5__6953_, data_stage_5__6952_, data_stage_5__6951_, data_stage_5__6950_, data_stage_5__6949_, data_stage_5__6948_, data_stage_5__6947_, data_stage_5__6946_, data_stage_5__6945_, data_stage_5__6944_, data_stage_5__6943_, data_stage_5__6942_, data_stage_5__6941_, data_stage_5__6940_, data_stage_5__6939_, data_stage_5__6938_, data_stage_5__6937_, data_stage_5__6936_, data_stage_5__6935_, data_stage_5__6934_, data_stage_5__6933_, data_stage_5__6932_, data_stage_5__6931_, data_stage_5__6930_, data_stage_5__6929_, data_stage_5__6928_, data_stage_5__6927_, data_stage_5__6926_, data_stage_5__6925_, data_stage_5__6924_, data_stage_5__6923_, data_stage_5__6922_, data_stage_5__6921_, data_stage_5__6920_, data_stage_5__6919_, data_stage_5__6918_, data_stage_5__6917_, data_stage_5__6916_, data_stage_5__6915_, data_stage_5__6914_, data_stage_5__6913_, data_stage_5__6912_, data_stage_5__6911_, data_stage_5__6910_, data_stage_5__6909_, data_stage_5__6908_, data_stage_5__6907_, data_stage_5__6906_, data_stage_5__6905_, data_stage_5__6904_, data_stage_5__6903_, data_stage_5__6902_, data_stage_5__6901_, data_stage_5__6900_, data_stage_5__6899_, data_stage_5__6898_, data_stage_5__6897_, data_stage_5__6896_, data_stage_5__6895_, data_stage_5__6894_, data_stage_5__6893_, data_stage_5__6892_, data_stage_5__6891_, data_stage_5__6890_, data_stage_5__6889_, data_stage_5__6888_, data_stage_5__6887_, data_stage_5__6886_, data_stage_5__6885_, data_stage_5__6884_, data_stage_5__6883_, data_stage_5__6882_, data_stage_5__6881_, data_stage_5__6880_, data_stage_5__6879_, data_stage_5__6878_, data_stage_5__6877_, data_stage_5__6876_, data_stage_5__6875_, data_stage_5__6874_, data_stage_5__6873_, data_stage_5__6872_, data_stage_5__6871_, data_stage_5__6870_, data_stage_5__6869_, data_stage_5__6868_, data_stage_5__6867_, data_stage_5__6866_, data_stage_5__6865_, data_stage_5__6864_, data_stage_5__6863_, data_stage_5__6862_, data_stage_5__6861_, data_stage_5__6860_, data_stage_5__6859_, data_stage_5__6858_, data_stage_5__6857_, data_stage_5__6856_, data_stage_5__6855_, data_stage_5__6854_, data_stage_5__6853_, data_stage_5__6852_, data_stage_5__6851_, data_stage_5__6850_, data_stage_5__6849_, data_stage_5__6848_, data_stage_5__6847_, data_stage_5__6846_, data_stage_5__6845_, data_stage_5__6844_, data_stage_5__6843_, data_stage_5__6842_, data_stage_5__6841_, data_stage_5__6840_, data_stage_5__6839_, data_stage_5__6838_, data_stage_5__6837_, data_stage_5__6836_, data_stage_5__6835_, data_stage_5__6834_, data_stage_5__6833_, data_stage_5__6832_, data_stage_5__6831_, data_stage_5__6830_, data_stage_5__6829_, data_stage_5__6828_, data_stage_5__6827_, data_stage_5__6826_, data_stage_5__6825_, data_stage_5__6824_, data_stage_5__6823_, data_stage_5__6822_, data_stage_5__6821_, data_stage_5__6820_, data_stage_5__6819_, data_stage_5__6818_, data_stage_5__6817_, data_stage_5__6816_, data_stage_5__6815_, data_stage_5__6814_, data_stage_5__6813_, data_stage_5__6812_, data_stage_5__6811_, data_stage_5__6810_, data_stage_5__6809_, data_stage_5__6808_, data_stage_5__6807_, data_stage_5__6806_, data_stage_5__6805_, data_stage_5__6804_, data_stage_5__6803_, data_stage_5__6802_, data_stage_5__6801_, data_stage_5__6800_, data_stage_5__6799_, data_stage_5__6798_, data_stage_5__6797_, data_stage_5__6796_, data_stage_5__6795_, data_stage_5__6794_, data_stage_5__6793_, data_stage_5__6792_, data_stage_5__6791_, data_stage_5__6790_, data_stage_5__6789_, data_stage_5__6788_, data_stage_5__6787_, data_stage_5__6786_, data_stage_5__6785_, data_stage_5__6784_, data_stage_5__6783_, data_stage_5__6782_, data_stage_5__6781_, data_stage_5__6780_, data_stage_5__6779_, data_stage_5__6778_, data_stage_5__6777_, data_stage_5__6776_, data_stage_5__6775_, data_stage_5__6774_, data_stage_5__6773_, data_stage_5__6772_, data_stage_5__6771_, data_stage_5__6770_, data_stage_5__6769_, data_stage_5__6768_, data_stage_5__6767_, data_stage_5__6766_, data_stage_5__6765_, data_stage_5__6764_, data_stage_5__6763_, data_stage_5__6762_, data_stage_5__6761_, data_stage_5__6760_, data_stage_5__6759_, data_stage_5__6758_, data_stage_5__6757_, data_stage_5__6756_, data_stage_5__6755_, data_stage_5__6754_, data_stage_5__6753_, data_stage_5__6752_, data_stage_5__6751_, data_stage_5__6750_, data_stage_5__6749_, data_stage_5__6748_, data_stage_5__6747_, data_stage_5__6746_, data_stage_5__6745_, data_stage_5__6744_, data_stage_5__6743_, data_stage_5__6742_, data_stage_5__6741_, data_stage_5__6740_, data_stage_5__6739_, data_stage_5__6738_, data_stage_5__6737_, data_stage_5__6736_, data_stage_5__6735_, data_stage_5__6734_, data_stage_5__6733_, data_stage_5__6732_, data_stage_5__6731_, data_stage_5__6730_, data_stage_5__6729_, data_stage_5__6728_, data_stage_5__6727_, data_stage_5__6726_, data_stage_5__6725_, data_stage_5__6724_, data_stage_5__6723_, data_stage_5__6722_, data_stage_5__6721_, data_stage_5__6720_, data_stage_5__6719_, data_stage_5__6718_, data_stage_5__6717_, data_stage_5__6716_, data_stage_5__6715_, data_stage_5__6714_, data_stage_5__6713_, data_stage_5__6712_, data_stage_5__6711_, data_stage_5__6710_, data_stage_5__6709_, data_stage_5__6708_, data_stage_5__6707_, data_stage_5__6706_, data_stage_5__6705_, data_stage_5__6704_, data_stage_5__6703_, data_stage_5__6702_, data_stage_5__6701_, data_stage_5__6700_, data_stage_5__6699_, data_stage_5__6698_, data_stage_5__6697_, data_stage_5__6696_, data_stage_5__6695_, data_stage_5__6694_, data_stage_5__6693_, data_stage_5__6692_, data_stage_5__6691_, data_stage_5__6690_, data_stage_5__6689_, data_stage_5__6688_, data_stage_5__6687_, data_stage_5__6686_, data_stage_5__6685_, data_stage_5__6684_, data_stage_5__6683_, data_stage_5__6682_, data_stage_5__6681_, data_stage_5__6680_, data_stage_5__6679_, data_stage_5__6678_, data_stage_5__6677_, data_stage_5__6676_, data_stage_5__6675_, data_stage_5__6674_, data_stage_5__6673_, data_stage_5__6672_, data_stage_5__6671_, data_stage_5__6670_, data_stage_5__6669_, data_stage_5__6668_, data_stage_5__6667_, data_stage_5__6666_, data_stage_5__6665_, data_stage_5__6664_, data_stage_5__6663_, data_stage_5__6662_, data_stage_5__6661_, data_stage_5__6660_, data_stage_5__6659_, data_stage_5__6658_, data_stage_5__6657_, data_stage_5__6656_, data_stage_5__6655_, data_stage_5__6654_, data_stage_5__6653_, data_stage_5__6652_, data_stage_5__6651_, data_stage_5__6650_, data_stage_5__6649_, data_stage_5__6648_, data_stage_5__6647_, data_stage_5__6646_, data_stage_5__6645_, data_stage_5__6644_, data_stage_5__6643_, data_stage_5__6642_, data_stage_5__6641_, data_stage_5__6640_, data_stage_5__6639_, data_stage_5__6638_, data_stage_5__6637_, data_stage_5__6636_, data_stage_5__6635_, data_stage_5__6634_, data_stage_5__6633_, data_stage_5__6632_, data_stage_5__6631_, data_stage_5__6630_, data_stage_5__6629_, data_stage_5__6628_, data_stage_5__6627_, data_stage_5__6626_, data_stage_5__6625_, data_stage_5__6624_, data_stage_5__6623_, data_stage_5__6622_, data_stage_5__6621_, data_stage_5__6620_, data_stage_5__6619_, data_stage_5__6618_, data_stage_5__6617_, data_stage_5__6616_, data_stage_5__6615_, data_stage_5__6614_, data_stage_5__6613_, data_stage_5__6612_, data_stage_5__6611_, data_stage_5__6610_, data_stage_5__6609_, data_stage_5__6608_, data_stage_5__6607_, data_stage_5__6606_, data_stage_5__6605_, data_stage_5__6604_, data_stage_5__6603_, data_stage_5__6602_, data_stage_5__6601_, data_stage_5__6600_, data_stage_5__6599_, data_stage_5__6598_, data_stage_5__6597_, data_stage_5__6596_, data_stage_5__6595_, data_stage_5__6594_, data_stage_5__6593_, data_stage_5__6592_, data_stage_5__6591_, data_stage_5__6590_, data_stage_5__6589_, data_stage_5__6588_, data_stage_5__6587_, data_stage_5__6586_, data_stage_5__6585_, data_stage_5__6584_, data_stage_5__6583_, data_stage_5__6582_, data_stage_5__6581_, data_stage_5__6580_, data_stage_5__6579_, data_stage_5__6578_, data_stage_5__6577_, data_stage_5__6576_, data_stage_5__6575_, data_stage_5__6574_, data_stage_5__6573_, data_stage_5__6572_, data_stage_5__6571_, data_stage_5__6570_, data_stage_5__6569_, data_stage_5__6568_, data_stage_5__6567_, data_stage_5__6566_, data_stage_5__6565_, data_stage_5__6564_, data_stage_5__6563_, data_stage_5__6562_, data_stage_5__6561_, data_stage_5__6560_, data_stage_5__6559_, data_stage_5__6558_, data_stage_5__6557_, data_stage_5__6556_, data_stage_5__6555_, data_stage_5__6554_, data_stage_5__6553_, data_stage_5__6552_, data_stage_5__6551_, data_stage_5__6550_, data_stage_5__6549_, data_stage_5__6548_, data_stage_5__6547_, data_stage_5__6546_, data_stage_5__6545_, data_stage_5__6544_, data_stage_5__6543_, data_stage_5__6542_, data_stage_5__6541_, data_stage_5__6540_, data_stage_5__6539_, data_stage_5__6538_, data_stage_5__6537_, data_stage_5__6536_, data_stage_5__6535_, data_stage_5__6534_, data_stage_5__6533_, data_stage_5__6532_, data_stage_5__6531_, data_stage_5__6530_, data_stage_5__6529_, data_stage_5__6528_, data_stage_5__6527_, data_stage_5__6526_, data_stage_5__6525_, data_stage_5__6524_, data_stage_5__6523_, data_stage_5__6522_, data_stage_5__6521_, data_stage_5__6520_, data_stage_5__6519_, data_stage_5__6518_, data_stage_5__6517_, data_stage_5__6516_, data_stage_5__6515_, data_stage_5__6514_, data_stage_5__6513_, data_stage_5__6512_, data_stage_5__6511_, data_stage_5__6510_, data_stage_5__6509_, data_stage_5__6508_, data_stage_5__6507_, data_stage_5__6506_, data_stage_5__6505_, data_stage_5__6504_, data_stage_5__6503_, data_stage_5__6502_, data_stage_5__6501_, data_stage_5__6500_, data_stage_5__6499_, data_stage_5__6498_, data_stage_5__6497_, data_stage_5__6496_, data_stage_5__6495_, data_stage_5__6494_, data_stage_5__6493_, data_stage_5__6492_, data_stage_5__6491_, data_stage_5__6490_, data_stage_5__6489_, data_stage_5__6488_, data_stage_5__6487_, data_stage_5__6486_, data_stage_5__6485_, data_stage_5__6484_, data_stage_5__6483_, data_stage_5__6482_, data_stage_5__6481_, data_stage_5__6480_, data_stage_5__6479_, data_stage_5__6478_, data_stage_5__6477_, data_stage_5__6476_, data_stage_5__6475_, data_stage_5__6474_, data_stage_5__6473_, data_stage_5__6472_, data_stage_5__6471_, data_stage_5__6470_, data_stage_5__6469_, data_stage_5__6468_, data_stage_5__6467_, data_stage_5__6466_, data_stage_5__6465_, data_stage_5__6464_, data_stage_5__6463_, data_stage_5__6462_, data_stage_5__6461_, data_stage_5__6460_, data_stage_5__6459_, data_stage_5__6458_, data_stage_5__6457_, data_stage_5__6456_, data_stage_5__6455_, data_stage_5__6454_, data_stage_5__6453_, data_stage_5__6452_, data_stage_5__6451_, data_stage_5__6450_, data_stage_5__6449_, data_stage_5__6448_, data_stage_5__6447_, data_stage_5__6446_, data_stage_5__6445_, data_stage_5__6444_, data_stage_5__6443_, data_stage_5__6442_, data_stage_5__6441_, data_stage_5__6440_, data_stage_5__6439_, data_stage_5__6438_, data_stage_5__6437_, data_stage_5__6436_, data_stage_5__6435_, data_stage_5__6434_, data_stage_5__6433_, data_stage_5__6432_, data_stage_5__6431_, data_stage_5__6430_, data_stage_5__6429_, data_stage_5__6428_, data_stage_5__6427_, data_stage_5__6426_, data_stage_5__6425_, data_stage_5__6424_, data_stage_5__6423_, data_stage_5__6422_, data_stage_5__6421_, data_stage_5__6420_, data_stage_5__6419_, data_stage_5__6418_, data_stage_5__6417_, data_stage_5__6416_, data_stage_5__6415_, data_stage_5__6414_, data_stage_5__6413_, data_stage_5__6412_, data_stage_5__6411_, data_stage_5__6410_, data_stage_5__6409_, data_stage_5__6408_, data_stage_5__6407_, data_stage_5__6406_, data_stage_5__6405_, data_stage_5__6404_, data_stage_5__6403_, data_stage_5__6402_, data_stage_5__6401_, data_stage_5__6400_, data_stage_5__6399_, data_stage_5__6398_, data_stage_5__6397_, data_stage_5__6396_, data_stage_5__6395_, data_stage_5__6394_, data_stage_5__6393_, data_stage_5__6392_, data_stage_5__6391_, data_stage_5__6390_, data_stage_5__6389_, data_stage_5__6388_, data_stage_5__6387_, data_stage_5__6386_, data_stage_5__6385_, data_stage_5__6384_, data_stage_5__6383_, data_stage_5__6382_, data_stage_5__6381_, data_stage_5__6380_, data_stage_5__6379_, data_stage_5__6378_, data_stage_5__6377_, data_stage_5__6376_, data_stage_5__6375_, data_stage_5__6374_, data_stage_5__6373_, data_stage_5__6372_, data_stage_5__6371_, data_stage_5__6370_, data_stage_5__6369_, data_stage_5__6368_, data_stage_5__6367_, data_stage_5__6366_, data_stage_5__6365_, data_stage_5__6364_, data_stage_5__6363_, data_stage_5__6362_, data_stage_5__6361_, data_stage_5__6360_, data_stage_5__6359_, data_stage_5__6358_, data_stage_5__6357_, data_stage_5__6356_, data_stage_5__6355_, data_stage_5__6354_, data_stage_5__6353_, data_stage_5__6352_, data_stage_5__6351_, data_stage_5__6350_, data_stage_5__6349_, data_stage_5__6348_, data_stage_5__6347_, data_stage_5__6346_, data_stage_5__6345_, data_stage_5__6344_, data_stage_5__6343_, data_stage_5__6342_, data_stage_5__6341_, data_stage_5__6340_, data_stage_5__6339_, data_stage_5__6338_, data_stage_5__6337_, data_stage_5__6336_, data_stage_5__6335_, data_stage_5__6334_, data_stage_5__6333_, data_stage_5__6332_, data_stage_5__6331_, data_stage_5__6330_, data_stage_5__6329_, data_stage_5__6328_, data_stage_5__6327_, data_stage_5__6326_, data_stage_5__6325_, data_stage_5__6324_, data_stage_5__6323_, data_stage_5__6322_, data_stage_5__6321_, data_stage_5__6320_, data_stage_5__6319_, data_stage_5__6318_, data_stage_5__6317_, data_stage_5__6316_, data_stage_5__6315_, data_stage_5__6314_, data_stage_5__6313_, data_stage_5__6312_, data_stage_5__6311_, data_stage_5__6310_, data_stage_5__6309_, data_stage_5__6308_, data_stage_5__6307_, data_stage_5__6306_, data_stage_5__6305_, data_stage_5__6304_, data_stage_5__6303_, data_stage_5__6302_, data_stage_5__6301_, data_stage_5__6300_, data_stage_5__6299_, data_stage_5__6298_, data_stage_5__6297_, data_stage_5__6296_, data_stage_5__6295_, data_stage_5__6294_, data_stage_5__6293_, data_stage_5__6292_, data_stage_5__6291_, data_stage_5__6290_, data_stage_5__6289_, data_stage_5__6288_, data_stage_5__6287_, data_stage_5__6286_, data_stage_5__6285_, data_stage_5__6284_, data_stage_5__6283_, data_stage_5__6282_, data_stage_5__6281_, data_stage_5__6280_, data_stage_5__6279_, data_stage_5__6278_, data_stage_5__6277_, data_stage_5__6276_, data_stage_5__6275_, data_stage_5__6274_, data_stage_5__6273_, data_stage_5__6272_, data_stage_5__6271_, data_stage_5__6270_, data_stage_5__6269_, data_stage_5__6268_, data_stage_5__6267_, data_stage_5__6266_, data_stage_5__6265_, data_stage_5__6264_, data_stage_5__6263_, data_stage_5__6262_, data_stage_5__6261_, data_stage_5__6260_, data_stage_5__6259_, data_stage_5__6258_, data_stage_5__6257_, data_stage_5__6256_, data_stage_5__6255_, data_stage_5__6254_, data_stage_5__6253_, data_stage_5__6252_, data_stage_5__6251_, data_stage_5__6250_, data_stage_5__6249_, data_stage_5__6248_, data_stage_5__6247_, data_stage_5__6246_, data_stage_5__6245_, data_stage_5__6244_, data_stage_5__6243_, data_stage_5__6242_, data_stage_5__6241_, data_stage_5__6240_, data_stage_5__6239_, data_stage_5__6238_, data_stage_5__6237_, data_stage_5__6236_, data_stage_5__6235_, data_stage_5__6234_, data_stage_5__6233_, data_stage_5__6232_, data_stage_5__6231_, data_stage_5__6230_, data_stage_5__6229_, data_stage_5__6228_, data_stage_5__6227_, data_stage_5__6226_, data_stage_5__6225_, data_stage_5__6224_, data_stage_5__6223_, data_stage_5__6222_, data_stage_5__6221_, data_stage_5__6220_, data_stage_5__6219_, data_stage_5__6218_, data_stage_5__6217_, data_stage_5__6216_, data_stage_5__6215_, data_stage_5__6214_, data_stage_5__6213_, data_stage_5__6212_, data_stage_5__6211_, data_stage_5__6210_, data_stage_5__6209_, data_stage_5__6208_, data_stage_5__6207_, data_stage_5__6206_, data_stage_5__6205_, data_stage_5__6204_, data_stage_5__6203_, data_stage_5__6202_, data_stage_5__6201_, data_stage_5__6200_, data_stage_5__6199_, data_stage_5__6198_, data_stage_5__6197_, data_stage_5__6196_, data_stage_5__6195_, data_stage_5__6194_, data_stage_5__6193_, data_stage_5__6192_, data_stage_5__6191_, data_stage_5__6190_, data_stage_5__6189_, data_stage_5__6188_, data_stage_5__6187_, data_stage_5__6186_, data_stage_5__6185_, data_stage_5__6184_, data_stage_5__6183_, data_stage_5__6182_, data_stage_5__6181_, data_stage_5__6180_, data_stage_5__6179_, data_stage_5__6178_, data_stage_5__6177_, data_stage_5__6176_, data_stage_5__6175_, data_stage_5__6174_, data_stage_5__6173_, data_stage_5__6172_, data_stage_5__6171_, data_stage_5__6170_, data_stage_5__6169_, data_stage_5__6168_, data_stage_5__6167_, data_stage_5__6166_, data_stage_5__6165_, data_stage_5__6164_, data_stage_5__6163_, data_stage_5__6162_, data_stage_5__6161_, data_stage_5__6160_, data_stage_5__6159_, data_stage_5__6158_, data_stage_5__6157_, data_stage_5__6156_, data_stage_5__6155_, data_stage_5__6154_, data_stage_5__6153_, data_stage_5__6152_, data_stage_5__6151_, data_stage_5__6150_, data_stage_5__6149_, data_stage_5__6148_, data_stage_5__6147_, data_stage_5__6146_, data_stage_5__6145_, data_stage_5__6144_, data_stage_5__6143_, data_stage_5__6142_, data_stage_5__6141_, data_stage_5__6140_, data_stage_5__6139_, data_stage_5__6138_, data_stage_5__6137_, data_stage_5__6136_, data_stage_5__6135_, data_stage_5__6134_, data_stage_5__6133_, data_stage_5__6132_, data_stage_5__6131_, data_stage_5__6130_, data_stage_5__6129_, data_stage_5__6128_, data_stage_5__6127_, data_stage_5__6126_, data_stage_5__6125_, data_stage_5__6124_, data_stage_5__6123_, data_stage_5__6122_, data_stage_5__6121_, data_stage_5__6120_, data_stage_5__6119_, data_stage_5__6118_, data_stage_5__6117_, data_stage_5__6116_, data_stage_5__6115_, data_stage_5__6114_, data_stage_5__6113_, data_stage_5__6112_, data_stage_5__6111_, data_stage_5__6110_, data_stage_5__6109_, data_stage_5__6108_, data_stage_5__6107_, data_stage_5__6106_, data_stage_5__6105_, data_stage_5__6104_, data_stage_5__6103_, data_stage_5__6102_, data_stage_5__6101_, data_stage_5__6100_, data_stage_5__6099_, data_stage_5__6098_, data_stage_5__6097_, data_stage_5__6096_, data_stage_5__6095_, data_stage_5__6094_, data_stage_5__6093_, data_stage_5__6092_, data_stage_5__6091_, data_stage_5__6090_, data_stage_5__6089_, data_stage_5__6088_, data_stage_5__6087_, data_stage_5__6086_, data_stage_5__6085_, data_stage_5__6084_, data_stage_5__6083_, data_stage_5__6082_, data_stage_5__6081_, data_stage_5__6080_, data_stage_5__6079_, data_stage_5__6078_, data_stage_5__6077_, data_stage_5__6076_, data_stage_5__6075_, data_stage_5__6074_, data_stage_5__6073_, data_stage_5__6072_, data_stage_5__6071_, data_stage_5__6070_, data_stage_5__6069_, data_stage_5__6068_, data_stage_5__6067_, data_stage_5__6066_, data_stage_5__6065_, data_stage_5__6064_, data_stage_5__6063_, data_stage_5__6062_, data_stage_5__6061_, data_stage_5__6060_, data_stage_5__6059_, data_stage_5__6058_, data_stage_5__6057_, data_stage_5__6056_, data_stage_5__6055_, data_stage_5__6054_, data_stage_5__6053_, data_stage_5__6052_, data_stage_5__6051_, data_stage_5__6050_, data_stage_5__6049_, data_stage_5__6048_, data_stage_5__6047_, data_stage_5__6046_, data_stage_5__6045_, data_stage_5__6044_, data_stage_5__6043_, data_stage_5__6042_, data_stage_5__6041_, data_stage_5__6040_, data_stage_5__6039_, data_stage_5__6038_, data_stage_5__6037_, data_stage_5__6036_, data_stage_5__6035_, data_stage_5__6034_, data_stage_5__6033_, data_stage_5__6032_, data_stage_5__6031_, data_stage_5__6030_, data_stage_5__6029_, data_stage_5__6028_, data_stage_5__6027_, data_stage_5__6026_, data_stage_5__6025_, data_stage_5__6024_, data_stage_5__6023_, data_stage_5__6022_, data_stage_5__6021_, data_stage_5__6020_, data_stage_5__6019_, data_stage_5__6018_, data_stage_5__6017_, data_stage_5__6016_, data_stage_5__6015_, data_stage_5__6014_, data_stage_5__6013_, data_stage_5__6012_, data_stage_5__6011_, data_stage_5__6010_, data_stage_5__6009_, data_stage_5__6008_, data_stage_5__6007_, data_stage_5__6006_, data_stage_5__6005_, data_stage_5__6004_, data_stage_5__6003_, data_stage_5__6002_, data_stage_5__6001_, data_stage_5__6000_, data_stage_5__5999_, data_stage_5__5998_, data_stage_5__5997_, data_stage_5__5996_, data_stage_5__5995_, data_stage_5__5994_, data_stage_5__5993_, data_stage_5__5992_, data_stage_5__5991_, data_stage_5__5990_, data_stage_5__5989_, data_stage_5__5988_, data_stage_5__5987_, data_stage_5__5986_, data_stage_5__5985_, data_stage_5__5984_, data_stage_5__5983_, data_stage_5__5982_, data_stage_5__5981_, data_stage_5__5980_, data_stage_5__5979_, data_stage_5__5978_, data_stage_5__5977_, data_stage_5__5976_, data_stage_5__5975_, data_stage_5__5974_, data_stage_5__5973_, data_stage_5__5972_, data_stage_5__5971_, data_stage_5__5970_, data_stage_5__5969_, data_stage_5__5968_, data_stage_5__5967_, data_stage_5__5966_, data_stage_5__5965_, data_stage_5__5964_, data_stage_5__5963_, data_stage_5__5962_, data_stage_5__5961_, data_stage_5__5960_, data_stage_5__5959_, data_stage_5__5958_, data_stage_5__5957_, data_stage_5__5956_, data_stage_5__5955_, data_stage_5__5954_, data_stage_5__5953_, data_stage_5__5952_, data_stage_5__5951_, data_stage_5__5950_, data_stage_5__5949_, data_stage_5__5948_, data_stage_5__5947_, data_stage_5__5946_, data_stage_5__5945_, data_stage_5__5944_, data_stage_5__5943_, data_stage_5__5942_, data_stage_5__5941_, data_stage_5__5940_, data_stage_5__5939_, data_stage_5__5938_, data_stage_5__5937_, data_stage_5__5936_, data_stage_5__5935_, data_stage_5__5934_, data_stage_5__5933_, data_stage_5__5932_, data_stage_5__5931_, data_stage_5__5930_, data_stage_5__5929_, data_stage_5__5928_, data_stage_5__5927_, data_stage_5__5926_, data_stage_5__5925_, data_stage_5__5924_, data_stage_5__5923_, data_stage_5__5922_, data_stage_5__5921_, data_stage_5__5920_, data_stage_5__5919_, data_stage_5__5918_, data_stage_5__5917_, data_stage_5__5916_, data_stage_5__5915_, data_stage_5__5914_, data_stage_5__5913_, data_stage_5__5912_, data_stage_5__5911_, data_stage_5__5910_, data_stage_5__5909_, data_stage_5__5908_, data_stage_5__5907_, data_stage_5__5906_, data_stage_5__5905_, data_stage_5__5904_, data_stage_5__5903_, data_stage_5__5902_, data_stage_5__5901_, data_stage_5__5900_, data_stage_5__5899_, data_stage_5__5898_, data_stage_5__5897_, data_stage_5__5896_, data_stage_5__5895_, data_stage_5__5894_, data_stage_5__5893_, data_stage_5__5892_, data_stage_5__5891_, data_stage_5__5890_, data_stage_5__5889_, data_stage_5__5888_, data_stage_5__5887_, data_stage_5__5886_, data_stage_5__5885_, data_stage_5__5884_, data_stage_5__5883_, data_stage_5__5882_, data_stage_5__5881_, data_stage_5__5880_, data_stage_5__5879_, data_stage_5__5878_, data_stage_5__5877_, data_stage_5__5876_, data_stage_5__5875_, data_stage_5__5874_, data_stage_5__5873_, data_stage_5__5872_, data_stage_5__5871_, data_stage_5__5870_, data_stage_5__5869_, data_stage_5__5868_, data_stage_5__5867_, data_stage_5__5866_, data_stage_5__5865_, data_stage_5__5864_, data_stage_5__5863_, data_stage_5__5862_, data_stage_5__5861_, data_stage_5__5860_, data_stage_5__5859_, data_stage_5__5858_, data_stage_5__5857_, data_stage_5__5856_, data_stage_5__5855_, data_stage_5__5854_, data_stage_5__5853_, data_stage_5__5852_, data_stage_5__5851_, data_stage_5__5850_, data_stage_5__5849_, data_stage_5__5848_, data_stage_5__5847_, data_stage_5__5846_, data_stage_5__5845_, data_stage_5__5844_, data_stage_5__5843_, data_stage_5__5842_, data_stage_5__5841_, data_stage_5__5840_, data_stage_5__5839_, data_stage_5__5838_, data_stage_5__5837_, data_stage_5__5836_, data_stage_5__5835_, data_stage_5__5834_, data_stage_5__5833_, data_stage_5__5832_, data_stage_5__5831_, data_stage_5__5830_, data_stage_5__5829_, data_stage_5__5828_, data_stage_5__5827_, data_stage_5__5826_, data_stage_5__5825_, data_stage_5__5824_, data_stage_5__5823_, data_stage_5__5822_, data_stage_5__5821_, data_stage_5__5820_, data_stage_5__5819_, data_stage_5__5818_, data_stage_5__5817_, data_stage_5__5816_, data_stage_5__5815_, data_stage_5__5814_, data_stage_5__5813_, data_stage_5__5812_, data_stage_5__5811_, data_stage_5__5810_, data_stage_5__5809_, data_stage_5__5808_, data_stage_5__5807_, data_stage_5__5806_, data_stage_5__5805_, data_stage_5__5804_, data_stage_5__5803_, data_stage_5__5802_, data_stage_5__5801_, data_stage_5__5800_, data_stage_5__5799_, data_stage_5__5798_, data_stage_5__5797_, data_stage_5__5796_, data_stage_5__5795_, data_stage_5__5794_, data_stage_5__5793_, data_stage_5__5792_, data_stage_5__5791_, data_stage_5__5790_, data_stage_5__5789_, data_stage_5__5788_, data_stage_5__5787_, data_stage_5__5786_, data_stage_5__5785_, data_stage_5__5784_, data_stage_5__5783_, data_stage_5__5782_, data_stage_5__5781_, data_stage_5__5780_, data_stage_5__5779_, data_stage_5__5778_, data_stage_5__5777_, data_stage_5__5776_, data_stage_5__5775_, data_stage_5__5774_, data_stage_5__5773_, data_stage_5__5772_, data_stage_5__5771_, data_stage_5__5770_, data_stage_5__5769_, data_stage_5__5768_, data_stage_5__5767_, data_stage_5__5766_, data_stage_5__5765_, data_stage_5__5764_, data_stage_5__5763_, data_stage_5__5762_, data_stage_5__5761_, data_stage_5__5760_, data_stage_5__5759_, data_stage_5__5758_, data_stage_5__5757_, data_stage_5__5756_, data_stage_5__5755_, data_stage_5__5754_, data_stage_5__5753_, data_stage_5__5752_, data_stage_5__5751_, data_stage_5__5750_, data_stage_5__5749_, data_stage_5__5748_, data_stage_5__5747_, data_stage_5__5746_, data_stage_5__5745_, data_stage_5__5744_, data_stage_5__5743_, data_stage_5__5742_, data_stage_5__5741_, data_stage_5__5740_, data_stage_5__5739_, data_stage_5__5738_, data_stage_5__5737_, data_stage_5__5736_, data_stage_5__5735_, data_stage_5__5734_, data_stage_5__5733_, data_stage_5__5732_, data_stage_5__5731_, data_stage_5__5730_, data_stage_5__5729_, data_stage_5__5728_, data_stage_5__5727_, data_stage_5__5726_, data_stage_5__5725_, data_stage_5__5724_, data_stage_5__5723_, data_stage_5__5722_, data_stage_5__5721_, data_stage_5__5720_, data_stage_5__5719_, data_stage_5__5718_, data_stage_5__5717_, data_stage_5__5716_, data_stage_5__5715_, data_stage_5__5714_, data_stage_5__5713_, data_stage_5__5712_, data_stage_5__5711_, data_stage_5__5710_, data_stage_5__5709_, data_stage_5__5708_, data_stage_5__5707_, data_stage_5__5706_, data_stage_5__5705_, data_stage_5__5704_, data_stage_5__5703_, data_stage_5__5702_, data_stage_5__5701_, data_stage_5__5700_, data_stage_5__5699_, data_stage_5__5698_, data_stage_5__5697_, data_stage_5__5696_, data_stage_5__5695_, data_stage_5__5694_, data_stage_5__5693_, data_stage_5__5692_, data_stage_5__5691_, data_stage_5__5690_, data_stage_5__5689_, data_stage_5__5688_, data_stage_5__5687_, data_stage_5__5686_, data_stage_5__5685_, data_stage_5__5684_, data_stage_5__5683_, data_stage_5__5682_, data_stage_5__5681_, data_stage_5__5680_, data_stage_5__5679_, data_stage_5__5678_, data_stage_5__5677_, data_stage_5__5676_, data_stage_5__5675_, data_stage_5__5674_, data_stage_5__5673_, data_stage_5__5672_, data_stage_5__5671_, data_stage_5__5670_, data_stage_5__5669_, data_stage_5__5668_, data_stage_5__5667_, data_stage_5__5666_, data_stage_5__5665_, data_stage_5__5664_, data_stage_5__5663_, data_stage_5__5662_, data_stage_5__5661_, data_stage_5__5660_, data_stage_5__5659_, data_stage_5__5658_, data_stage_5__5657_, data_stage_5__5656_, data_stage_5__5655_, data_stage_5__5654_, data_stage_5__5653_, data_stage_5__5652_, data_stage_5__5651_, data_stage_5__5650_, data_stage_5__5649_, data_stage_5__5648_, data_stage_5__5647_, data_stage_5__5646_, data_stage_5__5645_, data_stage_5__5644_, data_stage_5__5643_, data_stage_5__5642_, data_stage_5__5641_, data_stage_5__5640_, data_stage_5__5639_, data_stage_5__5638_, data_stage_5__5637_, data_stage_5__5636_, data_stage_5__5635_, data_stage_5__5634_, data_stage_5__5633_, data_stage_5__5632_, data_stage_5__5631_, data_stage_5__5630_, data_stage_5__5629_, data_stage_5__5628_, data_stage_5__5627_, data_stage_5__5626_, data_stage_5__5625_, data_stage_5__5624_, data_stage_5__5623_, data_stage_5__5622_, data_stage_5__5621_, data_stage_5__5620_, data_stage_5__5619_, data_stage_5__5618_, data_stage_5__5617_, data_stage_5__5616_, data_stage_5__5615_, data_stage_5__5614_, data_stage_5__5613_, data_stage_5__5612_, data_stage_5__5611_, data_stage_5__5610_, data_stage_5__5609_, data_stage_5__5608_, data_stage_5__5607_, data_stage_5__5606_, data_stage_5__5605_, data_stage_5__5604_, data_stage_5__5603_, data_stage_5__5602_, data_stage_5__5601_, data_stage_5__5600_, data_stage_5__5599_, data_stage_5__5598_, data_stage_5__5597_, data_stage_5__5596_, data_stage_5__5595_, data_stage_5__5594_, data_stage_5__5593_, data_stage_5__5592_, data_stage_5__5591_, data_stage_5__5590_, data_stage_5__5589_, data_stage_5__5588_, data_stage_5__5587_, data_stage_5__5586_, data_stage_5__5585_, data_stage_5__5584_, data_stage_5__5583_, data_stage_5__5582_, data_stage_5__5581_, data_stage_5__5580_, data_stage_5__5579_, data_stage_5__5578_, data_stage_5__5577_, data_stage_5__5576_, data_stage_5__5575_, data_stage_5__5574_, data_stage_5__5573_, data_stage_5__5572_, data_stage_5__5571_, data_stage_5__5570_, data_stage_5__5569_, data_stage_5__5568_, data_stage_5__5567_, data_stage_5__5566_, data_stage_5__5565_, data_stage_5__5564_, data_stage_5__5563_, data_stage_5__5562_, data_stage_5__5561_, data_stage_5__5560_, data_stage_5__5559_, data_stage_5__5558_, data_stage_5__5557_, data_stage_5__5556_, data_stage_5__5555_, data_stage_5__5554_, data_stage_5__5553_, data_stage_5__5552_, data_stage_5__5551_, data_stage_5__5550_, data_stage_5__5549_, data_stage_5__5548_, data_stage_5__5547_, data_stage_5__5546_, data_stage_5__5545_, data_stage_5__5544_, data_stage_5__5543_, data_stage_5__5542_, data_stage_5__5541_, data_stage_5__5540_, data_stage_5__5539_, data_stage_5__5538_, data_stage_5__5537_, data_stage_5__5536_, data_stage_5__5535_, data_stage_5__5534_, data_stage_5__5533_, data_stage_5__5532_, data_stage_5__5531_, data_stage_5__5530_, data_stage_5__5529_, data_stage_5__5528_, data_stage_5__5527_, data_stage_5__5526_, data_stage_5__5525_, data_stage_5__5524_, data_stage_5__5523_, data_stage_5__5522_, data_stage_5__5521_, data_stage_5__5520_, data_stage_5__5519_, data_stage_5__5518_, data_stage_5__5517_, data_stage_5__5516_, data_stage_5__5515_, data_stage_5__5514_, data_stage_5__5513_, data_stage_5__5512_, data_stage_5__5511_, data_stage_5__5510_, data_stage_5__5509_, data_stage_5__5508_, data_stage_5__5507_, data_stage_5__5506_, data_stage_5__5505_, data_stage_5__5504_, data_stage_5__5503_, data_stage_5__5502_, data_stage_5__5501_, data_stage_5__5500_, data_stage_5__5499_, data_stage_5__5498_, data_stage_5__5497_, data_stage_5__5496_, data_stage_5__5495_, data_stage_5__5494_, data_stage_5__5493_, data_stage_5__5492_, data_stage_5__5491_, data_stage_5__5490_, data_stage_5__5489_, data_stage_5__5488_, data_stage_5__5487_, data_stage_5__5486_, data_stage_5__5485_, data_stage_5__5484_, data_stage_5__5483_, data_stage_5__5482_, data_stage_5__5481_, data_stage_5__5480_, data_stage_5__5479_, data_stage_5__5478_, data_stage_5__5477_, data_stage_5__5476_, data_stage_5__5475_, data_stage_5__5474_, data_stage_5__5473_, data_stage_5__5472_, data_stage_5__5471_, data_stage_5__5470_, data_stage_5__5469_, data_stage_5__5468_, data_stage_5__5467_, data_stage_5__5466_, data_stage_5__5465_, data_stage_5__5464_, data_stage_5__5463_, data_stage_5__5462_, data_stage_5__5461_, data_stage_5__5460_, data_stage_5__5459_, data_stage_5__5458_, data_stage_5__5457_, data_stage_5__5456_, data_stage_5__5455_, data_stage_5__5454_, data_stage_5__5453_, data_stage_5__5452_, data_stage_5__5451_, data_stage_5__5450_, data_stage_5__5449_, data_stage_5__5448_, data_stage_5__5447_, data_stage_5__5446_, data_stage_5__5445_, data_stage_5__5444_, data_stage_5__5443_, data_stage_5__5442_, data_stage_5__5441_, data_stage_5__5440_, data_stage_5__5439_, data_stage_5__5438_, data_stage_5__5437_, data_stage_5__5436_, data_stage_5__5435_, data_stage_5__5434_, data_stage_5__5433_, data_stage_5__5432_, data_stage_5__5431_, data_stage_5__5430_, data_stage_5__5429_, data_stage_5__5428_, data_stage_5__5427_, data_stage_5__5426_, data_stage_5__5425_, data_stage_5__5424_, data_stage_5__5423_, data_stage_5__5422_, data_stage_5__5421_, data_stage_5__5420_, data_stage_5__5419_, data_stage_5__5418_, data_stage_5__5417_, data_stage_5__5416_, data_stage_5__5415_, data_stage_5__5414_, data_stage_5__5413_, data_stage_5__5412_, data_stage_5__5411_, data_stage_5__5410_, data_stage_5__5409_, data_stage_5__5408_, data_stage_5__5407_, data_stage_5__5406_, data_stage_5__5405_, data_stage_5__5404_, data_stage_5__5403_, data_stage_5__5402_, data_stage_5__5401_, data_stage_5__5400_, data_stage_5__5399_, data_stage_5__5398_, data_stage_5__5397_, data_stage_5__5396_, data_stage_5__5395_, data_stage_5__5394_, data_stage_5__5393_, data_stage_5__5392_, data_stage_5__5391_, data_stage_5__5390_, data_stage_5__5389_, data_stage_5__5388_, data_stage_5__5387_, data_stage_5__5386_, data_stage_5__5385_, data_stage_5__5384_, data_stage_5__5383_, data_stage_5__5382_, data_stage_5__5381_, data_stage_5__5380_, data_stage_5__5379_, data_stage_5__5378_, data_stage_5__5377_, data_stage_5__5376_, data_stage_5__5375_, data_stage_5__5374_, data_stage_5__5373_, data_stage_5__5372_, data_stage_5__5371_, data_stage_5__5370_, data_stage_5__5369_, data_stage_5__5368_, data_stage_5__5367_, data_stage_5__5366_, data_stage_5__5365_, data_stage_5__5364_, data_stage_5__5363_, data_stage_5__5362_, data_stage_5__5361_, data_stage_5__5360_, data_stage_5__5359_, data_stage_5__5358_, data_stage_5__5357_, data_stage_5__5356_, data_stage_5__5355_, data_stage_5__5354_, data_stage_5__5353_, data_stage_5__5352_, data_stage_5__5351_, data_stage_5__5350_, data_stage_5__5349_, data_stage_5__5348_, data_stage_5__5347_, data_stage_5__5346_, data_stage_5__5345_, data_stage_5__5344_, data_stage_5__5343_, data_stage_5__5342_, data_stage_5__5341_, data_stage_5__5340_, data_stage_5__5339_, data_stage_5__5338_, data_stage_5__5337_, data_stage_5__5336_, data_stage_5__5335_, data_stage_5__5334_, data_stage_5__5333_, data_stage_5__5332_, data_stage_5__5331_, data_stage_5__5330_, data_stage_5__5329_, data_stage_5__5328_, data_stage_5__5327_, data_stage_5__5326_, data_stage_5__5325_, data_stage_5__5324_, data_stage_5__5323_, data_stage_5__5322_, data_stage_5__5321_, data_stage_5__5320_, data_stage_5__5319_, data_stage_5__5318_, data_stage_5__5317_, data_stage_5__5316_, data_stage_5__5315_, data_stage_5__5314_, data_stage_5__5313_, data_stage_5__5312_, data_stage_5__5311_, data_stage_5__5310_, data_stage_5__5309_, data_stage_5__5308_, data_stage_5__5307_, data_stage_5__5306_, data_stage_5__5305_, data_stage_5__5304_, data_stage_5__5303_, data_stage_5__5302_, data_stage_5__5301_, data_stage_5__5300_, data_stage_5__5299_, data_stage_5__5298_, data_stage_5__5297_, data_stage_5__5296_, data_stage_5__5295_, data_stage_5__5294_, data_stage_5__5293_, data_stage_5__5292_, data_stage_5__5291_, data_stage_5__5290_, data_stage_5__5289_, data_stage_5__5288_, data_stage_5__5287_, data_stage_5__5286_, data_stage_5__5285_, data_stage_5__5284_, data_stage_5__5283_, data_stage_5__5282_, data_stage_5__5281_, data_stage_5__5280_, data_stage_5__5279_, data_stage_5__5278_, data_stage_5__5277_, data_stage_5__5276_, data_stage_5__5275_, data_stage_5__5274_, data_stage_5__5273_, data_stage_5__5272_, data_stage_5__5271_, data_stage_5__5270_, data_stage_5__5269_, data_stage_5__5268_, data_stage_5__5267_, data_stage_5__5266_, data_stage_5__5265_, data_stage_5__5264_, data_stage_5__5263_, data_stage_5__5262_, data_stage_5__5261_, data_stage_5__5260_, data_stage_5__5259_, data_stage_5__5258_, data_stage_5__5257_, data_stage_5__5256_, data_stage_5__5255_, data_stage_5__5254_, data_stage_5__5253_, data_stage_5__5252_, data_stage_5__5251_, data_stage_5__5250_, data_stage_5__5249_, data_stage_5__5248_, data_stage_5__5247_, data_stage_5__5246_, data_stage_5__5245_, data_stage_5__5244_, data_stage_5__5243_, data_stage_5__5242_, data_stage_5__5241_, data_stage_5__5240_, data_stage_5__5239_, data_stage_5__5238_, data_stage_5__5237_, data_stage_5__5236_, data_stage_5__5235_, data_stage_5__5234_, data_stage_5__5233_, data_stage_5__5232_, data_stage_5__5231_, data_stage_5__5230_, data_stage_5__5229_, data_stage_5__5228_, data_stage_5__5227_, data_stage_5__5226_, data_stage_5__5225_, data_stage_5__5224_, data_stage_5__5223_, data_stage_5__5222_, data_stage_5__5221_, data_stage_5__5220_, data_stage_5__5219_, data_stage_5__5218_, data_stage_5__5217_, data_stage_5__5216_, data_stage_5__5215_, data_stage_5__5214_, data_stage_5__5213_, data_stage_5__5212_, data_stage_5__5211_, data_stage_5__5210_, data_stage_5__5209_, data_stage_5__5208_, data_stage_5__5207_, data_stage_5__5206_, data_stage_5__5205_, data_stage_5__5204_, data_stage_5__5203_, data_stage_5__5202_, data_stage_5__5201_, data_stage_5__5200_, data_stage_5__5199_, data_stage_5__5198_, data_stage_5__5197_, data_stage_5__5196_, data_stage_5__5195_, data_stage_5__5194_, data_stage_5__5193_, data_stage_5__5192_, data_stage_5__5191_, data_stage_5__5190_, data_stage_5__5189_, data_stage_5__5188_, data_stage_5__5187_, data_stage_5__5186_, data_stage_5__5185_, data_stage_5__5184_, data_stage_5__5183_, data_stage_5__5182_, data_stage_5__5181_, data_stage_5__5180_, data_stage_5__5179_, data_stage_5__5178_, data_stage_5__5177_, data_stage_5__5176_, data_stage_5__5175_, data_stage_5__5174_, data_stage_5__5173_, data_stage_5__5172_, data_stage_5__5171_, data_stage_5__5170_, data_stage_5__5169_, data_stage_5__5168_, data_stage_5__5167_, data_stage_5__5166_, data_stage_5__5165_, data_stage_5__5164_, data_stage_5__5163_, data_stage_5__5162_, data_stage_5__5161_, data_stage_5__5160_, data_stage_5__5159_, data_stage_5__5158_, data_stage_5__5157_, data_stage_5__5156_, data_stage_5__5155_, data_stage_5__5154_, data_stage_5__5153_, data_stage_5__5152_, data_stage_5__5151_, data_stage_5__5150_, data_stage_5__5149_, data_stage_5__5148_, data_stage_5__5147_, data_stage_5__5146_, data_stage_5__5145_, data_stage_5__5144_, data_stage_5__5143_, data_stage_5__5142_, data_stage_5__5141_, data_stage_5__5140_, data_stage_5__5139_, data_stage_5__5138_, data_stage_5__5137_, data_stage_5__5136_, data_stage_5__5135_, data_stage_5__5134_, data_stage_5__5133_, data_stage_5__5132_, data_stage_5__5131_, data_stage_5__5130_, data_stage_5__5129_, data_stage_5__5128_, data_stage_5__5127_, data_stage_5__5126_, data_stage_5__5125_, data_stage_5__5124_, data_stage_5__5123_, data_stage_5__5122_, data_stage_5__5121_, data_stage_5__5120_, data_stage_5__5119_, data_stage_5__5118_, data_stage_5__5117_, data_stage_5__5116_, data_stage_5__5115_, data_stage_5__5114_, data_stage_5__5113_, data_stage_5__5112_, data_stage_5__5111_, data_stage_5__5110_, data_stage_5__5109_, data_stage_5__5108_, data_stage_5__5107_, data_stage_5__5106_, data_stage_5__5105_, data_stage_5__5104_, data_stage_5__5103_, data_stage_5__5102_, data_stage_5__5101_, data_stage_5__5100_, data_stage_5__5099_, data_stage_5__5098_, data_stage_5__5097_, data_stage_5__5096_, data_stage_5__5095_, data_stage_5__5094_, data_stage_5__5093_, data_stage_5__5092_, data_stage_5__5091_, data_stage_5__5090_, data_stage_5__5089_, data_stage_5__5088_, data_stage_5__5087_, data_stage_5__5086_, data_stage_5__5085_, data_stage_5__5084_, data_stage_5__5083_, data_stage_5__5082_, data_stage_5__5081_, data_stage_5__5080_, data_stage_5__5079_, data_stage_5__5078_, data_stage_5__5077_, data_stage_5__5076_, data_stage_5__5075_, data_stage_5__5074_, data_stage_5__5073_, data_stage_5__5072_, data_stage_5__5071_, data_stage_5__5070_, data_stage_5__5069_, data_stage_5__5068_, data_stage_5__5067_, data_stage_5__5066_, data_stage_5__5065_, data_stage_5__5064_, data_stage_5__5063_, data_stage_5__5062_, data_stage_5__5061_, data_stage_5__5060_, data_stage_5__5059_, data_stage_5__5058_, data_stage_5__5057_, data_stage_5__5056_, data_stage_5__5055_, data_stage_5__5054_, data_stage_5__5053_, data_stage_5__5052_, data_stage_5__5051_, data_stage_5__5050_, data_stage_5__5049_, data_stage_5__5048_, data_stage_5__5047_, data_stage_5__5046_, data_stage_5__5045_, data_stage_5__5044_, data_stage_5__5043_, data_stage_5__5042_, data_stage_5__5041_, data_stage_5__5040_, data_stage_5__5039_, data_stage_5__5038_, data_stage_5__5037_, data_stage_5__5036_, data_stage_5__5035_, data_stage_5__5034_, data_stage_5__5033_, data_stage_5__5032_, data_stage_5__5031_, data_stage_5__5030_, data_stage_5__5029_, data_stage_5__5028_, data_stage_5__5027_, data_stage_5__5026_, data_stage_5__5025_, data_stage_5__5024_, data_stage_5__5023_, data_stage_5__5022_, data_stage_5__5021_, data_stage_5__5020_, data_stage_5__5019_, data_stage_5__5018_, data_stage_5__5017_, data_stage_5__5016_, data_stage_5__5015_, data_stage_5__5014_, data_stage_5__5013_, data_stage_5__5012_, data_stage_5__5011_, data_stage_5__5010_, data_stage_5__5009_, data_stage_5__5008_, data_stage_5__5007_, data_stage_5__5006_, data_stage_5__5005_, data_stage_5__5004_, data_stage_5__5003_, data_stage_5__5002_, data_stage_5__5001_, data_stage_5__5000_, data_stage_5__4999_, data_stage_5__4998_, data_stage_5__4997_, data_stage_5__4996_, data_stage_5__4995_, data_stage_5__4994_, data_stage_5__4993_, data_stage_5__4992_, data_stage_5__4991_, data_stage_5__4990_, data_stage_5__4989_, data_stage_5__4988_, data_stage_5__4987_, data_stage_5__4986_, data_stage_5__4985_, data_stage_5__4984_, data_stage_5__4983_, data_stage_5__4982_, data_stage_5__4981_, data_stage_5__4980_, data_stage_5__4979_, data_stage_5__4978_, data_stage_5__4977_, data_stage_5__4976_, data_stage_5__4975_, data_stage_5__4974_, data_stage_5__4973_, data_stage_5__4972_, data_stage_5__4971_, data_stage_5__4970_, data_stage_5__4969_, data_stage_5__4968_, data_stage_5__4967_, data_stage_5__4966_, data_stage_5__4965_, data_stage_5__4964_, data_stage_5__4963_, data_stage_5__4962_, data_stage_5__4961_, data_stage_5__4960_, data_stage_5__4959_, data_stage_5__4958_, data_stage_5__4957_, data_stage_5__4956_, data_stage_5__4955_, data_stage_5__4954_, data_stage_5__4953_, data_stage_5__4952_, data_stage_5__4951_, data_stage_5__4950_, data_stage_5__4949_, data_stage_5__4948_, data_stage_5__4947_, data_stage_5__4946_, data_stage_5__4945_, data_stage_5__4944_, data_stage_5__4943_, data_stage_5__4942_, data_stage_5__4941_, data_stage_5__4940_, data_stage_5__4939_, data_stage_5__4938_, data_stage_5__4937_, data_stage_5__4936_, data_stage_5__4935_, data_stage_5__4934_, data_stage_5__4933_, data_stage_5__4932_, data_stage_5__4931_, data_stage_5__4930_, data_stage_5__4929_, data_stage_5__4928_, data_stage_5__4927_, data_stage_5__4926_, data_stage_5__4925_, data_stage_5__4924_, data_stage_5__4923_, data_stage_5__4922_, data_stage_5__4921_, data_stage_5__4920_, data_stage_5__4919_, data_stage_5__4918_, data_stage_5__4917_, data_stage_5__4916_, data_stage_5__4915_, data_stage_5__4914_, data_stage_5__4913_, data_stage_5__4912_, data_stage_5__4911_, data_stage_5__4910_, data_stage_5__4909_, data_stage_5__4908_, data_stage_5__4907_, data_stage_5__4906_, data_stage_5__4905_, data_stage_5__4904_, data_stage_5__4903_, data_stage_5__4902_, data_stage_5__4901_, data_stage_5__4900_, data_stage_5__4899_, data_stage_5__4898_, data_stage_5__4897_, data_stage_5__4896_, data_stage_5__4895_, data_stage_5__4894_, data_stage_5__4893_, data_stage_5__4892_, data_stage_5__4891_, data_stage_5__4890_, data_stage_5__4889_, data_stage_5__4888_, data_stage_5__4887_, data_stage_5__4886_, data_stage_5__4885_, data_stage_5__4884_, data_stage_5__4883_, data_stage_5__4882_, data_stage_5__4881_, data_stage_5__4880_, data_stage_5__4879_, data_stage_5__4878_, data_stage_5__4877_, data_stage_5__4876_, data_stage_5__4875_, data_stage_5__4874_, data_stage_5__4873_, data_stage_5__4872_, data_stage_5__4871_, data_stage_5__4870_, data_stage_5__4869_, data_stage_5__4868_, data_stage_5__4867_, data_stage_5__4866_, data_stage_5__4865_, data_stage_5__4864_, data_stage_5__4863_, data_stage_5__4862_, data_stage_5__4861_, data_stage_5__4860_, data_stage_5__4859_, data_stage_5__4858_, data_stage_5__4857_, data_stage_5__4856_, data_stage_5__4855_, data_stage_5__4854_, data_stage_5__4853_, data_stage_5__4852_, data_stage_5__4851_, data_stage_5__4850_, data_stage_5__4849_, data_stage_5__4848_, data_stage_5__4847_, data_stage_5__4846_, data_stage_5__4845_, data_stage_5__4844_, data_stage_5__4843_, data_stage_5__4842_, data_stage_5__4841_, data_stage_5__4840_, data_stage_5__4839_, data_stage_5__4838_, data_stage_5__4837_, data_stage_5__4836_, data_stage_5__4835_, data_stage_5__4834_, data_stage_5__4833_, data_stage_5__4832_, data_stage_5__4831_, data_stage_5__4830_, data_stage_5__4829_, data_stage_5__4828_, data_stage_5__4827_, data_stage_5__4826_, data_stage_5__4825_, data_stage_5__4824_, data_stage_5__4823_, data_stage_5__4822_, data_stage_5__4821_, data_stage_5__4820_, data_stage_5__4819_, data_stage_5__4818_, data_stage_5__4817_, data_stage_5__4816_, data_stage_5__4815_, data_stage_5__4814_, data_stage_5__4813_, data_stage_5__4812_, data_stage_5__4811_, data_stage_5__4810_, data_stage_5__4809_, data_stage_5__4808_, data_stage_5__4807_, data_stage_5__4806_, data_stage_5__4805_, data_stage_5__4804_, data_stage_5__4803_, data_stage_5__4802_, data_stage_5__4801_, data_stage_5__4800_, data_stage_5__4799_, data_stage_5__4798_, data_stage_5__4797_, data_stage_5__4796_, data_stage_5__4795_, data_stage_5__4794_, data_stage_5__4793_, data_stage_5__4792_, data_stage_5__4791_, data_stage_5__4790_, data_stage_5__4789_, data_stage_5__4788_, data_stage_5__4787_, data_stage_5__4786_, data_stage_5__4785_, data_stage_5__4784_, data_stage_5__4783_, data_stage_5__4782_, data_stage_5__4781_, data_stage_5__4780_, data_stage_5__4779_, data_stage_5__4778_, data_stage_5__4777_, data_stage_5__4776_, data_stage_5__4775_, data_stage_5__4774_, data_stage_5__4773_, data_stage_5__4772_, data_stage_5__4771_, data_stage_5__4770_, data_stage_5__4769_, data_stage_5__4768_, data_stage_5__4767_, data_stage_5__4766_, data_stage_5__4765_, data_stage_5__4764_, data_stage_5__4763_, data_stage_5__4762_, data_stage_5__4761_, data_stage_5__4760_, data_stage_5__4759_, data_stage_5__4758_, data_stage_5__4757_, data_stage_5__4756_, data_stage_5__4755_, data_stage_5__4754_, data_stage_5__4753_, data_stage_5__4752_, data_stage_5__4751_, data_stage_5__4750_, data_stage_5__4749_, data_stage_5__4748_, data_stage_5__4747_, data_stage_5__4746_, data_stage_5__4745_, data_stage_5__4744_, data_stage_5__4743_, data_stage_5__4742_, data_stage_5__4741_, data_stage_5__4740_, data_stage_5__4739_, data_stage_5__4738_, data_stage_5__4737_, data_stage_5__4736_, data_stage_5__4735_, data_stage_5__4734_, data_stage_5__4733_, data_stage_5__4732_, data_stage_5__4731_, data_stage_5__4730_, data_stage_5__4729_, data_stage_5__4728_, data_stage_5__4727_, data_stage_5__4726_, data_stage_5__4725_, data_stage_5__4724_, data_stage_5__4723_, data_stage_5__4722_, data_stage_5__4721_, data_stage_5__4720_, data_stage_5__4719_, data_stage_5__4718_, data_stage_5__4717_, data_stage_5__4716_, data_stage_5__4715_, data_stage_5__4714_, data_stage_5__4713_, data_stage_5__4712_, data_stage_5__4711_, data_stage_5__4710_, data_stage_5__4709_, data_stage_5__4708_, data_stage_5__4707_, data_stage_5__4706_, data_stage_5__4705_, data_stage_5__4704_, data_stage_5__4703_, data_stage_5__4702_, data_stage_5__4701_, data_stage_5__4700_, data_stage_5__4699_, data_stage_5__4698_, data_stage_5__4697_, data_stage_5__4696_, data_stage_5__4695_, data_stage_5__4694_, data_stage_5__4693_, data_stage_5__4692_, data_stage_5__4691_, data_stage_5__4690_, data_stage_5__4689_, data_stage_5__4688_, data_stage_5__4687_, data_stage_5__4686_, data_stage_5__4685_, data_stage_5__4684_, data_stage_5__4683_, data_stage_5__4682_, data_stage_5__4681_, data_stage_5__4680_, data_stage_5__4679_, data_stage_5__4678_, data_stage_5__4677_, data_stage_5__4676_, data_stage_5__4675_, data_stage_5__4674_, data_stage_5__4673_, data_stage_5__4672_, data_stage_5__4671_, data_stage_5__4670_, data_stage_5__4669_, data_stage_5__4668_, data_stage_5__4667_, data_stage_5__4666_, data_stage_5__4665_, data_stage_5__4664_, data_stage_5__4663_, data_stage_5__4662_, data_stage_5__4661_, data_stage_5__4660_, data_stage_5__4659_, data_stage_5__4658_, data_stage_5__4657_, data_stage_5__4656_, data_stage_5__4655_, data_stage_5__4654_, data_stage_5__4653_, data_stage_5__4652_, data_stage_5__4651_, data_stage_5__4650_, data_stage_5__4649_, data_stage_5__4648_, data_stage_5__4647_, data_stage_5__4646_, data_stage_5__4645_, data_stage_5__4644_, data_stage_5__4643_, data_stage_5__4642_, data_stage_5__4641_, data_stage_5__4640_, data_stage_5__4639_, data_stage_5__4638_, data_stage_5__4637_, data_stage_5__4636_, data_stage_5__4635_, data_stage_5__4634_, data_stage_5__4633_, data_stage_5__4632_, data_stage_5__4631_, data_stage_5__4630_, data_stage_5__4629_, data_stage_5__4628_, data_stage_5__4627_, data_stage_5__4626_, data_stage_5__4625_, data_stage_5__4624_, data_stage_5__4623_, data_stage_5__4622_, data_stage_5__4621_, data_stage_5__4620_, data_stage_5__4619_, data_stage_5__4618_, data_stage_5__4617_, data_stage_5__4616_, data_stage_5__4615_, data_stage_5__4614_, data_stage_5__4613_, data_stage_5__4612_, data_stage_5__4611_, data_stage_5__4610_, data_stage_5__4609_, data_stage_5__4608_, data_stage_5__4607_, data_stage_5__4606_, data_stage_5__4605_, data_stage_5__4604_, data_stage_5__4603_, data_stage_5__4602_, data_stage_5__4601_, data_stage_5__4600_, data_stage_5__4599_, data_stage_5__4598_, data_stage_5__4597_, data_stage_5__4596_, data_stage_5__4595_, data_stage_5__4594_, data_stage_5__4593_, data_stage_5__4592_, data_stage_5__4591_, data_stage_5__4590_, data_stage_5__4589_, data_stage_5__4588_, data_stage_5__4587_, data_stage_5__4586_, data_stage_5__4585_, data_stage_5__4584_, data_stage_5__4583_, data_stage_5__4582_, data_stage_5__4581_, data_stage_5__4580_, data_stage_5__4579_, data_stage_5__4578_, data_stage_5__4577_, data_stage_5__4576_, data_stage_5__4575_, data_stage_5__4574_, data_stage_5__4573_, data_stage_5__4572_, data_stage_5__4571_, data_stage_5__4570_, data_stage_5__4569_, data_stage_5__4568_, data_stage_5__4567_, data_stage_5__4566_, data_stage_5__4565_, data_stage_5__4564_, data_stage_5__4563_, data_stage_5__4562_, data_stage_5__4561_, data_stage_5__4560_, data_stage_5__4559_, data_stage_5__4558_, data_stage_5__4557_, data_stage_5__4556_, data_stage_5__4555_, data_stage_5__4554_, data_stage_5__4553_, data_stage_5__4552_, data_stage_5__4551_, data_stage_5__4550_, data_stage_5__4549_, data_stage_5__4548_, data_stage_5__4547_, data_stage_5__4546_, data_stage_5__4545_, data_stage_5__4544_, data_stage_5__4543_, data_stage_5__4542_, data_stage_5__4541_, data_stage_5__4540_, data_stage_5__4539_, data_stage_5__4538_, data_stage_5__4537_, data_stage_5__4536_, data_stage_5__4535_, data_stage_5__4534_, data_stage_5__4533_, data_stage_5__4532_, data_stage_5__4531_, data_stage_5__4530_, data_stage_5__4529_, data_stage_5__4528_, data_stage_5__4527_, data_stage_5__4526_, data_stage_5__4525_, data_stage_5__4524_, data_stage_5__4523_, data_stage_5__4522_, data_stage_5__4521_, data_stage_5__4520_, data_stage_5__4519_, data_stage_5__4518_, data_stage_5__4517_, data_stage_5__4516_, data_stage_5__4515_, data_stage_5__4514_, data_stage_5__4513_, data_stage_5__4512_, data_stage_5__4511_, data_stage_5__4510_, data_stage_5__4509_, data_stage_5__4508_, data_stage_5__4507_, data_stage_5__4506_, data_stage_5__4505_, data_stage_5__4504_, data_stage_5__4503_, data_stage_5__4502_, data_stage_5__4501_, data_stage_5__4500_, data_stage_5__4499_, data_stage_5__4498_, data_stage_5__4497_, data_stage_5__4496_, data_stage_5__4495_, data_stage_5__4494_, data_stage_5__4493_, data_stage_5__4492_, data_stage_5__4491_, data_stage_5__4490_, data_stage_5__4489_, data_stage_5__4488_, data_stage_5__4487_, data_stage_5__4486_, data_stage_5__4485_, data_stage_5__4484_, data_stage_5__4483_, data_stage_5__4482_, data_stage_5__4481_, data_stage_5__4480_, data_stage_5__4479_, data_stage_5__4478_, data_stage_5__4477_, data_stage_5__4476_, data_stage_5__4475_, data_stage_5__4474_, data_stage_5__4473_, data_stage_5__4472_, data_stage_5__4471_, data_stage_5__4470_, data_stage_5__4469_, data_stage_5__4468_, data_stage_5__4467_, data_stage_5__4466_, data_stage_5__4465_, data_stage_5__4464_, data_stage_5__4463_, data_stage_5__4462_, data_stage_5__4461_, data_stage_5__4460_, data_stage_5__4459_, data_stage_5__4458_, data_stage_5__4457_, data_stage_5__4456_, data_stage_5__4455_, data_stage_5__4454_, data_stage_5__4453_, data_stage_5__4452_, data_stage_5__4451_, data_stage_5__4450_, data_stage_5__4449_, data_stage_5__4448_, data_stage_5__4447_, data_stage_5__4446_, data_stage_5__4445_, data_stage_5__4444_, data_stage_5__4443_, data_stage_5__4442_, data_stage_5__4441_, data_stage_5__4440_, data_stage_5__4439_, data_stage_5__4438_, data_stage_5__4437_, data_stage_5__4436_, data_stage_5__4435_, data_stage_5__4434_, data_stage_5__4433_, data_stage_5__4432_, data_stage_5__4431_, data_stage_5__4430_, data_stage_5__4429_, data_stage_5__4428_, data_stage_5__4427_, data_stage_5__4426_, data_stage_5__4425_, data_stage_5__4424_, data_stage_5__4423_, data_stage_5__4422_, data_stage_5__4421_, data_stage_5__4420_, data_stage_5__4419_, data_stage_5__4418_, data_stage_5__4417_, data_stage_5__4416_, data_stage_5__4415_, data_stage_5__4414_, data_stage_5__4413_, data_stage_5__4412_, data_stage_5__4411_, data_stage_5__4410_, data_stage_5__4409_, data_stage_5__4408_, data_stage_5__4407_, data_stage_5__4406_, data_stage_5__4405_, data_stage_5__4404_, data_stage_5__4403_, data_stage_5__4402_, data_stage_5__4401_, data_stage_5__4400_, data_stage_5__4399_, data_stage_5__4398_, data_stage_5__4397_, data_stage_5__4396_, data_stage_5__4395_, data_stage_5__4394_, data_stage_5__4393_, data_stage_5__4392_, data_stage_5__4391_, data_stage_5__4390_, data_stage_5__4389_, data_stage_5__4388_, data_stage_5__4387_, data_stage_5__4386_, data_stage_5__4385_, data_stage_5__4384_, data_stage_5__4383_, data_stage_5__4382_, data_stage_5__4381_, data_stage_5__4380_, data_stage_5__4379_, data_stage_5__4378_, data_stage_5__4377_, data_stage_5__4376_, data_stage_5__4375_, data_stage_5__4374_, data_stage_5__4373_, data_stage_5__4372_, data_stage_5__4371_, data_stage_5__4370_, data_stage_5__4369_, data_stage_5__4368_, data_stage_5__4367_, data_stage_5__4366_, data_stage_5__4365_, data_stage_5__4364_, data_stage_5__4363_, data_stage_5__4362_, data_stage_5__4361_, data_stage_5__4360_, data_stage_5__4359_, data_stage_5__4358_, data_stage_5__4357_, data_stage_5__4356_, data_stage_5__4355_, data_stage_5__4354_, data_stage_5__4353_, data_stage_5__4352_, data_stage_5__4351_, data_stage_5__4350_, data_stage_5__4349_, data_stage_5__4348_, data_stage_5__4347_, data_stage_5__4346_, data_stage_5__4345_, data_stage_5__4344_, data_stage_5__4343_, data_stage_5__4342_, data_stage_5__4341_, data_stage_5__4340_, data_stage_5__4339_, data_stage_5__4338_, data_stage_5__4337_, data_stage_5__4336_, data_stage_5__4335_, data_stage_5__4334_, data_stage_5__4333_, data_stage_5__4332_, data_stage_5__4331_, data_stage_5__4330_, data_stage_5__4329_, data_stage_5__4328_, data_stage_5__4327_, data_stage_5__4326_, data_stage_5__4325_, data_stage_5__4324_, data_stage_5__4323_, data_stage_5__4322_, data_stage_5__4321_, data_stage_5__4320_, data_stage_5__4319_, data_stage_5__4318_, data_stage_5__4317_, data_stage_5__4316_, data_stage_5__4315_, data_stage_5__4314_, data_stage_5__4313_, data_stage_5__4312_, data_stage_5__4311_, data_stage_5__4310_, data_stage_5__4309_, data_stage_5__4308_, data_stage_5__4307_, data_stage_5__4306_, data_stage_5__4305_, data_stage_5__4304_, data_stage_5__4303_, data_stage_5__4302_, data_stage_5__4301_, data_stage_5__4300_, data_stage_5__4299_, data_stage_5__4298_, data_stage_5__4297_, data_stage_5__4296_, data_stage_5__4295_, data_stage_5__4294_, data_stage_5__4293_, data_stage_5__4292_, data_stage_5__4291_, data_stage_5__4290_, data_stage_5__4289_, data_stage_5__4288_, data_stage_5__4287_, data_stage_5__4286_, data_stage_5__4285_, data_stage_5__4284_, data_stage_5__4283_, data_stage_5__4282_, data_stage_5__4281_, data_stage_5__4280_, data_stage_5__4279_, data_stage_5__4278_, data_stage_5__4277_, data_stage_5__4276_, data_stage_5__4275_, data_stage_5__4274_, data_stage_5__4273_, data_stage_5__4272_, data_stage_5__4271_, data_stage_5__4270_, data_stage_5__4269_, data_stage_5__4268_, data_stage_5__4267_, data_stage_5__4266_, data_stage_5__4265_, data_stage_5__4264_, data_stage_5__4263_, data_stage_5__4262_, data_stage_5__4261_, data_stage_5__4260_, data_stage_5__4259_, data_stage_5__4258_, data_stage_5__4257_, data_stage_5__4256_, data_stage_5__4255_, data_stage_5__4254_, data_stage_5__4253_, data_stage_5__4252_, data_stage_5__4251_, data_stage_5__4250_, data_stage_5__4249_, data_stage_5__4248_, data_stage_5__4247_, data_stage_5__4246_, data_stage_5__4245_, data_stage_5__4244_, data_stage_5__4243_, data_stage_5__4242_, data_stage_5__4241_, data_stage_5__4240_, data_stage_5__4239_, data_stage_5__4238_, data_stage_5__4237_, data_stage_5__4236_, data_stage_5__4235_, data_stage_5__4234_, data_stage_5__4233_, data_stage_5__4232_, data_stage_5__4231_, data_stage_5__4230_, data_stage_5__4229_, data_stage_5__4228_, data_stage_5__4227_, data_stage_5__4226_, data_stage_5__4225_, data_stage_5__4224_, data_stage_5__4223_, data_stage_5__4222_, data_stage_5__4221_, data_stage_5__4220_, data_stage_5__4219_, data_stage_5__4218_, data_stage_5__4217_, data_stage_5__4216_, data_stage_5__4215_, data_stage_5__4214_, data_stage_5__4213_, data_stage_5__4212_, data_stage_5__4211_, data_stage_5__4210_, data_stage_5__4209_, data_stage_5__4208_, data_stage_5__4207_, data_stage_5__4206_, data_stage_5__4205_, data_stage_5__4204_, data_stage_5__4203_, data_stage_5__4202_, data_stage_5__4201_, data_stage_5__4200_, data_stage_5__4199_, data_stage_5__4198_, data_stage_5__4197_, data_stage_5__4196_, data_stage_5__4195_, data_stage_5__4194_, data_stage_5__4193_, data_stage_5__4192_, data_stage_5__4191_, data_stage_5__4190_, data_stage_5__4189_, data_stage_5__4188_, data_stage_5__4187_, data_stage_5__4186_, data_stage_5__4185_, data_stage_5__4184_, data_stage_5__4183_, data_stage_5__4182_, data_stage_5__4181_, data_stage_5__4180_, data_stage_5__4179_, data_stage_5__4178_, data_stage_5__4177_, data_stage_5__4176_, data_stage_5__4175_, data_stage_5__4174_, data_stage_5__4173_, data_stage_5__4172_, data_stage_5__4171_, data_stage_5__4170_, data_stage_5__4169_, data_stage_5__4168_, data_stage_5__4167_, data_stage_5__4166_, data_stage_5__4165_, data_stage_5__4164_, data_stage_5__4163_, data_stage_5__4162_, data_stage_5__4161_, data_stage_5__4160_, data_stage_5__4159_, data_stage_5__4158_, data_stage_5__4157_, data_stage_5__4156_, data_stage_5__4155_, data_stage_5__4154_, data_stage_5__4153_, data_stage_5__4152_, data_stage_5__4151_, data_stage_5__4150_, data_stage_5__4149_, data_stage_5__4148_, data_stage_5__4147_, data_stage_5__4146_, data_stage_5__4145_, data_stage_5__4144_, data_stage_5__4143_, data_stage_5__4142_, data_stage_5__4141_, data_stage_5__4140_, data_stage_5__4139_, data_stage_5__4138_, data_stage_5__4137_, data_stage_5__4136_, data_stage_5__4135_, data_stage_5__4134_, data_stage_5__4133_, data_stage_5__4132_, data_stage_5__4131_, data_stage_5__4130_, data_stage_5__4129_, data_stage_5__4128_, data_stage_5__4127_, data_stage_5__4126_, data_stage_5__4125_, data_stage_5__4124_, data_stage_5__4123_, data_stage_5__4122_, data_stage_5__4121_, data_stage_5__4120_, data_stage_5__4119_, data_stage_5__4118_, data_stage_5__4117_, data_stage_5__4116_, data_stage_5__4115_, data_stage_5__4114_, data_stage_5__4113_, data_stage_5__4112_, data_stage_5__4111_, data_stage_5__4110_, data_stage_5__4109_, data_stage_5__4108_, data_stage_5__4107_, data_stage_5__4106_, data_stage_5__4105_, data_stage_5__4104_, data_stage_5__4103_, data_stage_5__4102_, data_stage_5__4101_, data_stage_5__4100_, data_stage_5__4099_, data_stage_5__4098_, data_stage_5__4097_, data_stage_5__4096_ })
  );


  bsg_swap_width_p4096
  mux_stage_5__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_5__8191_, data_stage_5__8190_, data_stage_5__8189_, data_stage_5__8188_, data_stage_5__8187_, data_stage_5__8186_, data_stage_5__8185_, data_stage_5__8184_, data_stage_5__8183_, data_stage_5__8182_, data_stage_5__8181_, data_stage_5__8180_, data_stage_5__8179_, data_stage_5__8178_, data_stage_5__8177_, data_stage_5__8176_, data_stage_5__8175_, data_stage_5__8174_, data_stage_5__8173_, data_stage_5__8172_, data_stage_5__8171_, data_stage_5__8170_, data_stage_5__8169_, data_stage_5__8168_, data_stage_5__8167_, data_stage_5__8166_, data_stage_5__8165_, data_stage_5__8164_, data_stage_5__8163_, data_stage_5__8162_, data_stage_5__8161_, data_stage_5__8160_, data_stage_5__8159_, data_stage_5__8158_, data_stage_5__8157_, data_stage_5__8156_, data_stage_5__8155_, data_stage_5__8154_, data_stage_5__8153_, data_stage_5__8152_, data_stage_5__8151_, data_stage_5__8150_, data_stage_5__8149_, data_stage_5__8148_, data_stage_5__8147_, data_stage_5__8146_, data_stage_5__8145_, data_stage_5__8144_, data_stage_5__8143_, data_stage_5__8142_, data_stage_5__8141_, data_stage_5__8140_, data_stage_5__8139_, data_stage_5__8138_, data_stage_5__8137_, data_stage_5__8136_, data_stage_5__8135_, data_stage_5__8134_, data_stage_5__8133_, data_stage_5__8132_, data_stage_5__8131_, data_stage_5__8130_, data_stage_5__8129_, data_stage_5__8128_, data_stage_5__8127_, data_stage_5__8126_, data_stage_5__8125_, data_stage_5__8124_, data_stage_5__8123_, data_stage_5__8122_, data_stage_5__8121_, data_stage_5__8120_, data_stage_5__8119_, data_stage_5__8118_, data_stage_5__8117_, data_stage_5__8116_, data_stage_5__8115_, data_stage_5__8114_, data_stage_5__8113_, data_stage_5__8112_, data_stage_5__8111_, data_stage_5__8110_, data_stage_5__8109_, data_stage_5__8108_, data_stage_5__8107_, data_stage_5__8106_, data_stage_5__8105_, data_stage_5__8104_, data_stage_5__8103_, data_stage_5__8102_, data_stage_5__8101_, data_stage_5__8100_, data_stage_5__8099_, data_stage_5__8098_, data_stage_5__8097_, data_stage_5__8096_, data_stage_5__8095_, data_stage_5__8094_, data_stage_5__8093_, data_stage_5__8092_, data_stage_5__8091_, data_stage_5__8090_, data_stage_5__8089_, data_stage_5__8088_, data_stage_5__8087_, data_stage_5__8086_, data_stage_5__8085_, data_stage_5__8084_, data_stage_5__8083_, data_stage_5__8082_, data_stage_5__8081_, data_stage_5__8080_, data_stage_5__8079_, data_stage_5__8078_, data_stage_5__8077_, data_stage_5__8076_, data_stage_5__8075_, data_stage_5__8074_, data_stage_5__8073_, data_stage_5__8072_, data_stage_5__8071_, data_stage_5__8070_, data_stage_5__8069_, data_stage_5__8068_, data_stage_5__8067_, data_stage_5__8066_, data_stage_5__8065_, data_stage_5__8064_, data_stage_5__8063_, data_stage_5__8062_, data_stage_5__8061_, data_stage_5__8060_, data_stage_5__8059_, data_stage_5__8058_, data_stage_5__8057_, data_stage_5__8056_, data_stage_5__8055_, data_stage_5__8054_, data_stage_5__8053_, data_stage_5__8052_, data_stage_5__8051_, data_stage_5__8050_, data_stage_5__8049_, data_stage_5__8048_, data_stage_5__8047_, data_stage_5__8046_, data_stage_5__8045_, data_stage_5__8044_, data_stage_5__8043_, data_stage_5__8042_, data_stage_5__8041_, data_stage_5__8040_, data_stage_5__8039_, data_stage_5__8038_, data_stage_5__8037_, data_stage_5__8036_, data_stage_5__8035_, data_stage_5__8034_, data_stage_5__8033_, data_stage_5__8032_, data_stage_5__8031_, data_stage_5__8030_, data_stage_5__8029_, data_stage_5__8028_, data_stage_5__8027_, data_stage_5__8026_, data_stage_5__8025_, data_stage_5__8024_, data_stage_5__8023_, data_stage_5__8022_, data_stage_5__8021_, data_stage_5__8020_, data_stage_5__8019_, data_stage_5__8018_, data_stage_5__8017_, data_stage_5__8016_, data_stage_5__8015_, data_stage_5__8014_, data_stage_5__8013_, data_stage_5__8012_, data_stage_5__8011_, data_stage_5__8010_, data_stage_5__8009_, data_stage_5__8008_, data_stage_5__8007_, data_stage_5__8006_, data_stage_5__8005_, data_stage_5__8004_, data_stage_5__8003_, data_stage_5__8002_, data_stage_5__8001_, data_stage_5__8000_, data_stage_5__7999_, data_stage_5__7998_, data_stage_5__7997_, data_stage_5__7996_, data_stage_5__7995_, data_stage_5__7994_, data_stage_5__7993_, data_stage_5__7992_, data_stage_5__7991_, data_stage_5__7990_, data_stage_5__7989_, data_stage_5__7988_, data_stage_5__7987_, data_stage_5__7986_, data_stage_5__7985_, data_stage_5__7984_, data_stage_5__7983_, data_stage_5__7982_, data_stage_5__7981_, data_stage_5__7980_, data_stage_5__7979_, data_stage_5__7978_, data_stage_5__7977_, data_stage_5__7976_, data_stage_5__7975_, data_stage_5__7974_, data_stage_5__7973_, data_stage_5__7972_, data_stage_5__7971_, data_stage_5__7970_, data_stage_5__7969_, data_stage_5__7968_, data_stage_5__7967_, data_stage_5__7966_, data_stage_5__7965_, data_stage_5__7964_, data_stage_5__7963_, data_stage_5__7962_, data_stage_5__7961_, data_stage_5__7960_, data_stage_5__7959_, data_stage_5__7958_, data_stage_5__7957_, data_stage_5__7956_, data_stage_5__7955_, data_stage_5__7954_, data_stage_5__7953_, data_stage_5__7952_, data_stage_5__7951_, data_stage_5__7950_, data_stage_5__7949_, data_stage_5__7948_, data_stage_5__7947_, data_stage_5__7946_, data_stage_5__7945_, data_stage_5__7944_, data_stage_5__7943_, data_stage_5__7942_, data_stage_5__7941_, data_stage_5__7940_, data_stage_5__7939_, data_stage_5__7938_, data_stage_5__7937_, data_stage_5__7936_, data_stage_5__7935_, data_stage_5__7934_, data_stage_5__7933_, data_stage_5__7932_, data_stage_5__7931_, data_stage_5__7930_, data_stage_5__7929_, data_stage_5__7928_, data_stage_5__7927_, data_stage_5__7926_, data_stage_5__7925_, data_stage_5__7924_, data_stage_5__7923_, data_stage_5__7922_, data_stage_5__7921_, data_stage_5__7920_, data_stage_5__7919_, data_stage_5__7918_, data_stage_5__7917_, data_stage_5__7916_, data_stage_5__7915_, data_stage_5__7914_, data_stage_5__7913_, data_stage_5__7912_, data_stage_5__7911_, data_stage_5__7910_, data_stage_5__7909_, data_stage_5__7908_, data_stage_5__7907_, data_stage_5__7906_, data_stage_5__7905_, data_stage_5__7904_, data_stage_5__7903_, data_stage_5__7902_, data_stage_5__7901_, data_stage_5__7900_, data_stage_5__7899_, data_stage_5__7898_, data_stage_5__7897_, data_stage_5__7896_, data_stage_5__7895_, data_stage_5__7894_, data_stage_5__7893_, data_stage_5__7892_, data_stage_5__7891_, data_stage_5__7890_, data_stage_5__7889_, data_stage_5__7888_, data_stage_5__7887_, data_stage_5__7886_, data_stage_5__7885_, data_stage_5__7884_, data_stage_5__7883_, data_stage_5__7882_, data_stage_5__7881_, data_stage_5__7880_, data_stage_5__7879_, data_stage_5__7878_, data_stage_5__7877_, data_stage_5__7876_, data_stage_5__7875_, data_stage_5__7874_, data_stage_5__7873_, data_stage_5__7872_, data_stage_5__7871_, data_stage_5__7870_, data_stage_5__7869_, data_stage_5__7868_, data_stage_5__7867_, data_stage_5__7866_, data_stage_5__7865_, data_stage_5__7864_, data_stage_5__7863_, data_stage_5__7862_, data_stage_5__7861_, data_stage_5__7860_, data_stage_5__7859_, data_stage_5__7858_, data_stage_5__7857_, data_stage_5__7856_, data_stage_5__7855_, data_stage_5__7854_, data_stage_5__7853_, data_stage_5__7852_, data_stage_5__7851_, data_stage_5__7850_, data_stage_5__7849_, data_stage_5__7848_, data_stage_5__7847_, data_stage_5__7846_, data_stage_5__7845_, data_stage_5__7844_, data_stage_5__7843_, data_stage_5__7842_, data_stage_5__7841_, data_stage_5__7840_, data_stage_5__7839_, data_stage_5__7838_, data_stage_5__7837_, data_stage_5__7836_, data_stage_5__7835_, data_stage_5__7834_, data_stage_5__7833_, data_stage_5__7832_, data_stage_5__7831_, data_stage_5__7830_, data_stage_5__7829_, data_stage_5__7828_, data_stage_5__7827_, data_stage_5__7826_, data_stage_5__7825_, data_stage_5__7824_, data_stage_5__7823_, data_stage_5__7822_, data_stage_5__7821_, data_stage_5__7820_, data_stage_5__7819_, data_stage_5__7818_, data_stage_5__7817_, data_stage_5__7816_, data_stage_5__7815_, data_stage_5__7814_, data_stage_5__7813_, data_stage_5__7812_, data_stage_5__7811_, data_stage_5__7810_, data_stage_5__7809_, data_stage_5__7808_, data_stage_5__7807_, data_stage_5__7806_, data_stage_5__7805_, data_stage_5__7804_, data_stage_5__7803_, data_stage_5__7802_, data_stage_5__7801_, data_stage_5__7800_, data_stage_5__7799_, data_stage_5__7798_, data_stage_5__7797_, data_stage_5__7796_, data_stage_5__7795_, data_stage_5__7794_, data_stage_5__7793_, data_stage_5__7792_, data_stage_5__7791_, data_stage_5__7790_, data_stage_5__7789_, data_stage_5__7788_, data_stage_5__7787_, data_stage_5__7786_, data_stage_5__7785_, data_stage_5__7784_, data_stage_5__7783_, data_stage_5__7782_, data_stage_5__7781_, data_stage_5__7780_, data_stage_5__7779_, data_stage_5__7778_, data_stage_5__7777_, data_stage_5__7776_, data_stage_5__7775_, data_stage_5__7774_, data_stage_5__7773_, data_stage_5__7772_, data_stage_5__7771_, data_stage_5__7770_, data_stage_5__7769_, data_stage_5__7768_, data_stage_5__7767_, data_stage_5__7766_, data_stage_5__7765_, data_stage_5__7764_, data_stage_5__7763_, data_stage_5__7762_, data_stage_5__7761_, data_stage_5__7760_, data_stage_5__7759_, data_stage_5__7758_, data_stage_5__7757_, data_stage_5__7756_, data_stage_5__7755_, data_stage_5__7754_, data_stage_5__7753_, data_stage_5__7752_, data_stage_5__7751_, data_stage_5__7750_, data_stage_5__7749_, data_stage_5__7748_, data_stage_5__7747_, data_stage_5__7746_, data_stage_5__7745_, data_stage_5__7744_, data_stage_5__7743_, data_stage_5__7742_, data_stage_5__7741_, data_stage_5__7740_, data_stage_5__7739_, data_stage_5__7738_, data_stage_5__7737_, data_stage_5__7736_, data_stage_5__7735_, data_stage_5__7734_, data_stage_5__7733_, data_stage_5__7732_, data_stage_5__7731_, data_stage_5__7730_, data_stage_5__7729_, data_stage_5__7728_, data_stage_5__7727_, data_stage_5__7726_, data_stage_5__7725_, data_stage_5__7724_, data_stage_5__7723_, data_stage_5__7722_, data_stage_5__7721_, data_stage_5__7720_, data_stage_5__7719_, data_stage_5__7718_, data_stage_5__7717_, data_stage_5__7716_, data_stage_5__7715_, data_stage_5__7714_, data_stage_5__7713_, data_stage_5__7712_, data_stage_5__7711_, data_stage_5__7710_, data_stage_5__7709_, data_stage_5__7708_, data_stage_5__7707_, data_stage_5__7706_, data_stage_5__7705_, data_stage_5__7704_, data_stage_5__7703_, data_stage_5__7702_, data_stage_5__7701_, data_stage_5__7700_, data_stage_5__7699_, data_stage_5__7698_, data_stage_5__7697_, data_stage_5__7696_, data_stage_5__7695_, data_stage_5__7694_, data_stage_5__7693_, data_stage_5__7692_, data_stage_5__7691_, data_stage_5__7690_, data_stage_5__7689_, data_stage_5__7688_, data_stage_5__7687_, data_stage_5__7686_, data_stage_5__7685_, data_stage_5__7684_, data_stage_5__7683_, data_stage_5__7682_, data_stage_5__7681_, data_stage_5__7680_, data_stage_5__7679_, data_stage_5__7678_, data_stage_5__7677_, data_stage_5__7676_, data_stage_5__7675_, data_stage_5__7674_, data_stage_5__7673_, data_stage_5__7672_, data_stage_5__7671_, data_stage_5__7670_, data_stage_5__7669_, data_stage_5__7668_, data_stage_5__7667_, data_stage_5__7666_, data_stage_5__7665_, data_stage_5__7664_, data_stage_5__7663_, data_stage_5__7662_, data_stage_5__7661_, data_stage_5__7660_, data_stage_5__7659_, data_stage_5__7658_, data_stage_5__7657_, data_stage_5__7656_, data_stage_5__7655_, data_stage_5__7654_, data_stage_5__7653_, data_stage_5__7652_, data_stage_5__7651_, data_stage_5__7650_, data_stage_5__7649_, data_stage_5__7648_, data_stage_5__7647_, data_stage_5__7646_, data_stage_5__7645_, data_stage_5__7644_, data_stage_5__7643_, data_stage_5__7642_, data_stage_5__7641_, data_stage_5__7640_, data_stage_5__7639_, data_stage_5__7638_, data_stage_5__7637_, data_stage_5__7636_, data_stage_5__7635_, data_stage_5__7634_, data_stage_5__7633_, data_stage_5__7632_, data_stage_5__7631_, data_stage_5__7630_, data_stage_5__7629_, data_stage_5__7628_, data_stage_5__7627_, data_stage_5__7626_, data_stage_5__7625_, data_stage_5__7624_, data_stage_5__7623_, data_stage_5__7622_, data_stage_5__7621_, data_stage_5__7620_, data_stage_5__7619_, data_stage_5__7618_, data_stage_5__7617_, data_stage_5__7616_, data_stage_5__7615_, data_stage_5__7614_, data_stage_5__7613_, data_stage_5__7612_, data_stage_5__7611_, data_stage_5__7610_, data_stage_5__7609_, data_stage_5__7608_, data_stage_5__7607_, data_stage_5__7606_, data_stage_5__7605_, data_stage_5__7604_, data_stage_5__7603_, data_stage_5__7602_, data_stage_5__7601_, data_stage_5__7600_, data_stage_5__7599_, data_stage_5__7598_, data_stage_5__7597_, data_stage_5__7596_, data_stage_5__7595_, data_stage_5__7594_, data_stage_5__7593_, data_stage_5__7592_, data_stage_5__7591_, data_stage_5__7590_, data_stage_5__7589_, data_stage_5__7588_, data_stage_5__7587_, data_stage_5__7586_, data_stage_5__7585_, data_stage_5__7584_, data_stage_5__7583_, data_stage_5__7582_, data_stage_5__7581_, data_stage_5__7580_, data_stage_5__7579_, data_stage_5__7578_, data_stage_5__7577_, data_stage_5__7576_, data_stage_5__7575_, data_stage_5__7574_, data_stage_5__7573_, data_stage_5__7572_, data_stage_5__7571_, data_stage_5__7570_, data_stage_5__7569_, data_stage_5__7568_, data_stage_5__7567_, data_stage_5__7566_, data_stage_5__7565_, data_stage_5__7564_, data_stage_5__7563_, data_stage_5__7562_, data_stage_5__7561_, data_stage_5__7560_, data_stage_5__7559_, data_stage_5__7558_, data_stage_5__7557_, data_stage_5__7556_, data_stage_5__7555_, data_stage_5__7554_, data_stage_5__7553_, data_stage_5__7552_, data_stage_5__7551_, data_stage_5__7550_, data_stage_5__7549_, data_stage_5__7548_, data_stage_5__7547_, data_stage_5__7546_, data_stage_5__7545_, data_stage_5__7544_, data_stage_5__7543_, data_stage_5__7542_, data_stage_5__7541_, data_stage_5__7540_, data_stage_5__7539_, data_stage_5__7538_, data_stage_5__7537_, data_stage_5__7536_, data_stage_5__7535_, data_stage_5__7534_, data_stage_5__7533_, data_stage_5__7532_, data_stage_5__7531_, data_stage_5__7530_, data_stage_5__7529_, data_stage_5__7528_, data_stage_5__7527_, data_stage_5__7526_, data_stage_5__7525_, data_stage_5__7524_, data_stage_5__7523_, data_stage_5__7522_, data_stage_5__7521_, data_stage_5__7520_, data_stage_5__7519_, data_stage_5__7518_, data_stage_5__7517_, data_stage_5__7516_, data_stage_5__7515_, data_stage_5__7514_, data_stage_5__7513_, data_stage_5__7512_, data_stage_5__7511_, data_stage_5__7510_, data_stage_5__7509_, data_stage_5__7508_, data_stage_5__7507_, data_stage_5__7506_, data_stage_5__7505_, data_stage_5__7504_, data_stage_5__7503_, data_stage_5__7502_, data_stage_5__7501_, data_stage_5__7500_, data_stage_5__7499_, data_stage_5__7498_, data_stage_5__7497_, data_stage_5__7496_, data_stage_5__7495_, data_stage_5__7494_, data_stage_5__7493_, data_stage_5__7492_, data_stage_5__7491_, data_stage_5__7490_, data_stage_5__7489_, data_stage_5__7488_, data_stage_5__7487_, data_stage_5__7486_, data_stage_5__7485_, data_stage_5__7484_, data_stage_5__7483_, data_stage_5__7482_, data_stage_5__7481_, data_stage_5__7480_, data_stage_5__7479_, data_stage_5__7478_, data_stage_5__7477_, data_stage_5__7476_, data_stage_5__7475_, data_stage_5__7474_, data_stage_5__7473_, data_stage_5__7472_, data_stage_5__7471_, data_stage_5__7470_, data_stage_5__7469_, data_stage_5__7468_, data_stage_5__7467_, data_stage_5__7466_, data_stage_5__7465_, data_stage_5__7464_, data_stage_5__7463_, data_stage_5__7462_, data_stage_5__7461_, data_stage_5__7460_, data_stage_5__7459_, data_stage_5__7458_, data_stage_5__7457_, data_stage_5__7456_, data_stage_5__7455_, data_stage_5__7454_, data_stage_5__7453_, data_stage_5__7452_, data_stage_5__7451_, data_stage_5__7450_, data_stage_5__7449_, data_stage_5__7448_, data_stage_5__7447_, data_stage_5__7446_, data_stage_5__7445_, data_stage_5__7444_, data_stage_5__7443_, data_stage_5__7442_, data_stage_5__7441_, data_stage_5__7440_, data_stage_5__7439_, data_stage_5__7438_, data_stage_5__7437_, data_stage_5__7436_, data_stage_5__7435_, data_stage_5__7434_, data_stage_5__7433_, data_stage_5__7432_, data_stage_5__7431_, data_stage_5__7430_, data_stage_5__7429_, data_stage_5__7428_, data_stage_5__7427_, data_stage_5__7426_, data_stage_5__7425_, data_stage_5__7424_, data_stage_5__7423_, data_stage_5__7422_, data_stage_5__7421_, data_stage_5__7420_, data_stage_5__7419_, data_stage_5__7418_, data_stage_5__7417_, data_stage_5__7416_, data_stage_5__7415_, data_stage_5__7414_, data_stage_5__7413_, data_stage_5__7412_, data_stage_5__7411_, data_stage_5__7410_, data_stage_5__7409_, data_stage_5__7408_, data_stage_5__7407_, data_stage_5__7406_, data_stage_5__7405_, data_stage_5__7404_, data_stage_5__7403_, data_stage_5__7402_, data_stage_5__7401_, data_stage_5__7400_, data_stage_5__7399_, data_stage_5__7398_, data_stage_5__7397_, data_stage_5__7396_, data_stage_5__7395_, data_stage_5__7394_, data_stage_5__7393_, data_stage_5__7392_, data_stage_5__7391_, data_stage_5__7390_, data_stage_5__7389_, data_stage_5__7388_, data_stage_5__7387_, data_stage_5__7386_, data_stage_5__7385_, data_stage_5__7384_, data_stage_5__7383_, data_stage_5__7382_, data_stage_5__7381_, data_stage_5__7380_, data_stage_5__7379_, data_stage_5__7378_, data_stage_5__7377_, data_stage_5__7376_, data_stage_5__7375_, data_stage_5__7374_, data_stage_5__7373_, data_stage_5__7372_, data_stage_5__7371_, data_stage_5__7370_, data_stage_5__7369_, data_stage_5__7368_, data_stage_5__7367_, data_stage_5__7366_, data_stage_5__7365_, data_stage_5__7364_, data_stage_5__7363_, data_stage_5__7362_, data_stage_5__7361_, data_stage_5__7360_, data_stage_5__7359_, data_stage_5__7358_, data_stage_5__7357_, data_stage_5__7356_, data_stage_5__7355_, data_stage_5__7354_, data_stage_5__7353_, data_stage_5__7352_, data_stage_5__7351_, data_stage_5__7350_, data_stage_5__7349_, data_stage_5__7348_, data_stage_5__7347_, data_stage_5__7346_, data_stage_5__7345_, data_stage_5__7344_, data_stage_5__7343_, data_stage_5__7342_, data_stage_5__7341_, data_stage_5__7340_, data_stage_5__7339_, data_stage_5__7338_, data_stage_5__7337_, data_stage_5__7336_, data_stage_5__7335_, data_stage_5__7334_, data_stage_5__7333_, data_stage_5__7332_, data_stage_5__7331_, data_stage_5__7330_, data_stage_5__7329_, data_stage_5__7328_, data_stage_5__7327_, data_stage_5__7326_, data_stage_5__7325_, data_stage_5__7324_, data_stage_5__7323_, data_stage_5__7322_, data_stage_5__7321_, data_stage_5__7320_, data_stage_5__7319_, data_stage_5__7318_, data_stage_5__7317_, data_stage_5__7316_, data_stage_5__7315_, data_stage_5__7314_, data_stage_5__7313_, data_stage_5__7312_, data_stage_5__7311_, data_stage_5__7310_, data_stage_5__7309_, data_stage_5__7308_, data_stage_5__7307_, data_stage_5__7306_, data_stage_5__7305_, data_stage_5__7304_, data_stage_5__7303_, data_stage_5__7302_, data_stage_5__7301_, data_stage_5__7300_, data_stage_5__7299_, data_stage_5__7298_, data_stage_5__7297_, data_stage_5__7296_, data_stage_5__7295_, data_stage_5__7294_, data_stage_5__7293_, data_stage_5__7292_, data_stage_5__7291_, data_stage_5__7290_, data_stage_5__7289_, data_stage_5__7288_, data_stage_5__7287_, data_stage_5__7286_, data_stage_5__7285_, data_stage_5__7284_, data_stage_5__7283_, data_stage_5__7282_, data_stage_5__7281_, data_stage_5__7280_, data_stage_5__7279_, data_stage_5__7278_, data_stage_5__7277_, data_stage_5__7276_, data_stage_5__7275_, data_stage_5__7274_, data_stage_5__7273_, data_stage_5__7272_, data_stage_5__7271_, data_stage_5__7270_, data_stage_5__7269_, data_stage_5__7268_, data_stage_5__7267_, data_stage_5__7266_, data_stage_5__7265_, data_stage_5__7264_, data_stage_5__7263_, data_stage_5__7262_, data_stage_5__7261_, data_stage_5__7260_, data_stage_5__7259_, data_stage_5__7258_, data_stage_5__7257_, data_stage_5__7256_, data_stage_5__7255_, data_stage_5__7254_, data_stage_5__7253_, data_stage_5__7252_, data_stage_5__7251_, data_stage_5__7250_, data_stage_5__7249_, data_stage_5__7248_, data_stage_5__7247_, data_stage_5__7246_, data_stage_5__7245_, data_stage_5__7244_, data_stage_5__7243_, data_stage_5__7242_, data_stage_5__7241_, data_stage_5__7240_, data_stage_5__7239_, data_stage_5__7238_, data_stage_5__7237_, data_stage_5__7236_, data_stage_5__7235_, data_stage_5__7234_, data_stage_5__7233_, data_stage_5__7232_, data_stage_5__7231_, data_stage_5__7230_, data_stage_5__7229_, data_stage_5__7228_, data_stage_5__7227_, data_stage_5__7226_, data_stage_5__7225_, data_stage_5__7224_, data_stage_5__7223_, data_stage_5__7222_, data_stage_5__7221_, data_stage_5__7220_, data_stage_5__7219_, data_stage_5__7218_, data_stage_5__7217_, data_stage_5__7216_, data_stage_5__7215_, data_stage_5__7214_, data_stage_5__7213_, data_stage_5__7212_, data_stage_5__7211_, data_stage_5__7210_, data_stage_5__7209_, data_stage_5__7208_, data_stage_5__7207_, data_stage_5__7206_, data_stage_5__7205_, data_stage_5__7204_, data_stage_5__7203_, data_stage_5__7202_, data_stage_5__7201_, data_stage_5__7200_, data_stage_5__7199_, data_stage_5__7198_, data_stage_5__7197_, data_stage_5__7196_, data_stage_5__7195_, data_stage_5__7194_, data_stage_5__7193_, data_stage_5__7192_, data_stage_5__7191_, data_stage_5__7190_, data_stage_5__7189_, data_stage_5__7188_, data_stage_5__7187_, data_stage_5__7186_, data_stage_5__7185_, data_stage_5__7184_, data_stage_5__7183_, data_stage_5__7182_, data_stage_5__7181_, data_stage_5__7180_, data_stage_5__7179_, data_stage_5__7178_, data_stage_5__7177_, data_stage_5__7176_, data_stage_5__7175_, data_stage_5__7174_, data_stage_5__7173_, data_stage_5__7172_, data_stage_5__7171_, data_stage_5__7170_, data_stage_5__7169_, data_stage_5__7168_, data_stage_5__7167_, data_stage_5__7166_, data_stage_5__7165_, data_stage_5__7164_, data_stage_5__7163_, data_stage_5__7162_, data_stage_5__7161_, data_stage_5__7160_, data_stage_5__7159_, data_stage_5__7158_, data_stage_5__7157_, data_stage_5__7156_, data_stage_5__7155_, data_stage_5__7154_, data_stage_5__7153_, data_stage_5__7152_, data_stage_5__7151_, data_stage_5__7150_, data_stage_5__7149_, data_stage_5__7148_, data_stage_5__7147_, data_stage_5__7146_, data_stage_5__7145_, data_stage_5__7144_, data_stage_5__7143_, data_stage_5__7142_, data_stage_5__7141_, data_stage_5__7140_, data_stage_5__7139_, data_stage_5__7138_, data_stage_5__7137_, data_stage_5__7136_, data_stage_5__7135_, data_stage_5__7134_, data_stage_5__7133_, data_stage_5__7132_, data_stage_5__7131_, data_stage_5__7130_, data_stage_5__7129_, data_stage_5__7128_, data_stage_5__7127_, data_stage_5__7126_, data_stage_5__7125_, data_stage_5__7124_, data_stage_5__7123_, data_stage_5__7122_, data_stage_5__7121_, data_stage_5__7120_, data_stage_5__7119_, data_stage_5__7118_, data_stage_5__7117_, data_stage_5__7116_, data_stage_5__7115_, data_stage_5__7114_, data_stage_5__7113_, data_stage_5__7112_, data_stage_5__7111_, data_stage_5__7110_, data_stage_5__7109_, data_stage_5__7108_, data_stage_5__7107_, data_stage_5__7106_, data_stage_5__7105_, data_stage_5__7104_, data_stage_5__7103_, data_stage_5__7102_, data_stage_5__7101_, data_stage_5__7100_, data_stage_5__7099_, data_stage_5__7098_, data_stage_5__7097_, data_stage_5__7096_, data_stage_5__7095_, data_stage_5__7094_, data_stage_5__7093_, data_stage_5__7092_, data_stage_5__7091_, data_stage_5__7090_, data_stage_5__7089_, data_stage_5__7088_, data_stage_5__7087_, data_stage_5__7086_, data_stage_5__7085_, data_stage_5__7084_, data_stage_5__7083_, data_stage_5__7082_, data_stage_5__7081_, data_stage_5__7080_, data_stage_5__7079_, data_stage_5__7078_, data_stage_5__7077_, data_stage_5__7076_, data_stage_5__7075_, data_stage_5__7074_, data_stage_5__7073_, data_stage_5__7072_, data_stage_5__7071_, data_stage_5__7070_, data_stage_5__7069_, data_stage_5__7068_, data_stage_5__7067_, data_stage_5__7066_, data_stage_5__7065_, data_stage_5__7064_, data_stage_5__7063_, data_stage_5__7062_, data_stage_5__7061_, data_stage_5__7060_, data_stage_5__7059_, data_stage_5__7058_, data_stage_5__7057_, data_stage_5__7056_, data_stage_5__7055_, data_stage_5__7054_, data_stage_5__7053_, data_stage_5__7052_, data_stage_5__7051_, data_stage_5__7050_, data_stage_5__7049_, data_stage_5__7048_, data_stage_5__7047_, data_stage_5__7046_, data_stage_5__7045_, data_stage_5__7044_, data_stage_5__7043_, data_stage_5__7042_, data_stage_5__7041_, data_stage_5__7040_, data_stage_5__7039_, data_stage_5__7038_, data_stage_5__7037_, data_stage_5__7036_, data_stage_5__7035_, data_stage_5__7034_, data_stage_5__7033_, data_stage_5__7032_, data_stage_5__7031_, data_stage_5__7030_, data_stage_5__7029_, data_stage_5__7028_, data_stage_5__7027_, data_stage_5__7026_, data_stage_5__7025_, data_stage_5__7024_, data_stage_5__7023_, data_stage_5__7022_, data_stage_5__7021_, data_stage_5__7020_, data_stage_5__7019_, data_stage_5__7018_, data_stage_5__7017_, data_stage_5__7016_, data_stage_5__7015_, data_stage_5__7014_, data_stage_5__7013_, data_stage_5__7012_, data_stage_5__7011_, data_stage_5__7010_, data_stage_5__7009_, data_stage_5__7008_, data_stage_5__7007_, data_stage_5__7006_, data_stage_5__7005_, data_stage_5__7004_, data_stage_5__7003_, data_stage_5__7002_, data_stage_5__7001_, data_stage_5__7000_, data_stage_5__6999_, data_stage_5__6998_, data_stage_5__6997_, data_stage_5__6996_, data_stage_5__6995_, data_stage_5__6994_, data_stage_5__6993_, data_stage_5__6992_, data_stage_5__6991_, data_stage_5__6990_, data_stage_5__6989_, data_stage_5__6988_, data_stage_5__6987_, data_stage_5__6986_, data_stage_5__6985_, data_stage_5__6984_, data_stage_5__6983_, data_stage_5__6982_, data_stage_5__6981_, data_stage_5__6980_, data_stage_5__6979_, data_stage_5__6978_, data_stage_5__6977_, data_stage_5__6976_, data_stage_5__6975_, data_stage_5__6974_, data_stage_5__6973_, data_stage_5__6972_, data_stage_5__6971_, data_stage_5__6970_, data_stage_5__6969_, data_stage_5__6968_, data_stage_5__6967_, data_stage_5__6966_, data_stage_5__6965_, data_stage_5__6964_, data_stage_5__6963_, data_stage_5__6962_, data_stage_5__6961_, data_stage_5__6960_, data_stage_5__6959_, data_stage_5__6958_, data_stage_5__6957_, data_stage_5__6956_, data_stage_5__6955_, data_stage_5__6954_, data_stage_5__6953_, data_stage_5__6952_, data_stage_5__6951_, data_stage_5__6950_, data_stage_5__6949_, data_stage_5__6948_, data_stage_5__6947_, data_stage_5__6946_, data_stage_5__6945_, data_stage_5__6944_, data_stage_5__6943_, data_stage_5__6942_, data_stage_5__6941_, data_stage_5__6940_, data_stage_5__6939_, data_stage_5__6938_, data_stage_5__6937_, data_stage_5__6936_, data_stage_5__6935_, data_stage_5__6934_, data_stage_5__6933_, data_stage_5__6932_, data_stage_5__6931_, data_stage_5__6930_, data_stage_5__6929_, data_stage_5__6928_, data_stage_5__6927_, data_stage_5__6926_, data_stage_5__6925_, data_stage_5__6924_, data_stage_5__6923_, data_stage_5__6922_, data_stage_5__6921_, data_stage_5__6920_, data_stage_5__6919_, data_stage_5__6918_, data_stage_5__6917_, data_stage_5__6916_, data_stage_5__6915_, data_stage_5__6914_, data_stage_5__6913_, data_stage_5__6912_, data_stage_5__6911_, data_stage_5__6910_, data_stage_5__6909_, data_stage_5__6908_, data_stage_5__6907_, data_stage_5__6906_, data_stage_5__6905_, data_stage_5__6904_, data_stage_5__6903_, data_stage_5__6902_, data_stage_5__6901_, data_stage_5__6900_, data_stage_5__6899_, data_stage_5__6898_, data_stage_5__6897_, data_stage_5__6896_, data_stage_5__6895_, data_stage_5__6894_, data_stage_5__6893_, data_stage_5__6892_, data_stage_5__6891_, data_stage_5__6890_, data_stage_5__6889_, data_stage_5__6888_, data_stage_5__6887_, data_stage_5__6886_, data_stage_5__6885_, data_stage_5__6884_, data_stage_5__6883_, data_stage_5__6882_, data_stage_5__6881_, data_stage_5__6880_, data_stage_5__6879_, data_stage_5__6878_, data_stage_5__6877_, data_stage_5__6876_, data_stage_5__6875_, data_stage_5__6874_, data_stage_5__6873_, data_stage_5__6872_, data_stage_5__6871_, data_stage_5__6870_, data_stage_5__6869_, data_stage_5__6868_, data_stage_5__6867_, data_stage_5__6866_, data_stage_5__6865_, data_stage_5__6864_, data_stage_5__6863_, data_stage_5__6862_, data_stage_5__6861_, data_stage_5__6860_, data_stage_5__6859_, data_stage_5__6858_, data_stage_5__6857_, data_stage_5__6856_, data_stage_5__6855_, data_stage_5__6854_, data_stage_5__6853_, data_stage_5__6852_, data_stage_5__6851_, data_stage_5__6850_, data_stage_5__6849_, data_stage_5__6848_, data_stage_5__6847_, data_stage_5__6846_, data_stage_5__6845_, data_stage_5__6844_, data_stage_5__6843_, data_stage_5__6842_, data_stage_5__6841_, data_stage_5__6840_, data_stage_5__6839_, data_stage_5__6838_, data_stage_5__6837_, data_stage_5__6836_, data_stage_5__6835_, data_stage_5__6834_, data_stage_5__6833_, data_stage_5__6832_, data_stage_5__6831_, data_stage_5__6830_, data_stage_5__6829_, data_stage_5__6828_, data_stage_5__6827_, data_stage_5__6826_, data_stage_5__6825_, data_stage_5__6824_, data_stage_5__6823_, data_stage_5__6822_, data_stage_5__6821_, data_stage_5__6820_, data_stage_5__6819_, data_stage_5__6818_, data_stage_5__6817_, data_stage_5__6816_, data_stage_5__6815_, data_stage_5__6814_, data_stage_5__6813_, data_stage_5__6812_, data_stage_5__6811_, data_stage_5__6810_, data_stage_5__6809_, data_stage_5__6808_, data_stage_5__6807_, data_stage_5__6806_, data_stage_5__6805_, data_stage_5__6804_, data_stage_5__6803_, data_stage_5__6802_, data_stage_5__6801_, data_stage_5__6800_, data_stage_5__6799_, data_stage_5__6798_, data_stage_5__6797_, data_stage_5__6796_, data_stage_5__6795_, data_stage_5__6794_, data_stage_5__6793_, data_stage_5__6792_, data_stage_5__6791_, data_stage_5__6790_, data_stage_5__6789_, data_stage_5__6788_, data_stage_5__6787_, data_stage_5__6786_, data_stage_5__6785_, data_stage_5__6784_, data_stage_5__6783_, data_stage_5__6782_, data_stage_5__6781_, data_stage_5__6780_, data_stage_5__6779_, data_stage_5__6778_, data_stage_5__6777_, data_stage_5__6776_, data_stage_5__6775_, data_stage_5__6774_, data_stage_5__6773_, data_stage_5__6772_, data_stage_5__6771_, data_stage_5__6770_, data_stage_5__6769_, data_stage_5__6768_, data_stage_5__6767_, data_stage_5__6766_, data_stage_5__6765_, data_stage_5__6764_, data_stage_5__6763_, data_stage_5__6762_, data_stage_5__6761_, data_stage_5__6760_, data_stage_5__6759_, data_stage_5__6758_, data_stage_5__6757_, data_stage_5__6756_, data_stage_5__6755_, data_stage_5__6754_, data_stage_5__6753_, data_stage_5__6752_, data_stage_5__6751_, data_stage_5__6750_, data_stage_5__6749_, data_stage_5__6748_, data_stage_5__6747_, data_stage_5__6746_, data_stage_5__6745_, data_stage_5__6744_, data_stage_5__6743_, data_stage_5__6742_, data_stage_5__6741_, data_stage_5__6740_, data_stage_5__6739_, data_stage_5__6738_, data_stage_5__6737_, data_stage_5__6736_, data_stage_5__6735_, data_stage_5__6734_, data_stage_5__6733_, data_stage_5__6732_, data_stage_5__6731_, data_stage_5__6730_, data_stage_5__6729_, data_stage_5__6728_, data_stage_5__6727_, data_stage_5__6726_, data_stage_5__6725_, data_stage_5__6724_, data_stage_5__6723_, data_stage_5__6722_, data_stage_5__6721_, data_stage_5__6720_, data_stage_5__6719_, data_stage_5__6718_, data_stage_5__6717_, data_stage_5__6716_, data_stage_5__6715_, data_stage_5__6714_, data_stage_5__6713_, data_stage_5__6712_, data_stage_5__6711_, data_stage_5__6710_, data_stage_5__6709_, data_stage_5__6708_, data_stage_5__6707_, data_stage_5__6706_, data_stage_5__6705_, data_stage_5__6704_, data_stage_5__6703_, data_stage_5__6702_, data_stage_5__6701_, data_stage_5__6700_, data_stage_5__6699_, data_stage_5__6698_, data_stage_5__6697_, data_stage_5__6696_, data_stage_5__6695_, data_stage_5__6694_, data_stage_5__6693_, data_stage_5__6692_, data_stage_5__6691_, data_stage_5__6690_, data_stage_5__6689_, data_stage_5__6688_, data_stage_5__6687_, data_stage_5__6686_, data_stage_5__6685_, data_stage_5__6684_, data_stage_5__6683_, data_stage_5__6682_, data_stage_5__6681_, data_stage_5__6680_, data_stage_5__6679_, data_stage_5__6678_, data_stage_5__6677_, data_stage_5__6676_, data_stage_5__6675_, data_stage_5__6674_, data_stage_5__6673_, data_stage_5__6672_, data_stage_5__6671_, data_stage_5__6670_, data_stage_5__6669_, data_stage_5__6668_, data_stage_5__6667_, data_stage_5__6666_, data_stage_5__6665_, data_stage_5__6664_, data_stage_5__6663_, data_stage_5__6662_, data_stage_5__6661_, data_stage_5__6660_, data_stage_5__6659_, data_stage_5__6658_, data_stage_5__6657_, data_stage_5__6656_, data_stage_5__6655_, data_stage_5__6654_, data_stage_5__6653_, data_stage_5__6652_, data_stage_5__6651_, data_stage_5__6650_, data_stage_5__6649_, data_stage_5__6648_, data_stage_5__6647_, data_stage_5__6646_, data_stage_5__6645_, data_stage_5__6644_, data_stage_5__6643_, data_stage_5__6642_, data_stage_5__6641_, data_stage_5__6640_, data_stage_5__6639_, data_stage_5__6638_, data_stage_5__6637_, data_stage_5__6636_, data_stage_5__6635_, data_stage_5__6634_, data_stage_5__6633_, data_stage_5__6632_, data_stage_5__6631_, data_stage_5__6630_, data_stage_5__6629_, data_stage_5__6628_, data_stage_5__6627_, data_stage_5__6626_, data_stage_5__6625_, data_stage_5__6624_, data_stage_5__6623_, data_stage_5__6622_, data_stage_5__6621_, data_stage_5__6620_, data_stage_5__6619_, data_stage_5__6618_, data_stage_5__6617_, data_stage_5__6616_, data_stage_5__6615_, data_stage_5__6614_, data_stage_5__6613_, data_stage_5__6612_, data_stage_5__6611_, data_stage_5__6610_, data_stage_5__6609_, data_stage_5__6608_, data_stage_5__6607_, data_stage_5__6606_, data_stage_5__6605_, data_stage_5__6604_, data_stage_5__6603_, data_stage_5__6602_, data_stage_5__6601_, data_stage_5__6600_, data_stage_5__6599_, data_stage_5__6598_, data_stage_5__6597_, data_stage_5__6596_, data_stage_5__6595_, data_stage_5__6594_, data_stage_5__6593_, data_stage_5__6592_, data_stage_5__6591_, data_stage_5__6590_, data_stage_5__6589_, data_stage_5__6588_, data_stage_5__6587_, data_stage_5__6586_, data_stage_5__6585_, data_stage_5__6584_, data_stage_5__6583_, data_stage_5__6582_, data_stage_5__6581_, data_stage_5__6580_, data_stage_5__6579_, data_stage_5__6578_, data_stage_5__6577_, data_stage_5__6576_, data_stage_5__6575_, data_stage_5__6574_, data_stage_5__6573_, data_stage_5__6572_, data_stage_5__6571_, data_stage_5__6570_, data_stage_5__6569_, data_stage_5__6568_, data_stage_5__6567_, data_stage_5__6566_, data_stage_5__6565_, data_stage_5__6564_, data_stage_5__6563_, data_stage_5__6562_, data_stage_5__6561_, data_stage_5__6560_, data_stage_5__6559_, data_stage_5__6558_, data_stage_5__6557_, data_stage_5__6556_, data_stage_5__6555_, data_stage_5__6554_, data_stage_5__6553_, data_stage_5__6552_, data_stage_5__6551_, data_stage_5__6550_, data_stage_5__6549_, data_stage_5__6548_, data_stage_5__6547_, data_stage_5__6546_, data_stage_5__6545_, data_stage_5__6544_, data_stage_5__6543_, data_stage_5__6542_, data_stage_5__6541_, data_stage_5__6540_, data_stage_5__6539_, data_stage_5__6538_, data_stage_5__6537_, data_stage_5__6536_, data_stage_5__6535_, data_stage_5__6534_, data_stage_5__6533_, data_stage_5__6532_, data_stage_5__6531_, data_stage_5__6530_, data_stage_5__6529_, data_stage_5__6528_, data_stage_5__6527_, data_stage_5__6526_, data_stage_5__6525_, data_stage_5__6524_, data_stage_5__6523_, data_stage_5__6522_, data_stage_5__6521_, data_stage_5__6520_, data_stage_5__6519_, data_stage_5__6518_, data_stage_5__6517_, data_stage_5__6516_, data_stage_5__6515_, data_stage_5__6514_, data_stage_5__6513_, data_stage_5__6512_, data_stage_5__6511_, data_stage_5__6510_, data_stage_5__6509_, data_stage_5__6508_, data_stage_5__6507_, data_stage_5__6506_, data_stage_5__6505_, data_stage_5__6504_, data_stage_5__6503_, data_stage_5__6502_, data_stage_5__6501_, data_stage_5__6500_, data_stage_5__6499_, data_stage_5__6498_, data_stage_5__6497_, data_stage_5__6496_, data_stage_5__6495_, data_stage_5__6494_, data_stage_5__6493_, data_stage_5__6492_, data_stage_5__6491_, data_stage_5__6490_, data_stage_5__6489_, data_stage_5__6488_, data_stage_5__6487_, data_stage_5__6486_, data_stage_5__6485_, data_stage_5__6484_, data_stage_5__6483_, data_stage_5__6482_, data_stage_5__6481_, data_stage_5__6480_, data_stage_5__6479_, data_stage_5__6478_, data_stage_5__6477_, data_stage_5__6476_, data_stage_5__6475_, data_stage_5__6474_, data_stage_5__6473_, data_stage_5__6472_, data_stage_5__6471_, data_stage_5__6470_, data_stage_5__6469_, data_stage_5__6468_, data_stage_5__6467_, data_stage_5__6466_, data_stage_5__6465_, data_stage_5__6464_, data_stage_5__6463_, data_stage_5__6462_, data_stage_5__6461_, data_stage_5__6460_, data_stage_5__6459_, data_stage_5__6458_, data_stage_5__6457_, data_stage_5__6456_, data_stage_5__6455_, data_stage_5__6454_, data_stage_5__6453_, data_stage_5__6452_, data_stage_5__6451_, data_stage_5__6450_, data_stage_5__6449_, data_stage_5__6448_, data_stage_5__6447_, data_stage_5__6446_, data_stage_5__6445_, data_stage_5__6444_, data_stage_5__6443_, data_stage_5__6442_, data_stage_5__6441_, data_stage_5__6440_, data_stage_5__6439_, data_stage_5__6438_, data_stage_5__6437_, data_stage_5__6436_, data_stage_5__6435_, data_stage_5__6434_, data_stage_5__6433_, data_stage_5__6432_, data_stage_5__6431_, data_stage_5__6430_, data_stage_5__6429_, data_stage_5__6428_, data_stage_5__6427_, data_stage_5__6426_, data_stage_5__6425_, data_stage_5__6424_, data_stage_5__6423_, data_stage_5__6422_, data_stage_5__6421_, data_stage_5__6420_, data_stage_5__6419_, data_stage_5__6418_, data_stage_5__6417_, data_stage_5__6416_, data_stage_5__6415_, data_stage_5__6414_, data_stage_5__6413_, data_stage_5__6412_, data_stage_5__6411_, data_stage_5__6410_, data_stage_5__6409_, data_stage_5__6408_, data_stage_5__6407_, data_stage_5__6406_, data_stage_5__6405_, data_stage_5__6404_, data_stage_5__6403_, data_stage_5__6402_, data_stage_5__6401_, data_stage_5__6400_, data_stage_5__6399_, data_stage_5__6398_, data_stage_5__6397_, data_stage_5__6396_, data_stage_5__6395_, data_stage_5__6394_, data_stage_5__6393_, data_stage_5__6392_, data_stage_5__6391_, data_stage_5__6390_, data_stage_5__6389_, data_stage_5__6388_, data_stage_5__6387_, data_stage_5__6386_, data_stage_5__6385_, data_stage_5__6384_, data_stage_5__6383_, data_stage_5__6382_, data_stage_5__6381_, data_stage_5__6380_, data_stage_5__6379_, data_stage_5__6378_, data_stage_5__6377_, data_stage_5__6376_, data_stage_5__6375_, data_stage_5__6374_, data_stage_5__6373_, data_stage_5__6372_, data_stage_5__6371_, data_stage_5__6370_, data_stage_5__6369_, data_stage_5__6368_, data_stage_5__6367_, data_stage_5__6366_, data_stage_5__6365_, data_stage_5__6364_, data_stage_5__6363_, data_stage_5__6362_, data_stage_5__6361_, data_stage_5__6360_, data_stage_5__6359_, data_stage_5__6358_, data_stage_5__6357_, data_stage_5__6356_, data_stage_5__6355_, data_stage_5__6354_, data_stage_5__6353_, data_stage_5__6352_, data_stage_5__6351_, data_stage_5__6350_, data_stage_5__6349_, data_stage_5__6348_, data_stage_5__6347_, data_stage_5__6346_, data_stage_5__6345_, data_stage_5__6344_, data_stage_5__6343_, data_stage_5__6342_, data_stage_5__6341_, data_stage_5__6340_, data_stage_5__6339_, data_stage_5__6338_, data_stage_5__6337_, data_stage_5__6336_, data_stage_5__6335_, data_stage_5__6334_, data_stage_5__6333_, data_stage_5__6332_, data_stage_5__6331_, data_stage_5__6330_, data_stage_5__6329_, data_stage_5__6328_, data_stage_5__6327_, data_stage_5__6326_, data_stage_5__6325_, data_stage_5__6324_, data_stage_5__6323_, data_stage_5__6322_, data_stage_5__6321_, data_stage_5__6320_, data_stage_5__6319_, data_stage_5__6318_, data_stage_5__6317_, data_stage_5__6316_, data_stage_5__6315_, data_stage_5__6314_, data_stage_5__6313_, data_stage_5__6312_, data_stage_5__6311_, data_stage_5__6310_, data_stage_5__6309_, data_stage_5__6308_, data_stage_5__6307_, data_stage_5__6306_, data_stage_5__6305_, data_stage_5__6304_, data_stage_5__6303_, data_stage_5__6302_, data_stage_5__6301_, data_stage_5__6300_, data_stage_5__6299_, data_stage_5__6298_, data_stage_5__6297_, data_stage_5__6296_, data_stage_5__6295_, data_stage_5__6294_, data_stage_5__6293_, data_stage_5__6292_, data_stage_5__6291_, data_stage_5__6290_, data_stage_5__6289_, data_stage_5__6288_, data_stage_5__6287_, data_stage_5__6286_, data_stage_5__6285_, data_stage_5__6284_, data_stage_5__6283_, data_stage_5__6282_, data_stage_5__6281_, data_stage_5__6280_, data_stage_5__6279_, data_stage_5__6278_, data_stage_5__6277_, data_stage_5__6276_, data_stage_5__6275_, data_stage_5__6274_, data_stage_5__6273_, data_stage_5__6272_, data_stage_5__6271_, data_stage_5__6270_, data_stage_5__6269_, data_stage_5__6268_, data_stage_5__6267_, data_stage_5__6266_, data_stage_5__6265_, data_stage_5__6264_, data_stage_5__6263_, data_stage_5__6262_, data_stage_5__6261_, data_stage_5__6260_, data_stage_5__6259_, data_stage_5__6258_, data_stage_5__6257_, data_stage_5__6256_, data_stage_5__6255_, data_stage_5__6254_, data_stage_5__6253_, data_stage_5__6252_, data_stage_5__6251_, data_stage_5__6250_, data_stage_5__6249_, data_stage_5__6248_, data_stage_5__6247_, data_stage_5__6246_, data_stage_5__6245_, data_stage_5__6244_, data_stage_5__6243_, data_stage_5__6242_, data_stage_5__6241_, data_stage_5__6240_, data_stage_5__6239_, data_stage_5__6238_, data_stage_5__6237_, data_stage_5__6236_, data_stage_5__6235_, data_stage_5__6234_, data_stage_5__6233_, data_stage_5__6232_, data_stage_5__6231_, data_stage_5__6230_, data_stage_5__6229_, data_stage_5__6228_, data_stage_5__6227_, data_stage_5__6226_, data_stage_5__6225_, data_stage_5__6224_, data_stage_5__6223_, data_stage_5__6222_, data_stage_5__6221_, data_stage_5__6220_, data_stage_5__6219_, data_stage_5__6218_, data_stage_5__6217_, data_stage_5__6216_, data_stage_5__6215_, data_stage_5__6214_, data_stage_5__6213_, data_stage_5__6212_, data_stage_5__6211_, data_stage_5__6210_, data_stage_5__6209_, data_stage_5__6208_, data_stage_5__6207_, data_stage_5__6206_, data_stage_5__6205_, data_stage_5__6204_, data_stage_5__6203_, data_stage_5__6202_, data_stage_5__6201_, data_stage_5__6200_, data_stage_5__6199_, data_stage_5__6198_, data_stage_5__6197_, data_stage_5__6196_, data_stage_5__6195_, data_stage_5__6194_, data_stage_5__6193_, data_stage_5__6192_, data_stage_5__6191_, data_stage_5__6190_, data_stage_5__6189_, data_stage_5__6188_, data_stage_5__6187_, data_stage_5__6186_, data_stage_5__6185_, data_stage_5__6184_, data_stage_5__6183_, data_stage_5__6182_, data_stage_5__6181_, data_stage_5__6180_, data_stage_5__6179_, data_stage_5__6178_, data_stage_5__6177_, data_stage_5__6176_, data_stage_5__6175_, data_stage_5__6174_, data_stage_5__6173_, data_stage_5__6172_, data_stage_5__6171_, data_stage_5__6170_, data_stage_5__6169_, data_stage_5__6168_, data_stage_5__6167_, data_stage_5__6166_, data_stage_5__6165_, data_stage_5__6164_, data_stage_5__6163_, data_stage_5__6162_, data_stage_5__6161_, data_stage_5__6160_, data_stage_5__6159_, data_stage_5__6158_, data_stage_5__6157_, data_stage_5__6156_, data_stage_5__6155_, data_stage_5__6154_, data_stage_5__6153_, data_stage_5__6152_, data_stage_5__6151_, data_stage_5__6150_, data_stage_5__6149_, data_stage_5__6148_, data_stage_5__6147_, data_stage_5__6146_, data_stage_5__6145_, data_stage_5__6144_, data_stage_5__6143_, data_stage_5__6142_, data_stage_5__6141_, data_stage_5__6140_, data_stage_5__6139_, data_stage_5__6138_, data_stage_5__6137_, data_stage_5__6136_, data_stage_5__6135_, data_stage_5__6134_, data_stage_5__6133_, data_stage_5__6132_, data_stage_5__6131_, data_stage_5__6130_, data_stage_5__6129_, data_stage_5__6128_, data_stage_5__6127_, data_stage_5__6126_, data_stage_5__6125_, data_stage_5__6124_, data_stage_5__6123_, data_stage_5__6122_, data_stage_5__6121_, data_stage_5__6120_, data_stage_5__6119_, data_stage_5__6118_, data_stage_5__6117_, data_stage_5__6116_, data_stage_5__6115_, data_stage_5__6114_, data_stage_5__6113_, data_stage_5__6112_, data_stage_5__6111_, data_stage_5__6110_, data_stage_5__6109_, data_stage_5__6108_, data_stage_5__6107_, data_stage_5__6106_, data_stage_5__6105_, data_stage_5__6104_, data_stage_5__6103_, data_stage_5__6102_, data_stage_5__6101_, data_stage_5__6100_, data_stage_5__6099_, data_stage_5__6098_, data_stage_5__6097_, data_stage_5__6096_, data_stage_5__6095_, data_stage_5__6094_, data_stage_5__6093_, data_stage_5__6092_, data_stage_5__6091_, data_stage_5__6090_, data_stage_5__6089_, data_stage_5__6088_, data_stage_5__6087_, data_stage_5__6086_, data_stage_5__6085_, data_stage_5__6084_, data_stage_5__6083_, data_stage_5__6082_, data_stage_5__6081_, data_stage_5__6080_, data_stage_5__6079_, data_stage_5__6078_, data_stage_5__6077_, data_stage_5__6076_, data_stage_5__6075_, data_stage_5__6074_, data_stage_5__6073_, data_stage_5__6072_, data_stage_5__6071_, data_stage_5__6070_, data_stage_5__6069_, data_stage_5__6068_, data_stage_5__6067_, data_stage_5__6066_, data_stage_5__6065_, data_stage_5__6064_, data_stage_5__6063_, data_stage_5__6062_, data_stage_5__6061_, data_stage_5__6060_, data_stage_5__6059_, data_stage_5__6058_, data_stage_5__6057_, data_stage_5__6056_, data_stage_5__6055_, data_stage_5__6054_, data_stage_5__6053_, data_stage_5__6052_, data_stage_5__6051_, data_stage_5__6050_, data_stage_5__6049_, data_stage_5__6048_, data_stage_5__6047_, data_stage_5__6046_, data_stage_5__6045_, data_stage_5__6044_, data_stage_5__6043_, data_stage_5__6042_, data_stage_5__6041_, data_stage_5__6040_, data_stage_5__6039_, data_stage_5__6038_, data_stage_5__6037_, data_stage_5__6036_, data_stage_5__6035_, data_stage_5__6034_, data_stage_5__6033_, data_stage_5__6032_, data_stage_5__6031_, data_stage_5__6030_, data_stage_5__6029_, data_stage_5__6028_, data_stage_5__6027_, data_stage_5__6026_, data_stage_5__6025_, data_stage_5__6024_, data_stage_5__6023_, data_stage_5__6022_, data_stage_5__6021_, data_stage_5__6020_, data_stage_5__6019_, data_stage_5__6018_, data_stage_5__6017_, data_stage_5__6016_, data_stage_5__6015_, data_stage_5__6014_, data_stage_5__6013_, data_stage_5__6012_, data_stage_5__6011_, data_stage_5__6010_, data_stage_5__6009_, data_stage_5__6008_, data_stage_5__6007_, data_stage_5__6006_, data_stage_5__6005_, data_stage_5__6004_, data_stage_5__6003_, data_stage_5__6002_, data_stage_5__6001_, data_stage_5__6000_, data_stage_5__5999_, data_stage_5__5998_, data_stage_5__5997_, data_stage_5__5996_, data_stage_5__5995_, data_stage_5__5994_, data_stage_5__5993_, data_stage_5__5992_, data_stage_5__5991_, data_stage_5__5990_, data_stage_5__5989_, data_stage_5__5988_, data_stage_5__5987_, data_stage_5__5986_, data_stage_5__5985_, data_stage_5__5984_, data_stage_5__5983_, data_stage_5__5982_, data_stage_5__5981_, data_stage_5__5980_, data_stage_5__5979_, data_stage_5__5978_, data_stage_5__5977_, data_stage_5__5976_, data_stage_5__5975_, data_stage_5__5974_, data_stage_5__5973_, data_stage_5__5972_, data_stage_5__5971_, data_stage_5__5970_, data_stage_5__5969_, data_stage_5__5968_, data_stage_5__5967_, data_stage_5__5966_, data_stage_5__5965_, data_stage_5__5964_, data_stage_5__5963_, data_stage_5__5962_, data_stage_5__5961_, data_stage_5__5960_, data_stage_5__5959_, data_stage_5__5958_, data_stage_5__5957_, data_stage_5__5956_, data_stage_5__5955_, data_stage_5__5954_, data_stage_5__5953_, data_stage_5__5952_, data_stage_5__5951_, data_stage_5__5950_, data_stage_5__5949_, data_stage_5__5948_, data_stage_5__5947_, data_stage_5__5946_, data_stage_5__5945_, data_stage_5__5944_, data_stage_5__5943_, data_stage_5__5942_, data_stage_5__5941_, data_stage_5__5940_, data_stage_5__5939_, data_stage_5__5938_, data_stage_5__5937_, data_stage_5__5936_, data_stage_5__5935_, data_stage_5__5934_, data_stage_5__5933_, data_stage_5__5932_, data_stage_5__5931_, data_stage_5__5930_, data_stage_5__5929_, data_stage_5__5928_, data_stage_5__5927_, data_stage_5__5926_, data_stage_5__5925_, data_stage_5__5924_, data_stage_5__5923_, data_stage_5__5922_, data_stage_5__5921_, data_stage_5__5920_, data_stage_5__5919_, data_stage_5__5918_, data_stage_5__5917_, data_stage_5__5916_, data_stage_5__5915_, data_stage_5__5914_, data_stage_5__5913_, data_stage_5__5912_, data_stage_5__5911_, data_stage_5__5910_, data_stage_5__5909_, data_stage_5__5908_, data_stage_5__5907_, data_stage_5__5906_, data_stage_5__5905_, data_stage_5__5904_, data_stage_5__5903_, data_stage_5__5902_, data_stage_5__5901_, data_stage_5__5900_, data_stage_5__5899_, data_stage_5__5898_, data_stage_5__5897_, data_stage_5__5896_, data_stage_5__5895_, data_stage_5__5894_, data_stage_5__5893_, data_stage_5__5892_, data_stage_5__5891_, data_stage_5__5890_, data_stage_5__5889_, data_stage_5__5888_, data_stage_5__5887_, data_stage_5__5886_, data_stage_5__5885_, data_stage_5__5884_, data_stage_5__5883_, data_stage_5__5882_, data_stage_5__5881_, data_stage_5__5880_, data_stage_5__5879_, data_stage_5__5878_, data_stage_5__5877_, data_stage_5__5876_, data_stage_5__5875_, data_stage_5__5874_, data_stage_5__5873_, data_stage_5__5872_, data_stage_5__5871_, data_stage_5__5870_, data_stage_5__5869_, data_stage_5__5868_, data_stage_5__5867_, data_stage_5__5866_, data_stage_5__5865_, data_stage_5__5864_, data_stage_5__5863_, data_stage_5__5862_, data_stage_5__5861_, data_stage_5__5860_, data_stage_5__5859_, data_stage_5__5858_, data_stage_5__5857_, data_stage_5__5856_, data_stage_5__5855_, data_stage_5__5854_, data_stage_5__5853_, data_stage_5__5852_, data_stage_5__5851_, data_stage_5__5850_, data_stage_5__5849_, data_stage_5__5848_, data_stage_5__5847_, data_stage_5__5846_, data_stage_5__5845_, data_stage_5__5844_, data_stage_5__5843_, data_stage_5__5842_, data_stage_5__5841_, data_stage_5__5840_, data_stage_5__5839_, data_stage_5__5838_, data_stage_5__5837_, data_stage_5__5836_, data_stage_5__5835_, data_stage_5__5834_, data_stage_5__5833_, data_stage_5__5832_, data_stage_5__5831_, data_stage_5__5830_, data_stage_5__5829_, data_stage_5__5828_, data_stage_5__5827_, data_stage_5__5826_, data_stage_5__5825_, data_stage_5__5824_, data_stage_5__5823_, data_stage_5__5822_, data_stage_5__5821_, data_stage_5__5820_, data_stage_5__5819_, data_stage_5__5818_, data_stage_5__5817_, data_stage_5__5816_, data_stage_5__5815_, data_stage_5__5814_, data_stage_5__5813_, data_stage_5__5812_, data_stage_5__5811_, data_stage_5__5810_, data_stage_5__5809_, data_stage_5__5808_, data_stage_5__5807_, data_stage_5__5806_, data_stage_5__5805_, data_stage_5__5804_, data_stage_5__5803_, data_stage_5__5802_, data_stage_5__5801_, data_stage_5__5800_, data_stage_5__5799_, data_stage_5__5798_, data_stage_5__5797_, data_stage_5__5796_, data_stage_5__5795_, data_stage_5__5794_, data_stage_5__5793_, data_stage_5__5792_, data_stage_5__5791_, data_stage_5__5790_, data_stage_5__5789_, data_stage_5__5788_, data_stage_5__5787_, data_stage_5__5786_, data_stage_5__5785_, data_stage_5__5784_, data_stage_5__5783_, data_stage_5__5782_, data_stage_5__5781_, data_stage_5__5780_, data_stage_5__5779_, data_stage_5__5778_, data_stage_5__5777_, data_stage_5__5776_, data_stage_5__5775_, data_stage_5__5774_, data_stage_5__5773_, data_stage_5__5772_, data_stage_5__5771_, data_stage_5__5770_, data_stage_5__5769_, data_stage_5__5768_, data_stage_5__5767_, data_stage_5__5766_, data_stage_5__5765_, data_stage_5__5764_, data_stage_5__5763_, data_stage_5__5762_, data_stage_5__5761_, data_stage_5__5760_, data_stage_5__5759_, data_stage_5__5758_, data_stage_5__5757_, data_stage_5__5756_, data_stage_5__5755_, data_stage_5__5754_, data_stage_5__5753_, data_stage_5__5752_, data_stage_5__5751_, data_stage_5__5750_, data_stage_5__5749_, data_stage_5__5748_, data_stage_5__5747_, data_stage_5__5746_, data_stage_5__5745_, data_stage_5__5744_, data_stage_5__5743_, data_stage_5__5742_, data_stage_5__5741_, data_stage_5__5740_, data_stage_5__5739_, data_stage_5__5738_, data_stage_5__5737_, data_stage_5__5736_, data_stage_5__5735_, data_stage_5__5734_, data_stage_5__5733_, data_stage_5__5732_, data_stage_5__5731_, data_stage_5__5730_, data_stage_5__5729_, data_stage_5__5728_, data_stage_5__5727_, data_stage_5__5726_, data_stage_5__5725_, data_stage_5__5724_, data_stage_5__5723_, data_stage_5__5722_, data_stage_5__5721_, data_stage_5__5720_, data_stage_5__5719_, data_stage_5__5718_, data_stage_5__5717_, data_stage_5__5716_, data_stage_5__5715_, data_stage_5__5714_, data_stage_5__5713_, data_stage_5__5712_, data_stage_5__5711_, data_stage_5__5710_, data_stage_5__5709_, data_stage_5__5708_, data_stage_5__5707_, data_stage_5__5706_, data_stage_5__5705_, data_stage_5__5704_, data_stage_5__5703_, data_stage_5__5702_, data_stage_5__5701_, data_stage_5__5700_, data_stage_5__5699_, data_stage_5__5698_, data_stage_5__5697_, data_stage_5__5696_, data_stage_5__5695_, data_stage_5__5694_, data_stage_5__5693_, data_stage_5__5692_, data_stage_5__5691_, data_stage_5__5690_, data_stage_5__5689_, data_stage_5__5688_, data_stage_5__5687_, data_stage_5__5686_, data_stage_5__5685_, data_stage_5__5684_, data_stage_5__5683_, data_stage_5__5682_, data_stage_5__5681_, data_stage_5__5680_, data_stage_5__5679_, data_stage_5__5678_, data_stage_5__5677_, data_stage_5__5676_, data_stage_5__5675_, data_stage_5__5674_, data_stage_5__5673_, data_stage_5__5672_, data_stage_5__5671_, data_stage_5__5670_, data_stage_5__5669_, data_stage_5__5668_, data_stage_5__5667_, data_stage_5__5666_, data_stage_5__5665_, data_stage_5__5664_, data_stage_5__5663_, data_stage_5__5662_, data_stage_5__5661_, data_stage_5__5660_, data_stage_5__5659_, data_stage_5__5658_, data_stage_5__5657_, data_stage_5__5656_, data_stage_5__5655_, data_stage_5__5654_, data_stage_5__5653_, data_stage_5__5652_, data_stage_5__5651_, data_stage_5__5650_, data_stage_5__5649_, data_stage_5__5648_, data_stage_5__5647_, data_stage_5__5646_, data_stage_5__5645_, data_stage_5__5644_, data_stage_5__5643_, data_stage_5__5642_, data_stage_5__5641_, data_stage_5__5640_, data_stage_5__5639_, data_stage_5__5638_, data_stage_5__5637_, data_stage_5__5636_, data_stage_5__5635_, data_stage_5__5634_, data_stage_5__5633_, data_stage_5__5632_, data_stage_5__5631_, data_stage_5__5630_, data_stage_5__5629_, data_stage_5__5628_, data_stage_5__5627_, data_stage_5__5626_, data_stage_5__5625_, data_stage_5__5624_, data_stage_5__5623_, data_stage_5__5622_, data_stage_5__5621_, data_stage_5__5620_, data_stage_5__5619_, data_stage_5__5618_, data_stage_5__5617_, data_stage_5__5616_, data_stage_5__5615_, data_stage_5__5614_, data_stage_5__5613_, data_stage_5__5612_, data_stage_5__5611_, data_stage_5__5610_, data_stage_5__5609_, data_stage_5__5608_, data_stage_5__5607_, data_stage_5__5606_, data_stage_5__5605_, data_stage_5__5604_, data_stage_5__5603_, data_stage_5__5602_, data_stage_5__5601_, data_stage_5__5600_, data_stage_5__5599_, data_stage_5__5598_, data_stage_5__5597_, data_stage_5__5596_, data_stage_5__5595_, data_stage_5__5594_, data_stage_5__5593_, data_stage_5__5592_, data_stage_5__5591_, data_stage_5__5590_, data_stage_5__5589_, data_stage_5__5588_, data_stage_5__5587_, data_stage_5__5586_, data_stage_5__5585_, data_stage_5__5584_, data_stage_5__5583_, data_stage_5__5582_, data_stage_5__5581_, data_stage_5__5580_, data_stage_5__5579_, data_stage_5__5578_, data_stage_5__5577_, data_stage_5__5576_, data_stage_5__5575_, data_stage_5__5574_, data_stage_5__5573_, data_stage_5__5572_, data_stage_5__5571_, data_stage_5__5570_, data_stage_5__5569_, data_stage_5__5568_, data_stage_5__5567_, data_stage_5__5566_, data_stage_5__5565_, data_stage_5__5564_, data_stage_5__5563_, data_stage_5__5562_, data_stage_5__5561_, data_stage_5__5560_, data_stage_5__5559_, data_stage_5__5558_, data_stage_5__5557_, data_stage_5__5556_, data_stage_5__5555_, data_stage_5__5554_, data_stage_5__5553_, data_stage_5__5552_, data_stage_5__5551_, data_stage_5__5550_, data_stage_5__5549_, data_stage_5__5548_, data_stage_5__5547_, data_stage_5__5546_, data_stage_5__5545_, data_stage_5__5544_, data_stage_5__5543_, data_stage_5__5542_, data_stage_5__5541_, data_stage_5__5540_, data_stage_5__5539_, data_stage_5__5538_, data_stage_5__5537_, data_stage_5__5536_, data_stage_5__5535_, data_stage_5__5534_, data_stage_5__5533_, data_stage_5__5532_, data_stage_5__5531_, data_stage_5__5530_, data_stage_5__5529_, data_stage_5__5528_, data_stage_5__5527_, data_stage_5__5526_, data_stage_5__5525_, data_stage_5__5524_, data_stage_5__5523_, data_stage_5__5522_, data_stage_5__5521_, data_stage_5__5520_, data_stage_5__5519_, data_stage_5__5518_, data_stage_5__5517_, data_stage_5__5516_, data_stage_5__5515_, data_stage_5__5514_, data_stage_5__5513_, data_stage_5__5512_, data_stage_5__5511_, data_stage_5__5510_, data_stage_5__5509_, data_stage_5__5508_, data_stage_5__5507_, data_stage_5__5506_, data_stage_5__5505_, data_stage_5__5504_, data_stage_5__5503_, data_stage_5__5502_, data_stage_5__5501_, data_stage_5__5500_, data_stage_5__5499_, data_stage_5__5498_, data_stage_5__5497_, data_stage_5__5496_, data_stage_5__5495_, data_stage_5__5494_, data_stage_5__5493_, data_stage_5__5492_, data_stage_5__5491_, data_stage_5__5490_, data_stage_5__5489_, data_stage_5__5488_, data_stage_5__5487_, data_stage_5__5486_, data_stage_5__5485_, data_stage_5__5484_, data_stage_5__5483_, data_stage_5__5482_, data_stage_5__5481_, data_stage_5__5480_, data_stage_5__5479_, data_stage_5__5478_, data_stage_5__5477_, data_stage_5__5476_, data_stage_5__5475_, data_stage_5__5474_, data_stage_5__5473_, data_stage_5__5472_, data_stage_5__5471_, data_stage_5__5470_, data_stage_5__5469_, data_stage_5__5468_, data_stage_5__5467_, data_stage_5__5466_, data_stage_5__5465_, data_stage_5__5464_, data_stage_5__5463_, data_stage_5__5462_, data_stage_5__5461_, data_stage_5__5460_, data_stage_5__5459_, data_stage_5__5458_, data_stage_5__5457_, data_stage_5__5456_, data_stage_5__5455_, data_stage_5__5454_, data_stage_5__5453_, data_stage_5__5452_, data_stage_5__5451_, data_stage_5__5450_, data_stage_5__5449_, data_stage_5__5448_, data_stage_5__5447_, data_stage_5__5446_, data_stage_5__5445_, data_stage_5__5444_, data_stage_5__5443_, data_stage_5__5442_, data_stage_5__5441_, data_stage_5__5440_, data_stage_5__5439_, data_stage_5__5438_, data_stage_5__5437_, data_stage_5__5436_, data_stage_5__5435_, data_stage_5__5434_, data_stage_5__5433_, data_stage_5__5432_, data_stage_5__5431_, data_stage_5__5430_, data_stage_5__5429_, data_stage_5__5428_, data_stage_5__5427_, data_stage_5__5426_, data_stage_5__5425_, data_stage_5__5424_, data_stage_5__5423_, data_stage_5__5422_, data_stage_5__5421_, data_stage_5__5420_, data_stage_5__5419_, data_stage_5__5418_, data_stage_5__5417_, data_stage_5__5416_, data_stage_5__5415_, data_stage_5__5414_, data_stage_5__5413_, data_stage_5__5412_, data_stage_5__5411_, data_stage_5__5410_, data_stage_5__5409_, data_stage_5__5408_, data_stage_5__5407_, data_stage_5__5406_, data_stage_5__5405_, data_stage_5__5404_, data_stage_5__5403_, data_stage_5__5402_, data_stage_5__5401_, data_stage_5__5400_, data_stage_5__5399_, data_stage_5__5398_, data_stage_5__5397_, data_stage_5__5396_, data_stage_5__5395_, data_stage_5__5394_, data_stage_5__5393_, data_stage_5__5392_, data_stage_5__5391_, data_stage_5__5390_, data_stage_5__5389_, data_stage_5__5388_, data_stage_5__5387_, data_stage_5__5386_, data_stage_5__5385_, data_stage_5__5384_, data_stage_5__5383_, data_stage_5__5382_, data_stage_5__5381_, data_stage_5__5380_, data_stage_5__5379_, data_stage_5__5378_, data_stage_5__5377_, data_stage_5__5376_, data_stage_5__5375_, data_stage_5__5374_, data_stage_5__5373_, data_stage_5__5372_, data_stage_5__5371_, data_stage_5__5370_, data_stage_5__5369_, data_stage_5__5368_, data_stage_5__5367_, data_stage_5__5366_, data_stage_5__5365_, data_stage_5__5364_, data_stage_5__5363_, data_stage_5__5362_, data_stage_5__5361_, data_stage_5__5360_, data_stage_5__5359_, data_stage_5__5358_, data_stage_5__5357_, data_stage_5__5356_, data_stage_5__5355_, data_stage_5__5354_, data_stage_5__5353_, data_stage_5__5352_, data_stage_5__5351_, data_stage_5__5350_, data_stage_5__5349_, data_stage_5__5348_, data_stage_5__5347_, data_stage_5__5346_, data_stage_5__5345_, data_stage_5__5344_, data_stage_5__5343_, data_stage_5__5342_, data_stage_5__5341_, data_stage_5__5340_, data_stage_5__5339_, data_stage_5__5338_, data_stage_5__5337_, data_stage_5__5336_, data_stage_5__5335_, data_stage_5__5334_, data_stage_5__5333_, data_stage_5__5332_, data_stage_5__5331_, data_stage_5__5330_, data_stage_5__5329_, data_stage_5__5328_, data_stage_5__5327_, data_stage_5__5326_, data_stage_5__5325_, data_stage_5__5324_, data_stage_5__5323_, data_stage_5__5322_, data_stage_5__5321_, data_stage_5__5320_, data_stage_5__5319_, data_stage_5__5318_, data_stage_5__5317_, data_stage_5__5316_, data_stage_5__5315_, data_stage_5__5314_, data_stage_5__5313_, data_stage_5__5312_, data_stage_5__5311_, data_stage_5__5310_, data_stage_5__5309_, data_stage_5__5308_, data_stage_5__5307_, data_stage_5__5306_, data_stage_5__5305_, data_stage_5__5304_, data_stage_5__5303_, data_stage_5__5302_, data_stage_5__5301_, data_stage_5__5300_, data_stage_5__5299_, data_stage_5__5298_, data_stage_5__5297_, data_stage_5__5296_, data_stage_5__5295_, data_stage_5__5294_, data_stage_5__5293_, data_stage_5__5292_, data_stage_5__5291_, data_stage_5__5290_, data_stage_5__5289_, data_stage_5__5288_, data_stage_5__5287_, data_stage_5__5286_, data_stage_5__5285_, data_stage_5__5284_, data_stage_5__5283_, data_stage_5__5282_, data_stage_5__5281_, data_stage_5__5280_, data_stage_5__5279_, data_stage_5__5278_, data_stage_5__5277_, data_stage_5__5276_, data_stage_5__5275_, data_stage_5__5274_, data_stage_5__5273_, data_stage_5__5272_, data_stage_5__5271_, data_stage_5__5270_, data_stage_5__5269_, data_stage_5__5268_, data_stage_5__5267_, data_stage_5__5266_, data_stage_5__5265_, data_stage_5__5264_, data_stage_5__5263_, data_stage_5__5262_, data_stage_5__5261_, data_stage_5__5260_, data_stage_5__5259_, data_stage_5__5258_, data_stage_5__5257_, data_stage_5__5256_, data_stage_5__5255_, data_stage_5__5254_, data_stage_5__5253_, data_stage_5__5252_, data_stage_5__5251_, data_stage_5__5250_, data_stage_5__5249_, data_stage_5__5248_, data_stage_5__5247_, data_stage_5__5246_, data_stage_5__5245_, data_stage_5__5244_, data_stage_5__5243_, data_stage_5__5242_, data_stage_5__5241_, data_stage_5__5240_, data_stage_5__5239_, data_stage_5__5238_, data_stage_5__5237_, data_stage_5__5236_, data_stage_5__5235_, data_stage_5__5234_, data_stage_5__5233_, data_stage_5__5232_, data_stage_5__5231_, data_stage_5__5230_, data_stage_5__5229_, data_stage_5__5228_, data_stage_5__5227_, data_stage_5__5226_, data_stage_5__5225_, data_stage_5__5224_, data_stage_5__5223_, data_stage_5__5222_, data_stage_5__5221_, data_stage_5__5220_, data_stage_5__5219_, data_stage_5__5218_, data_stage_5__5217_, data_stage_5__5216_, data_stage_5__5215_, data_stage_5__5214_, data_stage_5__5213_, data_stage_5__5212_, data_stage_5__5211_, data_stage_5__5210_, data_stage_5__5209_, data_stage_5__5208_, data_stage_5__5207_, data_stage_5__5206_, data_stage_5__5205_, data_stage_5__5204_, data_stage_5__5203_, data_stage_5__5202_, data_stage_5__5201_, data_stage_5__5200_, data_stage_5__5199_, data_stage_5__5198_, data_stage_5__5197_, data_stage_5__5196_, data_stage_5__5195_, data_stage_5__5194_, data_stage_5__5193_, data_stage_5__5192_, data_stage_5__5191_, data_stage_5__5190_, data_stage_5__5189_, data_stage_5__5188_, data_stage_5__5187_, data_stage_5__5186_, data_stage_5__5185_, data_stage_5__5184_, data_stage_5__5183_, data_stage_5__5182_, data_stage_5__5181_, data_stage_5__5180_, data_stage_5__5179_, data_stage_5__5178_, data_stage_5__5177_, data_stage_5__5176_, data_stage_5__5175_, data_stage_5__5174_, data_stage_5__5173_, data_stage_5__5172_, data_stage_5__5171_, data_stage_5__5170_, data_stage_5__5169_, data_stage_5__5168_, data_stage_5__5167_, data_stage_5__5166_, data_stage_5__5165_, data_stage_5__5164_, data_stage_5__5163_, data_stage_5__5162_, data_stage_5__5161_, data_stage_5__5160_, data_stage_5__5159_, data_stage_5__5158_, data_stage_5__5157_, data_stage_5__5156_, data_stage_5__5155_, data_stage_5__5154_, data_stage_5__5153_, data_stage_5__5152_, data_stage_5__5151_, data_stage_5__5150_, data_stage_5__5149_, data_stage_5__5148_, data_stage_5__5147_, data_stage_5__5146_, data_stage_5__5145_, data_stage_5__5144_, data_stage_5__5143_, data_stage_5__5142_, data_stage_5__5141_, data_stage_5__5140_, data_stage_5__5139_, data_stage_5__5138_, data_stage_5__5137_, data_stage_5__5136_, data_stage_5__5135_, data_stage_5__5134_, data_stage_5__5133_, data_stage_5__5132_, data_stage_5__5131_, data_stage_5__5130_, data_stage_5__5129_, data_stage_5__5128_, data_stage_5__5127_, data_stage_5__5126_, data_stage_5__5125_, data_stage_5__5124_, data_stage_5__5123_, data_stage_5__5122_, data_stage_5__5121_, data_stage_5__5120_, data_stage_5__5119_, data_stage_5__5118_, data_stage_5__5117_, data_stage_5__5116_, data_stage_5__5115_, data_stage_5__5114_, data_stage_5__5113_, data_stage_5__5112_, data_stage_5__5111_, data_stage_5__5110_, data_stage_5__5109_, data_stage_5__5108_, data_stage_5__5107_, data_stage_5__5106_, data_stage_5__5105_, data_stage_5__5104_, data_stage_5__5103_, data_stage_5__5102_, data_stage_5__5101_, data_stage_5__5100_, data_stage_5__5099_, data_stage_5__5098_, data_stage_5__5097_, data_stage_5__5096_, data_stage_5__5095_, data_stage_5__5094_, data_stage_5__5093_, data_stage_5__5092_, data_stage_5__5091_, data_stage_5__5090_, data_stage_5__5089_, data_stage_5__5088_, data_stage_5__5087_, data_stage_5__5086_, data_stage_5__5085_, data_stage_5__5084_, data_stage_5__5083_, data_stage_5__5082_, data_stage_5__5081_, data_stage_5__5080_, data_stage_5__5079_, data_stage_5__5078_, data_stage_5__5077_, data_stage_5__5076_, data_stage_5__5075_, data_stage_5__5074_, data_stage_5__5073_, data_stage_5__5072_, data_stage_5__5071_, data_stage_5__5070_, data_stage_5__5069_, data_stage_5__5068_, data_stage_5__5067_, data_stage_5__5066_, data_stage_5__5065_, data_stage_5__5064_, data_stage_5__5063_, data_stage_5__5062_, data_stage_5__5061_, data_stage_5__5060_, data_stage_5__5059_, data_stage_5__5058_, data_stage_5__5057_, data_stage_5__5056_, data_stage_5__5055_, data_stage_5__5054_, data_stage_5__5053_, data_stage_5__5052_, data_stage_5__5051_, data_stage_5__5050_, data_stage_5__5049_, data_stage_5__5048_, data_stage_5__5047_, data_stage_5__5046_, data_stage_5__5045_, data_stage_5__5044_, data_stage_5__5043_, data_stage_5__5042_, data_stage_5__5041_, data_stage_5__5040_, data_stage_5__5039_, data_stage_5__5038_, data_stage_5__5037_, data_stage_5__5036_, data_stage_5__5035_, data_stage_5__5034_, data_stage_5__5033_, data_stage_5__5032_, data_stage_5__5031_, data_stage_5__5030_, data_stage_5__5029_, data_stage_5__5028_, data_stage_5__5027_, data_stage_5__5026_, data_stage_5__5025_, data_stage_5__5024_, data_stage_5__5023_, data_stage_5__5022_, data_stage_5__5021_, data_stage_5__5020_, data_stage_5__5019_, data_stage_5__5018_, data_stage_5__5017_, data_stage_5__5016_, data_stage_5__5015_, data_stage_5__5014_, data_stage_5__5013_, data_stage_5__5012_, data_stage_5__5011_, data_stage_5__5010_, data_stage_5__5009_, data_stage_5__5008_, data_stage_5__5007_, data_stage_5__5006_, data_stage_5__5005_, data_stage_5__5004_, data_stage_5__5003_, data_stage_5__5002_, data_stage_5__5001_, data_stage_5__5000_, data_stage_5__4999_, data_stage_5__4998_, data_stage_5__4997_, data_stage_5__4996_, data_stage_5__4995_, data_stage_5__4994_, data_stage_5__4993_, data_stage_5__4992_, data_stage_5__4991_, data_stage_5__4990_, data_stage_5__4989_, data_stage_5__4988_, data_stage_5__4987_, data_stage_5__4986_, data_stage_5__4985_, data_stage_5__4984_, data_stage_5__4983_, data_stage_5__4982_, data_stage_5__4981_, data_stage_5__4980_, data_stage_5__4979_, data_stage_5__4978_, data_stage_5__4977_, data_stage_5__4976_, data_stage_5__4975_, data_stage_5__4974_, data_stage_5__4973_, data_stage_5__4972_, data_stage_5__4971_, data_stage_5__4970_, data_stage_5__4969_, data_stage_5__4968_, data_stage_5__4967_, data_stage_5__4966_, data_stage_5__4965_, data_stage_5__4964_, data_stage_5__4963_, data_stage_5__4962_, data_stage_5__4961_, data_stage_5__4960_, data_stage_5__4959_, data_stage_5__4958_, data_stage_5__4957_, data_stage_5__4956_, data_stage_5__4955_, data_stage_5__4954_, data_stage_5__4953_, data_stage_5__4952_, data_stage_5__4951_, data_stage_5__4950_, data_stage_5__4949_, data_stage_5__4948_, data_stage_5__4947_, data_stage_5__4946_, data_stage_5__4945_, data_stage_5__4944_, data_stage_5__4943_, data_stage_5__4942_, data_stage_5__4941_, data_stage_5__4940_, data_stage_5__4939_, data_stage_5__4938_, data_stage_5__4937_, data_stage_5__4936_, data_stage_5__4935_, data_stage_5__4934_, data_stage_5__4933_, data_stage_5__4932_, data_stage_5__4931_, data_stage_5__4930_, data_stage_5__4929_, data_stage_5__4928_, data_stage_5__4927_, data_stage_5__4926_, data_stage_5__4925_, data_stage_5__4924_, data_stage_5__4923_, data_stage_5__4922_, data_stage_5__4921_, data_stage_5__4920_, data_stage_5__4919_, data_stage_5__4918_, data_stage_5__4917_, data_stage_5__4916_, data_stage_5__4915_, data_stage_5__4914_, data_stage_5__4913_, data_stage_5__4912_, data_stage_5__4911_, data_stage_5__4910_, data_stage_5__4909_, data_stage_5__4908_, data_stage_5__4907_, data_stage_5__4906_, data_stage_5__4905_, data_stage_5__4904_, data_stage_5__4903_, data_stage_5__4902_, data_stage_5__4901_, data_stage_5__4900_, data_stage_5__4899_, data_stage_5__4898_, data_stage_5__4897_, data_stage_5__4896_, data_stage_5__4895_, data_stage_5__4894_, data_stage_5__4893_, data_stage_5__4892_, data_stage_5__4891_, data_stage_5__4890_, data_stage_5__4889_, data_stage_5__4888_, data_stage_5__4887_, data_stage_5__4886_, data_stage_5__4885_, data_stage_5__4884_, data_stage_5__4883_, data_stage_5__4882_, data_stage_5__4881_, data_stage_5__4880_, data_stage_5__4879_, data_stage_5__4878_, data_stage_5__4877_, data_stage_5__4876_, data_stage_5__4875_, data_stage_5__4874_, data_stage_5__4873_, data_stage_5__4872_, data_stage_5__4871_, data_stage_5__4870_, data_stage_5__4869_, data_stage_5__4868_, data_stage_5__4867_, data_stage_5__4866_, data_stage_5__4865_, data_stage_5__4864_, data_stage_5__4863_, data_stage_5__4862_, data_stage_5__4861_, data_stage_5__4860_, data_stage_5__4859_, data_stage_5__4858_, data_stage_5__4857_, data_stage_5__4856_, data_stage_5__4855_, data_stage_5__4854_, data_stage_5__4853_, data_stage_5__4852_, data_stage_5__4851_, data_stage_5__4850_, data_stage_5__4849_, data_stage_5__4848_, data_stage_5__4847_, data_stage_5__4846_, data_stage_5__4845_, data_stage_5__4844_, data_stage_5__4843_, data_stage_5__4842_, data_stage_5__4841_, data_stage_5__4840_, data_stage_5__4839_, data_stage_5__4838_, data_stage_5__4837_, data_stage_5__4836_, data_stage_5__4835_, data_stage_5__4834_, data_stage_5__4833_, data_stage_5__4832_, data_stage_5__4831_, data_stage_5__4830_, data_stage_5__4829_, data_stage_5__4828_, data_stage_5__4827_, data_stage_5__4826_, data_stage_5__4825_, data_stage_5__4824_, data_stage_5__4823_, data_stage_5__4822_, data_stage_5__4821_, data_stage_5__4820_, data_stage_5__4819_, data_stage_5__4818_, data_stage_5__4817_, data_stage_5__4816_, data_stage_5__4815_, data_stage_5__4814_, data_stage_5__4813_, data_stage_5__4812_, data_stage_5__4811_, data_stage_5__4810_, data_stage_5__4809_, data_stage_5__4808_, data_stage_5__4807_, data_stage_5__4806_, data_stage_5__4805_, data_stage_5__4804_, data_stage_5__4803_, data_stage_5__4802_, data_stage_5__4801_, data_stage_5__4800_, data_stage_5__4799_, data_stage_5__4798_, data_stage_5__4797_, data_stage_5__4796_, data_stage_5__4795_, data_stage_5__4794_, data_stage_5__4793_, data_stage_5__4792_, data_stage_5__4791_, data_stage_5__4790_, data_stage_5__4789_, data_stage_5__4788_, data_stage_5__4787_, data_stage_5__4786_, data_stage_5__4785_, data_stage_5__4784_, data_stage_5__4783_, data_stage_5__4782_, data_stage_5__4781_, data_stage_5__4780_, data_stage_5__4779_, data_stage_5__4778_, data_stage_5__4777_, data_stage_5__4776_, data_stage_5__4775_, data_stage_5__4774_, data_stage_5__4773_, data_stage_5__4772_, data_stage_5__4771_, data_stage_5__4770_, data_stage_5__4769_, data_stage_5__4768_, data_stage_5__4767_, data_stage_5__4766_, data_stage_5__4765_, data_stage_5__4764_, data_stage_5__4763_, data_stage_5__4762_, data_stage_5__4761_, data_stage_5__4760_, data_stage_5__4759_, data_stage_5__4758_, data_stage_5__4757_, data_stage_5__4756_, data_stage_5__4755_, data_stage_5__4754_, data_stage_5__4753_, data_stage_5__4752_, data_stage_5__4751_, data_stage_5__4750_, data_stage_5__4749_, data_stage_5__4748_, data_stage_5__4747_, data_stage_5__4746_, data_stage_5__4745_, data_stage_5__4744_, data_stage_5__4743_, data_stage_5__4742_, data_stage_5__4741_, data_stage_5__4740_, data_stage_5__4739_, data_stage_5__4738_, data_stage_5__4737_, data_stage_5__4736_, data_stage_5__4735_, data_stage_5__4734_, data_stage_5__4733_, data_stage_5__4732_, data_stage_5__4731_, data_stage_5__4730_, data_stage_5__4729_, data_stage_5__4728_, data_stage_5__4727_, data_stage_5__4726_, data_stage_5__4725_, data_stage_5__4724_, data_stage_5__4723_, data_stage_5__4722_, data_stage_5__4721_, data_stage_5__4720_, data_stage_5__4719_, data_stage_5__4718_, data_stage_5__4717_, data_stage_5__4716_, data_stage_5__4715_, data_stage_5__4714_, data_stage_5__4713_, data_stage_5__4712_, data_stage_5__4711_, data_stage_5__4710_, data_stage_5__4709_, data_stage_5__4708_, data_stage_5__4707_, data_stage_5__4706_, data_stage_5__4705_, data_stage_5__4704_, data_stage_5__4703_, data_stage_5__4702_, data_stage_5__4701_, data_stage_5__4700_, data_stage_5__4699_, data_stage_5__4698_, data_stage_5__4697_, data_stage_5__4696_, data_stage_5__4695_, data_stage_5__4694_, data_stage_5__4693_, data_stage_5__4692_, data_stage_5__4691_, data_stage_5__4690_, data_stage_5__4689_, data_stage_5__4688_, data_stage_5__4687_, data_stage_5__4686_, data_stage_5__4685_, data_stage_5__4684_, data_stage_5__4683_, data_stage_5__4682_, data_stage_5__4681_, data_stage_5__4680_, data_stage_5__4679_, data_stage_5__4678_, data_stage_5__4677_, data_stage_5__4676_, data_stage_5__4675_, data_stage_5__4674_, data_stage_5__4673_, data_stage_5__4672_, data_stage_5__4671_, data_stage_5__4670_, data_stage_5__4669_, data_stage_5__4668_, data_stage_5__4667_, data_stage_5__4666_, data_stage_5__4665_, data_stage_5__4664_, data_stage_5__4663_, data_stage_5__4662_, data_stage_5__4661_, data_stage_5__4660_, data_stage_5__4659_, data_stage_5__4658_, data_stage_5__4657_, data_stage_5__4656_, data_stage_5__4655_, data_stage_5__4654_, data_stage_5__4653_, data_stage_5__4652_, data_stage_5__4651_, data_stage_5__4650_, data_stage_5__4649_, data_stage_5__4648_, data_stage_5__4647_, data_stage_5__4646_, data_stage_5__4645_, data_stage_5__4644_, data_stage_5__4643_, data_stage_5__4642_, data_stage_5__4641_, data_stage_5__4640_, data_stage_5__4639_, data_stage_5__4638_, data_stage_5__4637_, data_stage_5__4636_, data_stage_5__4635_, data_stage_5__4634_, data_stage_5__4633_, data_stage_5__4632_, data_stage_5__4631_, data_stage_5__4630_, data_stage_5__4629_, data_stage_5__4628_, data_stage_5__4627_, data_stage_5__4626_, data_stage_5__4625_, data_stage_5__4624_, data_stage_5__4623_, data_stage_5__4622_, data_stage_5__4621_, data_stage_5__4620_, data_stage_5__4619_, data_stage_5__4618_, data_stage_5__4617_, data_stage_5__4616_, data_stage_5__4615_, data_stage_5__4614_, data_stage_5__4613_, data_stage_5__4612_, data_stage_5__4611_, data_stage_5__4610_, data_stage_5__4609_, data_stage_5__4608_, data_stage_5__4607_, data_stage_5__4606_, data_stage_5__4605_, data_stage_5__4604_, data_stage_5__4603_, data_stage_5__4602_, data_stage_5__4601_, data_stage_5__4600_, data_stage_5__4599_, data_stage_5__4598_, data_stage_5__4597_, data_stage_5__4596_, data_stage_5__4595_, data_stage_5__4594_, data_stage_5__4593_, data_stage_5__4592_, data_stage_5__4591_, data_stage_5__4590_, data_stage_5__4589_, data_stage_5__4588_, data_stage_5__4587_, data_stage_5__4586_, data_stage_5__4585_, data_stage_5__4584_, data_stage_5__4583_, data_stage_5__4582_, data_stage_5__4581_, data_stage_5__4580_, data_stage_5__4579_, data_stage_5__4578_, data_stage_5__4577_, data_stage_5__4576_, data_stage_5__4575_, data_stage_5__4574_, data_stage_5__4573_, data_stage_5__4572_, data_stage_5__4571_, data_stage_5__4570_, data_stage_5__4569_, data_stage_5__4568_, data_stage_5__4567_, data_stage_5__4566_, data_stage_5__4565_, data_stage_5__4564_, data_stage_5__4563_, data_stage_5__4562_, data_stage_5__4561_, data_stage_5__4560_, data_stage_5__4559_, data_stage_5__4558_, data_stage_5__4557_, data_stage_5__4556_, data_stage_5__4555_, data_stage_5__4554_, data_stage_5__4553_, data_stage_5__4552_, data_stage_5__4551_, data_stage_5__4550_, data_stage_5__4549_, data_stage_5__4548_, data_stage_5__4547_, data_stage_5__4546_, data_stage_5__4545_, data_stage_5__4544_, data_stage_5__4543_, data_stage_5__4542_, data_stage_5__4541_, data_stage_5__4540_, data_stage_5__4539_, data_stage_5__4538_, data_stage_5__4537_, data_stage_5__4536_, data_stage_5__4535_, data_stage_5__4534_, data_stage_5__4533_, data_stage_5__4532_, data_stage_5__4531_, data_stage_5__4530_, data_stage_5__4529_, data_stage_5__4528_, data_stage_5__4527_, data_stage_5__4526_, data_stage_5__4525_, data_stage_5__4524_, data_stage_5__4523_, data_stage_5__4522_, data_stage_5__4521_, data_stage_5__4520_, data_stage_5__4519_, data_stage_5__4518_, data_stage_5__4517_, data_stage_5__4516_, data_stage_5__4515_, data_stage_5__4514_, data_stage_5__4513_, data_stage_5__4512_, data_stage_5__4511_, data_stage_5__4510_, data_stage_5__4509_, data_stage_5__4508_, data_stage_5__4507_, data_stage_5__4506_, data_stage_5__4505_, data_stage_5__4504_, data_stage_5__4503_, data_stage_5__4502_, data_stage_5__4501_, data_stage_5__4500_, data_stage_5__4499_, data_stage_5__4498_, data_stage_5__4497_, data_stage_5__4496_, data_stage_5__4495_, data_stage_5__4494_, data_stage_5__4493_, data_stage_5__4492_, data_stage_5__4491_, data_stage_5__4490_, data_stage_5__4489_, data_stage_5__4488_, data_stage_5__4487_, data_stage_5__4486_, data_stage_5__4485_, data_stage_5__4484_, data_stage_5__4483_, data_stage_5__4482_, data_stage_5__4481_, data_stage_5__4480_, data_stage_5__4479_, data_stage_5__4478_, data_stage_5__4477_, data_stage_5__4476_, data_stage_5__4475_, data_stage_5__4474_, data_stage_5__4473_, data_stage_5__4472_, data_stage_5__4471_, data_stage_5__4470_, data_stage_5__4469_, data_stage_5__4468_, data_stage_5__4467_, data_stage_5__4466_, data_stage_5__4465_, data_stage_5__4464_, data_stage_5__4463_, data_stage_5__4462_, data_stage_5__4461_, data_stage_5__4460_, data_stage_5__4459_, data_stage_5__4458_, data_stage_5__4457_, data_stage_5__4456_, data_stage_5__4455_, data_stage_5__4454_, data_stage_5__4453_, data_stage_5__4452_, data_stage_5__4451_, data_stage_5__4450_, data_stage_5__4449_, data_stage_5__4448_, data_stage_5__4447_, data_stage_5__4446_, data_stage_5__4445_, data_stage_5__4444_, data_stage_5__4443_, data_stage_5__4442_, data_stage_5__4441_, data_stage_5__4440_, data_stage_5__4439_, data_stage_5__4438_, data_stage_5__4437_, data_stage_5__4436_, data_stage_5__4435_, data_stage_5__4434_, data_stage_5__4433_, data_stage_5__4432_, data_stage_5__4431_, data_stage_5__4430_, data_stage_5__4429_, data_stage_5__4428_, data_stage_5__4427_, data_stage_5__4426_, data_stage_5__4425_, data_stage_5__4424_, data_stage_5__4423_, data_stage_5__4422_, data_stage_5__4421_, data_stage_5__4420_, data_stage_5__4419_, data_stage_5__4418_, data_stage_5__4417_, data_stage_5__4416_, data_stage_5__4415_, data_stage_5__4414_, data_stage_5__4413_, data_stage_5__4412_, data_stage_5__4411_, data_stage_5__4410_, data_stage_5__4409_, data_stage_5__4408_, data_stage_5__4407_, data_stage_5__4406_, data_stage_5__4405_, data_stage_5__4404_, data_stage_5__4403_, data_stage_5__4402_, data_stage_5__4401_, data_stage_5__4400_, data_stage_5__4399_, data_stage_5__4398_, data_stage_5__4397_, data_stage_5__4396_, data_stage_5__4395_, data_stage_5__4394_, data_stage_5__4393_, data_stage_5__4392_, data_stage_5__4391_, data_stage_5__4390_, data_stage_5__4389_, data_stage_5__4388_, data_stage_5__4387_, data_stage_5__4386_, data_stage_5__4385_, data_stage_5__4384_, data_stage_5__4383_, data_stage_5__4382_, data_stage_5__4381_, data_stage_5__4380_, data_stage_5__4379_, data_stage_5__4378_, data_stage_5__4377_, data_stage_5__4376_, data_stage_5__4375_, data_stage_5__4374_, data_stage_5__4373_, data_stage_5__4372_, data_stage_5__4371_, data_stage_5__4370_, data_stage_5__4369_, data_stage_5__4368_, data_stage_5__4367_, data_stage_5__4366_, data_stage_5__4365_, data_stage_5__4364_, data_stage_5__4363_, data_stage_5__4362_, data_stage_5__4361_, data_stage_5__4360_, data_stage_5__4359_, data_stage_5__4358_, data_stage_5__4357_, data_stage_5__4356_, data_stage_5__4355_, data_stage_5__4354_, data_stage_5__4353_, data_stage_5__4352_, data_stage_5__4351_, data_stage_5__4350_, data_stage_5__4349_, data_stage_5__4348_, data_stage_5__4347_, data_stage_5__4346_, data_stage_5__4345_, data_stage_5__4344_, data_stage_5__4343_, data_stage_5__4342_, data_stage_5__4341_, data_stage_5__4340_, data_stage_5__4339_, data_stage_5__4338_, data_stage_5__4337_, data_stage_5__4336_, data_stage_5__4335_, data_stage_5__4334_, data_stage_5__4333_, data_stage_5__4332_, data_stage_5__4331_, data_stage_5__4330_, data_stage_5__4329_, data_stage_5__4328_, data_stage_5__4327_, data_stage_5__4326_, data_stage_5__4325_, data_stage_5__4324_, data_stage_5__4323_, data_stage_5__4322_, data_stage_5__4321_, data_stage_5__4320_, data_stage_5__4319_, data_stage_5__4318_, data_stage_5__4317_, data_stage_5__4316_, data_stage_5__4315_, data_stage_5__4314_, data_stage_5__4313_, data_stage_5__4312_, data_stage_5__4311_, data_stage_5__4310_, data_stage_5__4309_, data_stage_5__4308_, data_stage_5__4307_, data_stage_5__4306_, data_stage_5__4305_, data_stage_5__4304_, data_stage_5__4303_, data_stage_5__4302_, data_stage_5__4301_, data_stage_5__4300_, data_stage_5__4299_, data_stage_5__4298_, data_stage_5__4297_, data_stage_5__4296_, data_stage_5__4295_, data_stage_5__4294_, data_stage_5__4293_, data_stage_5__4292_, data_stage_5__4291_, data_stage_5__4290_, data_stage_5__4289_, data_stage_5__4288_, data_stage_5__4287_, data_stage_5__4286_, data_stage_5__4285_, data_stage_5__4284_, data_stage_5__4283_, data_stage_5__4282_, data_stage_5__4281_, data_stage_5__4280_, data_stage_5__4279_, data_stage_5__4278_, data_stage_5__4277_, data_stage_5__4276_, data_stage_5__4275_, data_stage_5__4274_, data_stage_5__4273_, data_stage_5__4272_, data_stage_5__4271_, data_stage_5__4270_, data_stage_5__4269_, data_stage_5__4268_, data_stage_5__4267_, data_stage_5__4266_, data_stage_5__4265_, data_stage_5__4264_, data_stage_5__4263_, data_stage_5__4262_, data_stage_5__4261_, data_stage_5__4260_, data_stage_5__4259_, data_stage_5__4258_, data_stage_5__4257_, data_stage_5__4256_, data_stage_5__4255_, data_stage_5__4254_, data_stage_5__4253_, data_stage_5__4252_, data_stage_5__4251_, data_stage_5__4250_, data_stage_5__4249_, data_stage_5__4248_, data_stage_5__4247_, data_stage_5__4246_, data_stage_5__4245_, data_stage_5__4244_, data_stage_5__4243_, data_stage_5__4242_, data_stage_5__4241_, data_stage_5__4240_, data_stage_5__4239_, data_stage_5__4238_, data_stage_5__4237_, data_stage_5__4236_, data_stage_5__4235_, data_stage_5__4234_, data_stage_5__4233_, data_stage_5__4232_, data_stage_5__4231_, data_stage_5__4230_, data_stage_5__4229_, data_stage_5__4228_, data_stage_5__4227_, data_stage_5__4226_, data_stage_5__4225_, data_stage_5__4224_, data_stage_5__4223_, data_stage_5__4222_, data_stage_5__4221_, data_stage_5__4220_, data_stage_5__4219_, data_stage_5__4218_, data_stage_5__4217_, data_stage_5__4216_, data_stage_5__4215_, data_stage_5__4214_, data_stage_5__4213_, data_stage_5__4212_, data_stage_5__4211_, data_stage_5__4210_, data_stage_5__4209_, data_stage_5__4208_, data_stage_5__4207_, data_stage_5__4206_, data_stage_5__4205_, data_stage_5__4204_, data_stage_5__4203_, data_stage_5__4202_, data_stage_5__4201_, data_stage_5__4200_, data_stage_5__4199_, data_stage_5__4198_, data_stage_5__4197_, data_stage_5__4196_, data_stage_5__4195_, data_stage_5__4194_, data_stage_5__4193_, data_stage_5__4192_, data_stage_5__4191_, data_stage_5__4190_, data_stage_5__4189_, data_stage_5__4188_, data_stage_5__4187_, data_stage_5__4186_, data_stage_5__4185_, data_stage_5__4184_, data_stage_5__4183_, data_stage_5__4182_, data_stage_5__4181_, data_stage_5__4180_, data_stage_5__4179_, data_stage_5__4178_, data_stage_5__4177_, data_stage_5__4176_, data_stage_5__4175_, data_stage_5__4174_, data_stage_5__4173_, data_stage_5__4172_, data_stage_5__4171_, data_stage_5__4170_, data_stage_5__4169_, data_stage_5__4168_, data_stage_5__4167_, data_stage_5__4166_, data_stage_5__4165_, data_stage_5__4164_, data_stage_5__4163_, data_stage_5__4162_, data_stage_5__4161_, data_stage_5__4160_, data_stage_5__4159_, data_stage_5__4158_, data_stage_5__4157_, data_stage_5__4156_, data_stage_5__4155_, data_stage_5__4154_, data_stage_5__4153_, data_stage_5__4152_, data_stage_5__4151_, data_stage_5__4150_, data_stage_5__4149_, data_stage_5__4148_, data_stage_5__4147_, data_stage_5__4146_, data_stage_5__4145_, data_stage_5__4144_, data_stage_5__4143_, data_stage_5__4142_, data_stage_5__4141_, data_stage_5__4140_, data_stage_5__4139_, data_stage_5__4138_, data_stage_5__4137_, data_stage_5__4136_, data_stage_5__4135_, data_stage_5__4134_, data_stage_5__4133_, data_stage_5__4132_, data_stage_5__4131_, data_stage_5__4130_, data_stage_5__4129_, data_stage_5__4128_, data_stage_5__4127_, data_stage_5__4126_, data_stage_5__4125_, data_stage_5__4124_, data_stage_5__4123_, data_stage_5__4122_, data_stage_5__4121_, data_stage_5__4120_, data_stage_5__4119_, data_stage_5__4118_, data_stage_5__4117_, data_stage_5__4116_, data_stage_5__4115_, data_stage_5__4114_, data_stage_5__4113_, data_stage_5__4112_, data_stage_5__4111_, data_stage_5__4110_, data_stage_5__4109_, data_stage_5__4108_, data_stage_5__4107_, data_stage_5__4106_, data_stage_5__4105_, data_stage_5__4104_, data_stage_5__4103_, data_stage_5__4102_, data_stage_5__4101_, data_stage_5__4100_, data_stage_5__4099_, data_stage_5__4098_, data_stage_5__4097_, data_stage_5__4096_, data_stage_5__4095_, data_stage_5__4094_, data_stage_5__4093_, data_stage_5__4092_, data_stage_5__4091_, data_stage_5__4090_, data_stage_5__4089_, data_stage_5__4088_, data_stage_5__4087_, data_stage_5__4086_, data_stage_5__4085_, data_stage_5__4084_, data_stage_5__4083_, data_stage_5__4082_, data_stage_5__4081_, data_stage_5__4080_, data_stage_5__4079_, data_stage_5__4078_, data_stage_5__4077_, data_stage_5__4076_, data_stage_5__4075_, data_stage_5__4074_, data_stage_5__4073_, data_stage_5__4072_, data_stage_5__4071_, data_stage_5__4070_, data_stage_5__4069_, data_stage_5__4068_, data_stage_5__4067_, data_stage_5__4066_, data_stage_5__4065_, data_stage_5__4064_, data_stage_5__4063_, data_stage_5__4062_, data_stage_5__4061_, data_stage_5__4060_, data_stage_5__4059_, data_stage_5__4058_, data_stage_5__4057_, data_stage_5__4056_, data_stage_5__4055_, data_stage_5__4054_, data_stage_5__4053_, data_stage_5__4052_, data_stage_5__4051_, data_stage_5__4050_, data_stage_5__4049_, data_stage_5__4048_, data_stage_5__4047_, data_stage_5__4046_, data_stage_5__4045_, data_stage_5__4044_, data_stage_5__4043_, data_stage_5__4042_, data_stage_5__4041_, data_stage_5__4040_, data_stage_5__4039_, data_stage_5__4038_, data_stage_5__4037_, data_stage_5__4036_, data_stage_5__4035_, data_stage_5__4034_, data_stage_5__4033_, data_stage_5__4032_, data_stage_5__4031_, data_stage_5__4030_, data_stage_5__4029_, data_stage_5__4028_, data_stage_5__4027_, data_stage_5__4026_, data_stage_5__4025_, data_stage_5__4024_, data_stage_5__4023_, data_stage_5__4022_, data_stage_5__4021_, data_stage_5__4020_, data_stage_5__4019_, data_stage_5__4018_, data_stage_5__4017_, data_stage_5__4016_, data_stage_5__4015_, data_stage_5__4014_, data_stage_5__4013_, data_stage_5__4012_, data_stage_5__4011_, data_stage_5__4010_, data_stage_5__4009_, data_stage_5__4008_, data_stage_5__4007_, data_stage_5__4006_, data_stage_5__4005_, data_stage_5__4004_, data_stage_5__4003_, data_stage_5__4002_, data_stage_5__4001_, data_stage_5__4000_, data_stage_5__3999_, data_stage_5__3998_, data_stage_5__3997_, data_stage_5__3996_, data_stage_5__3995_, data_stage_5__3994_, data_stage_5__3993_, data_stage_5__3992_, data_stage_5__3991_, data_stage_5__3990_, data_stage_5__3989_, data_stage_5__3988_, data_stage_5__3987_, data_stage_5__3986_, data_stage_5__3985_, data_stage_5__3984_, data_stage_5__3983_, data_stage_5__3982_, data_stage_5__3981_, data_stage_5__3980_, data_stage_5__3979_, data_stage_5__3978_, data_stage_5__3977_, data_stage_5__3976_, data_stage_5__3975_, data_stage_5__3974_, data_stage_5__3973_, data_stage_5__3972_, data_stage_5__3971_, data_stage_5__3970_, data_stage_5__3969_, data_stage_5__3968_, data_stage_5__3967_, data_stage_5__3966_, data_stage_5__3965_, data_stage_5__3964_, data_stage_5__3963_, data_stage_5__3962_, data_stage_5__3961_, data_stage_5__3960_, data_stage_5__3959_, data_stage_5__3958_, data_stage_5__3957_, data_stage_5__3956_, data_stage_5__3955_, data_stage_5__3954_, data_stage_5__3953_, data_stage_5__3952_, data_stage_5__3951_, data_stage_5__3950_, data_stage_5__3949_, data_stage_5__3948_, data_stage_5__3947_, data_stage_5__3946_, data_stage_5__3945_, data_stage_5__3944_, data_stage_5__3943_, data_stage_5__3942_, data_stage_5__3941_, data_stage_5__3940_, data_stage_5__3939_, data_stage_5__3938_, data_stage_5__3937_, data_stage_5__3936_, data_stage_5__3935_, data_stage_5__3934_, data_stage_5__3933_, data_stage_5__3932_, data_stage_5__3931_, data_stage_5__3930_, data_stage_5__3929_, data_stage_5__3928_, data_stage_5__3927_, data_stage_5__3926_, data_stage_5__3925_, data_stage_5__3924_, data_stage_5__3923_, data_stage_5__3922_, data_stage_5__3921_, data_stage_5__3920_, data_stage_5__3919_, data_stage_5__3918_, data_stage_5__3917_, data_stage_5__3916_, data_stage_5__3915_, data_stage_5__3914_, data_stage_5__3913_, data_stage_5__3912_, data_stage_5__3911_, data_stage_5__3910_, data_stage_5__3909_, data_stage_5__3908_, data_stage_5__3907_, data_stage_5__3906_, data_stage_5__3905_, data_stage_5__3904_, data_stage_5__3903_, data_stage_5__3902_, data_stage_5__3901_, data_stage_5__3900_, data_stage_5__3899_, data_stage_5__3898_, data_stage_5__3897_, data_stage_5__3896_, data_stage_5__3895_, data_stage_5__3894_, data_stage_5__3893_, data_stage_5__3892_, data_stage_5__3891_, data_stage_5__3890_, data_stage_5__3889_, data_stage_5__3888_, data_stage_5__3887_, data_stage_5__3886_, data_stage_5__3885_, data_stage_5__3884_, data_stage_5__3883_, data_stage_5__3882_, data_stage_5__3881_, data_stage_5__3880_, data_stage_5__3879_, data_stage_5__3878_, data_stage_5__3877_, data_stage_5__3876_, data_stage_5__3875_, data_stage_5__3874_, data_stage_5__3873_, data_stage_5__3872_, data_stage_5__3871_, data_stage_5__3870_, data_stage_5__3869_, data_stage_5__3868_, data_stage_5__3867_, data_stage_5__3866_, data_stage_5__3865_, data_stage_5__3864_, data_stage_5__3863_, data_stage_5__3862_, data_stage_5__3861_, data_stage_5__3860_, data_stage_5__3859_, data_stage_5__3858_, data_stage_5__3857_, data_stage_5__3856_, data_stage_5__3855_, data_stage_5__3854_, data_stage_5__3853_, data_stage_5__3852_, data_stage_5__3851_, data_stage_5__3850_, data_stage_5__3849_, data_stage_5__3848_, data_stage_5__3847_, data_stage_5__3846_, data_stage_5__3845_, data_stage_5__3844_, data_stage_5__3843_, data_stage_5__3842_, data_stage_5__3841_, data_stage_5__3840_, data_stage_5__3839_, data_stage_5__3838_, data_stage_5__3837_, data_stage_5__3836_, data_stage_5__3835_, data_stage_5__3834_, data_stage_5__3833_, data_stage_5__3832_, data_stage_5__3831_, data_stage_5__3830_, data_stage_5__3829_, data_stage_5__3828_, data_stage_5__3827_, data_stage_5__3826_, data_stage_5__3825_, data_stage_5__3824_, data_stage_5__3823_, data_stage_5__3822_, data_stage_5__3821_, data_stage_5__3820_, data_stage_5__3819_, data_stage_5__3818_, data_stage_5__3817_, data_stage_5__3816_, data_stage_5__3815_, data_stage_5__3814_, data_stage_5__3813_, data_stage_5__3812_, data_stage_5__3811_, data_stage_5__3810_, data_stage_5__3809_, data_stage_5__3808_, data_stage_5__3807_, data_stage_5__3806_, data_stage_5__3805_, data_stage_5__3804_, data_stage_5__3803_, data_stage_5__3802_, data_stage_5__3801_, data_stage_5__3800_, data_stage_5__3799_, data_stage_5__3798_, data_stage_5__3797_, data_stage_5__3796_, data_stage_5__3795_, data_stage_5__3794_, data_stage_5__3793_, data_stage_5__3792_, data_stage_5__3791_, data_stage_5__3790_, data_stage_5__3789_, data_stage_5__3788_, data_stage_5__3787_, data_stage_5__3786_, data_stage_5__3785_, data_stage_5__3784_, data_stage_5__3783_, data_stage_5__3782_, data_stage_5__3781_, data_stage_5__3780_, data_stage_5__3779_, data_stage_5__3778_, data_stage_5__3777_, data_stage_5__3776_, data_stage_5__3775_, data_stage_5__3774_, data_stage_5__3773_, data_stage_5__3772_, data_stage_5__3771_, data_stage_5__3770_, data_stage_5__3769_, data_stage_5__3768_, data_stage_5__3767_, data_stage_5__3766_, data_stage_5__3765_, data_stage_5__3764_, data_stage_5__3763_, data_stage_5__3762_, data_stage_5__3761_, data_stage_5__3760_, data_stage_5__3759_, data_stage_5__3758_, data_stage_5__3757_, data_stage_5__3756_, data_stage_5__3755_, data_stage_5__3754_, data_stage_5__3753_, data_stage_5__3752_, data_stage_5__3751_, data_stage_5__3750_, data_stage_5__3749_, data_stage_5__3748_, data_stage_5__3747_, data_stage_5__3746_, data_stage_5__3745_, data_stage_5__3744_, data_stage_5__3743_, data_stage_5__3742_, data_stage_5__3741_, data_stage_5__3740_, data_stage_5__3739_, data_stage_5__3738_, data_stage_5__3737_, data_stage_5__3736_, data_stage_5__3735_, data_stage_5__3734_, data_stage_5__3733_, data_stage_5__3732_, data_stage_5__3731_, data_stage_5__3730_, data_stage_5__3729_, data_stage_5__3728_, data_stage_5__3727_, data_stage_5__3726_, data_stage_5__3725_, data_stage_5__3724_, data_stage_5__3723_, data_stage_5__3722_, data_stage_5__3721_, data_stage_5__3720_, data_stage_5__3719_, data_stage_5__3718_, data_stage_5__3717_, data_stage_5__3716_, data_stage_5__3715_, data_stage_5__3714_, data_stage_5__3713_, data_stage_5__3712_, data_stage_5__3711_, data_stage_5__3710_, data_stage_5__3709_, data_stage_5__3708_, data_stage_5__3707_, data_stage_5__3706_, data_stage_5__3705_, data_stage_5__3704_, data_stage_5__3703_, data_stage_5__3702_, data_stage_5__3701_, data_stage_5__3700_, data_stage_5__3699_, data_stage_5__3698_, data_stage_5__3697_, data_stage_5__3696_, data_stage_5__3695_, data_stage_5__3694_, data_stage_5__3693_, data_stage_5__3692_, data_stage_5__3691_, data_stage_5__3690_, data_stage_5__3689_, data_stage_5__3688_, data_stage_5__3687_, data_stage_5__3686_, data_stage_5__3685_, data_stage_5__3684_, data_stage_5__3683_, data_stage_5__3682_, data_stage_5__3681_, data_stage_5__3680_, data_stage_5__3679_, data_stage_5__3678_, data_stage_5__3677_, data_stage_5__3676_, data_stage_5__3675_, data_stage_5__3674_, data_stage_5__3673_, data_stage_5__3672_, data_stage_5__3671_, data_stage_5__3670_, data_stage_5__3669_, data_stage_5__3668_, data_stage_5__3667_, data_stage_5__3666_, data_stage_5__3665_, data_stage_5__3664_, data_stage_5__3663_, data_stage_5__3662_, data_stage_5__3661_, data_stage_5__3660_, data_stage_5__3659_, data_stage_5__3658_, data_stage_5__3657_, data_stage_5__3656_, data_stage_5__3655_, data_stage_5__3654_, data_stage_5__3653_, data_stage_5__3652_, data_stage_5__3651_, data_stage_5__3650_, data_stage_5__3649_, data_stage_5__3648_, data_stage_5__3647_, data_stage_5__3646_, data_stage_5__3645_, data_stage_5__3644_, data_stage_5__3643_, data_stage_5__3642_, data_stage_5__3641_, data_stage_5__3640_, data_stage_5__3639_, data_stage_5__3638_, data_stage_5__3637_, data_stage_5__3636_, data_stage_5__3635_, data_stage_5__3634_, data_stage_5__3633_, data_stage_5__3632_, data_stage_5__3631_, data_stage_5__3630_, data_stage_5__3629_, data_stage_5__3628_, data_stage_5__3627_, data_stage_5__3626_, data_stage_5__3625_, data_stage_5__3624_, data_stage_5__3623_, data_stage_5__3622_, data_stage_5__3621_, data_stage_5__3620_, data_stage_5__3619_, data_stage_5__3618_, data_stage_5__3617_, data_stage_5__3616_, data_stage_5__3615_, data_stage_5__3614_, data_stage_5__3613_, data_stage_5__3612_, data_stage_5__3611_, data_stage_5__3610_, data_stage_5__3609_, data_stage_5__3608_, data_stage_5__3607_, data_stage_5__3606_, data_stage_5__3605_, data_stage_5__3604_, data_stage_5__3603_, data_stage_5__3602_, data_stage_5__3601_, data_stage_5__3600_, data_stage_5__3599_, data_stage_5__3598_, data_stage_5__3597_, data_stage_5__3596_, data_stage_5__3595_, data_stage_5__3594_, data_stage_5__3593_, data_stage_5__3592_, data_stage_5__3591_, data_stage_5__3590_, data_stage_5__3589_, data_stage_5__3588_, data_stage_5__3587_, data_stage_5__3586_, data_stage_5__3585_, data_stage_5__3584_, data_stage_5__3583_, data_stage_5__3582_, data_stage_5__3581_, data_stage_5__3580_, data_stage_5__3579_, data_stage_5__3578_, data_stage_5__3577_, data_stage_5__3576_, data_stage_5__3575_, data_stage_5__3574_, data_stage_5__3573_, data_stage_5__3572_, data_stage_5__3571_, data_stage_5__3570_, data_stage_5__3569_, data_stage_5__3568_, data_stage_5__3567_, data_stage_5__3566_, data_stage_5__3565_, data_stage_5__3564_, data_stage_5__3563_, data_stage_5__3562_, data_stage_5__3561_, data_stage_5__3560_, data_stage_5__3559_, data_stage_5__3558_, data_stage_5__3557_, data_stage_5__3556_, data_stage_5__3555_, data_stage_5__3554_, data_stage_5__3553_, data_stage_5__3552_, data_stage_5__3551_, data_stage_5__3550_, data_stage_5__3549_, data_stage_5__3548_, data_stage_5__3547_, data_stage_5__3546_, data_stage_5__3545_, data_stage_5__3544_, data_stage_5__3543_, data_stage_5__3542_, data_stage_5__3541_, data_stage_5__3540_, data_stage_5__3539_, data_stage_5__3538_, data_stage_5__3537_, data_stage_5__3536_, data_stage_5__3535_, data_stage_5__3534_, data_stage_5__3533_, data_stage_5__3532_, data_stage_5__3531_, data_stage_5__3530_, data_stage_5__3529_, data_stage_5__3528_, data_stage_5__3527_, data_stage_5__3526_, data_stage_5__3525_, data_stage_5__3524_, data_stage_5__3523_, data_stage_5__3522_, data_stage_5__3521_, data_stage_5__3520_, data_stage_5__3519_, data_stage_5__3518_, data_stage_5__3517_, data_stage_5__3516_, data_stage_5__3515_, data_stage_5__3514_, data_stage_5__3513_, data_stage_5__3512_, data_stage_5__3511_, data_stage_5__3510_, data_stage_5__3509_, data_stage_5__3508_, data_stage_5__3507_, data_stage_5__3506_, data_stage_5__3505_, data_stage_5__3504_, data_stage_5__3503_, data_stage_5__3502_, data_stage_5__3501_, data_stage_5__3500_, data_stage_5__3499_, data_stage_5__3498_, data_stage_5__3497_, data_stage_5__3496_, data_stage_5__3495_, data_stage_5__3494_, data_stage_5__3493_, data_stage_5__3492_, data_stage_5__3491_, data_stage_5__3490_, data_stage_5__3489_, data_stage_5__3488_, data_stage_5__3487_, data_stage_5__3486_, data_stage_5__3485_, data_stage_5__3484_, data_stage_5__3483_, data_stage_5__3482_, data_stage_5__3481_, data_stage_5__3480_, data_stage_5__3479_, data_stage_5__3478_, data_stage_5__3477_, data_stage_5__3476_, data_stage_5__3475_, data_stage_5__3474_, data_stage_5__3473_, data_stage_5__3472_, data_stage_5__3471_, data_stage_5__3470_, data_stage_5__3469_, data_stage_5__3468_, data_stage_5__3467_, data_stage_5__3466_, data_stage_5__3465_, data_stage_5__3464_, data_stage_5__3463_, data_stage_5__3462_, data_stage_5__3461_, data_stage_5__3460_, data_stage_5__3459_, data_stage_5__3458_, data_stage_5__3457_, data_stage_5__3456_, data_stage_5__3455_, data_stage_5__3454_, data_stage_5__3453_, data_stage_5__3452_, data_stage_5__3451_, data_stage_5__3450_, data_stage_5__3449_, data_stage_5__3448_, data_stage_5__3447_, data_stage_5__3446_, data_stage_5__3445_, data_stage_5__3444_, data_stage_5__3443_, data_stage_5__3442_, data_stage_5__3441_, data_stage_5__3440_, data_stage_5__3439_, data_stage_5__3438_, data_stage_5__3437_, data_stage_5__3436_, data_stage_5__3435_, data_stage_5__3434_, data_stage_5__3433_, data_stage_5__3432_, data_stage_5__3431_, data_stage_5__3430_, data_stage_5__3429_, data_stage_5__3428_, data_stage_5__3427_, data_stage_5__3426_, data_stage_5__3425_, data_stage_5__3424_, data_stage_5__3423_, data_stage_5__3422_, data_stage_5__3421_, data_stage_5__3420_, data_stage_5__3419_, data_stage_5__3418_, data_stage_5__3417_, data_stage_5__3416_, data_stage_5__3415_, data_stage_5__3414_, data_stage_5__3413_, data_stage_5__3412_, data_stage_5__3411_, data_stage_5__3410_, data_stage_5__3409_, data_stage_5__3408_, data_stage_5__3407_, data_stage_5__3406_, data_stage_5__3405_, data_stage_5__3404_, data_stage_5__3403_, data_stage_5__3402_, data_stage_5__3401_, data_stage_5__3400_, data_stage_5__3399_, data_stage_5__3398_, data_stage_5__3397_, data_stage_5__3396_, data_stage_5__3395_, data_stage_5__3394_, data_stage_5__3393_, data_stage_5__3392_, data_stage_5__3391_, data_stage_5__3390_, data_stage_5__3389_, data_stage_5__3388_, data_stage_5__3387_, data_stage_5__3386_, data_stage_5__3385_, data_stage_5__3384_, data_stage_5__3383_, data_stage_5__3382_, data_stage_5__3381_, data_stage_5__3380_, data_stage_5__3379_, data_stage_5__3378_, data_stage_5__3377_, data_stage_5__3376_, data_stage_5__3375_, data_stage_5__3374_, data_stage_5__3373_, data_stage_5__3372_, data_stage_5__3371_, data_stage_5__3370_, data_stage_5__3369_, data_stage_5__3368_, data_stage_5__3367_, data_stage_5__3366_, data_stage_5__3365_, data_stage_5__3364_, data_stage_5__3363_, data_stage_5__3362_, data_stage_5__3361_, data_stage_5__3360_, data_stage_5__3359_, data_stage_5__3358_, data_stage_5__3357_, data_stage_5__3356_, data_stage_5__3355_, data_stage_5__3354_, data_stage_5__3353_, data_stage_5__3352_, data_stage_5__3351_, data_stage_5__3350_, data_stage_5__3349_, data_stage_5__3348_, data_stage_5__3347_, data_stage_5__3346_, data_stage_5__3345_, data_stage_5__3344_, data_stage_5__3343_, data_stage_5__3342_, data_stage_5__3341_, data_stage_5__3340_, data_stage_5__3339_, data_stage_5__3338_, data_stage_5__3337_, data_stage_5__3336_, data_stage_5__3335_, data_stage_5__3334_, data_stage_5__3333_, data_stage_5__3332_, data_stage_5__3331_, data_stage_5__3330_, data_stage_5__3329_, data_stage_5__3328_, data_stage_5__3327_, data_stage_5__3326_, data_stage_5__3325_, data_stage_5__3324_, data_stage_5__3323_, data_stage_5__3322_, data_stage_5__3321_, data_stage_5__3320_, data_stage_5__3319_, data_stage_5__3318_, data_stage_5__3317_, data_stage_5__3316_, data_stage_5__3315_, data_stage_5__3314_, data_stage_5__3313_, data_stage_5__3312_, data_stage_5__3311_, data_stage_5__3310_, data_stage_5__3309_, data_stage_5__3308_, data_stage_5__3307_, data_stage_5__3306_, data_stage_5__3305_, data_stage_5__3304_, data_stage_5__3303_, data_stage_5__3302_, data_stage_5__3301_, data_stage_5__3300_, data_stage_5__3299_, data_stage_5__3298_, data_stage_5__3297_, data_stage_5__3296_, data_stage_5__3295_, data_stage_5__3294_, data_stage_5__3293_, data_stage_5__3292_, data_stage_5__3291_, data_stage_5__3290_, data_stage_5__3289_, data_stage_5__3288_, data_stage_5__3287_, data_stage_5__3286_, data_stage_5__3285_, data_stage_5__3284_, data_stage_5__3283_, data_stage_5__3282_, data_stage_5__3281_, data_stage_5__3280_, data_stage_5__3279_, data_stage_5__3278_, data_stage_5__3277_, data_stage_5__3276_, data_stage_5__3275_, data_stage_5__3274_, data_stage_5__3273_, data_stage_5__3272_, data_stage_5__3271_, data_stage_5__3270_, data_stage_5__3269_, data_stage_5__3268_, data_stage_5__3267_, data_stage_5__3266_, data_stage_5__3265_, data_stage_5__3264_, data_stage_5__3263_, data_stage_5__3262_, data_stage_5__3261_, data_stage_5__3260_, data_stage_5__3259_, data_stage_5__3258_, data_stage_5__3257_, data_stage_5__3256_, data_stage_5__3255_, data_stage_5__3254_, data_stage_5__3253_, data_stage_5__3252_, data_stage_5__3251_, data_stage_5__3250_, data_stage_5__3249_, data_stage_5__3248_, data_stage_5__3247_, data_stage_5__3246_, data_stage_5__3245_, data_stage_5__3244_, data_stage_5__3243_, data_stage_5__3242_, data_stage_5__3241_, data_stage_5__3240_, data_stage_5__3239_, data_stage_5__3238_, data_stage_5__3237_, data_stage_5__3236_, data_stage_5__3235_, data_stage_5__3234_, data_stage_5__3233_, data_stage_5__3232_, data_stage_5__3231_, data_stage_5__3230_, data_stage_5__3229_, data_stage_5__3228_, data_stage_5__3227_, data_stage_5__3226_, data_stage_5__3225_, data_stage_5__3224_, data_stage_5__3223_, data_stage_5__3222_, data_stage_5__3221_, data_stage_5__3220_, data_stage_5__3219_, data_stage_5__3218_, data_stage_5__3217_, data_stage_5__3216_, data_stage_5__3215_, data_stage_5__3214_, data_stage_5__3213_, data_stage_5__3212_, data_stage_5__3211_, data_stage_5__3210_, data_stage_5__3209_, data_stage_5__3208_, data_stage_5__3207_, data_stage_5__3206_, data_stage_5__3205_, data_stage_5__3204_, data_stage_5__3203_, data_stage_5__3202_, data_stage_5__3201_, data_stage_5__3200_, data_stage_5__3199_, data_stage_5__3198_, data_stage_5__3197_, data_stage_5__3196_, data_stage_5__3195_, data_stage_5__3194_, data_stage_5__3193_, data_stage_5__3192_, data_stage_5__3191_, data_stage_5__3190_, data_stage_5__3189_, data_stage_5__3188_, data_stage_5__3187_, data_stage_5__3186_, data_stage_5__3185_, data_stage_5__3184_, data_stage_5__3183_, data_stage_5__3182_, data_stage_5__3181_, data_stage_5__3180_, data_stage_5__3179_, data_stage_5__3178_, data_stage_5__3177_, data_stage_5__3176_, data_stage_5__3175_, data_stage_5__3174_, data_stage_5__3173_, data_stage_5__3172_, data_stage_5__3171_, data_stage_5__3170_, data_stage_5__3169_, data_stage_5__3168_, data_stage_5__3167_, data_stage_5__3166_, data_stage_5__3165_, data_stage_5__3164_, data_stage_5__3163_, data_stage_5__3162_, data_stage_5__3161_, data_stage_5__3160_, data_stage_5__3159_, data_stage_5__3158_, data_stage_5__3157_, data_stage_5__3156_, data_stage_5__3155_, data_stage_5__3154_, data_stage_5__3153_, data_stage_5__3152_, data_stage_5__3151_, data_stage_5__3150_, data_stage_5__3149_, data_stage_5__3148_, data_stage_5__3147_, data_stage_5__3146_, data_stage_5__3145_, data_stage_5__3144_, data_stage_5__3143_, data_stage_5__3142_, data_stage_5__3141_, data_stage_5__3140_, data_stage_5__3139_, data_stage_5__3138_, data_stage_5__3137_, data_stage_5__3136_, data_stage_5__3135_, data_stage_5__3134_, data_stage_5__3133_, data_stage_5__3132_, data_stage_5__3131_, data_stage_5__3130_, data_stage_5__3129_, data_stage_5__3128_, data_stage_5__3127_, data_stage_5__3126_, data_stage_5__3125_, data_stage_5__3124_, data_stage_5__3123_, data_stage_5__3122_, data_stage_5__3121_, data_stage_5__3120_, data_stage_5__3119_, data_stage_5__3118_, data_stage_5__3117_, data_stage_5__3116_, data_stage_5__3115_, data_stage_5__3114_, data_stage_5__3113_, data_stage_5__3112_, data_stage_5__3111_, data_stage_5__3110_, data_stage_5__3109_, data_stage_5__3108_, data_stage_5__3107_, data_stage_5__3106_, data_stage_5__3105_, data_stage_5__3104_, data_stage_5__3103_, data_stage_5__3102_, data_stage_5__3101_, data_stage_5__3100_, data_stage_5__3099_, data_stage_5__3098_, data_stage_5__3097_, data_stage_5__3096_, data_stage_5__3095_, data_stage_5__3094_, data_stage_5__3093_, data_stage_5__3092_, data_stage_5__3091_, data_stage_5__3090_, data_stage_5__3089_, data_stage_5__3088_, data_stage_5__3087_, data_stage_5__3086_, data_stage_5__3085_, data_stage_5__3084_, data_stage_5__3083_, data_stage_5__3082_, data_stage_5__3081_, data_stage_5__3080_, data_stage_5__3079_, data_stage_5__3078_, data_stage_5__3077_, data_stage_5__3076_, data_stage_5__3075_, data_stage_5__3074_, data_stage_5__3073_, data_stage_5__3072_, data_stage_5__3071_, data_stage_5__3070_, data_stage_5__3069_, data_stage_5__3068_, data_stage_5__3067_, data_stage_5__3066_, data_stage_5__3065_, data_stage_5__3064_, data_stage_5__3063_, data_stage_5__3062_, data_stage_5__3061_, data_stage_5__3060_, data_stage_5__3059_, data_stage_5__3058_, data_stage_5__3057_, data_stage_5__3056_, data_stage_5__3055_, data_stage_5__3054_, data_stage_5__3053_, data_stage_5__3052_, data_stage_5__3051_, data_stage_5__3050_, data_stage_5__3049_, data_stage_5__3048_, data_stage_5__3047_, data_stage_5__3046_, data_stage_5__3045_, data_stage_5__3044_, data_stage_5__3043_, data_stage_5__3042_, data_stage_5__3041_, data_stage_5__3040_, data_stage_5__3039_, data_stage_5__3038_, data_stage_5__3037_, data_stage_5__3036_, data_stage_5__3035_, data_stage_5__3034_, data_stage_5__3033_, data_stage_5__3032_, data_stage_5__3031_, data_stage_5__3030_, data_stage_5__3029_, data_stage_5__3028_, data_stage_5__3027_, data_stage_5__3026_, data_stage_5__3025_, data_stage_5__3024_, data_stage_5__3023_, data_stage_5__3022_, data_stage_5__3021_, data_stage_5__3020_, data_stage_5__3019_, data_stage_5__3018_, data_stage_5__3017_, data_stage_5__3016_, data_stage_5__3015_, data_stage_5__3014_, data_stage_5__3013_, data_stage_5__3012_, data_stage_5__3011_, data_stage_5__3010_, data_stage_5__3009_, data_stage_5__3008_, data_stage_5__3007_, data_stage_5__3006_, data_stage_5__3005_, data_stage_5__3004_, data_stage_5__3003_, data_stage_5__3002_, data_stage_5__3001_, data_stage_5__3000_, data_stage_5__2999_, data_stage_5__2998_, data_stage_5__2997_, data_stage_5__2996_, data_stage_5__2995_, data_stage_5__2994_, data_stage_5__2993_, data_stage_5__2992_, data_stage_5__2991_, data_stage_5__2990_, data_stage_5__2989_, data_stage_5__2988_, data_stage_5__2987_, data_stage_5__2986_, data_stage_5__2985_, data_stage_5__2984_, data_stage_5__2983_, data_stage_5__2982_, data_stage_5__2981_, data_stage_5__2980_, data_stage_5__2979_, data_stage_5__2978_, data_stage_5__2977_, data_stage_5__2976_, data_stage_5__2975_, data_stage_5__2974_, data_stage_5__2973_, data_stage_5__2972_, data_stage_5__2971_, data_stage_5__2970_, data_stage_5__2969_, data_stage_5__2968_, data_stage_5__2967_, data_stage_5__2966_, data_stage_5__2965_, data_stage_5__2964_, data_stage_5__2963_, data_stage_5__2962_, data_stage_5__2961_, data_stage_5__2960_, data_stage_5__2959_, data_stage_5__2958_, data_stage_5__2957_, data_stage_5__2956_, data_stage_5__2955_, data_stage_5__2954_, data_stage_5__2953_, data_stage_5__2952_, data_stage_5__2951_, data_stage_5__2950_, data_stage_5__2949_, data_stage_5__2948_, data_stage_5__2947_, data_stage_5__2946_, data_stage_5__2945_, data_stage_5__2944_, data_stage_5__2943_, data_stage_5__2942_, data_stage_5__2941_, data_stage_5__2940_, data_stage_5__2939_, data_stage_5__2938_, data_stage_5__2937_, data_stage_5__2936_, data_stage_5__2935_, data_stage_5__2934_, data_stage_5__2933_, data_stage_5__2932_, data_stage_5__2931_, data_stage_5__2930_, data_stage_5__2929_, data_stage_5__2928_, data_stage_5__2927_, data_stage_5__2926_, data_stage_5__2925_, data_stage_5__2924_, data_stage_5__2923_, data_stage_5__2922_, data_stage_5__2921_, data_stage_5__2920_, data_stage_5__2919_, data_stage_5__2918_, data_stage_5__2917_, data_stage_5__2916_, data_stage_5__2915_, data_stage_5__2914_, data_stage_5__2913_, data_stage_5__2912_, data_stage_5__2911_, data_stage_5__2910_, data_stage_5__2909_, data_stage_5__2908_, data_stage_5__2907_, data_stage_5__2906_, data_stage_5__2905_, data_stage_5__2904_, data_stage_5__2903_, data_stage_5__2902_, data_stage_5__2901_, data_stage_5__2900_, data_stage_5__2899_, data_stage_5__2898_, data_stage_5__2897_, data_stage_5__2896_, data_stage_5__2895_, data_stage_5__2894_, data_stage_5__2893_, data_stage_5__2892_, data_stage_5__2891_, data_stage_5__2890_, data_stage_5__2889_, data_stage_5__2888_, data_stage_5__2887_, data_stage_5__2886_, data_stage_5__2885_, data_stage_5__2884_, data_stage_5__2883_, data_stage_5__2882_, data_stage_5__2881_, data_stage_5__2880_, data_stage_5__2879_, data_stage_5__2878_, data_stage_5__2877_, data_stage_5__2876_, data_stage_5__2875_, data_stage_5__2874_, data_stage_5__2873_, data_stage_5__2872_, data_stage_5__2871_, data_stage_5__2870_, data_stage_5__2869_, data_stage_5__2868_, data_stage_5__2867_, data_stage_5__2866_, data_stage_5__2865_, data_stage_5__2864_, data_stage_5__2863_, data_stage_5__2862_, data_stage_5__2861_, data_stage_5__2860_, data_stage_5__2859_, data_stage_5__2858_, data_stage_5__2857_, data_stage_5__2856_, data_stage_5__2855_, data_stage_5__2854_, data_stage_5__2853_, data_stage_5__2852_, data_stage_5__2851_, data_stage_5__2850_, data_stage_5__2849_, data_stage_5__2848_, data_stage_5__2847_, data_stage_5__2846_, data_stage_5__2845_, data_stage_5__2844_, data_stage_5__2843_, data_stage_5__2842_, data_stage_5__2841_, data_stage_5__2840_, data_stage_5__2839_, data_stage_5__2838_, data_stage_5__2837_, data_stage_5__2836_, data_stage_5__2835_, data_stage_5__2834_, data_stage_5__2833_, data_stage_5__2832_, data_stage_5__2831_, data_stage_5__2830_, data_stage_5__2829_, data_stage_5__2828_, data_stage_5__2827_, data_stage_5__2826_, data_stage_5__2825_, data_stage_5__2824_, data_stage_5__2823_, data_stage_5__2822_, data_stage_5__2821_, data_stage_5__2820_, data_stage_5__2819_, data_stage_5__2818_, data_stage_5__2817_, data_stage_5__2816_, data_stage_5__2815_, data_stage_5__2814_, data_stage_5__2813_, data_stage_5__2812_, data_stage_5__2811_, data_stage_5__2810_, data_stage_5__2809_, data_stage_5__2808_, data_stage_5__2807_, data_stage_5__2806_, data_stage_5__2805_, data_stage_5__2804_, data_stage_5__2803_, data_stage_5__2802_, data_stage_5__2801_, data_stage_5__2800_, data_stage_5__2799_, data_stage_5__2798_, data_stage_5__2797_, data_stage_5__2796_, data_stage_5__2795_, data_stage_5__2794_, data_stage_5__2793_, data_stage_5__2792_, data_stage_5__2791_, data_stage_5__2790_, data_stage_5__2789_, data_stage_5__2788_, data_stage_5__2787_, data_stage_5__2786_, data_stage_5__2785_, data_stage_5__2784_, data_stage_5__2783_, data_stage_5__2782_, data_stage_5__2781_, data_stage_5__2780_, data_stage_5__2779_, data_stage_5__2778_, data_stage_5__2777_, data_stage_5__2776_, data_stage_5__2775_, data_stage_5__2774_, data_stage_5__2773_, data_stage_5__2772_, data_stage_5__2771_, data_stage_5__2770_, data_stage_5__2769_, data_stage_5__2768_, data_stage_5__2767_, data_stage_5__2766_, data_stage_5__2765_, data_stage_5__2764_, data_stage_5__2763_, data_stage_5__2762_, data_stage_5__2761_, data_stage_5__2760_, data_stage_5__2759_, data_stage_5__2758_, data_stage_5__2757_, data_stage_5__2756_, data_stage_5__2755_, data_stage_5__2754_, data_stage_5__2753_, data_stage_5__2752_, data_stage_5__2751_, data_stage_5__2750_, data_stage_5__2749_, data_stage_5__2748_, data_stage_5__2747_, data_stage_5__2746_, data_stage_5__2745_, data_stage_5__2744_, data_stage_5__2743_, data_stage_5__2742_, data_stage_5__2741_, data_stage_5__2740_, data_stage_5__2739_, data_stage_5__2738_, data_stage_5__2737_, data_stage_5__2736_, data_stage_5__2735_, data_stage_5__2734_, data_stage_5__2733_, data_stage_5__2732_, data_stage_5__2731_, data_stage_5__2730_, data_stage_5__2729_, data_stage_5__2728_, data_stage_5__2727_, data_stage_5__2726_, data_stage_5__2725_, data_stage_5__2724_, data_stage_5__2723_, data_stage_5__2722_, data_stage_5__2721_, data_stage_5__2720_, data_stage_5__2719_, data_stage_5__2718_, data_stage_5__2717_, data_stage_5__2716_, data_stage_5__2715_, data_stage_5__2714_, data_stage_5__2713_, data_stage_5__2712_, data_stage_5__2711_, data_stage_5__2710_, data_stage_5__2709_, data_stage_5__2708_, data_stage_5__2707_, data_stage_5__2706_, data_stage_5__2705_, data_stage_5__2704_, data_stage_5__2703_, data_stage_5__2702_, data_stage_5__2701_, data_stage_5__2700_, data_stage_5__2699_, data_stage_5__2698_, data_stage_5__2697_, data_stage_5__2696_, data_stage_5__2695_, data_stage_5__2694_, data_stage_5__2693_, data_stage_5__2692_, data_stage_5__2691_, data_stage_5__2690_, data_stage_5__2689_, data_stage_5__2688_, data_stage_5__2687_, data_stage_5__2686_, data_stage_5__2685_, data_stage_5__2684_, data_stage_5__2683_, data_stage_5__2682_, data_stage_5__2681_, data_stage_5__2680_, data_stage_5__2679_, data_stage_5__2678_, data_stage_5__2677_, data_stage_5__2676_, data_stage_5__2675_, data_stage_5__2674_, data_stage_5__2673_, data_stage_5__2672_, data_stage_5__2671_, data_stage_5__2670_, data_stage_5__2669_, data_stage_5__2668_, data_stage_5__2667_, data_stage_5__2666_, data_stage_5__2665_, data_stage_5__2664_, data_stage_5__2663_, data_stage_5__2662_, data_stage_5__2661_, data_stage_5__2660_, data_stage_5__2659_, data_stage_5__2658_, data_stage_5__2657_, data_stage_5__2656_, data_stage_5__2655_, data_stage_5__2654_, data_stage_5__2653_, data_stage_5__2652_, data_stage_5__2651_, data_stage_5__2650_, data_stage_5__2649_, data_stage_5__2648_, data_stage_5__2647_, data_stage_5__2646_, data_stage_5__2645_, data_stage_5__2644_, data_stage_5__2643_, data_stage_5__2642_, data_stage_5__2641_, data_stage_5__2640_, data_stage_5__2639_, data_stage_5__2638_, data_stage_5__2637_, data_stage_5__2636_, data_stage_5__2635_, data_stage_5__2634_, data_stage_5__2633_, data_stage_5__2632_, data_stage_5__2631_, data_stage_5__2630_, data_stage_5__2629_, data_stage_5__2628_, data_stage_5__2627_, data_stage_5__2626_, data_stage_5__2625_, data_stage_5__2624_, data_stage_5__2623_, data_stage_5__2622_, data_stage_5__2621_, data_stage_5__2620_, data_stage_5__2619_, data_stage_5__2618_, data_stage_5__2617_, data_stage_5__2616_, data_stage_5__2615_, data_stage_5__2614_, data_stage_5__2613_, data_stage_5__2612_, data_stage_5__2611_, data_stage_5__2610_, data_stage_5__2609_, data_stage_5__2608_, data_stage_5__2607_, data_stage_5__2606_, data_stage_5__2605_, data_stage_5__2604_, data_stage_5__2603_, data_stage_5__2602_, data_stage_5__2601_, data_stage_5__2600_, data_stage_5__2599_, data_stage_5__2598_, data_stage_5__2597_, data_stage_5__2596_, data_stage_5__2595_, data_stage_5__2594_, data_stage_5__2593_, data_stage_5__2592_, data_stage_5__2591_, data_stage_5__2590_, data_stage_5__2589_, data_stage_5__2588_, data_stage_5__2587_, data_stage_5__2586_, data_stage_5__2585_, data_stage_5__2584_, data_stage_5__2583_, data_stage_5__2582_, data_stage_5__2581_, data_stage_5__2580_, data_stage_5__2579_, data_stage_5__2578_, data_stage_5__2577_, data_stage_5__2576_, data_stage_5__2575_, data_stage_5__2574_, data_stage_5__2573_, data_stage_5__2572_, data_stage_5__2571_, data_stage_5__2570_, data_stage_5__2569_, data_stage_5__2568_, data_stage_5__2567_, data_stage_5__2566_, data_stage_5__2565_, data_stage_5__2564_, data_stage_5__2563_, data_stage_5__2562_, data_stage_5__2561_, data_stage_5__2560_, data_stage_5__2559_, data_stage_5__2558_, data_stage_5__2557_, data_stage_5__2556_, data_stage_5__2555_, data_stage_5__2554_, data_stage_5__2553_, data_stage_5__2552_, data_stage_5__2551_, data_stage_5__2550_, data_stage_5__2549_, data_stage_5__2548_, data_stage_5__2547_, data_stage_5__2546_, data_stage_5__2545_, data_stage_5__2544_, data_stage_5__2543_, data_stage_5__2542_, data_stage_5__2541_, data_stage_5__2540_, data_stage_5__2539_, data_stage_5__2538_, data_stage_5__2537_, data_stage_5__2536_, data_stage_5__2535_, data_stage_5__2534_, data_stage_5__2533_, data_stage_5__2532_, data_stage_5__2531_, data_stage_5__2530_, data_stage_5__2529_, data_stage_5__2528_, data_stage_5__2527_, data_stage_5__2526_, data_stage_5__2525_, data_stage_5__2524_, data_stage_5__2523_, data_stage_5__2522_, data_stage_5__2521_, data_stage_5__2520_, data_stage_5__2519_, data_stage_5__2518_, data_stage_5__2517_, data_stage_5__2516_, data_stage_5__2515_, data_stage_5__2514_, data_stage_5__2513_, data_stage_5__2512_, data_stage_5__2511_, data_stage_5__2510_, data_stage_5__2509_, data_stage_5__2508_, data_stage_5__2507_, data_stage_5__2506_, data_stage_5__2505_, data_stage_5__2504_, data_stage_5__2503_, data_stage_5__2502_, data_stage_5__2501_, data_stage_5__2500_, data_stage_5__2499_, data_stage_5__2498_, data_stage_5__2497_, data_stage_5__2496_, data_stage_5__2495_, data_stage_5__2494_, data_stage_5__2493_, data_stage_5__2492_, data_stage_5__2491_, data_stage_5__2490_, data_stage_5__2489_, data_stage_5__2488_, data_stage_5__2487_, data_stage_5__2486_, data_stage_5__2485_, data_stage_5__2484_, data_stage_5__2483_, data_stage_5__2482_, data_stage_5__2481_, data_stage_5__2480_, data_stage_5__2479_, data_stage_5__2478_, data_stage_5__2477_, data_stage_5__2476_, data_stage_5__2475_, data_stage_5__2474_, data_stage_5__2473_, data_stage_5__2472_, data_stage_5__2471_, data_stage_5__2470_, data_stage_5__2469_, data_stage_5__2468_, data_stage_5__2467_, data_stage_5__2466_, data_stage_5__2465_, data_stage_5__2464_, data_stage_5__2463_, data_stage_5__2462_, data_stage_5__2461_, data_stage_5__2460_, data_stage_5__2459_, data_stage_5__2458_, data_stage_5__2457_, data_stage_5__2456_, data_stage_5__2455_, data_stage_5__2454_, data_stage_5__2453_, data_stage_5__2452_, data_stage_5__2451_, data_stage_5__2450_, data_stage_5__2449_, data_stage_5__2448_, data_stage_5__2447_, data_stage_5__2446_, data_stage_5__2445_, data_stage_5__2444_, data_stage_5__2443_, data_stage_5__2442_, data_stage_5__2441_, data_stage_5__2440_, data_stage_5__2439_, data_stage_5__2438_, data_stage_5__2437_, data_stage_5__2436_, data_stage_5__2435_, data_stage_5__2434_, data_stage_5__2433_, data_stage_5__2432_, data_stage_5__2431_, data_stage_5__2430_, data_stage_5__2429_, data_stage_5__2428_, data_stage_5__2427_, data_stage_5__2426_, data_stage_5__2425_, data_stage_5__2424_, data_stage_5__2423_, data_stage_5__2422_, data_stage_5__2421_, data_stage_5__2420_, data_stage_5__2419_, data_stage_5__2418_, data_stage_5__2417_, data_stage_5__2416_, data_stage_5__2415_, data_stage_5__2414_, data_stage_5__2413_, data_stage_5__2412_, data_stage_5__2411_, data_stage_5__2410_, data_stage_5__2409_, data_stage_5__2408_, data_stage_5__2407_, data_stage_5__2406_, data_stage_5__2405_, data_stage_5__2404_, data_stage_5__2403_, data_stage_5__2402_, data_stage_5__2401_, data_stage_5__2400_, data_stage_5__2399_, data_stage_5__2398_, data_stage_5__2397_, data_stage_5__2396_, data_stage_5__2395_, data_stage_5__2394_, data_stage_5__2393_, data_stage_5__2392_, data_stage_5__2391_, data_stage_5__2390_, data_stage_5__2389_, data_stage_5__2388_, data_stage_5__2387_, data_stage_5__2386_, data_stage_5__2385_, data_stage_5__2384_, data_stage_5__2383_, data_stage_5__2382_, data_stage_5__2381_, data_stage_5__2380_, data_stage_5__2379_, data_stage_5__2378_, data_stage_5__2377_, data_stage_5__2376_, data_stage_5__2375_, data_stage_5__2374_, data_stage_5__2373_, data_stage_5__2372_, data_stage_5__2371_, data_stage_5__2370_, data_stage_5__2369_, data_stage_5__2368_, data_stage_5__2367_, data_stage_5__2366_, data_stage_5__2365_, data_stage_5__2364_, data_stage_5__2363_, data_stage_5__2362_, data_stage_5__2361_, data_stage_5__2360_, data_stage_5__2359_, data_stage_5__2358_, data_stage_5__2357_, data_stage_5__2356_, data_stage_5__2355_, data_stage_5__2354_, data_stage_5__2353_, data_stage_5__2352_, data_stage_5__2351_, data_stage_5__2350_, data_stage_5__2349_, data_stage_5__2348_, data_stage_5__2347_, data_stage_5__2346_, data_stage_5__2345_, data_stage_5__2344_, data_stage_5__2343_, data_stage_5__2342_, data_stage_5__2341_, data_stage_5__2340_, data_stage_5__2339_, data_stage_5__2338_, data_stage_5__2337_, data_stage_5__2336_, data_stage_5__2335_, data_stage_5__2334_, data_stage_5__2333_, data_stage_5__2332_, data_stage_5__2331_, data_stage_5__2330_, data_stage_5__2329_, data_stage_5__2328_, data_stage_5__2327_, data_stage_5__2326_, data_stage_5__2325_, data_stage_5__2324_, data_stage_5__2323_, data_stage_5__2322_, data_stage_5__2321_, data_stage_5__2320_, data_stage_5__2319_, data_stage_5__2318_, data_stage_5__2317_, data_stage_5__2316_, data_stage_5__2315_, data_stage_5__2314_, data_stage_5__2313_, data_stage_5__2312_, data_stage_5__2311_, data_stage_5__2310_, data_stage_5__2309_, data_stage_5__2308_, data_stage_5__2307_, data_stage_5__2306_, data_stage_5__2305_, data_stage_5__2304_, data_stage_5__2303_, data_stage_5__2302_, data_stage_5__2301_, data_stage_5__2300_, data_stage_5__2299_, data_stage_5__2298_, data_stage_5__2297_, data_stage_5__2296_, data_stage_5__2295_, data_stage_5__2294_, data_stage_5__2293_, data_stage_5__2292_, data_stage_5__2291_, data_stage_5__2290_, data_stage_5__2289_, data_stage_5__2288_, data_stage_5__2287_, data_stage_5__2286_, data_stage_5__2285_, data_stage_5__2284_, data_stage_5__2283_, data_stage_5__2282_, data_stage_5__2281_, data_stage_5__2280_, data_stage_5__2279_, data_stage_5__2278_, data_stage_5__2277_, data_stage_5__2276_, data_stage_5__2275_, data_stage_5__2274_, data_stage_5__2273_, data_stage_5__2272_, data_stage_5__2271_, data_stage_5__2270_, data_stage_5__2269_, data_stage_5__2268_, data_stage_5__2267_, data_stage_5__2266_, data_stage_5__2265_, data_stage_5__2264_, data_stage_5__2263_, data_stage_5__2262_, data_stage_5__2261_, data_stage_5__2260_, data_stage_5__2259_, data_stage_5__2258_, data_stage_5__2257_, data_stage_5__2256_, data_stage_5__2255_, data_stage_5__2254_, data_stage_5__2253_, data_stage_5__2252_, data_stage_5__2251_, data_stage_5__2250_, data_stage_5__2249_, data_stage_5__2248_, data_stage_5__2247_, data_stage_5__2246_, data_stage_5__2245_, data_stage_5__2244_, data_stage_5__2243_, data_stage_5__2242_, data_stage_5__2241_, data_stage_5__2240_, data_stage_5__2239_, data_stage_5__2238_, data_stage_5__2237_, data_stage_5__2236_, data_stage_5__2235_, data_stage_5__2234_, data_stage_5__2233_, data_stage_5__2232_, data_stage_5__2231_, data_stage_5__2230_, data_stage_5__2229_, data_stage_5__2228_, data_stage_5__2227_, data_stage_5__2226_, data_stage_5__2225_, data_stage_5__2224_, data_stage_5__2223_, data_stage_5__2222_, data_stage_5__2221_, data_stage_5__2220_, data_stage_5__2219_, data_stage_5__2218_, data_stage_5__2217_, data_stage_5__2216_, data_stage_5__2215_, data_stage_5__2214_, data_stage_5__2213_, data_stage_5__2212_, data_stage_5__2211_, data_stage_5__2210_, data_stage_5__2209_, data_stage_5__2208_, data_stage_5__2207_, data_stage_5__2206_, data_stage_5__2205_, data_stage_5__2204_, data_stage_5__2203_, data_stage_5__2202_, data_stage_5__2201_, data_stage_5__2200_, data_stage_5__2199_, data_stage_5__2198_, data_stage_5__2197_, data_stage_5__2196_, data_stage_5__2195_, data_stage_5__2194_, data_stage_5__2193_, data_stage_5__2192_, data_stage_5__2191_, data_stage_5__2190_, data_stage_5__2189_, data_stage_5__2188_, data_stage_5__2187_, data_stage_5__2186_, data_stage_5__2185_, data_stage_5__2184_, data_stage_5__2183_, data_stage_5__2182_, data_stage_5__2181_, data_stage_5__2180_, data_stage_5__2179_, data_stage_5__2178_, data_stage_5__2177_, data_stage_5__2176_, data_stage_5__2175_, data_stage_5__2174_, data_stage_5__2173_, data_stage_5__2172_, data_stage_5__2171_, data_stage_5__2170_, data_stage_5__2169_, data_stage_5__2168_, data_stage_5__2167_, data_stage_5__2166_, data_stage_5__2165_, data_stage_5__2164_, data_stage_5__2163_, data_stage_5__2162_, data_stage_5__2161_, data_stage_5__2160_, data_stage_5__2159_, data_stage_5__2158_, data_stage_5__2157_, data_stage_5__2156_, data_stage_5__2155_, data_stage_5__2154_, data_stage_5__2153_, data_stage_5__2152_, data_stage_5__2151_, data_stage_5__2150_, data_stage_5__2149_, data_stage_5__2148_, data_stage_5__2147_, data_stage_5__2146_, data_stage_5__2145_, data_stage_5__2144_, data_stage_5__2143_, data_stage_5__2142_, data_stage_5__2141_, data_stage_5__2140_, data_stage_5__2139_, data_stage_5__2138_, data_stage_5__2137_, data_stage_5__2136_, data_stage_5__2135_, data_stage_5__2134_, data_stage_5__2133_, data_stage_5__2132_, data_stage_5__2131_, data_stage_5__2130_, data_stage_5__2129_, data_stage_5__2128_, data_stage_5__2127_, data_stage_5__2126_, data_stage_5__2125_, data_stage_5__2124_, data_stage_5__2123_, data_stage_5__2122_, data_stage_5__2121_, data_stage_5__2120_, data_stage_5__2119_, data_stage_5__2118_, data_stage_5__2117_, data_stage_5__2116_, data_stage_5__2115_, data_stage_5__2114_, data_stage_5__2113_, data_stage_5__2112_, data_stage_5__2111_, data_stage_5__2110_, data_stage_5__2109_, data_stage_5__2108_, data_stage_5__2107_, data_stage_5__2106_, data_stage_5__2105_, data_stage_5__2104_, data_stage_5__2103_, data_stage_5__2102_, data_stage_5__2101_, data_stage_5__2100_, data_stage_5__2099_, data_stage_5__2098_, data_stage_5__2097_, data_stage_5__2096_, data_stage_5__2095_, data_stage_5__2094_, data_stage_5__2093_, data_stage_5__2092_, data_stage_5__2091_, data_stage_5__2090_, data_stage_5__2089_, data_stage_5__2088_, data_stage_5__2087_, data_stage_5__2086_, data_stage_5__2085_, data_stage_5__2084_, data_stage_5__2083_, data_stage_5__2082_, data_stage_5__2081_, data_stage_5__2080_, data_stage_5__2079_, data_stage_5__2078_, data_stage_5__2077_, data_stage_5__2076_, data_stage_5__2075_, data_stage_5__2074_, data_stage_5__2073_, data_stage_5__2072_, data_stage_5__2071_, data_stage_5__2070_, data_stage_5__2069_, data_stage_5__2068_, data_stage_5__2067_, data_stage_5__2066_, data_stage_5__2065_, data_stage_5__2064_, data_stage_5__2063_, data_stage_5__2062_, data_stage_5__2061_, data_stage_5__2060_, data_stage_5__2059_, data_stage_5__2058_, data_stage_5__2057_, data_stage_5__2056_, data_stage_5__2055_, data_stage_5__2054_, data_stage_5__2053_, data_stage_5__2052_, data_stage_5__2051_, data_stage_5__2050_, data_stage_5__2049_, data_stage_5__2048_, data_stage_5__2047_, data_stage_5__2046_, data_stage_5__2045_, data_stage_5__2044_, data_stage_5__2043_, data_stage_5__2042_, data_stage_5__2041_, data_stage_5__2040_, data_stage_5__2039_, data_stage_5__2038_, data_stage_5__2037_, data_stage_5__2036_, data_stage_5__2035_, data_stage_5__2034_, data_stage_5__2033_, data_stage_5__2032_, data_stage_5__2031_, data_stage_5__2030_, data_stage_5__2029_, data_stage_5__2028_, data_stage_5__2027_, data_stage_5__2026_, data_stage_5__2025_, data_stage_5__2024_, data_stage_5__2023_, data_stage_5__2022_, data_stage_5__2021_, data_stage_5__2020_, data_stage_5__2019_, data_stage_5__2018_, data_stage_5__2017_, data_stage_5__2016_, data_stage_5__2015_, data_stage_5__2014_, data_stage_5__2013_, data_stage_5__2012_, data_stage_5__2011_, data_stage_5__2010_, data_stage_5__2009_, data_stage_5__2008_, data_stage_5__2007_, data_stage_5__2006_, data_stage_5__2005_, data_stage_5__2004_, data_stage_5__2003_, data_stage_5__2002_, data_stage_5__2001_, data_stage_5__2000_, data_stage_5__1999_, data_stage_5__1998_, data_stage_5__1997_, data_stage_5__1996_, data_stage_5__1995_, data_stage_5__1994_, data_stage_5__1993_, data_stage_5__1992_, data_stage_5__1991_, data_stage_5__1990_, data_stage_5__1989_, data_stage_5__1988_, data_stage_5__1987_, data_stage_5__1986_, data_stage_5__1985_, data_stage_5__1984_, data_stage_5__1983_, data_stage_5__1982_, data_stage_5__1981_, data_stage_5__1980_, data_stage_5__1979_, data_stage_5__1978_, data_stage_5__1977_, data_stage_5__1976_, data_stage_5__1975_, data_stage_5__1974_, data_stage_5__1973_, data_stage_5__1972_, data_stage_5__1971_, data_stage_5__1970_, data_stage_5__1969_, data_stage_5__1968_, data_stage_5__1967_, data_stage_5__1966_, data_stage_5__1965_, data_stage_5__1964_, data_stage_5__1963_, data_stage_5__1962_, data_stage_5__1961_, data_stage_5__1960_, data_stage_5__1959_, data_stage_5__1958_, data_stage_5__1957_, data_stage_5__1956_, data_stage_5__1955_, data_stage_5__1954_, data_stage_5__1953_, data_stage_5__1952_, data_stage_5__1951_, data_stage_5__1950_, data_stage_5__1949_, data_stage_5__1948_, data_stage_5__1947_, data_stage_5__1946_, data_stage_5__1945_, data_stage_5__1944_, data_stage_5__1943_, data_stage_5__1942_, data_stage_5__1941_, data_stage_5__1940_, data_stage_5__1939_, data_stage_5__1938_, data_stage_5__1937_, data_stage_5__1936_, data_stage_5__1935_, data_stage_5__1934_, data_stage_5__1933_, data_stage_5__1932_, data_stage_5__1931_, data_stage_5__1930_, data_stage_5__1929_, data_stage_5__1928_, data_stage_5__1927_, data_stage_5__1926_, data_stage_5__1925_, data_stage_5__1924_, data_stage_5__1923_, data_stage_5__1922_, data_stage_5__1921_, data_stage_5__1920_, data_stage_5__1919_, data_stage_5__1918_, data_stage_5__1917_, data_stage_5__1916_, data_stage_5__1915_, data_stage_5__1914_, data_stage_5__1913_, data_stage_5__1912_, data_stage_5__1911_, data_stage_5__1910_, data_stage_5__1909_, data_stage_5__1908_, data_stage_5__1907_, data_stage_5__1906_, data_stage_5__1905_, data_stage_5__1904_, data_stage_5__1903_, data_stage_5__1902_, data_stage_5__1901_, data_stage_5__1900_, data_stage_5__1899_, data_stage_5__1898_, data_stage_5__1897_, data_stage_5__1896_, data_stage_5__1895_, data_stage_5__1894_, data_stage_5__1893_, data_stage_5__1892_, data_stage_5__1891_, data_stage_5__1890_, data_stage_5__1889_, data_stage_5__1888_, data_stage_5__1887_, data_stage_5__1886_, data_stage_5__1885_, data_stage_5__1884_, data_stage_5__1883_, data_stage_5__1882_, data_stage_5__1881_, data_stage_5__1880_, data_stage_5__1879_, data_stage_5__1878_, data_stage_5__1877_, data_stage_5__1876_, data_stage_5__1875_, data_stage_5__1874_, data_stage_5__1873_, data_stage_5__1872_, data_stage_5__1871_, data_stage_5__1870_, data_stage_5__1869_, data_stage_5__1868_, data_stage_5__1867_, data_stage_5__1866_, data_stage_5__1865_, data_stage_5__1864_, data_stage_5__1863_, data_stage_5__1862_, data_stage_5__1861_, data_stage_5__1860_, data_stage_5__1859_, data_stage_5__1858_, data_stage_5__1857_, data_stage_5__1856_, data_stage_5__1855_, data_stage_5__1854_, data_stage_5__1853_, data_stage_5__1852_, data_stage_5__1851_, data_stage_5__1850_, data_stage_5__1849_, data_stage_5__1848_, data_stage_5__1847_, data_stage_5__1846_, data_stage_5__1845_, data_stage_5__1844_, data_stage_5__1843_, data_stage_5__1842_, data_stage_5__1841_, data_stage_5__1840_, data_stage_5__1839_, data_stage_5__1838_, data_stage_5__1837_, data_stage_5__1836_, data_stage_5__1835_, data_stage_5__1834_, data_stage_5__1833_, data_stage_5__1832_, data_stage_5__1831_, data_stage_5__1830_, data_stage_5__1829_, data_stage_5__1828_, data_stage_5__1827_, data_stage_5__1826_, data_stage_5__1825_, data_stage_5__1824_, data_stage_5__1823_, data_stage_5__1822_, data_stage_5__1821_, data_stage_5__1820_, data_stage_5__1819_, data_stage_5__1818_, data_stage_5__1817_, data_stage_5__1816_, data_stage_5__1815_, data_stage_5__1814_, data_stage_5__1813_, data_stage_5__1812_, data_stage_5__1811_, data_stage_5__1810_, data_stage_5__1809_, data_stage_5__1808_, data_stage_5__1807_, data_stage_5__1806_, data_stage_5__1805_, data_stage_5__1804_, data_stage_5__1803_, data_stage_5__1802_, data_stage_5__1801_, data_stage_5__1800_, data_stage_5__1799_, data_stage_5__1798_, data_stage_5__1797_, data_stage_5__1796_, data_stage_5__1795_, data_stage_5__1794_, data_stage_5__1793_, data_stage_5__1792_, data_stage_5__1791_, data_stage_5__1790_, data_stage_5__1789_, data_stage_5__1788_, data_stage_5__1787_, data_stage_5__1786_, data_stage_5__1785_, data_stage_5__1784_, data_stage_5__1783_, data_stage_5__1782_, data_stage_5__1781_, data_stage_5__1780_, data_stage_5__1779_, data_stage_5__1778_, data_stage_5__1777_, data_stage_5__1776_, data_stage_5__1775_, data_stage_5__1774_, data_stage_5__1773_, data_stage_5__1772_, data_stage_5__1771_, data_stage_5__1770_, data_stage_5__1769_, data_stage_5__1768_, data_stage_5__1767_, data_stage_5__1766_, data_stage_5__1765_, data_stage_5__1764_, data_stage_5__1763_, data_stage_5__1762_, data_stage_5__1761_, data_stage_5__1760_, data_stage_5__1759_, data_stage_5__1758_, data_stage_5__1757_, data_stage_5__1756_, data_stage_5__1755_, data_stage_5__1754_, data_stage_5__1753_, data_stage_5__1752_, data_stage_5__1751_, data_stage_5__1750_, data_stage_5__1749_, data_stage_5__1748_, data_stage_5__1747_, data_stage_5__1746_, data_stage_5__1745_, data_stage_5__1744_, data_stage_5__1743_, data_stage_5__1742_, data_stage_5__1741_, data_stage_5__1740_, data_stage_5__1739_, data_stage_5__1738_, data_stage_5__1737_, data_stage_5__1736_, data_stage_5__1735_, data_stage_5__1734_, data_stage_5__1733_, data_stage_5__1732_, data_stage_5__1731_, data_stage_5__1730_, data_stage_5__1729_, data_stage_5__1728_, data_stage_5__1727_, data_stage_5__1726_, data_stage_5__1725_, data_stage_5__1724_, data_stage_5__1723_, data_stage_5__1722_, data_stage_5__1721_, data_stage_5__1720_, data_stage_5__1719_, data_stage_5__1718_, data_stage_5__1717_, data_stage_5__1716_, data_stage_5__1715_, data_stage_5__1714_, data_stage_5__1713_, data_stage_5__1712_, data_stage_5__1711_, data_stage_5__1710_, data_stage_5__1709_, data_stage_5__1708_, data_stage_5__1707_, data_stage_5__1706_, data_stage_5__1705_, data_stage_5__1704_, data_stage_5__1703_, data_stage_5__1702_, data_stage_5__1701_, data_stage_5__1700_, data_stage_5__1699_, data_stage_5__1698_, data_stage_5__1697_, data_stage_5__1696_, data_stage_5__1695_, data_stage_5__1694_, data_stage_5__1693_, data_stage_5__1692_, data_stage_5__1691_, data_stage_5__1690_, data_stage_5__1689_, data_stage_5__1688_, data_stage_5__1687_, data_stage_5__1686_, data_stage_5__1685_, data_stage_5__1684_, data_stage_5__1683_, data_stage_5__1682_, data_stage_5__1681_, data_stage_5__1680_, data_stage_5__1679_, data_stage_5__1678_, data_stage_5__1677_, data_stage_5__1676_, data_stage_5__1675_, data_stage_5__1674_, data_stage_5__1673_, data_stage_5__1672_, data_stage_5__1671_, data_stage_5__1670_, data_stage_5__1669_, data_stage_5__1668_, data_stage_5__1667_, data_stage_5__1666_, data_stage_5__1665_, data_stage_5__1664_, data_stage_5__1663_, data_stage_5__1662_, data_stage_5__1661_, data_stage_5__1660_, data_stage_5__1659_, data_stage_5__1658_, data_stage_5__1657_, data_stage_5__1656_, data_stage_5__1655_, data_stage_5__1654_, data_stage_5__1653_, data_stage_5__1652_, data_stage_5__1651_, data_stage_5__1650_, data_stage_5__1649_, data_stage_5__1648_, data_stage_5__1647_, data_stage_5__1646_, data_stage_5__1645_, data_stage_5__1644_, data_stage_5__1643_, data_stage_5__1642_, data_stage_5__1641_, data_stage_5__1640_, data_stage_5__1639_, data_stage_5__1638_, data_stage_5__1637_, data_stage_5__1636_, data_stage_5__1635_, data_stage_5__1634_, data_stage_5__1633_, data_stage_5__1632_, data_stage_5__1631_, data_stage_5__1630_, data_stage_5__1629_, data_stage_5__1628_, data_stage_5__1627_, data_stage_5__1626_, data_stage_5__1625_, data_stage_5__1624_, data_stage_5__1623_, data_stage_5__1622_, data_stage_5__1621_, data_stage_5__1620_, data_stage_5__1619_, data_stage_5__1618_, data_stage_5__1617_, data_stage_5__1616_, data_stage_5__1615_, data_stage_5__1614_, data_stage_5__1613_, data_stage_5__1612_, data_stage_5__1611_, data_stage_5__1610_, data_stage_5__1609_, data_stage_5__1608_, data_stage_5__1607_, data_stage_5__1606_, data_stage_5__1605_, data_stage_5__1604_, data_stage_5__1603_, data_stage_5__1602_, data_stage_5__1601_, data_stage_5__1600_, data_stage_5__1599_, data_stage_5__1598_, data_stage_5__1597_, data_stage_5__1596_, data_stage_5__1595_, data_stage_5__1594_, data_stage_5__1593_, data_stage_5__1592_, data_stage_5__1591_, data_stage_5__1590_, data_stage_5__1589_, data_stage_5__1588_, data_stage_5__1587_, data_stage_5__1586_, data_stage_5__1585_, data_stage_5__1584_, data_stage_5__1583_, data_stage_5__1582_, data_stage_5__1581_, data_stage_5__1580_, data_stage_5__1579_, data_stage_5__1578_, data_stage_5__1577_, data_stage_5__1576_, data_stage_5__1575_, data_stage_5__1574_, data_stage_5__1573_, data_stage_5__1572_, data_stage_5__1571_, data_stage_5__1570_, data_stage_5__1569_, data_stage_5__1568_, data_stage_5__1567_, data_stage_5__1566_, data_stage_5__1565_, data_stage_5__1564_, data_stage_5__1563_, data_stage_5__1562_, data_stage_5__1561_, data_stage_5__1560_, data_stage_5__1559_, data_stage_5__1558_, data_stage_5__1557_, data_stage_5__1556_, data_stage_5__1555_, data_stage_5__1554_, data_stage_5__1553_, data_stage_5__1552_, data_stage_5__1551_, data_stage_5__1550_, data_stage_5__1549_, data_stage_5__1548_, data_stage_5__1547_, data_stage_5__1546_, data_stage_5__1545_, data_stage_5__1544_, data_stage_5__1543_, data_stage_5__1542_, data_stage_5__1541_, data_stage_5__1540_, data_stage_5__1539_, data_stage_5__1538_, data_stage_5__1537_, data_stage_5__1536_, data_stage_5__1535_, data_stage_5__1534_, data_stage_5__1533_, data_stage_5__1532_, data_stage_5__1531_, data_stage_5__1530_, data_stage_5__1529_, data_stage_5__1528_, data_stage_5__1527_, data_stage_5__1526_, data_stage_5__1525_, data_stage_5__1524_, data_stage_5__1523_, data_stage_5__1522_, data_stage_5__1521_, data_stage_5__1520_, data_stage_5__1519_, data_stage_5__1518_, data_stage_5__1517_, data_stage_5__1516_, data_stage_5__1515_, data_stage_5__1514_, data_stage_5__1513_, data_stage_5__1512_, data_stage_5__1511_, data_stage_5__1510_, data_stage_5__1509_, data_stage_5__1508_, data_stage_5__1507_, data_stage_5__1506_, data_stage_5__1505_, data_stage_5__1504_, data_stage_5__1503_, data_stage_5__1502_, data_stage_5__1501_, data_stage_5__1500_, data_stage_5__1499_, data_stage_5__1498_, data_stage_5__1497_, data_stage_5__1496_, data_stage_5__1495_, data_stage_5__1494_, data_stage_5__1493_, data_stage_5__1492_, data_stage_5__1491_, data_stage_5__1490_, data_stage_5__1489_, data_stage_5__1488_, data_stage_5__1487_, data_stage_5__1486_, data_stage_5__1485_, data_stage_5__1484_, data_stage_5__1483_, data_stage_5__1482_, data_stage_5__1481_, data_stage_5__1480_, data_stage_5__1479_, data_stage_5__1478_, data_stage_5__1477_, data_stage_5__1476_, data_stage_5__1475_, data_stage_5__1474_, data_stage_5__1473_, data_stage_5__1472_, data_stage_5__1471_, data_stage_5__1470_, data_stage_5__1469_, data_stage_5__1468_, data_stage_5__1467_, data_stage_5__1466_, data_stage_5__1465_, data_stage_5__1464_, data_stage_5__1463_, data_stage_5__1462_, data_stage_5__1461_, data_stage_5__1460_, data_stage_5__1459_, data_stage_5__1458_, data_stage_5__1457_, data_stage_5__1456_, data_stage_5__1455_, data_stage_5__1454_, data_stage_5__1453_, data_stage_5__1452_, data_stage_5__1451_, data_stage_5__1450_, data_stage_5__1449_, data_stage_5__1448_, data_stage_5__1447_, data_stage_5__1446_, data_stage_5__1445_, data_stage_5__1444_, data_stage_5__1443_, data_stage_5__1442_, data_stage_5__1441_, data_stage_5__1440_, data_stage_5__1439_, data_stage_5__1438_, data_stage_5__1437_, data_stage_5__1436_, data_stage_5__1435_, data_stage_5__1434_, data_stage_5__1433_, data_stage_5__1432_, data_stage_5__1431_, data_stage_5__1430_, data_stage_5__1429_, data_stage_5__1428_, data_stage_5__1427_, data_stage_5__1426_, data_stage_5__1425_, data_stage_5__1424_, data_stage_5__1423_, data_stage_5__1422_, data_stage_5__1421_, data_stage_5__1420_, data_stage_5__1419_, data_stage_5__1418_, data_stage_5__1417_, data_stage_5__1416_, data_stage_5__1415_, data_stage_5__1414_, data_stage_5__1413_, data_stage_5__1412_, data_stage_5__1411_, data_stage_5__1410_, data_stage_5__1409_, data_stage_5__1408_, data_stage_5__1407_, data_stage_5__1406_, data_stage_5__1405_, data_stage_5__1404_, data_stage_5__1403_, data_stage_5__1402_, data_stage_5__1401_, data_stage_5__1400_, data_stage_5__1399_, data_stage_5__1398_, data_stage_5__1397_, data_stage_5__1396_, data_stage_5__1395_, data_stage_5__1394_, data_stage_5__1393_, data_stage_5__1392_, data_stage_5__1391_, data_stage_5__1390_, data_stage_5__1389_, data_stage_5__1388_, data_stage_5__1387_, data_stage_5__1386_, data_stage_5__1385_, data_stage_5__1384_, data_stage_5__1383_, data_stage_5__1382_, data_stage_5__1381_, data_stage_5__1380_, data_stage_5__1379_, data_stage_5__1378_, data_stage_5__1377_, data_stage_5__1376_, data_stage_5__1375_, data_stage_5__1374_, data_stage_5__1373_, data_stage_5__1372_, data_stage_5__1371_, data_stage_5__1370_, data_stage_5__1369_, data_stage_5__1368_, data_stage_5__1367_, data_stage_5__1366_, data_stage_5__1365_, data_stage_5__1364_, data_stage_5__1363_, data_stage_5__1362_, data_stage_5__1361_, data_stage_5__1360_, data_stage_5__1359_, data_stage_5__1358_, data_stage_5__1357_, data_stage_5__1356_, data_stage_5__1355_, data_stage_5__1354_, data_stage_5__1353_, data_stage_5__1352_, data_stage_5__1351_, data_stage_5__1350_, data_stage_5__1349_, data_stage_5__1348_, data_stage_5__1347_, data_stage_5__1346_, data_stage_5__1345_, data_stage_5__1344_, data_stage_5__1343_, data_stage_5__1342_, data_stage_5__1341_, data_stage_5__1340_, data_stage_5__1339_, data_stage_5__1338_, data_stage_5__1337_, data_stage_5__1336_, data_stage_5__1335_, data_stage_5__1334_, data_stage_5__1333_, data_stage_5__1332_, data_stage_5__1331_, data_stage_5__1330_, data_stage_5__1329_, data_stage_5__1328_, data_stage_5__1327_, data_stage_5__1326_, data_stage_5__1325_, data_stage_5__1324_, data_stage_5__1323_, data_stage_5__1322_, data_stage_5__1321_, data_stage_5__1320_, data_stage_5__1319_, data_stage_5__1318_, data_stage_5__1317_, data_stage_5__1316_, data_stage_5__1315_, data_stage_5__1314_, data_stage_5__1313_, data_stage_5__1312_, data_stage_5__1311_, data_stage_5__1310_, data_stage_5__1309_, data_stage_5__1308_, data_stage_5__1307_, data_stage_5__1306_, data_stage_5__1305_, data_stage_5__1304_, data_stage_5__1303_, data_stage_5__1302_, data_stage_5__1301_, data_stage_5__1300_, data_stage_5__1299_, data_stage_5__1298_, data_stage_5__1297_, data_stage_5__1296_, data_stage_5__1295_, data_stage_5__1294_, data_stage_5__1293_, data_stage_5__1292_, data_stage_5__1291_, data_stage_5__1290_, data_stage_5__1289_, data_stage_5__1288_, data_stage_5__1287_, data_stage_5__1286_, data_stage_5__1285_, data_stage_5__1284_, data_stage_5__1283_, data_stage_5__1282_, data_stage_5__1281_, data_stage_5__1280_, data_stage_5__1279_, data_stage_5__1278_, data_stage_5__1277_, data_stage_5__1276_, data_stage_5__1275_, data_stage_5__1274_, data_stage_5__1273_, data_stage_5__1272_, data_stage_5__1271_, data_stage_5__1270_, data_stage_5__1269_, data_stage_5__1268_, data_stage_5__1267_, data_stage_5__1266_, data_stage_5__1265_, data_stage_5__1264_, data_stage_5__1263_, data_stage_5__1262_, data_stage_5__1261_, data_stage_5__1260_, data_stage_5__1259_, data_stage_5__1258_, data_stage_5__1257_, data_stage_5__1256_, data_stage_5__1255_, data_stage_5__1254_, data_stage_5__1253_, data_stage_5__1252_, data_stage_5__1251_, data_stage_5__1250_, data_stage_5__1249_, data_stage_5__1248_, data_stage_5__1247_, data_stage_5__1246_, data_stage_5__1245_, data_stage_5__1244_, data_stage_5__1243_, data_stage_5__1242_, data_stage_5__1241_, data_stage_5__1240_, data_stage_5__1239_, data_stage_5__1238_, data_stage_5__1237_, data_stage_5__1236_, data_stage_5__1235_, data_stage_5__1234_, data_stage_5__1233_, data_stage_5__1232_, data_stage_5__1231_, data_stage_5__1230_, data_stage_5__1229_, data_stage_5__1228_, data_stage_5__1227_, data_stage_5__1226_, data_stage_5__1225_, data_stage_5__1224_, data_stage_5__1223_, data_stage_5__1222_, data_stage_5__1221_, data_stage_5__1220_, data_stage_5__1219_, data_stage_5__1218_, data_stage_5__1217_, data_stage_5__1216_, data_stage_5__1215_, data_stage_5__1214_, data_stage_5__1213_, data_stage_5__1212_, data_stage_5__1211_, data_stage_5__1210_, data_stage_5__1209_, data_stage_5__1208_, data_stage_5__1207_, data_stage_5__1206_, data_stage_5__1205_, data_stage_5__1204_, data_stage_5__1203_, data_stage_5__1202_, data_stage_5__1201_, data_stage_5__1200_, data_stage_5__1199_, data_stage_5__1198_, data_stage_5__1197_, data_stage_5__1196_, data_stage_5__1195_, data_stage_5__1194_, data_stage_5__1193_, data_stage_5__1192_, data_stage_5__1191_, data_stage_5__1190_, data_stage_5__1189_, data_stage_5__1188_, data_stage_5__1187_, data_stage_5__1186_, data_stage_5__1185_, data_stage_5__1184_, data_stage_5__1183_, data_stage_5__1182_, data_stage_5__1181_, data_stage_5__1180_, data_stage_5__1179_, data_stage_5__1178_, data_stage_5__1177_, data_stage_5__1176_, data_stage_5__1175_, data_stage_5__1174_, data_stage_5__1173_, data_stage_5__1172_, data_stage_5__1171_, data_stage_5__1170_, data_stage_5__1169_, data_stage_5__1168_, data_stage_5__1167_, data_stage_5__1166_, data_stage_5__1165_, data_stage_5__1164_, data_stage_5__1163_, data_stage_5__1162_, data_stage_5__1161_, data_stage_5__1160_, data_stage_5__1159_, data_stage_5__1158_, data_stage_5__1157_, data_stage_5__1156_, data_stage_5__1155_, data_stage_5__1154_, data_stage_5__1153_, data_stage_5__1152_, data_stage_5__1151_, data_stage_5__1150_, data_stage_5__1149_, data_stage_5__1148_, data_stage_5__1147_, data_stage_5__1146_, data_stage_5__1145_, data_stage_5__1144_, data_stage_5__1143_, data_stage_5__1142_, data_stage_5__1141_, data_stage_5__1140_, data_stage_5__1139_, data_stage_5__1138_, data_stage_5__1137_, data_stage_5__1136_, data_stage_5__1135_, data_stage_5__1134_, data_stage_5__1133_, data_stage_5__1132_, data_stage_5__1131_, data_stage_5__1130_, data_stage_5__1129_, data_stage_5__1128_, data_stage_5__1127_, data_stage_5__1126_, data_stage_5__1125_, data_stage_5__1124_, data_stage_5__1123_, data_stage_5__1122_, data_stage_5__1121_, data_stage_5__1120_, data_stage_5__1119_, data_stage_5__1118_, data_stage_5__1117_, data_stage_5__1116_, data_stage_5__1115_, data_stage_5__1114_, data_stage_5__1113_, data_stage_5__1112_, data_stage_5__1111_, data_stage_5__1110_, data_stage_5__1109_, data_stage_5__1108_, data_stage_5__1107_, data_stage_5__1106_, data_stage_5__1105_, data_stage_5__1104_, data_stage_5__1103_, data_stage_5__1102_, data_stage_5__1101_, data_stage_5__1100_, data_stage_5__1099_, data_stage_5__1098_, data_stage_5__1097_, data_stage_5__1096_, data_stage_5__1095_, data_stage_5__1094_, data_stage_5__1093_, data_stage_5__1092_, data_stage_5__1091_, data_stage_5__1090_, data_stage_5__1089_, data_stage_5__1088_, data_stage_5__1087_, data_stage_5__1086_, data_stage_5__1085_, data_stage_5__1084_, data_stage_5__1083_, data_stage_5__1082_, data_stage_5__1081_, data_stage_5__1080_, data_stage_5__1079_, data_stage_5__1078_, data_stage_5__1077_, data_stage_5__1076_, data_stage_5__1075_, data_stage_5__1074_, data_stage_5__1073_, data_stage_5__1072_, data_stage_5__1071_, data_stage_5__1070_, data_stage_5__1069_, data_stage_5__1068_, data_stage_5__1067_, data_stage_5__1066_, data_stage_5__1065_, data_stage_5__1064_, data_stage_5__1063_, data_stage_5__1062_, data_stage_5__1061_, data_stage_5__1060_, data_stage_5__1059_, data_stage_5__1058_, data_stage_5__1057_, data_stage_5__1056_, data_stage_5__1055_, data_stage_5__1054_, data_stage_5__1053_, data_stage_5__1052_, data_stage_5__1051_, data_stage_5__1050_, data_stage_5__1049_, data_stage_5__1048_, data_stage_5__1047_, data_stage_5__1046_, data_stage_5__1045_, data_stage_5__1044_, data_stage_5__1043_, data_stage_5__1042_, data_stage_5__1041_, data_stage_5__1040_, data_stage_5__1039_, data_stage_5__1038_, data_stage_5__1037_, data_stage_5__1036_, data_stage_5__1035_, data_stage_5__1034_, data_stage_5__1033_, data_stage_5__1032_, data_stage_5__1031_, data_stage_5__1030_, data_stage_5__1029_, data_stage_5__1028_, data_stage_5__1027_, data_stage_5__1026_, data_stage_5__1025_, data_stage_5__1024_, data_stage_5__1023_, data_stage_5__1022_, data_stage_5__1021_, data_stage_5__1020_, data_stage_5__1019_, data_stage_5__1018_, data_stage_5__1017_, data_stage_5__1016_, data_stage_5__1015_, data_stage_5__1014_, data_stage_5__1013_, data_stage_5__1012_, data_stage_5__1011_, data_stage_5__1010_, data_stage_5__1009_, data_stage_5__1008_, data_stage_5__1007_, data_stage_5__1006_, data_stage_5__1005_, data_stage_5__1004_, data_stage_5__1003_, data_stage_5__1002_, data_stage_5__1001_, data_stage_5__1000_, data_stage_5__999_, data_stage_5__998_, data_stage_5__997_, data_stage_5__996_, data_stage_5__995_, data_stage_5__994_, data_stage_5__993_, data_stage_5__992_, data_stage_5__991_, data_stage_5__990_, data_stage_5__989_, data_stage_5__988_, data_stage_5__987_, data_stage_5__986_, data_stage_5__985_, data_stage_5__984_, data_stage_5__983_, data_stage_5__982_, data_stage_5__981_, data_stage_5__980_, data_stage_5__979_, data_stage_5__978_, data_stage_5__977_, data_stage_5__976_, data_stage_5__975_, data_stage_5__974_, data_stage_5__973_, data_stage_5__972_, data_stage_5__971_, data_stage_5__970_, data_stage_5__969_, data_stage_5__968_, data_stage_5__967_, data_stage_5__966_, data_stage_5__965_, data_stage_5__964_, data_stage_5__963_, data_stage_5__962_, data_stage_5__961_, data_stage_5__960_, data_stage_5__959_, data_stage_5__958_, data_stage_5__957_, data_stage_5__956_, data_stage_5__955_, data_stage_5__954_, data_stage_5__953_, data_stage_5__952_, data_stage_5__951_, data_stage_5__950_, data_stage_5__949_, data_stage_5__948_, data_stage_5__947_, data_stage_5__946_, data_stage_5__945_, data_stage_5__944_, data_stage_5__943_, data_stage_5__942_, data_stage_5__941_, data_stage_5__940_, data_stage_5__939_, data_stage_5__938_, data_stage_5__937_, data_stage_5__936_, data_stage_5__935_, data_stage_5__934_, data_stage_5__933_, data_stage_5__932_, data_stage_5__931_, data_stage_5__930_, data_stage_5__929_, data_stage_5__928_, data_stage_5__927_, data_stage_5__926_, data_stage_5__925_, data_stage_5__924_, data_stage_5__923_, data_stage_5__922_, data_stage_5__921_, data_stage_5__920_, data_stage_5__919_, data_stage_5__918_, data_stage_5__917_, data_stage_5__916_, data_stage_5__915_, data_stage_5__914_, data_stage_5__913_, data_stage_5__912_, data_stage_5__911_, data_stage_5__910_, data_stage_5__909_, data_stage_5__908_, data_stage_5__907_, data_stage_5__906_, data_stage_5__905_, data_stage_5__904_, data_stage_5__903_, data_stage_5__902_, data_stage_5__901_, data_stage_5__900_, data_stage_5__899_, data_stage_5__898_, data_stage_5__897_, data_stage_5__896_, data_stage_5__895_, data_stage_5__894_, data_stage_5__893_, data_stage_5__892_, data_stage_5__891_, data_stage_5__890_, data_stage_5__889_, data_stage_5__888_, data_stage_5__887_, data_stage_5__886_, data_stage_5__885_, data_stage_5__884_, data_stage_5__883_, data_stage_5__882_, data_stage_5__881_, data_stage_5__880_, data_stage_5__879_, data_stage_5__878_, data_stage_5__877_, data_stage_5__876_, data_stage_5__875_, data_stage_5__874_, data_stage_5__873_, data_stage_5__872_, data_stage_5__871_, data_stage_5__870_, data_stage_5__869_, data_stage_5__868_, data_stage_5__867_, data_stage_5__866_, data_stage_5__865_, data_stage_5__864_, data_stage_5__863_, data_stage_5__862_, data_stage_5__861_, data_stage_5__860_, data_stage_5__859_, data_stage_5__858_, data_stage_5__857_, data_stage_5__856_, data_stage_5__855_, data_stage_5__854_, data_stage_5__853_, data_stage_5__852_, data_stage_5__851_, data_stage_5__850_, data_stage_5__849_, data_stage_5__848_, data_stage_5__847_, data_stage_5__846_, data_stage_5__845_, data_stage_5__844_, data_stage_5__843_, data_stage_5__842_, data_stage_5__841_, data_stage_5__840_, data_stage_5__839_, data_stage_5__838_, data_stage_5__837_, data_stage_5__836_, data_stage_5__835_, data_stage_5__834_, data_stage_5__833_, data_stage_5__832_, data_stage_5__831_, data_stage_5__830_, data_stage_5__829_, data_stage_5__828_, data_stage_5__827_, data_stage_5__826_, data_stage_5__825_, data_stage_5__824_, data_stage_5__823_, data_stage_5__822_, data_stage_5__821_, data_stage_5__820_, data_stage_5__819_, data_stage_5__818_, data_stage_5__817_, data_stage_5__816_, data_stage_5__815_, data_stage_5__814_, data_stage_5__813_, data_stage_5__812_, data_stage_5__811_, data_stage_5__810_, data_stage_5__809_, data_stage_5__808_, data_stage_5__807_, data_stage_5__806_, data_stage_5__805_, data_stage_5__804_, data_stage_5__803_, data_stage_5__802_, data_stage_5__801_, data_stage_5__800_, data_stage_5__799_, data_stage_5__798_, data_stage_5__797_, data_stage_5__796_, data_stage_5__795_, data_stage_5__794_, data_stage_5__793_, data_stage_5__792_, data_stage_5__791_, data_stage_5__790_, data_stage_5__789_, data_stage_5__788_, data_stage_5__787_, data_stage_5__786_, data_stage_5__785_, data_stage_5__784_, data_stage_5__783_, data_stage_5__782_, data_stage_5__781_, data_stage_5__780_, data_stage_5__779_, data_stage_5__778_, data_stage_5__777_, data_stage_5__776_, data_stage_5__775_, data_stage_5__774_, data_stage_5__773_, data_stage_5__772_, data_stage_5__771_, data_stage_5__770_, data_stage_5__769_, data_stage_5__768_, data_stage_5__767_, data_stage_5__766_, data_stage_5__765_, data_stage_5__764_, data_stage_5__763_, data_stage_5__762_, data_stage_5__761_, data_stage_5__760_, data_stage_5__759_, data_stage_5__758_, data_stage_5__757_, data_stage_5__756_, data_stage_5__755_, data_stage_5__754_, data_stage_5__753_, data_stage_5__752_, data_stage_5__751_, data_stage_5__750_, data_stage_5__749_, data_stage_5__748_, data_stage_5__747_, data_stage_5__746_, data_stage_5__745_, data_stage_5__744_, data_stage_5__743_, data_stage_5__742_, data_stage_5__741_, data_stage_5__740_, data_stage_5__739_, data_stage_5__738_, data_stage_5__737_, data_stage_5__736_, data_stage_5__735_, data_stage_5__734_, data_stage_5__733_, data_stage_5__732_, data_stage_5__731_, data_stage_5__730_, data_stage_5__729_, data_stage_5__728_, data_stage_5__727_, data_stage_5__726_, data_stage_5__725_, data_stage_5__724_, data_stage_5__723_, data_stage_5__722_, data_stage_5__721_, data_stage_5__720_, data_stage_5__719_, data_stage_5__718_, data_stage_5__717_, data_stage_5__716_, data_stage_5__715_, data_stage_5__714_, data_stage_5__713_, data_stage_5__712_, data_stage_5__711_, data_stage_5__710_, data_stage_5__709_, data_stage_5__708_, data_stage_5__707_, data_stage_5__706_, data_stage_5__705_, data_stage_5__704_, data_stage_5__703_, data_stage_5__702_, data_stage_5__701_, data_stage_5__700_, data_stage_5__699_, data_stage_5__698_, data_stage_5__697_, data_stage_5__696_, data_stage_5__695_, data_stage_5__694_, data_stage_5__693_, data_stage_5__692_, data_stage_5__691_, data_stage_5__690_, data_stage_5__689_, data_stage_5__688_, data_stage_5__687_, data_stage_5__686_, data_stage_5__685_, data_stage_5__684_, data_stage_5__683_, data_stage_5__682_, data_stage_5__681_, data_stage_5__680_, data_stage_5__679_, data_stage_5__678_, data_stage_5__677_, data_stage_5__676_, data_stage_5__675_, data_stage_5__674_, data_stage_5__673_, data_stage_5__672_, data_stage_5__671_, data_stage_5__670_, data_stage_5__669_, data_stage_5__668_, data_stage_5__667_, data_stage_5__666_, data_stage_5__665_, data_stage_5__664_, data_stage_5__663_, data_stage_5__662_, data_stage_5__661_, data_stage_5__660_, data_stage_5__659_, data_stage_5__658_, data_stage_5__657_, data_stage_5__656_, data_stage_5__655_, data_stage_5__654_, data_stage_5__653_, data_stage_5__652_, data_stage_5__651_, data_stage_5__650_, data_stage_5__649_, data_stage_5__648_, data_stage_5__647_, data_stage_5__646_, data_stage_5__645_, data_stage_5__644_, data_stage_5__643_, data_stage_5__642_, data_stage_5__641_, data_stage_5__640_, data_stage_5__639_, data_stage_5__638_, data_stage_5__637_, data_stage_5__636_, data_stage_5__635_, data_stage_5__634_, data_stage_5__633_, data_stage_5__632_, data_stage_5__631_, data_stage_5__630_, data_stage_5__629_, data_stage_5__628_, data_stage_5__627_, data_stage_5__626_, data_stage_5__625_, data_stage_5__624_, data_stage_5__623_, data_stage_5__622_, data_stage_5__621_, data_stage_5__620_, data_stage_5__619_, data_stage_5__618_, data_stage_5__617_, data_stage_5__616_, data_stage_5__615_, data_stage_5__614_, data_stage_5__613_, data_stage_5__612_, data_stage_5__611_, data_stage_5__610_, data_stage_5__609_, data_stage_5__608_, data_stage_5__607_, data_stage_5__606_, data_stage_5__605_, data_stage_5__604_, data_stage_5__603_, data_stage_5__602_, data_stage_5__601_, data_stage_5__600_, data_stage_5__599_, data_stage_5__598_, data_stage_5__597_, data_stage_5__596_, data_stage_5__595_, data_stage_5__594_, data_stage_5__593_, data_stage_5__592_, data_stage_5__591_, data_stage_5__590_, data_stage_5__589_, data_stage_5__588_, data_stage_5__587_, data_stage_5__586_, data_stage_5__585_, data_stage_5__584_, data_stage_5__583_, data_stage_5__582_, data_stage_5__581_, data_stage_5__580_, data_stage_5__579_, data_stage_5__578_, data_stage_5__577_, data_stage_5__576_, data_stage_5__575_, data_stage_5__574_, data_stage_5__573_, data_stage_5__572_, data_stage_5__571_, data_stage_5__570_, data_stage_5__569_, data_stage_5__568_, data_stage_5__567_, data_stage_5__566_, data_stage_5__565_, data_stage_5__564_, data_stage_5__563_, data_stage_5__562_, data_stage_5__561_, data_stage_5__560_, data_stage_5__559_, data_stage_5__558_, data_stage_5__557_, data_stage_5__556_, data_stage_5__555_, data_stage_5__554_, data_stage_5__553_, data_stage_5__552_, data_stage_5__551_, data_stage_5__550_, data_stage_5__549_, data_stage_5__548_, data_stage_5__547_, data_stage_5__546_, data_stage_5__545_, data_stage_5__544_, data_stage_5__543_, data_stage_5__542_, data_stage_5__541_, data_stage_5__540_, data_stage_5__539_, data_stage_5__538_, data_stage_5__537_, data_stage_5__536_, data_stage_5__535_, data_stage_5__534_, data_stage_5__533_, data_stage_5__532_, data_stage_5__531_, data_stage_5__530_, data_stage_5__529_, data_stage_5__528_, data_stage_5__527_, data_stage_5__526_, data_stage_5__525_, data_stage_5__524_, data_stage_5__523_, data_stage_5__522_, data_stage_5__521_, data_stage_5__520_, data_stage_5__519_, data_stage_5__518_, data_stage_5__517_, data_stage_5__516_, data_stage_5__515_, data_stage_5__514_, data_stage_5__513_, data_stage_5__512_, data_stage_5__511_, data_stage_5__510_, data_stage_5__509_, data_stage_5__508_, data_stage_5__507_, data_stage_5__506_, data_stage_5__505_, data_stage_5__504_, data_stage_5__503_, data_stage_5__502_, data_stage_5__501_, data_stage_5__500_, data_stage_5__499_, data_stage_5__498_, data_stage_5__497_, data_stage_5__496_, data_stage_5__495_, data_stage_5__494_, data_stage_5__493_, data_stage_5__492_, data_stage_5__491_, data_stage_5__490_, data_stage_5__489_, data_stage_5__488_, data_stage_5__487_, data_stage_5__486_, data_stage_5__485_, data_stage_5__484_, data_stage_5__483_, data_stage_5__482_, data_stage_5__481_, data_stage_5__480_, data_stage_5__479_, data_stage_5__478_, data_stage_5__477_, data_stage_5__476_, data_stage_5__475_, data_stage_5__474_, data_stage_5__473_, data_stage_5__472_, data_stage_5__471_, data_stage_5__470_, data_stage_5__469_, data_stage_5__468_, data_stage_5__467_, data_stage_5__466_, data_stage_5__465_, data_stage_5__464_, data_stage_5__463_, data_stage_5__462_, data_stage_5__461_, data_stage_5__460_, data_stage_5__459_, data_stage_5__458_, data_stage_5__457_, data_stage_5__456_, data_stage_5__455_, data_stage_5__454_, data_stage_5__453_, data_stage_5__452_, data_stage_5__451_, data_stage_5__450_, data_stage_5__449_, data_stage_5__448_, data_stage_5__447_, data_stage_5__446_, data_stage_5__445_, data_stage_5__444_, data_stage_5__443_, data_stage_5__442_, data_stage_5__441_, data_stage_5__440_, data_stage_5__439_, data_stage_5__438_, data_stage_5__437_, data_stage_5__436_, data_stage_5__435_, data_stage_5__434_, data_stage_5__433_, data_stage_5__432_, data_stage_5__431_, data_stage_5__430_, data_stage_5__429_, data_stage_5__428_, data_stage_5__427_, data_stage_5__426_, data_stage_5__425_, data_stage_5__424_, data_stage_5__423_, data_stage_5__422_, data_stage_5__421_, data_stage_5__420_, data_stage_5__419_, data_stage_5__418_, data_stage_5__417_, data_stage_5__416_, data_stage_5__415_, data_stage_5__414_, data_stage_5__413_, data_stage_5__412_, data_stage_5__411_, data_stage_5__410_, data_stage_5__409_, data_stage_5__408_, data_stage_5__407_, data_stage_5__406_, data_stage_5__405_, data_stage_5__404_, data_stage_5__403_, data_stage_5__402_, data_stage_5__401_, data_stage_5__400_, data_stage_5__399_, data_stage_5__398_, data_stage_5__397_, data_stage_5__396_, data_stage_5__395_, data_stage_5__394_, data_stage_5__393_, data_stage_5__392_, data_stage_5__391_, data_stage_5__390_, data_stage_5__389_, data_stage_5__388_, data_stage_5__387_, data_stage_5__386_, data_stage_5__385_, data_stage_5__384_, data_stage_5__383_, data_stage_5__382_, data_stage_5__381_, data_stage_5__380_, data_stage_5__379_, data_stage_5__378_, data_stage_5__377_, data_stage_5__376_, data_stage_5__375_, data_stage_5__374_, data_stage_5__373_, data_stage_5__372_, data_stage_5__371_, data_stage_5__370_, data_stage_5__369_, data_stage_5__368_, data_stage_5__367_, data_stage_5__366_, data_stage_5__365_, data_stage_5__364_, data_stage_5__363_, data_stage_5__362_, data_stage_5__361_, data_stage_5__360_, data_stage_5__359_, data_stage_5__358_, data_stage_5__357_, data_stage_5__356_, data_stage_5__355_, data_stage_5__354_, data_stage_5__353_, data_stage_5__352_, data_stage_5__351_, data_stage_5__350_, data_stage_5__349_, data_stage_5__348_, data_stage_5__347_, data_stage_5__346_, data_stage_5__345_, data_stage_5__344_, data_stage_5__343_, data_stage_5__342_, data_stage_5__341_, data_stage_5__340_, data_stage_5__339_, data_stage_5__338_, data_stage_5__337_, data_stage_5__336_, data_stage_5__335_, data_stage_5__334_, data_stage_5__333_, data_stage_5__332_, data_stage_5__331_, data_stage_5__330_, data_stage_5__329_, data_stage_5__328_, data_stage_5__327_, data_stage_5__326_, data_stage_5__325_, data_stage_5__324_, data_stage_5__323_, data_stage_5__322_, data_stage_5__321_, data_stage_5__320_, data_stage_5__319_, data_stage_5__318_, data_stage_5__317_, data_stage_5__316_, data_stage_5__315_, data_stage_5__314_, data_stage_5__313_, data_stage_5__312_, data_stage_5__311_, data_stage_5__310_, data_stage_5__309_, data_stage_5__308_, data_stage_5__307_, data_stage_5__306_, data_stage_5__305_, data_stage_5__304_, data_stage_5__303_, data_stage_5__302_, data_stage_5__301_, data_stage_5__300_, data_stage_5__299_, data_stage_5__298_, data_stage_5__297_, data_stage_5__296_, data_stage_5__295_, data_stage_5__294_, data_stage_5__293_, data_stage_5__292_, data_stage_5__291_, data_stage_5__290_, data_stage_5__289_, data_stage_5__288_, data_stage_5__287_, data_stage_5__286_, data_stage_5__285_, data_stage_5__284_, data_stage_5__283_, data_stage_5__282_, data_stage_5__281_, data_stage_5__280_, data_stage_5__279_, data_stage_5__278_, data_stage_5__277_, data_stage_5__276_, data_stage_5__275_, data_stage_5__274_, data_stage_5__273_, data_stage_5__272_, data_stage_5__271_, data_stage_5__270_, data_stage_5__269_, data_stage_5__268_, data_stage_5__267_, data_stage_5__266_, data_stage_5__265_, data_stage_5__264_, data_stage_5__263_, data_stage_5__262_, data_stage_5__261_, data_stage_5__260_, data_stage_5__259_, data_stage_5__258_, data_stage_5__257_, data_stage_5__256_, data_stage_5__255_, data_stage_5__254_, data_stage_5__253_, data_stage_5__252_, data_stage_5__251_, data_stage_5__250_, data_stage_5__249_, data_stage_5__248_, data_stage_5__247_, data_stage_5__246_, data_stage_5__245_, data_stage_5__244_, data_stage_5__243_, data_stage_5__242_, data_stage_5__241_, data_stage_5__240_, data_stage_5__239_, data_stage_5__238_, data_stage_5__237_, data_stage_5__236_, data_stage_5__235_, data_stage_5__234_, data_stage_5__233_, data_stage_5__232_, data_stage_5__231_, data_stage_5__230_, data_stage_5__229_, data_stage_5__228_, data_stage_5__227_, data_stage_5__226_, data_stage_5__225_, data_stage_5__224_, data_stage_5__223_, data_stage_5__222_, data_stage_5__221_, data_stage_5__220_, data_stage_5__219_, data_stage_5__218_, data_stage_5__217_, data_stage_5__216_, data_stage_5__215_, data_stage_5__214_, data_stage_5__213_, data_stage_5__212_, data_stage_5__211_, data_stage_5__210_, data_stage_5__209_, data_stage_5__208_, data_stage_5__207_, data_stage_5__206_, data_stage_5__205_, data_stage_5__204_, data_stage_5__203_, data_stage_5__202_, data_stage_5__201_, data_stage_5__200_, data_stage_5__199_, data_stage_5__198_, data_stage_5__197_, data_stage_5__196_, data_stage_5__195_, data_stage_5__194_, data_stage_5__193_, data_stage_5__192_, data_stage_5__191_, data_stage_5__190_, data_stage_5__189_, data_stage_5__188_, data_stage_5__187_, data_stage_5__186_, data_stage_5__185_, data_stage_5__184_, data_stage_5__183_, data_stage_5__182_, data_stage_5__181_, data_stage_5__180_, data_stage_5__179_, data_stage_5__178_, data_stage_5__177_, data_stage_5__176_, data_stage_5__175_, data_stage_5__174_, data_stage_5__173_, data_stage_5__172_, data_stage_5__171_, data_stage_5__170_, data_stage_5__169_, data_stage_5__168_, data_stage_5__167_, data_stage_5__166_, data_stage_5__165_, data_stage_5__164_, data_stage_5__163_, data_stage_5__162_, data_stage_5__161_, data_stage_5__160_, data_stage_5__159_, data_stage_5__158_, data_stage_5__157_, data_stage_5__156_, data_stage_5__155_, data_stage_5__154_, data_stage_5__153_, data_stage_5__152_, data_stage_5__151_, data_stage_5__150_, data_stage_5__149_, data_stage_5__148_, data_stage_5__147_, data_stage_5__146_, data_stage_5__145_, data_stage_5__144_, data_stage_5__143_, data_stage_5__142_, data_stage_5__141_, data_stage_5__140_, data_stage_5__139_, data_stage_5__138_, data_stage_5__137_, data_stage_5__136_, data_stage_5__135_, data_stage_5__134_, data_stage_5__133_, data_stage_5__132_, data_stage_5__131_, data_stage_5__130_, data_stage_5__129_, data_stage_5__128_, data_stage_5__127_, data_stage_5__126_, data_stage_5__125_, data_stage_5__124_, data_stage_5__123_, data_stage_5__122_, data_stage_5__121_, data_stage_5__120_, data_stage_5__119_, data_stage_5__118_, data_stage_5__117_, data_stage_5__116_, data_stage_5__115_, data_stage_5__114_, data_stage_5__113_, data_stage_5__112_, data_stage_5__111_, data_stage_5__110_, data_stage_5__109_, data_stage_5__108_, data_stage_5__107_, data_stage_5__106_, data_stage_5__105_, data_stage_5__104_, data_stage_5__103_, data_stage_5__102_, data_stage_5__101_, data_stage_5__100_, data_stage_5__99_, data_stage_5__98_, data_stage_5__97_, data_stage_5__96_, data_stage_5__95_, data_stage_5__94_, data_stage_5__93_, data_stage_5__92_, data_stage_5__91_, data_stage_5__90_, data_stage_5__89_, data_stage_5__88_, data_stage_5__87_, data_stage_5__86_, data_stage_5__85_, data_stage_5__84_, data_stage_5__83_, data_stage_5__82_, data_stage_5__81_, data_stage_5__80_, data_stage_5__79_, data_stage_5__78_, data_stage_5__77_, data_stage_5__76_, data_stage_5__75_, data_stage_5__74_, data_stage_5__73_, data_stage_5__72_, data_stage_5__71_, data_stage_5__70_, data_stage_5__69_, data_stage_5__68_, data_stage_5__67_, data_stage_5__66_, data_stage_5__65_, data_stage_5__64_, data_stage_5__63_, data_stage_5__62_, data_stage_5__61_, data_stage_5__60_, data_stage_5__59_, data_stage_5__58_, data_stage_5__57_, data_stage_5__56_, data_stage_5__55_, data_stage_5__54_, data_stage_5__53_, data_stage_5__52_, data_stage_5__51_, data_stage_5__50_, data_stage_5__49_, data_stage_5__48_, data_stage_5__47_, data_stage_5__46_, data_stage_5__45_, data_stage_5__44_, data_stage_5__43_, data_stage_5__42_, data_stage_5__41_, data_stage_5__40_, data_stage_5__39_, data_stage_5__38_, data_stage_5__37_, data_stage_5__36_, data_stage_5__35_, data_stage_5__34_, data_stage_5__33_, data_stage_5__32_, data_stage_5__31_, data_stage_5__30_, data_stage_5__29_, data_stage_5__28_, data_stage_5__27_, data_stage_5__26_, data_stage_5__25_, data_stage_5__24_, data_stage_5__23_, data_stage_5__22_, data_stage_5__21_, data_stage_5__20_, data_stage_5__19_, data_stage_5__18_, data_stage_5__17_, data_stage_5__16_, data_stage_5__15_, data_stage_5__14_, data_stage_5__13_, data_stage_5__12_, data_stage_5__11_, data_stage_5__10_, data_stage_5__9_, data_stage_5__8_, data_stage_5__7_, data_stage_5__6_, data_stage_5__5_, data_stage_5__4_, data_stage_5__3_, data_stage_5__2_, data_stage_5__1_, data_stage_5__0_ }),
    .swap_i(sel_i[5]),
    .data_o(data_o)
  );


endmodule

