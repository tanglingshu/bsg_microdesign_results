

module top
(
  clk_i,
  reset_i,
  v_i,
  len_i,
  data_i,
  ready_o,
  v_o,
  len_v_o,
  data_o,
  yumi_i
);

  input [5:0] len_i;
  input [1599:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  output len_v_o;

  bsg_parallel_in_serial_out_dynamic
  wrapper
  (
    .len_i(len_i),
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_i(yumi_i),
    .ready_o(ready_o),
    .v_o(v_o),
    .len_v_o(len_v_o)
  );


endmodule



module bsg_mem_1r1w_synth_width_p6_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [5:0] w_data_i;
  input [0:0] r_addr_i;
  output [5:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [5:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8;
  reg [11:0] mem;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[11] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[10] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[9] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[8] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[7] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[6] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N8, N7 } = (N1)? { w_addr_i[0:0], N5 } : 
                      (N2)? { 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N8) begin
      { mem[11:6] } <= { w_data_i[5:0] };
    end 
    if(N7) begin
      { mem[5:0] } <= { w_data_i[5:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p6_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [5:0] w_data_i;
  input [0:0] r_addr_i;
  output [5:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [5:0] r_data_o;

  bsg_mem_1r1w_synth_width_p6_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p6
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [5:0] data_i;
  output [5:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [5:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p6_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bsg_mem_1r1w_synth_width_p1600_els_p2_read_write_same_addr_p0_harden_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [1599:0] w_data_i;
  input [0:0] r_addr_i;
  output [1599:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [1599:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,N22,
  N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38;
  reg [3199:0] mem;
  assign r_data_o[1599] = (N3)? mem[1599] : 
                          (N0)? mem[3199] : 1'b0;
  assign N0 = r_addr_i[0];
  assign r_data_o[1598] = (N3)? mem[1598] : 
                          (N0)? mem[3198] : 1'b0;
  assign r_data_o[1597] = (N3)? mem[1597] : 
                          (N0)? mem[3197] : 1'b0;
  assign r_data_o[1596] = (N3)? mem[1596] : 
                          (N0)? mem[3196] : 1'b0;
  assign r_data_o[1595] = (N3)? mem[1595] : 
                          (N0)? mem[3195] : 1'b0;
  assign r_data_o[1594] = (N3)? mem[1594] : 
                          (N0)? mem[3194] : 1'b0;
  assign r_data_o[1593] = (N3)? mem[1593] : 
                          (N0)? mem[3193] : 1'b0;
  assign r_data_o[1592] = (N3)? mem[1592] : 
                          (N0)? mem[3192] : 1'b0;
  assign r_data_o[1591] = (N3)? mem[1591] : 
                          (N0)? mem[3191] : 1'b0;
  assign r_data_o[1590] = (N3)? mem[1590] : 
                          (N0)? mem[3190] : 1'b0;
  assign r_data_o[1589] = (N3)? mem[1589] : 
                          (N0)? mem[3189] : 1'b0;
  assign r_data_o[1588] = (N3)? mem[1588] : 
                          (N0)? mem[3188] : 1'b0;
  assign r_data_o[1587] = (N3)? mem[1587] : 
                          (N0)? mem[3187] : 1'b0;
  assign r_data_o[1586] = (N3)? mem[1586] : 
                          (N0)? mem[3186] : 1'b0;
  assign r_data_o[1585] = (N3)? mem[1585] : 
                          (N0)? mem[3185] : 1'b0;
  assign r_data_o[1584] = (N3)? mem[1584] : 
                          (N0)? mem[3184] : 1'b0;
  assign r_data_o[1583] = (N3)? mem[1583] : 
                          (N0)? mem[3183] : 1'b0;
  assign r_data_o[1582] = (N3)? mem[1582] : 
                          (N0)? mem[3182] : 1'b0;
  assign r_data_o[1581] = (N3)? mem[1581] : 
                          (N0)? mem[3181] : 1'b0;
  assign r_data_o[1580] = (N3)? mem[1580] : 
                          (N0)? mem[3180] : 1'b0;
  assign r_data_o[1579] = (N3)? mem[1579] : 
                          (N0)? mem[3179] : 1'b0;
  assign r_data_o[1578] = (N3)? mem[1578] : 
                          (N0)? mem[3178] : 1'b0;
  assign r_data_o[1577] = (N3)? mem[1577] : 
                          (N0)? mem[3177] : 1'b0;
  assign r_data_o[1576] = (N3)? mem[1576] : 
                          (N0)? mem[3176] : 1'b0;
  assign r_data_o[1575] = (N3)? mem[1575] : 
                          (N0)? mem[3175] : 1'b0;
  assign r_data_o[1574] = (N3)? mem[1574] : 
                          (N0)? mem[3174] : 1'b0;
  assign r_data_o[1573] = (N3)? mem[1573] : 
                          (N0)? mem[3173] : 1'b0;
  assign r_data_o[1572] = (N3)? mem[1572] : 
                          (N0)? mem[3172] : 1'b0;
  assign r_data_o[1571] = (N3)? mem[1571] : 
                          (N0)? mem[3171] : 1'b0;
  assign r_data_o[1570] = (N3)? mem[1570] : 
                          (N0)? mem[3170] : 1'b0;
  assign r_data_o[1569] = (N3)? mem[1569] : 
                          (N0)? mem[3169] : 1'b0;
  assign r_data_o[1568] = (N3)? mem[1568] : 
                          (N0)? mem[3168] : 1'b0;
  assign r_data_o[1567] = (N3)? mem[1567] : 
                          (N0)? mem[3167] : 1'b0;
  assign r_data_o[1566] = (N3)? mem[1566] : 
                          (N0)? mem[3166] : 1'b0;
  assign r_data_o[1565] = (N3)? mem[1565] : 
                          (N0)? mem[3165] : 1'b0;
  assign r_data_o[1564] = (N3)? mem[1564] : 
                          (N0)? mem[3164] : 1'b0;
  assign r_data_o[1563] = (N3)? mem[1563] : 
                          (N0)? mem[3163] : 1'b0;
  assign r_data_o[1562] = (N3)? mem[1562] : 
                          (N0)? mem[3162] : 1'b0;
  assign r_data_o[1561] = (N3)? mem[1561] : 
                          (N0)? mem[3161] : 1'b0;
  assign r_data_o[1560] = (N3)? mem[1560] : 
                          (N0)? mem[3160] : 1'b0;
  assign r_data_o[1559] = (N3)? mem[1559] : 
                          (N0)? mem[3159] : 1'b0;
  assign r_data_o[1558] = (N3)? mem[1558] : 
                          (N0)? mem[3158] : 1'b0;
  assign r_data_o[1557] = (N3)? mem[1557] : 
                          (N0)? mem[3157] : 1'b0;
  assign r_data_o[1556] = (N3)? mem[1556] : 
                          (N0)? mem[3156] : 1'b0;
  assign r_data_o[1555] = (N3)? mem[1555] : 
                          (N0)? mem[3155] : 1'b0;
  assign r_data_o[1554] = (N3)? mem[1554] : 
                          (N0)? mem[3154] : 1'b0;
  assign r_data_o[1553] = (N3)? mem[1553] : 
                          (N0)? mem[3153] : 1'b0;
  assign r_data_o[1552] = (N3)? mem[1552] : 
                          (N0)? mem[3152] : 1'b0;
  assign r_data_o[1551] = (N3)? mem[1551] : 
                          (N0)? mem[3151] : 1'b0;
  assign r_data_o[1550] = (N3)? mem[1550] : 
                          (N0)? mem[3150] : 1'b0;
  assign r_data_o[1549] = (N3)? mem[1549] : 
                          (N0)? mem[3149] : 1'b0;
  assign r_data_o[1548] = (N3)? mem[1548] : 
                          (N0)? mem[3148] : 1'b0;
  assign r_data_o[1547] = (N3)? mem[1547] : 
                          (N0)? mem[3147] : 1'b0;
  assign r_data_o[1546] = (N3)? mem[1546] : 
                          (N0)? mem[3146] : 1'b0;
  assign r_data_o[1545] = (N3)? mem[1545] : 
                          (N0)? mem[3145] : 1'b0;
  assign r_data_o[1544] = (N3)? mem[1544] : 
                          (N0)? mem[3144] : 1'b0;
  assign r_data_o[1543] = (N3)? mem[1543] : 
                          (N0)? mem[3143] : 1'b0;
  assign r_data_o[1542] = (N3)? mem[1542] : 
                          (N0)? mem[3142] : 1'b0;
  assign r_data_o[1541] = (N3)? mem[1541] : 
                          (N0)? mem[3141] : 1'b0;
  assign r_data_o[1540] = (N3)? mem[1540] : 
                          (N0)? mem[3140] : 1'b0;
  assign r_data_o[1539] = (N3)? mem[1539] : 
                          (N0)? mem[3139] : 1'b0;
  assign r_data_o[1538] = (N3)? mem[1538] : 
                          (N0)? mem[3138] : 1'b0;
  assign r_data_o[1537] = (N3)? mem[1537] : 
                          (N0)? mem[3137] : 1'b0;
  assign r_data_o[1536] = (N3)? mem[1536] : 
                          (N0)? mem[3136] : 1'b0;
  assign r_data_o[1535] = (N3)? mem[1535] : 
                          (N0)? mem[3135] : 1'b0;
  assign r_data_o[1534] = (N3)? mem[1534] : 
                          (N0)? mem[3134] : 1'b0;
  assign r_data_o[1533] = (N3)? mem[1533] : 
                          (N0)? mem[3133] : 1'b0;
  assign r_data_o[1532] = (N3)? mem[1532] : 
                          (N0)? mem[3132] : 1'b0;
  assign r_data_o[1531] = (N3)? mem[1531] : 
                          (N0)? mem[3131] : 1'b0;
  assign r_data_o[1530] = (N3)? mem[1530] : 
                          (N0)? mem[3130] : 1'b0;
  assign r_data_o[1529] = (N3)? mem[1529] : 
                          (N0)? mem[3129] : 1'b0;
  assign r_data_o[1528] = (N3)? mem[1528] : 
                          (N0)? mem[3128] : 1'b0;
  assign r_data_o[1527] = (N3)? mem[1527] : 
                          (N0)? mem[3127] : 1'b0;
  assign r_data_o[1526] = (N3)? mem[1526] : 
                          (N0)? mem[3126] : 1'b0;
  assign r_data_o[1525] = (N3)? mem[1525] : 
                          (N0)? mem[3125] : 1'b0;
  assign r_data_o[1524] = (N3)? mem[1524] : 
                          (N0)? mem[3124] : 1'b0;
  assign r_data_o[1523] = (N3)? mem[1523] : 
                          (N0)? mem[3123] : 1'b0;
  assign r_data_o[1522] = (N3)? mem[1522] : 
                          (N0)? mem[3122] : 1'b0;
  assign r_data_o[1521] = (N3)? mem[1521] : 
                          (N0)? mem[3121] : 1'b0;
  assign r_data_o[1520] = (N3)? mem[1520] : 
                          (N0)? mem[3120] : 1'b0;
  assign r_data_o[1519] = (N3)? mem[1519] : 
                          (N0)? mem[3119] : 1'b0;
  assign r_data_o[1518] = (N3)? mem[1518] : 
                          (N0)? mem[3118] : 1'b0;
  assign r_data_o[1517] = (N3)? mem[1517] : 
                          (N0)? mem[3117] : 1'b0;
  assign r_data_o[1516] = (N3)? mem[1516] : 
                          (N0)? mem[3116] : 1'b0;
  assign r_data_o[1515] = (N3)? mem[1515] : 
                          (N0)? mem[3115] : 1'b0;
  assign r_data_o[1514] = (N3)? mem[1514] : 
                          (N0)? mem[3114] : 1'b0;
  assign r_data_o[1513] = (N3)? mem[1513] : 
                          (N0)? mem[3113] : 1'b0;
  assign r_data_o[1512] = (N3)? mem[1512] : 
                          (N0)? mem[3112] : 1'b0;
  assign r_data_o[1511] = (N3)? mem[1511] : 
                          (N0)? mem[3111] : 1'b0;
  assign r_data_o[1510] = (N3)? mem[1510] : 
                          (N0)? mem[3110] : 1'b0;
  assign r_data_o[1509] = (N3)? mem[1509] : 
                          (N0)? mem[3109] : 1'b0;
  assign r_data_o[1508] = (N3)? mem[1508] : 
                          (N0)? mem[3108] : 1'b0;
  assign r_data_o[1507] = (N3)? mem[1507] : 
                          (N0)? mem[3107] : 1'b0;
  assign r_data_o[1506] = (N3)? mem[1506] : 
                          (N0)? mem[3106] : 1'b0;
  assign r_data_o[1505] = (N3)? mem[1505] : 
                          (N0)? mem[3105] : 1'b0;
  assign r_data_o[1504] = (N3)? mem[1504] : 
                          (N0)? mem[3104] : 1'b0;
  assign r_data_o[1503] = (N3)? mem[1503] : 
                          (N0)? mem[3103] : 1'b0;
  assign r_data_o[1502] = (N3)? mem[1502] : 
                          (N0)? mem[3102] : 1'b0;
  assign r_data_o[1501] = (N3)? mem[1501] : 
                          (N0)? mem[3101] : 1'b0;
  assign r_data_o[1500] = (N3)? mem[1500] : 
                          (N0)? mem[3100] : 1'b0;
  assign r_data_o[1499] = (N3)? mem[1499] : 
                          (N0)? mem[3099] : 1'b0;
  assign r_data_o[1498] = (N3)? mem[1498] : 
                          (N0)? mem[3098] : 1'b0;
  assign r_data_o[1497] = (N3)? mem[1497] : 
                          (N0)? mem[3097] : 1'b0;
  assign r_data_o[1496] = (N3)? mem[1496] : 
                          (N0)? mem[3096] : 1'b0;
  assign r_data_o[1495] = (N3)? mem[1495] : 
                          (N0)? mem[3095] : 1'b0;
  assign r_data_o[1494] = (N3)? mem[1494] : 
                          (N0)? mem[3094] : 1'b0;
  assign r_data_o[1493] = (N3)? mem[1493] : 
                          (N0)? mem[3093] : 1'b0;
  assign r_data_o[1492] = (N3)? mem[1492] : 
                          (N0)? mem[3092] : 1'b0;
  assign r_data_o[1491] = (N3)? mem[1491] : 
                          (N0)? mem[3091] : 1'b0;
  assign r_data_o[1490] = (N3)? mem[1490] : 
                          (N0)? mem[3090] : 1'b0;
  assign r_data_o[1489] = (N3)? mem[1489] : 
                          (N0)? mem[3089] : 1'b0;
  assign r_data_o[1488] = (N3)? mem[1488] : 
                          (N0)? mem[3088] : 1'b0;
  assign r_data_o[1487] = (N3)? mem[1487] : 
                          (N0)? mem[3087] : 1'b0;
  assign r_data_o[1486] = (N3)? mem[1486] : 
                          (N0)? mem[3086] : 1'b0;
  assign r_data_o[1485] = (N3)? mem[1485] : 
                          (N0)? mem[3085] : 1'b0;
  assign r_data_o[1484] = (N3)? mem[1484] : 
                          (N0)? mem[3084] : 1'b0;
  assign r_data_o[1483] = (N3)? mem[1483] : 
                          (N0)? mem[3083] : 1'b0;
  assign r_data_o[1482] = (N3)? mem[1482] : 
                          (N0)? mem[3082] : 1'b0;
  assign r_data_o[1481] = (N3)? mem[1481] : 
                          (N0)? mem[3081] : 1'b0;
  assign r_data_o[1480] = (N3)? mem[1480] : 
                          (N0)? mem[3080] : 1'b0;
  assign r_data_o[1479] = (N3)? mem[1479] : 
                          (N0)? mem[3079] : 1'b0;
  assign r_data_o[1478] = (N3)? mem[1478] : 
                          (N0)? mem[3078] : 1'b0;
  assign r_data_o[1477] = (N3)? mem[1477] : 
                          (N0)? mem[3077] : 1'b0;
  assign r_data_o[1476] = (N3)? mem[1476] : 
                          (N0)? mem[3076] : 1'b0;
  assign r_data_o[1475] = (N3)? mem[1475] : 
                          (N0)? mem[3075] : 1'b0;
  assign r_data_o[1474] = (N3)? mem[1474] : 
                          (N0)? mem[3074] : 1'b0;
  assign r_data_o[1473] = (N3)? mem[1473] : 
                          (N0)? mem[3073] : 1'b0;
  assign r_data_o[1472] = (N3)? mem[1472] : 
                          (N0)? mem[3072] : 1'b0;
  assign r_data_o[1471] = (N3)? mem[1471] : 
                          (N0)? mem[3071] : 1'b0;
  assign r_data_o[1470] = (N3)? mem[1470] : 
                          (N0)? mem[3070] : 1'b0;
  assign r_data_o[1469] = (N3)? mem[1469] : 
                          (N0)? mem[3069] : 1'b0;
  assign r_data_o[1468] = (N3)? mem[1468] : 
                          (N0)? mem[3068] : 1'b0;
  assign r_data_o[1467] = (N3)? mem[1467] : 
                          (N0)? mem[3067] : 1'b0;
  assign r_data_o[1466] = (N3)? mem[1466] : 
                          (N0)? mem[3066] : 1'b0;
  assign r_data_o[1465] = (N3)? mem[1465] : 
                          (N0)? mem[3065] : 1'b0;
  assign r_data_o[1464] = (N3)? mem[1464] : 
                          (N0)? mem[3064] : 1'b0;
  assign r_data_o[1463] = (N3)? mem[1463] : 
                          (N0)? mem[3063] : 1'b0;
  assign r_data_o[1462] = (N3)? mem[1462] : 
                          (N0)? mem[3062] : 1'b0;
  assign r_data_o[1461] = (N3)? mem[1461] : 
                          (N0)? mem[3061] : 1'b0;
  assign r_data_o[1460] = (N3)? mem[1460] : 
                          (N0)? mem[3060] : 1'b0;
  assign r_data_o[1459] = (N3)? mem[1459] : 
                          (N0)? mem[3059] : 1'b0;
  assign r_data_o[1458] = (N3)? mem[1458] : 
                          (N0)? mem[3058] : 1'b0;
  assign r_data_o[1457] = (N3)? mem[1457] : 
                          (N0)? mem[3057] : 1'b0;
  assign r_data_o[1456] = (N3)? mem[1456] : 
                          (N0)? mem[3056] : 1'b0;
  assign r_data_o[1455] = (N3)? mem[1455] : 
                          (N0)? mem[3055] : 1'b0;
  assign r_data_o[1454] = (N3)? mem[1454] : 
                          (N0)? mem[3054] : 1'b0;
  assign r_data_o[1453] = (N3)? mem[1453] : 
                          (N0)? mem[3053] : 1'b0;
  assign r_data_o[1452] = (N3)? mem[1452] : 
                          (N0)? mem[3052] : 1'b0;
  assign r_data_o[1451] = (N3)? mem[1451] : 
                          (N0)? mem[3051] : 1'b0;
  assign r_data_o[1450] = (N3)? mem[1450] : 
                          (N0)? mem[3050] : 1'b0;
  assign r_data_o[1449] = (N3)? mem[1449] : 
                          (N0)? mem[3049] : 1'b0;
  assign r_data_o[1448] = (N3)? mem[1448] : 
                          (N0)? mem[3048] : 1'b0;
  assign r_data_o[1447] = (N3)? mem[1447] : 
                          (N0)? mem[3047] : 1'b0;
  assign r_data_o[1446] = (N3)? mem[1446] : 
                          (N0)? mem[3046] : 1'b0;
  assign r_data_o[1445] = (N3)? mem[1445] : 
                          (N0)? mem[3045] : 1'b0;
  assign r_data_o[1444] = (N3)? mem[1444] : 
                          (N0)? mem[3044] : 1'b0;
  assign r_data_o[1443] = (N3)? mem[1443] : 
                          (N0)? mem[3043] : 1'b0;
  assign r_data_o[1442] = (N3)? mem[1442] : 
                          (N0)? mem[3042] : 1'b0;
  assign r_data_o[1441] = (N3)? mem[1441] : 
                          (N0)? mem[3041] : 1'b0;
  assign r_data_o[1440] = (N3)? mem[1440] : 
                          (N0)? mem[3040] : 1'b0;
  assign r_data_o[1439] = (N3)? mem[1439] : 
                          (N0)? mem[3039] : 1'b0;
  assign r_data_o[1438] = (N3)? mem[1438] : 
                          (N0)? mem[3038] : 1'b0;
  assign r_data_o[1437] = (N3)? mem[1437] : 
                          (N0)? mem[3037] : 1'b0;
  assign r_data_o[1436] = (N3)? mem[1436] : 
                          (N0)? mem[3036] : 1'b0;
  assign r_data_o[1435] = (N3)? mem[1435] : 
                          (N0)? mem[3035] : 1'b0;
  assign r_data_o[1434] = (N3)? mem[1434] : 
                          (N0)? mem[3034] : 1'b0;
  assign r_data_o[1433] = (N3)? mem[1433] : 
                          (N0)? mem[3033] : 1'b0;
  assign r_data_o[1432] = (N3)? mem[1432] : 
                          (N0)? mem[3032] : 1'b0;
  assign r_data_o[1431] = (N3)? mem[1431] : 
                          (N0)? mem[3031] : 1'b0;
  assign r_data_o[1430] = (N3)? mem[1430] : 
                          (N0)? mem[3030] : 1'b0;
  assign r_data_o[1429] = (N3)? mem[1429] : 
                          (N0)? mem[3029] : 1'b0;
  assign r_data_o[1428] = (N3)? mem[1428] : 
                          (N0)? mem[3028] : 1'b0;
  assign r_data_o[1427] = (N3)? mem[1427] : 
                          (N0)? mem[3027] : 1'b0;
  assign r_data_o[1426] = (N3)? mem[1426] : 
                          (N0)? mem[3026] : 1'b0;
  assign r_data_o[1425] = (N3)? mem[1425] : 
                          (N0)? mem[3025] : 1'b0;
  assign r_data_o[1424] = (N3)? mem[1424] : 
                          (N0)? mem[3024] : 1'b0;
  assign r_data_o[1423] = (N3)? mem[1423] : 
                          (N0)? mem[3023] : 1'b0;
  assign r_data_o[1422] = (N3)? mem[1422] : 
                          (N0)? mem[3022] : 1'b0;
  assign r_data_o[1421] = (N3)? mem[1421] : 
                          (N0)? mem[3021] : 1'b0;
  assign r_data_o[1420] = (N3)? mem[1420] : 
                          (N0)? mem[3020] : 1'b0;
  assign r_data_o[1419] = (N3)? mem[1419] : 
                          (N0)? mem[3019] : 1'b0;
  assign r_data_o[1418] = (N3)? mem[1418] : 
                          (N0)? mem[3018] : 1'b0;
  assign r_data_o[1417] = (N3)? mem[1417] : 
                          (N0)? mem[3017] : 1'b0;
  assign r_data_o[1416] = (N3)? mem[1416] : 
                          (N0)? mem[3016] : 1'b0;
  assign r_data_o[1415] = (N3)? mem[1415] : 
                          (N0)? mem[3015] : 1'b0;
  assign r_data_o[1414] = (N3)? mem[1414] : 
                          (N0)? mem[3014] : 1'b0;
  assign r_data_o[1413] = (N3)? mem[1413] : 
                          (N0)? mem[3013] : 1'b0;
  assign r_data_o[1412] = (N3)? mem[1412] : 
                          (N0)? mem[3012] : 1'b0;
  assign r_data_o[1411] = (N3)? mem[1411] : 
                          (N0)? mem[3011] : 1'b0;
  assign r_data_o[1410] = (N3)? mem[1410] : 
                          (N0)? mem[3010] : 1'b0;
  assign r_data_o[1409] = (N3)? mem[1409] : 
                          (N0)? mem[3009] : 1'b0;
  assign r_data_o[1408] = (N3)? mem[1408] : 
                          (N0)? mem[3008] : 1'b0;
  assign r_data_o[1407] = (N3)? mem[1407] : 
                          (N0)? mem[3007] : 1'b0;
  assign r_data_o[1406] = (N3)? mem[1406] : 
                          (N0)? mem[3006] : 1'b0;
  assign r_data_o[1405] = (N3)? mem[1405] : 
                          (N0)? mem[3005] : 1'b0;
  assign r_data_o[1404] = (N3)? mem[1404] : 
                          (N0)? mem[3004] : 1'b0;
  assign r_data_o[1403] = (N3)? mem[1403] : 
                          (N0)? mem[3003] : 1'b0;
  assign r_data_o[1402] = (N3)? mem[1402] : 
                          (N0)? mem[3002] : 1'b0;
  assign r_data_o[1401] = (N3)? mem[1401] : 
                          (N0)? mem[3001] : 1'b0;
  assign r_data_o[1400] = (N3)? mem[1400] : 
                          (N0)? mem[3000] : 1'b0;
  assign r_data_o[1399] = (N3)? mem[1399] : 
                          (N0)? mem[2999] : 1'b0;
  assign r_data_o[1398] = (N3)? mem[1398] : 
                          (N0)? mem[2998] : 1'b0;
  assign r_data_o[1397] = (N3)? mem[1397] : 
                          (N0)? mem[2997] : 1'b0;
  assign r_data_o[1396] = (N3)? mem[1396] : 
                          (N0)? mem[2996] : 1'b0;
  assign r_data_o[1395] = (N3)? mem[1395] : 
                          (N0)? mem[2995] : 1'b0;
  assign r_data_o[1394] = (N3)? mem[1394] : 
                          (N0)? mem[2994] : 1'b0;
  assign r_data_o[1393] = (N3)? mem[1393] : 
                          (N0)? mem[2993] : 1'b0;
  assign r_data_o[1392] = (N3)? mem[1392] : 
                          (N0)? mem[2992] : 1'b0;
  assign r_data_o[1391] = (N3)? mem[1391] : 
                          (N0)? mem[2991] : 1'b0;
  assign r_data_o[1390] = (N3)? mem[1390] : 
                          (N0)? mem[2990] : 1'b0;
  assign r_data_o[1389] = (N3)? mem[1389] : 
                          (N0)? mem[2989] : 1'b0;
  assign r_data_o[1388] = (N3)? mem[1388] : 
                          (N0)? mem[2988] : 1'b0;
  assign r_data_o[1387] = (N3)? mem[1387] : 
                          (N0)? mem[2987] : 1'b0;
  assign r_data_o[1386] = (N3)? mem[1386] : 
                          (N0)? mem[2986] : 1'b0;
  assign r_data_o[1385] = (N3)? mem[1385] : 
                          (N0)? mem[2985] : 1'b0;
  assign r_data_o[1384] = (N3)? mem[1384] : 
                          (N0)? mem[2984] : 1'b0;
  assign r_data_o[1383] = (N3)? mem[1383] : 
                          (N0)? mem[2983] : 1'b0;
  assign r_data_o[1382] = (N3)? mem[1382] : 
                          (N0)? mem[2982] : 1'b0;
  assign r_data_o[1381] = (N3)? mem[1381] : 
                          (N0)? mem[2981] : 1'b0;
  assign r_data_o[1380] = (N3)? mem[1380] : 
                          (N0)? mem[2980] : 1'b0;
  assign r_data_o[1379] = (N3)? mem[1379] : 
                          (N0)? mem[2979] : 1'b0;
  assign r_data_o[1378] = (N3)? mem[1378] : 
                          (N0)? mem[2978] : 1'b0;
  assign r_data_o[1377] = (N3)? mem[1377] : 
                          (N0)? mem[2977] : 1'b0;
  assign r_data_o[1376] = (N3)? mem[1376] : 
                          (N0)? mem[2976] : 1'b0;
  assign r_data_o[1375] = (N3)? mem[1375] : 
                          (N0)? mem[2975] : 1'b0;
  assign r_data_o[1374] = (N3)? mem[1374] : 
                          (N0)? mem[2974] : 1'b0;
  assign r_data_o[1373] = (N3)? mem[1373] : 
                          (N0)? mem[2973] : 1'b0;
  assign r_data_o[1372] = (N3)? mem[1372] : 
                          (N0)? mem[2972] : 1'b0;
  assign r_data_o[1371] = (N3)? mem[1371] : 
                          (N0)? mem[2971] : 1'b0;
  assign r_data_o[1370] = (N3)? mem[1370] : 
                          (N0)? mem[2970] : 1'b0;
  assign r_data_o[1369] = (N3)? mem[1369] : 
                          (N0)? mem[2969] : 1'b0;
  assign r_data_o[1368] = (N3)? mem[1368] : 
                          (N0)? mem[2968] : 1'b0;
  assign r_data_o[1367] = (N3)? mem[1367] : 
                          (N0)? mem[2967] : 1'b0;
  assign r_data_o[1366] = (N3)? mem[1366] : 
                          (N0)? mem[2966] : 1'b0;
  assign r_data_o[1365] = (N3)? mem[1365] : 
                          (N0)? mem[2965] : 1'b0;
  assign r_data_o[1364] = (N3)? mem[1364] : 
                          (N0)? mem[2964] : 1'b0;
  assign r_data_o[1363] = (N3)? mem[1363] : 
                          (N0)? mem[2963] : 1'b0;
  assign r_data_o[1362] = (N3)? mem[1362] : 
                          (N0)? mem[2962] : 1'b0;
  assign r_data_o[1361] = (N3)? mem[1361] : 
                          (N0)? mem[2961] : 1'b0;
  assign r_data_o[1360] = (N3)? mem[1360] : 
                          (N0)? mem[2960] : 1'b0;
  assign r_data_o[1359] = (N3)? mem[1359] : 
                          (N0)? mem[2959] : 1'b0;
  assign r_data_o[1358] = (N3)? mem[1358] : 
                          (N0)? mem[2958] : 1'b0;
  assign r_data_o[1357] = (N3)? mem[1357] : 
                          (N0)? mem[2957] : 1'b0;
  assign r_data_o[1356] = (N3)? mem[1356] : 
                          (N0)? mem[2956] : 1'b0;
  assign r_data_o[1355] = (N3)? mem[1355] : 
                          (N0)? mem[2955] : 1'b0;
  assign r_data_o[1354] = (N3)? mem[1354] : 
                          (N0)? mem[2954] : 1'b0;
  assign r_data_o[1353] = (N3)? mem[1353] : 
                          (N0)? mem[2953] : 1'b0;
  assign r_data_o[1352] = (N3)? mem[1352] : 
                          (N0)? mem[2952] : 1'b0;
  assign r_data_o[1351] = (N3)? mem[1351] : 
                          (N0)? mem[2951] : 1'b0;
  assign r_data_o[1350] = (N3)? mem[1350] : 
                          (N0)? mem[2950] : 1'b0;
  assign r_data_o[1349] = (N3)? mem[1349] : 
                          (N0)? mem[2949] : 1'b0;
  assign r_data_o[1348] = (N3)? mem[1348] : 
                          (N0)? mem[2948] : 1'b0;
  assign r_data_o[1347] = (N3)? mem[1347] : 
                          (N0)? mem[2947] : 1'b0;
  assign r_data_o[1346] = (N3)? mem[1346] : 
                          (N0)? mem[2946] : 1'b0;
  assign r_data_o[1345] = (N3)? mem[1345] : 
                          (N0)? mem[2945] : 1'b0;
  assign r_data_o[1344] = (N3)? mem[1344] : 
                          (N0)? mem[2944] : 1'b0;
  assign r_data_o[1343] = (N3)? mem[1343] : 
                          (N0)? mem[2943] : 1'b0;
  assign r_data_o[1342] = (N3)? mem[1342] : 
                          (N0)? mem[2942] : 1'b0;
  assign r_data_o[1341] = (N3)? mem[1341] : 
                          (N0)? mem[2941] : 1'b0;
  assign r_data_o[1340] = (N3)? mem[1340] : 
                          (N0)? mem[2940] : 1'b0;
  assign r_data_o[1339] = (N3)? mem[1339] : 
                          (N0)? mem[2939] : 1'b0;
  assign r_data_o[1338] = (N3)? mem[1338] : 
                          (N0)? mem[2938] : 1'b0;
  assign r_data_o[1337] = (N3)? mem[1337] : 
                          (N0)? mem[2937] : 1'b0;
  assign r_data_o[1336] = (N3)? mem[1336] : 
                          (N0)? mem[2936] : 1'b0;
  assign r_data_o[1335] = (N3)? mem[1335] : 
                          (N0)? mem[2935] : 1'b0;
  assign r_data_o[1334] = (N3)? mem[1334] : 
                          (N0)? mem[2934] : 1'b0;
  assign r_data_o[1333] = (N3)? mem[1333] : 
                          (N0)? mem[2933] : 1'b0;
  assign r_data_o[1332] = (N3)? mem[1332] : 
                          (N0)? mem[2932] : 1'b0;
  assign r_data_o[1331] = (N3)? mem[1331] : 
                          (N0)? mem[2931] : 1'b0;
  assign r_data_o[1330] = (N3)? mem[1330] : 
                          (N0)? mem[2930] : 1'b0;
  assign r_data_o[1329] = (N3)? mem[1329] : 
                          (N0)? mem[2929] : 1'b0;
  assign r_data_o[1328] = (N3)? mem[1328] : 
                          (N0)? mem[2928] : 1'b0;
  assign r_data_o[1327] = (N3)? mem[1327] : 
                          (N0)? mem[2927] : 1'b0;
  assign r_data_o[1326] = (N3)? mem[1326] : 
                          (N0)? mem[2926] : 1'b0;
  assign r_data_o[1325] = (N3)? mem[1325] : 
                          (N0)? mem[2925] : 1'b0;
  assign r_data_o[1324] = (N3)? mem[1324] : 
                          (N0)? mem[2924] : 1'b0;
  assign r_data_o[1323] = (N3)? mem[1323] : 
                          (N0)? mem[2923] : 1'b0;
  assign r_data_o[1322] = (N3)? mem[1322] : 
                          (N0)? mem[2922] : 1'b0;
  assign r_data_o[1321] = (N3)? mem[1321] : 
                          (N0)? mem[2921] : 1'b0;
  assign r_data_o[1320] = (N3)? mem[1320] : 
                          (N0)? mem[2920] : 1'b0;
  assign r_data_o[1319] = (N3)? mem[1319] : 
                          (N0)? mem[2919] : 1'b0;
  assign r_data_o[1318] = (N3)? mem[1318] : 
                          (N0)? mem[2918] : 1'b0;
  assign r_data_o[1317] = (N3)? mem[1317] : 
                          (N0)? mem[2917] : 1'b0;
  assign r_data_o[1316] = (N3)? mem[1316] : 
                          (N0)? mem[2916] : 1'b0;
  assign r_data_o[1315] = (N3)? mem[1315] : 
                          (N0)? mem[2915] : 1'b0;
  assign r_data_o[1314] = (N3)? mem[1314] : 
                          (N0)? mem[2914] : 1'b0;
  assign r_data_o[1313] = (N3)? mem[1313] : 
                          (N0)? mem[2913] : 1'b0;
  assign r_data_o[1312] = (N3)? mem[1312] : 
                          (N0)? mem[2912] : 1'b0;
  assign r_data_o[1311] = (N3)? mem[1311] : 
                          (N0)? mem[2911] : 1'b0;
  assign r_data_o[1310] = (N3)? mem[1310] : 
                          (N0)? mem[2910] : 1'b0;
  assign r_data_o[1309] = (N3)? mem[1309] : 
                          (N0)? mem[2909] : 1'b0;
  assign r_data_o[1308] = (N3)? mem[1308] : 
                          (N0)? mem[2908] : 1'b0;
  assign r_data_o[1307] = (N3)? mem[1307] : 
                          (N0)? mem[2907] : 1'b0;
  assign r_data_o[1306] = (N3)? mem[1306] : 
                          (N0)? mem[2906] : 1'b0;
  assign r_data_o[1305] = (N3)? mem[1305] : 
                          (N0)? mem[2905] : 1'b0;
  assign r_data_o[1304] = (N3)? mem[1304] : 
                          (N0)? mem[2904] : 1'b0;
  assign r_data_o[1303] = (N3)? mem[1303] : 
                          (N0)? mem[2903] : 1'b0;
  assign r_data_o[1302] = (N3)? mem[1302] : 
                          (N0)? mem[2902] : 1'b0;
  assign r_data_o[1301] = (N3)? mem[1301] : 
                          (N0)? mem[2901] : 1'b0;
  assign r_data_o[1300] = (N3)? mem[1300] : 
                          (N0)? mem[2900] : 1'b0;
  assign r_data_o[1299] = (N3)? mem[1299] : 
                          (N0)? mem[2899] : 1'b0;
  assign r_data_o[1298] = (N3)? mem[1298] : 
                          (N0)? mem[2898] : 1'b0;
  assign r_data_o[1297] = (N3)? mem[1297] : 
                          (N0)? mem[2897] : 1'b0;
  assign r_data_o[1296] = (N3)? mem[1296] : 
                          (N0)? mem[2896] : 1'b0;
  assign r_data_o[1295] = (N3)? mem[1295] : 
                          (N0)? mem[2895] : 1'b0;
  assign r_data_o[1294] = (N3)? mem[1294] : 
                          (N0)? mem[2894] : 1'b0;
  assign r_data_o[1293] = (N3)? mem[1293] : 
                          (N0)? mem[2893] : 1'b0;
  assign r_data_o[1292] = (N3)? mem[1292] : 
                          (N0)? mem[2892] : 1'b0;
  assign r_data_o[1291] = (N3)? mem[1291] : 
                          (N0)? mem[2891] : 1'b0;
  assign r_data_o[1290] = (N3)? mem[1290] : 
                          (N0)? mem[2890] : 1'b0;
  assign r_data_o[1289] = (N3)? mem[1289] : 
                          (N0)? mem[2889] : 1'b0;
  assign r_data_o[1288] = (N3)? mem[1288] : 
                          (N0)? mem[2888] : 1'b0;
  assign r_data_o[1287] = (N3)? mem[1287] : 
                          (N0)? mem[2887] : 1'b0;
  assign r_data_o[1286] = (N3)? mem[1286] : 
                          (N0)? mem[2886] : 1'b0;
  assign r_data_o[1285] = (N3)? mem[1285] : 
                          (N0)? mem[2885] : 1'b0;
  assign r_data_o[1284] = (N3)? mem[1284] : 
                          (N0)? mem[2884] : 1'b0;
  assign r_data_o[1283] = (N3)? mem[1283] : 
                          (N0)? mem[2883] : 1'b0;
  assign r_data_o[1282] = (N3)? mem[1282] : 
                          (N0)? mem[2882] : 1'b0;
  assign r_data_o[1281] = (N3)? mem[1281] : 
                          (N0)? mem[2881] : 1'b0;
  assign r_data_o[1280] = (N3)? mem[1280] : 
                          (N0)? mem[2880] : 1'b0;
  assign r_data_o[1279] = (N3)? mem[1279] : 
                          (N0)? mem[2879] : 1'b0;
  assign r_data_o[1278] = (N3)? mem[1278] : 
                          (N0)? mem[2878] : 1'b0;
  assign r_data_o[1277] = (N3)? mem[1277] : 
                          (N0)? mem[2877] : 1'b0;
  assign r_data_o[1276] = (N3)? mem[1276] : 
                          (N0)? mem[2876] : 1'b0;
  assign r_data_o[1275] = (N3)? mem[1275] : 
                          (N0)? mem[2875] : 1'b0;
  assign r_data_o[1274] = (N3)? mem[1274] : 
                          (N0)? mem[2874] : 1'b0;
  assign r_data_o[1273] = (N3)? mem[1273] : 
                          (N0)? mem[2873] : 1'b0;
  assign r_data_o[1272] = (N3)? mem[1272] : 
                          (N0)? mem[2872] : 1'b0;
  assign r_data_o[1271] = (N3)? mem[1271] : 
                          (N0)? mem[2871] : 1'b0;
  assign r_data_o[1270] = (N3)? mem[1270] : 
                          (N0)? mem[2870] : 1'b0;
  assign r_data_o[1269] = (N3)? mem[1269] : 
                          (N0)? mem[2869] : 1'b0;
  assign r_data_o[1268] = (N3)? mem[1268] : 
                          (N0)? mem[2868] : 1'b0;
  assign r_data_o[1267] = (N3)? mem[1267] : 
                          (N0)? mem[2867] : 1'b0;
  assign r_data_o[1266] = (N3)? mem[1266] : 
                          (N0)? mem[2866] : 1'b0;
  assign r_data_o[1265] = (N3)? mem[1265] : 
                          (N0)? mem[2865] : 1'b0;
  assign r_data_o[1264] = (N3)? mem[1264] : 
                          (N0)? mem[2864] : 1'b0;
  assign r_data_o[1263] = (N3)? mem[1263] : 
                          (N0)? mem[2863] : 1'b0;
  assign r_data_o[1262] = (N3)? mem[1262] : 
                          (N0)? mem[2862] : 1'b0;
  assign r_data_o[1261] = (N3)? mem[1261] : 
                          (N0)? mem[2861] : 1'b0;
  assign r_data_o[1260] = (N3)? mem[1260] : 
                          (N0)? mem[2860] : 1'b0;
  assign r_data_o[1259] = (N3)? mem[1259] : 
                          (N0)? mem[2859] : 1'b0;
  assign r_data_o[1258] = (N3)? mem[1258] : 
                          (N0)? mem[2858] : 1'b0;
  assign r_data_o[1257] = (N3)? mem[1257] : 
                          (N0)? mem[2857] : 1'b0;
  assign r_data_o[1256] = (N3)? mem[1256] : 
                          (N0)? mem[2856] : 1'b0;
  assign r_data_o[1255] = (N3)? mem[1255] : 
                          (N0)? mem[2855] : 1'b0;
  assign r_data_o[1254] = (N3)? mem[1254] : 
                          (N0)? mem[2854] : 1'b0;
  assign r_data_o[1253] = (N3)? mem[1253] : 
                          (N0)? mem[2853] : 1'b0;
  assign r_data_o[1252] = (N3)? mem[1252] : 
                          (N0)? mem[2852] : 1'b0;
  assign r_data_o[1251] = (N3)? mem[1251] : 
                          (N0)? mem[2851] : 1'b0;
  assign r_data_o[1250] = (N3)? mem[1250] : 
                          (N0)? mem[2850] : 1'b0;
  assign r_data_o[1249] = (N3)? mem[1249] : 
                          (N0)? mem[2849] : 1'b0;
  assign r_data_o[1248] = (N3)? mem[1248] : 
                          (N0)? mem[2848] : 1'b0;
  assign r_data_o[1247] = (N3)? mem[1247] : 
                          (N0)? mem[2847] : 1'b0;
  assign r_data_o[1246] = (N3)? mem[1246] : 
                          (N0)? mem[2846] : 1'b0;
  assign r_data_o[1245] = (N3)? mem[1245] : 
                          (N0)? mem[2845] : 1'b0;
  assign r_data_o[1244] = (N3)? mem[1244] : 
                          (N0)? mem[2844] : 1'b0;
  assign r_data_o[1243] = (N3)? mem[1243] : 
                          (N0)? mem[2843] : 1'b0;
  assign r_data_o[1242] = (N3)? mem[1242] : 
                          (N0)? mem[2842] : 1'b0;
  assign r_data_o[1241] = (N3)? mem[1241] : 
                          (N0)? mem[2841] : 1'b0;
  assign r_data_o[1240] = (N3)? mem[1240] : 
                          (N0)? mem[2840] : 1'b0;
  assign r_data_o[1239] = (N3)? mem[1239] : 
                          (N0)? mem[2839] : 1'b0;
  assign r_data_o[1238] = (N3)? mem[1238] : 
                          (N0)? mem[2838] : 1'b0;
  assign r_data_o[1237] = (N3)? mem[1237] : 
                          (N0)? mem[2837] : 1'b0;
  assign r_data_o[1236] = (N3)? mem[1236] : 
                          (N0)? mem[2836] : 1'b0;
  assign r_data_o[1235] = (N3)? mem[1235] : 
                          (N0)? mem[2835] : 1'b0;
  assign r_data_o[1234] = (N3)? mem[1234] : 
                          (N0)? mem[2834] : 1'b0;
  assign r_data_o[1233] = (N3)? mem[1233] : 
                          (N0)? mem[2833] : 1'b0;
  assign r_data_o[1232] = (N3)? mem[1232] : 
                          (N0)? mem[2832] : 1'b0;
  assign r_data_o[1231] = (N3)? mem[1231] : 
                          (N0)? mem[2831] : 1'b0;
  assign r_data_o[1230] = (N3)? mem[1230] : 
                          (N0)? mem[2830] : 1'b0;
  assign r_data_o[1229] = (N3)? mem[1229] : 
                          (N0)? mem[2829] : 1'b0;
  assign r_data_o[1228] = (N3)? mem[1228] : 
                          (N0)? mem[2828] : 1'b0;
  assign r_data_o[1227] = (N3)? mem[1227] : 
                          (N0)? mem[2827] : 1'b0;
  assign r_data_o[1226] = (N3)? mem[1226] : 
                          (N0)? mem[2826] : 1'b0;
  assign r_data_o[1225] = (N3)? mem[1225] : 
                          (N0)? mem[2825] : 1'b0;
  assign r_data_o[1224] = (N3)? mem[1224] : 
                          (N0)? mem[2824] : 1'b0;
  assign r_data_o[1223] = (N3)? mem[1223] : 
                          (N0)? mem[2823] : 1'b0;
  assign r_data_o[1222] = (N3)? mem[1222] : 
                          (N0)? mem[2822] : 1'b0;
  assign r_data_o[1221] = (N3)? mem[1221] : 
                          (N0)? mem[2821] : 1'b0;
  assign r_data_o[1220] = (N3)? mem[1220] : 
                          (N0)? mem[2820] : 1'b0;
  assign r_data_o[1219] = (N3)? mem[1219] : 
                          (N0)? mem[2819] : 1'b0;
  assign r_data_o[1218] = (N3)? mem[1218] : 
                          (N0)? mem[2818] : 1'b0;
  assign r_data_o[1217] = (N3)? mem[1217] : 
                          (N0)? mem[2817] : 1'b0;
  assign r_data_o[1216] = (N3)? mem[1216] : 
                          (N0)? mem[2816] : 1'b0;
  assign r_data_o[1215] = (N3)? mem[1215] : 
                          (N0)? mem[2815] : 1'b0;
  assign r_data_o[1214] = (N3)? mem[1214] : 
                          (N0)? mem[2814] : 1'b0;
  assign r_data_o[1213] = (N3)? mem[1213] : 
                          (N0)? mem[2813] : 1'b0;
  assign r_data_o[1212] = (N3)? mem[1212] : 
                          (N0)? mem[2812] : 1'b0;
  assign r_data_o[1211] = (N3)? mem[1211] : 
                          (N0)? mem[2811] : 1'b0;
  assign r_data_o[1210] = (N3)? mem[1210] : 
                          (N0)? mem[2810] : 1'b0;
  assign r_data_o[1209] = (N3)? mem[1209] : 
                          (N0)? mem[2809] : 1'b0;
  assign r_data_o[1208] = (N3)? mem[1208] : 
                          (N0)? mem[2808] : 1'b0;
  assign r_data_o[1207] = (N3)? mem[1207] : 
                          (N0)? mem[2807] : 1'b0;
  assign r_data_o[1206] = (N3)? mem[1206] : 
                          (N0)? mem[2806] : 1'b0;
  assign r_data_o[1205] = (N3)? mem[1205] : 
                          (N0)? mem[2805] : 1'b0;
  assign r_data_o[1204] = (N3)? mem[1204] : 
                          (N0)? mem[2804] : 1'b0;
  assign r_data_o[1203] = (N3)? mem[1203] : 
                          (N0)? mem[2803] : 1'b0;
  assign r_data_o[1202] = (N3)? mem[1202] : 
                          (N0)? mem[2802] : 1'b0;
  assign r_data_o[1201] = (N3)? mem[1201] : 
                          (N0)? mem[2801] : 1'b0;
  assign r_data_o[1200] = (N3)? mem[1200] : 
                          (N0)? mem[2800] : 1'b0;
  assign r_data_o[1199] = (N3)? mem[1199] : 
                          (N0)? mem[2799] : 1'b0;
  assign r_data_o[1198] = (N3)? mem[1198] : 
                          (N0)? mem[2798] : 1'b0;
  assign r_data_o[1197] = (N3)? mem[1197] : 
                          (N0)? mem[2797] : 1'b0;
  assign r_data_o[1196] = (N3)? mem[1196] : 
                          (N0)? mem[2796] : 1'b0;
  assign r_data_o[1195] = (N3)? mem[1195] : 
                          (N0)? mem[2795] : 1'b0;
  assign r_data_o[1194] = (N3)? mem[1194] : 
                          (N0)? mem[2794] : 1'b0;
  assign r_data_o[1193] = (N3)? mem[1193] : 
                          (N0)? mem[2793] : 1'b0;
  assign r_data_o[1192] = (N3)? mem[1192] : 
                          (N0)? mem[2792] : 1'b0;
  assign r_data_o[1191] = (N3)? mem[1191] : 
                          (N0)? mem[2791] : 1'b0;
  assign r_data_o[1190] = (N3)? mem[1190] : 
                          (N0)? mem[2790] : 1'b0;
  assign r_data_o[1189] = (N3)? mem[1189] : 
                          (N0)? mem[2789] : 1'b0;
  assign r_data_o[1188] = (N3)? mem[1188] : 
                          (N0)? mem[2788] : 1'b0;
  assign r_data_o[1187] = (N3)? mem[1187] : 
                          (N0)? mem[2787] : 1'b0;
  assign r_data_o[1186] = (N3)? mem[1186] : 
                          (N0)? mem[2786] : 1'b0;
  assign r_data_o[1185] = (N3)? mem[1185] : 
                          (N0)? mem[2785] : 1'b0;
  assign r_data_o[1184] = (N3)? mem[1184] : 
                          (N0)? mem[2784] : 1'b0;
  assign r_data_o[1183] = (N3)? mem[1183] : 
                          (N0)? mem[2783] : 1'b0;
  assign r_data_o[1182] = (N3)? mem[1182] : 
                          (N0)? mem[2782] : 1'b0;
  assign r_data_o[1181] = (N3)? mem[1181] : 
                          (N0)? mem[2781] : 1'b0;
  assign r_data_o[1180] = (N3)? mem[1180] : 
                          (N0)? mem[2780] : 1'b0;
  assign r_data_o[1179] = (N3)? mem[1179] : 
                          (N0)? mem[2779] : 1'b0;
  assign r_data_o[1178] = (N3)? mem[1178] : 
                          (N0)? mem[2778] : 1'b0;
  assign r_data_o[1177] = (N3)? mem[1177] : 
                          (N0)? mem[2777] : 1'b0;
  assign r_data_o[1176] = (N3)? mem[1176] : 
                          (N0)? mem[2776] : 1'b0;
  assign r_data_o[1175] = (N3)? mem[1175] : 
                          (N0)? mem[2775] : 1'b0;
  assign r_data_o[1174] = (N3)? mem[1174] : 
                          (N0)? mem[2774] : 1'b0;
  assign r_data_o[1173] = (N3)? mem[1173] : 
                          (N0)? mem[2773] : 1'b0;
  assign r_data_o[1172] = (N3)? mem[1172] : 
                          (N0)? mem[2772] : 1'b0;
  assign r_data_o[1171] = (N3)? mem[1171] : 
                          (N0)? mem[2771] : 1'b0;
  assign r_data_o[1170] = (N3)? mem[1170] : 
                          (N0)? mem[2770] : 1'b0;
  assign r_data_o[1169] = (N3)? mem[1169] : 
                          (N0)? mem[2769] : 1'b0;
  assign r_data_o[1168] = (N3)? mem[1168] : 
                          (N0)? mem[2768] : 1'b0;
  assign r_data_o[1167] = (N3)? mem[1167] : 
                          (N0)? mem[2767] : 1'b0;
  assign r_data_o[1166] = (N3)? mem[1166] : 
                          (N0)? mem[2766] : 1'b0;
  assign r_data_o[1165] = (N3)? mem[1165] : 
                          (N0)? mem[2765] : 1'b0;
  assign r_data_o[1164] = (N3)? mem[1164] : 
                          (N0)? mem[2764] : 1'b0;
  assign r_data_o[1163] = (N3)? mem[1163] : 
                          (N0)? mem[2763] : 1'b0;
  assign r_data_o[1162] = (N3)? mem[1162] : 
                          (N0)? mem[2762] : 1'b0;
  assign r_data_o[1161] = (N3)? mem[1161] : 
                          (N0)? mem[2761] : 1'b0;
  assign r_data_o[1160] = (N3)? mem[1160] : 
                          (N0)? mem[2760] : 1'b0;
  assign r_data_o[1159] = (N3)? mem[1159] : 
                          (N0)? mem[2759] : 1'b0;
  assign r_data_o[1158] = (N3)? mem[1158] : 
                          (N0)? mem[2758] : 1'b0;
  assign r_data_o[1157] = (N3)? mem[1157] : 
                          (N0)? mem[2757] : 1'b0;
  assign r_data_o[1156] = (N3)? mem[1156] : 
                          (N0)? mem[2756] : 1'b0;
  assign r_data_o[1155] = (N3)? mem[1155] : 
                          (N0)? mem[2755] : 1'b0;
  assign r_data_o[1154] = (N3)? mem[1154] : 
                          (N0)? mem[2754] : 1'b0;
  assign r_data_o[1153] = (N3)? mem[1153] : 
                          (N0)? mem[2753] : 1'b0;
  assign r_data_o[1152] = (N3)? mem[1152] : 
                          (N0)? mem[2752] : 1'b0;
  assign r_data_o[1151] = (N3)? mem[1151] : 
                          (N0)? mem[2751] : 1'b0;
  assign r_data_o[1150] = (N3)? mem[1150] : 
                          (N0)? mem[2750] : 1'b0;
  assign r_data_o[1149] = (N3)? mem[1149] : 
                          (N0)? mem[2749] : 1'b0;
  assign r_data_o[1148] = (N3)? mem[1148] : 
                          (N0)? mem[2748] : 1'b0;
  assign r_data_o[1147] = (N3)? mem[1147] : 
                          (N0)? mem[2747] : 1'b0;
  assign r_data_o[1146] = (N3)? mem[1146] : 
                          (N0)? mem[2746] : 1'b0;
  assign r_data_o[1145] = (N3)? mem[1145] : 
                          (N0)? mem[2745] : 1'b0;
  assign r_data_o[1144] = (N3)? mem[1144] : 
                          (N0)? mem[2744] : 1'b0;
  assign r_data_o[1143] = (N3)? mem[1143] : 
                          (N0)? mem[2743] : 1'b0;
  assign r_data_o[1142] = (N3)? mem[1142] : 
                          (N0)? mem[2742] : 1'b0;
  assign r_data_o[1141] = (N3)? mem[1141] : 
                          (N0)? mem[2741] : 1'b0;
  assign r_data_o[1140] = (N3)? mem[1140] : 
                          (N0)? mem[2740] : 1'b0;
  assign r_data_o[1139] = (N3)? mem[1139] : 
                          (N0)? mem[2739] : 1'b0;
  assign r_data_o[1138] = (N3)? mem[1138] : 
                          (N0)? mem[2738] : 1'b0;
  assign r_data_o[1137] = (N3)? mem[1137] : 
                          (N0)? mem[2737] : 1'b0;
  assign r_data_o[1136] = (N3)? mem[1136] : 
                          (N0)? mem[2736] : 1'b0;
  assign r_data_o[1135] = (N3)? mem[1135] : 
                          (N0)? mem[2735] : 1'b0;
  assign r_data_o[1134] = (N3)? mem[1134] : 
                          (N0)? mem[2734] : 1'b0;
  assign r_data_o[1133] = (N3)? mem[1133] : 
                          (N0)? mem[2733] : 1'b0;
  assign r_data_o[1132] = (N3)? mem[1132] : 
                          (N0)? mem[2732] : 1'b0;
  assign r_data_o[1131] = (N3)? mem[1131] : 
                          (N0)? mem[2731] : 1'b0;
  assign r_data_o[1130] = (N3)? mem[1130] : 
                          (N0)? mem[2730] : 1'b0;
  assign r_data_o[1129] = (N3)? mem[1129] : 
                          (N0)? mem[2729] : 1'b0;
  assign r_data_o[1128] = (N3)? mem[1128] : 
                          (N0)? mem[2728] : 1'b0;
  assign r_data_o[1127] = (N3)? mem[1127] : 
                          (N0)? mem[2727] : 1'b0;
  assign r_data_o[1126] = (N3)? mem[1126] : 
                          (N0)? mem[2726] : 1'b0;
  assign r_data_o[1125] = (N3)? mem[1125] : 
                          (N0)? mem[2725] : 1'b0;
  assign r_data_o[1124] = (N3)? mem[1124] : 
                          (N0)? mem[2724] : 1'b0;
  assign r_data_o[1123] = (N3)? mem[1123] : 
                          (N0)? mem[2723] : 1'b0;
  assign r_data_o[1122] = (N3)? mem[1122] : 
                          (N0)? mem[2722] : 1'b0;
  assign r_data_o[1121] = (N3)? mem[1121] : 
                          (N0)? mem[2721] : 1'b0;
  assign r_data_o[1120] = (N3)? mem[1120] : 
                          (N0)? mem[2720] : 1'b0;
  assign r_data_o[1119] = (N3)? mem[1119] : 
                          (N0)? mem[2719] : 1'b0;
  assign r_data_o[1118] = (N3)? mem[1118] : 
                          (N0)? mem[2718] : 1'b0;
  assign r_data_o[1117] = (N3)? mem[1117] : 
                          (N0)? mem[2717] : 1'b0;
  assign r_data_o[1116] = (N3)? mem[1116] : 
                          (N0)? mem[2716] : 1'b0;
  assign r_data_o[1115] = (N3)? mem[1115] : 
                          (N0)? mem[2715] : 1'b0;
  assign r_data_o[1114] = (N3)? mem[1114] : 
                          (N0)? mem[2714] : 1'b0;
  assign r_data_o[1113] = (N3)? mem[1113] : 
                          (N0)? mem[2713] : 1'b0;
  assign r_data_o[1112] = (N3)? mem[1112] : 
                          (N0)? mem[2712] : 1'b0;
  assign r_data_o[1111] = (N3)? mem[1111] : 
                          (N0)? mem[2711] : 1'b0;
  assign r_data_o[1110] = (N3)? mem[1110] : 
                          (N0)? mem[2710] : 1'b0;
  assign r_data_o[1109] = (N3)? mem[1109] : 
                          (N0)? mem[2709] : 1'b0;
  assign r_data_o[1108] = (N3)? mem[1108] : 
                          (N0)? mem[2708] : 1'b0;
  assign r_data_o[1107] = (N3)? mem[1107] : 
                          (N0)? mem[2707] : 1'b0;
  assign r_data_o[1106] = (N3)? mem[1106] : 
                          (N0)? mem[2706] : 1'b0;
  assign r_data_o[1105] = (N3)? mem[1105] : 
                          (N0)? mem[2705] : 1'b0;
  assign r_data_o[1104] = (N3)? mem[1104] : 
                          (N0)? mem[2704] : 1'b0;
  assign r_data_o[1103] = (N3)? mem[1103] : 
                          (N0)? mem[2703] : 1'b0;
  assign r_data_o[1102] = (N3)? mem[1102] : 
                          (N0)? mem[2702] : 1'b0;
  assign r_data_o[1101] = (N3)? mem[1101] : 
                          (N0)? mem[2701] : 1'b0;
  assign r_data_o[1100] = (N3)? mem[1100] : 
                          (N0)? mem[2700] : 1'b0;
  assign r_data_o[1099] = (N3)? mem[1099] : 
                          (N0)? mem[2699] : 1'b0;
  assign r_data_o[1098] = (N3)? mem[1098] : 
                          (N0)? mem[2698] : 1'b0;
  assign r_data_o[1097] = (N3)? mem[1097] : 
                          (N0)? mem[2697] : 1'b0;
  assign r_data_o[1096] = (N3)? mem[1096] : 
                          (N0)? mem[2696] : 1'b0;
  assign r_data_o[1095] = (N3)? mem[1095] : 
                          (N0)? mem[2695] : 1'b0;
  assign r_data_o[1094] = (N3)? mem[1094] : 
                          (N0)? mem[2694] : 1'b0;
  assign r_data_o[1093] = (N3)? mem[1093] : 
                          (N0)? mem[2693] : 1'b0;
  assign r_data_o[1092] = (N3)? mem[1092] : 
                          (N0)? mem[2692] : 1'b0;
  assign r_data_o[1091] = (N3)? mem[1091] : 
                          (N0)? mem[2691] : 1'b0;
  assign r_data_o[1090] = (N3)? mem[1090] : 
                          (N0)? mem[2690] : 1'b0;
  assign r_data_o[1089] = (N3)? mem[1089] : 
                          (N0)? mem[2689] : 1'b0;
  assign r_data_o[1088] = (N3)? mem[1088] : 
                          (N0)? mem[2688] : 1'b0;
  assign r_data_o[1087] = (N3)? mem[1087] : 
                          (N0)? mem[2687] : 1'b0;
  assign r_data_o[1086] = (N3)? mem[1086] : 
                          (N0)? mem[2686] : 1'b0;
  assign r_data_o[1085] = (N3)? mem[1085] : 
                          (N0)? mem[2685] : 1'b0;
  assign r_data_o[1084] = (N3)? mem[1084] : 
                          (N0)? mem[2684] : 1'b0;
  assign r_data_o[1083] = (N3)? mem[1083] : 
                          (N0)? mem[2683] : 1'b0;
  assign r_data_o[1082] = (N3)? mem[1082] : 
                          (N0)? mem[2682] : 1'b0;
  assign r_data_o[1081] = (N3)? mem[1081] : 
                          (N0)? mem[2681] : 1'b0;
  assign r_data_o[1080] = (N3)? mem[1080] : 
                          (N0)? mem[2680] : 1'b0;
  assign r_data_o[1079] = (N3)? mem[1079] : 
                          (N0)? mem[2679] : 1'b0;
  assign r_data_o[1078] = (N3)? mem[1078] : 
                          (N0)? mem[2678] : 1'b0;
  assign r_data_o[1077] = (N3)? mem[1077] : 
                          (N0)? mem[2677] : 1'b0;
  assign r_data_o[1076] = (N3)? mem[1076] : 
                          (N0)? mem[2676] : 1'b0;
  assign r_data_o[1075] = (N3)? mem[1075] : 
                          (N0)? mem[2675] : 1'b0;
  assign r_data_o[1074] = (N3)? mem[1074] : 
                          (N0)? mem[2674] : 1'b0;
  assign r_data_o[1073] = (N3)? mem[1073] : 
                          (N0)? mem[2673] : 1'b0;
  assign r_data_o[1072] = (N3)? mem[1072] : 
                          (N0)? mem[2672] : 1'b0;
  assign r_data_o[1071] = (N3)? mem[1071] : 
                          (N0)? mem[2671] : 1'b0;
  assign r_data_o[1070] = (N3)? mem[1070] : 
                          (N0)? mem[2670] : 1'b0;
  assign r_data_o[1069] = (N3)? mem[1069] : 
                          (N0)? mem[2669] : 1'b0;
  assign r_data_o[1068] = (N3)? mem[1068] : 
                          (N0)? mem[2668] : 1'b0;
  assign r_data_o[1067] = (N3)? mem[1067] : 
                          (N0)? mem[2667] : 1'b0;
  assign r_data_o[1066] = (N3)? mem[1066] : 
                          (N0)? mem[2666] : 1'b0;
  assign r_data_o[1065] = (N3)? mem[1065] : 
                          (N0)? mem[2665] : 1'b0;
  assign r_data_o[1064] = (N3)? mem[1064] : 
                          (N0)? mem[2664] : 1'b0;
  assign r_data_o[1063] = (N3)? mem[1063] : 
                          (N0)? mem[2663] : 1'b0;
  assign r_data_o[1062] = (N3)? mem[1062] : 
                          (N0)? mem[2662] : 1'b0;
  assign r_data_o[1061] = (N3)? mem[1061] : 
                          (N0)? mem[2661] : 1'b0;
  assign r_data_o[1060] = (N3)? mem[1060] : 
                          (N0)? mem[2660] : 1'b0;
  assign r_data_o[1059] = (N3)? mem[1059] : 
                          (N0)? mem[2659] : 1'b0;
  assign r_data_o[1058] = (N3)? mem[1058] : 
                          (N0)? mem[2658] : 1'b0;
  assign r_data_o[1057] = (N3)? mem[1057] : 
                          (N0)? mem[2657] : 1'b0;
  assign r_data_o[1056] = (N3)? mem[1056] : 
                          (N0)? mem[2656] : 1'b0;
  assign r_data_o[1055] = (N3)? mem[1055] : 
                          (N0)? mem[2655] : 1'b0;
  assign r_data_o[1054] = (N3)? mem[1054] : 
                          (N0)? mem[2654] : 1'b0;
  assign r_data_o[1053] = (N3)? mem[1053] : 
                          (N0)? mem[2653] : 1'b0;
  assign r_data_o[1052] = (N3)? mem[1052] : 
                          (N0)? mem[2652] : 1'b0;
  assign r_data_o[1051] = (N3)? mem[1051] : 
                          (N0)? mem[2651] : 1'b0;
  assign r_data_o[1050] = (N3)? mem[1050] : 
                          (N0)? mem[2650] : 1'b0;
  assign r_data_o[1049] = (N3)? mem[1049] : 
                          (N0)? mem[2649] : 1'b0;
  assign r_data_o[1048] = (N3)? mem[1048] : 
                          (N0)? mem[2648] : 1'b0;
  assign r_data_o[1047] = (N3)? mem[1047] : 
                          (N0)? mem[2647] : 1'b0;
  assign r_data_o[1046] = (N3)? mem[1046] : 
                          (N0)? mem[2646] : 1'b0;
  assign r_data_o[1045] = (N3)? mem[1045] : 
                          (N0)? mem[2645] : 1'b0;
  assign r_data_o[1044] = (N3)? mem[1044] : 
                          (N0)? mem[2644] : 1'b0;
  assign r_data_o[1043] = (N3)? mem[1043] : 
                          (N0)? mem[2643] : 1'b0;
  assign r_data_o[1042] = (N3)? mem[1042] : 
                          (N0)? mem[2642] : 1'b0;
  assign r_data_o[1041] = (N3)? mem[1041] : 
                          (N0)? mem[2641] : 1'b0;
  assign r_data_o[1040] = (N3)? mem[1040] : 
                          (N0)? mem[2640] : 1'b0;
  assign r_data_o[1039] = (N3)? mem[1039] : 
                          (N0)? mem[2639] : 1'b0;
  assign r_data_o[1038] = (N3)? mem[1038] : 
                          (N0)? mem[2638] : 1'b0;
  assign r_data_o[1037] = (N3)? mem[1037] : 
                          (N0)? mem[2637] : 1'b0;
  assign r_data_o[1036] = (N3)? mem[1036] : 
                          (N0)? mem[2636] : 1'b0;
  assign r_data_o[1035] = (N3)? mem[1035] : 
                          (N0)? mem[2635] : 1'b0;
  assign r_data_o[1034] = (N3)? mem[1034] : 
                          (N0)? mem[2634] : 1'b0;
  assign r_data_o[1033] = (N3)? mem[1033] : 
                          (N0)? mem[2633] : 1'b0;
  assign r_data_o[1032] = (N3)? mem[1032] : 
                          (N0)? mem[2632] : 1'b0;
  assign r_data_o[1031] = (N3)? mem[1031] : 
                          (N0)? mem[2631] : 1'b0;
  assign r_data_o[1030] = (N3)? mem[1030] : 
                          (N0)? mem[2630] : 1'b0;
  assign r_data_o[1029] = (N3)? mem[1029] : 
                          (N0)? mem[2629] : 1'b0;
  assign r_data_o[1028] = (N3)? mem[1028] : 
                          (N0)? mem[2628] : 1'b0;
  assign r_data_o[1027] = (N3)? mem[1027] : 
                          (N0)? mem[2627] : 1'b0;
  assign r_data_o[1026] = (N3)? mem[1026] : 
                          (N0)? mem[2626] : 1'b0;
  assign r_data_o[1025] = (N3)? mem[1025] : 
                          (N0)? mem[2625] : 1'b0;
  assign r_data_o[1024] = (N3)? mem[1024] : 
                          (N0)? mem[2624] : 1'b0;
  assign r_data_o[1023] = (N3)? mem[1023] : 
                          (N0)? mem[2623] : 1'b0;
  assign r_data_o[1022] = (N3)? mem[1022] : 
                          (N0)? mem[2622] : 1'b0;
  assign r_data_o[1021] = (N3)? mem[1021] : 
                          (N0)? mem[2621] : 1'b0;
  assign r_data_o[1020] = (N3)? mem[1020] : 
                          (N0)? mem[2620] : 1'b0;
  assign r_data_o[1019] = (N3)? mem[1019] : 
                          (N0)? mem[2619] : 1'b0;
  assign r_data_o[1018] = (N3)? mem[1018] : 
                          (N0)? mem[2618] : 1'b0;
  assign r_data_o[1017] = (N3)? mem[1017] : 
                          (N0)? mem[2617] : 1'b0;
  assign r_data_o[1016] = (N3)? mem[1016] : 
                          (N0)? mem[2616] : 1'b0;
  assign r_data_o[1015] = (N3)? mem[1015] : 
                          (N0)? mem[2615] : 1'b0;
  assign r_data_o[1014] = (N3)? mem[1014] : 
                          (N0)? mem[2614] : 1'b0;
  assign r_data_o[1013] = (N3)? mem[1013] : 
                          (N0)? mem[2613] : 1'b0;
  assign r_data_o[1012] = (N3)? mem[1012] : 
                          (N0)? mem[2612] : 1'b0;
  assign r_data_o[1011] = (N3)? mem[1011] : 
                          (N0)? mem[2611] : 1'b0;
  assign r_data_o[1010] = (N3)? mem[1010] : 
                          (N0)? mem[2610] : 1'b0;
  assign r_data_o[1009] = (N3)? mem[1009] : 
                          (N0)? mem[2609] : 1'b0;
  assign r_data_o[1008] = (N3)? mem[1008] : 
                          (N0)? mem[2608] : 1'b0;
  assign r_data_o[1007] = (N3)? mem[1007] : 
                          (N0)? mem[2607] : 1'b0;
  assign r_data_o[1006] = (N3)? mem[1006] : 
                          (N0)? mem[2606] : 1'b0;
  assign r_data_o[1005] = (N3)? mem[1005] : 
                          (N0)? mem[2605] : 1'b0;
  assign r_data_o[1004] = (N3)? mem[1004] : 
                          (N0)? mem[2604] : 1'b0;
  assign r_data_o[1003] = (N3)? mem[1003] : 
                          (N0)? mem[2603] : 1'b0;
  assign r_data_o[1002] = (N3)? mem[1002] : 
                          (N0)? mem[2602] : 1'b0;
  assign r_data_o[1001] = (N3)? mem[1001] : 
                          (N0)? mem[2601] : 1'b0;
  assign r_data_o[1000] = (N3)? mem[1000] : 
                          (N0)? mem[2600] : 1'b0;
  assign r_data_o[999] = (N3)? mem[999] : 
                         (N0)? mem[2599] : 1'b0;
  assign r_data_o[998] = (N3)? mem[998] : 
                         (N0)? mem[2598] : 1'b0;
  assign r_data_o[997] = (N3)? mem[997] : 
                         (N0)? mem[2597] : 1'b0;
  assign r_data_o[996] = (N3)? mem[996] : 
                         (N0)? mem[2596] : 1'b0;
  assign r_data_o[995] = (N3)? mem[995] : 
                         (N0)? mem[2595] : 1'b0;
  assign r_data_o[994] = (N3)? mem[994] : 
                         (N0)? mem[2594] : 1'b0;
  assign r_data_o[993] = (N3)? mem[993] : 
                         (N0)? mem[2593] : 1'b0;
  assign r_data_o[992] = (N3)? mem[992] : 
                         (N0)? mem[2592] : 1'b0;
  assign r_data_o[991] = (N3)? mem[991] : 
                         (N0)? mem[2591] : 1'b0;
  assign r_data_o[990] = (N3)? mem[990] : 
                         (N0)? mem[2590] : 1'b0;
  assign r_data_o[989] = (N3)? mem[989] : 
                         (N0)? mem[2589] : 1'b0;
  assign r_data_o[988] = (N3)? mem[988] : 
                         (N0)? mem[2588] : 1'b0;
  assign r_data_o[987] = (N3)? mem[987] : 
                         (N0)? mem[2587] : 1'b0;
  assign r_data_o[986] = (N3)? mem[986] : 
                         (N0)? mem[2586] : 1'b0;
  assign r_data_o[985] = (N3)? mem[985] : 
                         (N0)? mem[2585] : 1'b0;
  assign r_data_o[984] = (N3)? mem[984] : 
                         (N0)? mem[2584] : 1'b0;
  assign r_data_o[983] = (N3)? mem[983] : 
                         (N0)? mem[2583] : 1'b0;
  assign r_data_o[982] = (N3)? mem[982] : 
                         (N0)? mem[2582] : 1'b0;
  assign r_data_o[981] = (N3)? mem[981] : 
                         (N0)? mem[2581] : 1'b0;
  assign r_data_o[980] = (N3)? mem[980] : 
                         (N0)? mem[2580] : 1'b0;
  assign r_data_o[979] = (N3)? mem[979] : 
                         (N0)? mem[2579] : 1'b0;
  assign r_data_o[978] = (N3)? mem[978] : 
                         (N0)? mem[2578] : 1'b0;
  assign r_data_o[977] = (N3)? mem[977] : 
                         (N0)? mem[2577] : 1'b0;
  assign r_data_o[976] = (N3)? mem[976] : 
                         (N0)? mem[2576] : 1'b0;
  assign r_data_o[975] = (N3)? mem[975] : 
                         (N0)? mem[2575] : 1'b0;
  assign r_data_o[974] = (N3)? mem[974] : 
                         (N0)? mem[2574] : 1'b0;
  assign r_data_o[973] = (N3)? mem[973] : 
                         (N0)? mem[2573] : 1'b0;
  assign r_data_o[972] = (N3)? mem[972] : 
                         (N0)? mem[2572] : 1'b0;
  assign r_data_o[971] = (N3)? mem[971] : 
                         (N0)? mem[2571] : 1'b0;
  assign r_data_o[970] = (N3)? mem[970] : 
                         (N0)? mem[2570] : 1'b0;
  assign r_data_o[969] = (N3)? mem[969] : 
                         (N0)? mem[2569] : 1'b0;
  assign r_data_o[968] = (N3)? mem[968] : 
                         (N0)? mem[2568] : 1'b0;
  assign r_data_o[967] = (N3)? mem[967] : 
                         (N0)? mem[2567] : 1'b0;
  assign r_data_o[966] = (N3)? mem[966] : 
                         (N0)? mem[2566] : 1'b0;
  assign r_data_o[965] = (N3)? mem[965] : 
                         (N0)? mem[2565] : 1'b0;
  assign r_data_o[964] = (N3)? mem[964] : 
                         (N0)? mem[2564] : 1'b0;
  assign r_data_o[963] = (N3)? mem[963] : 
                         (N0)? mem[2563] : 1'b0;
  assign r_data_o[962] = (N3)? mem[962] : 
                         (N0)? mem[2562] : 1'b0;
  assign r_data_o[961] = (N3)? mem[961] : 
                         (N0)? mem[2561] : 1'b0;
  assign r_data_o[960] = (N3)? mem[960] : 
                         (N0)? mem[2560] : 1'b0;
  assign r_data_o[959] = (N3)? mem[959] : 
                         (N0)? mem[2559] : 1'b0;
  assign r_data_o[958] = (N3)? mem[958] : 
                         (N0)? mem[2558] : 1'b0;
  assign r_data_o[957] = (N3)? mem[957] : 
                         (N0)? mem[2557] : 1'b0;
  assign r_data_o[956] = (N3)? mem[956] : 
                         (N0)? mem[2556] : 1'b0;
  assign r_data_o[955] = (N3)? mem[955] : 
                         (N0)? mem[2555] : 1'b0;
  assign r_data_o[954] = (N3)? mem[954] : 
                         (N0)? mem[2554] : 1'b0;
  assign r_data_o[953] = (N3)? mem[953] : 
                         (N0)? mem[2553] : 1'b0;
  assign r_data_o[952] = (N3)? mem[952] : 
                         (N0)? mem[2552] : 1'b0;
  assign r_data_o[951] = (N3)? mem[951] : 
                         (N0)? mem[2551] : 1'b0;
  assign r_data_o[950] = (N3)? mem[950] : 
                         (N0)? mem[2550] : 1'b0;
  assign r_data_o[949] = (N3)? mem[949] : 
                         (N0)? mem[2549] : 1'b0;
  assign r_data_o[948] = (N3)? mem[948] : 
                         (N0)? mem[2548] : 1'b0;
  assign r_data_o[947] = (N3)? mem[947] : 
                         (N0)? mem[2547] : 1'b0;
  assign r_data_o[946] = (N3)? mem[946] : 
                         (N0)? mem[2546] : 1'b0;
  assign r_data_o[945] = (N3)? mem[945] : 
                         (N0)? mem[2545] : 1'b0;
  assign r_data_o[944] = (N3)? mem[944] : 
                         (N0)? mem[2544] : 1'b0;
  assign r_data_o[943] = (N3)? mem[943] : 
                         (N0)? mem[2543] : 1'b0;
  assign r_data_o[942] = (N3)? mem[942] : 
                         (N0)? mem[2542] : 1'b0;
  assign r_data_o[941] = (N3)? mem[941] : 
                         (N0)? mem[2541] : 1'b0;
  assign r_data_o[940] = (N3)? mem[940] : 
                         (N0)? mem[2540] : 1'b0;
  assign r_data_o[939] = (N3)? mem[939] : 
                         (N0)? mem[2539] : 1'b0;
  assign r_data_o[938] = (N3)? mem[938] : 
                         (N0)? mem[2538] : 1'b0;
  assign r_data_o[937] = (N3)? mem[937] : 
                         (N0)? mem[2537] : 1'b0;
  assign r_data_o[936] = (N3)? mem[936] : 
                         (N0)? mem[2536] : 1'b0;
  assign r_data_o[935] = (N3)? mem[935] : 
                         (N0)? mem[2535] : 1'b0;
  assign r_data_o[934] = (N3)? mem[934] : 
                         (N0)? mem[2534] : 1'b0;
  assign r_data_o[933] = (N3)? mem[933] : 
                         (N0)? mem[2533] : 1'b0;
  assign r_data_o[932] = (N3)? mem[932] : 
                         (N0)? mem[2532] : 1'b0;
  assign r_data_o[931] = (N3)? mem[931] : 
                         (N0)? mem[2531] : 1'b0;
  assign r_data_o[930] = (N3)? mem[930] : 
                         (N0)? mem[2530] : 1'b0;
  assign r_data_o[929] = (N3)? mem[929] : 
                         (N0)? mem[2529] : 1'b0;
  assign r_data_o[928] = (N3)? mem[928] : 
                         (N0)? mem[2528] : 1'b0;
  assign r_data_o[927] = (N3)? mem[927] : 
                         (N0)? mem[2527] : 1'b0;
  assign r_data_o[926] = (N3)? mem[926] : 
                         (N0)? mem[2526] : 1'b0;
  assign r_data_o[925] = (N3)? mem[925] : 
                         (N0)? mem[2525] : 1'b0;
  assign r_data_o[924] = (N3)? mem[924] : 
                         (N0)? mem[2524] : 1'b0;
  assign r_data_o[923] = (N3)? mem[923] : 
                         (N0)? mem[2523] : 1'b0;
  assign r_data_o[922] = (N3)? mem[922] : 
                         (N0)? mem[2522] : 1'b0;
  assign r_data_o[921] = (N3)? mem[921] : 
                         (N0)? mem[2521] : 1'b0;
  assign r_data_o[920] = (N3)? mem[920] : 
                         (N0)? mem[2520] : 1'b0;
  assign r_data_o[919] = (N3)? mem[919] : 
                         (N0)? mem[2519] : 1'b0;
  assign r_data_o[918] = (N3)? mem[918] : 
                         (N0)? mem[2518] : 1'b0;
  assign r_data_o[917] = (N3)? mem[917] : 
                         (N0)? mem[2517] : 1'b0;
  assign r_data_o[916] = (N3)? mem[916] : 
                         (N0)? mem[2516] : 1'b0;
  assign r_data_o[915] = (N3)? mem[915] : 
                         (N0)? mem[2515] : 1'b0;
  assign r_data_o[914] = (N3)? mem[914] : 
                         (N0)? mem[2514] : 1'b0;
  assign r_data_o[913] = (N3)? mem[913] : 
                         (N0)? mem[2513] : 1'b0;
  assign r_data_o[912] = (N3)? mem[912] : 
                         (N0)? mem[2512] : 1'b0;
  assign r_data_o[911] = (N3)? mem[911] : 
                         (N0)? mem[2511] : 1'b0;
  assign r_data_o[910] = (N3)? mem[910] : 
                         (N0)? mem[2510] : 1'b0;
  assign r_data_o[909] = (N3)? mem[909] : 
                         (N0)? mem[2509] : 1'b0;
  assign r_data_o[908] = (N3)? mem[908] : 
                         (N0)? mem[2508] : 1'b0;
  assign r_data_o[907] = (N3)? mem[907] : 
                         (N0)? mem[2507] : 1'b0;
  assign r_data_o[906] = (N3)? mem[906] : 
                         (N0)? mem[2506] : 1'b0;
  assign r_data_o[905] = (N3)? mem[905] : 
                         (N0)? mem[2505] : 1'b0;
  assign r_data_o[904] = (N3)? mem[904] : 
                         (N0)? mem[2504] : 1'b0;
  assign r_data_o[903] = (N3)? mem[903] : 
                         (N0)? mem[2503] : 1'b0;
  assign r_data_o[902] = (N3)? mem[902] : 
                         (N0)? mem[2502] : 1'b0;
  assign r_data_o[901] = (N3)? mem[901] : 
                         (N0)? mem[2501] : 1'b0;
  assign r_data_o[900] = (N3)? mem[900] : 
                         (N0)? mem[2500] : 1'b0;
  assign r_data_o[899] = (N3)? mem[899] : 
                         (N0)? mem[2499] : 1'b0;
  assign r_data_o[898] = (N3)? mem[898] : 
                         (N0)? mem[2498] : 1'b0;
  assign r_data_o[897] = (N3)? mem[897] : 
                         (N0)? mem[2497] : 1'b0;
  assign r_data_o[896] = (N3)? mem[896] : 
                         (N0)? mem[2496] : 1'b0;
  assign r_data_o[895] = (N3)? mem[895] : 
                         (N0)? mem[2495] : 1'b0;
  assign r_data_o[894] = (N3)? mem[894] : 
                         (N0)? mem[2494] : 1'b0;
  assign r_data_o[893] = (N3)? mem[893] : 
                         (N0)? mem[2493] : 1'b0;
  assign r_data_o[892] = (N3)? mem[892] : 
                         (N0)? mem[2492] : 1'b0;
  assign r_data_o[891] = (N3)? mem[891] : 
                         (N0)? mem[2491] : 1'b0;
  assign r_data_o[890] = (N3)? mem[890] : 
                         (N0)? mem[2490] : 1'b0;
  assign r_data_o[889] = (N3)? mem[889] : 
                         (N0)? mem[2489] : 1'b0;
  assign r_data_o[888] = (N3)? mem[888] : 
                         (N0)? mem[2488] : 1'b0;
  assign r_data_o[887] = (N3)? mem[887] : 
                         (N0)? mem[2487] : 1'b0;
  assign r_data_o[886] = (N3)? mem[886] : 
                         (N0)? mem[2486] : 1'b0;
  assign r_data_o[885] = (N3)? mem[885] : 
                         (N0)? mem[2485] : 1'b0;
  assign r_data_o[884] = (N3)? mem[884] : 
                         (N0)? mem[2484] : 1'b0;
  assign r_data_o[883] = (N3)? mem[883] : 
                         (N0)? mem[2483] : 1'b0;
  assign r_data_o[882] = (N3)? mem[882] : 
                         (N0)? mem[2482] : 1'b0;
  assign r_data_o[881] = (N3)? mem[881] : 
                         (N0)? mem[2481] : 1'b0;
  assign r_data_o[880] = (N3)? mem[880] : 
                         (N0)? mem[2480] : 1'b0;
  assign r_data_o[879] = (N3)? mem[879] : 
                         (N0)? mem[2479] : 1'b0;
  assign r_data_o[878] = (N3)? mem[878] : 
                         (N0)? mem[2478] : 1'b0;
  assign r_data_o[877] = (N3)? mem[877] : 
                         (N0)? mem[2477] : 1'b0;
  assign r_data_o[876] = (N3)? mem[876] : 
                         (N0)? mem[2476] : 1'b0;
  assign r_data_o[875] = (N3)? mem[875] : 
                         (N0)? mem[2475] : 1'b0;
  assign r_data_o[874] = (N3)? mem[874] : 
                         (N0)? mem[2474] : 1'b0;
  assign r_data_o[873] = (N3)? mem[873] : 
                         (N0)? mem[2473] : 1'b0;
  assign r_data_o[872] = (N3)? mem[872] : 
                         (N0)? mem[2472] : 1'b0;
  assign r_data_o[871] = (N3)? mem[871] : 
                         (N0)? mem[2471] : 1'b0;
  assign r_data_o[870] = (N3)? mem[870] : 
                         (N0)? mem[2470] : 1'b0;
  assign r_data_o[869] = (N3)? mem[869] : 
                         (N0)? mem[2469] : 1'b0;
  assign r_data_o[868] = (N3)? mem[868] : 
                         (N0)? mem[2468] : 1'b0;
  assign r_data_o[867] = (N3)? mem[867] : 
                         (N0)? mem[2467] : 1'b0;
  assign r_data_o[866] = (N3)? mem[866] : 
                         (N0)? mem[2466] : 1'b0;
  assign r_data_o[865] = (N3)? mem[865] : 
                         (N0)? mem[2465] : 1'b0;
  assign r_data_o[864] = (N3)? mem[864] : 
                         (N0)? mem[2464] : 1'b0;
  assign r_data_o[863] = (N3)? mem[863] : 
                         (N0)? mem[2463] : 1'b0;
  assign r_data_o[862] = (N3)? mem[862] : 
                         (N0)? mem[2462] : 1'b0;
  assign r_data_o[861] = (N3)? mem[861] : 
                         (N0)? mem[2461] : 1'b0;
  assign r_data_o[860] = (N3)? mem[860] : 
                         (N0)? mem[2460] : 1'b0;
  assign r_data_o[859] = (N3)? mem[859] : 
                         (N0)? mem[2459] : 1'b0;
  assign r_data_o[858] = (N3)? mem[858] : 
                         (N0)? mem[2458] : 1'b0;
  assign r_data_o[857] = (N3)? mem[857] : 
                         (N0)? mem[2457] : 1'b0;
  assign r_data_o[856] = (N3)? mem[856] : 
                         (N0)? mem[2456] : 1'b0;
  assign r_data_o[855] = (N3)? mem[855] : 
                         (N0)? mem[2455] : 1'b0;
  assign r_data_o[854] = (N3)? mem[854] : 
                         (N0)? mem[2454] : 1'b0;
  assign r_data_o[853] = (N3)? mem[853] : 
                         (N0)? mem[2453] : 1'b0;
  assign r_data_o[852] = (N3)? mem[852] : 
                         (N0)? mem[2452] : 1'b0;
  assign r_data_o[851] = (N3)? mem[851] : 
                         (N0)? mem[2451] : 1'b0;
  assign r_data_o[850] = (N3)? mem[850] : 
                         (N0)? mem[2450] : 1'b0;
  assign r_data_o[849] = (N3)? mem[849] : 
                         (N0)? mem[2449] : 1'b0;
  assign r_data_o[848] = (N3)? mem[848] : 
                         (N0)? mem[2448] : 1'b0;
  assign r_data_o[847] = (N3)? mem[847] : 
                         (N0)? mem[2447] : 1'b0;
  assign r_data_o[846] = (N3)? mem[846] : 
                         (N0)? mem[2446] : 1'b0;
  assign r_data_o[845] = (N3)? mem[845] : 
                         (N0)? mem[2445] : 1'b0;
  assign r_data_o[844] = (N3)? mem[844] : 
                         (N0)? mem[2444] : 1'b0;
  assign r_data_o[843] = (N3)? mem[843] : 
                         (N0)? mem[2443] : 1'b0;
  assign r_data_o[842] = (N3)? mem[842] : 
                         (N0)? mem[2442] : 1'b0;
  assign r_data_o[841] = (N3)? mem[841] : 
                         (N0)? mem[2441] : 1'b0;
  assign r_data_o[840] = (N3)? mem[840] : 
                         (N0)? mem[2440] : 1'b0;
  assign r_data_o[839] = (N3)? mem[839] : 
                         (N0)? mem[2439] : 1'b0;
  assign r_data_o[838] = (N3)? mem[838] : 
                         (N0)? mem[2438] : 1'b0;
  assign r_data_o[837] = (N3)? mem[837] : 
                         (N0)? mem[2437] : 1'b0;
  assign r_data_o[836] = (N3)? mem[836] : 
                         (N0)? mem[2436] : 1'b0;
  assign r_data_o[835] = (N3)? mem[835] : 
                         (N0)? mem[2435] : 1'b0;
  assign r_data_o[834] = (N3)? mem[834] : 
                         (N0)? mem[2434] : 1'b0;
  assign r_data_o[833] = (N3)? mem[833] : 
                         (N0)? mem[2433] : 1'b0;
  assign r_data_o[832] = (N3)? mem[832] : 
                         (N0)? mem[2432] : 1'b0;
  assign r_data_o[831] = (N3)? mem[831] : 
                         (N0)? mem[2431] : 1'b0;
  assign r_data_o[830] = (N3)? mem[830] : 
                         (N0)? mem[2430] : 1'b0;
  assign r_data_o[829] = (N3)? mem[829] : 
                         (N0)? mem[2429] : 1'b0;
  assign r_data_o[828] = (N3)? mem[828] : 
                         (N0)? mem[2428] : 1'b0;
  assign r_data_o[827] = (N3)? mem[827] : 
                         (N0)? mem[2427] : 1'b0;
  assign r_data_o[826] = (N3)? mem[826] : 
                         (N0)? mem[2426] : 1'b0;
  assign r_data_o[825] = (N3)? mem[825] : 
                         (N0)? mem[2425] : 1'b0;
  assign r_data_o[824] = (N3)? mem[824] : 
                         (N0)? mem[2424] : 1'b0;
  assign r_data_o[823] = (N3)? mem[823] : 
                         (N0)? mem[2423] : 1'b0;
  assign r_data_o[822] = (N3)? mem[822] : 
                         (N0)? mem[2422] : 1'b0;
  assign r_data_o[821] = (N3)? mem[821] : 
                         (N0)? mem[2421] : 1'b0;
  assign r_data_o[820] = (N3)? mem[820] : 
                         (N0)? mem[2420] : 1'b0;
  assign r_data_o[819] = (N3)? mem[819] : 
                         (N0)? mem[2419] : 1'b0;
  assign r_data_o[818] = (N3)? mem[818] : 
                         (N0)? mem[2418] : 1'b0;
  assign r_data_o[817] = (N3)? mem[817] : 
                         (N0)? mem[2417] : 1'b0;
  assign r_data_o[816] = (N3)? mem[816] : 
                         (N0)? mem[2416] : 1'b0;
  assign r_data_o[815] = (N3)? mem[815] : 
                         (N0)? mem[2415] : 1'b0;
  assign r_data_o[814] = (N3)? mem[814] : 
                         (N0)? mem[2414] : 1'b0;
  assign r_data_o[813] = (N3)? mem[813] : 
                         (N0)? mem[2413] : 1'b0;
  assign r_data_o[812] = (N3)? mem[812] : 
                         (N0)? mem[2412] : 1'b0;
  assign r_data_o[811] = (N3)? mem[811] : 
                         (N0)? mem[2411] : 1'b0;
  assign r_data_o[810] = (N3)? mem[810] : 
                         (N0)? mem[2410] : 1'b0;
  assign r_data_o[809] = (N3)? mem[809] : 
                         (N0)? mem[2409] : 1'b0;
  assign r_data_o[808] = (N3)? mem[808] : 
                         (N0)? mem[2408] : 1'b0;
  assign r_data_o[807] = (N3)? mem[807] : 
                         (N0)? mem[2407] : 1'b0;
  assign r_data_o[806] = (N3)? mem[806] : 
                         (N0)? mem[2406] : 1'b0;
  assign r_data_o[805] = (N3)? mem[805] : 
                         (N0)? mem[2405] : 1'b0;
  assign r_data_o[804] = (N3)? mem[804] : 
                         (N0)? mem[2404] : 1'b0;
  assign r_data_o[803] = (N3)? mem[803] : 
                         (N0)? mem[2403] : 1'b0;
  assign r_data_o[802] = (N3)? mem[802] : 
                         (N0)? mem[2402] : 1'b0;
  assign r_data_o[801] = (N3)? mem[801] : 
                         (N0)? mem[2401] : 1'b0;
  assign r_data_o[800] = (N3)? mem[800] : 
                         (N0)? mem[2400] : 1'b0;
  assign r_data_o[799] = (N3)? mem[799] : 
                         (N0)? mem[2399] : 1'b0;
  assign r_data_o[798] = (N3)? mem[798] : 
                         (N0)? mem[2398] : 1'b0;
  assign r_data_o[797] = (N3)? mem[797] : 
                         (N0)? mem[2397] : 1'b0;
  assign r_data_o[796] = (N3)? mem[796] : 
                         (N0)? mem[2396] : 1'b0;
  assign r_data_o[795] = (N3)? mem[795] : 
                         (N0)? mem[2395] : 1'b0;
  assign r_data_o[794] = (N3)? mem[794] : 
                         (N0)? mem[2394] : 1'b0;
  assign r_data_o[793] = (N3)? mem[793] : 
                         (N0)? mem[2393] : 1'b0;
  assign r_data_o[792] = (N3)? mem[792] : 
                         (N0)? mem[2392] : 1'b0;
  assign r_data_o[791] = (N3)? mem[791] : 
                         (N0)? mem[2391] : 1'b0;
  assign r_data_o[790] = (N3)? mem[790] : 
                         (N0)? mem[2390] : 1'b0;
  assign r_data_o[789] = (N3)? mem[789] : 
                         (N0)? mem[2389] : 1'b0;
  assign r_data_o[788] = (N3)? mem[788] : 
                         (N0)? mem[2388] : 1'b0;
  assign r_data_o[787] = (N3)? mem[787] : 
                         (N0)? mem[2387] : 1'b0;
  assign r_data_o[786] = (N3)? mem[786] : 
                         (N0)? mem[2386] : 1'b0;
  assign r_data_o[785] = (N3)? mem[785] : 
                         (N0)? mem[2385] : 1'b0;
  assign r_data_o[784] = (N3)? mem[784] : 
                         (N0)? mem[2384] : 1'b0;
  assign r_data_o[783] = (N3)? mem[783] : 
                         (N0)? mem[2383] : 1'b0;
  assign r_data_o[782] = (N3)? mem[782] : 
                         (N0)? mem[2382] : 1'b0;
  assign r_data_o[781] = (N3)? mem[781] : 
                         (N0)? mem[2381] : 1'b0;
  assign r_data_o[780] = (N3)? mem[780] : 
                         (N0)? mem[2380] : 1'b0;
  assign r_data_o[779] = (N3)? mem[779] : 
                         (N0)? mem[2379] : 1'b0;
  assign r_data_o[778] = (N3)? mem[778] : 
                         (N0)? mem[2378] : 1'b0;
  assign r_data_o[777] = (N3)? mem[777] : 
                         (N0)? mem[2377] : 1'b0;
  assign r_data_o[776] = (N3)? mem[776] : 
                         (N0)? mem[2376] : 1'b0;
  assign r_data_o[775] = (N3)? mem[775] : 
                         (N0)? mem[2375] : 1'b0;
  assign r_data_o[774] = (N3)? mem[774] : 
                         (N0)? mem[2374] : 1'b0;
  assign r_data_o[773] = (N3)? mem[773] : 
                         (N0)? mem[2373] : 1'b0;
  assign r_data_o[772] = (N3)? mem[772] : 
                         (N0)? mem[2372] : 1'b0;
  assign r_data_o[771] = (N3)? mem[771] : 
                         (N0)? mem[2371] : 1'b0;
  assign r_data_o[770] = (N3)? mem[770] : 
                         (N0)? mem[2370] : 1'b0;
  assign r_data_o[769] = (N3)? mem[769] : 
                         (N0)? mem[2369] : 1'b0;
  assign r_data_o[768] = (N3)? mem[768] : 
                         (N0)? mem[2368] : 1'b0;
  assign r_data_o[767] = (N3)? mem[767] : 
                         (N0)? mem[2367] : 1'b0;
  assign r_data_o[766] = (N3)? mem[766] : 
                         (N0)? mem[2366] : 1'b0;
  assign r_data_o[765] = (N3)? mem[765] : 
                         (N0)? mem[2365] : 1'b0;
  assign r_data_o[764] = (N3)? mem[764] : 
                         (N0)? mem[2364] : 1'b0;
  assign r_data_o[763] = (N3)? mem[763] : 
                         (N0)? mem[2363] : 1'b0;
  assign r_data_o[762] = (N3)? mem[762] : 
                         (N0)? mem[2362] : 1'b0;
  assign r_data_o[761] = (N3)? mem[761] : 
                         (N0)? mem[2361] : 1'b0;
  assign r_data_o[760] = (N3)? mem[760] : 
                         (N0)? mem[2360] : 1'b0;
  assign r_data_o[759] = (N3)? mem[759] : 
                         (N0)? mem[2359] : 1'b0;
  assign r_data_o[758] = (N3)? mem[758] : 
                         (N0)? mem[2358] : 1'b0;
  assign r_data_o[757] = (N3)? mem[757] : 
                         (N0)? mem[2357] : 1'b0;
  assign r_data_o[756] = (N3)? mem[756] : 
                         (N0)? mem[2356] : 1'b0;
  assign r_data_o[755] = (N3)? mem[755] : 
                         (N0)? mem[2355] : 1'b0;
  assign r_data_o[754] = (N3)? mem[754] : 
                         (N0)? mem[2354] : 1'b0;
  assign r_data_o[753] = (N3)? mem[753] : 
                         (N0)? mem[2353] : 1'b0;
  assign r_data_o[752] = (N3)? mem[752] : 
                         (N0)? mem[2352] : 1'b0;
  assign r_data_o[751] = (N3)? mem[751] : 
                         (N0)? mem[2351] : 1'b0;
  assign r_data_o[750] = (N3)? mem[750] : 
                         (N0)? mem[2350] : 1'b0;
  assign r_data_o[749] = (N3)? mem[749] : 
                         (N0)? mem[2349] : 1'b0;
  assign r_data_o[748] = (N3)? mem[748] : 
                         (N0)? mem[2348] : 1'b0;
  assign r_data_o[747] = (N3)? mem[747] : 
                         (N0)? mem[2347] : 1'b0;
  assign r_data_o[746] = (N3)? mem[746] : 
                         (N0)? mem[2346] : 1'b0;
  assign r_data_o[745] = (N3)? mem[745] : 
                         (N0)? mem[2345] : 1'b0;
  assign r_data_o[744] = (N3)? mem[744] : 
                         (N0)? mem[2344] : 1'b0;
  assign r_data_o[743] = (N3)? mem[743] : 
                         (N0)? mem[2343] : 1'b0;
  assign r_data_o[742] = (N3)? mem[742] : 
                         (N0)? mem[2342] : 1'b0;
  assign r_data_o[741] = (N3)? mem[741] : 
                         (N0)? mem[2341] : 1'b0;
  assign r_data_o[740] = (N3)? mem[740] : 
                         (N0)? mem[2340] : 1'b0;
  assign r_data_o[739] = (N3)? mem[739] : 
                         (N0)? mem[2339] : 1'b0;
  assign r_data_o[738] = (N3)? mem[738] : 
                         (N0)? mem[2338] : 1'b0;
  assign r_data_o[737] = (N3)? mem[737] : 
                         (N0)? mem[2337] : 1'b0;
  assign r_data_o[736] = (N3)? mem[736] : 
                         (N0)? mem[2336] : 1'b0;
  assign r_data_o[735] = (N3)? mem[735] : 
                         (N0)? mem[2335] : 1'b0;
  assign r_data_o[734] = (N3)? mem[734] : 
                         (N0)? mem[2334] : 1'b0;
  assign r_data_o[733] = (N3)? mem[733] : 
                         (N0)? mem[2333] : 1'b0;
  assign r_data_o[732] = (N3)? mem[732] : 
                         (N0)? mem[2332] : 1'b0;
  assign r_data_o[731] = (N3)? mem[731] : 
                         (N0)? mem[2331] : 1'b0;
  assign r_data_o[730] = (N3)? mem[730] : 
                         (N0)? mem[2330] : 1'b0;
  assign r_data_o[729] = (N3)? mem[729] : 
                         (N0)? mem[2329] : 1'b0;
  assign r_data_o[728] = (N3)? mem[728] : 
                         (N0)? mem[2328] : 1'b0;
  assign r_data_o[727] = (N3)? mem[727] : 
                         (N0)? mem[2327] : 1'b0;
  assign r_data_o[726] = (N3)? mem[726] : 
                         (N0)? mem[2326] : 1'b0;
  assign r_data_o[725] = (N3)? mem[725] : 
                         (N0)? mem[2325] : 1'b0;
  assign r_data_o[724] = (N3)? mem[724] : 
                         (N0)? mem[2324] : 1'b0;
  assign r_data_o[723] = (N3)? mem[723] : 
                         (N0)? mem[2323] : 1'b0;
  assign r_data_o[722] = (N3)? mem[722] : 
                         (N0)? mem[2322] : 1'b0;
  assign r_data_o[721] = (N3)? mem[721] : 
                         (N0)? mem[2321] : 1'b0;
  assign r_data_o[720] = (N3)? mem[720] : 
                         (N0)? mem[2320] : 1'b0;
  assign r_data_o[719] = (N3)? mem[719] : 
                         (N0)? mem[2319] : 1'b0;
  assign r_data_o[718] = (N3)? mem[718] : 
                         (N0)? mem[2318] : 1'b0;
  assign r_data_o[717] = (N3)? mem[717] : 
                         (N0)? mem[2317] : 1'b0;
  assign r_data_o[716] = (N3)? mem[716] : 
                         (N0)? mem[2316] : 1'b0;
  assign r_data_o[715] = (N3)? mem[715] : 
                         (N0)? mem[2315] : 1'b0;
  assign r_data_o[714] = (N3)? mem[714] : 
                         (N0)? mem[2314] : 1'b0;
  assign r_data_o[713] = (N3)? mem[713] : 
                         (N0)? mem[2313] : 1'b0;
  assign r_data_o[712] = (N3)? mem[712] : 
                         (N0)? mem[2312] : 1'b0;
  assign r_data_o[711] = (N3)? mem[711] : 
                         (N0)? mem[2311] : 1'b0;
  assign r_data_o[710] = (N3)? mem[710] : 
                         (N0)? mem[2310] : 1'b0;
  assign r_data_o[709] = (N3)? mem[709] : 
                         (N0)? mem[2309] : 1'b0;
  assign r_data_o[708] = (N3)? mem[708] : 
                         (N0)? mem[2308] : 1'b0;
  assign r_data_o[707] = (N3)? mem[707] : 
                         (N0)? mem[2307] : 1'b0;
  assign r_data_o[706] = (N3)? mem[706] : 
                         (N0)? mem[2306] : 1'b0;
  assign r_data_o[705] = (N3)? mem[705] : 
                         (N0)? mem[2305] : 1'b0;
  assign r_data_o[704] = (N3)? mem[704] : 
                         (N0)? mem[2304] : 1'b0;
  assign r_data_o[703] = (N3)? mem[703] : 
                         (N0)? mem[2303] : 1'b0;
  assign r_data_o[702] = (N3)? mem[702] : 
                         (N0)? mem[2302] : 1'b0;
  assign r_data_o[701] = (N3)? mem[701] : 
                         (N0)? mem[2301] : 1'b0;
  assign r_data_o[700] = (N3)? mem[700] : 
                         (N0)? mem[2300] : 1'b0;
  assign r_data_o[699] = (N3)? mem[699] : 
                         (N0)? mem[2299] : 1'b0;
  assign r_data_o[698] = (N3)? mem[698] : 
                         (N0)? mem[2298] : 1'b0;
  assign r_data_o[697] = (N3)? mem[697] : 
                         (N0)? mem[2297] : 1'b0;
  assign r_data_o[696] = (N3)? mem[696] : 
                         (N0)? mem[2296] : 1'b0;
  assign r_data_o[695] = (N3)? mem[695] : 
                         (N0)? mem[2295] : 1'b0;
  assign r_data_o[694] = (N3)? mem[694] : 
                         (N0)? mem[2294] : 1'b0;
  assign r_data_o[693] = (N3)? mem[693] : 
                         (N0)? mem[2293] : 1'b0;
  assign r_data_o[692] = (N3)? mem[692] : 
                         (N0)? mem[2292] : 1'b0;
  assign r_data_o[691] = (N3)? mem[691] : 
                         (N0)? mem[2291] : 1'b0;
  assign r_data_o[690] = (N3)? mem[690] : 
                         (N0)? mem[2290] : 1'b0;
  assign r_data_o[689] = (N3)? mem[689] : 
                         (N0)? mem[2289] : 1'b0;
  assign r_data_o[688] = (N3)? mem[688] : 
                         (N0)? mem[2288] : 1'b0;
  assign r_data_o[687] = (N3)? mem[687] : 
                         (N0)? mem[2287] : 1'b0;
  assign r_data_o[686] = (N3)? mem[686] : 
                         (N0)? mem[2286] : 1'b0;
  assign r_data_o[685] = (N3)? mem[685] : 
                         (N0)? mem[2285] : 1'b0;
  assign r_data_o[684] = (N3)? mem[684] : 
                         (N0)? mem[2284] : 1'b0;
  assign r_data_o[683] = (N3)? mem[683] : 
                         (N0)? mem[2283] : 1'b0;
  assign r_data_o[682] = (N3)? mem[682] : 
                         (N0)? mem[2282] : 1'b0;
  assign r_data_o[681] = (N3)? mem[681] : 
                         (N0)? mem[2281] : 1'b0;
  assign r_data_o[680] = (N3)? mem[680] : 
                         (N0)? mem[2280] : 1'b0;
  assign r_data_o[679] = (N3)? mem[679] : 
                         (N0)? mem[2279] : 1'b0;
  assign r_data_o[678] = (N3)? mem[678] : 
                         (N0)? mem[2278] : 1'b0;
  assign r_data_o[677] = (N3)? mem[677] : 
                         (N0)? mem[2277] : 1'b0;
  assign r_data_o[676] = (N3)? mem[676] : 
                         (N0)? mem[2276] : 1'b0;
  assign r_data_o[675] = (N3)? mem[675] : 
                         (N0)? mem[2275] : 1'b0;
  assign r_data_o[674] = (N3)? mem[674] : 
                         (N0)? mem[2274] : 1'b0;
  assign r_data_o[673] = (N3)? mem[673] : 
                         (N0)? mem[2273] : 1'b0;
  assign r_data_o[672] = (N3)? mem[672] : 
                         (N0)? mem[2272] : 1'b0;
  assign r_data_o[671] = (N3)? mem[671] : 
                         (N0)? mem[2271] : 1'b0;
  assign r_data_o[670] = (N3)? mem[670] : 
                         (N0)? mem[2270] : 1'b0;
  assign r_data_o[669] = (N3)? mem[669] : 
                         (N0)? mem[2269] : 1'b0;
  assign r_data_o[668] = (N3)? mem[668] : 
                         (N0)? mem[2268] : 1'b0;
  assign r_data_o[667] = (N3)? mem[667] : 
                         (N0)? mem[2267] : 1'b0;
  assign r_data_o[666] = (N3)? mem[666] : 
                         (N0)? mem[2266] : 1'b0;
  assign r_data_o[665] = (N3)? mem[665] : 
                         (N0)? mem[2265] : 1'b0;
  assign r_data_o[664] = (N3)? mem[664] : 
                         (N0)? mem[2264] : 1'b0;
  assign r_data_o[663] = (N3)? mem[663] : 
                         (N0)? mem[2263] : 1'b0;
  assign r_data_o[662] = (N3)? mem[662] : 
                         (N0)? mem[2262] : 1'b0;
  assign r_data_o[661] = (N3)? mem[661] : 
                         (N0)? mem[2261] : 1'b0;
  assign r_data_o[660] = (N3)? mem[660] : 
                         (N0)? mem[2260] : 1'b0;
  assign r_data_o[659] = (N3)? mem[659] : 
                         (N0)? mem[2259] : 1'b0;
  assign r_data_o[658] = (N3)? mem[658] : 
                         (N0)? mem[2258] : 1'b0;
  assign r_data_o[657] = (N3)? mem[657] : 
                         (N0)? mem[2257] : 1'b0;
  assign r_data_o[656] = (N3)? mem[656] : 
                         (N0)? mem[2256] : 1'b0;
  assign r_data_o[655] = (N3)? mem[655] : 
                         (N0)? mem[2255] : 1'b0;
  assign r_data_o[654] = (N3)? mem[654] : 
                         (N0)? mem[2254] : 1'b0;
  assign r_data_o[653] = (N3)? mem[653] : 
                         (N0)? mem[2253] : 1'b0;
  assign r_data_o[652] = (N3)? mem[652] : 
                         (N0)? mem[2252] : 1'b0;
  assign r_data_o[651] = (N3)? mem[651] : 
                         (N0)? mem[2251] : 1'b0;
  assign r_data_o[650] = (N3)? mem[650] : 
                         (N0)? mem[2250] : 1'b0;
  assign r_data_o[649] = (N3)? mem[649] : 
                         (N0)? mem[2249] : 1'b0;
  assign r_data_o[648] = (N3)? mem[648] : 
                         (N0)? mem[2248] : 1'b0;
  assign r_data_o[647] = (N3)? mem[647] : 
                         (N0)? mem[2247] : 1'b0;
  assign r_data_o[646] = (N3)? mem[646] : 
                         (N0)? mem[2246] : 1'b0;
  assign r_data_o[645] = (N3)? mem[645] : 
                         (N0)? mem[2245] : 1'b0;
  assign r_data_o[644] = (N3)? mem[644] : 
                         (N0)? mem[2244] : 1'b0;
  assign r_data_o[643] = (N3)? mem[643] : 
                         (N0)? mem[2243] : 1'b0;
  assign r_data_o[642] = (N3)? mem[642] : 
                         (N0)? mem[2242] : 1'b0;
  assign r_data_o[641] = (N3)? mem[641] : 
                         (N0)? mem[2241] : 1'b0;
  assign r_data_o[640] = (N3)? mem[640] : 
                         (N0)? mem[2240] : 1'b0;
  assign r_data_o[639] = (N3)? mem[639] : 
                         (N0)? mem[2239] : 1'b0;
  assign r_data_o[638] = (N3)? mem[638] : 
                         (N0)? mem[2238] : 1'b0;
  assign r_data_o[637] = (N3)? mem[637] : 
                         (N0)? mem[2237] : 1'b0;
  assign r_data_o[636] = (N3)? mem[636] : 
                         (N0)? mem[2236] : 1'b0;
  assign r_data_o[635] = (N3)? mem[635] : 
                         (N0)? mem[2235] : 1'b0;
  assign r_data_o[634] = (N3)? mem[634] : 
                         (N0)? mem[2234] : 1'b0;
  assign r_data_o[633] = (N3)? mem[633] : 
                         (N0)? mem[2233] : 1'b0;
  assign r_data_o[632] = (N3)? mem[632] : 
                         (N0)? mem[2232] : 1'b0;
  assign r_data_o[631] = (N3)? mem[631] : 
                         (N0)? mem[2231] : 1'b0;
  assign r_data_o[630] = (N3)? mem[630] : 
                         (N0)? mem[2230] : 1'b0;
  assign r_data_o[629] = (N3)? mem[629] : 
                         (N0)? mem[2229] : 1'b0;
  assign r_data_o[628] = (N3)? mem[628] : 
                         (N0)? mem[2228] : 1'b0;
  assign r_data_o[627] = (N3)? mem[627] : 
                         (N0)? mem[2227] : 1'b0;
  assign r_data_o[626] = (N3)? mem[626] : 
                         (N0)? mem[2226] : 1'b0;
  assign r_data_o[625] = (N3)? mem[625] : 
                         (N0)? mem[2225] : 1'b0;
  assign r_data_o[624] = (N3)? mem[624] : 
                         (N0)? mem[2224] : 1'b0;
  assign r_data_o[623] = (N3)? mem[623] : 
                         (N0)? mem[2223] : 1'b0;
  assign r_data_o[622] = (N3)? mem[622] : 
                         (N0)? mem[2222] : 1'b0;
  assign r_data_o[621] = (N3)? mem[621] : 
                         (N0)? mem[2221] : 1'b0;
  assign r_data_o[620] = (N3)? mem[620] : 
                         (N0)? mem[2220] : 1'b0;
  assign r_data_o[619] = (N3)? mem[619] : 
                         (N0)? mem[2219] : 1'b0;
  assign r_data_o[618] = (N3)? mem[618] : 
                         (N0)? mem[2218] : 1'b0;
  assign r_data_o[617] = (N3)? mem[617] : 
                         (N0)? mem[2217] : 1'b0;
  assign r_data_o[616] = (N3)? mem[616] : 
                         (N0)? mem[2216] : 1'b0;
  assign r_data_o[615] = (N3)? mem[615] : 
                         (N0)? mem[2215] : 1'b0;
  assign r_data_o[614] = (N3)? mem[614] : 
                         (N0)? mem[2214] : 1'b0;
  assign r_data_o[613] = (N3)? mem[613] : 
                         (N0)? mem[2213] : 1'b0;
  assign r_data_o[612] = (N3)? mem[612] : 
                         (N0)? mem[2212] : 1'b0;
  assign r_data_o[611] = (N3)? mem[611] : 
                         (N0)? mem[2211] : 1'b0;
  assign r_data_o[610] = (N3)? mem[610] : 
                         (N0)? mem[2210] : 1'b0;
  assign r_data_o[609] = (N3)? mem[609] : 
                         (N0)? mem[2209] : 1'b0;
  assign r_data_o[608] = (N3)? mem[608] : 
                         (N0)? mem[2208] : 1'b0;
  assign r_data_o[607] = (N3)? mem[607] : 
                         (N0)? mem[2207] : 1'b0;
  assign r_data_o[606] = (N3)? mem[606] : 
                         (N0)? mem[2206] : 1'b0;
  assign r_data_o[605] = (N3)? mem[605] : 
                         (N0)? mem[2205] : 1'b0;
  assign r_data_o[604] = (N3)? mem[604] : 
                         (N0)? mem[2204] : 1'b0;
  assign r_data_o[603] = (N3)? mem[603] : 
                         (N0)? mem[2203] : 1'b0;
  assign r_data_o[602] = (N3)? mem[602] : 
                         (N0)? mem[2202] : 1'b0;
  assign r_data_o[601] = (N3)? mem[601] : 
                         (N0)? mem[2201] : 1'b0;
  assign r_data_o[600] = (N3)? mem[600] : 
                         (N0)? mem[2200] : 1'b0;
  assign r_data_o[599] = (N3)? mem[599] : 
                         (N0)? mem[2199] : 1'b0;
  assign r_data_o[598] = (N3)? mem[598] : 
                         (N0)? mem[2198] : 1'b0;
  assign r_data_o[597] = (N3)? mem[597] : 
                         (N0)? mem[2197] : 1'b0;
  assign r_data_o[596] = (N3)? mem[596] : 
                         (N0)? mem[2196] : 1'b0;
  assign r_data_o[595] = (N3)? mem[595] : 
                         (N0)? mem[2195] : 1'b0;
  assign r_data_o[594] = (N3)? mem[594] : 
                         (N0)? mem[2194] : 1'b0;
  assign r_data_o[593] = (N3)? mem[593] : 
                         (N0)? mem[2193] : 1'b0;
  assign r_data_o[592] = (N3)? mem[592] : 
                         (N0)? mem[2192] : 1'b0;
  assign r_data_o[591] = (N3)? mem[591] : 
                         (N0)? mem[2191] : 1'b0;
  assign r_data_o[590] = (N3)? mem[590] : 
                         (N0)? mem[2190] : 1'b0;
  assign r_data_o[589] = (N3)? mem[589] : 
                         (N0)? mem[2189] : 1'b0;
  assign r_data_o[588] = (N3)? mem[588] : 
                         (N0)? mem[2188] : 1'b0;
  assign r_data_o[587] = (N3)? mem[587] : 
                         (N0)? mem[2187] : 1'b0;
  assign r_data_o[586] = (N3)? mem[586] : 
                         (N0)? mem[2186] : 1'b0;
  assign r_data_o[585] = (N3)? mem[585] : 
                         (N0)? mem[2185] : 1'b0;
  assign r_data_o[584] = (N3)? mem[584] : 
                         (N0)? mem[2184] : 1'b0;
  assign r_data_o[583] = (N3)? mem[583] : 
                         (N0)? mem[2183] : 1'b0;
  assign r_data_o[582] = (N3)? mem[582] : 
                         (N0)? mem[2182] : 1'b0;
  assign r_data_o[581] = (N3)? mem[581] : 
                         (N0)? mem[2181] : 1'b0;
  assign r_data_o[580] = (N3)? mem[580] : 
                         (N0)? mem[2180] : 1'b0;
  assign r_data_o[579] = (N3)? mem[579] : 
                         (N0)? mem[2179] : 1'b0;
  assign r_data_o[578] = (N3)? mem[578] : 
                         (N0)? mem[2178] : 1'b0;
  assign r_data_o[577] = (N3)? mem[577] : 
                         (N0)? mem[2177] : 1'b0;
  assign r_data_o[576] = (N3)? mem[576] : 
                         (N0)? mem[2176] : 1'b0;
  assign r_data_o[575] = (N3)? mem[575] : 
                         (N0)? mem[2175] : 1'b0;
  assign r_data_o[574] = (N3)? mem[574] : 
                         (N0)? mem[2174] : 1'b0;
  assign r_data_o[573] = (N3)? mem[573] : 
                         (N0)? mem[2173] : 1'b0;
  assign r_data_o[572] = (N3)? mem[572] : 
                         (N0)? mem[2172] : 1'b0;
  assign r_data_o[571] = (N3)? mem[571] : 
                         (N0)? mem[2171] : 1'b0;
  assign r_data_o[570] = (N3)? mem[570] : 
                         (N0)? mem[2170] : 1'b0;
  assign r_data_o[569] = (N3)? mem[569] : 
                         (N0)? mem[2169] : 1'b0;
  assign r_data_o[568] = (N3)? mem[568] : 
                         (N0)? mem[2168] : 1'b0;
  assign r_data_o[567] = (N3)? mem[567] : 
                         (N0)? mem[2167] : 1'b0;
  assign r_data_o[566] = (N3)? mem[566] : 
                         (N0)? mem[2166] : 1'b0;
  assign r_data_o[565] = (N3)? mem[565] : 
                         (N0)? mem[2165] : 1'b0;
  assign r_data_o[564] = (N3)? mem[564] : 
                         (N0)? mem[2164] : 1'b0;
  assign r_data_o[563] = (N3)? mem[563] : 
                         (N0)? mem[2163] : 1'b0;
  assign r_data_o[562] = (N3)? mem[562] : 
                         (N0)? mem[2162] : 1'b0;
  assign r_data_o[561] = (N3)? mem[561] : 
                         (N0)? mem[2161] : 1'b0;
  assign r_data_o[560] = (N3)? mem[560] : 
                         (N0)? mem[2160] : 1'b0;
  assign r_data_o[559] = (N3)? mem[559] : 
                         (N0)? mem[2159] : 1'b0;
  assign r_data_o[558] = (N3)? mem[558] : 
                         (N0)? mem[2158] : 1'b0;
  assign r_data_o[557] = (N3)? mem[557] : 
                         (N0)? mem[2157] : 1'b0;
  assign r_data_o[556] = (N3)? mem[556] : 
                         (N0)? mem[2156] : 1'b0;
  assign r_data_o[555] = (N3)? mem[555] : 
                         (N0)? mem[2155] : 1'b0;
  assign r_data_o[554] = (N3)? mem[554] : 
                         (N0)? mem[2154] : 1'b0;
  assign r_data_o[553] = (N3)? mem[553] : 
                         (N0)? mem[2153] : 1'b0;
  assign r_data_o[552] = (N3)? mem[552] : 
                         (N0)? mem[2152] : 1'b0;
  assign r_data_o[551] = (N3)? mem[551] : 
                         (N0)? mem[2151] : 1'b0;
  assign r_data_o[550] = (N3)? mem[550] : 
                         (N0)? mem[2150] : 1'b0;
  assign r_data_o[549] = (N3)? mem[549] : 
                         (N0)? mem[2149] : 1'b0;
  assign r_data_o[548] = (N3)? mem[548] : 
                         (N0)? mem[2148] : 1'b0;
  assign r_data_o[547] = (N3)? mem[547] : 
                         (N0)? mem[2147] : 1'b0;
  assign r_data_o[546] = (N3)? mem[546] : 
                         (N0)? mem[2146] : 1'b0;
  assign r_data_o[545] = (N3)? mem[545] : 
                         (N0)? mem[2145] : 1'b0;
  assign r_data_o[544] = (N3)? mem[544] : 
                         (N0)? mem[2144] : 1'b0;
  assign r_data_o[543] = (N3)? mem[543] : 
                         (N0)? mem[2143] : 1'b0;
  assign r_data_o[542] = (N3)? mem[542] : 
                         (N0)? mem[2142] : 1'b0;
  assign r_data_o[541] = (N3)? mem[541] : 
                         (N0)? mem[2141] : 1'b0;
  assign r_data_o[540] = (N3)? mem[540] : 
                         (N0)? mem[2140] : 1'b0;
  assign r_data_o[539] = (N3)? mem[539] : 
                         (N0)? mem[2139] : 1'b0;
  assign r_data_o[538] = (N3)? mem[538] : 
                         (N0)? mem[2138] : 1'b0;
  assign r_data_o[537] = (N3)? mem[537] : 
                         (N0)? mem[2137] : 1'b0;
  assign r_data_o[536] = (N3)? mem[536] : 
                         (N0)? mem[2136] : 1'b0;
  assign r_data_o[535] = (N3)? mem[535] : 
                         (N0)? mem[2135] : 1'b0;
  assign r_data_o[534] = (N3)? mem[534] : 
                         (N0)? mem[2134] : 1'b0;
  assign r_data_o[533] = (N3)? mem[533] : 
                         (N0)? mem[2133] : 1'b0;
  assign r_data_o[532] = (N3)? mem[532] : 
                         (N0)? mem[2132] : 1'b0;
  assign r_data_o[531] = (N3)? mem[531] : 
                         (N0)? mem[2131] : 1'b0;
  assign r_data_o[530] = (N3)? mem[530] : 
                         (N0)? mem[2130] : 1'b0;
  assign r_data_o[529] = (N3)? mem[529] : 
                         (N0)? mem[2129] : 1'b0;
  assign r_data_o[528] = (N3)? mem[528] : 
                         (N0)? mem[2128] : 1'b0;
  assign r_data_o[527] = (N3)? mem[527] : 
                         (N0)? mem[2127] : 1'b0;
  assign r_data_o[526] = (N3)? mem[526] : 
                         (N0)? mem[2126] : 1'b0;
  assign r_data_o[525] = (N3)? mem[525] : 
                         (N0)? mem[2125] : 1'b0;
  assign r_data_o[524] = (N3)? mem[524] : 
                         (N0)? mem[2124] : 1'b0;
  assign r_data_o[523] = (N3)? mem[523] : 
                         (N0)? mem[2123] : 1'b0;
  assign r_data_o[522] = (N3)? mem[522] : 
                         (N0)? mem[2122] : 1'b0;
  assign r_data_o[521] = (N3)? mem[521] : 
                         (N0)? mem[2121] : 1'b0;
  assign r_data_o[520] = (N3)? mem[520] : 
                         (N0)? mem[2120] : 1'b0;
  assign r_data_o[519] = (N3)? mem[519] : 
                         (N0)? mem[2119] : 1'b0;
  assign r_data_o[518] = (N3)? mem[518] : 
                         (N0)? mem[2118] : 1'b0;
  assign r_data_o[517] = (N3)? mem[517] : 
                         (N0)? mem[2117] : 1'b0;
  assign r_data_o[516] = (N3)? mem[516] : 
                         (N0)? mem[2116] : 1'b0;
  assign r_data_o[515] = (N3)? mem[515] : 
                         (N0)? mem[2115] : 1'b0;
  assign r_data_o[514] = (N3)? mem[514] : 
                         (N0)? mem[2114] : 1'b0;
  assign r_data_o[513] = (N3)? mem[513] : 
                         (N0)? mem[2113] : 1'b0;
  assign r_data_o[512] = (N3)? mem[512] : 
                         (N0)? mem[2112] : 1'b0;
  assign r_data_o[511] = (N3)? mem[511] : 
                         (N0)? mem[2111] : 1'b0;
  assign r_data_o[510] = (N3)? mem[510] : 
                         (N0)? mem[2110] : 1'b0;
  assign r_data_o[509] = (N3)? mem[509] : 
                         (N0)? mem[2109] : 1'b0;
  assign r_data_o[508] = (N3)? mem[508] : 
                         (N0)? mem[2108] : 1'b0;
  assign r_data_o[507] = (N3)? mem[507] : 
                         (N0)? mem[2107] : 1'b0;
  assign r_data_o[506] = (N3)? mem[506] : 
                         (N0)? mem[2106] : 1'b0;
  assign r_data_o[505] = (N3)? mem[505] : 
                         (N0)? mem[2105] : 1'b0;
  assign r_data_o[504] = (N3)? mem[504] : 
                         (N0)? mem[2104] : 1'b0;
  assign r_data_o[503] = (N3)? mem[503] : 
                         (N0)? mem[2103] : 1'b0;
  assign r_data_o[502] = (N3)? mem[502] : 
                         (N0)? mem[2102] : 1'b0;
  assign r_data_o[501] = (N3)? mem[501] : 
                         (N0)? mem[2101] : 1'b0;
  assign r_data_o[500] = (N3)? mem[500] : 
                         (N0)? mem[2100] : 1'b0;
  assign r_data_o[499] = (N3)? mem[499] : 
                         (N0)? mem[2099] : 1'b0;
  assign r_data_o[498] = (N3)? mem[498] : 
                         (N0)? mem[2098] : 1'b0;
  assign r_data_o[497] = (N3)? mem[497] : 
                         (N0)? mem[2097] : 1'b0;
  assign r_data_o[496] = (N3)? mem[496] : 
                         (N0)? mem[2096] : 1'b0;
  assign r_data_o[495] = (N3)? mem[495] : 
                         (N0)? mem[2095] : 1'b0;
  assign r_data_o[494] = (N3)? mem[494] : 
                         (N0)? mem[2094] : 1'b0;
  assign r_data_o[493] = (N3)? mem[493] : 
                         (N0)? mem[2093] : 1'b0;
  assign r_data_o[492] = (N3)? mem[492] : 
                         (N0)? mem[2092] : 1'b0;
  assign r_data_o[491] = (N3)? mem[491] : 
                         (N0)? mem[2091] : 1'b0;
  assign r_data_o[490] = (N3)? mem[490] : 
                         (N0)? mem[2090] : 1'b0;
  assign r_data_o[489] = (N3)? mem[489] : 
                         (N0)? mem[2089] : 1'b0;
  assign r_data_o[488] = (N3)? mem[488] : 
                         (N0)? mem[2088] : 1'b0;
  assign r_data_o[487] = (N3)? mem[487] : 
                         (N0)? mem[2087] : 1'b0;
  assign r_data_o[486] = (N3)? mem[486] : 
                         (N0)? mem[2086] : 1'b0;
  assign r_data_o[485] = (N3)? mem[485] : 
                         (N0)? mem[2085] : 1'b0;
  assign r_data_o[484] = (N3)? mem[484] : 
                         (N0)? mem[2084] : 1'b0;
  assign r_data_o[483] = (N3)? mem[483] : 
                         (N0)? mem[2083] : 1'b0;
  assign r_data_o[482] = (N3)? mem[482] : 
                         (N0)? mem[2082] : 1'b0;
  assign r_data_o[481] = (N3)? mem[481] : 
                         (N0)? mem[2081] : 1'b0;
  assign r_data_o[480] = (N3)? mem[480] : 
                         (N0)? mem[2080] : 1'b0;
  assign r_data_o[479] = (N3)? mem[479] : 
                         (N0)? mem[2079] : 1'b0;
  assign r_data_o[478] = (N3)? mem[478] : 
                         (N0)? mem[2078] : 1'b0;
  assign r_data_o[477] = (N3)? mem[477] : 
                         (N0)? mem[2077] : 1'b0;
  assign r_data_o[476] = (N3)? mem[476] : 
                         (N0)? mem[2076] : 1'b0;
  assign r_data_o[475] = (N3)? mem[475] : 
                         (N0)? mem[2075] : 1'b0;
  assign r_data_o[474] = (N3)? mem[474] : 
                         (N0)? mem[2074] : 1'b0;
  assign r_data_o[473] = (N3)? mem[473] : 
                         (N0)? mem[2073] : 1'b0;
  assign r_data_o[472] = (N3)? mem[472] : 
                         (N0)? mem[2072] : 1'b0;
  assign r_data_o[471] = (N3)? mem[471] : 
                         (N0)? mem[2071] : 1'b0;
  assign r_data_o[470] = (N3)? mem[470] : 
                         (N0)? mem[2070] : 1'b0;
  assign r_data_o[469] = (N3)? mem[469] : 
                         (N0)? mem[2069] : 1'b0;
  assign r_data_o[468] = (N3)? mem[468] : 
                         (N0)? mem[2068] : 1'b0;
  assign r_data_o[467] = (N3)? mem[467] : 
                         (N0)? mem[2067] : 1'b0;
  assign r_data_o[466] = (N3)? mem[466] : 
                         (N0)? mem[2066] : 1'b0;
  assign r_data_o[465] = (N3)? mem[465] : 
                         (N0)? mem[2065] : 1'b0;
  assign r_data_o[464] = (N3)? mem[464] : 
                         (N0)? mem[2064] : 1'b0;
  assign r_data_o[463] = (N3)? mem[463] : 
                         (N0)? mem[2063] : 1'b0;
  assign r_data_o[462] = (N3)? mem[462] : 
                         (N0)? mem[2062] : 1'b0;
  assign r_data_o[461] = (N3)? mem[461] : 
                         (N0)? mem[2061] : 1'b0;
  assign r_data_o[460] = (N3)? mem[460] : 
                         (N0)? mem[2060] : 1'b0;
  assign r_data_o[459] = (N3)? mem[459] : 
                         (N0)? mem[2059] : 1'b0;
  assign r_data_o[458] = (N3)? mem[458] : 
                         (N0)? mem[2058] : 1'b0;
  assign r_data_o[457] = (N3)? mem[457] : 
                         (N0)? mem[2057] : 1'b0;
  assign r_data_o[456] = (N3)? mem[456] : 
                         (N0)? mem[2056] : 1'b0;
  assign r_data_o[455] = (N3)? mem[455] : 
                         (N0)? mem[2055] : 1'b0;
  assign r_data_o[454] = (N3)? mem[454] : 
                         (N0)? mem[2054] : 1'b0;
  assign r_data_o[453] = (N3)? mem[453] : 
                         (N0)? mem[2053] : 1'b0;
  assign r_data_o[452] = (N3)? mem[452] : 
                         (N0)? mem[2052] : 1'b0;
  assign r_data_o[451] = (N3)? mem[451] : 
                         (N0)? mem[2051] : 1'b0;
  assign r_data_o[450] = (N3)? mem[450] : 
                         (N0)? mem[2050] : 1'b0;
  assign r_data_o[449] = (N3)? mem[449] : 
                         (N0)? mem[2049] : 1'b0;
  assign r_data_o[448] = (N3)? mem[448] : 
                         (N0)? mem[2048] : 1'b0;
  assign r_data_o[447] = (N3)? mem[447] : 
                         (N0)? mem[2047] : 1'b0;
  assign r_data_o[446] = (N3)? mem[446] : 
                         (N0)? mem[2046] : 1'b0;
  assign r_data_o[445] = (N3)? mem[445] : 
                         (N0)? mem[2045] : 1'b0;
  assign r_data_o[444] = (N3)? mem[444] : 
                         (N0)? mem[2044] : 1'b0;
  assign r_data_o[443] = (N3)? mem[443] : 
                         (N0)? mem[2043] : 1'b0;
  assign r_data_o[442] = (N3)? mem[442] : 
                         (N0)? mem[2042] : 1'b0;
  assign r_data_o[441] = (N3)? mem[441] : 
                         (N0)? mem[2041] : 1'b0;
  assign r_data_o[440] = (N3)? mem[440] : 
                         (N0)? mem[2040] : 1'b0;
  assign r_data_o[439] = (N3)? mem[439] : 
                         (N0)? mem[2039] : 1'b0;
  assign r_data_o[438] = (N3)? mem[438] : 
                         (N0)? mem[2038] : 1'b0;
  assign r_data_o[437] = (N3)? mem[437] : 
                         (N0)? mem[2037] : 1'b0;
  assign r_data_o[436] = (N3)? mem[436] : 
                         (N0)? mem[2036] : 1'b0;
  assign r_data_o[435] = (N3)? mem[435] : 
                         (N0)? mem[2035] : 1'b0;
  assign r_data_o[434] = (N3)? mem[434] : 
                         (N0)? mem[2034] : 1'b0;
  assign r_data_o[433] = (N3)? mem[433] : 
                         (N0)? mem[2033] : 1'b0;
  assign r_data_o[432] = (N3)? mem[432] : 
                         (N0)? mem[2032] : 1'b0;
  assign r_data_o[431] = (N3)? mem[431] : 
                         (N0)? mem[2031] : 1'b0;
  assign r_data_o[430] = (N3)? mem[430] : 
                         (N0)? mem[2030] : 1'b0;
  assign r_data_o[429] = (N3)? mem[429] : 
                         (N0)? mem[2029] : 1'b0;
  assign r_data_o[428] = (N3)? mem[428] : 
                         (N0)? mem[2028] : 1'b0;
  assign r_data_o[427] = (N3)? mem[427] : 
                         (N0)? mem[2027] : 1'b0;
  assign r_data_o[426] = (N3)? mem[426] : 
                         (N0)? mem[2026] : 1'b0;
  assign r_data_o[425] = (N3)? mem[425] : 
                         (N0)? mem[2025] : 1'b0;
  assign r_data_o[424] = (N3)? mem[424] : 
                         (N0)? mem[2024] : 1'b0;
  assign r_data_o[423] = (N3)? mem[423] : 
                         (N0)? mem[2023] : 1'b0;
  assign r_data_o[422] = (N3)? mem[422] : 
                         (N0)? mem[2022] : 1'b0;
  assign r_data_o[421] = (N3)? mem[421] : 
                         (N0)? mem[2021] : 1'b0;
  assign r_data_o[420] = (N3)? mem[420] : 
                         (N0)? mem[2020] : 1'b0;
  assign r_data_o[419] = (N3)? mem[419] : 
                         (N0)? mem[2019] : 1'b0;
  assign r_data_o[418] = (N3)? mem[418] : 
                         (N0)? mem[2018] : 1'b0;
  assign r_data_o[417] = (N3)? mem[417] : 
                         (N0)? mem[2017] : 1'b0;
  assign r_data_o[416] = (N3)? mem[416] : 
                         (N0)? mem[2016] : 1'b0;
  assign r_data_o[415] = (N3)? mem[415] : 
                         (N0)? mem[2015] : 1'b0;
  assign r_data_o[414] = (N3)? mem[414] : 
                         (N0)? mem[2014] : 1'b0;
  assign r_data_o[413] = (N3)? mem[413] : 
                         (N0)? mem[2013] : 1'b0;
  assign r_data_o[412] = (N3)? mem[412] : 
                         (N0)? mem[2012] : 1'b0;
  assign r_data_o[411] = (N3)? mem[411] : 
                         (N0)? mem[2011] : 1'b0;
  assign r_data_o[410] = (N3)? mem[410] : 
                         (N0)? mem[2010] : 1'b0;
  assign r_data_o[409] = (N3)? mem[409] : 
                         (N0)? mem[2009] : 1'b0;
  assign r_data_o[408] = (N3)? mem[408] : 
                         (N0)? mem[2008] : 1'b0;
  assign r_data_o[407] = (N3)? mem[407] : 
                         (N0)? mem[2007] : 1'b0;
  assign r_data_o[406] = (N3)? mem[406] : 
                         (N0)? mem[2006] : 1'b0;
  assign r_data_o[405] = (N3)? mem[405] : 
                         (N0)? mem[2005] : 1'b0;
  assign r_data_o[404] = (N3)? mem[404] : 
                         (N0)? mem[2004] : 1'b0;
  assign r_data_o[403] = (N3)? mem[403] : 
                         (N0)? mem[2003] : 1'b0;
  assign r_data_o[402] = (N3)? mem[402] : 
                         (N0)? mem[2002] : 1'b0;
  assign r_data_o[401] = (N3)? mem[401] : 
                         (N0)? mem[2001] : 1'b0;
  assign r_data_o[400] = (N3)? mem[400] : 
                         (N0)? mem[2000] : 1'b0;
  assign r_data_o[399] = (N3)? mem[399] : 
                         (N0)? mem[1999] : 1'b0;
  assign r_data_o[398] = (N3)? mem[398] : 
                         (N0)? mem[1998] : 1'b0;
  assign r_data_o[397] = (N3)? mem[397] : 
                         (N0)? mem[1997] : 1'b0;
  assign r_data_o[396] = (N3)? mem[396] : 
                         (N0)? mem[1996] : 1'b0;
  assign r_data_o[395] = (N3)? mem[395] : 
                         (N0)? mem[1995] : 1'b0;
  assign r_data_o[394] = (N3)? mem[394] : 
                         (N0)? mem[1994] : 1'b0;
  assign r_data_o[393] = (N3)? mem[393] : 
                         (N0)? mem[1993] : 1'b0;
  assign r_data_o[392] = (N3)? mem[392] : 
                         (N0)? mem[1992] : 1'b0;
  assign r_data_o[391] = (N3)? mem[391] : 
                         (N0)? mem[1991] : 1'b0;
  assign r_data_o[390] = (N3)? mem[390] : 
                         (N0)? mem[1990] : 1'b0;
  assign r_data_o[389] = (N3)? mem[389] : 
                         (N0)? mem[1989] : 1'b0;
  assign r_data_o[388] = (N3)? mem[388] : 
                         (N0)? mem[1988] : 1'b0;
  assign r_data_o[387] = (N3)? mem[387] : 
                         (N0)? mem[1987] : 1'b0;
  assign r_data_o[386] = (N3)? mem[386] : 
                         (N0)? mem[1986] : 1'b0;
  assign r_data_o[385] = (N3)? mem[385] : 
                         (N0)? mem[1985] : 1'b0;
  assign r_data_o[384] = (N3)? mem[384] : 
                         (N0)? mem[1984] : 1'b0;
  assign r_data_o[383] = (N3)? mem[383] : 
                         (N0)? mem[1983] : 1'b0;
  assign r_data_o[382] = (N3)? mem[382] : 
                         (N0)? mem[1982] : 1'b0;
  assign r_data_o[381] = (N3)? mem[381] : 
                         (N0)? mem[1981] : 1'b0;
  assign r_data_o[380] = (N3)? mem[380] : 
                         (N0)? mem[1980] : 1'b0;
  assign r_data_o[379] = (N3)? mem[379] : 
                         (N0)? mem[1979] : 1'b0;
  assign r_data_o[378] = (N3)? mem[378] : 
                         (N0)? mem[1978] : 1'b0;
  assign r_data_o[377] = (N3)? mem[377] : 
                         (N0)? mem[1977] : 1'b0;
  assign r_data_o[376] = (N3)? mem[376] : 
                         (N0)? mem[1976] : 1'b0;
  assign r_data_o[375] = (N3)? mem[375] : 
                         (N0)? mem[1975] : 1'b0;
  assign r_data_o[374] = (N3)? mem[374] : 
                         (N0)? mem[1974] : 1'b0;
  assign r_data_o[373] = (N3)? mem[373] : 
                         (N0)? mem[1973] : 1'b0;
  assign r_data_o[372] = (N3)? mem[372] : 
                         (N0)? mem[1972] : 1'b0;
  assign r_data_o[371] = (N3)? mem[371] : 
                         (N0)? mem[1971] : 1'b0;
  assign r_data_o[370] = (N3)? mem[370] : 
                         (N0)? mem[1970] : 1'b0;
  assign r_data_o[369] = (N3)? mem[369] : 
                         (N0)? mem[1969] : 1'b0;
  assign r_data_o[368] = (N3)? mem[368] : 
                         (N0)? mem[1968] : 1'b0;
  assign r_data_o[367] = (N3)? mem[367] : 
                         (N0)? mem[1967] : 1'b0;
  assign r_data_o[366] = (N3)? mem[366] : 
                         (N0)? mem[1966] : 1'b0;
  assign r_data_o[365] = (N3)? mem[365] : 
                         (N0)? mem[1965] : 1'b0;
  assign r_data_o[364] = (N3)? mem[364] : 
                         (N0)? mem[1964] : 1'b0;
  assign r_data_o[363] = (N3)? mem[363] : 
                         (N0)? mem[1963] : 1'b0;
  assign r_data_o[362] = (N3)? mem[362] : 
                         (N0)? mem[1962] : 1'b0;
  assign r_data_o[361] = (N3)? mem[361] : 
                         (N0)? mem[1961] : 1'b0;
  assign r_data_o[360] = (N3)? mem[360] : 
                         (N0)? mem[1960] : 1'b0;
  assign r_data_o[359] = (N3)? mem[359] : 
                         (N0)? mem[1959] : 1'b0;
  assign r_data_o[358] = (N3)? mem[358] : 
                         (N0)? mem[1958] : 1'b0;
  assign r_data_o[357] = (N3)? mem[357] : 
                         (N0)? mem[1957] : 1'b0;
  assign r_data_o[356] = (N3)? mem[356] : 
                         (N0)? mem[1956] : 1'b0;
  assign r_data_o[355] = (N3)? mem[355] : 
                         (N0)? mem[1955] : 1'b0;
  assign r_data_o[354] = (N3)? mem[354] : 
                         (N0)? mem[1954] : 1'b0;
  assign r_data_o[353] = (N3)? mem[353] : 
                         (N0)? mem[1953] : 1'b0;
  assign r_data_o[352] = (N3)? mem[352] : 
                         (N0)? mem[1952] : 1'b0;
  assign r_data_o[351] = (N3)? mem[351] : 
                         (N0)? mem[1951] : 1'b0;
  assign r_data_o[350] = (N3)? mem[350] : 
                         (N0)? mem[1950] : 1'b0;
  assign r_data_o[349] = (N3)? mem[349] : 
                         (N0)? mem[1949] : 1'b0;
  assign r_data_o[348] = (N3)? mem[348] : 
                         (N0)? mem[1948] : 1'b0;
  assign r_data_o[347] = (N3)? mem[347] : 
                         (N0)? mem[1947] : 1'b0;
  assign r_data_o[346] = (N3)? mem[346] : 
                         (N0)? mem[1946] : 1'b0;
  assign r_data_o[345] = (N3)? mem[345] : 
                         (N0)? mem[1945] : 1'b0;
  assign r_data_o[344] = (N3)? mem[344] : 
                         (N0)? mem[1944] : 1'b0;
  assign r_data_o[343] = (N3)? mem[343] : 
                         (N0)? mem[1943] : 1'b0;
  assign r_data_o[342] = (N3)? mem[342] : 
                         (N0)? mem[1942] : 1'b0;
  assign r_data_o[341] = (N3)? mem[341] : 
                         (N0)? mem[1941] : 1'b0;
  assign r_data_o[340] = (N3)? mem[340] : 
                         (N0)? mem[1940] : 1'b0;
  assign r_data_o[339] = (N3)? mem[339] : 
                         (N0)? mem[1939] : 1'b0;
  assign r_data_o[338] = (N3)? mem[338] : 
                         (N0)? mem[1938] : 1'b0;
  assign r_data_o[337] = (N3)? mem[337] : 
                         (N0)? mem[1937] : 1'b0;
  assign r_data_o[336] = (N3)? mem[336] : 
                         (N0)? mem[1936] : 1'b0;
  assign r_data_o[335] = (N3)? mem[335] : 
                         (N0)? mem[1935] : 1'b0;
  assign r_data_o[334] = (N3)? mem[334] : 
                         (N0)? mem[1934] : 1'b0;
  assign r_data_o[333] = (N3)? mem[333] : 
                         (N0)? mem[1933] : 1'b0;
  assign r_data_o[332] = (N3)? mem[332] : 
                         (N0)? mem[1932] : 1'b0;
  assign r_data_o[331] = (N3)? mem[331] : 
                         (N0)? mem[1931] : 1'b0;
  assign r_data_o[330] = (N3)? mem[330] : 
                         (N0)? mem[1930] : 1'b0;
  assign r_data_o[329] = (N3)? mem[329] : 
                         (N0)? mem[1929] : 1'b0;
  assign r_data_o[328] = (N3)? mem[328] : 
                         (N0)? mem[1928] : 1'b0;
  assign r_data_o[327] = (N3)? mem[327] : 
                         (N0)? mem[1927] : 1'b0;
  assign r_data_o[326] = (N3)? mem[326] : 
                         (N0)? mem[1926] : 1'b0;
  assign r_data_o[325] = (N3)? mem[325] : 
                         (N0)? mem[1925] : 1'b0;
  assign r_data_o[324] = (N3)? mem[324] : 
                         (N0)? mem[1924] : 1'b0;
  assign r_data_o[323] = (N3)? mem[323] : 
                         (N0)? mem[1923] : 1'b0;
  assign r_data_o[322] = (N3)? mem[322] : 
                         (N0)? mem[1922] : 1'b0;
  assign r_data_o[321] = (N3)? mem[321] : 
                         (N0)? mem[1921] : 1'b0;
  assign r_data_o[320] = (N3)? mem[320] : 
                         (N0)? mem[1920] : 1'b0;
  assign r_data_o[319] = (N3)? mem[319] : 
                         (N0)? mem[1919] : 1'b0;
  assign r_data_o[318] = (N3)? mem[318] : 
                         (N0)? mem[1918] : 1'b0;
  assign r_data_o[317] = (N3)? mem[317] : 
                         (N0)? mem[1917] : 1'b0;
  assign r_data_o[316] = (N3)? mem[316] : 
                         (N0)? mem[1916] : 1'b0;
  assign r_data_o[315] = (N3)? mem[315] : 
                         (N0)? mem[1915] : 1'b0;
  assign r_data_o[314] = (N3)? mem[314] : 
                         (N0)? mem[1914] : 1'b0;
  assign r_data_o[313] = (N3)? mem[313] : 
                         (N0)? mem[1913] : 1'b0;
  assign r_data_o[312] = (N3)? mem[312] : 
                         (N0)? mem[1912] : 1'b0;
  assign r_data_o[311] = (N3)? mem[311] : 
                         (N0)? mem[1911] : 1'b0;
  assign r_data_o[310] = (N3)? mem[310] : 
                         (N0)? mem[1910] : 1'b0;
  assign r_data_o[309] = (N3)? mem[309] : 
                         (N0)? mem[1909] : 1'b0;
  assign r_data_o[308] = (N3)? mem[308] : 
                         (N0)? mem[1908] : 1'b0;
  assign r_data_o[307] = (N3)? mem[307] : 
                         (N0)? mem[1907] : 1'b0;
  assign r_data_o[306] = (N3)? mem[306] : 
                         (N0)? mem[1906] : 1'b0;
  assign r_data_o[305] = (N3)? mem[305] : 
                         (N0)? mem[1905] : 1'b0;
  assign r_data_o[304] = (N3)? mem[304] : 
                         (N0)? mem[1904] : 1'b0;
  assign r_data_o[303] = (N3)? mem[303] : 
                         (N0)? mem[1903] : 1'b0;
  assign r_data_o[302] = (N3)? mem[302] : 
                         (N0)? mem[1902] : 1'b0;
  assign r_data_o[301] = (N3)? mem[301] : 
                         (N0)? mem[1901] : 1'b0;
  assign r_data_o[300] = (N3)? mem[300] : 
                         (N0)? mem[1900] : 1'b0;
  assign r_data_o[299] = (N3)? mem[299] : 
                         (N0)? mem[1899] : 1'b0;
  assign r_data_o[298] = (N3)? mem[298] : 
                         (N0)? mem[1898] : 1'b0;
  assign r_data_o[297] = (N3)? mem[297] : 
                         (N0)? mem[1897] : 1'b0;
  assign r_data_o[296] = (N3)? mem[296] : 
                         (N0)? mem[1896] : 1'b0;
  assign r_data_o[295] = (N3)? mem[295] : 
                         (N0)? mem[1895] : 1'b0;
  assign r_data_o[294] = (N3)? mem[294] : 
                         (N0)? mem[1894] : 1'b0;
  assign r_data_o[293] = (N3)? mem[293] : 
                         (N0)? mem[1893] : 1'b0;
  assign r_data_o[292] = (N3)? mem[292] : 
                         (N0)? mem[1892] : 1'b0;
  assign r_data_o[291] = (N3)? mem[291] : 
                         (N0)? mem[1891] : 1'b0;
  assign r_data_o[290] = (N3)? mem[290] : 
                         (N0)? mem[1890] : 1'b0;
  assign r_data_o[289] = (N3)? mem[289] : 
                         (N0)? mem[1889] : 1'b0;
  assign r_data_o[288] = (N3)? mem[288] : 
                         (N0)? mem[1888] : 1'b0;
  assign r_data_o[287] = (N3)? mem[287] : 
                         (N0)? mem[1887] : 1'b0;
  assign r_data_o[286] = (N3)? mem[286] : 
                         (N0)? mem[1886] : 1'b0;
  assign r_data_o[285] = (N3)? mem[285] : 
                         (N0)? mem[1885] : 1'b0;
  assign r_data_o[284] = (N3)? mem[284] : 
                         (N0)? mem[1884] : 1'b0;
  assign r_data_o[283] = (N3)? mem[283] : 
                         (N0)? mem[1883] : 1'b0;
  assign r_data_o[282] = (N3)? mem[282] : 
                         (N0)? mem[1882] : 1'b0;
  assign r_data_o[281] = (N3)? mem[281] : 
                         (N0)? mem[1881] : 1'b0;
  assign r_data_o[280] = (N3)? mem[280] : 
                         (N0)? mem[1880] : 1'b0;
  assign r_data_o[279] = (N3)? mem[279] : 
                         (N0)? mem[1879] : 1'b0;
  assign r_data_o[278] = (N3)? mem[278] : 
                         (N0)? mem[1878] : 1'b0;
  assign r_data_o[277] = (N3)? mem[277] : 
                         (N0)? mem[1877] : 1'b0;
  assign r_data_o[276] = (N3)? mem[276] : 
                         (N0)? mem[1876] : 1'b0;
  assign r_data_o[275] = (N3)? mem[275] : 
                         (N0)? mem[1875] : 1'b0;
  assign r_data_o[274] = (N3)? mem[274] : 
                         (N0)? mem[1874] : 1'b0;
  assign r_data_o[273] = (N3)? mem[273] : 
                         (N0)? mem[1873] : 1'b0;
  assign r_data_o[272] = (N3)? mem[272] : 
                         (N0)? mem[1872] : 1'b0;
  assign r_data_o[271] = (N3)? mem[271] : 
                         (N0)? mem[1871] : 1'b0;
  assign r_data_o[270] = (N3)? mem[270] : 
                         (N0)? mem[1870] : 1'b0;
  assign r_data_o[269] = (N3)? mem[269] : 
                         (N0)? mem[1869] : 1'b0;
  assign r_data_o[268] = (N3)? mem[268] : 
                         (N0)? mem[1868] : 1'b0;
  assign r_data_o[267] = (N3)? mem[267] : 
                         (N0)? mem[1867] : 1'b0;
  assign r_data_o[266] = (N3)? mem[266] : 
                         (N0)? mem[1866] : 1'b0;
  assign r_data_o[265] = (N3)? mem[265] : 
                         (N0)? mem[1865] : 1'b0;
  assign r_data_o[264] = (N3)? mem[264] : 
                         (N0)? mem[1864] : 1'b0;
  assign r_data_o[263] = (N3)? mem[263] : 
                         (N0)? mem[1863] : 1'b0;
  assign r_data_o[262] = (N3)? mem[262] : 
                         (N0)? mem[1862] : 1'b0;
  assign r_data_o[261] = (N3)? mem[261] : 
                         (N0)? mem[1861] : 1'b0;
  assign r_data_o[260] = (N3)? mem[260] : 
                         (N0)? mem[1860] : 1'b0;
  assign r_data_o[259] = (N3)? mem[259] : 
                         (N0)? mem[1859] : 1'b0;
  assign r_data_o[258] = (N3)? mem[258] : 
                         (N0)? mem[1858] : 1'b0;
  assign r_data_o[257] = (N3)? mem[257] : 
                         (N0)? mem[1857] : 1'b0;
  assign r_data_o[256] = (N3)? mem[256] : 
                         (N0)? mem[1856] : 1'b0;
  assign r_data_o[255] = (N3)? mem[255] : 
                         (N0)? mem[1855] : 1'b0;
  assign r_data_o[254] = (N3)? mem[254] : 
                         (N0)? mem[1854] : 1'b0;
  assign r_data_o[253] = (N3)? mem[253] : 
                         (N0)? mem[1853] : 1'b0;
  assign r_data_o[252] = (N3)? mem[252] : 
                         (N0)? mem[1852] : 1'b0;
  assign r_data_o[251] = (N3)? mem[251] : 
                         (N0)? mem[1851] : 1'b0;
  assign r_data_o[250] = (N3)? mem[250] : 
                         (N0)? mem[1850] : 1'b0;
  assign r_data_o[249] = (N3)? mem[249] : 
                         (N0)? mem[1849] : 1'b0;
  assign r_data_o[248] = (N3)? mem[248] : 
                         (N0)? mem[1848] : 1'b0;
  assign r_data_o[247] = (N3)? mem[247] : 
                         (N0)? mem[1847] : 1'b0;
  assign r_data_o[246] = (N3)? mem[246] : 
                         (N0)? mem[1846] : 1'b0;
  assign r_data_o[245] = (N3)? mem[245] : 
                         (N0)? mem[1845] : 1'b0;
  assign r_data_o[244] = (N3)? mem[244] : 
                         (N0)? mem[1844] : 1'b0;
  assign r_data_o[243] = (N3)? mem[243] : 
                         (N0)? mem[1843] : 1'b0;
  assign r_data_o[242] = (N3)? mem[242] : 
                         (N0)? mem[1842] : 1'b0;
  assign r_data_o[241] = (N3)? mem[241] : 
                         (N0)? mem[1841] : 1'b0;
  assign r_data_o[240] = (N3)? mem[240] : 
                         (N0)? mem[1840] : 1'b0;
  assign r_data_o[239] = (N3)? mem[239] : 
                         (N0)? mem[1839] : 1'b0;
  assign r_data_o[238] = (N3)? mem[238] : 
                         (N0)? mem[1838] : 1'b0;
  assign r_data_o[237] = (N3)? mem[237] : 
                         (N0)? mem[1837] : 1'b0;
  assign r_data_o[236] = (N3)? mem[236] : 
                         (N0)? mem[1836] : 1'b0;
  assign r_data_o[235] = (N3)? mem[235] : 
                         (N0)? mem[1835] : 1'b0;
  assign r_data_o[234] = (N3)? mem[234] : 
                         (N0)? mem[1834] : 1'b0;
  assign r_data_o[233] = (N3)? mem[233] : 
                         (N0)? mem[1833] : 1'b0;
  assign r_data_o[232] = (N3)? mem[232] : 
                         (N0)? mem[1832] : 1'b0;
  assign r_data_o[231] = (N3)? mem[231] : 
                         (N0)? mem[1831] : 1'b0;
  assign r_data_o[230] = (N3)? mem[230] : 
                         (N0)? mem[1830] : 1'b0;
  assign r_data_o[229] = (N3)? mem[229] : 
                         (N0)? mem[1829] : 1'b0;
  assign r_data_o[228] = (N3)? mem[228] : 
                         (N0)? mem[1828] : 1'b0;
  assign r_data_o[227] = (N3)? mem[227] : 
                         (N0)? mem[1827] : 1'b0;
  assign r_data_o[226] = (N3)? mem[226] : 
                         (N0)? mem[1826] : 1'b0;
  assign r_data_o[225] = (N3)? mem[225] : 
                         (N0)? mem[1825] : 1'b0;
  assign r_data_o[224] = (N3)? mem[224] : 
                         (N0)? mem[1824] : 1'b0;
  assign r_data_o[223] = (N3)? mem[223] : 
                         (N0)? mem[1823] : 1'b0;
  assign r_data_o[222] = (N3)? mem[222] : 
                         (N0)? mem[1822] : 1'b0;
  assign r_data_o[221] = (N3)? mem[221] : 
                         (N0)? mem[1821] : 1'b0;
  assign r_data_o[220] = (N3)? mem[220] : 
                         (N0)? mem[1820] : 1'b0;
  assign r_data_o[219] = (N3)? mem[219] : 
                         (N0)? mem[1819] : 1'b0;
  assign r_data_o[218] = (N3)? mem[218] : 
                         (N0)? mem[1818] : 1'b0;
  assign r_data_o[217] = (N3)? mem[217] : 
                         (N0)? mem[1817] : 1'b0;
  assign r_data_o[216] = (N3)? mem[216] : 
                         (N0)? mem[1816] : 1'b0;
  assign r_data_o[215] = (N3)? mem[215] : 
                         (N0)? mem[1815] : 1'b0;
  assign r_data_o[214] = (N3)? mem[214] : 
                         (N0)? mem[1814] : 1'b0;
  assign r_data_o[213] = (N3)? mem[213] : 
                         (N0)? mem[1813] : 1'b0;
  assign r_data_o[212] = (N3)? mem[212] : 
                         (N0)? mem[1812] : 1'b0;
  assign r_data_o[211] = (N3)? mem[211] : 
                         (N0)? mem[1811] : 1'b0;
  assign r_data_o[210] = (N3)? mem[210] : 
                         (N0)? mem[1810] : 1'b0;
  assign r_data_o[209] = (N3)? mem[209] : 
                         (N0)? mem[1809] : 1'b0;
  assign r_data_o[208] = (N3)? mem[208] : 
                         (N0)? mem[1808] : 1'b0;
  assign r_data_o[207] = (N3)? mem[207] : 
                         (N0)? mem[1807] : 1'b0;
  assign r_data_o[206] = (N3)? mem[206] : 
                         (N0)? mem[1806] : 1'b0;
  assign r_data_o[205] = (N3)? mem[205] : 
                         (N0)? mem[1805] : 1'b0;
  assign r_data_o[204] = (N3)? mem[204] : 
                         (N0)? mem[1804] : 1'b0;
  assign r_data_o[203] = (N3)? mem[203] : 
                         (N0)? mem[1803] : 1'b0;
  assign r_data_o[202] = (N3)? mem[202] : 
                         (N0)? mem[1802] : 1'b0;
  assign r_data_o[201] = (N3)? mem[201] : 
                         (N0)? mem[1801] : 1'b0;
  assign r_data_o[200] = (N3)? mem[200] : 
                         (N0)? mem[1800] : 1'b0;
  assign r_data_o[199] = (N3)? mem[199] : 
                         (N0)? mem[1799] : 1'b0;
  assign r_data_o[198] = (N3)? mem[198] : 
                         (N0)? mem[1798] : 1'b0;
  assign r_data_o[197] = (N3)? mem[197] : 
                         (N0)? mem[1797] : 1'b0;
  assign r_data_o[196] = (N3)? mem[196] : 
                         (N0)? mem[1796] : 1'b0;
  assign r_data_o[195] = (N3)? mem[195] : 
                         (N0)? mem[1795] : 1'b0;
  assign r_data_o[194] = (N3)? mem[194] : 
                         (N0)? mem[1794] : 1'b0;
  assign r_data_o[193] = (N3)? mem[193] : 
                         (N0)? mem[1793] : 1'b0;
  assign r_data_o[192] = (N3)? mem[192] : 
                         (N0)? mem[1792] : 1'b0;
  assign r_data_o[191] = (N3)? mem[191] : 
                         (N0)? mem[1791] : 1'b0;
  assign r_data_o[190] = (N3)? mem[190] : 
                         (N0)? mem[1790] : 1'b0;
  assign r_data_o[189] = (N3)? mem[189] : 
                         (N0)? mem[1789] : 1'b0;
  assign r_data_o[188] = (N3)? mem[188] : 
                         (N0)? mem[1788] : 1'b0;
  assign r_data_o[187] = (N3)? mem[187] : 
                         (N0)? mem[1787] : 1'b0;
  assign r_data_o[186] = (N3)? mem[186] : 
                         (N0)? mem[1786] : 1'b0;
  assign r_data_o[185] = (N3)? mem[185] : 
                         (N0)? mem[1785] : 1'b0;
  assign r_data_o[184] = (N3)? mem[184] : 
                         (N0)? mem[1784] : 1'b0;
  assign r_data_o[183] = (N3)? mem[183] : 
                         (N0)? mem[1783] : 1'b0;
  assign r_data_o[182] = (N3)? mem[182] : 
                         (N0)? mem[1782] : 1'b0;
  assign r_data_o[181] = (N3)? mem[181] : 
                         (N0)? mem[1781] : 1'b0;
  assign r_data_o[180] = (N3)? mem[180] : 
                         (N0)? mem[1780] : 1'b0;
  assign r_data_o[179] = (N3)? mem[179] : 
                         (N0)? mem[1779] : 1'b0;
  assign r_data_o[178] = (N3)? mem[178] : 
                         (N0)? mem[1778] : 1'b0;
  assign r_data_o[177] = (N3)? mem[177] : 
                         (N0)? mem[1777] : 1'b0;
  assign r_data_o[176] = (N3)? mem[176] : 
                         (N0)? mem[1776] : 1'b0;
  assign r_data_o[175] = (N3)? mem[175] : 
                         (N0)? mem[1775] : 1'b0;
  assign r_data_o[174] = (N3)? mem[174] : 
                         (N0)? mem[1774] : 1'b0;
  assign r_data_o[173] = (N3)? mem[173] : 
                         (N0)? mem[1773] : 1'b0;
  assign r_data_o[172] = (N3)? mem[172] : 
                         (N0)? mem[1772] : 1'b0;
  assign r_data_o[171] = (N3)? mem[171] : 
                         (N0)? mem[1771] : 1'b0;
  assign r_data_o[170] = (N3)? mem[170] : 
                         (N0)? mem[1770] : 1'b0;
  assign r_data_o[169] = (N3)? mem[169] : 
                         (N0)? mem[1769] : 1'b0;
  assign r_data_o[168] = (N3)? mem[168] : 
                         (N0)? mem[1768] : 1'b0;
  assign r_data_o[167] = (N3)? mem[167] : 
                         (N0)? mem[1767] : 1'b0;
  assign r_data_o[166] = (N3)? mem[166] : 
                         (N0)? mem[1766] : 1'b0;
  assign r_data_o[165] = (N3)? mem[165] : 
                         (N0)? mem[1765] : 1'b0;
  assign r_data_o[164] = (N3)? mem[164] : 
                         (N0)? mem[1764] : 1'b0;
  assign r_data_o[163] = (N3)? mem[163] : 
                         (N0)? mem[1763] : 1'b0;
  assign r_data_o[162] = (N3)? mem[162] : 
                         (N0)? mem[1762] : 1'b0;
  assign r_data_o[161] = (N3)? mem[161] : 
                         (N0)? mem[1761] : 1'b0;
  assign r_data_o[160] = (N3)? mem[160] : 
                         (N0)? mem[1760] : 1'b0;
  assign r_data_o[159] = (N3)? mem[159] : 
                         (N0)? mem[1759] : 1'b0;
  assign r_data_o[158] = (N3)? mem[158] : 
                         (N0)? mem[1758] : 1'b0;
  assign r_data_o[157] = (N3)? mem[157] : 
                         (N0)? mem[1757] : 1'b0;
  assign r_data_o[156] = (N3)? mem[156] : 
                         (N0)? mem[1756] : 1'b0;
  assign r_data_o[155] = (N3)? mem[155] : 
                         (N0)? mem[1755] : 1'b0;
  assign r_data_o[154] = (N3)? mem[154] : 
                         (N0)? mem[1754] : 1'b0;
  assign r_data_o[153] = (N3)? mem[153] : 
                         (N0)? mem[1753] : 1'b0;
  assign r_data_o[152] = (N3)? mem[152] : 
                         (N0)? mem[1752] : 1'b0;
  assign r_data_o[151] = (N3)? mem[151] : 
                         (N0)? mem[1751] : 1'b0;
  assign r_data_o[150] = (N3)? mem[150] : 
                         (N0)? mem[1750] : 1'b0;
  assign r_data_o[149] = (N3)? mem[149] : 
                         (N0)? mem[1749] : 1'b0;
  assign r_data_o[148] = (N3)? mem[148] : 
                         (N0)? mem[1748] : 1'b0;
  assign r_data_o[147] = (N3)? mem[147] : 
                         (N0)? mem[1747] : 1'b0;
  assign r_data_o[146] = (N3)? mem[146] : 
                         (N0)? mem[1746] : 1'b0;
  assign r_data_o[145] = (N3)? mem[145] : 
                         (N0)? mem[1745] : 1'b0;
  assign r_data_o[144] = (N3)? mem[144] : 
                         (N0)? mem[1744] : 1'b0;
  assign r_data_o[143] = (N3)? mem[143] : 
                         (N0)? mem[1743] : 1'b0;
  assign r_data_o[142] = (N3)? mem[142] : 
                         (N0)? mem[1742] : 1'b0;
  assign r_data_o[141] = (N3)? mem[141] : 
                         (N0)? mem[1741] : 1'b0;
  assign r_data_o[140] = (N3)? mem[140] : 
                         (N0)? mem[1740] : 1'b0;
  assign r_data_o[139] = (N3)? mem[139] : 
                         (N0)? mem[1739] : 1'b0;
  assign r_data_o[138] = (N3)? mem[138] : 
                         (N0)? mem[1738] : 1'b0;
  assign r_data_o[137] = (N3)? mem[137] : 
                         (N0)? mem[1737] : 1'b0;
  assign r_data_o[136] = (N3)? mem[136] : 
                         (N0)? mem[1736] : 1'b0;
  assign r_data_o[135] = (N3)? mem[135] : 
                         (N0)? mem[1735] : 1'b0;
  assign r_data_o[134] = (N3)? mem[134] : 
                         (N0)? mem[1734] : 1'b0;
  assign r_data_o[133] = (N3)? mem[133] : 
                         (N0)? mem[1733] : 1'b0;
  assign r_data_o[132] = (N3)? mem[132] : 
                         (N0)? mem[1732] : 1'b0;
  assign r_data_o[131] = (N3)? mem[131] : 
                         (N0)? mem[1731] : 1'b0;
  assign r_data_o[130] = (N3)? mem[130] : 
                         (N0)? mem[1730] : 1'b0;
  assign r_data_o[129] = (N3)? mem[129] : 
                         (N0)? mem[1729] : 1'b0;
  assign r_data_o[128] = (N3)? mem[128] : 
                         (N0)? mem[1728] : 1'b0;
  assign r_data_o[127] = (N3)? mem[127] : 
                         (N0)? mem[1727] : 1'b0;
  assign r_data_o[126] = (N3)? mem[126] : 
                         (N0)? mem[1726] : 1'b0;
  assign r_data_o[125] = (N3)? mem[125] : 
                         (N0)? mem[1725] : 1'b0;
  assign r_data_o[124] = (N3)? mem[124] : 
                         (N0)? mem[1724] : 1'b0;
  assign r_data_o[123] = (N3)? mem[123] : 
                         (N0)? mem[1723] : 1'b0;
  assign r_data_o[122] = (N3)? mem[122] : 
                         (N0)? mem[1722] : 1'b0;
  assign r_data_o[121] = (N3)? mem[121] : 
                         (N0)? mem[1721] : 1'b0;
  assign r_data_o[120] = (N3)? mem[120] : 
                         (N0)? mem[1720] : 1'b0;
  assign r_data_o[119] = (N3)? mem[119] : 
                         (N0)? mem[1719] : 1'b0;
  assign r_data_o[118] = (N3)? mem[118] : 
                         (N0)? mem[1718] : 1'b0;
  assign r_data_o[117] = (N3)? mem[117] : 
                         (N0)? mem[1717] : 1'b0;
  assign r_data_o[116] = (N3)? mem[116] : 
                         (N0)? mem[1716] : 1'b0;
  assign r_data_o[115] = (N3)? mem[115] : 
                         (N0)? mem[1715] : 1'b0;
  assign r_data_o[114] = (N3)? mem[114] : 
                         (N0)? mem[1714] : 1'b0;
  assign r_data_o[113] = (N3)? mem[113] : 
                         (N0)? mem[1713] : 1'b0;
  assign r_data_o[112] = (N3)? mem[112] : 
                         (N0)? mem[1712] : 1'b0;
  assign r_data_o[111] = (N3)? mem[111] : 
                         (N0)? mem[1711] : 1'b0;
  assign r_data_o[110] = (N3)? mem[110] : 
                         (N0)? mem[1710] : 1'b0;
  assign r_data_o[109] = (N3)? mem[109] : 
                         (N0)? mem[1709] : 1'b0;
  assign r_data_o[108] = (N3)? mem[108] : 
                         (N0)? mem[1708] : 1'b0;
  assign r_data_o[107] = (N3)? mem[107] : 
                         (N0)? mem[1707] : 1'b0;
  assign r_data_o[106] = (N3)? mem[106] : 
                         (N0)? mem[1706] : 1'b0;
  assign r_data_o[105] = (N3)? mem[105] : 
                         (N0)? mem[1705] : 1'b0;
  assign r_data_o[104] = (N3)? mem[104] : 
                         (N0)? mem[1704] : 1'b0;
  assign r_data_o[103] = (N3)? mem[103] : 
                         (N0)? mem[1703] : 1'b0;
  assign r_data_o[102] = (N3)? mem[102] : 
                         (N0)? mem[1702] : 1'b0;
  assign r_data_o[101] = (N3)? mem[101] : 
                         (N0)? mem[1701] : 1'b0;
  assign r_data_o[100] = (N3)? mem[100] : 
                         (N0)? mem[1700] : 1'b0;
  assign r_data_o[99] = (N3)? mem[99] : 
                        (N0)? mem[1699] : 1'b0;
  assign r_data_o[98] = (N3)? mem[98] : 
                        (N0)? mem[1698] : 1'b0;
  assign r_data_o[97] = (N3)? mem[97] : 
                        (N0)? mem[1697] : 1'b0;
  assign r_data_o[96] = (N3)? mem[96] : 
                        (N0)? mem[1696] : 1'b0;
  assign r_data_o[95] = (N3)? mem[95] : 
                        (N0)? mem[1695] : 1'b0;
  assign r_data_o[94] = (N3)? mem[94] : 
                        (N0)? mem[1694] : 1'b0;
  assign r_data_o[93] = (N3)? mem[93] : 
                        (N0)? mem[1693] : 1'b0;
  assign r_data_o[92] = (N3)? mem[92] : 
                        (N0)? mem[1692] : 1'b0;
  assign r_data_o[91] = (N3)? mem[91] : 
                        (N0)? mem[1691] : 1'b0;
  assign r_data_o[90] = (N3)? mem[90] : 
                        (N0)? mem[1690] : 1'b0;
  assign r_data_o[89] = (N3)? mem[89] : 
                        (N0)? mem[1689] : 1'b0;
  assign r_data_o[88] = (N3)? mem[88] : 
                        (N0)? mem[1688] : 1'b0;
  assign r_data_o[87] = (N3)? mem[87] : 
                        (N0)? mem[1687] : 1'b0;
  assign r_data_o[86] = (N3)? mem[86] : 
                        (N0)? mem[1686] : 1'b0;
  assign r_data_o[85] = (N3)? mem[85] : 
                        (N0)? mem[1685] : 1'b0;
  assign r_data_o[84] = (N3)? mem[84] : 
                        (N0)? mem[1684] : 1'b0;
  assign r_data_o[83] = (N3)? mem[83] : 
                        (N0)? mem[1683] : 1'b0;
  assign r_data_o[82] = (N3)? mem[82] : 
                        (N0)? mem[1682] : 1'b0;
  assign r_data_o[81] = (N3)? mem[81] : 
                        (N0)? mem[1681] : 1'b0;
  assign r_data_o[80] = (N3)? mem[80] : 
                        (N0)? mem[1680] : 1'b0;
  assign r_data_o[79] = (N3)? mem[79] : 
                        (N0)? mem[1679] : 1'b0;
  assign r_data_o[78] = (N3)? mem[78] : 
                        (N0)? mem[1678] : 1'b0;
  assign r_data_o[77] = (N3)? mem[77] : 
                        (N0)? mem[1677] : 1'b0;
  assign r_data_o[76] = (N3)? mem[76] : 
                        (N0)? mem[1676] : 1'b0;
  assign r_data_o[75] = (N3)? mem[75] : 
                        (N0)? mem[1675] : 1'b0;
  assign r_data_o[74] = (N3)? mem[74] : 
                        (N0)? mem[1674] : 1'b0;
  assign r_data_o[73] = (N3)? mem[73] : 
                        (N0)? mem[1673] : 1'b0;
  assign r_data_o[72] = (N3)? mem[72] : 
                        (N0)? mem[1672] : 1'b0;
  assign r_data_o[71] = (N3)? mem[71] : 
                        (N0)? mem[1671] : 1'b0;
  assign r_data_o[70] = (N3)? mem[70] : 
                        (N0)? mem[1670] : 1'b0;
  assign r_data_o[69] = (N3)? mem[69] : 
                        (N0)? mem[1669] : 1'b0;
  assign r_data_o[68] = (N3)? mem[68] : 
                        (N0)? mem[1668] : 1'b0;
  assign r_data_o[67] = (N3)? mem[67] : 
                        (N0)? mem[1667] : 1'b0;
  assign r_data_o[66] = (N3)? mem[66] : 
                        (N0)? mem[1666] : 1'b0;
  assign r_data_o[65] = (N3)? mem[65] : 
                        (N0)? mem[1665] : 1'b0;
  assign r_data_o[64] = (N3)? mem[64] : 
                        (N0)? mem[1664] : 1'b0;
  assign r_data_o[63] = (N3)? mem[63] : 
                        (N0)? mem[1663] : 1'b0;
  assign r_data_o[62] = (N3)? mem[62] : 
                        (N0)? mem[1662] : 1'b0;
  assign r_data_o[61] = (N3)? mem[61] : 
                        (N0)? mem[1661] : 1'b0;
  assign r_data_o[60] = (N3)? mem[60] : 
                        (N0)? mem[1660] : 1'b0;
  assign r_data_o[59] = (N3)? mem[59] : 
                        (N0)? mem[1659] : 1'b0;
  assign r_data_o[58] = (N3)? mem[58] : 
                        (N0)? mem[1658] : 1'b0;
  assign r_data_o[57] = (N3)? mem[57] : 
                        (N0)? mem[1657] : 1'b0;
  assign r_data_o[56] = (N3)? mem[56] : 
                        (N0)? mem[1656] : 1'b0;
  assign r_data_o[55] = (N3)? mem[55] : 
                        (N0)? mem[1655] : 1'b0;
  assign r_data_o[54] = (N3)? mem[54] : 
                        (N0)? mem[1654] : 1'b0;
  assign r_data_o[53] = (N3)? mem[53] : 
                        (N0)? mem[1653] : 1'b0;
  assign r_data_o[52] = (N3)? mem[52] : 
                        (N0)? mem[1652] : 1'b0;
  assign r_data_o[51] = (N3)? mem[51] : 
                        (N0)? mem[1651] : 1'b0;
  assign r_data_o[50] = (N3)? mem[50] : 
                        (N0)? mem[1650] : 1'b0;
  assign r_data_o[49] = (N3)? mem[49] : 
                        (N0)? mem[1649] : 1'b0;
  assign r_data_o[48] = (N3)? mem[48] : 
                        (N0)? mem[1648] : 1'b0;
  assign r_data_o[47] = (N3)? mem[47] : 
                        (N0)? mem[1647] : 1'b0;
  assign r_data_o[46] = (N3)? mem[46] : 
                        (N0)? mem[1646] : 1'b0;
  assign r_data_o[45] = (N3)? mem[45] : 
                        (N0)? mem[1645] : 1'b0;
  assign r_data_o[44] = (N3)? mem[44] : 
                        (N0)? mem[1644] : 1'b0;
  assign r_data_o[43] = (N3)? mem[43] : 
                        (N0)? mem[1643] : 1'b0;
  assign r_data_o[42] = (N3)? mem[42] : 
                        (N0)? mem[1642] : 1'b0;
  assign r_data_o[41] = (N3)? mem[41] : 
                        (N0)? mem[1641] : 1'b0;
  assign r_data_o[40] = (N3)? mem[40] : 
                        (N0)? mem[1640] : 1'b0;
  assign r_data_o[39] = (N3)? mem[39] : 
                        (N0)? mem[1639] : 1'b0;
  assign r_data_o[38] = (N3)? mem[38] : 
                        (N0)? mem[1638] : 1'b0;
  assign r_data_o[37] = (N3)? mem[37] : 
                        (N0)? mem[1637] : 1'b0;
  assign r_data_o[36] = (N3)? mem[36] : 
                        (N0)? mem[1636] : 1'b0;
  assign r_data_o[35] = (N3)? mem[35] : 
                        (N0)? mem[1635] : 1'b0;
  assign r_data_o[34] = (N3)? mem[34] : 
                        (N0)? mem[1634] : 1'b0;
  assign r_data_o[33] = (N3)? mem[33] : 
                        (N0)? mem[1633] : 1'b0;
  assign r_data_o[32] = (N3)? mem[32] : 
                        (N0)? mem[1632] : 1'b0;
  assign r_data_o[31] = (N3)? mem[31] : 
                        (N0)? mem[1631] : 1'b0;
  assign r_data_o[30] = (N3)? mem[30] : 
                        (N0)? mem[1630] : 1'b0;
  assign r_data_o[29] = (N3)? mem[29] : 
                        (N0)? mem[1629] : 1'b0;
  assign r_data_o[28] = (N3)? mem[28] : 
                        (N0)? mem[1628] : 1'b0;
  assign r_data_o[27] = (N3)? mem[27] : 
                        (N0)? mem[1627] : 1'b0;
  assign r_data_o[26] = (N3)? mem[26] : 
                        (N0)? mem[1626] : 1'b0;
  assign r_data_o[25] = (N3)? mem[25] : 
                        (N0)? mem[1625] : 1'b0;
  assign r_data_o[24] = (N3)? mem[24] : 
                        (N0)? mem[1624] : 1'b0;
  assign r_data_o[23] = (N3)? mem[23] : 
                        (N0)? mem[1623] : 1'b0;
  assign r_data_o[22] = (N3)? mem[22] : 
                        (N0)? mem[1622] : 1'b0;
  assign r_data_o[21] = (N3)? mem[21] : 
                        (N0)? mem[1621] : 1'b0;
  assign r_data_o[20] = (N3)? mem[20] : 
                        (N0)? mem[1620] : 1'b0;
  assign r_data_o[19] = (N3)? mem[19] : 
                        (N0)? mem[1619] : 1'b0;
  assign r_data_o[18] = (N3)? mem[18] : 
                        (N0)? mem[1618] : 1'b0;
  assign r_data_o[17] = (N3)? mem[17] : 
                        (N0)? mem[1617] : 1'b0;
  assign r_data_o[16] = (N3)? mem[16] : 
                        (N0)? mem[1616] : 1'b0;
  assign r_data_o[15] = (N3)? mem[15] : 
                        (N0)? mem[1615] : 1'b0;
  assign r_data_o[14] = (N3)? mem[14] : 
                        (N0)? mem[1614] : 1'b0;
  assign r_data_o[13] = (N3)? mem[13] : 
                        (N0)? mem[1613] : 1'b0;
  assign r_data_o[12] = (N3)? mem[12] : 
                        (N0)? mem[1612] : 1'b0;
  assign r_data_o[11] = (N3)? mem[11] : 
                        (N0)? mem[1611] : 1'b0;
  assign r_data_o[10] = (N3)? mem[10] : 
                        (N0)? mem[1610] : 1'b0;
  assign r_data_o[9] = (N3)? mem[9] : 
                       (N0)? mem[1609] : 1'b0;
  assign r_data_o[8] = (N3)? mem[8] : 
                       (N0)? mem[1608] : 1'b0;
  assign r_data_o[7] = (N3)? mem[7] : 
                       (N0)? mem[1607] : 1'b0;
  assign r_data_o[6] = (N3)? mem[6] : 
                       (N0)? mem[1606] : 1'b0;
  assign r_data_o[5] = (N3)? mem[5] : 
                       (N0)? mem[1605] : 1'b0;
  assign r_data_o[4] = (N3)? mem[4] : 
                       (N0)? mem[1604] : 1'b0;
  assign r_data_o[3] = (N3)? mem[3] : 
                       (N0)? mem[1603] : 1'b0;
  assign r_data_o[2] = (N3)? mem[2] : 
                       (N0)? mem[1602] : 1'b0;
  assign r_data_o[1] = (N3)? mem[1] : 
                       (N0)? mem[1601] : 1'b0;
  assign r_data_o[0] = (N3)? mem[0] : 
                       (N0)? mem[1600] : 1'b0;
  assign N5 = ~w_addr_i[0];
  assign { N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, N12, N11, N10, N9, N8, N7 } = (N1)? { w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], w_addr_i[0:0], N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5, N5 } : 
                                                                                                                                                                           (N2)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N1 = w_v_i;
  assign N2 = N4;
  assign N3 = ~r_addr_i[0];
  assign N4 = ~w_v_i;

  always @(posedge w_clk_i) begin
    if(N23) begin
      { mem[3199:3101], mem[1600:1600] } <= { w_data_i[1599:1501], w_data_i[0:0] };
    end 
    if(N24) begin
      { mem[3100:3002], mem[1601:1601] } <= { w_data_i[1500:1402], w_data_i[1:1] };
    end 
    if(N25) begin
      { mem[3001:2903], mem[1602:1602] } <= { w_data_i[1401:1303], w_data_i[2:2] };
    end 
    if(N26) begin
      { mem[2902:2804], mem[1603:1603] } <= { w_data_i[1302:1204], w_data_i[3:3] };
    end 
    if(N27) begin
      { mem[2803:2705], mem[1604:1604] } <= { w_data_i[1203:1105], w_data_i[4:4] };
    end 
    if(N28) begin
      { mem[2704:2606], mem[1605:1605] } <= { w_data_i[1104:1006], w_data_i[5:5] };
    end 
    if(N29) begin
      { mem[2605:2507], mem[1606:1606] } <= { w_data_i[1005:907], w_data_i[6:6] };
    end 
    if(N30) begin
      { mem[2506:2408], mem[1607:1607] } <= { w_data_i[906:808], w_data_i[7:7] };
    end 
    if(N31) begin
      { mem[2407:2309], mem[1608:1608] } <= { w_data_i[807:709], w_data_i[8:8] };
    end 
    if(N32) begin
      { mem[2308:2210], mem[1609:1609] } <= { w_data_i[708:610], w_data_i[9:9] };
    end 
    if(N33) begin
      { mem[2209:2111], mem[1610:1610] } <= { w_data_i[609:511], w_data_i[10:10] };
    end 
    if(N34) begin
      { mem[2110:2012], mem[1611:1611] } <= { w_data_i[510:412], w_data_i[11:11] };
    end 
    if(N35) begin
      { mem[2011:1913], mem[1612:1612] } <= { w_data_i[411:313], w_data_i[12:12] };
    end 
    if(N36) begin
      { mem[1912:1814], mem[1613:1613] } <= { w_data_i[312:214], w_data_i[13:13] };
    end 
    if(N37) begin
      { mem[1813:1715], mem[1614:1614] } <= { w_data_i[213:115], w_data_i[14:14] };
    end 
    if(N38) begin
      { mem[1714:1615] } <= { w_data_i[114:15] };
    end 
    if(N7) begin
      { mem[1599:1501], mem[0:0] } <= { w_data_i[1599:1501], w_data_i[0:0] };
    end 
    if(N8) begin
      { mem[1500:1402], mem[1:1] } <= { w_data_i[1500:1402], w_data_i[1:1] };
    end 
    if(N9) begin
      { mem[1401:1303], mem[2:2] } <= { w_data_i[1401:1303], w_data_i[2:2] };
    end 
    if(N10) begin
      { mem[1302:1204], mem[3:3] } <= { w_data_i[1302:1204], w_data_i[3:3] };
    end 
    if(N11) begin
      { mem[1203:1105], mem[4:4] } <= { w_data_i[1203:1105], w_data_i[4:4] };
    end 
    if(N12) begin
      { mem[1104:1006], mem[5:5] } <= { w_data_i[1104:1006], w_data_i[5:5] };
    end 
    if(N13) begin
      { mem[1005:907], mem[6:6] } <= { w_data_i[1005:907], w_data_i[6:6] };
    end 
    if(N14) begin
      { mem[906:808], mem[7:7] } <= { w_data_i[906:808], w_data_i[7:7] };
    end 
    if(N15) begin
      { mem[807:709], mem[8:8] } <= { w_data_i[807:709], w_data_i[8:8] };
    end 
    if(N16) begin
      { mem[708:610], mem[9:9] } <= { w_data_i[708:610], w_data_i[9:9] };
    end 
    if(N17) begin
      { mem[609:511], mem[10:10] } <= { w_data_i[609:511], w_data_i[10:10] };
    end 
    if(N18) begin
      { mem[510:412], mem[11:11] } <= { w_data_i[510:412], w_data_i[11:11] };
    end 
    if(N19) begin
      { mem[411:313], mem[12:12] } <= { w_data_i[411:313], w_data_i[12:12] };
    end 
    if(N20) begin
      { mem[312:214], mem[13:13] } <= { w_data_i[312:214], w_data_i[13:13] };
    end 
    if(N21) begin
      { mem[213:115], mem[14:14] } <= { w_data_i[213:115], w_data_i[14:14] };
    end 
    if(N22) begin
      { mem[114:15] } <= { w_data_i[114:15] };
    end 
  end


endmodule



module bsg_mem_1r1w_width_p1600_els_p2_read_write_same_addr_p0
(
  w_clk_i,
  w_reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [0:0] w_addr_i;
  input [1599:0] w_data_i;
  input [0:0] r_addr_i;
  output [1599:0] r_data_o;
  input w_clk_i;
  input w_reset_i;
  input w_v_i;
  input r_v_i;
  wire [1599:0] r_data_o;

  bsg_mem_1r1w_synth_width_p1600_els_p2_read_write_same_addr_p0_harden_p0
  synth
  (
    .w_clk_i(w_clk_i),
    .w_reset_i(w_reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i[0]),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i[0]),
    .r_data_o(r_data_o)
  );


endmodule



module bsg_two_fifo_width_p1600
(
  clk_i,
  reset_i,
  ready_o,
  data_i,
  v_i,
  v_o,
  data_o,
  yumi_i
);

  input [1599:0] data_i;
  output [1599:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [1599:0] data_o;
  wire ready_o,v_o,N0,N1,enq_i,n_0_net_,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,
  N15,N16,N17,N18,N19,N20,N21,N22,N23,N24;
  reg full_r,tail_r,head_r,empty_r;

  bsg_mem_1r1w_width_p1600_els_p2_read_write_same_addr_p0
  mem_1r1w
  (
    .w_clk_i(clk_i),
    .w_reset_i(reset_i),
    .w_v_i(enq_i),
    .w_addr_i(tail_r),
    .w_data_i(data_i),
    .r_v_i(n_0_net_),
    .r_addr_i(head_r),
    .r_data_o(data_o)
  );

  assign N9 = (N0)? 1'b1 : 
              (N1)? N5 : 1'b0;
  assign N0 = N3;
  assign N1 = N2;
  assign N10 = (N0)? 1'b0 : 
               (N1)? N4 : 1'b0;
  assign N11 = (N0)? 1'b1 : 
               (N1)? yumi_i : 1'b0;
  assign N12 = (N0)? 1'b0 : 
               (N1)? N6 : 1'b0;
  assign N13 = (N0)? 1'b1 : 
               (N1)? N7 : 1'b0;
  assign N14 = (N0)? 1'b0 : 
               (N1)? N8 : 1'b0;
  assign n_0_net_ = ~empty_r;
  assign v_o = ~empty_r;
  assign ready_o = ~full_r;
  assign enq_i = v_i & N15;
  assign N15 = ~full_r;
  assign N2 = ~reset_i;
  assign N3 = reset_i;
  assign N5 = enq_i;
  assign N4 = ~tail_r;
  assign N6 = ~head_r;
  assign N7 = N17 | N19;
  assign N17 = empty_r & N16;
  assign N16 = ~enq_i;
  assign N19 = N18 & N16;
  assign N18 = N15 & yumi_i;
  assign N8 = N23 | N24;
  assign N23 = N21 & N22;
  assign N21 = N20 & enq_i;
  assign N20 = ~empty_r;
  assign N22 = ~yumi_i;
  assign N24 = full_r & N22;

  always @(posedge clk_i) begin
    if(1'b1) begin
      full_r <= N14;
      empty_r <= N13;
    end 
    if(N9) begin
      tail_r <= N10;
    end 
    if(N11) begin
      head_r <= N12;
    end 
  end


endmodule



module bsg_counter_clear_up_max_val_p49_init_val_p0
(
  clk_i,
  reset_i,
  clear_i,
  up_i,
  count_o
);

  output [5:0] count_o;
  input clk_i;
  input reset_i;
  input clear_i;
  input up_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23;
  reg [5:0] count_o;
  assign { N11, N10, N9, N8, N7, N6 } = { N23, N22, N21, N20, N19, N18 } + up_i;
  assign { N17, N16, N15, N14, N13, N12 } = (N0)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                            (N1)? { N11, N10, N9, N8, N7, N6 } : 1'b0;
  assign N0 = reset_i;
  assign N1 = N2;
  assign { N23, N22, N21, N20, N19, N18 } = count_o * N4;
  assign N2 = ~reset_i;
  assign N3 = N2;
  assign N4 = ~clear_i;
  assign N5 = N3 & N4;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { count_o[5:0] } <= { N17, N16, N15, N14, N13, N12 };
    end 
  end


endmodule



module bsg_mux_width_p32_els_p50
(
  data_i,
  sel_i,
  data_o
);

  input [1599:0] data_i;
  input [5:0] sel_i;
  output [31:0] data_o;
  wire [31:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312;
  assign N0 = N4 & N5;
  assign N1 = N0 & N6;
  assign N2 = N1 & N7;
  assign N3 = N2 & N8;
  assign N263 = N3 & N9;
  assign N4 = ~sel_i[5];
  assign N5 = ~sel_i[4];
  assign N6 = ~sel_i[3];
  assign N7 = ~sel_i[2];
  assign N8 = ~sel_i[0];
  assign N9 = ~sel_i[1];
  assign N10 = sel_i[5] & N14;
  assign N11 = N10 & N15;
  assign N12 = N11 & N16;
  assign N13 = N12 & N17;
  assign N264 = N13 & N18;
  assign N14 = ~sel_i[4];
  assign N15 = ~sel_i[3];
  assign N16 = ~sel_i[2];
  assign N17 = ~sel_i[0];
  assign N18 = ~sel_i[1];
  assign N19 = N23 & N24;
  assign N20 = N19 & N25;
  assign N21 = N20 & N26;
  assign N22 = N21 & sel_i[0];
  assign N265 = N22 & N27;
  assign N23 = ~sel_i[5];
  assign N24 = ~sel_i[4];
  assign N25 = ~sel_i[3];
  assign N26 = ~sel_i[2];
  assign N27 = ~sel_i[1];
  assign N28 = N32 & N33;
  assign N29 = N28 & N34;
  assign N30 = N29 & N35;
  assign N31 = N30 & N36;
  assign N267 = N31 & sel_i[1];
  assign N32 = ~sel_i[5];
  assign N33 = ~sel_i[4];
  assign N34 = ~sel_i[3];
  assign N35 = ~sel_i[2];
  assign N36 = ~sel_i[0];
  assign N37 = N41 & N42;
  assign N38 = N37 & N43;
  assign N39 = N38 & N44;
  assign N40 = N39 & sel_i[0];
  assign N269 = N40 & sel_i[1];
  assign N41 = ~sel_i[5];
  assign N42 = ~sel_i[4];
  assign N43 = ~sel_i[3];
  assign N44 = ~sel_i[2];
  assign N45 = N49 & N50;
  assign N46 = N45 & N51;
  assign N47 = N46 & sel_i[2];
  assign N48 = N47 & N52;
  assign N271 = N48 & N53;
  assign N49 = ~sel_i[5];
  assign N50 = ~sel_i[4];
  assign N51 = ~sel_i[3];
  assign N52 = ~sel_i[0];
  assign N53 = ~sel_i[1];
  assign N54 = N58 & N59;
  assign N55 = N54 & N60;
  assign N56 = N55 & sel_i[2];
  assign N57 = N56 & sel_i[0];
  assign N273 = N57 & N61;
  assign N58 = ~sel_i[5];
  assign N59 = ~sel_i[4];
  assign N60 = ~sel_i[3];
  assign N61 = ~sel_i[1];
  assign N62 = N66 & N67;
  assign N63 = N62 & N68;
  assign N64 = N63 & sel_i[2];
  assign N65 = N64 & N69;
  assign N275 = N65 & sel_i[1];
  assign N66 = ~sel_i[5];
  assign N67 = ~sel_i[4];
  assign N68 = ~sel_i[3];
  assign N69 = ~sel_i[0];
  assign N70 = N74 & N75;
  assign N71 = N70 & N76;
  assign N72 = N71 & sel_i[2];
  assign N73 = N72 & sel_i[0];
  assign N277 = N73 & sel_i[1];
  assign N74 = ~sel_i[5];
  assign N75 = ~sel_i[4];
  assign N76 = ~sel_i[3];
  assign N77 = N81 & N82;
  assign N78 = N77 & sel_i[3];
  assign N79 = N78 & N83;
  assign N80 = N79 & N84;
  assign N279 = N80 & N85;
  assign N81 = ~sel_i[5];
  assign N82 = ~sel_i[4];
  assign N83 = ~sel_i[2];
  assign N84 = ~sel_i[0];
  assign N85 = ~sel_i[1];
  assign N86 = N90 & N91;
  assign N87 = N86 & sel_i[3];
  assign N88 = N87 & N92;
  assign N89 = N88 & sel_i[0];
  assign N281 = N89 & N93;
  assign N90 = ~sel_i[5];
  assign N91 = ~sel_i[4];
  assign N92 = ~sel_i[2];
  assign N93 = ~sel_i[1];
  assign N94 = N98 & N99;
  assign N95 = N94 & sel_i[3];
  assign N96 = N95 & N100;
  assign N97 = N96 & N101;
  assign N283 = N97 & sel_i[1];
  assign N98 = ~sel_i[5];
  assign N99 = ~sel_i[4];
  assign N100 = ~sel_i[2];
  assign N101 = ~sel_i[0];
  assign N102 = N106 & N107;
  assign N103 = N102 & sel_i[3];
  assign N104 = N103 & N108;
  assign N105 = N104 & sel_i[0];
  assign N285 = N105 & sel_i[1];
  assign N106 = ~sel_i[5];
  assign N107 = ~sel_i[4];
  assign N108 = ~sel_i[2];
  assign N109 = N113 & N114;
  assign N110 = N109 & sel_i[3];
  assign N111 = N110 & sel_i[2];
  assign N112 = N111 & N115;
  assign N287 = N112 & N116;
  assign N113 = ~sel_i[5];
  assign N114 = ~sel_i[4];
  assign N115 = ~sel_i[0];
  assign N116 = ~sel_i[1];
  assign N117 = N121 & N122;
  assign N118 = N117 & sel_i[3];
  assign N119 = N118 & sel_i[2];
  assign N120 = N119 & sel_i[0];
  assign N289 = N120 & N123;
  assign N121 = ~sel_i[5];
  assign N122 = ~sel_i[4];
  assign N123 = ~sel_i[1];
  assign N124 = N128 & N129;
  assign N125 = N124 & sel_i[3];
  assign N126 = N125 & sel_i[2];
  assign N127 = N126 & N130;
  assign N291 = N127 & sel_i[1];
  assign N128 = ~sel_i[5];
  assign N129 = ~sel_i[4];
  assign N130 = ~sel_i[0];
  assign N131 = N135 & N136;
  assign N132 = N131 & sel_i[3];
  assign N133 = N132 & sel_i[2];
  assign N134 = N133 & sel_i[0];
  assign N293 = N134 & sel_i[1];
  assign N135 = ~sel_i[5];
  assign N136 = ~sel_i[4];
  assign N137 = N141 & sel_i[4];
  assign N138 = N137 & N142;
  assign N139 = N138 & N143;
  assign N140 = N139 & N144;
  assign N295 = N140 & N145;
  assign N141 = ~sel_i[5];
  assign N142 = ~sel_i[3];
  assign N143 = ~sel_i[2];
  assign N144 = ~sel_i[0];
  assign N145 = ~sel_i[1];
  assign N146 = N150 & sel_i[4];
  assign N147 = N146 & N151;
  assign N148 = N147 & N152;
  assign N149 = N148 & sel_i[0];
  assign N297 = N149 & N153;
  assign N150 = ~sel_i[5];
  assign N151 = ~sel_i[3];
  assign N152 = ~sel_i[2];
  assign N153 = ~sel_i[1];
  assign N299 = sel_i[4] & N154 & (N155 & N156) & sel_i[1];
  assign N154 = ~sel_i[3];
  assign N155 = ~sel_i[2];
  assign N156 = ~sel_i[0];
  assign N300 = sel_i[4] & N157 & (N158 & sel_i[0]) & sel_i[1];
  assign N157 = ~sel_i[3];
  assign N158 = ~sel_i[2];
  assign N301 = sel_i[4] & N159 & (sel_i[2] & N160) & N161;
  assign N159 = ~sel_i[3];
  assign N160 = ~sel_i[0];
  assign N161 = ~sel_i[1];
  assign N302 = sel_i[4] & N162 & (sel_i[2] & sel_i[0]) & N163;
  assign N162 = ~sel_i[3];
  assign N163 = ~sel_i[1];
  assign N303 = sel_i[4] & N164 & (sel_i[2] & N165) & sel_i[1];
  assign N164 = ~sel_i[3];
  assign N165 = ~sel_i[0];
  assign N304 = sel_i[4] & N166 & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N166 = ~sel_i[3];
  assign N305 = sel_i[4] & sel_i[3] & (N167 & N168) & N169;
  assign N167 = ~sel_i[2];
  assign N168 = ~sel_i[0];
  assign N169 = ~sel_i[1];
  assign N306 = sel_i[4] & sel_i[3] & (N170 & sel_i[0]) & N171;
  assign N170 = ~sel_i[2];
  assign N171 = ~sel_i[1];
  assign N307 = sel_i[4] & sel_i[3] & (N172 & N173) & sel_i[1];
  assign N172 = ~sel_i[2];
  assign N173 = ~sel_i[0];
  assign N308 = sel_i[4] & sel_i[3] & (N174 & sel_i[0]) & sel_i[1];
  assign N174 = ~sel_i[2];
  assign N309 = sel_i[4] & sel_i[3] & (sel_i[2] & N175) & N176;
  assign N175 = ~sel_i[0];
  assign N176 = ~sel_i[1];
  assign N310 = sel_i[4] & sel_i[3] & (sel_i[2] & sel_i[0]) & N177;
  assign N177 = ~sel_i[1];
  assign N311 = sel_i[4] & sel_i[3] & (sel_i[2] & N178) & sel_i[1];
  assign N178 = ~sel_i[0];
  assign N312 = sel_i[4] & sel_i[3] & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N179 = sel_i[5] & N183;
  assign N180 = N179 & N184;
  assign N181 = N180 & N185;
  assign N182 = N181 & sel_i[0];
  assign N266 = N182 & N186;
  assign N183 = ~sel_i[4];
  assign N184 = ~sel_i[3];
  assign N185 = ~sel_i[2];
  assign N186 = ~sel_i[1];
  assign N268 = sel_i[5] & N187 & (N188 & N189) & sel_i[1];
  assign N187 = ~sel_i[3];
  assign N188 = ~sel_i[2];
  assign N189 = ~sel_i[0];
  assign N270 = sel_i[5] & N190 & (N191 & sel_i[0]) & sel_i[1];
  assign N190 = ~sel_i[3];
  assign N191 = ~sel_i[2];
  assign N272 = sel_i[5] & N192 & (sel_i[2] & N193) & N194;
  assign N192 = ~sel_i[3];
  assign N193 = ~sel_i[0];
  assign N194 = ~sel_i[1];
  assign N274 = sel_i[5] & N195 & (sel_i[2] & sel_i[0]) & N196;
  assign N195 = ~sel_i[3];
  assign N196 = ~sel_i[1];
  assign N276 = sel_i[5] & N197 & (sel_i[2] & N198) & sel_i[1];
  assign N197 = ~sel_i[3];
  assign N198 = ~sel_i[0];
  assign N278 = sel_i[5] & N199 & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N199 = ~sel_i[3];
  assign N280 = sel_i[5] & sel_i[3] & (N200 & N201) & N202;
  assign N200 = ~sel_i[2];
  assign N201 = ~sel_i[0];
  assign N202 = ~sel_i[1];
  assign N282 = sel_i[5] & sel_i[3] & (N203 & sel_i[0]) & N204;
  assign N203 = ~sel_i[2];
  assign N204 = ~sel_i[1];
  assign N284 = sel_i[5] & sel_i[3] & (N205 & N206) & sel_i[1];
  assign N205 = ~sel_i[2];
  assign N206 = ~sel_i[0];
  assign N286 = sel_i[5] & sel_i[3] & (N207 & sel_i[0]) & sel_i[1];
  assign N207 = ~sel_i[2];
  assign N288 = sel_i[5] & sel_i[3] & (sel_i[2] & N208) & N209;
  assign N208 = ~sel_i[0];
  assign N209 = ~sel_i[1];
  assign N290 = sel_i[5] & sel_i[3] & (sel_i[2] & sel_i[0]) & N210;
  assign N210 = ~sel_i[1];
  assign N292 = sel_i[5] & sel_i[3] & (sel_i[2] & N211) & sel_i[1];
  assign N211 = ~sel_i[0];
  assign N294 = sel_i[5] & sel_i[3] & (sel_i[2] & sel_i[0]) & sel_i[1];
  assign N296 = sel_i[5] & sel_i[4] & N212;
  assign N212 = ~sel_i[0];
  assign N298 = sel_i[5] & sel_i[4] & sel_i[0];
  assign data_o[31] = (N213)? data_i[31] : 
                      (N214)? data_i[63] : 
                      (N215)? data_i[95] : 
                      (N216)? data_i[127] : 
                      (N217)? data_i[159] : 
                      (N218)? data_i[191] : 
                      (N219)? data_i[223] : 
                      (N220)? data_i[255] : 
                      (N221)? data_i[287] : 
                      (N222)? data_i[319] : 
                      (N223)? data_i[351] : 
                      (N224)? data_i[383] : 
                      (N225)? data_i[415] : 
                      (N226)? data_i[447] : 
                      (N227)? data_i[479] : 
                      (N228)? data_i[511] : 
                      (N229)? data_i[543] : 
                      (N230)? data_i[575] : 
                      (N231)? data_i[607] : 
                      (N232)? data_i[639] : 
                      (N233)? data_i[671] : 
                      (N234)? data_i[703] : 
                      (N235)? data_i[735] : 
                      (N236)? data_i[767] : 
                      (N237)? data_i[799] : 
                      (N238)? data_i[831] : 
                      (N239)? data_i[863] : 
                      (N240)? data_i[895] : 
                      (N241)? data_i[927] : 
                      (N242)? data_i[959] : 
                      (N243)? data_i[991] : 
                      (N244)? data_i[1023] : 
                      (N245)? data_i[1055] : 
                      (N246)? data_i[1087] : 
                      (N247)? data_i[1119] : 
                      (N248)? data_i[1151] : 
                      (N249)? data_i[1183] : 
                      (N250)? data_i[1215] : 
                      (N251)? data_i[1247] : 
                      (N252)? data_i[1279] : 
                      (N253)? data_i[1311] : 
                      (N254)? data_i[1343] : 
                      (N255)? data_i[1375] : 
                      (N256)? data_i[1407] : 
                      (N257)? data_i[1439] : 
                      (N258)? data_i[1471] : 
                      (N259)? data_i[1503] : 
                      (N260)? data_i[1535] : 
                      (N261)? data_i[1567] : 
                      (N262)? data_i[1599] : 1'b0;
  assign N213 = N263;
  assign N214 = N265;
  assign N215 = N267;
  assign N216 = N269;
  assign N217 = N271;
  assign N218 = N273;
  assign N219 = N275;
  assign N220 = N277;
  assign N221 = N279;
  assign N222 = N281;
  assign N223 = N283;
  assign N224 = N285;
  assign N225 = N287;
  assign N226 = N289;
  assign N227 = N291;
  assign N228 = N293;
  assign N229 = N295;
  assign N230 = N297;
  assign N231 = N299;
  assign N232 = N300;
  assign N233 = N301;
  assign N234 = N302;
  assign N235 = N303;
  assign N236 = N304;
  assign N237 = N305;
  assign N238 = N306;
  assign N239 = N307;
  assign N240 = N308;
  assign N241 = N309;
  assign N242 = N310;
  assign N243 = N311;
  assign N244 = N312;
  assign N245 = N264;
  assign N246 = N266;
  assign N247 = N268;
  assign N248 = N270;
  assign N249 = N272;
  assign N250 = N274;
  assign N251 = N276;
  assign N252 = N278;
  assign N253 = N280;
  assign N254 = N282;
  assign N255 = N284;
  assign N256 = N286;
  assign N257 = N288;
  assign N258 = N290;
  assign N259 = N292;
  assign N260 = N294;
  assign N261 = N296;
  assign N262 = N298;
  assign data_o[30] = (N213)? data_i[30] : 
                      (N214)? data_i[62] : 
                      (N215)? data_i[94] : 
                      (N216)? data_i[126] : 
                      (N217)? data_i[158] : 
                      (N218)? data_i[190] : 
                      (N219)? data_i[222] : 
                      (N220)? data_i[254] : 
                      (N221)? data_i[286] : 
                      (N222)? data_i[318] : 
                      (N223)? data_i[350] : 
                      (N224)? data_i[382] : 
                      (N225)? data_i[414] : 
                      (N226)? data_i[446] : 
                      (N227)? data_i[478] : 
                      (N228)? data_i[510] : 
                      (N229)? data_i[542] : 
                      (N230)? data_i[574] : 
                      (N231)? data_i[606] : 
                      (N232)? data_i[638] : 
                      (N233)? data_i[670] : 
                      (N234)? data_i[702] : 
                      (N235)? data_i[734] : 
                      (N236)? data_i[766] : 
                      (N237)? data_i[798] : 
                      (N238)? data_i[830] : 
                      (N239)? data_i[862] : 
                      (N240)? data_i[894] : 
                      (N241)? data_i[926] : 
                      (N242)? data_i[958] : 
                      (N243)? data_i[990] : 
                      (N244)? data_i[1022] : 
                      (N245)? data_i[1054] : 
                      (N246)? data_i[1086] : 
                      (N247)? data_i[1118] : 
                      (N248)? data_i[1150] : 
                      (N249)? data_i[1182] : 
                      (N250)? data_i[1214] : 
                      (N251)? data_i[1246] : 
                      (N252)? data_i[1278] : 
                      (N253)? data_i[1310] : 
                      (N254)? data_i[1342] : 
                      (N255)? data_i[1374] : 
                      (N256)? data_i[1406] : 
                      (N257)? data_i[1438] : 
                      (N258)? data_i[1470] : 
                      (N259)? data_i[1502] : 
                      (N260)? data_i[1534] : 
                      (N261)? data_i[1566] : 
                      (N262)? data_i[1598] : 1'b0;
  assign data_o[29] = (N213)? data_i[29] : 
                      (N214)? data_i[61] : 
                      (N215)? data_i[93] : 
                      (N216)? data_i[125] : 
                      (N217)? data_i[157] : 
                      (N218)? data_i[189] : 
                      (N219)? data_i[221] : 
                      (N220)? data_i[253] : 
                      (N221)? data_i[285] : 
                      (N222)? data_i[317] : 
                      (N223)? data_i[349] : 
                      (N224)? data_i[381] : 
                      (N225)? data_i[413] : 
                      (N226)? data_i[445] : 
                      (N227)? data_i[477] : 
                      (N228)? data_i[509] : 
                      (N229)? data_i[541] : 
                      (N230)? data_i[573] : 
                      (N231)? data_i[605] : 
                      (N232)? data_i[637] : 
                      (N233)? data_i[669] : 
                      (N234)? data_i[701] : 
                      (N235)? data_i[733] : 
                      (N236)? data_i[765] : 
                      (N237)? data_i[797] : 
                      (N238)? data_i[829] : 
                      (N239)? data_i[861] : 
                      (N240)? data_i[893] : 
                      (N241)? data_i[925] : 
                      (N242)? data_i[957] : 
                      (N243)? data_i[989] : 
                      (N244)? data_i[1021] : 
                      (N245)? data_i[1053] : 
                      (N246)? data_i[1085] : 
                      (N247)? data_i[1117] : 
                      (N248)? data_i[1149] : 
                      (N249)? data_i[1181] : 
                      (N250)? data_i[1213] : 
                      (N251)? data_i[1245] : 
                      (N252)? data_i[1277] : 
                      (N253)? data_i[1309] : 
                      (N254)? data_i[1341] : 
                      (N255)? data_i[1373] : 
                      (N256)? data_i[1405] : 
                      (N257)? data_i[1437] : 
                      (N258)? data_i[1469] : 
                      (N259)? data_i[1501] : 
                      (N260)? data_i[1533] : 
                      (N261)? data_i[1565] : 
                      (N262)? data_i[1597] : 1'b0;
  assign data_o[28] = (N213)? data_i[28] : 
                      (N214)? data_i[60] : 
                      (N215)? data_i[92] : 
                      (N216)? data_i[124] : 
                      (N217)? data_i[156] : 
                      (N218)? data_i[188] : 
                      (N219)? data_i[220] : 
                      (N220)? data_i[252] : 
                      (N221)? data_i[284] : 
                      (N222)? data_i[316] : 
                      (N223)? data_i[348] : 
                      (N224)? data_i[380] : 
                      (N225)? data_i[412] : 
                      (N226)? data_i[444] : 
                      (N227)? data_i[476] : 
                      (N228)? data_i[508] : 
                      (N229)? data_i[540] : 
                      (N230)? data_i[572] : 
                      (N231)? data_i[604] : 
                      (N232)? data_i[636] : 
                      (N233)? data_i[668] : 
                      (N234)? data_i[700] : 
                      (N235)? data_i[732] : 
                      (N236)? data_i[764] : 
                      (N237)? data_i[796] : 
                      (N238)? data_i[828] : 
                      (N239)? data_i[860] : 
                      (N240)? data_i[892] : 
                      (N241)? data_i[924] : 
                      (N242)? data_i[956] : 
                      (N243)? data_i[988] : 
                      (N244)? data_i[1020] : 
                      (N245)? data_i[1052] : 
                      (N246)? data_i[1084] : 
                      (N247)? data_i[1116] : 
                      (N248)? data_i[1148] : 
                      (N249)? data_i[1180] : 
                      (N250)? data_i[1212] : 
                      (N251)? data_i[1244] : 
                      (N252)? data_i[1276] : 
                      (N253)? data_i[1308] : 
                      (N254)? data_i[1340] : 
                      (N255)? data_i[1372] : 
                      (N256)? data_i[1404] : 
                      (N257)? data_i[1436] : 
                      (N258)? data_i[1468] : 
                      (N259)? data_i[1500] : 
                      (N260)? data_i[1532] : 
                      (N261)? data_i[1564] : 
                      (N262)? data_i[1596] : 1'b0;
  assign data_o[27] = (N213)? data_i[27] : 
                      (N214)? data_i[59] : 
                      (N215)? data_i[91] : 
                      (N216)? data_i[123] : 
                      (N217)? data_i[155] : 
                      (N218)? data_i[187] : 
                      (N219)? data_i[219] : 
                      (N220)? data_i[251] : 
                      (N221)? data_i[283] : 
                      (N222)? data_i[315] : 
                      (N223)? data_i[347] : 
                      (N224)? data_i[379] : 
                      (N225)? data_i[411] : 
                      (N226)? data_i[443] : 
                      (N227)? data_i[475] : 
                      (N228)? data_i[507] : 
                      (N229)? data_i[539] : 
                      (N230)? data_i[571] : 
                      (N231)? data_i[603] : 
                      (N232)? data_i[635] : 
                      (N233)? data_i[667] : 
                      (N234)? data_i[699] : 
                      (N235)? data_i[731] : 
                      (N236)? data_i[763] : 
                      (N237)? data_i[795] : 
                      (N238)? data_i[827] : 
                      (N239)? data_i[859] : 
                      (N240)? data_i[891] : 
                      (N241)? data_i[923] : 
                      (N242)? data_i[955] : 
                      (N243)? data_i[987] : 
                      (N244)? data_i[1019] : 
                      (N245)? data_i[1051] : 
                      (N246)? data_i[1083] : 
                      (N247)? data_i[1115] : 
                      (N248)? data_i[1147] : 
                      (N249)? data_i[1179] : 
                      (N250)? data_i[1211] : 
                      (N251)? data_i[1243] : 
                      (N252)? data_i[1275] : 
                      (N253)? data_i[1307] : 
                      (N254)? data_i[1339] : 
                      (N255)? data_i[1371] : 
                      (N256)? data_i[1403] : 
                      (N257)? data_i[1435] : 
                      (N258)? data_i[1467] : 
                      (N259)? data_i[1499] : 
                      (N260)? data_i[1531] : 
                      (N261)? data_i[1563] : 
                      (N262)? data_i[1595] : 1'b0;
  assign data_o[26] = (N213)? data_i[26] : 
                      (N214)? data_i[58] : 
                      (N215)? data_i[90] : 
                      (N216)? data_i[122] : 
                      (N217)? data_i[154] : 
                      (N218)? data_i[186] : 
                      (N219)? data_i[218] : 
                      (N220)? data_i[250] : 
                      (N221)? data_i[282] : 
                      (N222)? data_i[314] : 
                      (N223)? data_i[346] : 
                      (N224)? data_i[378] : 
                      (N225)? data_i[410] : 
                      (N226)? data_i[442] : 
                      (N227)? data_i[474] : 
                      (N228)? data_i[506] : 
                      (N229)? data_i[538] : 
                      (N230)? data_i[570] : 
                      (N231)? data_i[602] : 
                      (N232)? data_i[634] : 
                      (N233)? data_i[666] : 
                      (N234)? data_i[698] : 
                      (N235)? data_i[730] : 
                      (N236)? data_i[762] : 
                      (N237)? data_i[794] : 
                      (N238)? data_i[826] : 
                      (N239)? data_i[858] : 
                      (N240)? data_i[890] : 
                      (N241)? data_i[922] : 
                      (N242)? data_i[954] : 
                      (N243)? data_i[986] : 
                      (N244)? data_i[1018] : 
                      (N245)? data_i[1050] : 
                      (N246)? data_i[1082] : 
                      (N247)? data_i[1114] : 
                      (N248)? data_i[1146] : 
                      (N249)? data_i[1178] : 
                      (N250)? data_i[1210] : 
                      (N251)? data_i[1242] : 
                      (N252)? data_i[1274] : 
                      (N253)? data_i[1306] : 
                      (N254)? data_i[1338] : 
                      (N255)? data_i[1370] : 
                      (N256)? data_i[1402] : 
                      (N257)? data_i[1434] : 
                      (N258)? data_i[1466] : 
                      (N259)? data_i[1498] : 
                      (N260)? data_i[1530] : 
                      (N261)? data_i[1562] : 
                      (N262)? data_i[1594] : 1'b0;
  assign data_o[25] = (N213)? data_i[25] : 
                      (N214)? data_i[57] : 
                      (N215)? data_i[89] : 
                      (N216)? data_i[121] : 
                      (N217)? data_i[153] : 
                      (N218)? data_i[185] : 
                      (N219)? data_i[217] : 
                      (N220)? data_i[249] : 
                      (N221)? data_i[281] : 
                      (N222)? data_i[313] : 
                      (N223)? data_i[345] : 
                      (N224)? data_i[377] : 
                      (N225)? data_i[409] : 
                      (N226)? data_i[441] : 
                      (N227)? data_i[473] : 
                      (N228)? data_i[505] : 
                      (N229)? data_i[537] : 
                      (N230)? data_i[569] : 
                      (N231)? data_i[601] : 
                      (N232)? data_i[633] : 
                      (N233)? data_i[665] : 
                      (N234)? data_i[697] : 
                      (N235)? data_i[729] : 
                      (N236)? data_i[761] : 
                      (N237)? data_i[793] : 
                      (N238)? data_i[825] : 
                      (N239)? data_i[857] : 
                      (N240)? data_i[889] : 
                      (N241)? data_i[921] : 
                      (N242)? data_i[953] : 
                      (N243)? data_i[985] : 
                      (N244)? data_i[1017] : 
                      (N245)? data_i[1049] : 
                      (N246)? data_i[1081] : 
                      (N247)? data_i[1113] : 
                      (N248)? data_i[1145] : 
                      (N249)? data_i[1177] : 
                      (N250)? data_i[1209] : 
                      (N251)? data_i[1241] : 
                      (N252)? data_i[1273] : 
                      (N253)? data_i[1305] : 
                      (N254)? data_i[1337] : 
                      (N255)? data_i[1369] : 
                      (N256)? data_i[1401] : 
                      (N257)? data_i[1433] : 
                      (N258)? data_i[1465] : 
                      (N259)? data_i[1497] : 
                      (N260)? data_i[1529] : 
                      (N261)? data_i[1561] : 
                      (N262)? data_i[1593] : 1'b0;
  assign data_o[24] = (N213)? data_i[24] : 
                      (N214)? data_i[56] : 
                      (N215)? data_i[88] : 
                      (N216)? data_i[120] : 
                      (N217)? data_i[152] : 
                      (N218)? data_i[184] : 
                      (N219)? data_i[216] : 
                      (N220)? data_i[248] : 
                      (N221)? data_i[280] : 
                      (N222)? data_i[312] : 
                      (N223)? data_i[344] : 
                      (N224)? data_i[376] : 
                      (N225)? data_i[408] : 
                      (N226)? data_i[440] : 
                      (N227)? data_i[472] : 
                      (N228)? data_i[504] : 
                      (N229)? data_i[536] : 
                      (N230)? data_i[568] : 
                      (N231)? data_i[600] : 
                      (N232)? data_i[632] : 
                      (N233)? data_i[664] : 
                      (N234)? data_i[696] : 
                      (N235)? data_i[728] : 
                      (N236)? data_i[760] : 
                      (N237)? data_i[792] : 
                      (N238)? data_i[824] : 
                      (N239)? data_i[856] : 
                      (N240)? data_i[888] : 
                      (N241)? data_i[920] : 
                      (N242)? data_i[952] : 
                      (N243)? data_i[984] : 
                      (N244)? data_i[1016] : 
                      (N245)? data_i[1048] : 
                      (N246)? data_i[1080] : 
                      (N247)? data_i[1112] : 
                      (N248)? data_i[1144] : 
                      (N249)? data_i[1176] : 
                      (N250)? data_i[1208] : 
                      (N251)? data_i[1240] : 
                      (N252)? data_i[1272] : 
                      (N253)? data_i[1304] : 
                      (N254)? data_i[1336] : 
                      (N255)? data_i[1368] : 
                      (N256)? data_i[1400] : 
                      (N257)? data_i[1432] : 
                      (N258)? data_i[1464] : 
                      (N259)? data_i[1496] : 
                      (N260)? data_i[1528] : 
                      (N261)? data_i[1560] : 
                      (N262)? data_i[1592] : 1'b0;
  assign data_o[23] = (N213)? data_i[23] : 
                      (N214)? data_i[55] : 
                      (N215)? data_i[87] : 
                      (N216)? data_i[119] : 
                      (N217)? data_i[151] : 
                      (N218)? data_i[183] : 
                      (N219)? data_i[215] : 
                      (N220)? data_i[247] : 
                      (N221)? data_i[279] : 
                      (N222)? data_i[311] : 
                      (N223)? data_i[343] : 
                      (N224)? data_i[375] : 
                      (N225)? data_i[407] : 
                      (N226)? data_i[439] : 
                      (N227)? data_i[471] : 
                      (N228)? data_i[503] : 
                      (N229)? data_i[535] : 
                      (N230)? data_i[567] : 
                      (N231)? data_i[599] : 
                      (N232)? data_i[631] : 
                      (N233)? data_i[663] : 
                      (N234)? data_i[695] : 
                      (N235)? data_i[727] : 
                      (N236)? data_i[759] : 
                      (N237)? data_i[791] : 
                      (N238)? data_i[823] : 
                      (N239)? data_i[855] : 
                      (N240)? data_i[887] : 
                      (N241)? data_i[919] : 
                      (N242)? data_i[951] : 
                      (N243)? data_i[983] : 
                      (N244)? data_i[1015] : 
                      (N245)? data_i[1047] : 
                      (N246)? data_i[1079] : 
                      (N247)? data_i[1111] : 
                      (N248)? data_i[1143] : 
                      (N249)? data_i[1175] : 
                      (N250)? data_i[1207] : 
                      (N251)? data_i[1239] : 
                      (N252)? data_i[1271] : 
                      (N253)? data_i[1303] : 
                      (N254)? data_i[1335] : 
                      (N255)? data_i[1367] : 
                      (N256)? data_i[1399] : 
                      (N257)? data_i[1431] : 
                      (N258)? data_i[1463] : 
                      (N259)? data_i[1495] : 
                      (N260)? data_i[1527] : 
                      (N261)? data_i[1559] : 
                      (N262)? data_i[1591] : 1'b0;
  assign data_o[22] = (N213)? data_i[22] : 
                      (N214)? data_i[54] : 
                      (N215)? data_i[86] : 
                      (N216)? data_i[118] : 
                      (N217)? data_i[150] : 
                      (N218)? data_i[182] : 
                      (N219)? data_i[214] : 
                      (N220)? data_i[246] : 
                      (N221)? data_i[278] : 
                      (N222)? data_i[310] : 
                      (N223)? data_i[342] : 
                      (N224)? data_i[374] : 
                      (N225)? data_i[406] : 
                      (N226)? data_i[438] : 
                      (N227)? data_i[470] : 
                      (N228)? data_i[502] : 
                      (N229)? data_i[534] : 
                      (N230)? data_i[566] : 
                      (N231)? data_i[598] : 
                      (N232)? data_i[630] : 
                      (N233)? data_i[662] : 
                      (N234)? data_i[694] : 
                      (N235)? data_i[726] : 
                      (N236)? data_i[758] : 
                      (N237)? data_i[790] : 
                      (N238)? data_i[822] : 
                      (N239)? data_i[854] : 
                      (N240)? data_i[886] : 
                      (N241)? data_i[918] : 
                      (N242)? data_i[950] : 
                      (N243)? data_i[982] : 
                      (N244)? data_i[1014] : 
                      (N245)? data_i[1046] : 
                      (N246)? data_i[1078] : 
                      (N247)? data_i[1110] : 
                      (N248)? data_i[1142] : 
                      (N249)? data_i[1174] : 
                      (N250)? data_i[1206] : 
                      (N251)? data_i[1238] : 
                      (N252)? data_i[1270] : 
                      (N253)? data_i[1302] : 
                      (N254)? data_i[1334] : 
                      (N255)? data_i[1366] : 
                      (N256)? data_i[1398] : 
                      (N257)? data_i[1430] : 
                      (N258)? data_i[1462] : 
                      (N259)? data_i[1494] : 
                      (N260)? data_i[1526] : 
                      (N261)? data_i[1558] : 
                      (N262)? data_i[1590] : 1'b0;
  assign data_o[21] = (N213)? data_i[21] : 
                      (N214)? data_i[53] : 
                      (N215)? data_i[85] : 
                      (N216)? data_i[117] : 
                      (N217)? data_i[149] : 
                      (N218)? data_i[181] : 
                      (N219)? data_i[213] : 
                      (N220)? data_i[245] : 
                      (N221)? data_i[277] : 
                      (N222)? data_i[309] : 
                      (N223)? data_i[341] : 
                      (N224)? data_i[373] : 
                      (N225)? data_i[405] : 
                      (N226)? data_i[437] : 
                      (N227)? data_i[469] : 
                      (N228)? data_i[501] : 
                      (N229)? data_i[533] : 
                      (N230)? data_i[565] : 
                      (N231)? data_i[597] : 
                      (N232)? data_i[629] : 
                      (N233)? data_i[661] : 
                      (N234)? data_i[693] : 
                      (N235)? data_i[725] : 
                      (N236)? data_i[757] : 
                      (N237)? data_i[789] : 
                      (N238)? data_i[821] : 
                      (N239)? data_i[853] : 
                      (N240)? data_i[885] : 
                      (N241)? data_i[917] : 
                      (N242)? data_i[949] : 
                      (N243)? data_i[981] : 
                      (N244)? data_i[1013] : 
                      (N245)? data_i[1045] : 
                      (N246)? data_i[1077] : 
                      (N247)? data_i[1109] : 
                      (N248)? data_i[1141] : 
                      (N249)? data_i[1173] : 
                      (N250)? data_i[1205] : 
                      (N251)? data_i[1237] : 
                      (N252)? data_i[1269] : 
                      (N253)? data_i[1301] : 
                      (N254)? data_i[1333] : 
                      (N255)? data_i[1365] : 
                      (N256)? data_i[1397] : 
                      (N257)? data_i[1429] : 
                      (N258)? data_i[1461] : 
                      (N259)? data_i[1493] : 
                      (N260)? data_i[1525] : 
                      (N261)? data_i[1557] : 
                      (N262)? data_i[1589] : 1'b0;
  assign data_o[20] = (N213)? data_i[20] : 
                      (N214)? data_i[52] : 
                      (N215)? data_i[84] : 
                      (N216)? data_i[116] : 
                      (N217)? data_i[148] : 
                      (N218)? data_i[180] : 
                      (N219)? data_i[212] : 
                      (N220)? data_i[244] : 
                      (N221)? data_i[276] : 
                      (N222)? data_i[308] : 
                      (N223)? data_i[340] : 
                      (N224)? data_i[372] : 
                      (N225)? data_i[404] : 
                      (N226)? data_i[436] : 
                      (N227)? data_i[468] : 
                      (N228)? data_i[500] : 
                      (N229)? data_i[532] : 
                      (N230)? data_i[564] : 
                      (N231)? data_i[596] : 
                      (N232)? data_i[628] : 
                      (N233)? data_i[660] : 
                      (N234)? data_i[692] : 
                      (N235)? data_i[724] : 
                      (N236)? data_i[756] : 
                      (N237)? data_i[788] : 
                      (N238)? data_i[820] : 
                      (N239)? data_i[852] : 
                      (N240)? data_i[884] : 
                      (N241)? data_i[916] : 
                      (N242)? data_i[948] : 
                      (N243)? data_i[980] : 
                      (N244)? data_i[1012] : 
                      (N245)? data_i[1044] : 
                      (N246)? data_i[1076] : 
                      (N247)? data_i[1108] : 
                      (N248)? data_i[1140] : 
                      (N249)? data_i[1172] : 
                      (N250)? data_i[1204] : 
                      (N251)? data_i[1236] : 
                      (N252)? data_i[1268] : 
                      (N253)? data_i[1300] : 
                      (N254)? data_i[1332] : 
                      (N255)? data_i[1364] : 
                      (N256)? data_i[1396] : 
                      (N257)? data_i[1428] : 
                      (N258)? data_i[1460] : 
                      (N259)? data_i[1492] : 
                      (N260)? data_i[1524] : 
                      (N261)? data_i[1556] : 
                      (N262)? data_i[1588] : 1'b0;
  assign data_o[19] = (N213)? data_i[19] : 
                      (N214)? data_i[51] : 
                      (N215)? data_i[83] : 
                      (N216)? data_i[115] : 
                      (N217)? data_i[147] : 
                      (N218)? data_i[179] : 
                      (N219)? data_i[211] : 
                      (N220)? data_i[243] : 
                      (N221)? data_i[275] : 
                      (N222)? data_i[307] : 
                      (N223)? data_i[339] : 
                      (N224)? data_i[371] : 
                      (N225)? data_i[403] : 
                      (N226)? data_i[435] : 
                      (N227)? data_i[467] : 
                      (N228)? data_i[499] : 
                      (N229)? data_i[531] : 
                      (N230)? data_i[563] : 
                      (N231)? data_i[595] : 
                      (N232)? data_i[627] : 
                      (N233)? data_i[659] : 
                      (N234)? data_i[691] : 
                      (N235)? data_i[723] : 
                      (N236)? data_i[755] : 
                      (N237)? data_i[787] : 
                      (N238)? data_i[819] : 
                      (N239)? data_i[851] : 
                      (N240)? data_i[883] : 
                      (N241)? data_i[915] : 
                      (N242)? data_i[947] : 
                      (N243)? data_i[979] : 
                      (N244)? data_i[1011] : 
                      (N245)? data_i[1043] : 
                      (N246)? data_i[1075] : 
                      (N247)? data_i[1107] : 
                      (N248)? data_i[1139] : 
                      (N249)? data_i[1171] : 
                      (N250)? data_i[1203] : 
                      (N251)? data_i[1235] : 
                      (N252)? data_i[1267] : 
                      (N253)? data_i[1299] : 
                      (N254)? data_i[1331] : 
                      (N255)? data_i[1363] : 
                      (N256)? data_i[1395] : 
                      (N257)? data_i[1427] : 
                      (N258)? data_i[1459] : 
                      (N259)? data_i[1491] : 
                      (N260)? data_i[1523] : 
                      (N261)? data_i[1555] : 
                      (N262)? data_i[1587] : 1'b0;
  assign data_o[18] = (N213)? data_i[18] : 
                      (N214)? data_i[50] : 
                      (N215)? data_i[82] : 
                      (N216)? data_i[114] : 
                      (N217)? data_i[146] : 
                      (N218)? data_i[178] : 
                      (N219)? data_i[210] : 
                      (N220)? data_i[242] : 
                      (N221)? data_i[274] : 
                      (N222)? data_i[306] : 
                      (N223)? data_i[338] : 
                      (N224)? data_i[370] : 
                      (N225)? data_i[402] : 
                      (N226)? data_i[434] : 
                      (N227)? data_i[466] : 
                      (N228)? data_i[498] : 
                      (N229)? data_i[530] : 
                      (N230)? data_i[562] : 
                      (N231)? data_i[594] : 
                      (N232)? data_i[626] : 
                      (N233)? data_i[658] : 
                      (N234)? data_i[690] : 
                      (N235)? data_i[722] : 
                      (N236)? data_i[754] : 
                      (N237)? data_i[786] : 
                      (N238)? data_i[818] : 
                      (N239)? data_i[850] : 
                      (N240)? data_i[882] : 
                      (N241)? data_i[914] : 
                      (N242)? data_i[946] : 
                      (N243)? data_i[978] : 
                      (N244)? data_i[1010] : 
                      (N245)? data_i[1042] : 
                      (N246)? data_i[1074] : 
                      (N247)? data_i[1106] : 
                      (N248)? data_i[1138] : 
                      (N249)? data_i[1170] : 
                      (N250)? data_i[1202] : 
                      (N251)? data_i[1234] : 
                      (N252)? data_i[1266] : 
                      (N253)? data_i[1298] : 
                      (N254)? data_i[1330] : 
                      (N255)? data_i[1362] : 
                      (N256)? data_i[1394] : 
                      (N257)? data_i[1426] : 
                      (N258)? data_i[1458] : 
                      (N259)? data_i[1490] : 
                      (N260)? data_i[1522] : 
                      (N261)? data_i[1554] : 
                      (N262)? data_i[1586] : 1'b0;
  assign data_o[17] = (N213)? data_i[17] : 
                      (N214)? data_i[49] : 
                      (N215)? data_i[81] : 
                      (N216)? data_i[113] : 
                      (N217)? data_i[145] : 
                      (N218)? data_i[177] : 
                      (N219)? data_i[209] : 
                      (N220)? data_i[241] : 
                      (N221)? data_i[273] : 
                      (N222)? data_i[305] : 
                      (N223)? data_i[337] : 
                      (N224)? data_i[369] : 
                      (N225)? data_i[401] : 
                      (N226)? data_i[433] : 
                      (N227)? data_i[465] : 
                      (N228)? data_i[497] : 
                      (N229)? data_i[529] : 
                      (N230)? data_i[561] : 
                      (N231)? data_i[593] : 
                      (N232)? data_i[625] : 
                      (N233)? data_i[657] : 
                      (N234)? data_i[689] : 
                      (N235)? data_i[721] : 
                      (N236)? data_i[753] : 
                      (N237)? data_i[785] : 
                      (N238)? data_i[817] : 
                      (N239)? data_i[849] : 
                      (N240)? data_i[881] : 
                      (N241)? data_i[913] : 
                      (N242)? data_i[945] : 
                      (N243)? data_i[977] : 
                      (N244)? data_i[1009] : 
                      (N245)? data_i[1041] : 
                      (N246)? data_i[1073] : 
                      (N247)? data_i[1105] : 
                      (N248)? data_i[1137] : 
                      (N249)? data_i[1169] : 
                      (N250)? data_i[1201] : 
                      (N251)? data_i[1233] : 
                      (N252)? data_i[1265] : 
                      (N253)? data_i[1297] : 
                      (N254)? data_i[1329] : 
                      (N255)? data_i[1361] : 
                      (N256)? data_i[1393] : 
                      (N257)? data_i[1425] : 
                      (N258)? data_i[1457] : 
                      (N259)? data_i[1489] : 
                      (N260)? data_i[1521] : 
                      (N261)? data_i[1553] : 
                      (N262)? data_i[1585] : 1'b0;
  assign data_o[16] = (N213)? data_i[16] : 
                      (N214)? data_i[48] : 
                      (N215)? data_i[80] : 
                      (N216)? data_i[112] : 
                      (N217)? data_i[144] : 
                      (N218)? data_i[176] : 
                      (N219)? data_i[208] : 
                      (N220)? data_i[240] : 
                      (N221)? data_i[272] : 
                      (N222)? data_i[304] : 
                      (N223)? data_i[336] : 
                      (N224)? data_i[368] : 
                      (N225)? data_i[400] : 
                      (N226)? data_i[432] : 
                      (N227)? data_i[464] : 
                      (N228)? data_i[496] : 
                      (N229)? data_i[528] : 
                      (N230)? data_i[560] : 
                      (N231)? data_i[592] : 
                      (N232)? data_i[624] : 
                      (N233)? data_i[656] : 
                      (N234)? data_i[688] : 
                      (N235)? data_i[720] : 
                      (N236)? data_i[752] : 
                      (N237)? data_i[784] : 
                      (N238)? data_i[816] : 
                      (N239)? data_i[848] : 
                      (N240)? data_i[880] : 
                      (N241)? data_i[912] : 
                      (N242)? data_i[944] : 
                      (N243)? data_i[976] : 
                      (N244)? data_i[1008] : 
                      (N245)? data_i[1040] : 
                      (N246)? data_i[1072] : 
                      (N247)? data_i[1104] : 
                      (N248)? data_i[1136] : 
                      (N249)? data_i[1168] : 
                      (N250)? data_i[1200] : 
                      (N251)? data_i[1232] : 
                      (N252)? data_i[1264] : 
                      (N253)? data_i[1296] : 
                      (N254)? data_i[1328] : 
                      (N255)? data_i[1360] : 
                      (N256)? data_i[1392] : 
                      (N257)? data_i[1424] : 
                      (N258)? data_i[1456] : 
                      (N259)? data_i[1488] : 
                      (N260)? data_i[1520] : 
                      (N261)? data_i[1552] : 
                      (N262)? data_i[1584] : 1'b0;
  assign data_o[15] = (N213)? data_i[15] : 
                      (N214)? data_i[47] : 
                      (N215)? data_i[79] : 
                      (N216)? data_i[111] : 
                      (N217)? data_i[143] : 
                      (N218)? data_i[175] : 
                      (N219)? data_i[207] : 
                      (N220)? data_i[239] : 
                      (N221)? data_i[271] : 
                      (N222)? data_i[303] : 
                      (N223)? data_i[335] : 
                      (N224)? data_i[367] : 
                      (N225)? data_i[399] : 
                      (N226)? data_i[431] : 
                      (N227)? data_i[463] : 
                      (N228)? data_i[495] : 
                      (N229)? data_i[527] : 
                      (N230)? data_i[559] : 
                      (N231)? data_i[591] : 
                      (N232)? data_i[623] : 
                      (N233)? data_i[655] : 
                      (N234)? data_i[687] : 
                      (N235)? data_i[719] : 
                      (N236)? data_i[751] : 
                      (N237)? data_i[783] : 
                      (N238)? data_i[815] : 
                      (N239)? data_i[847] : 
                      (N240)? data_i[879] : 
                      (N241)? data_i[911] : 
                      (N242)? data_i[943] : 
                      (N243)? data_i[975] : 
                      (N244)? data_i[1007] : 
                      (N245)? data_i[1039] : 
                      (N246)? data_i[1071] : 
                      (N247)? data_i[1103] : 
                      (N248)? data_i[1135] : 
                      (N249)? data_i[1167] : 
                      (N250)? data_i[1199] : 
                      (N251)? data_i[1231] : 
                      (N252)? data_i[1263] : 
                      (N253)? data_i[1295] : 
                      (N254)? data_i[1327] : 
                      (N255)? data_i[1359] : 
                      (N256)? data_i[1391] : 
                      (N257)? data_i[1423] : 
                      (N258)? data_i[1455] : 
                      (N259)? data_i[1487] : 
                      (N260)? data_i[1519] : 
                      (N261)? data_i[1551] : 
                      (N262)? data_i[1583] : 1'b0;
  assign data_o[14] = (N213)? data_i[14] : 
                      (N214)? data_i[46] : 
                      (N215)? data_i[78] : 
                      (N216)? data_i[110] : 
                      (N217)? data_i[142] : 
                      (N218)? data_i[174] : 
                      (N219)? data_i[206] : 
                      (N220)? data_i[238] : 
                      (N221)? data_i[270] : 
                      (N222)? data_i[302] : 
                      (N223)? data_i[334] : 
                      (N224)? data_i[366] : 
                      (N225)? data_i[398] : 
                      (N226)? data_i[430] : 
                      (N227)? data_i[462] : 
                      (N228)? data_i[494] : 
                      (N229)? data_i[526] : 
                      (N230)? data_i[558] : 
                      (N231)? data_i[590] : 
                      (N232)? data_i[622] : 
                      (N233)? data_i[654] : 
                      (N234)? data_i[686] : 
                      (N235)? data_i[718] : 
                      (N236)? data_i[750] : 
                      (N237)? data_i[782] : 
                      (N238)? data_i[814] : 
                      (N239)? data_i[846] : 
                      (N240)? data_i[878] : 
                      (N241)? data_i[910] : 
                      (N242)? data_i[942] : 
                      (N243)? data_i[974] : 
                      (N244)? data_i[1006] : 
                      (N245)? data_i[1038] : 
                      (N246)? data_i[1070] : 
                      (N247)? data_i[1102] : 
                      (N248)? data_i[1134] : 
                      (N249)? data_i[1166] : 
                      (N250)? data_i[1198] : 
                      (N251)? data_i[1230] : 
                      (N252)? data_i[1262] : 
                      (N253)? data_i[1294] : 
                      (N254)? data_i[1326] : 
                      (N255)? data_i[1358] : 
                      (N256)? data_i[1390] : 
                      (N257)? data_i[1422] : 
                      (N258)? data_i[1454] : 
                      (N259)? data_i[1486] : 
                      (N260)? data_i[1518] : 
                      (N261)? data_i[1550] : 
                      (N262)? data_i[1582] : 1'b0;
  assign data_o[13] = (N213)? data_i[13] : 
                      (N214)? data_i[45] : 
                      (N215)? data_i[77] : 
                      (N216)? data_i[109] : 
                      (N217)? data_i[141] : 
                      (N218)? data_i[173] : 
                      (N219)? data_i[205] : 
                      (N220)? data_i[237] : 
                      (N221)? data_i[269] : 
                      (N222)? data_i[301] : 
                      (N223)? data_i[333] : 
                      (N224)? data_i[365] : 
                      (N225)? data_i[397] : 
                      (N226)? data_i[429] : 
                      (N227)? data_i[461] : 
                      (N228)? data_i[493] : 
                      (N229)? data_i[525] : 
                      (N230)? data_i[557] : 
                      (N231)? data_i[589] : 
                      (N232)? data_i[621] : 
                      (N233)? data_i[653] : 
                      (N234)? data_i[685] : 
                      (N235)? data_i[717] : 
                      (N236)? data_i[749] : 
                      (N237)? data_i[781] : 
                      (N238)? data_i[813] : 
                      (N239)? data_i[845] : 
                      (N240)? data_i[877] : 
                      (N241)? data_i[909] : 
                      (N242)? data_i[941] : 
                      (N243)? data_i[973] : 
                      (N244)? data_i[1005] : 
                      (N245)? data_i[1037] : 
                      (N246)? data_i[1069] : 
                      (N247)? data_i[1101] : 
                      (N248)? data_i[1133] : 
                      (N249)? data_i[1165] : 
                      (N250)? data_i[1197] : 
                      (N251)? data_i[1229] : 
                      (N252)? data_i[1261] : 
                      (N253)? data_i[1293] : 
                      (N254)? data_i[1325] : 
                      (N255)? data_i[1357] : 
                      (N256)? data_i[1389] : 
                      (N257)? data_i[1421] : 
                      (N258)? data_i[1453] : 
                      (N259)? data_i[1485] : 
                      (N260)? data_i[1517] : 
                      (N261)? data_i[1549] : 
                      (N262)? data_i[1581] : 1'b0;
  assign data_o[12] = (N213)? data_i[12] : 
                      (N214)? data_i[44] : 
                      (N215)? data_i[76] : 
                      (N216)? data_i[108] : 
                      (N217)? data_i[140] : 
                      (N218)? data_i[172] : 
                      (N219)? data_i[204] : 
                      (N220)? data_i[236] : 
                      (N221)? data_i[268] : 
                      (N222)? data_i[300] : 
                      (N223)? data_i[332] : 
                      (N224)? data_i[364] : 
                      (N225)? data_i[396] : 
                      (N226)? data_i[428] : 
                      (N227)? data_i[460] : 
                      (N228)? data_i[492] : 
                      (N229)? data_i[524] : 
                      (N230)? data_i[556] : 
                      (N231)? data_i[588] : 
                      (N232)? data_i[620] : 
                      (N233)? data_i[652] : 
                      (N234)? data_i[684] : 
                      (N235)? data_i[716] : 
                      (N236)? data_i[748] : 
                      (N237)? data_i[780] : 
                      (N238)? data_i[812] : 
                      (N239)? data_i[844] : 
                      (N240)? data_i[876] : 
                      (N241)? data_i[908] : 
                      (N242)? data_i[940] : 
                      (N243)? data_i[972] : 
                      (N244)? data_i[1004] : 
                      (N245)? data_i[1036] : 
                      (N246)? data_i[1068] : 
                      (N247)? data_i[1100] : 
                      (N248)? data_i[1132] : 
                      (N249)? data_i[1164] : 
                      (N250)? data_i[1196] : 
                      (N251)? data_i[1228] : 
                      (N252)? data_i[1260] : 
                      (N253)? data_i[1292] : 
                      (N254)? data_i[1324] : 
                      (N255)? data_i[1356] : 
                      (N256)? data_i[1388] : 
                      (N257)? data_i[1420] : 
                      (N258)? data_i[1452] : 
                      (N259)? data_i[1484] : 
                      (N260)? data_i[1516] : 
                      (N261)? data_i[1548] : 
                      (N262)? data_i[1580] : 1'b0;
  assign data_o[11] = (N213)? data_i[11] : 
                      (N214)? data_i[43] : 
                      (N215)? data_i[75] : 
                      (N216)? data_i[107] : 
                      (N217)? data_i[139] : 
                      (N218)? data_i[171] : 
                      (N219)? data_i[203] : 
                      (N220)? data_i[235] : 
                      (N221)? data_i[267] : 
                      (N222)? data_i[299] : 
                      (N223)? data_i[331] : 
                      (N224)? data_i[363] : 
                      (N225)? data_i[395] : 
                      (N226)? data_i[427] : 
                      (N227)? data_i[459] : 
                      (N228)? data_i[491] : 
                      (N229)? data_i[523] : 
                      (N230)? data_i[555] : 
                      (N231)? data_i[587] : 
                      (N232)? data_i[619] : 
                      (N233)? data_i[651] : 
                      (N234)? data_i[683] : 
                      (N235)? data_i[715] : 
                      (N236)? data_i[747] : 
                      (N237)? data_i[779] : 
                      (N238)? data_i[811] : 
                      (N239)? data_i[843] : 
                      (N240)? data_i[875] : 
                      (N241)? data_i[907] : 
                      (N242)? data_i[939] : 
                      (N243)? data_i[971] : 
                      (N244)? data_i[1003] : 
                      (N245)? data_i[1035] : 
                      (N246)? data_i[1067] : 
                      (N247)? data_i[1099] : 
                      (N248)? data_i[1131] : 
                      (N249)? data_i[1163] : 
                      (N250)? data_i[1195] : 
                      (N251)? data_i[1227] : 
                      (N252)? data_i[1259] : 
                      (N253)? data_i[1291] : 
                      (N254)? data_i[1323] : 
                      (N255)? data_i[1355] : 
                      (N256)? data_i[1387] : 
                      (N257)? data_i[1419] : 
                      (N258)? data_i[1451] : 
                      (N259)? data_i[1483] : 
                      (N260)? data_i[1515] : 
                      (N261)? data_i[1547] : 
                      (N262)? data_i[1579] : 1'b0;
  assign data_o[10] = (N213)? data_i[10] : 
                      (N214)? data_i[42] : 
                      (N215)? data_i[74] : 
                      (N216)? data_i[106] : 
                      (N217)? data_i[138] : 
                      (N218)? data_i[170] : 
                      (N219)? data_i[202] : 
                      (N220)? data_i[234] : 
                      (N221)? data_i[266] : 
                      (N222)? data_i[298] : 
                      (N223)? data_i[330] : 
                      (N224)? data_i[362] : 
                      (N225)? data_i[394] : 
                      (N226)? data_i[426] : 
                      (N227)? data_i[458] : 
                      (N228)? data_i[490] : 
                      (N229)? data_i[522] : 
                      (N230)? data_i[554] : 
                      (N231)? data_i[586] : 
                      (N232)? data_i[618] : 
                      (N233)? data_i[650] : 
                      (N234)? data_i[682] : 
                      (N235)? data_i[714] : 
                      (N236)? data_i[746] : 
                      (N237)? data_i[778] : 
                      (N238)? data_i[810] : 
                      (N239)? data_i[842] : 
                      (N240)? data_i[874] : 
                      (N241)? data_i[906] : 
                      (N242)? data_i[938] : 
                      (N243)? data_i[970] : 
                      (N244)? data_i[1002] : 
                      (N245)? data_i[1034] : 
                      (N246)? data_i[1066] : 
                      (N247)? data_i[1098] : 
                      (N248)? data_i[1130] : 
                      (N249)? data_i[1162] : 
                      (N250)? data_i[1194] : 
                      (N251)? data_i[1226] : 
                      (N252)? data_i[1258] : 
                      (N253)? data_i[1290] : 
                      (N254)? data_i[1322] : 
                      (N255)? data_i[1354] : 
                      (N256)? data_i[1386] : 
                      (N257)? data_i[1418] : 
                      (N258)? data_i[1450] : 
                      (N259)? data_i[1482] : 
                      (N260)? data_i[1514] : 
                      (N261)? data_i[1546] : 
                      (N262)? data_i[1578] : 1'b0;
  assign data_o[9] = (N213)? data_i[9] : 
                     (N214)? data_i[41] : 
                     (N215)? data_i[73] : 
                     (N216)? data_i[105] : 
                     (N217)? data_i[137] : 
                     (N218)? data_i[169] : 
                     (N219)? data_i[201] : 
                     (N220)? data_i[233] : 
                     (N221)? data_i[265] : 
                     (N222)? data_i[297] : 
                     (N223)? data_i[329] : 
                     (N224)? data_i[361] : 
                     (N225)? data_i[393] : 
                     (N226)? data_i[425] : 
                     (N227)? data_i[457] : 
                     (N228)? data_i[489] : 
                     (N229)? data_i[521] : 
                     (N230)? data_i[553] : 
                     (N231)? data_i[585] : 
                     (N232)? data_i[617] : 
                     (N233)? data_i[649] : 
                     (N234)? data_i[681] : 
                     (N235)? data_i[713] : 
                     (N236)? data_i[745] : 
                     (N237)? data_i[777] : 
                     (N238)? data_i[809] : 
                     (N239)? data_i[841] : 
                     (N240)? data_i[873] : 
                     (N241)? data_i[905] : 
                     (N242)? data_i[937] : 
                     (N243)? data_i[969] : 
                     (N244)? data_i[1001] : 
                     (N245)? data_i[1033] : 
                     (N246)? data_i[1065] : 
                     (N247)? data_i[1097] : 
                     (N248)? data_i[1129] : 
                     (N249)? data_i[1161] : 
                     (N250)? data_i[1193] : 
                     (N251)? data_i[1225] : 
                     (N252)? data_i[1257] : 
                     (N253)? data_i[1289] : 
                     (N254)? data_i[1321] : 
                     (N255)? data_i[1353] : 
                     (N256)? data_i[1385] : 
                     (N257)? data_i[1417] : 
                     (N258)? data_i[1449] : 
                     (N259)? data_i[1481] : 
                     (N260)? data_i[1513] : 
                     (N261)? data_i[1545] : 
                     (N262)? data_i[1577] : 1'b0;
  assign data_o[8] = (N213)? data_i[8] : 
                     (N214)? data_i[40] : 
                     (N215)? data_i[72] : 
                     (N216)? data_i[104] : 
                     (N217)? data_i[136] : 
                     (N218)? data_i[168] : 
                     (N219)? data_i[200] : 
                     (N220)? data_i[232] : 
                     (N221)? data_i[264] : 
                     (N222)? data_i[296] : 
                     (N223)? data_i[328] : 
                     (N224)? data_i[360] : 
                     (N225)? data_i[392] : 
                     (N226)? data_i[424] : 
                     (N227)? data_i[456] : 
                     (N228)? data_i[488] : 
                     (N229)? data_i[520] : 
                     (N230)? data_i[552] : 
                     (N231)? data_i[584] : 
                     (N232)? data_i[616] : 
                     (N233)? data_i[648] : 
                     (N234)? data_i[680] : 
                     (N235)? data_i[712] : 
                     (N236)? data_i[744] : 
                     (N237)? data_i[776] : 
                     (N238)? data_i[808] : 
                     (N239)? data_i[840] : 
                     (N240)? data_i[872] : 
                     (N241)? data_i[904] : 
                     (N242)? data_i[936] : 
                     (N243)? data_i[968] : 
                     (N244)? data_i[1000] : 
                     (N245)? data_i[1032] : 
                     (N246)? data_i[1064] : 
                     (N247)? data_i[1096] : 
                     (N248)? data_i[1128] : 
                     (N249)? data_i[1160] : 
                     (N250)? data_i[1192] : 
                     (N251)? data_i[1224] : 
                     (N252)? data_i[1256] : 
                     (N253)? data_i[1288] : 
                     (N254)? data_i[1320] : 
                     (N255)? data_i[1352] : 
                     (N256)? data_i[1384] : 
                     (N257)? data_i[1416] : 
                     (N258)? data_i[1448] : 
                     (N259)? data_i[1480] : 
                     (N260)? data_i[1512] : 
                     (N261)? data_i[1544] : 
                     (N262)? data_i[1576] : 1'b0;
  assign data_o[7] = (N213)? data_i[7] : 
                     (N214)? data_i[39] : 
                     (N215)? data_i[71] : 
                     (N216)? data_i[103] : 
                     (N217)? data_i[135] : 
                     (N218)? data_i[167] : 
                     (N219)? data_i[199] : 
                     (N220)? data_i[231] : 
                     (N221)? data_i[263] : 
                     (N222)? data_i[295] : 
                     (N223)? data_i[327] : 
                     (N224)? data_i[359] : 
                     (N225)? data_i[391] : 
                     (N226)? data_i[423] : 
                     (N227)? data_i[455] : 
                     (N228)? data_i[487] : 
                     (N229)? data_i[519] : 
                     (N230)? data_i[551] : 
                     (N231)? data_i[583] : 
                     (N232)? data_i[615] : 
                     (N233)? data_i[647] : 
                     (N234)? data_i[679] : 
                     (N235)? data_i[711] : 
                     (N236)? data_i[743] : 
                     (N237)? data_i[775] : 
                     (N238)? data_i[807] : 
                     (N239)? data_i[839] : 
                     (N240)? data_i[871] : 
                     (N241)? data_i[903] : 
                     (N242)? data_i[935] : 
                     (N243)? data_i[967] : 
                     (N244)? data_i[999] : 
                     (N245)? data_i[1031] : 
                     (N246)? data_i[1063] : 
                     (N247)? data_i[1095] : 
                     (N248)? data_i[1127] : 
                     (N249)? data_i[1159] : 
                     (N250)? data_i[1191] : 
                     (N251)? data_i[1223] : 
                     (N252)? data_i[1255] : 
                     (N253)? data_i[1287] : 
                     (N254)? data_i[1319] : 
                     (N255)? data_i[1351] : 
                     (N256)? data_i[1383] : 
                     (N257)? data_i[1415] : 
                     (N258)? data_i[1447] : 
                     (N259)? data_i[1479] : 
                     (N260)? data_i[1511] : 
                     (N261)? data_i[1543] : 
                     (N262)? data_i[1575] : 1'b0;
  assign data_o[6] = (N213)? data_i[6] : 
                     (N214)? data_i[38] : 
                     (N215)? data_i[70] : 
                     (N216)? data_i[102] : 
                     (N217)? data_i[134] : 
                     (N218)? data_i[166] : 
                     (N219)? data_i[198] : 
                     (N220)? data_i[230] : 
                     (N221)? data_i[262] : 
                     (N222)? data_i[294] : 
                     (N223)? data_i[326] : 
                     (N224)? data_i[358] : 
                     (N225)? data_i[390] : 
                     (N226)? data_i[422] : 
                     (N227)? data_i[454] : 
                     (N228)? data_i[486] : 
                     (N229)? data_i[518] : 
                     (N230)? data_i[550] : 
                     (N231)? data_i[582] : 
                     (N232)? data_i[614] : 
                     (N233)? data_i[646] : 
                     (N234)? data_i[678] : 
                     (N235)? data_i[710] : 
                     (N236)? data_i[742] : 
                     (N237)? data_i[774] : 
                     (N238)? data_i[806] : 
                     (N239)? data_i[838] : 
                     (N240)? data_i[870] : 
                     (N241)? data_i[902] : 
                     (N242)? data_i[934] : 
                     (N243)? data_i[966] : 
                     (N244)? data_i[998] : 
                     (N245)? data_i[1030] : 
                     (N246)? data_i[1062] : 
                     (N247)? data_i[1094] : 
                     (N248)? data_i[1126] : 
                     (N249)? data_i[1158] : 
                     (N250)? data_i[1190] : 
                     (N251)? data_i[1222] : 
                     (N252)? data_i[1254] : 
                     (N253)? data_i[1286] : 
                     (N254)? data_i[1318] : 
                     (N255)? data_i[1350] : 
                     (N256)? data_i[1382] : 
                     (N257)? data_i[1414] : 
                     (N258)? data_i[1446] : 
                     (N259)? data_i[1478] : 
                     (N260)? data_i[1510] : 
                     (N261)? data_i[1542] : 
                     (N262)? data_i[1574] : 1'b0;
  assign data_o[5] = (N213)? data_i[5] : 
                     (N214)? data_i[37] : 
                     (N215)? data_i[69] : 
                     (N216)? data_i[101] : 
                     (N217)? data_i[133] : 
                     (N218)? data_i[165] : 
                     (N219)? data_i[197] : 
                     (N220)? data_i[229] : 
                     (N221)? data_i[261] : 
                     (N222)? data_i[293] : 
                     (N223)? data_i[325] : 
                     (N224)? data_i[357] : 
                     (N225)? data_i[389] : 
                     (N226)? data_i[421] : 
                     (N227)? data_i[453] : 
                     (N228)? data_i[485] : 
                     (N229)? data_i[517] : 
                     (N230)? data_i[549] : 
                     (N231)? data_i[581] : 
                     (N232)? data_i[613] : 
                     (N233)? data_i[645] : 
                     (N234)? data_i[677] : 
                     (N235)? data_i[709] : 
                     (N236)? data_i[741] : 
                     (N237)? data_i[773] : 
                     (N238)? data_i[805] : 
                     (N239)? data_i[837] : 
                     (N240)? data_i[869] : 
                     (N241)? data_i[901] : 
                     (N242)? data_i[933] : 
                     (N243)? data_i[965] : 
                     (N244)? data_i[997] : 
                     (N245)? data_i[1029] : 
                     (N246)? data_i[1061] : 
                     (N247)? data_i[1093] : 
                     (N248)? data_i[1125] : 
                     (N249)? data_i[1157] : 
                     (N250)? data_i[1189] : 
                     (N251)? data_i[1221] : 
                     (N252)? data_i[1253] : 
                     (N253)? data_i[1285] : 
                     (N254)? data_i[1317] : 
                     (N255)? data_i[1349] : 
                     (N256)? data_i[1381] : 
                     (N257)? data_i[1413] : 
                     (N258)? data_i[1445] : 
                     (N259)? data_i[1477] : 
                     (N260)? data_i[1509] : 
                     (N261)? data_i[1541] : 
                     (N262)? data_i[1573] : 1'b0;
  assign data_o[4] = (N213)? data_i[4] : 
                     (N214)? data_i[36] : 
                     (N215)? data_i[68] : 
                     (N216)? data_i[100] : 
                     (N217)? data_i[132] : 
                     (N218)? data_i[164] : 
                     (N219)? data_i[196] : 
                     (N220)? data_i[228] : 
                     (N221)? data_i[260] : 
                     (N222)? data_i[292] : 
                     (N223)? data_i[324] : 
                     (N224)? data_i[356] : 
                     (N225)? data_i[388] : 
                     (N226)? data_i[420] : 
                     (N227)? data_i[452] : 
                     (N228)? data_i[484] : 
                     (N229)? data_i[516] : 
                     (N230)? data_i[548] : 
                     (N231)? data_i[580] : 
                     (N232)? data_i[612] : 
                     (N233)? data_i[644] : 
                     (N234)? data_i[676] : 
                     (N235)? data_i[708] : 
                     (N236)? data_i[740] : 
                     (N237)? data_i[772] : 
                     (N238)? data_i[804] : 
                     (N239)? data_i[836] : 
                     (N240)? data_i[868] : 
                     (N241)? data_i[900] : 
                     (N242)? data_i[932] : 
                     (N243)? data_i[964] : 
                     (N244)? data_i[996] : 
                     (N245)? data_i[1028] : 
                     (N246)? data_i[1060] : 
                     (N247)? data_i[1092] : 
                     (N248)? data_i[1124] : 
                     (N249)? data_i[1156] : 
                     (N250)? data_i[1188] : 
                     (N251)? data_i[1220] : 
                     (N252)? data_i[1252] : 
                     (N253)? data_i[1284] : 
                     (N254)? data_i[1316] : 
                     (N255)? data_i[1348] : 
                     (N256)? data_i[1380] : 
                     (N257)? data_i[1412] : 
                     (N258)? data_i[1444] : 
                     (N259)? data_i[1476] : 
                     (N260)? data_i[1508] : 
                     (N261)? data_i[1540] : 
                     (N262)? data_i[1572] : 1'b0;
  assign data_o[3] = (N213)? data_i[3] : 
                     (N214)? data_i[35] : 
                     (N215)? data_i[67] : 
                     (N216)? data_i[99] : 
                     (N217)? data_i[131] : 
                     (N218)? data_i[163] : 
                     (N219)? data_i[195] : 
                     (N220)? data_i[227] : 
                     (N221)? data_i[259] : 
                     (N222)? data_i[291] : 
                     (N223)? data_i[323] : 
                     (N224)? data_i[355] : 
                     (N225)? data_i[387] : 
                     (N226)? data_i[419] : 
                     (N227)? data_i[451] : 
                     (N228)? data_i[483] : 
                     (N229)? data_i[515] : 
                     (N230)? data_i[547] : 
                     (N231)? data_i[579] : 
                     (N232)? data_i[611] : 
                     (N233)? data_i[643] : 
                     (N234)? data_i[675] : 
                     (N235)? data_i[707] : 
                     (N236)? data_i[739] : 
                     (N237)? data_i[771] : 
                     (N238)? data_i[803] : 
                     (N239)? data_i[835] : 
                     (N240)? data_i[867] : 
                     (N241)? data_i[899] : 
                     (N242)? data_i[931] : 
                     (N243)? data_i[963] : 
                     (N244)? data_i[995] : 
                     (N245)? data_i[1027] : 
                     (N246)? data_i[1059] : 
                     (N247)? data_i[1091] : 
                     (N248)? data_i[1123] : 
                     (N249)? data_i[1155] : 
                     (N250)? data_i[1187] : 
                     (N251)? data_i[1219] : 
                     (N252)? data_i[1251] : 
                     (N253)? data_i[1283] : 
                     (N254)? data_i[1315] : 
                     (N255)? data_i[1347] : 
                     (N256)? data_i[1379] : 
                     (N257)? data_i[1411] : 
                     (N258)? data_i[1443] : 
                     (N259)? data_i[1475] : 
                     (N260)? data_i[1507] : 
                     (N261)? data_i[1539] : 
                     (N262)? data_i[1571] : 1'b0;
  assign data_o[2] = (N213)? data_i[2] : 
                     (N214)? data_i[34] : 
                     (N215)? data_i[66] : 
                     (N216)? data_i[98] : 
                     (N217)? data_i[130] : 
                     (N218)? data_i[162] : 
                     (N219)? data_i[194] : 
                     (N220)? data_i[226] : 
                     (N221)? data_i[258] : 
                     (N222)? data_i[290] : 
                     (N223)? data_i[322] : 
                     (N224)? data_i[354] : 
                     (N225)? data_i[386] : 
                     (N226)? data_i[418] : 
                     (N227)? data_i[450] : 
                     (N228)? data_i[482] : 
                     (N229)? data_i[514] : 
                     (N230)? data_i[546] : 
                     (N231)? data_i[578] : 
                     (N232)? data_i[610] : 
                     (N233)? data_i[642] : 
                     (N234)? data_i[674] : 
                     (N235)? data_i[706] : 
                     (N236)? data_i[738] : 
                     (N237)? data_i[770] : 
                     (N238)? data_i[802] : 
                     (N239)? data_i[834] : 
                     (N240)? data_i[866] : 
                     (N241)? data_i[898] : 
                     (N242)? data_i[930] : 
                     (N243)? data_i[962] : 
                     (N244)? data_i[994] : 
                     (N245)? data_i[1026] : 
                     (N246)? data_i[1058] : 
                     (N247)? data_i[1090] : 
                     (N248)? data_i[1122] : 
                     (N249)? data_i[1154] : 
                     (N250)? data_i[1186] : 
                     (N251)? data_i[1218] : 
                     (N252)? data_i[1250] : 
                     (N253)? data_i[1282] : 
                     (N254)? data_i[1314] : 
                     (N255)? data_i[1346] : 
                     (N256)? data_i[1378] : 
                     (N257)? data_i[1410] : 
                     (N258)? data_i[1442] : 
                     (N259)? data_i[1474] : 
                     (N260)? data_i[1506] : 
                     (N261)? data_i[1538] : 
                     (N262)? data_i[1570] : 1'b0;
  assign data_o[1] = (N213)? data_i[1] : 
                     (N214)? data_i[33] : 
                     (N215)? data_i[65] : 
                     (N216)? data_i[97] : 
                     (N217)? data_i[129] : 
                     (N218)? data_i[161] : 
                     (N219)? data_i[193] : 
                     (N220)? data_i[225] : 
                     (N221)? data_i[257] : 
                     (N222)? data_i[289] : 
                     (N223)? data_i[321] : 
                     (N224)? data_i[353] : 
                     (N225)? data_i[385] : 
                     (N226)? data_i[417] : 
                     (N227)? data_i[449] : 
                     (N228)? data_i[481] : 
                     (N229)? data_i[513] : 
                     (N230)? data_i[545] : 
                     (N231)? data_i[577] : 
                     (N232)? data_i[609] : 
                     (N233)? data_i[641] : 
                     (N234)? data_i[673] : 
                     (N235)? data_i[705] : 
                     (N236)? data_i[737] : 
                     (N237)? data_i[769] : 
                     (N238)? data_i[801] : 
                     (N239)? data_i[833] : 
                     (N240)? data_i[865] : 
                     (N241)? data_i[897] : 
                     (N242)? data_i[929] : 
                     (N243)? data_i[961] : 
                     (N244)? data_i[993] : 
                     (N245)? data_i[1025] : 
                     (N246)? data_i[1057] : 
                     (N247)? data_i[1089] : 
                     (N248)? data_i[1121] : 
                     (N249)? data_i[1153] : 
                     (N250)? data_i[1185] : 
                     (N251)? data_i[1217] : 
                     (N252)? data_i[1249] : 
                     (N253)? data_i[1281] : 
                     (N254)? data_i[1313] : 
                     (N255)? data_i[1345] : 
                     (N256)? data_i[1377] : 
                     (N257)? data_i[1409] : 
                     (N258)? data_i[1441] : 
                     (N259)? data_i[1473] : 
                     (N260)? data_i[1505] : 
                     (N261)? data_i[1537] : 
                     (N262)? data_i[1569] : 1'b0;
  assign data_o[0] = (N213)? data_i[0] : 
                     (N214)? data_i[32] : 
                     (N215)? data_i[64] : 
                     (N216)? data_i[96] : 
                     (N217)? data_i[128] : 
                     (N218)? data_i[160] : 
                     (N219)? data_i[192] : 
                     (N220)? data_i[224] : 
                     (N221)? data_i[256] : 
                     (N222)? data_i[288] : 
                     (N223)? data_i[320] : 
                     (N224)? data_i[352] : 
                     (N225)? data_i[384] : 
                     (N226)? data_i[416] : 
                     (N227)? data_i[448] : 
                     (N228)? data_i[480] : 
                     (N229)? data_i[512] : 
                     (N230)? data_i[544] : 
                     (N231)? data_i[576] : 
                     (N232)? data_i[608] : 
                     (N233)? data_i[640] : 
                     (N234)? data_i[672] : 
                     (N235)? data_i[704] : 
                     (N236)? data_i[736] : 
                     (N237)? data_i[768] : 
                     (N238)? data_i[800] : 
                     (N239)? data_i[832] : 
                     (N240)? data_i[864] : 
                     (N241)? data_i[896] : 
                     (N242)? data_i[928] : 
                     (N243)? data_i[960] : 
                     (N244)? data_i[992] : 
                     (N245)? data_i[1024] : 
                     (N246)? data_i[1056] : 
                     (N247)? data_i[1088] : 
                     (N248)? data_i[1120] : 
                     (N249)? data_i[1152] : 
                     (N250)? data_i[1184] : 
                     (N251)? data_i[1216] : 
                     (N252)? data_i[1248] : 
                     (N253)? data_i[1280] : 
                     (N254)? data_i[1312] : 
                     (N255)? data_i[1344] : 
                     (N256)? data_i[1376] : 
                     (N257)? data_i[1408] : 
                     (N258)? data_i[1440] : 
                     (N259)? data_i[1472] : 
                     (N260)? data_i[1504] : 
                     (N261)? data_i[1536] : 
                     (N262)? data_i[1568] : 1'b0;

endmodule



module bsg_parallel_in_serial_out_dynamic
(
  clk_i,
  reset_i,
  v_i,
  len_i,
  data_i,
  ready_o,
  v_o,
  len_v_o,
  data_o,
  yumi_i
);

  input [5:0] len_i;
  input [1599:0] data_i;
  output [31:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  output len_v_o;
  wire [31:0] data_o;
  wire ready_o,v_o,len_v_o,count_r_is_last,up_li,clear_li,N0,N1,N2,N3,N4,N6;
  wire [5:0] len_lo,count_lo;
  wire [1599:0] fifo_data_lo;

  bsg_two_fifo_width_p6
  go_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(ready_o),
    .data_i(len_i),
    .v_i(v_i),
    .v_o(v_o),
    .data_o(len_lo),
    .yumi_i(clear_li)
  );


  bsg_two_fifo_width_p1600
  data_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(v_i),
    .data_o(fifo_data_lo),
    .yumi_i(clear_li)
  );

  assign count_r_is_last = count_lo == len_lo;

  bsg_counter_clear_up_max_val_p49_init_val_p0
  ctr
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .clear_i(clear_li),
    .up_i(up_li),
    .count_o(count_lo)
  );


  bsg_mux_width_p32_els_p50
  data_mux
  (
    .data_i(fifo_data_lo),
    .sel_i(count_lo),
    .data_o(data_o)
  );

  assign N0 = count_lo[4] | count_lo[5];
  assign N1 = count_lo[3] | N0;
  assign N2 = count_lo[2] | N1;
  assign N3 = count_lo[1] | N2;
  assign N4 = count_lo[0] | N3;
  assign len_v_o = ~N4;
  assign up_li = yumi_i & N6;
  assign N6 = ~count_r_is_last;
  assign clear_li = yumi_i & count_r_is_last;

endmodule

