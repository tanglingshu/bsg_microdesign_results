

module bsg_mem_1r1w_sync_synth_width_p16_els_p512_read_write_same_addr_p0_harden_p0
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [8:0] w_addr_i;
  input [15:0] w_data_i;
  input [8:0] r_addr_i;
  output [15:0] r_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r_v_i;
  wire [15:0] r_data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144;
  reg [8:0] r_addr_r;
  reg [8191:0] mem;
  assign r_data_o[15] = (N535)? mem[15] : 
                        (N537)? mem[31] : 
                        (N539)? mem[47] : 
                        (N541)? mem[63] : 
                        (N543)? mem[79] : 
                        (N545)? mem[95] : 
                        (N547)? mem[111] : 
                        (N549)? mem[127] : 
                        (N551)? mem[143] : 
                        (N553)? mem[159] : 
                        (N555)? mem[175] : 
                        (N557)? mem[191] : 
                        (N559)? mem[207] : 
                        (N561)? mem[223] : 
                        (N563)? mem[239] : 
                        (N565)? mem[255] : 
                        (N567)? mem[271] : 
                        (N569)? mem[287] : 
                        (N571)? mem[303] : 
                        (N573)? mem[319] : 
                        (N575)? mem[335] : 
                        (N577)? mem[351] : 
                        (N579)? mem[367] : 
                        (N581)? mem[383] : 
                        (N583)? mem[399] : 
                        (N585)? mem[415] : 
                        (N587)? mem[431] : 
                        (N589)? mem[447] : 
                        (N591)? mem[463] : 
                        (N593)? mem[479] : 
                        (N595)? mem[495] : 
                        (N597)? mem[511] : 
                        (N599)? mem[527] : 
                        (N601)? mem[543] : 
                        (N603)? mem[559] : 
                        (N605)? mem[575] : 
                        (N607)? mem[591] : 
                        (N609)? mem[607] : 
                        (N611)? mem[623] : 
                        (N613)? mem[639] : 
                        (N615)? mem[655] : 
                        (N617)? mem[671] : 
                        (N619)? mem[687] : 
                        (N621)? mem[703] : 
                        (N623)? mem[719] : 
                        (N625)? mem[735] : 
                        (N627)? mem[751] : 
                        (N629)? mem[767] : 
                        (N631)? mem[783] : 
                        (N633)? mem[799] : 
                        (N635)? mem[815] : 
                        (N637)? mem[831] : 
                        (N639)? mem[847] : 
                        (N641)? mem[863] : 
                        (N643)? mem[879] : 
                        (N645)? mem[895] : 
                        (N647)? mem[911] : 
                        (N649)? mem[927] : 
                        (N651)? mem[943] : 
                        (N653)? mem[959] : 
                        (N655)? mem[975] : 
                        (N657)? mem[991] : 
                        (N659)? mem[1007] : 
                        (N661)? mem[1023] : 
                        (N663)? mem[1039] : 
                        (N665)? mem[1055] : 
                        (N667)? mem[1071] : 
                        (N669)? mem[1087] : 
                        (N671)? mem[1103] : 
                        (N673)? mem[1119] : 
                        (N675)? mem[1135] : 
                        (N677)? mem[1151] : 
                        (N679)? mem[1167] : 
                        (N681)? mem[1183] : 
                        (N683)? mem[1199] : 
                        (N685)? mem[1215] : 
                        (N687)? mem[1231] : 
                        (N689)? mem[1247] : 
                        (N691)? mem[1263] : 
                        (N693)? mem[1279] : 
                        (N695)? mem[1295] : 
                        (N697)? mem[1311] : 
                        (N699)? mem[1327] : 
                        (N701)? mem[1343] : 
                        (N703)? mem[1359] : 
                        (N705)? mem[1375] : 
                        (N707)? mem[1391] : 
                        (N709)? mem[1407] : 
                        (N711)? mem[1423] : 
                        (N713)? mem[1439] : 
                        (N715)? mem[1455] : 
                        (N717)? mem[1471] : 
                        (N719)? mem[1487] : 
                        (N721)? mem[1503] : 
                        (N723)? mem[1519] : 
                        (N725)? mem[1535] : 
                        (N727)? mem[1551] : 
                        (N729)? mem[1567] : 
                        (N731)? mem[1583] : 
                        (N733)? mem[1599] : 
                        (N735)? mem[1615] : 
                        (N737)? mem[1631] : 
                        (N739)? mem[1647] : 
                        (N741)? mem[1663] : 
                        (N743)? mem[1679] : 
                        (N745)? mem[1695] : 
                        (N747)? mem[1711] : 
                        (N749)? mem[1727] : 
                        (N751)? mem[1743] : 
                        (N753)? mem[1759] : 
                        (N755)? mem[1775] : 
                        (N757)? mem[1791] : 
                        (N759)? mem[1807] : 
                        (N761)? mem[1823] : 
                        (N763)? mem[1839] : 
                        (N765)? mem[1855] : 
                        (N767)? mem[1871] : 
                        (N769)? mem[1887] : 
                        (N771)? mem[1903] : 
                        (N773)? mem[1919] : 
                        (N775)? mem[1935] : 
                        (N777)? mem[1951] : 
                        (N779)? mem[1967] : 
                        (N781)? mem[1983] : 
                        (N783)? mem[1999] : 
                        (N785)? mem[2015] : 
                        (N787)? mem[2031] : 
                        (N789)? mem[2047] : 
                        (N791)? mem[2063] : 
                        (N793)? mem[2079] : 
                        (N795)? mem[2095] : 
                        (N797)? mem[2111] : 
                        (N799)? mem[2127] : 
                        (N801)? mem[2143] : 
                        (N803)? mem[2159] : 
                        (N805)? mem[2175] : 
                        (N807)? mem[2191] : 
                        (N809)? mem[2207] : 
                        (N811)? mem[2223] : 
                        (N813)? mem[2239] : 
                        (N815)? mem[2255] : 
                        (N817)? mem[2271] : 
                        (N819)? mem[2287] : 
                        (N821)? mem[2303] : 
                        (N823)? mem[2319] : 
                        (N825)? mem[2335] : 
                        (N827)? mem[2351] : 
                        (N829)? mem[2367] : 
                        (N831)? mem[2383] : 
                        (N833)? mem[2399] : 
                        (N835)? mem[2415] : 
                        (N837)? mem[2431] : 
                        (N839)? mem[2447] : 
                        (N841)? mem[2463] : 
                        (N843)? mem[2479] : 
                        (N845)? mem[2495] : 
                        (N847)? mem[2511] : 
                        (N849)? mem[2527] : 
                        (N851)? mem[2543] : 
                        (N853)? mem[2559] : 
                        (N855)? mem[2575] : 
                        (N857)? mem[2591] : 
                        (N859)? mem[2607] : 
                        (N861)? mem[2623] : 
                        (N863)? mem[2639] : 
                        (N865)? mem[2655] : 
                        (N867)? mem[2671] : 
                        (N869)? mem[2687] : 
                        (N871)? mem[2703] : 
                        (N873)? mem[2719] : 
                        (N875)? mem[2735] : 
                        (N877)? mem[2751] : 
                        (N879)? mem[2767] : 
                        (N881)? mem[2783] : 
                        (N883)? mem[2799] : 
                        (N885)? mem[2815] : 
                        (N887)? mem[2831] : 
                        (N889)? mem[2847] : 
                        (N891)? mem[2863] : 
                        (N893)? mem[2879] : 
                        (N895)? mem[2895] : 
                        (N897)? mem[2911] : 
                        (N899)? mem[2927] : 
                        (N901)? mem[2943] : 
                        (N903)? mem[2959] : 
                        (N905)? mem[2975] : 
                        (N907)? mem[2991] : 
                        (N909)? mem[3007] : 
                        (N911)? mem[3023] : 
                        (N913)? mem[3039] : 
                        (N915)? mem[3055] : 
                        (N917)? mem[3071] : 
                        (N919)? mem[3087] : 
                        (N921)? mem[3103] : 
                        (N923)? mem[3119] : 
                        (N925)? mem[3135] : 
                        (N927)? mem[3151] : 
                        (N929)? mem[3167] : 
                        (N931)? mem[3183] : 
                        (N933)? mem[3199] : 
                        (N935)? mem[3215] : 
                        (N937)? mem[3231] : 
                        (N939)? mem[3247] : 
                        (N941)? mem[3263] : 
                        (N943)? mem[3279] : 
                        (N945)? mem[3295] : 
                        (N947)? mem[3311] : 
                        (N949)? mem[3327] : 
                        (N951)? mem[3343] : 
                        (N953)? mem[3359] : 
                        (N955)? mem[3375] : 
                        (N957)? mem[3391] : 
                        (N959)? mem[3407] : 
                        (N961)? mem[3423] : 
                        (N963)? mem[3439] : 
                        (N965)? mem[3455] : 
                        (N967)? mem[3471] : 
                        (N969)? mem[3487] : 
                        (N971)? mem[3503] : 
                        (N973)? mem[3519] : 
                        (N975)? mem[3535] : 
                        (N977)? mem[3551] : 
                        (N979)? mem[3567] : 
                        (N981)? mem[3583] : 
                        (N983)? mem[3599] : 
                        (N985)? mem[3615] : 
                        (N987)? mem[3631] : 
                        (N989)? mem[3647] : 
                        (N991)? mem[3663] : 
                        (N993)? mem[3679] : 
                        (N995)? mem[3695] : 
                        (N997)? mem[3711] : 
                        (N999)? mem[3727] : 
                        (N1001)? mem[3743] : 
                        (N1003)? mem[3759] : 
                        (N1005)? mem[3775] : 
                        (N1007)? mem[3791] : 
                        (N1009)? mem[3807] : 
                        (N1011)? mem[3823] : 
                        (N1013)? mem[3839] : 
                        (N1015)? mem[3855] : 
                        (N1017)? mem[3871] : 
                        (N1019)? mem[3887] : 
                        (N1021)? mem[3903] : 
                        (N1023)? mem[3919] : 
                        (N1025)? mem[3935] : 
                        (N1027)? mem[3951] : 
                        (N1029)? mem[3967] : 
                        (N1031)? mem[3983] : 
                        (N1033)? mem[3999] : 
                        (N1035)? mem[4015] : 
                        (N1037)? mem[4031] : 
                        (N1039)? mem[4047] : 
                        (N1041)? mem[4063] : 
                        (N1043)? mem[4079] : 
                        (N1045)? mem[4095] : 
                        (N536)? mem[4111] : 
                        (N538)? mem[4127] : 
                        (N540)? mem[4143] : 
                        (N542)? mem[4159] : 
                        (N544)? mem[4175] : 
                        (N546)? mem[4191] : 
                        (N548)? mem[4207] : 
                        (N550)? mem[4223] : 
                        (N552)? mem[4239] : 
                        (N554)? mem[4255] : 
                        (N556)? mem[4271] : 
                        (N558)? mem[4287] : 
                        (N560)? mem[4303] : 
                        (N562)? mem[4319] : 
                        (N564)? mem[4335] : 
                        (N566)? mem[4351] : 
                        (N568)? mem[4367] : 
                        (N570)? mem[4383] : 
                        (N572)? mem[4399] : 
                        (N574)? mem[4415] : 
                        (N576)? mem[4431] : 
                        (N578)? mem[4447] : 
                        (N580)? mem[4463] : 
                        (N582)? mem[4479] : 
                        (N584)? mem[4495] : 
                        (N586)? mem[4511] : 
                        (N588)? mem[4527] : 
                        (N590)? mem[4543] : 
                        (N592)? mem[4559] : 
                        (N594)? mem[4575] : 
                        (N596)? mem[4591] : 
                        (N598)? mem[4607] : 
                        (N600)? mem[4623] : 
                        (N602)? mem[4639] : 
                        (N604)? mem[4655] : 
                        (N606)? mem[4671] : 
                        (N608)? mem[4687] : 
                        (N610)? mem[4703] : 
                        (N612)? mem[4719] : 
                        (N614)? mem[4735] : 
                        (N616)? mem[4751] : 
                        (N618)? mem[4767] : 
                        (N620)? mem[4783] : 
                        (N622)? mem[4799] : 
                        (N624)? mem[4815] : 
                        (N626)? mem[4831] : 
                        (N628)? mem[4847] : 
                        (N630)? mem[4863] : 
                        (N632)? mem[4879] : 
                        (N634)? mem[4895] : 
                        (N636)? mem[4911] : 
                        (N638)? mem[4927] : 
                        (N640)? mem[4943] : 
                        (N642)? mem[4959] : 
                        (N644)? mem[4975] : 
                        (N646)? mem[4991] : 
                        (N648)? mem[5007] : 
                        (N650)? mem[5023] : 
                        (N652)? mem[5039] : 
                        (N654)? mem[5055] : 
                        (N656)? mem[5071] : 
                        (N658)? mem[5087] : 
                        (N660)? mem[5103] : 
                        (N662)? mem[5119] : 
                        (N664)? mem[5135] : 
                        (N666)? mem[5151] : 
                        (N668)? mem[5167] : 
                        (N670)? mem[5183] : 
                        (N672)? mem[5199] : 
                        (N674)? mem[5215] : 
                        (N676)? mem[5231] : 
                        (N678)? mem[5247] : 
                        (N680)? mem[5263] : 
                        (N682)? mem[5279] : 
                        (N684)? mem[5295] : 
                        (N686)? mem[5311] : 
                        (N688)? mem[5327] : 
                        (N690)? mem[5343] : 
                        (N692)? mem[5359] : 
                        (N694)? mem[5375] : 
                        (N696)? mem[5391] : 
                        (N698)? mem[5407] : 
                        (N700)? mem[5423] : 
                        (N702)? mem[5439] : 
                        (N704)? mem[5455] : 
                        (N706)? mem[5471] : 
                        (N708)? mem[5487] : 
                        (N710)? mem[5503] : 
                        (N712)? mem[5519] : 
                        (N714)? mem[5535] : 
                        (N716)? mem[5551] : 
                        (N718)? mem[5567] : 
                        (N720)? mem[5583] : 
                        (N722)? mem[5599] : 
                        (N724)? mem[5615] : 
                        (N726)? mem[5631] : 
                        (N728)? mem[5647] : 
                        (N730)? mem[5663] : 
                        (N732)? mem[5679] : 
                        (N734)? mem[5695] : 
                        (N736)? mem[5711] : 
                        (N738)? mem[5727] : 
                        (N740)? mem[5743] : 
                        (N742)? mem[5759] : 
                        (N744)? mem[5775] : 
                        (N746)? mem[5791] : 
                        (N748)? mem[5807] : 
                        (N750)? mem[5823] : 
                        (N752)? mem[5839] : 
                        (N754)? mem[5855] : 
                        (N756)? mem[5871] : 
                        (N758)? mem[5887] : 
                        (N760)? mem[5903] : 
                        (N762)? mem[5919] : 
                        (N764)? mem[5935] : 
                        (N766)? mem[5951] : 
                        (N768)? mem[5967] : 
                        (N770)? mem[5983] : 
                        (N772)? mem[5999] : 
                        (N774)? mem[6015] : 
                        (N776)? mem[6031] : 
                        (N778)? mem[6047] : 
                        (N780)? mem[6063] : 
                        (N782)? mem[6079] : 
                        (N784)? mem[6095] : 
                        (N786)? mem[6111] : 
                        (N788)? mem[6127] : 
                        (N790)? mem[6143] : 
                        (N792)? mem[6159] : 
                        (N794)? mem[6175] : 
                        (N796)? mem[6191] : 
                        (N798)? mem[6207] : 
                        (N800)? mem[6223] : 
                        (N802)? mem[6239] : 
                        (N804)? mem[6255] : 
                        (N806)? mem[6271] : 
                        (N808)? mem[6287] : 
                        (N810)? mem[6303] : 
                        (N812)? mem[6319] : 
                        (N814)? mem[6335] : 
                        (N816)? mem[6351] : 
                        (N818)? mem[6367] : 
                        (N820)? mem[6383] : 
                        (N822)? mem[6399] : 
                        (N824)? mem[6415] : 
                        (N826)? mem[6431] : 
                        (N828)? mem[6447] : 
                        (N830)? mem[6463] : 
                        (N832)? mem[6479] : 
                        (N834)? mem[6495] : 
                        (N836)? mem[6511] : 
                        (N838)? mem[6527] : 
                        (N840)? mem[6543] : 
                        (N842)? mem[6559] : 
                        (N844)? mem[6575] : 
                        (N846)? mem[6591] : 
                        (N848)? mem[6607] : 
                        (N850)? mem[6623] : 
                        (N852)? mem[6639] : 
                        (N854)? mem[6655] : 
                        (N856)? mem[6671] : 
                        (N858)? mem[6687] : 
                        (N860)? mem[6703] : 
                        (N862)? mem[6719] : 
                        (N864)? mem[6735] : 
                        (N866)? mem[6751] : 
                        (N868)? mem[6767] : 
                        (N870)? mem[6783] : 
                        (N872)? mem[6799] : 
                        (N874)? mem[6815] : 
                        (N876)? mem[6831] : 
                        (N878)? mem[6847] : 
                        (N880)? mem[6863] : 
                        (N882)? mem[6879] : 
                        (N884)? mem[6895] : 
                        (N886)? mem[6911] : 
                        (N888)? mem[6927] : 
                        (N890)? mem[6943] : 
                        (N892)? mem[6959] : 
                        (N894)? mem[6975] : 
                        (N896)? mem[6991] : 
                        (N898)? mem[7007] : 
                        (N900)? mem[7023] : 
                        (N902)? mem[7039] : 
                        (N904)? mem[7055] : 
                        (N906)? mem[7071] : 
                        (N908)? mem[7087] : 
                        (N910)? mem[7103] : 
                        (N912)? mem[7119] : 
                        (N914)? mem[7135] : 
                        (N916)? mem[7151] : 
                        (N918)? mem[7167] : 
                        (N920)? mem[7183] : 
                        (N922)? mem[7199] : 
                        (N924)? mem[7215] : 
                        (N926)? mem[7231] : 
                        (N928)? mem[7247] : 
                        (N930)? mem[7263] : 
                        (N932)? mem[7279] : 
                        (N934)? mem[7295] : 
                        (N936)? mem[7311] : 
                        (N938)? mem[7327] : 
                        (N940)? mem[7343] : 
                        (N942)? mem[7359] : 
                        (N944)? mem[7375] : 
                        (N946)? mem[7391] : 
                        (N948)? mem[7407] : 
                        (N950)? mem[7423] : 
                        (N952)? mem[7439] : 
                        (N954)? mem[7455] : 
                        (N956)? mem[7471] : 
                        (N958)? mem[7487] : 
                        (N960)? mem[7503] : 
                        (N962)? mem[7519] : 
                        (N964)? mem[7535] : 
                        (N966)? mem[7551] : 
                        (N968)? mem[7567] : 
                        (N970)? mem[7583] : 
                        (N972)? mem[7599] : 
                        (N974)? mem[7615] : 
                        (N976)? mem[7631] : 
                        (N978)? mem[7647] : 
                        (N980)? mem[7663] : 
                        (N982)? mem[7679] : 
                        (N984)? mem[7695] : 
                        (N986)? mem[7711] : 
                        (N988)? mem[7727] : 
                        (N990)? mem[7743] : 
                        (N992)? mem[7759] : 
                        (N994)? mem[7775] : 
                        (N996)? mem[7791] : 
                        (N998)? mem[7807] : 
                        (N1000)? mem[7823] : 
                        (N1002)? mem[7839] : 
                        (N1004)? mem[7855] : 
                        (N1006)? mem[7871] : 
                        (N1008)? mem[7887] : 
                        (N1010)? mem[7903] : 
                        (N1012)? mem[7919] : 
                        (N1014)? mem[7935] : 
                        (N1016)? mem[7951] : 
                        (N1018)? mem[7967] : 
                        (N1020)? mem[7983] : 
                        (N1022)? mem[7999] : 
                        (N1024)? mem[8015] : 
                        (N1026)? mem[8031] : 
                        (N1028)? mem[8047] : 
                        (N1030)? mem[8063] : 
                        (N1032)? mem[8079] : 
                        (N1034)? mem[8095] : 
                        (N1036)? mem[8111] : 
                        (N1038)? mem[8127] : 
                        (N1040)? mem[8143] : 
                        (N1042)? mem[8159] : 
                        (N1044)? mem[8175] : 
                        (N1046)? mem[8191] : 1'b0;
  assign r_data_o[14] = (N535)? mem[14] : 
                        (N537)? mem[30] : 
                        (N539)? mem[46] : 
                        (N541)? mem[62] : 
                        (N543)? mem[78] : 
                        (N545)? mem[94] : 
                        (N547)? mem[110] : 
                        (N549)? mem[126] : 
                        (N551)? mem[142] : 
                        (N553)? mem[158] : 
                        (N555)? mem[174] : 
                        (N557)? mem[190] : 
                        (N559)? mem[206] : 
                        (N561)? mem[222] : 
                        (N563)? mem[238] : 
                        (N565)? mem[254] : 
                        (N567)? mem[270] : 
                        (N569)? mem[286] : 
                        (N571)? mem[302] : 
                        (N573)? mem[318] : 
                        (N575)? mem[334] : 
                        (N577)? mem[350] : 
                        (N579)? mem[366] : 
                        (N581)? mem[382] : 
                        (N583)? mem[398] : 
                        (N585)? mem[414] : 
                        (N587)? mem[430] : 
                        (N589)? mem[446] : 
                        (N591)? mem[462] : 
                        (N593)? mem[478] : 
                        (N595)? mem[494] : 
                        (N597)? mem[510] : 
                        (N599)? mem[526] : 
                        (N601)? mem[542] : 
                        (N603)? mem[558] : 
                        (N605)? mem[574] : 
                        (N607)? mem[590] : 
                        (N609)? mem[606] : 
                        (N611)? mem[622] : 
                        (N613)? mem[638] : 
                        (N615)? mem[654] : 
                        (N617)? mem[670] : 
                        (N619)? mem[686] : 
                        (N621)? mem[702] : 
                        (N623)? mem[718] : 
                        (N625)? mem[734] : 
                        (N627)? mem[750] : 
                        (N629)? mem[766] : 
                        (N631)? mem[782] : 
                        (N633)? mem[798] : 
                        (N635)? mem[814] : 
                        (N637)? mem[830] : 
                        (N639)? mem[846] : 
                        (N641)? mem[862] : 
                        (N643)? mem[878] : 
                        (N645)? mem[894] : 
                        (N647)? mem[910] : 
                        (N649)? mem[926] : 
                        (N651)? mem[942] : 
                        (N653)? mem[958] : 
                        (N655)? mem[974] : 
                        (N657)? mem[990] : 
                        (N659)? mem[1006] : 
                        (N661)? mem[1022] : 
                        (N663)? mem[1038] : 
                        (N665)? mem[1054] : 
                        (N667)? mem[1070] : 
                        (N669)? mem[1086] : 
                        (N671)? mem[1102] : 
                        (N673)? mem[1118] : 
                        (N675)? mem[1134] : 
                        (N677)? mem[1150] : 
                        (N679)? mem[1166] : 
                        (N681)? mem[1182] : 
                        (N683)? mem[1198] : 
                        (N685)? mem[1214] : 
                        (N687)? mem[1230] : 
                        (N689)? mem[1246] : 
                        (N691)? mem[1262] : 
                        (N693)? mem[1278] : 
                        (N695)? mem[1294] : 
                        (N697)? mem[1310] : 
                        (N699)? mem[1326] : 
                        (N701)? mem[1342] : 
                        (N703)? mem[1358] : 
                        (N705)? mem[1374] : 
                        (N707)? mem[1390] : 
                        (N709)? mem[1406] : 
                        (N711)? mem[1422] : 
                        (N713)? mem[1438] : 
                        (N715)? mem[1454] : 
                        (N717)? mem[1470] : 
                        (N719)? mem[1486] : 
                        (N721)? mem[1502] : 
                        (N723)? mem[1518] : 
                        (N725)? mem[1534] : 
                        (N727)? mem[1550] : 
                        (N729)? mem[1566] : 
                        (N731)? mem[1582] : 
                        (N733)? mem[1598] : 
                        (N735)? mem[1614] : 
                        (N737)? mem[1630] : 
                        (N739)? mem[1646] : 
                        (N741)? mem[1662] : 
                        (N743)? mem[1678] : 
                        (N745)? mem[1694] : 
                        (N747)? mem[1710] : 
                        (N749)? mem[1726] : 
                        (N751)? mem[1742] : 
                        (N753)? mem[1758] : 
                        (N755)? mem[1774] : 
                        (N757)? mem[1790] : 
                        (N759)? mem[1806] : 
                        (N761)? mem[1822] : 
                        (N763)? mem[1838] : 
                        (N765)? mem[1854] : 
                        (N767)? mem[1870] : 
                        (N769)? mem[1886] : 
                        (N771)? mem[1902] : 
                        (N773)? mem[1918] : 
                        (N775)? mem[1934] : 
                        (N777)? mem[1950] : 
                        (N779)? mem[1966] : 
                        (N781)? mem[1982] : 
                        (N783)? mem[1998] : 
                        (N785)? mem[2014] : 
                        (N787)? mem[2030] : 
                        (N789)? mem[2046] : 
                        (N791)? mem[2062] : 
                        (N793)? mem[2078] : 
                        (N795)? mem[2094] : 
                        (N797)? mem[2110] : 
                        (N799)? mem[2126] : 
                        (N801)? mem[2142] : 
                        (N803)? mem[2158] : 
                        (N805)? mem[2174] : 
                        (N807)? mem[2190] : 
                        (N809)? mem[2206] : 
                        (N811)? mem[2222] : 
                        (N813)? mem[2238] : 
                        (N815)? mem[2254] : 
                        (N817)? mem[2270] : 
                        (N819)? mem[2286] : 
                        (N821)? mem[2302] : 
                        (N823)? mem[2318] : 
                        (N825)? mem[2334] : 
                        (N827)? mem[2350] : 
                        (N829)? mem[2366] : 
                        (N831)? mem[2382] : 
                        (N833)? mem[2398] : 
                        (N835)? mem[2414] : 
                        (N837)? mem[2430] : 
                        (N839)? mem[2446] : 
                        (N841)? mem[2462] : 
                        (N843)? mem[2478] : 
                        (N845)? mem[2494] : 
                        (N847)? mem[2510] : 
                        (N849)? mem[2526] : 
                        (N851)? mem[2542] : 
                        (N853)? mem[2558] : 
                        (N855)? mem[2574] : 
                        (N857)? mem[2590] : 
                        (N859)? mem[2606] : 
                        (N861)? mem[2622] : 
                        (N863)? mem[2638] : 
                        (N865)? mem[2654] : 
                        (N867)? mem[2670] : 
                        (N869)? mem[2686] : 
                        (N871)? mem[2702] : 
                        (N873)? mem[2718] : 
                        (N875)? mem[2734] : 
                        (N877)? mem[2750] : 
                        (N879)? mem[2766] : 
                        (N881)? mem[2782] : 
                        (N883)? mem[2798] : 
                        (N885)? mem[2814] : 
                        (N887)? mem[2830] : 
                        (N889)? mem[2846] : 
                        (N891)? mem[2862] : 
                        (N893)? mem[2878] : 
                        (N895)? mem[2894] : 
                        (N897)? mem[2910] : 
                        (N899)? mem[2926] : 
                        (N901)? mem[2942] : 
                        (N903)? mem[2958] : 
                        (N905)? mem[2974] : 
                        (N907)? mem[2990] : 
                        (N909)? mem[3006] : 
                        (N911)? mem[3022] : 
                        (N913)? mem[3038] : 
                        (N915)? mem[3054] : 
                        (N917)? mem[3070] : 
                        (N919)? mem[3086] : 
                        (N921)? mem[3102] : 
                        (N923)? mem[3118] : 
                        (N925)? mem[3134] : 
                        (N927)? mem[3150] : 
                        (N929)? mem[3166] : 
                        (N931)? mem[3182] : 
                        (N933)? mem[3198] : 
                        (N935)? mem[3214] : 
                        (N937)? mem[3230] : 
                        (N939)? mem[3246] : 
                        (N941)? mem[3262] : 
                        (N943)? mem[3278] : 
                        (N945)? mem[3294] : 
                        (N947)? mem[3310] : 
                        (N949)? mem[3326] : 
                        (N951)? mem[3342] : 
                        (N953)? mem[3358] : 
                        (N955)? mem[3374] : 
                        (N957)? mem[3390] : 
                        (N959)? mem[3406] : 
                        (N961)? mem[3422] : 
                        (N963)? mem[3438] : 
                        (N965)? mem[3454] : 
                        (N967)? mem[3470] : 
                        (N969)? mem[3486] : 
                        (N971)? mem[3502] : 
                        (N973)? mem[3518] : 
                        (N975)? mem[3534] : 
                        (N977)? mem[3550] : 
                        (N979)? mem[3566] : 
                        (N981)? mem[3582] : 
                        (N983)? mem[3598] : 
                        (N985)? mem[3614] : 
                        (N987)? mem[3630] : 
                        (N989)? mem[3646] : 
                        (N991)? mem[3662] : 
                        (N993)? mem[3678] : 
                        (N995)? mem[3694] : 
                        (N997)? mem[3710] : 
                        (N999)? mem[3726] : 
                        (N1001)? mem[3742] : 
                        (N1003)? mem[3758] : 
                        (N1005)? mem[3774] : 
                        (N1007)? mem[3790] : 
                        (N1009)? mem[3806] : 
                        (N1011)? mem[3822] : 
                        (N1013)? mem[3838] : 
                        (N1015)? mem[3854] : 
                        (N1017)? mem[3870] : 
                        (N1019)? mem[3886] : 
                        (N1021)? mem[3902] : 
                        (N1023)? mem[3918] : 
                        (N1025)? mem[3934] : 
                        (N1027)? mem[3950] : 
                        (N1029)? mem[3966] : 
                        (N1031)? mem[3982] : 
                        (N1033)? mem[3998] : 
                        (N1035)? mem[4014] : 
                        (N1037)? mem[4030] : 
                        (N1039)? mem[4046] : 
                        (N1041)? mem[4062] : 
                        (N1043)? mem[4078] : 
                        (N1045)? mem[4094] : 
                        (N536)? mem[4110] : 
                        (N538)? mem[4126] : 
                        (N540)? mem[4142] : 
                        (N542)? mem[4158] : 
                        (N544)? mem[4174] : 
                        (N546)? mem[4190] : 
                        (N548)? mem[4206] : 
                        (N550)? mem[4222] : 
                        (N552)? mem[4238] : 
                        (N554)? mem[4254] : 
                        (N556)? mem[4270] : 
                        (N558)? mem[4286] : 
                        (N560)? mem[4302] : 
                        (N562)? mem[4318] : 
                        (N564)? mem[4334] : 
                        (N566)? mem[4350] : 
                        (N568)? mem[4366] : 
                        (N570)? mem[4382] : 
                        (N572)? mem[4398] : 
                        (N574)? mem[4414] : 
                        (N576)? mem[4430] : 
                        (N578)? mem[4446] : 
                        (N580)? mem[4462] : 
                        (N582)? mem[4478] : 
                        (N584)? mem[4494] : 
                        (N586)? mem[4510] : 
                        (N588)? mem[4526] : 
                        (N590)? mem[4542] : 
                        (N592)? mem[4558] : 
                        (N594)? mem[4574] : 
                        (N596)? mem[4590] : 
                        (N598)? mem[4606] : 
                        (N600)? mem[4622] : 
                        (N602)? mem[4638] : 
                        (N604)? mem[4654] : 
                        (N606)? mem[4670] : 
                        (N608)? mem[4686] : 
                        (N610)? mem[4702] : 
                        (N612)? mem[4718] : 
                        (N614)? mem[4734] : 
                        (N616)? mem[4750] : 
                        (N618)? mem[4766] : 
                        (N620)? mem[4782] : 
                        (N622)? mem[4798] : 
                        (N624)? mem[4814] : 
                        (N626)? mem[4830] : 
                        (N628)? mem[4846] : 
                        (N630)? mem[4862] : 
                        (N632)? mem[4878] : 
                        (N634)? mem[4894] : 
                        (N636)? mem[4910] : 
                        (N638)? mem[4926] : 
                        (N640)? mem[4942] : 
                        (N642)? mem[4958] : 
                        (N644)? mem[4974] : 
                        (N646)? mem[4990] : 
                        (N648)? mem[5006] : 
                        (N650)? mem[5022] : 
                        (N652)? mem[5038] : 
                        (N654)? mem[5054] : 
                        (N656)? mem[5070] : 
                        (N658)? mem[5086] : 
                        (N660)? mem[5102] : 
                        (N662)? mem[5118] : 
                        (N664)? mem[5134] : 
                        (N666)? mem[5150] : 
                        (N668)? mem[5166] : 
                        (N670)? mem[5182] : 
                        (N672)? mem[5198] : 
                        (N674)? mem[5214] : 
                        (N676)? mem[5230] : 
                        (N678)? mem[5246] : 
                        (N680)? mem[5262] : 
                        (N682)? mem[5278] : 
                        (N684)? mem[5294] : 
                        (N686)? mem[5310] : 
                        (N688)? mem[5326] : 
                        (N690)? mem[5342] : 
                        (N692)? mem[5358] : 
                        (N694)? mem[5374] : 
                        (N696)? mem[5390] : 
                        (N698)? mem[5406] : 
                        (N700)? mem[5422] : 
                        (N702)? mem[5438] : 
                        (N704)? mem[5454] : 
                        (N706)? mem[5470] : 
                        (N708)? mem[5486] : 
                        (N710)? mem[5502] : 
                        (N712)? mem[5518] : 
                        (N714)? mem[5534] : 
                        (N716)? mem[5550] : 
                        (N718)? mem[5566] : 
                        (N720)? mem[5582] : 
                        (N722)? mem[5598] : 
                        (N724)? mem[5614] : 
                        (N726)? mem[5630] : 
                        (N728)? mem[5646] : 
                        (N730)? mem[5662] : 
                        (N732)? mem[5678] : 
                        (N734)? mem[5694] : 
                        (N736)? mem[5710] : 
                        (N738)? mem[5726] : 
                        (N740)? mem[5742] : 
                        (N742)? mem[5758] : 
                        (N744)? mem[5774] : 
                        (N746)? mem[5790] : 
                        (N748)? mem[5806] : 
                        (N750)? mem[5822] : 
                        (N752)? mem[5838] : 
                        (N754)? mem[5854] : 
                        (N756)? mem[5870] : 
                        (N758)? mem[5886] : 
                        (N760)? mem[5902] : 
                        (N762)? mem[5918] : 
                        (N764)? mem[5934] : 
                        (N766)? mem[5950] : 
                        (N768)? mem[5966] : 
                        (N770)? mem[5982] : 
                        (N772)? mem[5998] : 
                        (N774)? mem[6014] : 
                        (N776)? mem[6030] : 
                        (N778)? mem[6046] : 
                        (N780)? mem[6062] : 
                        (N782)? mem[6078] : 
                        (N784)? mem[6094] : 
                        (N786)? mem[6110] : 
                        (N788)? mem[6126] : 
                        (N790)? mem[6142] : 
                        (N792)? mem[6158] : 
                        (N794)? mem[6174] : 
                        (N796)? mem[6190] : 
                        (N798)? mem[6206] : 
                        (N800)? mem[6222] : 
                        (N802)? mem[6238] : 
                        (N804)? mem[6254] : 
                        (N806)? mem[6270] : 
                        (N808)? mem[6286] : 
                        (N810)? mem[6302] : 
                        (N812)? mem[6318] : 
                        (N814)? mem[6334] : 
                        (N816)? mem[6350] : 
                        (N818)? mem[6366] : 
                        (N820)? mem[6382] : 
                        (N822)? mem[6398] : 
                        (N824)? mem[6414] : 
                        (N826)? mem[6430] : 
                        (N828)? mem[6446] : 
                        (N830)? mem[6462] : 
                        (N832)? mem[6478] : 
                        (N834)? mem[6494] : 
                        (N836)? mem[6510] : 
                        (N838)? mem[6526] : 
                        (N840)? mem[6542] : 
                        (N842)? mem[6558] : 
                        (N844)? mem[6574] : 
                        (N846)? mem[6590] : 
                        (N848)? mem[6606] : 
                        (N850)? mem[6622] : 
                        (N852)? mem[6638] : 
                        (N854)? mem[6654] : 
                        (N856)? mem[6670] : 
                        (N858)? mem[6686] : 
                        (N860)? mem[6702] : 
                        (N862)? mem[6718] : 
                        (N864)? mem[6734] : 
                        (N866)? mem[6750] : 
                        (N868)? mem[6766] : 
                        (N870)? mem[6782] : 
                        (N872)? mem[6798] : 
                        (N874)? mem[6814] : 
                        (N876)? mem[6830] : 
                        (N878)? mem[6846] : 
                        (N880)? mem[6862] : 
                        (N882)? mem[6878] : 
                        (N884)? mem[6894] : 
                        (N886)? mem[6910] : 
                        (N888)? mem[6926] : 
                        (N890)? mem[6942] : 
                        (N892)? mem[6958] : 
                        (N894)? mem[6974] : 
                        (N896)? mem[6990] : 
                        (N898)? mem[7006] : 
                        (N900)? mem[7022] : 
                        (N902)? mem[7038] : 
                        (N904)? mem[7054] : 
                        (N906)? mem[7070] : 
                        (N908)? mem[7086] : 
                        (N910)? mem[7102] : 
                        (N912)? mem[7118] : 
                        (N914)? mem[7134] : 
                        (N916)? mem[7150] : 
                        (N918)? mem[7166] : 
                        (N920)? mem[7182] : 
                        (N922)? mem[7198] : 
                        (N924)? mem[7214] : 
                        (N926)? mem[7230] : 
                        (N928)? mem[7246] : 
                        (N930)? mem[7262] : 
                        (N932)? mem[7278] : 
                        (N934)? mem[7294] : 
                        (N936)? mem[7310] : 
                        (N938)? mem[7326] : 
                        (N940)? mem[7342] : 
                        (N942)? mem[7358] : 
                        (N944)? mem[7374] : 
                        (N946)? mem[7390] : 
                        (N948)? mem[7406] : 
                        (N950)? mem[7422] : 
                        (N952)? mem[7438] : 
                        (N954)? mem[7454] : 
                        (N956)? mem[7470] : 
                        (N958)? mem[7486] : 
                        (N960)? mem[7502] : 
                        (N962)? mem[7518] : 
                        (N964)? mem[7534] : 
                        (N966)? mem[7550] : 
                        (N968)? mem[7566] : 
                        (N970)? mem[7582] : 
                        (N972)? mem[7598] : 
                        (N974)? mem[7614] : 
                        (N976)? mem[7630] : 
                        (N978)? mem[7646] : 
                        (N980)? mem[7662] : 
                        (N982)? mem[7678] : 
                        (N984)? mem[7694] : 
                        (N986)? mem[7710] : 
                        (N988)? mem[7726] : 
                        (N990)? mem[7742] : 
                        (N992)? mem[7758] : 
                        (N994)? mem[7774] : 
                        (N996)? mem[7790] : 
                        (N998)? mem[7806] : 
                        (N1000)? mem[7822] : 
                        (N1002)? mem[7838] : 
                        (N1004)? mem[7854] : 
                        (N1006)? mem[7870] : 
                        (N1008)? mem[7886] : 
                        (N1010)? mem[7902] : 
                        (N1012)? mem[7918] : 
                        (N1014)? mem[7934] : 
                        (N1016)? mem[7950] : 
                        (N1018)? mem[7966] : 
                        (N1020)? mem[7982] : 
                        (N1022)? mem[7998] : 
                        (N1024)? mem[8014] : 
                        (N1026)? mem[8030] : 
                        (N1028)? mem[8046] : 
                        (N1030)? mem[8062] : 
                        (N1032)? mem[8078] : 
                        (N1034)? mem[8094] : 
                        (N1036)? mem[8110] : 
                        (N1038)? mem[8126] : 
                        (N1040)? mem[8142] : 
                        (N1042)? mem[8158] : 
                        (N1044)? mem[8174] : 
                        (N1046)? mem[8190] : 1'b0;
  assign r_data_o[13] = (N535)? mem[13] : 
                        (N537)? mem[29] : 
                        (N539)? mem[45] : 
                        (N541)? mem[61] : 
                        (N543)? mem[77] : 
                        (N545)? mem[93] : 
                        (N547)? mem[109] : 
                        (N549)? mem[125] : 
                        (N551)? mem[141] : 
                        (N553)? mem[157] : 
                        (N555)? mem[173] : 
                        (N557)? mem[189] : 
                        (N559)? mem[205] : 
                        (N561)? mem[221] : 
                        (N563)? mem[237] : 
                        (N565)? mem[253] : 
                        (N567)? mem[269] : 
                        (N569)? mem[285] : 
                        (N571)? mem[301] : 
                        (N573)? mem[317] : 
                        (N575)? mem[333] : 
                        (N577)? mem[349] : 
                        (N579)? mem[365] : 
                        (N581)? mem[381] : 
                        (N583)? mem[397] : 
                        (N585)? mem[413] : 
                        (N587)? mem[429] : 
                        (N589)? mem[445] : 
                        (N591)? mem[461] : 
                        (N593)? mem[477] : 
                        (N595)? mem[493] : 
                        (N597)? mem[509] : 
                        (N599)? mem[525] : 
                        (N601)? mem[541] : 
                        (N603)? mem[557] : 
                        (N605)? mem[573] : 
                        (N607)? mem[589] : 
                        (N609)? mem[605] : 
                        (N611)? mem[621] : 
                        (N613)? mem[637] : 
                        (N615)? mem[653] : 
                        (N617)? mem[669] : 
                        (N619)? mem[685] : 
                        (N621)? mem[701] : 
                        (N623)? mem[717] : 
                        (N625)? mem[733] : 
                        (N627)? mem[749] : 
                        (N629)? mem[765] : 
                        (N631)? mem[781] : 
                        (N633)? mem[797] : 
                        (N635)? mem[813] : 
                        (N637)? mem[829] : 
                        (N639)? mem[845] : 
                        (N641)? mem[861] : 
                        (N643)? mem[877] : 
                        (N645)? mem[893] : 
                        (N647)? mem[909] : 
                        (N649)? mem[925] : 
                        (N651)? mem[941] : 
                        (N653)? mem[957] : 
                        (N655)? mem[973] : 
                        (N657)? mem[989] : 
                        (N659)? mem[1005] : 
                        (N661)? mem[1021] : 
                        (N663)? mem[1037] : 
                        (N665)? mem[1053] : 
                        (N667)? mem[1069] : 
                        (N669)? mem[1085] : 
                        (N671)? mem[1101] : 
                        (N673)? mem[1117] : 
                        (N675)? mem[1133] : 
                        (N677)? mem[1149] : 
                        (N679)? mem[1165] : 
                        (N681)? mem[1181] : 
                        (N683)? mem[1197] : 
                        (N685)? mem[1213] : 
                        (N687)? mem[1229] : 
                        (N689)? mem[1245] : 
                        (N691)? mem[1261] : 
                        (N693)? mem[1277] : 
                        (N695)? mem[1293] : 
                        (N697)? mem[1309] : 
                        (N699)? mem[1325] : 
                        (N701)? mem[1341] : 
                        (N703)? mem[1357] : 
                        (N705)? mem[1373] : 
                        (N707)? mem[1389] : 
                        (N709)? mem[1405] : 
                        (N711)? mem[1421] : 
                        (N713)? mem[1437] : 
                        (N715)? mem[1453] : 
                        (N717)? mem[1469] : 
                        (N719)? mem[1485] : 
                        (N721)? mem[1501] : 
                        (N723)? mem[1517] : 
                        (N725)? mem[1533] : 
                        (N727)? mem[1549] : 
                        (N729)? mem[1565] : 
                        (N731)? mem[1581] : 
                        (N733)? mem[1597] : 
                        (N735)? mem[1613] : 
                        (N737)? mem[1629] : 
                        (N739)? mem[1645] : 
                        (N741)? mem[1661] : 
                        (N743)? mem[1677] : 
                        (N745)? mem[1693] : 
                        (N747)? mem[1709] : 
                        (N749)? mem[1725] : 
                        (N751)? mem[1741] : 
                        (N753)? mem[1757] : 
                        (N755)? mem[1773] : 
                        (N757)? mem[1789] : 
                        (N759)? mem[1805] : 
                        (N761)? mem[1821] : 
                        (N763)? mem[1837] : 
                        (N765)? mem[1853] : 
                        (N767)? mem[1869] : 
                        (N769)? mem[1885] : 
                        (N771)? mem[1901] : 
                        (N773)? mem[1917] : 
                        (N775)? mem[1933] : 
                        (N777)? mem[1949] : 
                        (N779)? mem[1965] : 
                        (N781)? mem[1981] : 
                        (N783)? mem[1997] : 
                        (N785)? mem[2013] : 
                        (N787)? mem[2029] : 
                        (N789)? mem[2045] : 
                        (N791)? mem[2061] : 
                        (N793)? mem[2077] : 
                        (N795)? mem[2093] : 
                        (N797)? mem[2109] : 
                        (N799)? mem[2125] : 
                        (N801)? mem[2141] : 
                        (N803)? mem[2157] : 
                        (N805)? mem[2173] : 
                        (N807)? mem[2189] : 
                        (N809)? mem[2205] : 
                        (N811)? mem[2221] : 
                        (N813)? mem[2237] : 
                        (N815)? mem[2253] : 
                        (N817)? mem[2269] : 
                        (N819)? mem[2285] : 
                        (N821)? mem[2301] : 
                        (N823)? mem[2317] : 
                        (N825)? mem[2333] : 
                        (N827)? mem[2349] : 
                        (N829)? mem[2365] : 
                        (N831)? mem[2381] : 
                        (N833)? mem[2397] : 
                        (N835)? mem[2413] : 
                        (N837)? mem[2429] : 
                        (N839)? mem[2445] : 
                        (N841)? mem[2461] : 
                        (N843)? mem[2477] : 
                        (N845)? mem[2493] : 
                        (N847)? mem[2509] : 
                        (N849)? mem[2525] : 
                        (N851)? mem[2541] : 
                        (N853)? mem[2557] : 
                        (N855)? mem[2573] : 
                        (N857)? mem[2589] : 
                        (N859)? mem[2605] : 
                        (N861)? mem[2621] : 
                        (N863)? mem[2637] : 
                        (N865)? mem[2653] : 
                        (N867)? mem[2669] : 
                        (N869)? mem[2685] : 
                        (N871)? mem[2701] : 
                        (N873)? mem[2717] : 
                        (N875)? mem[2733] : 
                        (N877)? mem[2749] : 
                        (N879)? mem[2765] : 
                        (N881)? mem[2781] : 
                        (N883)? mem[2797] : 
                        (N885)? mem[2813] : 
                        (N887)? mem[2829] : 
                        (N889)? mem[2845] : 
                        (N891)? mem[2861] : 
                        (N893)? mem[2877] : 
                        (N895)? mem[2893] : 
                        (N897)? mem[2909] : 
                        (N899)? mem[2925] : 
                        (N901)? mem[2941] : 
                        (N903)? mem[2957] : 
                        (N905)? mem[2973] : 
                        (N907)? mem[2989] : 
                        (N909)? mem[3005] : 
                        (N911)? mem[3021] : 
                        (N913)? mem[3037] : 
                        (N915)? mem[3053] : 
                        (N917)? mem[3069] : 
                        (N919)? mem[3085] : 
                        (N921)? mem[3101] : 
                        (N923)? mem[3117] : 
                        (N925)? mem[3133] : 
                        (N927)? mem[3149] : 
                        (N929)? mem[3165] : 
                        (N931)? mem[3181] : 
                        (N933)? mem[3197] : 
                        (N935)? mem[3213] : 
                        (N937)? mem[3229] : 
                        (N939)? mem[3245] : 
                        (N941)? mem[3261] : 
                        (N943)? mem[3277] : 
                        (N945)? mem[3293] : 
                        (N947)? mem[3309] : 
                        (N949)? mem[3325] : 
                        (N951)? mem[3341] : 
                        (N953)? mem[3357] : 
                        (N955)? mem[3373] : 
                        (N957)? mem[3389] : 
                        (N959)? mem[3405] : 
                        (N961)? mem[3421] : 
                        (N963)? mem[3437] : 
                        (N965)? mem[3453] : 
                        (N967)? mem[3469] : 
                        (N969)? mem[3485] : 
                        (N971)? mem[3501] : 
                        (N973)? mem[3517] : 
                        (N975)? mem[3533] : 
                        (N977)? mem[3549] : 
                        (N979)? mem[3565] : 
                        (N981)? mem[3581] : 
                        (N983)? mem[3597] : 
                        (N985)? mem[3613] : 
                        (N987)? mem[3629] : 
                        (N989)? mem[3645] : 
                        (N991)? mem[3661] : 
                        (N993)? mem[3677] : 
                        (N995)? mem[3693] : 
                        (N997)? mem[3709] : 
                        (N999)? mem[3725] : 
                        (N1001)? mem[3741] : 
                        (N1003)? mem[3757] : 
                        (N1005)? mem[3773] : 
                        (N1007)? mem[3789] : 
                        (N1009)? mem[3805] : 
                        (N1011)? mem[3821] : 
                        (N1013)? mem[3837] : 
                        (N1015)? mem[3853] : 
                        (N1017)? mem[3869] : 
                        (N1019)? mem[3885] : 
                        (N1021)? mem[3901] : 
                        (N1023)? mem[3917] : 
                        (N1025)? mem[3933] : 
                        (N1027)? mem[3949] : 
                        (N1029)? mem[3965] : 
                        (N1031)? mem[3981] : 
                        (N1033)? mem[3997] : 
                        (N1035)? mem[4013] : 
                        (N1037)? mem[4029] : 
                        (N1039)? mem[4045] : 
                        (N1041)? mem[4061] : 
                        (N1043)? mem[4077] : 
                        (N1045)? mem[4093] : 
                        (N536)? mem[4109] : 
                        (N538)? mem[4125] : 
                        (N540)? mem[4141] : 
                        (N542)? mem[4157] : 
                        (N544)? mem[4173] : 
                        (N546)? mem[4189] : 
                        (N548)? mem[4205] : 
                        (N550)? mem[4221] : 
                        (N552)? mem[4237] : 
                        (N554)? mem[4253] : 
                        (N556)? mem[4269] : 
                        (N558)? mem[4285] : 
                        (N560)? mem[4301] : 
                        (N562)? mem[4317] : 
                        (N564)? mem[4333] : 
                        (N566)? mem[4349] : 
                        (N568)? mem[4365] : 
                        (N570)? mem[4381] : 
                        (N572)? mem[4397] : 
                        (N574)? mem[4413] : 
                        (N576)? mem[4429] : 
                        (N578)? mem[4445] : 
                        (N580)? mem[4461] : 
                        (N582)? mem[4477] : 
                        (N584)? mem[4493] : 
                        (N586)? mem[4509] : 
                        (N588)? mem[4525] : 
                        (N590)? mem[4541] : 
                        (N592)? mem[4557] : 
                        (N594)? mem[4573] : 
                        (N596)? mem[4589] : 
                        (N598)? mem[4605] : 
                        (N600)? mem[4621] : 
                        (N602)? mem[4637] : 
                        (N604)? mem[4653] : 
                        (N606)? mem[4669] : 
                        (N608)? mem[4685] : 
                        (N610)? mem[4701] : 
                        (N612)? mem[4717] : 
                        (N614)? mem[4733] : 
                        (N616)? mem[4749] : 
                        (N618)? mem[4765] : 
                        (N620)? mem[4781] : 
                        (N622)? mem[4797] : 
                        (N624)? mem[4813] : 
                        (N626)? mem[4829] : 
                        (N628)? mem[4845] : 
                        (N630)? mem[4861] : 
                        (N632)? mem[4877] : 
                        (N634)? mem[4893] : 
                        (N636)? mem[4909] : 
                        (N638)? mem[4925] : 
                        (N640)? mem[4941] : 
                        (N642)? mem[4957] : 
                        (N644)? mem[4973] : 
                        (N646)? mem[4989] : 
                        (N648)? mem[5005] : 
                        (N650)? mem[5021] : 
                        (N652)? mem[5037] : 
                        (N654)? mem[5053] : 
                        (N656)? mem[5069] : 
                        (N658)? mem[5085] : 
                        (N660)? mem[5101] : 
                        (N662)? mem[5117] : 
                        (N664)? mem[5133] : 
                        (N666)? mem[5149] : 
                        (N668)? mem[5165] : 
                        (N670)? mem[5181] : 
                        (N672)? mem[5197] : 
                        (N674)? mem[5213] : 
                        (N676)? mem[5229] : 
                        (N678)? mem[5245] : 
                        (N680)? mem[5261] : 
                        (N682)? mem[5277] : 
                        (N684)? mem[5293] : 
                        (N686)? mem[5309] : 
                        (N688)? mem[5325] : 
                        (N690)? mem[5341] : 
                        (N692)? mem[5357] : 
                        (N694)? mem[5373] : 
                        (N696)? mem[5389] : 
                        (N698)? mem[5405] : 
                        (N700)? mem[5421] : 
                        (N702)? mem[5437] : 
                        (N704)? mem[5453] : 
                        (N706)? mem[5469] : 
                        (N708)? mem[5485] : 
                        (N710)? mem[5501] : 
                        (N712)? mem[5517] : 
                        (N714)? mem[5533] : 
                        (N716)? mem[5549] : 
                        (N718)? mem[5565] : 
                        (N720)? mem[5581] : 
                        (N722)? mem[5597] : 
                        (N724)? mem[5613] : 
                        (N726)? mem[5629] : 
                        (N728)? mem[5645] : 
                        (N730)? mem[5661] : 
                        (N732)? mem[5677] : 
                        (N734)? mem[5693] : 
                        (N736)? mem[5709] : 
                        (N738)? mem[5725] : 
                        (N740)? mem[5741] : 
                        (N742)? mem[5757] : 
                        (N744)? mem[5773] : 
                        (N746)? mem[5789] : 
                        (N748)? mem[5805] : 
                        (N750)? mem[5821] : 
                        (N752)? mem[5837] : 
                        (N754)? mem[5853] : 
                        (N756)? mem[5869] : 
                        (N758)? mem[5885] : 
                        (N760)? mem[5901] : 
                        (N762)? mem[5917] : 
                        (N764)? mem[5933] : 
                        (N766)? mem[5949] : 
                        (N768)? mem[5965] : 
                        (N770)? mem[5981] : 
                        (N772)? mem[5997] : 
                        (N774)? mem[6013] : 
                        (N776)? mem[6029] : 
                        (N778)? mem[6045] : 
                        (N780)? mem[6061] : 
                        (N782)? mem[6077] : 
                        (N784)? mem[6093] : 
                        (N786)? mem[6109] : 
                        (N788)? mem[6125] : 
                        (N790)? mem[6141] : 
                        (N792)? mem[6157] : 
                        (N794)? mem[6173] : 
                        (N796)? mem[6189] : 
                        (N798)? mem[6205] : 
                        (N800)? mem[6221] : 
                        (N802)? mem[6237] : 
                        (N804)? mem[6253] : 
                        (N806)? mem[6269] : 
                        (N808)? mem[6285] : 
                        (N810)? mem[6301] : 
                        (N812)? mem[6317] : 
                        (N814)? mem[6333] : 
                        (N816)? mem[6349] : 
                        (N818)? mem[6365] : 
                        (N820)? mem[6381] : 
                        (N822)? mem[6397] : 
                        (N824)? mem[6413] : 
                        (N826)? mem[6429] : 
                        (N828)? mem[6445] : 
                        (N830)? mem[6461] : 
                        (N832)? mem[6477] : 
                        (N834)? mem[6493] : 
                        (N836)? mem[6509] : 
                        (N838)? mem[6525] : 
                        (N840)? mem[6541] : 
                        (N842)? mem[6557] : 
                        (N844)? mem[6573] : 
                        (N846)? mem[6589] : 
                        (N848)? mem[6605] : 
                        (N850)? mem[6621] : 
                        (N852)? mem[6637] : 
                        (N854)? mem[6653] : 
                        (N856)? mem[6669] : 
                        (N858)? mem[6685] : 
                        (N860)? mem[6701] : 
                        (N862)? mem[6717] : 
                        (N864)? mem[6733] : 
                        (N866)? mem[6749] : 
                        (N868)? mem[6765] : 
                        (N870)? mem[6781] : 
                        (N872)? mem[6797] : 
                        (N874)? mem[6813] : 
                        (N876)? mem[6829] : 
                        (N878)? mem[6845] : 
                        (N880)? mem[6861] : 
                        (N882)? mem[6877] : 
                        (N884)? mem[6893] : 
                        (N886)? mem[6909] : 
                        (N888)? mem[6925] : 
                        (N890)? mem[6941] : 
                        (N892)? mem[6957] : 
                        (N894)? mem[6973] : 
                        (N896)? mem[6989] : 
                        (N898)? mem[7005] : 
                        (N900)? mem[7021] : 
                        (N902)? mem[7037] : 
                        (N904)? mem[7053] : 
                        (N906)? mem[7069] : 
                        (N908)? mem[7085] : 
                        (N910)? mem[7101] : 
                        (N912)? mem[7117] : 
                        (N914)? mem[7133] : 
                        (N916)? mem[7149] : 
                        (N918)? mem[7165] : 
                        (N920)? mem[7181] : 
                        (N922)? mem[7197] : 
                        (N924)? mem[7213] : 
                        (N926)? mem[7229] : 
                        (N928)? mem[7245] : 
                        (N930)? mem[7261] : 
                        (N932)? mem[7277] : 
                        (N934)? mem[7293] : 
                        (N936)? mem[7309] : 
                        (N938)? mem[7325] : 
                        (N940)? mem[7341] : 
                        (N942)? mem[7357] : 
                        (N944)? mem[7373] : 
                        (N946)? mem[7389] : 
                        (N948)? mem[7405] : 
                        (N950)? mem[7421] : 
                        (N952)? mem[7437] : 
                        (N954)? mem[7453] : 
                        (N956)? mem[7469] : 
                        (N958)? mem[7485] : 
                        (N960)? mem[7501] : 
                        (N962)? mem[7517] : 
                        (N964)? mem[7533] : 
                        (N966)? mem[7549] : 
                        (N968)? mem[7565] : 
                        (N970)? mem[7581] : 
                        (N972)? mem[7597] : 
                        (N974)? mem[7613] : 
                        (N976)? mem[7629] : 
                        (N978)? mem[7645] : 
                        (N980)? mem[7661] : 
                        (N982)? mem[7677] : 
                        (N984)? mem[7693] : 
                        (N986)? mem[7709] : 
                        (N988)? mem[7725] : 
                        (N990)? mem[7741] : 
                        (N992)? mem[7757] : 
                        (N994)? mem[7773] : 
                        (N996)? mem[7789] : 
                        (N998)? mem[7805] : 
                        (N1000)? mem[7821] : 
                        (N1002)? mem[7837] : 
                        (N1004)? mem[7853] : 
                        (N1006)? mem[7869] : 
                        (N1008)? mem[7885] : 
                        (N1010)? mem[7901] : 
                        (N1012)? mem[7917] : 
                        (N1014)? mem[7933] : 
                        (N1016)? mem[7949] : 
                        (N1018)? mem[7965] : 
                        (N1020)? mem[7981] : 
                        (N1022)? mem[7997] : 
                        (N1024)? mem[8013] : 
                        (N1026)? mem[8029] : 
                        (N1028)? mem[8045] : 
                        (N1030)? mem[8061] : 
                        (N1032)? mem[8077] : 
                        (N1034)? mem[8093] : 
                        (N1036)? mem[8109] : 
                        (N1038)? mem[8125] : 
                        (N1040)? mem[8141] : 
                        (N1042)? mem[8157] : 
                        (N1044)? mem[8173] : 
                        (N1046)? mem[8189] : 1'b0;
  assign r_data_o[12] = (N535)? mem[12] : 
                        (N537)? mem[28] : 
                        (N539)? mem[44] : 
                        (N541)? mem[60] : 
                        (N543)? mem[76] : 
                        (N545)? mem[92] : 
                        (N547)? mem[108] : 
                        (N549)? mem[124] : 
                        (N551)? mem[140] : 
                        (N553)? mem[156] : 
                        (N555)? mem[172] : 
                        (N557)? mem[188] : 
                        (N559)? mem[204] : 
                        (N561)? mem[220] : 
                        (N563)? mem[236] : 
                        (N565)? mem[252] : 
                        (N567)? mem[268] : 
                        (N569)? mem[284] : 
                        (N571)? mem[300] : 
                        (N573)? mem[316] : 
                        (N575)? mem[332] : 
                        (N577)? mem[348] : 
                        (N579)? mem[364] : 
                        (N581)? mem[380] : 
                        (N583)? mem[396] : 
                        (N585)? mem[412] : 
                        (N587)? mem[428] : 
                        (N589)? mem[444] : 
                        (N591)? mem[460] : 
                        (N593)? mem[476] : 
                        (N595)? mem[492] : 
                        (N597)? mem[508] : 
                        (N599)? mem[524] : 
                        (N601)? mem[540] : 
                        (N603)? mem[556] : 
                        (N605)? mem[572] : 
                        (N607)? mem[588] : 
                        (N609)? mem[604] : 
                        (N611)? mem[620] : 
                        (N613)? mem[636] : 
                        (N615)? mem[652] : 
                        (N617)? mem[668] : 
                        (N619)? mem[684] : 
                        (N621)? mem[700] : 
                        (N623)? mem[716] : 
                        (N625)? mem[732] : 
                        (N627)? mem[748] : 
                        (N629)? mem[764] : 
                        (N631)? mem[780] : 
                        (N633)? mem[796] : 
                        (N635)? mem[812] : 
                        (N637)? mem[828] : 
                        (N639)? mem[844] : 
                        (N641)? mem[860] : 
                        (N643)? mem[876] : 
                        (N645)? mem[892] : 
                        (N647)? mem[908] : 
                        (N649)? mem[924] : 
                        (N651)? mem[940] : 
                        (N653)? mem[956] : 
                        (N655)? mem[972] : 
                        (N657)? mem[988] : 
                        (N659)? mem[1004] : 
                        (N661)? mem[1020] : 
                        (N663)? mem[1036] : 
                        (N665)? mem[1052] : 
                        (N667)? mem[1068] : 
                        (N669)? mem[1084] : 
                        (N671)? mem[1100] : 
                        (N673)? mem[1116] : 
                        (N675)? mem[1132] : 
                        (N677)? mem[1148] : 
                        (N679)? mem[1164] : 
                        (N681)? mem[1180] : 
                        (N683)? mem[1196] : 
                        (N685)? mem[1212] : 
                        (N687)? mem[1228] : 
                        (N689)? mem[1244] : 
                        (N691)? mem[1260] : 
                        (N693)? mem[1276] : 
                        (N695)? mem[1292] : 
                        (N697)? mem[1308] : 
                        (N699)? mem[1324] : 
                        (N701)? mem[1340] : 
                        (N703)? mem[1356] : 
                        (N705)? mem[1372] : 
                        (N707)? mem[1388] : 
                        (N709)? mem[1404] : 
                        (N711)? mem[1420] : 
                        (N713)? mem[1436] : 
                        (N715)? mem[1452] : 
                        (N717)? mem[1468] : 
                        (N719)? mem[1484] : 
                        (N721)? mem[1500] : 
                        (N723)? mem[1516] : 
                        (N725)? mem[1532] : 
                        (N727)? mem[1548] : 
                        (N729)? mem[1564] : 
                        (N731)? mem[1580] : 
                        (N733)? mem[1596] : 
                        (N735)? mem[1612] : 
                        (N737)? mem[1628] : 
                        (N739)? mem[1644] : 
                        (N741)? mem[1660] : 
                        (N743)? mem[1676] : 
                        (N745)? mem[1692] : 
                        (N747)? mem[1708] : 
                        (N749)? mem[1724] : 
                        (N751)? mem[1740] : 
                        (N753)? mem[1756] : 
                        (N755)? mem[1772] : 
                        (N757)? mem[1788] : 
                        (N759)? mem[1804] : 
                        (N761)? mem[1820] : 
                        (N763)? mem[1836] : 
                        (N765)? mem[1852] : 
                        (N767)? mem[1868] : 
                        (N769)? mem[1884] : 
                        (N771)? mem[1900] : 
                        (N773)? mem[1916] : 
                        (N775)? mem[1932] : 
                        (N777)? mem[1948] : 
                        (N779)? mem[1964] : 
                        (N781)? mem[1980] : 
                        (N783)? mem[1996] : 
                        (N785)? mem[2012] : 
                        (N787)? mem[2028] : 
                        (N789)? mem[2044] : 
                        (N791)? mem[2060] : 
                        (N793)? mem[2076] : 
                        (N795)? mem[2092] : 
                        (N797)? mem[2108] : 
                        (N799)? mem[2124] : 
                        (N801)? mem[2140] : 
                        (N803)? mem[2156] : 
                        (N805)? mem[2172] : 
                        (N807)? mem[2188] : 
                        (N809)? mem[2204] : 
                        (N811)? mem[2220] : 
                        (N813)? mem[2236] : 
                        (N815)? mem[2252] : 
                        (N817)? mem[2268] : 
                        (N819)? mem[2284] : 
                        (N821)? mem[2300] : 
                        (N823)? mem[2316] : 
                        (N825)? mem[2332] : 
                        (N827)? mem[2348] : 
                        (N829)? mem[2364] : 
                        (N831)? mem[2380] : 
                        (N833)? mem[2396] : 
                        (N835)? mem[2412] : 
                        (N837)? mem[2428] : 
                        (N839)? mem[2444] : 
                        (N841)? mem[2460] : 
                        (N843)? mem[2476] : 
                        (N845)? mem[2492] : 
                        (N847)? mem[2508] : 
                        (N849)? mem[2524] : 
                        (N851)? mem[2540] : 
                        (N853)? mem[2556] : 
                        (N855)? mem[2572] : 
                        (N857)? mem[2588] : 
                        (N859)? mem[2604] : 
                        (N861)? mem[2620] : 
                        (N863)? mem[2636] : 
                        (N865)? mem[2652] : 
                        (N867)? mem[2668] : 
                        (N869)? mem[2684] : 
                        (N871)? mem[2700] : 
                        (N873)? mem[2716] : 
                        (N875)? mem[2732] : 
                        (N877)? mem[2748] : 
                        (N879)? mem[2764] : 
                        (N881)? mem[2780] : 
                        (N883)? mem[2796] : 
                        (N885)? mem[2812] : 
                        (N887)? mem[2828] : 
                        (N889)? mem[2844] : 
                        (N891)? mem[2860] : 
                        (N893)? mem[2876] : 
                        (N895)? mem[2892] : 
                        (N897)? mem[2908] : 
                        (N899)? mem[2924] : 
                        (N901)? mem[2940] : 
                        (N903)? mem[2956] : 
                        (N905)? mem[2972] : 
                        (N907)? mem[2988] : 
                        (N909)? mem[3004] : 
                        (N911)? mem[3020] : 
                        (N913)? mem[3036] : 
                        (N915)? mem[3052] : 
                        (N917)? mem[3068] : 
                        (N919)? mem[3084] : 
                        (N921)? mem[3100] : 
                        (N923)? mem[3116] : 
                        (N925)? mem[3132] : 
                        (N927)? mem[3148] : 
                        (N929)? mem[3164] : 
                        (N931)? mem[3180] : 
                        (N933)? mem[3196] : 
                        (N935)? mem[3212] : 
                        (N937)? mem[3228] : 
                        (N939)? mem[3244] : 
                        (N941)? mem[3260] : 
                        (N943)? mem[3276] : 
                        (N945)? mem[3292] : 
                        (N947)? mem[3308] : 
                        (N949)? mem[3324] : 
                        (N951)? mem[3340] : 
                        (N953)? mem[3356] : 
                        (N955)? mem[3372] : 
                        (N957)? mem[3388] : 
                        (N959)? mem[3404] : 
                        (N961)? mem[3420] : 
                        (N963)? mem[3436] : 
                        (N965)? mem[3452] : 
                        (N967)? mem[3468] : 
                        (N969)? mem[3484] : 
                        (N971)? mem[3500] : 
                        (N973)? mem[3516] : 
                        (N975)? mem[3532] : 
                        (N977)? mem[3548] : 
                        (N979)? mem[3564] : 
                        (N981)? mem[3580] : 
                        (N983)? mem[3596] : 
                        (N985)? mem[3612] : 
                        (N987)? mem[3628] : 
                        (N989)? mem[3644] : 
                        (N991)? mem[3660] : 
                        (N993)? mem[3676] : 
                        (N995)? mem[3692] : 
                        (N997)? mem[3708] : 
                        (N999)? mem[3724] : 
                        (N1001)? mem[3740] : 
                        (N1003)? mem[3756] : 
                        (N1005)? mem[3772] : 
                        (N1007)? mem[3788] : 
                        (N1009)? mem[3804] : 
                        (N1011)? mem[3820] : 
                        (N1013)? mem[3836] : 
                        (N1015)? mem[3852] : 
                        (N1017)? mem[3868] : 
                        (N1019)? mem[3884] : 
                        (N1021)? mem[3900] : 
                        (N1023)? mem[3916] : 
                        (N1025)? mem[3932] : 
                        (N1027)? mem[3948] : 
                        (N1029)? mem[3964] : 
                        (N1031)? mem[3980] : 
                        (N1033)? mem[3996] : 
                        (N1035)? mem[4012] : 
                        (N1037)? mem[4028] : 
                        (N1039)? mem[4044] : 
                        (N1041)? mem[4060] : 
                        (N1043)? mem[4076] : 
                        (N1045)? mem[4092] : 
                        (N536)? mem[4108] : 
                        (N538)? mem[4124] : 
                        (N540)? mem[4140] : 
                        (N542)? mem[4156] : 
                        (N544)? mem[4172] : 
                        (N546)? mem[4188] : 
                        (N548)? mem[4204] : 
                        (N550)? mem[4220] : 
                        (N552)? mem[4236] : 
                        (N554)? mem[4252] : 
                        (N556)? mem[4268] : 
                        (N558)? mem[4284] : 
                        (N560)? mem[4300] : 
                        (N562)? mem[4316] : 
                        (N564)? mem[4332] : 
                        (N566)? mem[4348] : 
                        (N568)? mem[4364] : 
                        (N570)? mem[4380] : 
                        (N572)? mem[4396] : 
                        (N574)? mem[4412] : 
                        (N576)? mem[4428] : 
                        (N578)? mem[4444] : 
                        (N580)? mem[4460] : 
                        (N582)? mem[4476] : 
                        (N584)? mem[4492] : 
                        (N586)? mem[4508] : 
                        (N588)? mem[4524] : 
                        (N590)? mem[4540] : 
                        (N592)? mem[4556] : 
                        (N594)? mem[4572] : 
                        (N596)? mem[4588] : 
                        (N598)? mem[4604] : 
                        (N600)? mem[4620] : 
                        (N602)? mem[4636] : 
                        (N604)? mem[4652] : 
                        (N606)? mem[4668] : 
                        (N608)? mem[4684] : 
                        (N610)? mem[4700] : 
                        (N612)? mem[4716] : 
                        (N614)? mem[4732] : 
                        (N616)? mem[4748] : 
                        (N618)? mem[4764] : 
                        (N620)? mem[4780] : 
                        (N622)? mem[4796] : 
                        (N624)? mem[4812] : 
                        (N626)? mem[4828] : 
                        (N628)? mem[4844] : 
                        (N630)? mem[4860] : 
                        (N632)? mem[4876] : 
                        (N634)? mem[4892] : 
                        (N636)? mem[4908] : 
                        (N638)? mem[4924] : 
                        (N640)? mem[4940] : 
                        (N642)? mem[4956] : 
                        (N644)? mem[4972] : 
                        (N646)? mem[4988] : 
                        (N648)? mem[5004] : 
                        (N650)? mem[5020] : 
                        (N652)? mem[5036] : 
                        (N654)? mem[5052] : 
                        (N656)? mem[5068] : 
                        (N658)? mem[5084] : 
                        (N660)? mem[5100] : 
                        (N662)? mem[5116] : 
                        (N664)? mem[5132] : 
                        (N666)? mem[5148] : 
                        (N668)? mem[5164] : 
                        (N670)? mem[5180] : 
                        (N672)? mem[5196] : 
                        (N674)? mem[5212] : 
                        (N676)? mem[5228] : 
                        (N678)? mem[5244] : 
                        (N680)? mem[5260] : 
                        (N682)? mem[5276] : 
                        (N684)? mem[5292] : 
                        (N686)? mem[5308] : 
                        (N688)? mem[5324] : 
                        (N690)? mem[5340] : 
                        (N692)? mem[5356] : 
                        (N694)? mem[5372] : 
                        (N696)? mem[5388] : 
                        (N698)? mem[5404] : 
                        (N700)? mem[5420] : 
                        (N702)? mem[5436] : 
                        (N704)? mem[5452] : 
                        (N706)? mem[5468] : 
                        (N708)? mem[5484] : 
                        (N710)? mem[5500] : 
                        (N712)? mem[5516] : 
                        (N714)? mem[5532] : 
                        (N716)? mem[5548] : 
                        (N718)? mem[5564] : 
                        (N720)? mem[5580] : 
                        (N722)? mem[5596] : 
                        (N724)? mem[5612] : 
                        (N726)? mem[5628] : 
                        (N728)? mem[5644] : 
                        (N730)? mem[5660] : 
                        (N732)? mem[5676] : 
                        (N734)? mem[5692] : 
                        (N736)? mem[5708] : 
                        (N738)? mem[5724] : 
                        (N740)? mem[5740] : 
                        (N742)? mem[5756] : 
                        (N744)? mem[5772] : 
                        (N746)? mem[5788] : 
                        (N748)? mem[5804] : 
                        (N750)? mem[5820] : 
                        (N752)? mem[5836] : 
                        (N754)? mem[5852] : 
                        (N756)? mem[5868] : 
                        (N758)? mem[5884] : 
                        (N760)? mem[5900] : 
                        (N762)? mem[5916] : 
                        (N764)? mem[5932] : 
                        (N766)? mem[5948] : 
                        (N768)? mem[5964] : 
                        (N770)? mem[5980] : 
                        (N772)? mem[5996] : 
                        (N774)? mem[6012] : 
                        (N776)? mem[6028] : 
                        (N778)? mem[6044] : 
                        (N780)? mem[6060] : 
                        (N782)? mem[6076] : 
                        (N784)? mem[6092] : 
                        (N786)? mem[6108] : 
                        (N788)? mem[6124] : 
                        (N790)? mem[6140] : 
                        (N792)? mem[6156] : 
                        (N794)? mem[6172] : 
                        (N796)? mem[6188] : 
                        (N798)? mem[6204] : 
                        (N800)? mem[6220] : 
                        (N802)? mem[6236] : 
                        (N804)? mem[6252] : 
                        (N806)? mem[6268] : 
                        (N808)? mem[6284] : 
                        (N810)? mem[6300] : 
                        (N812)? mem[6316] : 
                        (N814)? mem[6332] : 
                        (N816)? mem[6348] : 
                        (N818)? mem[6364] : 
                        (N820)? mem[6380] : 
                        (N822)? mem[6396] : 
                        (N824)? mem[6412] : 
                        (N826)? mem[6428] : 
                        (N828)? mem[6444] : 
                        (N830)? mem[6460] : 
                        (N832)? mem[6476] : 
                        (N834)? mem[6492] : 
                        (N836)? mem[6508] : 
                        (N838)? mem[6524] : 
                        (N840)? mem[6540] : 
                        (N842)? mem[6556] : 
                        (N844)? mem[6572] : 
                        (N846)? mem[6588] : 
                        (N848)? mem[6604] : 
                        (N850)? mem[6620] : 
                        (N852)? mem[6636] : 
                        (N854)? mem[6652] : 
                        (N856)? mem[6668] : 
                        (N858)? mem[6684] : 
                        (N860)? mem[6700] : 
                        (N862)? mem[6716] : 
                        (N864)? mem[6732] : 
                        (N866)? mem[6748] : 
                        (N868)? mem[6764] : 
                        (N870)? mem[6780] : 
                        (N872)? mem[6796] : 
                        (N874)? mem[6812] : 
                        (N876)? mem[6828] : 
                        (N878)? mem[6844] : 
                        (N880)? mem[6860] : 
                        (N882)? mem[6876] : 
                        (N884)? mem[6892] : 
                        (N886)? mem[6908] : 
                        (N888)? mem[6924] : 
                        (N890)? mem[6940] : 
                        (N892)? mem[6956] : 
                        (N894)? mem[6972] : 
                        (N896)? mem[6988] : 
                        (N898)? mem[7004] : 
                        (N900)? mem[7020] : 
                        (N902)? mem[7036] : 
                        (N904)? mem[7052] : 
                        (N906)? mem[7068] : 
                        (N908)? mem[7084] : 
                        (N910)? mem[7100] : 
                        (N912)? mem[7116] : 
                        (N914)? mem[7132] : 
                        (N916)? mem[7148] : 
                        (N918)? mem[7164] : 
                        (N920)? mem[7180] : 
                        (N922)? mem[7196] : 
                        (N924)? mem[7212] : 
                        (N926)? mem[7228] : 
                        (N928)? mem[7244] : 
                        (N930)? mem[7260] : 
                        (N932)? mem[7276] : 
                        (N934)? mem[7292] : 
                        (N936)? mem[7308] : 
                        (N938)? mem[7324] : 
                        (N940)? mem[7340] : 
                        (N942)? mem[7356] : 
                        (N944)? mem[7372] : 
                        (N946)? mem[7388] : 
                        (N948)? mem[7404] : 
                        (N950)? mem[7420] : 
                        (N952)? mem[7436] : 
                        (N954)? mem[7452] : 
                        (N956)? mem[7468] : 
                        (N958)? mem[7484] : 
                        (N960)? mem[7500] : 
                        (N962)? mem[7516] : 
                        (N964)? mem[7532] : 
                        (N966)? mem[7548] : 
                        (N968)? mem[7564] : 
                        (N970)? mem[7580] : 
                        (N972)? mem[7596] : 
                        (N974)? mem[7612] : 
                        (N976)? mem[7628] : 
                        (N978)? mem[7644] : 
                        (N980)? mem[7660] : 
                        (N982)? mem[7676] : 
                        (N984)? mem[7692] : 
                        (N986)? mem[7708] : 
                        (N988)? mem[7724] : 
                        (N990)? mem[7740] : 
                        (N992)? mem[7756] : 
                        (N994)? mem[7772] : 
                        (N996)? mem[7788] : 
                        (N998)? mem[7804] : 
                        (N1000)? mem[7820] : 
                        (N1002)? mem[7836] : 
                        (N1004)? mem[7852] : 
                        (N1006)? mem[7868] : 
                        (N1008)? mem[7884] : 
                        (N1010)? mem[7900] : 
                        (N1012)? mem[7916] : 
                        (N1014)? mem[7932] : 
                        (N1016)? mem[7948] : 
                        (N1018)? mem[7964] : 
                        (N1020)? mem[7980] : 
                        (N1022)? mem[7996] : 
                        (N1024)? mem[8012] : 
                        (N1026)? mem[8028] : 
                        (N1028)? mem[8044] : 
                        (N1030)? mem[8060] : 
                        (N1032)? mem[8076] : 
                        (N1034)? mem[8092] : 
                        (N1036)? mem[8108] : 
                        (N1038)? mem[8124] : 
                        (N1040)? mem[8140] : 
                        (N1042)? mem[8156] : 
                        (N1044)? mem[8172] : 
                        (N1046)? mem[8188] : 1'b0;
  assign r_data_o[11] = (N535)? mem[11] : 
                        (N537)? mem[27] : 
                        (N539)? mem[43] : 
                        (N541)? mem[59] : 
                        (N543)? mem[75] : 
                        (N545)? mem[91] : 
                        (N547)? mem[107] : 
                        (N549)? mem[123] : 
                        (N551)? mem[139] : 
                        (N553)? mem[155] : 
                        (N555)? mem[171] : 
                        (N557)? mem[187] : 
                        (N559)? mem[203] : 
                        (N561)? mem[219] : 
                        (N563)? mem[235] : 
                        (N565)? mem[251] : 
                        (N567)? mem[267] : 
                        (N569)? mem[283] : 
                        (N571)? mem[299] : 
                        (N573)? mem[315] : 
                        (N575)? mem[331] : 
                        (N577)? mem[347] : 
                        (N579)? mem[363] : 
                        (N581)? mem[379] : 
                        (N583)? mem[395] : 
                        (N585)? mem[411] : 
                        (N587)? mem[427] : 
                        (N589)? mem[443] : 
                        (N591)? mem[459] : 
                        (N593)? mem[475] : 
                        (N595)? mem[491] : 
                        (N597)? mem[507] : 
                        (N599)? mem[523] : 
                        (N601)? mem[539] : 
                        (N603)? mem[555] : 
                        (N605)? mem[571] : 
                        (N607)? mem[587] : 
                        (N609)? mem[603] : 
                        (N611)? mem[619] : 
                        (N613)? mem[635] : 
                        (N615)? mem[651] : 
                        (N617)? mem[667] : 
                        (N619)? mem[683] : 
                        (N621)? mem[699] : 
                        (N623)? mem[715] : 
                        (N625)? mem[731] : 
                        (N627)? mem[747] : 
                        (N629)? mem[763] : 
                        (N631)? mem[779] : 
                        (N633)? mem[795] : 
                        (N635)? mem[811] : 
                        (N637)? mem[827] : 
                        (N639)? mem[843] : 
                        (N641)? mem[859] : 
                        (N643)? mem[875] : 
                        (N645)? mem[891] : 
                        (N647)? mem[907] : 
                        (N649)? mem[923] : 
                        (N651)? mem[939] : 
                        (N653)? mem[955] : 
                        (N655)? mem[971] : 
                        (N657)? mem[987] : 
                        (N659)? mem[1003] : 
                        (N661)? mem[1019] : 
                        (N663)? mem[1035] : 
                        (N665)? mem[1051] : 
                        (N667)? mem[1067] : 
                        (N669)? mem[1083] : 
                        (N671)? mem[1099] : 
                        (N673)? mem[1115] : 
                        (N675)? mem[1131] : 
                        (N677)? mem[1147] : 
                        (N679)? mem[1163] : 
                        (N681)? mem[1179] : 
                        (N683)? mem[1195] : 
                        (N685)? mem[1211] : 
                        (N687)? mem[1227] : 
                        (N689)? mem[1243] : 
                        (N691)? mem[1259] : 
                        (N693)? mem[1275] : 
                        (N695)? mem[1291] : 
                        (N697)? mem[1307] : 
                        (N699)? mem[1323] : 
                        (N701)? mem[1339] : 
                        (N703)? mem[1355] : 
                        (N705)? mem[1371] : 
                        (N707)? mem[1387] : 
                        (N709)? mem[1403] : 
                        (N711)? mem[1419] : 
                        (N713)? mem[1435] : 
                        (N715)? mem[1451] : 
                        (N717)? mem[1467] : 
                        (N719)? mem[1483] : 
                        (N721)? mem[1499] : 
                        (N723)? mem[1515] : 
                        (N725)? mem[1531] : 
                        (N727)? mem[1547] : 
                        (N729)? mem[1563] : 
                        (N731)? mem[1579] : 
                        (N733)? mem[1595] : 
                        (N735)? mem[1611] : 
                        (N737)? mem[1627] : 
                        (N739)? mem[1643] : 
                        (N741)? mem[1659] : 
                        (N743)? mem[1675] : 
                        (N745)? mem[1691] : 
                        (N747)? mem[1707] : 
                        (N749)? mem[1723] : 
                        (N751)? mem[1739] : 
                        (N753)? mem[1755] : 
                        (N755)? mem[1771] : 
                        (N757)? mem[1787] : 
                        (N759)? mem[1803] : 
                        (N761)? mem[1819] : 
                        (N763)? mem[1835] : 
                        (N765)? mem[1851] : 
                        (N767)? mem[1867] : 
                        (N769)? mem[1883] : 
                        (N771)? mem[1899] : 
                        (N773)? mem[1915] : 
                        (N775)? mem[1931] : 
                        (N777)? mem[1947] : 
                        (N779)? mem[1963] : 
                        (N781)? mem[1979] : 
                        (N783)? mem[1995] : 
                        (N785)? mem[2011] : 
                        (N787)? mem[2027] : 
                        (N789)? mem[2043] : 
                        (N791)? mem[2059] : 
                        (N793)? mem[2075] : 
                        (N795)? mem[2091] : 
                        (N797)? mem[2107] : 
                        (N799)? mem[2123] : 
                        (N801)? mem[2139] : 
                        (N803)? mem[2155] : 
                        (N805)? mem[2171] : 
                        (N807)? mem[2187] : 
                        (N809)? mem[2203] : 
                        (N811)? mem[2219] : 
                        (N813)? mem[2235] : 
                        (N815)? mem[2251] : 
                        (N817)? mem[2267] : 
                        (N819)? mem[2283] : 
                        (N821)? mem[2299] : 
                        (N823)? mem[2315] : 
                        (N825)? mem[2331] : 
                        (N827)? mem[2347] : 
                        (N829)? mem[2363] : 
                        (N831)? mem[2379] : 
                        (N833)? mem[2395] : 
                        (N835)? mem[2411] : 
                        (N837)? mem[2427] : 
                        (N839)? mem[2443] : 
                        (N841)? mem[2459] : 
                        (N843)? mem[2475] : 
                        (N845)? mem[2491] : 
                        (N847)? mem[2507] : 
                        (N849)? mem[2523] : 
                        (N851)? mem[2539] : 
                        (N853)? mem[2555] : 
                        (N855)? mem[2571] : 
                        (N857)? mem[2587] : 
                        (N859)? mem[2603] : 
                        (N861)? mem[2619] : 
                        (N863)? mem[2635] : 
                        (N865)? mem[2651] : 
                        (N867)? mem[2667] : 
                        (N869)? mem[2683] : 
                        (N871)? mem[2699] : 
                        (N873)? mem[2715] : 
                        (N875)? mem[2731] : 
                        (N877)? mem[2747] : 
                        (N879)? mem[2763] : 
                        (N881)? mem[2779] : 
                        (N883)? mem[2795] : 
                        (N885)? mem[2811] : 
                        (N887)? mem[2827] : 
                        (N889)? mem[2843] : 
                        (N891)? mem[2859] : 
                        (N893)? mem[2875] : 
                        (N895)? mem[2891] : 
                        (N897)? mem[2907] : 
                        (N899)? mem[2923] : 
                        (N901)? mem[2939] : 
                        (N903)? mem[2955] : 
                        (N905)? mem[2971] : 
                        (N907)? mem[2987] : 
                        (N909)? mem[3003] : 
                        (N911)? mem[3019] : 
                        (N913)? mem[3035] : 
                        (N915)? mem[3051] : 
                        (N917)? mem[3067] : 
                        (N919)? mem[3083] : 
                        (N921)? mem[3099] : 
                        (N923)? mem[3115] : 
                        (N925)? mem[3131] : 
                        (N927)? mem[3147] : 
                        (N929)? mem[3163] : 
                        (N931)? mem[3179] : 
                        (N933)? mem[3195] : 
                        (N935)? mem[3211] : 
                        (N937)? mem[3227] : 
                        (N939)? mem[3243] : 
                        (N941)? mem[3259] : 
                        (N943)? mem[3275] : 
                        (N945)? mem[3291] : 
                        (N947)? mem[3307] : 
                        (N949)? mem[3323] : 
                        (N951)? mem[3339] : 
                        (N953)? mem[3355] : 
                        (N955)? mem[3371] : 
                        (N957)? mem[3387] : 
                        (N959)? mem[3403] : 
                        (N961)? mem[3419] : 
                        (N963)? mem[3435] : 
                        (N965)? mem[3451] : 
                        (N967)? mem[3467] : 
                        (N969)? mem[3483] : 
                        (N971)? mem[3499] : 
                        (N973)? mem[3515] : 
                        (N975)? mem[3531] : 
                        (N977)? mem[3547] : 
                        (N979)? mem[3563] : 
                        (N981)? mem[3579] : 
                        (N983)? mem[3595] : 
                        (N985)? mem[3611] : 
                        (N987)? mem[3627] : 
                        (N989)? mem[3643] : 
                        (N991)? mem[3659] : 
                        (N993)? mem[3675] : 
                        (N995)? mem[3691] : 
                        (N997)? mem[3707] : 
                        (N999)? mem[3723] : 
                        (N1001)? mem[3739] : 
                        (N1003)? mem[3755] : 
                        (N1005)? mem[3771] : 
                        (N1007)? mem[3787] : 
                        (N1009)? mem[3803] : 
                        (N1011)? mem[3819] : 
                        (N1013)? mem[3835] : 
                        (N1015)? mem[3851] : 
                        (N1017)? mem[3867] : 
                        (N1019)? mem[3883] : 
                        (N1021)? mem[3899] : 
                        (N1023)? mem[3915] : 
                        (N1025)? mem[3931] : 
                        (N1027)? mem[3947] : 
                        (N1029)? mem[3963] : 
                        (N1031)? mem[3979] : 
                        (N1033)? mem[3995] : 
                        (N1035)? mem[4011] : 
                        (N1037)? mem[4027] : 
                        (N1039)? mem[4043] : 
                        (N1041)? mem[4059] : 
                        (N1043)? mem[4075] : 
                        (N1045)? mem[4091] : 
                        (N536)? mem[4107] : 
                        (N538)? mem[4123] : 
                        (N540)? mem[4139] : 
                        (N542)? mem[4155] : 
                        (N544)? mem[4171] : 
                        (N546)? mem[4187] : 
                        (N548)? mem[4203] : 
                        (N550)? mem[4219] : 
                        (N552)? mem[4235] : 
                        (N554)? mem[4251] : 
                        (N556)? mem[4267] : 
                        (N558)? mem[4283] : 
                        (N560)? mem[4299] : 
                        (N562)? mem[4315] : 
                        (N564)? mem[4331] : 
                        (N566)? mem[4347] : 
                        (N568)? mem[4363] : 
                        (N570)? mem[4379] : 
                        (N572)? mem[4395] : 
                        (N574)? mem[4411] : 
                        (N576)? mem[4427] : 
                        (N578)? mem[4443] : 
                        (N580)? mem[4459] : 
                        (N582)? mem[4475] : 
                        (N584)? mem[4491] : 
                        (N586)? mem[4507] : 
                        (N588)? mem[4523] : 
                        (N590)? mem[4539] : 
                        (N592)? mem[4555] : 
                        (N594)? mem[4571] : 
                        (N596)? mem[4587] : 
                        (N598)? mem[4603] : 
                        (N600)? mem[4619] : 
                        (N602)? mem[4635] : 
                        (N604)? mem[4651] : 
                        (N606)? mem[4667] : 
                        (N608)? mem[4683] : 
                        (N610)? mem[4699] : 
                        (N612)? mem[4715] : 
                        (N614)? mem[4731] : 
                        (N616)? mem[4747] : 
                        (N618)? mem[4763] : 
                        (N620)? mem[4779] : 
                        (N622)? mem[4795] : 
                        (N624)? mem[4811] : 
                        (N626)? mem[4827] : 
                        (N628)? mem[4843] : 
                        (N630)? mem[4859] : 
                        (N632)? mem[4875] : 
                        (N634)? mem[4891] : 
                        (N636)? mem[4907] : 
                        (N638)? mem[4923] : 
                        (N640)? mem[4939] : 
                        (N642)? mem[4955] : 
                        (N644)? mem[4971] : 
                        (N646)? mem[4987] : 
                        (N648)? mem[5003] : 
                        (N650)? mem[5019] : 
                        (N652)? mem[5035] : 
                        (N654)? mem[5051] : 
                        (N656)? mem[5067] : 
                        (N658)? mem[5083] : 
                        (N660)? mem[5099] : 
                        (N662)? mem[5115] : 
                        (N664)? mem[5131] : 
                        (N666)? mem[5147] : 
                        (N668)? mem[5163] : 
                        (N670)? mem[5179] : 
                        (N672)? mem[5195] : 
                        (N674)? mem[5211] : 
                        (N676)? mem[5227] : 
                        (N678)? mem[5243] : 
                        (N680)? mem[5259] : 
                        (N682)? mem[5275] : 
                        (N684)? mem[5291] : 
                        (N686)? mem[5307] : 
                        (N688)? mem[5323] : 
                        (N690)? mem[5339] : 
                        (N692)? mem[5355] : 
                        (N694)? mem[5371] : 
                        (N696)? mem[5387] : 
                        (N698)? mem[5403] : 
                        (N700)? mem[5419] : 
                        (N702)? mem[5435] : 
                        (N704)? mem[5451] : 
                        (N706)? mem[5467] : 
                        (N708)? mem[5483] : 
                        (N710)? mem[5499] : 
                        (N712)? mem[5515] : 
                        (N714)? mem[5531] : 
                        (N716)? mem[5547] : 
                        (N718)? mem[5563] : 
                        (N720)? mem[5579] : 
                        (N722)? mem[5595] : 
                        (N724)? mem[5611] : 
                        (N726)? mem[5627] : 
                        (N728)? mem[5643] : 
                        (N730)? mem[5659] : 
                        (N732)? mem[5675] : 
                        (N734)? mem[5691] : 
                        (N736)? mem[5707] : 
                        (N738)? mem[5723] : 
                        (N740)? mem[5739] : 
                        (N742)? mem[5755] : 
                        (N744)? mem[5771] : 
                        (N746)? mem[5787] : 
                        (N748)? mem[5803] : 
                        (N750)? mem[5819] : 
                        (N752)? mem[5835] : 
                        (N754)? mem[5851] : 
                        (N756)? mem[5867] : 
                        (N758)? mem[5883] : 
                        (N760)? mem[5899] : 
                        (N762)? mem[5915] : 
                        (N764)? mem[5931] : 
                        (N766)? mem[5947] : 
                        (N768)? mem[5963] : 
                        (N770)? mem[5979] : 
                        (N772)? mem[5995] : 
                        (N774)? mem[6011] : 
                        (N776)? mem[6027] : 
                        (N778)? mem[6043] : 
                        (N780)? mem[6059] : 
                        (N782)? mem[6075] : 
                        (N784)? mem[6091] : 
                        (N786)? mem[6107] : 
                        (N788)? mem[6123] : 
                        (N790)? mem[6139] : 
                        (N792)? mem[6155] : 
                        (N794)? mem[6171] : 
                        (N796)? mem[6187] : 
                        (N798)? mem[6203] : 
                        (N800)? mem[6219] : 
                        (N802)? mem[6235] : 
                        (N804)? mem[6251] : 
                        (N806)? mem[6267] : 
                        (N808)? mem[6283] : 
                        (N810)? mem[6299] : 
                        (N812)? mem[6315] : 
                        (N814)? mem[6331] : 
                        (N816)? mem[6347] : 
                        (N818)? mem[6363] : 
                        (N820)? mem[6379] : 
                        (N822)? mem[6395] : 
                        (N824)? mem[6411] : 
                        (N826)? mem[6427] : 
                        (N828)? mem[6443] : 
                        (N830)? mem[6459] : 
                        (N832)? mem[6475] : 
                        (N834)? mem[6491] : 
                        (N836)? mem[6507] : 
                        (N838)? mem[6523] : 
                        (N840)? mem[6539] : 
                        (N842)? mem[6555] : 
                        (N844)? mem[6571] : 
                        (N846)? mem[6587] : 
                        (N848)? mem[6603] : 
                        (N850)? mem[6619] : 
                        (N852)? mem[6635] : 
                        (N854)? mem[6651] : 
                        (N856)? mem[6667] : 
                        (N858)? mem[6683] : 
                        (N860)? mem[6699] : 
                        (N862)? mem[6715] : 
                        (N864)? mem[6731] : 
                        (N866)? mem[6747] : 
                        (N868)? mem[6763] : 
                        (N870)? mem[6779] : 
                        (N872)? mem[6795] : 
                        (N874)? mem[6811] : 
                        (N876)? mem[6827] : 
                        (N878)? mem[6843] : 
                        (N880)? mem[6859] : 
                        (N882)? mem[6875] : 
                        (N884)? mem[6891] : 
                        (N886)? mem[6907] : 
                        (N888)? mem[6923] : 
                        (N890)? mem[6939] : 
                        (N892)? mem[6955] : 
                        (N894)? mem[6971] : 
                        (N896)? mem[6987] : 
                        (N898)? mem[7003] : 
                        (N900)? mem[7019] : 
                        (N902)? mem[7035] : 
                        (N904)? mem[7051] : 
                        (N906)? mem[7067] : 
                        (N908)? mem[7083] : 
                        (N910)? mem[7099] : 
                        (N912)? mem[7115] : 
                        (N914)? mem[7131] : 
                        (N916)? mem[7147] : 
                        (N918)? mem[7163] : 
                        (N920)? mem[7179] : 
                        (N922)? mem[7195] : 
                        (N924)? mem[7211] : 
                        (N926)? mem[7227] : 
                        (N928)? mem[7243] : 
                        (N930)? mem[7259] : 
                        (N932)? mem[7275] : 
                        (N934)? mem[7291] : 
                        (N936)? mem[7307] : 
                        (N938)? mem[7323] : 
                        (N940)? mem[7339] : 
                        (N942)? mem[7355] : 
                        (N944)? mem[7371] : 
                        (N946)? mem[7387] : 
                        (N948)? mem[7403] : 
                        (N950)? mem[7419] : 
                        (N952)? mem[7435] : 
                        (N954)? mem[7451] : 
                        (N956)? mem[7467] : 
                        (N958)? mem[7483] : 
                        (N960)? mem[7499] : 
                        (N962)? mem[7515] : 
                        (N964)? mem[7531] : 
                        (N966)? mem[7547] : 
                        (N968)? mem[7563] : 
                        (N970)? mem[7579] : 
                        (N972)? mem[7595] : 
                        (N974)? mem[7611] : 
                        (N976)? mem[7627] : 
                        (N978)? mem[7643] : 
                        (N980)? mem[7659] : 
                        (N982)? mem[7675] : 
                        (N984)? mem[7691] : 
                        (N986)? mem[7707] : 
                        (N988)? mem[7723] : 
                        (N990)? mem[7739] : 
                        (N992)? mem[7755] : 
                        (N994)? mem[7771] : 
                        (N996)? mem[7787] : 
                        (N998)? mem[7803] : 
                        (N1000)? mem[7819] : 
                        (N1002)? mem[7835] : 
                        (N1004)? mem[7851] : 
                        (N1006)? mem[7867] : 
                        (N1008)? mem[7883] : 
                        (N1010)? mem[7899] : 
                        (N1012)? mem[7915] : 
                        (N1014)? mem[7931] : 
                        (N1016)? mem[7947] : 
                        (N1018)? mem[7963] : 
                        (N1020)? mem[7979] : 
                        (N1022)? mem[7995] : 
                        (N1024)? mem[8011] : 
                        (N1026)? mem[8027] : 
                        (N1028)? mem[8043] : 
                        (N1030)? mem[8059] : 
                        (N1032)? mem[8075] : 
                        (N1034)? mem[8091] : 
                        (N1036)? mem[8107] : 
                        (N1038)? mem[8123] : 
                        (N1040)? mem[8139] : 
                        (N1042)? mem[8155] : 
                        (N1044)? mem[8171] : 
                        (N1046)? mem[8187] : 1'b0;
  assign r_data_o[10] = (N535)? mem[10] : 
                        (N537)? mem[26] : 
                        (N539)? mem[42] : 
                        (N541)? mem[58] : 
                        (N543)? mem[74] : 
                        (N545)? mem[90] : 
                        (N547)? mem[106] : 
                        (N549)? mem[122] : 
                        (N551)? mem[138] : 
                        (N553)? mem[154] : 
                        (N555)? mem[170] : 
                        (N557)? mem[186] : 
                        (N559)? mem[202] : 
                        (N561)? mem[218] : 
                        (N563)? mem[234] : 
                        (N565)? mem[250] : 
                        (N567)? mem[266] : 
                        (N569)? mem[282] : 
                        (N571)? mem[298] : 
                        (N573)? mem[314] : 
                        (N575)? mem[330] : 
                        (N577)? mem[346] : 
                        (N579)? mem[362] : 
                        (N581)? mem[378] : 
                        (N583)? mem[394] : 
                        (N585)? mem[410] : 
                        (N587)? mem[426] : 
                        (N589)? mem[442] : 
                        (N591)? mem[458] : 
                        (N593)? mem[474] : 
                        (N595)? mem[490] : 
                        (N597)? mem[506] : 
                        (N599)? mem[522] : 
                        (N601)? mem[538] : 
                        (N603)? mem[554] : 
                        (N605)? mem[570] : 
                        (N607)? mem[586] : 
                        (N609)? mem[602] : 
                        (N611)? mem[618] : 
                        (N613)? mem[634] : 
                        (N615)? mem[650] : 
                        (N617)? mem[666] : 
                        (N619)? mem[682] : 
                        (N621)? mem[698] : 
                        (N623)? mem[714] : 
                        (N625)? mem[730] : 
                        (N627)? mem[746] : 
                        (N629)? mem[762] : 
                        (N631)? mem[778] : 
                        (N633)? mem[794] : 
                        (N635)? mem[810] : 
                        (N637)? mem[826] : 
                        (N639)? mem[842] : 
                        (N641)? mem[858] : 
                        (N643)? mem[874] : 
                        (N645)? mem[890] : 
                        (N647)? mem[906] : 
                        (N649)? mem[922] : 
                        (N651)? mem[938] : 
                        (N653)? mem[954] : 
                        (N655)? mem[970] : 
                        (N657)? mem[986] : 
                        (N659)? mem[1002] : 
                        (N661)? mem[1018] : 
                        (N663)? mem[1034] : 
                        (N665)? mem[1050] : 
                        (N667)? mem[1066] : 
                        (N669)? mem[1082] : 
                        (N671)? mem[1098] : 
                        (N673)? mem[1114] : 
                        (N675)? mem[1130] : 
                        (N677)? mem[1146] : 
                        (N679)? mem[1162] : 
                        (N681)? mem[1178] : 
                        (N683)? mem[1194] : 
                        (N685)? mem[1210] : 
                        (N687)? mem[1226] : 
                        (N689)? mem[1242] : 
                        (N691)? mem[1258] : 
                        (N693)? mem[1274] : 
                        (N695)? mem[1290] : 
                        (N697)? mem[1306] : 
                        (N699)? mem[1322] : 
                        (N701)? mem[1338] : 
                        (N703)? mem[1354] : 
                        (N705)? mem[1370] : 
                        (N707)? mem[1386] : 
                        (N709)? mem[1402] : 
                        (N711)? mem[1418] : 
                        (N713)? mem[1434] : 
                        (N715)? mem[1450] : 
                        (N717)? mem[1466] : 
                        (N719)? mem[1482] : 
                        (N721)? mem[1498] : 
                        (N723)? mem[1514] : 
                        (N725)? mem[1530] : 
                        (N727)? mem[1546] : 
                        (N729)? mem[1562] : 
                        (N731)? mem[1578] : 
                        (N733)? mem[1594] : 
                        (N735)? mem[1610] : 
                        (N737)? mem[1626] : 
                        (N739)? mem[1642] : 
                        (N741)? mem[1658] : 
                        (N743)? mem[1674] : 
                        (N745)? mem[1690] : 
                        (N747)? mem[1706] : 
                        (N749)? mem[1722] : 
                        (N751)? mem[1738] : 
                        (N753)? mem[1754] : 
                        (N755)? mem[1770] : 
                        (N757)? mem[1786] : 
                        (N759)? mem[1802] : 
                        (N761)? mem[1818] : 
                        (N763)? mem[1834] : 
                        (N765)? mem[1850] : 
                        (N767)? mem[1866] : 
                        (N769)? mem[1882] : 
                        (N771)? mem[1898] : 
                        (N773)? mem[1914] : 
                        (N775)? mem[1930] : 
                        (N777)? mem[1946] : 
                        (N779)? mem[1962] : 
                        (N781)? mem[1978] : 
                        (N783)? mem[1994] : 
                        (N785)? mem[2010] : 
                        (N787)? mem[2026] : 
                        (N789)? mem[2042] : 
                        (N791)? mem[2058] : 
                        (N793)? mem[2074] : 
                        (N795)? mem[2090] : 
                        (N797)? mem[2106] : 
                        (N799)? mem[2122] : 
                        (N801)? mem[2138] : 
                        (N803)? mem[2154] : 
                        (N805)? mem[2170] : 
                        (N807)? mem[2186] : 
                        (N809)? mem[2202] : 
                        (N811)? mem[2218] : 
                        (N813)? mem[2234] : 
                        (N815)? mem[2250] : 
                        (N817)? mem[2266] : 
                        (N819)? mem[2282] : 
                        (N821)? mem[2298] : 
                        (N823)? mem[2314] : 
                        (N825)? mem[2330] : 
                        (N827)? mem[2346] : 
                        (N829)? mem[2362] : 
                        (N831)? mem[2378] : 
                        (N833)? mem[2394] : 
                        (N835)? mem[2410] : 
                        (N837)? mem[2426] : 
                        (N839)? mem[2442] : 
                        (N841)? mem[2458] : 
                        (N843)? mem[2474] : 
                        (N845)? mem[2490] : 
                        (N847)? mem[2506] : 
                        (N849)? mem[2522] : 
                        (N851)? mem[2538] : 
                        (N853)? mem[2554] : 
                        (N855)? mem[2570] : 
                        (N857)? mem[2586] : 
                        (N859)? mem[2602] : 
                        (N861)? mem[2618] : 
                        (N863)? mem[2634] : 
                        (N865)? mem[2650] : 
                        (N867)? mem[2666] : 
                        (N869)? mem[2682] : 
                        (N871)? mem[2698] : 
                        (N873)? mem[2714] : 
                        (N875)? mem[2730] : 
                        (N877)? mem[2746] : 
                        (N879)? mem[2762] : 
                        (N881)? mem[2778] : 
                        (N883)? mem[2794] : 
                        (N885)? mem[2810] : 
                        (N887)? mem[2826] : 
                        (N889)? mem[2842] : 
                        (N891)? mem[2858] : 
                        (N893)? mem[2874] : 
                        (N895)? mem[2890] : 
                        (N897)? mem[2906] : 
                        (N899)? mem[2922] : 
                        (N901)? mem[2938] : 
                        (N903)? mem[2954] : 
                        (N905)? mem[2970] : 
                        (N907)? mem[2986] : 
                        (N909)? mem[3002] : 
                        (N911)? mem[3018] : 
                        (N913)? mem[3034] : 
                        (N915)? mem[3050] : 
                        (N917)? mem[3066] : 
                        (N919)? mem[3082] : 
                        (N921)? mem[3098] : 
                        (N923)? mem[3114] : 
                        (N925)? mem[3130] : 
                        (N927)? mem[3146] : 
                        (N929)? mem[3162] : 
                        (N931)? mem[3178] : 
                        (N933)? mem[3194] : 
                        (N935)? mem[3210] : 
                        (N937)? mem[3226] : 
                        (N939)? mem[3242] : 
                        (N941)? mem[3258] : 
                        (N943)? mem[3274] : 
                        (N945)? mem[3290] : 
                        (N947)? mem[3306] : 
                        (N949)? mem[3322] : 
                        (N951)? mem[3338] : 
                        (N953)? mem[3354] : 
                        (N955)? mem[3370] : 
                        (N957)? mem[3386] : 
                        (N959)? mem[3402] : 
                        (N961)? mem[3418] : 
                        (N963)? mem[3434] : 
                        (N965)? mem[3450] : 
                        (N967)? mem[3466] : 
                        (N969)? mem[3482] : 
                        (N971)? mem[3498] : 
                        (N973)? mem[3514] : 
                        (N975)? mem[3530] : 
                        (N977)? mem[3546] : 
                        (N979)? mem[3562] : 
                        (N981)? mem[3578] : 
                        (N983)? mem[3594] : 
                        (N985)? mem[3610] : 
                        (N987)? mem[3626] : 
                        (N989)? mem[3642] : 
                        (N991)? mem[3658] : 
                        (N993)? mem[3674] : 
                        (N995)? mem[3690] : 
                        (N997)? mem[3706] : 
                        (N999)? mem[3722] : 
                        (N1001)? mem[3738] : 
                        (N1003)? mem[3754] : 
                        (N1005)? mem[3770] : 
                        (N1007)? mem[3786] : 
                        (N1009)? mem[3802] : 
                        (N1011)? mem[3818] : 
                        (N1013)? mem[3834] : 
                        (N1015)? mem[3850] : 
                        (N1017)? mem[3866] : 
                        (N1019)? mem[3882] : 
                        (N1021)? mem[3898] : 
                        (N1023)? mem[3914] : 
                        (N1025)? mem[3930] : 
                        (N1027)? mem[3946] : 
                        (N1029)? mem[3962] : 
                        (N1031)? mem[3978] : 
                        (N1033)? mem[3994] : 
                        (N1035)? mem[4010] : 
                        (N1037)? mem[4026] : 
                        (N1039)? mem[4042] : 
                        (N1041)? mem[4058] : 
                        (N1043)? mem[4074] : 
                        (N1045)? mem[4090] : 
                        (N536)? mem[4106] : 
                        (N538)? mem[4122] : 
                        (N540)? mem[4138] : 
                        (N542)? mem[4154] : 
                        (N544)? mem[4170] : 
                        (N546)? mem[4186] : 
                        (N548)? mem[4202] : 
                        (N550)? mem[4218] : 
                        (N552)? mem[4234] : 
                        (N554)? mem[4250] : 
                        (N556)? mem[4266] : 
                        (N558)? mem[4282] : 
                        (N560)? mem[4298] : 
                        (N562)? mem[4314] : 
                        (N564)? mem[4330] : 
                        (N566)? mem[4346] : 
                        (N568)? mem[4362] : 
                        (N570)? mem[4378] : 
                        (N572)? mem[4394] : 
                        (N574)? mem[4410] : 
                        (N576)? mem[4426] : 
                        (N578)? mem[4442] : 
                        (N580)? mem[4458] : 
                        (N582)? mem[4474] : 
                        (N584)? mem[4490] : 
                        (N586)? mem[4506] : 
                        (N588)? mem[4522] : 
                        (N590)? mem[4538] : 
                        (N592)? mem[4554] : 
                        (N594)? mem[4570] : 
                        (N596)? mem[4586] : 
                        (N598)? mem[4602] : 
                        (N600)? mem[4618] : 
                        (N602)? mem[4634] : 
                        (N604)? mem[4650] : 
                        (N606)? mem[4666] : 
                        (N608)? mem[4682] : 
                        (N610)? mem[4698] : 
                        (N612)? mem[4714] : 
                        (N614)? mem[4730] : 
                        (N616)? mem[4746] : 
                        (N618)? mem[4762] : 
                        (N620)? mem[4778] : 
                        (N622)? mem[4794] : 
                        (N624)? mem[4810] : 
                        (N626)? mem[4826] : 
                        (N628)? mem[4842] : 
                        (N630)? mem[4858] : 
                        (N632)? mem[4874] : 
                        (N634)? mem[4890] : 
                        (N636)? mem[4906] : 
                        (N638)? mem[4922] : 
                        (N640)? mem[4938] : 
                        (N642)? mem[4954] : 
                        (N644)? mem[4970] : 
                        (N646)? mem[4986] : 
                        (N648)? mem[5002] : 
                        (N650)? mem[5018] : 
                        (N652)? mem[5034] : 
                        (N654)? mem[5050] : 
                        (N656)? mem[5066] : 
                        (N658)? mem[5082] : 
                        (N660)? mem[5098] : 
                        (N662)? mem[5114] : 
                        (N664)? mem[5130] : 
                        (N666)? mem[5146] : 
                        (N668)? mem[5162] : 
                        (N670)? mem[5178] : 
                        (N672)? mem[5194] : 
                        (N674)? mem[5210] : 
                        (N676)? mem[5226] : 
                        (N678)? mem[5242] : 
                        (N680)? mem[5258] : 
                        (N682)? mem[5274] : 
                        (N684)? mem[5290] : 
                        (N686)? mem[5306] : 
                        (N688)? mem[5322] : 
                        (N690)? mem[5338] : 
                        (N692)? mem[5354] : 
                        (N694)? mem[5370] : 
                        (N696)? mem[5386] : 
                        (N698)? mem[5402] : 
                        (N700)? mem[5418] : 
                        (N702)? mem[5434] : 
                        (N704)? mem[5450] : 
                        (N706)? mem[5466] : 
                        (N708)? mem[5482] : 
                        (N710)? mem[5498] : 
                        (N712)? mem[5514] : 
                        (N714)? mem[5530] : 
                        (N716)? mem[5546] : 
                        (N718)? mem[5562] : 
                        (N720)? mem[5578] : 
                        (N722)? mem[5594] : 
                        (N724)? mem[5610] : 
                        (N726)? mem[5626] : 
                        (N728)? mem[5642] : 
                        (N730)? mem[5658] : 
                        (N732)? mem[5674] : 
                        (N734)? mem[5690] : 
                        (N736)? mem[5706] : 
                        (N738)? mem[5722] : 
                        (N740)? mem[5738] : 
                        (N742)? mem[5754] : 
                        (N744)? mem[5770] : 
                        (N746)? mem[5786] : 
                        (N748)? mem[5802] : 
                        (N750)? mem[5818] : 
                        (N752)? mem[5834] : 
                        (N754)? mem[5850] : 
                        (N756)? mem[5866] : 
                        (N758)? mem[5882] : 
                        (N760)? mem[5898] : 
                        (N762)? mem[5914] : 
                        (N764)? mem[5930] : 
                        (N766)? mem[5946] : 
                        (N768)? mem[5962] : 
                        (N770)? mem[5978] : 
                        (N772)? mem[5994] : 
                        (N774)? mem[6010] : 
                        (N776)? mem[6026] : 
                        (N778)? mem[6042] : 
                        (N780)? mem[6058] : 
                        (N782)? mem[6074] : 
                        (N784)? mem[6090] : 
                        (N786)? mem[6106] : 
                        (N788)? mem[6122] : 
                        (N790)? mem[6138] : 
                        (N792)? mem[6154] : 
                        (N794)? mem[6170] : 
                        (N796)? mem[6186] : 
                        (N798)? mem[6202] : 
                        (N800)? mem[6218] : 
                        (N802)? mem[6234] : 
                        (N804)? mem[6250] : 
                        (N806)? mem[6266] : 
                        (N808)? mem[6282] : 
                        (N810)? mem[6298] : 
                        (N812)? mem[6314] : 
                        (N814)? mem[6330] : 
                        (N816)? mem[6346] : 
                        (N818)? mem[6362] : 
                        (N820)? mem[6378] : 
                        (N822)? mem[6394] : 
                        (N824)? mem[6410] : 
                        (N826)? mem[6426] : 
                        (N828)? mem[6442] : 
                        (N830)? mem[6458] : 
                        (N832)? mem[6474] : 
                        (N834)? mem[6490] : 
                        (N836)? mem[6506] : 
                        (N838)? mem[6522] : 
                        (N840)? mem[6538] : 
                        (N842)? mem[6554] : 
                        (N844)? mem[6570] : 
                        (N846)? mem[6586] : 
                        (N848)? mem[6602] : 
                        (N850)? mem[6618] : 
                        (N852)? mem[6634] : 
                        (N854)? mem[6650] : 
                        (N856)? mem[6666] : 
                        (N858)? mem[6682] : 
                        (N860)? mem[6698] : 
                        (N862)? mem[6714] : 
                        (N864)? mem[6730] : 
                        (N866)? mem[6746] : 
                        (N868)? mem[6762] : 
                        (N870)? mem[6778] : 
                        (N872)? mem[6794] : 
                        (N874)? mem[6810] : 
                        (N876)? mem[6826] : 
                        (N878)? mem[6842] : 
                        (N880)? mem[6858] : 
                        (N882)? mem[6874] : 
                        (N884)? mem[6890] : 
                        (N886)? mem[6906] : 
                        (N888)? mem[6922] : 
                        (N890)? mem[6938] : 
                        (N892)? mem[6954] : 
                        (N894)? mem[6970] : 
                        (N896)? mem[6986] : 
                        (N898)? mem[7002] : 
                        (N900)? mem[7018] : 
                        (N902)? mem[7034] : 
                        (N904)? mem[7050] : 
                        (N906)? mem[7066] : 
                        (N908)? mem[7082] : 
                        (N910)? mem[7098] : 
                        (N912)? mem[7114] : 
                        (N914)? mem[7130] : 
                        (N916)? mem[7146] : 
                        (N918)? mem[7162] : 
                        (N920)? mem[7178] : 
                        (N922)? mem[7194] : 
                        (N924)? mem[7210] : 
                        (N926)? mem[7226] : 
                        (N928)? mem[7242] : 
                        (N930)? mem[7258] : 
                        (N932)? mem[7274] : 
                        (N934)? mem[7290] : 
                        (N936)? mem[7306] : 
                        (N938)? mem[7322] : 
                        (N940)? mem[7338] : 
                        (N942)? mem[7354] : 
                        (N944)? mem[7370] : 
                        (N946)? mem[7386] : 
                        (N948)? mem[7402] : 
                        (N950)? mem[7418] : 
                        (N952)? mem[7434] : 
                        (N954)? mem[7450] : 
                        (N956)? mem[7466] : 
                        (N958)? mem[7482] : 
                        (N960)? mem[7498] : 
                        (N962)? mem[7514] : 
                        (N964)? mem[7530] : 
                        (N966)? mem[7546] : 
                        (N968)? mem[7562] : 
                        (N970)? mem[7578] : 
                        (N972)? mem[7594] : 
                        (N974)? mem[7610] : 
                        (N976)? mem[7626] : 
                        (N978)? mem[7642] : 
                        (N980)? mem[7658] : 
                        (N982)? mem[7674] : 
                        (N984)? mem[7690] : 
                        (N986)? mem[7706] : 
                        (N988)? mem[7722] : 
                        (N990)? mem[7738] : 
                        (N992)? mem[7754] : 
                        (N994)? mem[7770] : 
                        (N996)? mem[7786] : 
                        (N998)? mem[7802] : 
                        (N1000)? mem[7818] : 
                        (N1002)? mem[7834] : 
                        (N1004)? mem[7850] : 
                        (N1006)? mem[7866] : 
                        (N1008)? mem[7882] : 
                        (N1010)? mem[7898] : 
                        (N1012)? mem[7914] : 
                        (N1014)? mem[7930] : 
                        (N1016)? mem[7946] : 
                        (N1018)? mem[7962] : 
                        (N1020)? mem[7978] : 
                        (N1022)? mem[7994] : 
                        (N1024)? mem[8010] : 
                        (N1026)? mem[8026] : 
                        (N1028)? mem[8042] : 
                        (N1030)? mem[8058] : 
                        (N1032)? mem[8074] : 
                        (N1034)? mem[8090] : 
                        (N1036)? mem[8106] : 
                        (N1038)? mem[8122] : 
                        (N1040)? mem[8138] : 
                        (N1042)? mem[8154] : 
                        (N1044)? mem[8170] : 
                        (N1046)? mem[8186] : 1'b0;
  assign r_data_o[9] = (N535)? mem[9] : 
                       (N537)? mem[25] : 
                       (N539)? mem[41] : 
                       (N541)? mem[57] : 
                       (N543)? mem[73] : 
                       (N545)? mem[89] : 
                       (N547)? mem[105] : 
                       (N549)? mem[121] : 
                       (N551)? mem[137] : 
                       (N553)? mem[153] : 
                       (N555)? mem[169] : 
                       (N557)? mem[185] : 
                       (N559)? mem[201] : 
                       (N561)? mem[217] : 
                       (N563)? mem[233] : 
                       (N565)? mem[249] : 
                       (N567)? mem[265] : 
                       (N569)? mem[281] : 
                       (N571)? mem[297] : 
                       (N573)? mem[313] : 
                       (N575)? mem[329] : 
                       (N577)? mem[345] : 
                       (N579)? mem[361] : 
                       (N581)? mem[377] : 
                       (N583)? mem[393] : 
                       (N585)? mem[409] : 
                       (N587)? mem[425] : 
                       (N589)? mem[441] : 
                       (N591)? mem[457] : 
                       (N593)? mem[473] : 
                       (N595)? mem[489] : 
                       (N597)? mem[505] : 
                       (N599)? mem[521] : 
                       (N601)? mem[537] : 
                       (N603)? mem[553] : 
                       (N605)? mem[569] : 
                       (N607)? mem[585] : 
                       (N609)? mem[601] : 
                       (N611)? mem[617] : 
                       (N613)? mem[633] : 
                       (N615)? mem[649] : 
                       (N617)? mem[665] : 
                       (N619)? mem[681] : 
                       (N621)? mem[697] : 
                       (N623)? mem[713] : 
                       (N625)? mem[729] : 
                       (N627)? mem[745] : 
                       (N629)? mem[761] : 
                       (N631)? mem[777] : 
                       (N633)? mem[793] : 
                       (N635)? mem[809] : 
                       (N637)? mem[825] : 
                       (N639)? mem[841] : 
                       (N641)? mem[857] : 
                       (N643)? mem[873] : 
                       (N645)? mem[889] : 
                       (N647)? mem[905] : 
                       (N649)? mem[921] : 
                       (N651)? mem[937] : 
                       (N653)? mem[953] : 
                       (N655)? mem[969] : 
                       (N657)? mem[985] : 
                       (N659)? mem[1001] : 
                       (N661)? mem[1017] : 
                       (N663)? mem[1033] : 
                       (N665)? mem[1049] : 
                       (N667)? mem[1065] : 
                       (N669)? mem[1081] : 
                       (N671)? mem[1097] : 
                       (N673)? mem[1113] : 
                       (N675)? mem[1129] : 
                       (N677)? mem[1145] : 
                       (N679)? mem[1161] : 
                       (N681)? mem[1177] : 
                       (N683)? mem[1193] : 
                       (N685)? mem[1209] : 
                       (N687)? mem[1225] : 
                       (N689)? mem[1241] : 
                       (N691)? mem[1257] : 
                       (N693)? mem[1273] : 
                       (N695)? mem[1289] : 
                       (N697)? mem[1305] : 
                       (N699)? mem[1321] : 
                       (N701)? mem[1337] : 
                       (N703)? mem[1353] : 
                       (N705)? mem[1369] : 
                       (N707)? mem[1385] : 
                       (N709)? mem[1401] : 
                       (N711)? mem[1417] : 
                       (N713)? mem[1433] : 
                       (N715)? mem[1449] : 
                       (N717)? mem[1465] : 
                       (N719)? mem[1481] : 
                       (N721)? mem[1497] : 
                       (N723)? mem[1513] : 
                       (N725)? mem[1529] : 
                       (N727)? mem[1545] : 
                       (N729)? mem[1561] : 
                       (N731)? mem[1577] : 
                       (N733)? mem[1593] : 
                       (N735)? mem[1609] : 
                       (N737)? mem[1625] : 
                       (N739)? mem[1641] : 
                       (N741)? mem[1657] : 
                       (N743)? mem[1673] : 
                       (N745)? mem[1689] : 
                       (N747)? mem[1705] : 
                       (N749)? mem[1721] : 
                       (N751)? mem[1737] : 
                       (N753)? mem[1753] : 
                       (N755)? mem[1769] : 
                       (N757)? mem[1785] : 
                       (N759)? mem[1801] : 
                       (N761)? mem[1817] : 
                       (N763)? mem[1833] : 
                       (N765)? mem[1849] : 
                       (N767)? mem[1865] : 
                       (N769)? mem[1881] : 
                       (N771)? mem[1897] : 
                       (N773)? mem[1913] : 
                       (N775)? mem[1929] : 
                       (N777)? mem[1945] : 
                       (N779)? mem[1961] : 
                       (N781)? mem[1977] : 
                       (N783)? mem[1993] : 
                       (N785)? mem[2009] : 
                       (N787)? mem[2025] : 
                       (N789)? mem[2041] : 
                       (N791)? mem[2057] : 
                       (N793)? mem[2073] : 
                       (N795)? mem[2089] : 
                       (N797)? mem[2105] : 
                       (N799)? mem[2121] : 
                       (N801)? mem[2137] : 
                       (N803)? mem[2153] : 
                       (N805)? mem[2169] : 
                       (N807)? mem[2185] : 
                       (N809)? mem[2201] : 
                       (N811)? mem[2217] : 
                       (N813)? mem[2233] : 
                       (N815)? mem[2249] : 
                       (N817)? mem[2265] : 
                       (N819)? mem[2281] : 
                       (N821)? mem[2297] : 
                       (N823)? mem[2313] : 
                       (N825)? mem[2329] : 
                       (N827)? mem[2345] : 
                       (N829)? mem[2361] : 
                       (N831)? mem[2377] : 
                       (N833)? mem[2393] : 
                       (N835)? mem[2409] : 
                       (N837)? mem[2425] : 
                       (N839)? mem[2441] : 
                       (N841)? mem[2457] : 
                       (N843)? mem[2473] : 
                       (N845)? mem[2489] : 
                       (N847)? mem[2505] : 
                       (N849)? mem[2521] : 
                       (N851)? mem[2537] : 
                       (N853)? mem[2553] : 
                       (N855)? mem[2569] : 
                       (N857)? mem[2585] : 
                       (N859)? mem[2601] : 
                       (N861)? mem[2617] : 
                       (N863)? mem[2633] : 
                       (N865)? mem[2649] : 
                       (N867)? mem[2665] : 
                       (N869)? mem[2681] : 
                       (N871)? mem[2697] : 
                       (N873)? mem[2713] : 
                       (N875)? mem[2729] : 
                       (N877)? mem[2745] : 
                       (N879)? mem[2761] : 
                       (N881)? mem[2777] : 
                       (N883)? mem[2793] : 
                       (N885)? mem[2809] : 
                       (N887)? mem[2825] : 
                       (N889)? mem[2841] : 
                       (N891)? mem[2857] : 
                       (N893)? mem[2873] : 
                       (N895)? mem[2889] : 
                       (N897)? mem[2905] : 
                       (N899)? mem[2921] : 
                       (N901)? mem[2937] : 
                       (N903)? mem[2953] : 
                       (N905)? mem[2969] : 
                       (N907)? mem[2985] : 
                       (N909)? mem[3001] : 
                       (N911)? mem[3017] : 
                       (N913)? mem[3033] : 
                       (N915)? mem[3049] : 
                       (N917)? mem[3065] : 
                       (N919)? mem[3081] : 
                       (N921)? mem[3097] : 
                       (N923)? mem[3113] : 
                       (N925)? mem[3129] : 
                       (N927)? mem[3145] : 
                       (N929)? mem[3161] : 
                       (N931)? mem[3177] : 
                       (N933)? mem[3193] : 
                       (N935)? mem[3209] : 
                       (N937)? mem[3225] : 
                       (N939)? mem[3241] : 
                       (N941)? mem[3257] : 
                       (N943)? mem[3273] : 
                       (N945)? mem[3289] : 
                       (N947)? mem[3305] : 
                       (N949)? mem[3321] : 
                       (N951)? mem[3337] : 
                       (N953)? mem[3353] : 
                       (N955)? mem[3369] : 
                       (N957)? mem[3385] : 
                       (N959)? mem[3401] : 
                       (N961)? mem[3417] : 
                       (N963)? mem[3433] : 
                       (N965)? mem[3449] : 
                       (N967)? mem[3465] : 
                       (N969)? mem[3481] : 
                       (N971)? mem[3497] : 
                       (N973)? mem[3513] : 
                       (N975)? mem[3529] : 
                       (N977)? mem[3545] : 
                       (N979)? mem[3561] : 
                       (N981)? mem[3577] : 
                       (N983)? mem[3593] : 
                       (N985)? mem[3609] : 
                       (N987)? mem[3625] : 
                       (N989)? mem[3641] : 
                       (N991)? mem[3657] : 
                       (N993)? mem[3673] : 
                       (N995)? mem[3689] : 
                       (N997)? mem[3705] : 
                       (N999)? mem[3721] : 
                       (N1001)? mem[3737] : 
                       (N1003)? mem[3753] : 
                       (N1005)? mem[3769] : 
                       (N1007)? mem[3785] : 
                       (N1009)? mem[3801] : 
                       (N1011)? mem[3817] : 
                       (N1013)? mem[3833] : 
                       (N1015)? mem[3849] : 
                       (N1017)? mem[3865] : 
                       (N1019)? mem[3881] : 
                       (N1021)? mem[3897] : 
                       (N1023)? mem[3913] : 
                       (N1025)? mem[3929] : 
                       (N1027)? mem[3945] : 
                       (N1029)? mem[3961] : 
                       (N1031)? mem[3977] : 
                       (N1033)? mem[3993] : 
                       (N1035)? mem[4009] : 
                       (N1037)? mem[4025] : 
                       (N1039)? mem[4041] : 
                       (N1041)? mem[4057] : 
                       (N1043)? mem[4073] : 
                       (N1045)? mem[4089] : 
                       (N536)? mem[4105] : 
                       (N538)? mem[4121] : 
                       (N540)? mem[4137] : 
                       (N542)? mem[4153] : 
                       (N544)? mem[4169] : 
                       (N546)? mem[4185] : 
                       (N548)? mem[4201] : 
                       (N550)? mem[4217] : 
                       (N552)? mem[4233] : 
                       (N554)? mem[4249] : 
                       (N556)? mem[4265] : 
                       (N558)? mem[4281] : 
                       (N560)? mem[4297] : 
                       (N562)? mem[4313] : 
                       (N564)? mem[4329] : 
                       (N566)? mem[4345] : 
                       (N568)? mem[4361] : 
                       (N570)? mem[4377] : 
                       (N572)? mem[4393] : 
                       (N574)? mem[4409] : 
                       (N576)? mem[4425] : 
                       (N578)? mem[4441] : 
                       (N580)? mem[4457] : 
                       (N582)? mem[4473] : 
                       (N584)? mem[4489] : 
                       (N586)? mem[4505] : 
                       (N588)? mem[4521] : 
                       (N590)? mem[4537] : 
                       (N592)? mem[4553] : 
                       (N594)? mem[4569] : 
                       (N596)? mem[4585] : 
                       (N598)? mem[4601] : 
                       (N600)? mem[4617] : 
                       (N602)? mem[4633] : 
                       (N604)? mem[4649] : 
                       (N606)? mem[4665] : 
                       (N608)? mem[4681] : 
                       (N610)? mem[4697] : 
                       (N612)? mem[4713] : 
                       (N614)? mem[4729] : 
                       (N616)? mem[4745] : 
                       (N618)? mem[4761] : 
                       (N620)? mem[4777] : 
                       (N622)? mem[4793] : 
                       (N624)? mem[4809] : 
                       (N626)? mem[4825] : 
                       (N628)? mem[4841] : 
                       (N630)? mem[4857] : 
                       (N632)? mem[4873] : 
                       (N634)? mem[4889] : 
                       (N636)? mem[4905] : 
                       (N638)? mem[4921] : 
                       (N640)? mem[4937] : 
                       (N642)? mem[4953] : 
                       (N644)? mem[4969] : 
                       (N646)? mem[4985] : 
                       (N648)? mem[5001] : 
                       (N650)? mem[5017] : 
                       (N652)? mem[5033] : 
                       (N654)? mem[5049] : 
                       (N656)? mem[5065] : 
                       (N658)? mem[5081] : 
                       (N660)? mem[5097] : 
                       (N662)? mem[5113] : 
                       (N664)? mem[5129] : 
                       (N666)? mem[5145] : 
                       (N668)? mem[5161] : 
                       (N670)? mem[5177] : 
                       (N672)? mem[5193] : 
                       (N674)? mem[5209] : 
                       (N676)? mem[5225] : 
                       (N678)? mem[5241] : 
                       (N680)? mem[5257] : 
                       (N682)? mem[5273] : 
                       (N684)? mem[5289] : 
                       (N686)? mem[5305] : 
                       (N688)? mem[5321] : 
                       (N690)? mem[5337] : 
                       (N692)? mem[5353] : 
                       (N694)? mem[5369] : 
                       (N696)? mem[5385] : 
                       (N698)? mem[5401] : 
                       (N700)? mem[5417] : 
                       (N702)? mem[5433] : 
                       (N704)? mem[5449] : 
                       (N706)? mem[5465] : 
                       (N708)? mem[5481] : 
                       (N710)? mem[5497] : 
                       (N712)? mem[5513] : 
                       (N714)? mem[5529] : 
                       (N716)? mem[5545] : 
                       (N718)? mem[5561] : 
                       (N720)? mem[5577] : 
                       (N722)? mem[5593] : 
                       (N724)? mem[5609] : 
                       (N726)? mem[5625] : 
                       (N728)? mem[5641] : 
                       (N730)? mem[5657] : 
                       (N732)? mem[5673] : 
                       (N734)? mem[5689] : 
                       (N736)? mem[5705] : 
                       (N738)? mem[5721] : 
                       (N740)? mem[5737] : 
                       (N742)? mem[5753] : 
                       (N744)? mem[5769] : 
                       (N746)? mem[5785] : 
                       (N748)? mem[5801] : 
                       (N750)? mem[5817] : 
                       (N752)? mem[5833] : 
                       (N754)? mem[5849] : 
                       (N756)? mem[5865] : 
                       (N758)? mem[5881] : 
                       (N760)? mem[5897] : 
                       (N762)? mem[5913] : 
                       (N764)? mem[5929] : 
                       (N766)? mem[5945] : 
                       (N768)? mem[5961] : 
                       (N770)? mem[5977] : 
                       (N772)? mem[5993] : 
                       (N774)? mem[6009] : 
                       (N776)? mem[6025] : 
                       (N778)? mem[6041] : 
                       (N780)? mem[6057] : 
                       (N782)? mem[6073] : 
                       (N784)? mem[6089] : 
                       (N786)? mem[6105] : 
                       (N788)? mem[6121] : 
                       (N790)? mem[6137] : 
                       (N792)? mem[6153] : 
                       (N794)? mem[6169] : 
                       (N796)? mem[6185] : 
                       (N798)? mem[6201] : 
                       (N800)? mem[6217] : 
                       (N802)? mem[6233] : 
                       (N804)? mem[6249] : 
                       (N806)? mem[6265] : 
                       (N808)? mem[6281] : 
                       (N810)? mem[6297] : 
                       (N812)? mem[6313] : 
                       (N814)? mem[6329] : 
                       (N816)? mem[6345] : 
                       (N818)? mem[6361] : 
                       (N820)? mem[6377] : 
                       (N822)? mem[6393] : 
                       (N824)? mem[6409] : 
                       (N826)? mem[6425] : 
                       (N828)? mem[6441] : 
                       (N830)? mem[6457] : 
                       (N832)? mem[6473] : 
                       (N834)? mem[6489] : 
                       (N836)? mem[6505] : 
                       (N838)? mem[6521] : 
                       (N840)? mem[6537] : 
                       (N842)? mem[6553] : 
                       (N844)? mem[6569] : 
                       (N846)? mem[6585] : 
                       (N848)? mem[6601] : 
                       (N850)? mem[6617] : 
                       (N852)? mem[6633] : 
                       (N854)? mem[6649] : 
                       (N856)? mem[6665] : 
                       (N858)? mem[6681] : 
                       (N860)? mem[6697] : 
                       (N862)? mem[6713] : 
                       (N864)? mem[6729] : 
                       (N866)? mem[6745] : 
                       (N868)? mem[6761] : 
                       (N870)? mem[6777] : 
                       (N872)? mem[6793] : 
                       (N874)? mem[6809] : 
                       (N876)? mem[6825] : 
                       (N878)? mem[6841] : 
                       (N880)? mem[6857] : 
                       (N882)? mem[6873] : 
                       (N884)? mem[6889] : 
                       (N886)? mem[6905] : 
                       (N888)? mem[6921] : 
                       (N890)? mem[6937] : 
                       (N892)? mem[6953] : 
                       (N894)? mem[6969] : 
                       (N896)? mem[6985] : 
                       (N898)? mem[7001] : 
                       (N900)? mem[7017] : 
                       (N902)? mem[7033] : 
                       (N904)? mem[7049] : 
                       (N906)? mem[7065] : 
                       (N908)? mem[7081] : 
                       (N910)? mem[7097] : 
                       (N912)? mem[7113] : 
                       (N914)? mem[7129] : 
                       (N916)? mem[7145] : 
                       (N918)? mem[7161] : 
                       (N920)? mem[7177] : 
                       (N922)? mem[7193] : 
                       (N924)? mem[7209] : 
                       (N926)? mem[7225] : 
                       (N928)? mem[7241] : 
                       (N930)? mem[7257] : 
                       (N932)? mem[7273] : 
                       (N934)? mem[7289] : 
                       (N936)? mem[7305] : 
                       (N938)? mem[7321] : 
                       (N940)? mem[7337] : 
                       (N942)? mem[7353] : 
                       (N944)? mem[7369] : 
                       (N946)? mem[7385] : 
                       (N948)? mem[7401] : 
                       (N950)? mem[7417] : 
                       (N952)? mem[7433] : 
                       (N954)? mem[7449] : 
                       (N956)? mem[7465] : 
                       (N958)? mem[7481] : 
                       (N960)? mem[7497] : 
                       (N962)? mem[7513] : 
                       (N964)? mem[7529] : 
                       (N966)? mem[7545] : 
                       (N968)? mem[7561] : 
                       (N970)? mem[7577] : 
                       (N972)? mem[7593] : 
                       (N974)? mem[7609] : 
                       (N976)? mem[7625] : 
                       (N978)? mem[7641] : 
                       (N980)? mem[7657] : 
                       (N982)? mem[7673] : 
                       (N984)? mem[7689] : 
                       (N986)? mem[7705] : 
                       (N988)? mem[7721] : 
                       (N990)? mem[7737] : 
                       (N992)? mem[7753] : 
                       (N994)? mem[7769] : 
                       (N996)? mem[7785] : 
                       (N998)? mem[7801] : 
                       (N1000)? mem[7817] : 
                       (N1002)? mem[7833] : 
                       (N1004)? mem[7849] : 
                       (N1006)? mem[7865] : 
                       (N1008)? mem[7881] : 
                       (N1010)? mem[7897] : 
                       (N1012)? mem[7913] : 
                       (N1014)? mem[7929] : 
                       (N1016)? mem[7945] : 
                       (N1018)? mem[7961] : 
                       (N1020)? mem[7977] : 
                       (N1022)? mem[7993] : 
                       (N1024)? mem[8009] : 
                       (N1026)? mem[8025] : 
                       (N1028)? mem[8041] : 
                       (N1030)? mem[8057] : 
                       (N1032)? mem[8073] : 
                       (N1034)? mem[8089] : 
                       (N1036)? mem[8105] : 
                       (N1038)? mem[8121] : 
                       (N1040)? mem[8137] : 
                       (N1042)? mem[8153] : 
                       (N1044)? mem[8169] : 
                       (N1046)? mem[8185] : 1'b0;
  assign r_data_o[8] = (N535)? mem[8] : 
                       (N537)? mem[24] : 
                       (N539)? mem[40] : 
                       (N541)? mem[56] : 
                       (N543)? mem[72] : 
                       (N545)? mem[88] : 
                       (N547)? mem[104] : 
                       (N549)? mem[120] : 
                       (N551)? mem[136] : 
                       (N553)? mem[152] : 
                       (N555)? mem[168] : 
                       (N557)? mem[184] : 
                       (N559)? mem[200] : 
                       (N561)? mem[216] : 
                       (N563)? mem[232] : 
                       (N565)? mem[248] : 
                       (N567)? mem[264] : 
                       (N569)? mem[280] : 
                       (N571)? mem[296] : 
                       (N573)? mem[312] : 
                       (N575)? mem[328] : 
                       (N577)? mem[344] : 
                       (N579)? mem[360] : 
                       (N581)? mem[376] : 
                       (N583)? mem[392] : 
                       (N585)? mem[408] : 
                       (N587)? mem[424] : 
                       (N589)? mem[440] : 
                       (N591)? mem[456] : 
                       (N593)? mem[472] : 
                       (N595)? mem[488] : 
                       (N597)? mem[504] : 
                       (N599)? mem[520] : 
                       (N601)? mem[536] : 
                       (N603)? mem[552] : 
                       (N605)? mem[568] : 
                       (N607)? mem[584] : 
                       (N609)? mem[600] : 
                       (N611)? mem[616] : 
                       (N613)? mem[632] : 
                       (N615)? mem[648] : 
                       (N617)? mem[664] : 
                       (N619)? mem[680] : 
                       (N621)? mem[696] : 
                       (N623)? mem[712] : 
                       (N625)? mem[728] : 
                       (N627)? mem[744] : 
                       (N629)? mem[760] : 
                       (N631)? mem[776] : 
                       (N633)? mem[792] : 
                       (N635)? mem[808] : 
                       (N637)? mem[824] : 
                       (N639)? mem[840] : 
                       (N641)? mem[856] : 
                       (N643)? mem[872] : 
                       (N645)? mem[888] : 
                       (N647)? mem[904] : 
                       (N649)? mem[920] : 
                       (N651)? mem[936] : 
                       (N653)? mem[952] : 
                       (N655)? mem[968] : 
                       (N657)? mem[984] : 
                       (N659)? mem[1000] : 
                       (N661)? mem[1016] : 
                       (N663)? mem[1032] : 
                       (N665)? mem[1048] : 
                       (N667)? mem[1064] : 
                       (N669)? mem[1080] : 
                       (N671)? mem[1096] : 
                       (N673)? mem[1112] : 
                       (N675)? mem[1128] : 
                       (N677)? mem[1144] : 
                       (N679)? mem[1160] : 
                       (N681)? mem[1176] : 
                       (N683)? mem[1192] : 
                       (N685)? mem[1208] : 
                       (N687)? mem[1224] : 
                       (N689)? mem[1240] : 
                       (N691)? mem[1256] : 
                       (N693)? mem[1272] : 
                       (N695)? mem[1288] : 
                       (N697)? mem[1304] : 
                       (N699)? mem[1320] : 
                       (N701)? mem[1336] : 
                       (N703)? mem[1352] : 
                       (N705)? mem[1368] : 
                       (N707)? mem[1384] : 
                       (N709)? mem[1400] : 
                       (N711)? mem[1416] : 
                       (N713)? mem[1432] : 
                       (N715)? mem[1448] : 
                       (N717)? mem[1464] : 
                       (N719)? mem[1480] : 
                       (N721)? mem[1496] : 
                       (N723)? mem[1512] : 
                       (N725)? mem[1528] : 
                       (N727)? mem[1544] : 
                       (N729)? mem[1560] : 
                       (N731)? mem[1576] : 
                       (N733)? mem[1592] : 
                       (N735)? mem[1608] : 
                       (N737)? mem[1624] : 
                       (N739)? mem[1640] : 
                       (N741)? mem[1656] : 
                       (N743)? mem[1672] : 
                       (N745)? mem[1688] : 
                       (N747)? mem[1704] : 
                       (N749)? mem[1720] : 
                       (N751)? mem[1736] : 
                       (N753)? mem[1752] : 
                       (N755)? mem[1768] : 
                       (N757)? mem[1784] : 
                       (N759)? mem[1800] : 
                       (N761)? mem[1816] : 
                       (N763)? mem[1832] : 
                       (N765)? mem[1848] : 
                       (N767)? mem[1864] : 
                       (N769)? mem[1880] : 
                       (N771)? mem[1896] : 
                       (N773)? mem[1912] : 
                       (N775)? mem[1928] : 
                       (N777)? mem[1944] : 
                       (N779)? mem[1960] : 
                       (N781)? mem[1976] : 
                       (N783)? mem[1992] : 
                       (N785)? mem[2008] : 
                       (N787)? mem[2024] : 
                       (N789)? mem[2040] : 
                       (N791)? mem[2056] : 
                       (N793)? mem[2072] : 
                       (N795)? mem[2088] : 
                       (N797)? mem[2104] : 
                       (N799)? mem[2120] : 
                       (N801)? mem[2136] : 
                       (N803)? mem[2152] : 
                       (N805)? mem[2168] : 
                       (N807)? mem[2184] : 
                       (N809)? mem[2200] : 
                       (N811)? mem[2216] : 
                       (N813)? mem[2232] : 
                       (N815)? mem[2248] : 
                       (N817)? mem[2264] : 
                       (N819)? mem[2280] : 
                       (N821)? mem[2296] : 
                       (N823)? mem[2312] : 
                       (N825)? mem[2328] : 
                       (N827)? mem[2344] : 
                       (N829)? mem[2360] : 
                       (N831)? mem[2376] : 
                       (N833)? mem[2392] : 
                       (N835)? mem[2408] : 
                       (N837)? mem[2424] : 
                       (N839)? mem[2440] : 
                       (N841)? mem[2456] : 
                       (N843)? mem[2472] : 
                       (N845)? mem[2488] : 
                       (N847)? mem[2504] : 
                       (N849)? mem[2520] : 
                       (N851)? mem[2536] : 
                       (N853)? mem[2552] : 
                       (N855)? mem[2568] : 
                       (N857)? mem[2584] : 
                       (N859)? mem[2600] : 
                       (N861)? mem[2616] : 
                       (N863)? mem[2632] : 
                       (N865)? mem[2648] : 
                       (N867)? mem[2664] : 
                       (N869)? mem[2680] : 
                       (N871)? mem[2696] : 
                       (N873)? mem[2712] : 
                       (N875)? mem[2728] : 
                       (N877)? mem[2744] : 
                       (N879)? mem[2760] : 
                       (N881)? mem[2776] : 
                       (N883)? mem[2792] : 
                       (N885)? mem[2808] : 
                       (N887)? mem[2824] : 
                       (N889)? mem[2840] : 
                       (N891)? mem[2856] : 
                       (N893)? mem[2872] : 
                       (N895)? mem[2888] : 
                       (N897)? mem[2904] : 
                       (N899)? mem[2920] : 
                       (N901)? mem[2936] : 
                       (N903)? mem[2952] : 
                       (N905)? mem[2968] : 
                       (N907)? mem[2984] : 
                       (N909)? mem[3000] : 
                       (N911)? mem[3016] : 
                       (N913)? mem[3032] : 
                       (N915)? mem[3048] : 
                       (N917)? mem[3064] : 
                       (N919)? mem[3080] : 
                       (N921)? mem[3096] : 
                       (N923)? mem[3112] : 
                       (N925)? mem[3128] : 
                       (N927)? mem[3144] : 
                       (N929)? mem[3160] : 
                       (N931)? mem[3176] : 
                       (N933)? mem[3192] : 
                       (N935)? mem[3208] : 
                       (N937)? mem[3224] : 
                       (N939)? mem[3240] : 
                       (N941)? mem[3256] : 
                       (N943)? mem[3272] : 
                       (N945)? mem[3288] : 
                       (N947)? mem[3304] : 
                       (N949)? mem[3320] : 
                       (N951)? mem[3336] : 
                       (N953)? mem[3352] : 
                       (N955)? mem[3368] : 
                       (N957)? mem[3384] : 
                       (N959)? mem[3400] : 
                       (N961)? mem[3416] : 
                       (N963)? mem[3432] : 
                       (N965)? mem[3448] : 
                       (N967)? mem[3464] : 
                       (N969)? mem[3480] : 
                       (N971)? mem[3496] : 
                       (N973)? mem[3512] : 
                       (N975)? mem[3528] : 
                       (N977)? mem[3544] : 
                       (N979)? mem[3560] : 
                       (N981)? mem[3576] : 
                       (N983)? mem[3592] : 
                       (N985)? mem[3608] : 
                       (N987)? mem[3624] : 
                       (N989)? mem[3640] : 
                       (N991)? mem[3656] : 
                       (N993)? mem[3672] : 
                       (N995)? mem[3688] : 
                       (N997)? mem[3704] : 
                       (N999)? mem[3720] : 
                       (N1001)? mem[3736] : 
                       (N1003)? mem[3752] : 
                       (N1005)? mem[3768] : 
                       (N1007)? mem[3784] : 
                       (N1009)? mem[3800] : 
                       (N1011)? mem[3816] : 
                       (N1013)? mem[3832] : 
                       (N1015)? mem[3848] : 
                       (N1017)? mem[3864] : 
                       (N1019)? mem[3880] : 
                       (N1021)? mem[3896] : 
                       (N1023)? mem[3912] : 
                       (N1025)? mem[3928] : 
                       (N1027)? mem[3944] : 
                       (N1029)? mem[3960] : 
                       (N1031)? mem[3976] : 
                       (N1033)? mem[3992] : 
                       (N1035)? mem[4008] : 
                       (N1037)? mem[4024] : 
                       (N1039)? mem[4040] : 
                       (N1041)? mem[4056] : 
                       (N1043)? mem[4072] : 
                       (N1045)? mem[4088] : 
                       (N536)? mem[4104] : 
                       (N538)? mem[4120] : 
                       (N540)? mem[4136] : 
                       (N542)? mem[4152] : 
                       (N544)? mem[4168] : 
                       (N546)? mem[4184] : 
                       (N548)? mem[4200] : 
                       (N550)? mem[4216] : 
                       (N552)? mem[4232] : 
                       (N554)? mem[4248] : 
                       (N556)? mem[4264] : 
                       (N558)? mem[4280] : 
                       (N560)? mem[4296] : 
                       (N562)? mem[4312] : 
                       (N564)? mem[4328] : 
                       (N566)? mem[4344] : 
                       (N568)? mem[4360] : 
                       (N570)? mem[4376] : 
                       (N572)? mem[4392] : 
                       (N574)? mem[4408] : 
                       (N576)? mem[4424] : 
                       (N578)? mem[4440] : 
                       (N580)? mem[4456] : 
                       (N582)? mem[4472] : 
                       (N584)? mem[4488] : 
                       (N586)? mem[4504] : 
                       (N588)? mem[4520] : 
                       (N590)? mem[4536] : 
                       (N592)? mem[4552] : 
                       (N594)? mem[4568] : 
                       (N596)? mem[4584] : 
                       (N598)? mem[4600] : 
                       (N600)? mem[4616] : 
                       (N602)? mem[4632] : 
                       (N604)? mem[4648] : 
                       (N606)? mem[4664] : 
                       (N608)? mem[4680] : 
                       (N610)? mem[4696] : 
                       (N612)? mem[4712] : 
                       (N614)? mem[4728] : 
                       (N616)? mem[4744] : 
                       (N618)? mem[4760] : 
                       (N620)? mem[4776] : 
                       (N622)? mem[4792] : 
                       (N624)? mem[4808] : 
                       (N626)? mem[4824] : 
                       (N628)? mem[4840] : 
                       (N630)? mem[4856] : 
                       (N632)? mem[4872] : 
                       (N634)? mem[4888] : 
                       (N636)? mem[4904] : 
                       (N638)? mem[4920] : 
                       (N640)? mem[4936] : 
                       (N642)? mem[4952] : 
                       (N644)? mem[4968] : 
                       (N646)? mem[4984] : 
                       (N648)? mem[5000] : 
                       (N650)? mem[5016] : 
                       (N652)? mem[5032] : 
                       (N654)? mem[5048] : 
                       (N656)? mem[5064] : 
                       (N658)? mem[5080] : 
                       (N660)? mem[5096] : 
                       (N662)? mem[5112] : 
                       (N664)? mem[5128] : 
                       (N666)? mem[5144] : 
                       (N668)? mem[5160] : 
                       (N670)? mem[5176] : 
                       (N672)? mem[5192] : 
                       (N674)? mem[5208] : 
                       (N676)? mem[5224] : 
                       (N678)? mem[5240] : 
                       (N680)? mem[5256] : 
                       (N682)? mem[5272] : 
                       (N684)? mem[5288] : 
                       (N686)? mem[5304] : 
                       (N688)? mem[5320] : 
                       (N690)? mem[5336] : 
                       (N692)? mem[5352] : 
                       (N694)? mem[5368] : 
                       (N696)? mem[5384] : 
                       (N698)? mem[5400] : 
                       (N700)? mem[5416] : 
                       (N702)? mem[5432] : 
                       (N704)? mem[5448] : 
                       (N706)? mem[5464] : 
                       (N708)? mem[5480] : 
                       (N710)? mem[5496] : 
                       (N712)? mem[5512] : 
                       (N714)? mem[5528] : 
                       (N716)? mem[5544] : 
                       (N718)? mem[5560] : 
                       (N720)? mem[5576] : 
                       (N722)? mem[5592] : 
                       (N724)? mem[5608] : 
                       (N726)? mem[5624] : 
                       (N728)? mem[5640] : 
                       (N730)? mem[5656] : 
                       (N732)? mem[5672] : 
                       (N734)? mem[5688] : 
                       (N736)? mem[5704] : 
                       (N738)? mem[5720] : 
                       (N740)? mem[5736] : 
                       (N742)? mem[5752] : 
                       (N744)? mem[5768] : 
                       (N746)? mem[5784] : 
                       (N748)? mem[5800] : 
                       (N750)? mem[5816] : 
                       (N752)? mem[5832] : 
                       (N754)? mem[5848] : 
                       (N756)? mem[5864] : 
                       (N758)? mem[5880] : 
                       (N760)? mem[5896] : 
                       (N762)? mem[5912] : 
                       (N764)? mem[5928] : 
                       (N766)? mem[5944] : 
                       (N768)? mem[5960] : 
                       (N770)? mem[5976] : 
                       (N772)? mem[5992] : 
                       (N774)? mem[6008] : 
                       (N776)? mem[6024] : 
                       (N778)? mem[6040] : 
                       (N780)? mem[6056] : 
                       (N782)? mem[6072] : 
                       (N784)? mem[6088] : 
                       (N786)? mem[6104] : 
                       (N788)? mem[6120] : 
                       (N790)? mem[6136] : 
                       (N792)? mem[6152] : 
                       (N794)? mem[6168] : 
                       (N796)? mem[6184] : 
                       (N798)? mem[6200] : 
                       (N800)? mem[6216] : 
                       (N802)? mem[6232] : 
                       (N804)? mem[6248] : 
                       (N806)? mem[6264] : 
                       (N808)? mem[6280] : 
                       (N810)? mem[6296] : 
                       (N812)? mem[6312] : 
                       (N814)? mem[6328] : 
                       (N816)? mem[6344] : 
                       (N818)? mem[6360] : 
                       (N820)? mem[6376] : 
                       (N822)? mem[6392] : 
                       (N824)? mem[6408] : 
                       (N826)? mem[6424] : 
                       (N828)? mem[6440] : 
                       (N830)? mem[6456] : 
                       (N832)? mem[6472] : 
                       (N834)? mem[6488] : 
                       (N836)? mem[6504] : 
                       (N838)? mem[6520] : 
                       (N840)? mem[6536] : 
                       (N842)? mem[6552] : 
                       (N844)? mem[6568] : 
                       (N846)? mem[6584] : 
                       (N848)? mem[6600] : 
                       (N850)? mem[6616] : 
                       (N852)? mem[6632] : 
                       (N854)? mem[6648] : 
                       (N856)? mem[6664] : 
                       (N858)? mem[6680] : 
                       (N860)? mem[6696] : 
                       (N862)? mem[6712] : 
                       (N864)? mem[6728] : 
                       (N866)? mem[6744] : 
                       (N868)? mem[6760] : 
                       (N870)? mem[6776] : 
                       (N872)? mem[6792] : 
                       (N874)? mem[6808] : 
                       (N876)? mem[6824] : 
                       (N878)? mem[6840] : 
                       (N880)? mem[6856] : 
                       (N882)? mem[6872] : 
                       (N884)? mem[6888] : 
                       (N886)? mem[6904] : 
                       (N888)? mem[6920] : 
                       (N890)? mem[6936] : 
                       (N892)? mem[6952] : 
                       (N894)? mem[6968] : 
                       (N896)? mem[6984] : 
                       (N898)? mem[7000] : 
                       (N900)? mem[7016] : 
                       (N902)? mem[7032] : 
                       (N904)? mem[7048] : 
                       (N906)? mem[7064] : 
                       (N908)? mem[7080] : 
                       (N910)? mem[7096] : 
                       (N912)? mem[7112] : 
                       (N914)? mem[7128] : 
                       (N916)? mem[7144] : 
                       (N918)? mem[7160] : 
                       (N920)? mem[7176] : 
                       (N922)? mem[7192] : 
                       (N924)? mem[7208] : 
                       (N926)? mem[7224] : 
                       (N928)? mem[7240] : 
                       (N930)? mem[7256] : 
                       (N932)? mem[7272] : 
                       (N934)? mem[7288] : 
                       (N936)? mem[7304] : 
                       (N938)? mem[7320] : 
                       (N940)? mem[7336] : 
                       (N942)? mem[7352] : 
                       (N944)? mem[7368] : 
                       (N946)? mem[7384] : 
                       (N948)? mem[7400] : 
                       (N950)? mem[7416] : 
                       (N952)? mem[7432] : 
                       (N954)? mem[7448] : 
                       (N956)? mem[7464] : 
                       (N958)? mem[7480] : 
                       (N960)? mem[7496] : 
                       (N962)? mem[7512] : 
                       (N964)? mem[7528] : 
                       (N966)? mem[7544] : 
                       (N968)? mem[7560] : 
                       (N970)? mem[7576] : 
                       (N972)? mem[7592] : 
                       (N974)? mem[7608] : 
                       (N976)? mem[7624] : 
                       (N978)? mem[7640] : 
                       (N980)? mem[7656] : 
                       (N982)? mem[7672] : 
                       (N984)? mem[7688] : 
                       (N986)? mem[7704] : 
                       (N988)? mem[7720] : 
                       (N990)? mem[7736] : 
                       (N992)? mem[7752] : 
                       (N994)? mem[7768] : 
                       (N996)? mem[7784] : 
                       (N998)? mem[7800] : 
                       (N1000)? mem[7816] : 
                       (N1002)? mem[7832] : 
                       (N1004)? mem[7848] : 
                       (N1006)? mem[7864] : 
                       (N1008)? mem[7880] : 
                       (N1010)? mem[7896] : 
                       (N1012)? mem[7912] : 
                       (N1014)? mem[7928] : 
                       (N1016)? mem[7944] : 
                       (N1018)? mem[7960] : 
                       (N1020)? mem[7976] : 
                       (N1022)? mem[7992] : 
                       (N1024)? mem[8008] : 
                       (N1026)? mem[8024] : 
                       (N1028)? mem[8040] : 
                       (N1030)? mem[8056] : 
                       (N1032)? mem[8072] : 
                       (N1034)? mem[8088] : 
                       (N1036)? mem[8104] : 
                       (N1038)? mem[8120] : 
                       (N1040)? mem[8136] : 
                       (N1042)? mem[8152] : 
                       (N1044)? mem[8168] : 
                       (N1046)? mem[8184] : 1'b0;
  assign r_data_o[7] = (N535)? mem[7] : 
                       (N537)? mem[23] : 
                       (N539)? mem[39] : 
                       (N541)? mem[55] : 
                       (N543)? mem[71] : 
                       (N545)? mem[87] : 
                       (N547)? mem[103] : 
                       (N549)? mem[119] : 
                       (N551)? mem[135] : 
                       (N553)? mem[151] : 
                       (N555)? mem[167] : 
                       (N557)? mem[183] : 
                       (N559)? mem[199] : 
                       (N561)? mem[215] : 
                       (N563)? mem[231] : 
                       (N565)? mem[247] : 
                       (N567)? mem[263] : 
                       (N569)? mem[279] : 
                       (N571)? mem[295] : 
                       (N573)? mem[311] : 
                       (N575)? mem[327] : 
                       (N577)? mem[343] : 
                       (N579)? mem[359] : 
                       (N581)? mem[375] : 
                       (N583)? mem[391] : 
                       (N585)? mem[407] : 
                       (N587)? mem[423] : 
                       (N589)? mem[439] : 
                       (N591)? mem[455] : 
                       (N593)? mem[471] : 
                       (N595)? mem[487] : 
                       (N597)? mem[503] : 
                       (N599)? mem[519] : 
                       (N601)? mem[535] : 
                       (N603)? mem[551] : 
                       (N605)? mem[567] : 
                       (N607)? mem[583] : 
                       (N609)? mem[599] : 
                       (N611)? mem[615] : 
                       (N613)? mem[631] : 
                       (N615)? mem[647] : 
                       (N617)? mem[663] : 
                       (N619)? mem[679] : 
                       (N621)? mem[695] : 
                       (N623)? mem[711] : 
                       (N625)? mem[727] : 
                       (N627)? mem[743] : 
                       (N629)? mem[759] : 
                       (N631)? mem[775] : 
                       (N633)? mem[791] : 
                       (N635)? mem[807] : 
                       (N637)? mem[823] : 
                       (N639)? mem[839] : 
                       (N641)? mem[855] : 
                       (N643)? mem[871] : 
                       (N645)? mem[887] : 
                       (N647)? mem[903] : 
                       (N649)? mem[919] : 
                       (N651)? mem[935] : 
                       (N653)? mem[951] : 
                       (N655)? mem[967] : 
                       (N657)? mem[983] : 
                       (N659)? mem[999] : 
                       (N661)? mem[1015] : 
                       (N663)? mem[1031] : 
                       (N665)? mem[1047] : 
                       (N667)? mem[1063] : 
                       (N669)? mem[1079] : 
                       (N671)? mem[1095] : 
                       (N673)? mem[1111] : 
                       (N675)? mem[1127] : 
                       (N677)? mem[1143] : 
                       (N679)? mem[1159] : 
                       (N681)? mem[1175] : 
                       (N683)? mem[1191] : 
                       (N685)? mem[1207] : 
                       (N687)? mem[1223] : 
                       (N689)? mem[1239] : 
                       (N691)? mem[1255] : 
                       (N693)? mem[1271] : 
                       (N695)? mem[1287] : 
                       (N697)? mem[1303] : 
                       (N699)? mem[1319] : 
                       (N701)? mem[1335] : 
                       (N703)? mem[1351] : 
                       (N705)? mem[1367] : 
                       (N707)? mem[1383] : 
                       (N709)? mem[1399] : 
                       (N711)? mem[1415] : 
                       (N713)? mem[1431] : 
                       (N715)? mem[1447] : 
                       (N717)? mem[1463] : 
                       (N719)? mem[1479] : 
                       (N721)? mem[1495] : 
                       (N723)? mem[1511] : 
                       (N725)? mem[1527] : 
                       (N727)? mem[1543] : 
                       (N729)? mem[1559] : 
                       (N731)? mem[1575] : 
                       (N733)? mem[1591] : 
                       (N735)? mem[1607] : 
                       (N737)? mem[1623] : 
                       (N739)? mem[1639] : 
                       (N741)? mem[1655] : 
                       (N743)? mem[1671] : 
                       (N745)? mem[1687] : 
                       (N747)? mem[1703] : 
                       (N749)? mem[1719] : 
                       (N751)? mem[1735] : 
                       (N753)? mem[1751] : 
                       (N755)? mem[1767] : 
                       (N757)? mem[1783] : 
                       (N759)? mem[1799] : 
                       (N761)? mem[1815] : 
                       (N763)? mem[1831] : 
                       (N765)? mem[1847] : 
                       (N767)? mem[1863] : 
                       (N769)? mem[1879] : 
                       (N771)? mem[1895] : 
                       (N773)? mem[1911] : 
                       (N775)? mem[1927] : 
                       (N777)? mem[1943] : 
                       (N779)? mem[1959] : 
                       (N781)? mem[1975] : 
                       (N783)? mem[1991] : 
                       (N785)? mem[2007] : 
                       (N787)? mem[2023] : 
                       (N789)? mem[2039] : 
                       (N791)? mem[2055] : 
                       (N793)? mem[2071] : 
                       (N795)? mem[2087] : 
                       (N797)? mem[2103] : 
                       (N799)? mem[2119] : 
                       (N801)? mem[2135] : 
                       (N803)? mem[2151] : 
                       (N805)? mem[2167] : 
                       (N807)? mem[2183] : 
                       (N809)? mem[2199] : 
                       (N811)? mem[2215] : 
                       (N813)? mem[2231] : 
                       (N815)? mem[2247] : 
                       (N817)? mem[2263] : 
                       (N819)? mem[2279] : 
                       (N821)? mem[2295] : 
                       (N823)? mem[2311] : 
                       (N825)? mem[2327] : 
                       (N827)? mem[2343] : 
                       (N829)? mem[2359] : 
                       (N831)? mem[2375] : 
                       (N833)? mem[2391] : 
                       (N835)? mem[2407] : 
                       (N837)? mem[2423] : 
                       (N839)? mem[2439] : 
                       (N841)? mem[2455] : 
                       (N843)? mem[2471] : 
                       (N845)? mem[2487] : 
                       (N847)? mem[2503] : 
                       (N849)? mem[2519] : 
                       (N851)? mem[2535] : 
                       (N853)? mem[2551] : 
                       (N855)? mem[2567] : 
                       (N857)? mem[2583] : 
                       (N859)? mem[2599] : 
                       (N861)? mem[2615] : 
                       (N863)? mem[2631] : 
                       (N865)? mem[2647] : 
                       (N867)? mem[2663] : 
                       (N869)? mem[2679] : 
                       (N871)? mem[2695] : 
                       (N873)? mem[2711] : 
                       (N875)? mem[2727] : 
                       (N877)? mem[2743] : 
                       (N879)? mem[2759] : 
                       (N881)? mem[2775] : 
                       (N883)? mem[2791] : 
                       (N885)? mem[2807] : 
                       (N887)? mem[2823] : 
                       (N889)? mem[2839] : 
                       (N891)? mem[2855] : 
                       (N893)? mem[2871] : 
                       (N895)? mem[2887] : 
                       (N897)? mem[2903] : 
                       (N899)? mem[2919] : 
                       (N901)? mem[2935] : 
                       (N903)? mem[2951] : 
                       (N905)? mem[2967] : 
                       (N907)? mem[2983] : 
                       (N909)? mem[2999] : 
                       (N911)? mem[3015] : 
                       (N913)? mem[3031] : 
                       (N915)? mem[3047] : 
                       (N917)? mem[3063] : 
                       (N919)? mem[3079] : 
                       (N921)? mem[3095] : 
                       (N923)? mem[3111] : 
                       (N925)? mem[3127] : 
                       (N927)? mem[3143] : 
                       (N929)? mem[3159] : 
                       (N931)? mem[3175] : 
                       (N933)? mem[3191] : 
                       (N935)? mem[3207] : 
                       (N937)? mem[3223] : 
                       (N939)? mem[3239] : 
                       (N941)? mem[3255] : 
                       (N943)? mem[3271] : 
                       (N945)? mem[3287] : 
                       (N947)? mem[3303] : 
                       (N949)? mem[3319] : 
                       (N951)? mem[3335] : 
                       (N953)? mem[3351] : 
                       (N955)? mem[3367] : 
                       (N957)? mem[3383] : 
                       (N959)? mem[3399] : 
                       (N961)? mem[3415] : 
                       (N963)? mem[3431] : 
                       (N965)? mem[3447] : 
                       (N967)? mem[3463] : 
                       (N969)? mem[3479] : 
                       (N971)? mem[3495] : 
                       (N973)? mem[3511] : 
                       (N975)? mem[3527] : 
                       (N977)? mem[3543] : 
                       (N979)? mem[3559] : 
                       (N981)? mem[3575] : 
                       (N983)? mem[3591] : 
                       (N985)? mem[3607] : 
                       (N987)? mem[3623] : 
                       (N989)? mem[3639] : 
                       (N991)? mem[3655] : 
                       (N993)? mem[3671] : 
                       (N995)? mem[3687] : 
                       (N997)? mem[3703] : 
                       (N999)? mem[3719] : 
                       (N1001)? mem[3735] : 
                       (N1003)? mem[3751] : 
                       (N1005)? mem[3767] : 
                       (N1007)? mem[3783] : 
                       (N1009)? mem[3799] : 
                       (N1011)? mem[3815] : 
                       (N1013)? mem[3831] : 
                       (N1015)? mem[3847] : 
                       (N1017)? mem[3863] : 
                       (N1019)? mem[3879] : 
                       (N1021)? mem[3895] : 
                       (N1023)? mem[3911] : 
                       (N1025)? mem[3927] : 
                       (N1027)? mem[3943] : 
                       (N1029)? mem[3959] : 
                       (N1031)? mem[3975] : 
                       (N1033)? mem[3991] : 
                       (N1035)? mem[4007] : 
                       (N1037)? mem[4023] : 
                       (N1039)? mem[4039] : 
                       (N1041)? mem[4055] : 
                       (N1043)? mem[4071] : 
                       (N1045)? mem[4087] : 
                       (N536)? mem[4103] : 
                       (N538)? mem[4119] : 
                       (N540)? mem[4135] : 
                       (N542)? mem[4151] : 
                       (N544)? mem[4167] : 
                       (N546)? mem[4183] : 
                       (N548)? mem[4199] : 
                       (N550)? mem[4215] : 
                       (N552)? mem[4231] : 
                       (N554)? mem[4247] : 
                       (N556)? mem[4263] : 
                       (N558)? mem[4279] : 
                       (N560)? mem[4295] : 
                       (N562)? mem[4311] : 
                       (N564)? mem[4327] : 
                       (N566)? mem[4343] : 
                       (N568)? mem[4359] : 
                       (N570)? mem[4375] : 
                       (N572)? mem[4391] : 
                       (N574)? mem[4407] : 
                       (N576)? mem[4423] : 
                       (N578)? mem[4439] : 
                       (N580)? mem[4455] : 
                       (N582)? mem[4471] : 
                       (N584)? mem[4487] : 
                       (N586)? mem[4503] : 
                       (N588)? mem[4519] : 
                       (N590)? mem[4535] : 
                       (N592)? mem[4551] : 
                       (N594)? mem[4567] : 
                       (N596)? mem[4583] : 
                       (N598)? mem[4599] : 
                       (N600)? mem[4615] : 
                       (N602)? mem[4631] : 
                       (N604)? mem[4647] : 
                       (N606)? mem[4663] : 
                       (N608)? mem[4679] : 
                       (N610)? mem[4695] : 
                       (N612)? mem[4711] : 
                       (N614)? mem[4727] : 
                       (N616)? mem[4743] : 
                       (N618)? mem[4759] : 
                       (N620)? mem[4775] : 
                       (N622)? mem[4791] : 
                       (N624)? mem[4807] : 
                       (N626)? mem[4823] : 
                       (N628)? mem[4839] : 
                       (N630)? mem[4855] : 
                       (N632)? mem[4871] : 
                       (N634)? mem[4887] : 
                       (N636)? mem[4903] : 
                       (N638)? mem[4919] : 
                       (N640)? mem[4935] : 
                       (N642)? mem[4951] : 
                       (N644)? mem[4967] : 
                       (N646)? mem[4983] : 
                       (N648)? mem[4999] : 
                       (N650)? mem[5015] : 
                       (N652)? mem[5031] : 
                       (N654)? mem[5047] : 
                       (N656)? mem[5063] : 
                       (N658)? mem[5079] : 
                       (N660)? mem[5095] : 
                       (N662)? mem[5111] : 
                       (N664)? mem[5127] : 
                       (N666)? mem[5143] : 
                       (N668)? mem[5159] : 
                       (N670)? mem[5175] : 
                       (N672)? mem[5191] : 
                       (N674)? mem[5207] : 
                       (N676)? mem[5223] : 
                       (N678)? mem[5239] : 
                       (N680)? mem[5255] : 
                       (N682)? mem[5271] : 
                       (N684)? mem[5287] : 
                       (N686)? mem[5303] : 
                       (N688)? mem[5319] : 
                       (N690)? mem[5335] : 
                       (N692)? mem[5351] : 
                       (N694)? mem[5367] : 
                       (N696)? mem[5383] : 
                       (N698)? mem[5399] : 
                       (N700)? mem[5415] : 
                       (N702)? mem[5431] : 
                       (N704)? mem[5447] : 
                       (N706)? mem[5463] : 
                       (N708)? mem[5479] : 
                       (N710)? mem[5495] : 
                       (N712)? mem[5511] : 
                       (N714)? mem[5527] : 
                       (N716)? mem[5543] : 
                       (N718)? mem[5559] : 
                       (N720)? mem[5575] : 
                       (N722)? mem[5591] : 
                       (N724)? mem[5607] : 
                       (N726)? mem[5623] : 
                       (N728)? mem[5639] : 
                       (N730)? mem[5655] : 
                       (N732)? mem[5671] : 
                       (N734)? mem[5687] : 
                       (N736)? mem[5703] : 
                       (N738)? mem[5719] : 
                       (N740)? mem[5735] : 
                       (N742)? mem[5751] : 
                       (N744)? mem[5767] : 
                       (N746)? mem[5783] : 
                       (N748)? mem[5799] : 
                       (N750)? mem[5815] : 
                       (N752)? mem[5831] : 
                       (N754)? mem[5847] : 
                       (N756)? mem[5863] : 
                       (N758)? mem[5879] : 
                       (N760)? mem[5895] : 
                       (N762)? mem[5911] : 
                       (N764)? mem[5927] : 
                       (N766)? mem[5943] : 
                       (N768)? mem[5959] : 
                       (N770)? mem[5975] : 
                       (N772)? mem[5991] : 
                       (N774)? mem[6007] : 
                       (N776)? mem[6023] : 
                       (N778)? mem[6039] : 
                       (N780)? mem[6055] : 
                       (N782)? mem[6071] : 
                       (N784)? mem[6087] : 
                       (N786)? mem[6103] : 
                       (N788)? mem[6119] : 
                       (N790)? mem[6135] : 
                       (N792)? mem[6151] : 
                       (N794)? mem[6167] : 
                       (N796)? mem[6183] : 
                       (N798)? mem[6199] : 
                       (N800)? mem[6215] : 
                       (N802)? mem[6231] : 
                       (N804)? mem[6247] : 
                       (N806)? mem[6263] : 
                       (N808)? mem[6279] : 
                       (N810)? mem[6295] : 
                       (N812)? mem[6311] : 
                       (N814)? mem[6327] : 
                       (N816)? mem[6343] : 
                       (N818)? mem[6359] : 
                       (N820)? mem[6375] : 
                       (N822)? mem[6391] : 
                       (N824)? mem[6407] : 
                       (N826)? mem[6423] : 
                       (N828)? mem[6439] : 
                       (N830)? mem[6455] : 
                       (N832)? mem[6471] : 
                       (N834)? mem[6487] : 
                       (N836)? mem[6503] : 
                       (N838)? mem[6519] : 
                       (N840)? mem[6535] : 
                       (N842)? mem[6551] : 
                       (N844)? mem[6567] : 
                       (N846)? mem[6583] : 
                       (N848)? mem[6599] : 
                       (N850)? mem[6615] : 
                       (N852)? mem[6631] : 
                       (N854)? mem[6647] : 
                       (N856)? mem[6663] : 
                       (N858)? mem[6679] : 
                       (N860)? mem[6695] : 
                       (N862)? mem[6711] : 
                       (N864)? mem[6727] : 
                       (N866)? mem[6743] : 
                       (N868)? mem[6759] : 
                       (N870)? mem[6775] : 
                       (N872)? mem[6791] : 
                       (N874)? mem[6807] : 
                       (N876)? mem[6823] : 
                       (N878)? mem[6839] : 
                       (N880)? mem[6855] : 
                       (N882)? mem[6871] : 
                       (N884)? mem[6887] : 
                       (N886)? mem[6903] : 
                       (N888)? mem[6919] : 
                       (N890)? mem[6935] : 
                       (N892)? mem[6951] : 
                       (N894)? mem[6967] : 
                       (N896)? mem[6983] : 
                       (N898)? mem[6999] : 
                       (N900)? mem[7015] : 
                       (N902)? mem[7031] : 
                       (N904)? mem[7047] : 
                       (N906)? mem[7063] : 
                       (N908)? mem[7079] : 
                       (N910)? mem[7095] : 
                       (N912)? mem[7111] : 
                       (N914)? mem[7127] : 
                       (N916)? mem[7143] : 
                       (N918)? mem[7159] : 
                       (N920)? mem[7175] : 
                       (N922)? mem[7191] : 
                       (N924)? mem[7207] : 
                       (N926)? mem[7223] : 
                       (N928)? mem[7239] : 
                       (N930)? mem[7255] : 
                       (N932)? mem[7271] : 
                       (N934)? mem[7287] : 
                       (N936)? mem[7303] : 
                       (N938)? mem[7319] : 
                       (N940)? mem[7335] : 
                       (N942)? mem[7351] : 
                       (N944)? mem[7367] : 
                       (N946)? mem[7383] : 
                       (N948)? mem[7399] : 
                       (N950)? mem[7415] : 
                       (N952)? mem[7431] : 
                       (N954)? mem[7447] : 
                       (N956)? mem[7463] : 
                       (N958)? mem[7479] : 
                       (N960)? mem[7495] : 
                       (N962)? mem[7511] : 
                       (N964)? mem[7527] : 
                       (N966)? mem[7543] : 
                       (N968)? mem[7559] : 
                       (N970)? mem[7575] : 
                       (N972)? mem[7591] : 
                       (N974)? mem[7607] : 
                       (N976)? mem[7623] : 
                       (N978)? mem[7639] : 
                       (N980)? mem[7655] : 
                       (N982)? mem[7671] : 
                       (N984)? mem[7687] : 
                       (N986)? mem[7703] : 
                       (N988)? mem[7719] : 
                       (N990)? mem[7735] : 
                       (N992)? mem[7751] : 
                       (N994)? mem[7767] : 
                       (N996)? mem[7783] : 
                       (N998)? mem[7799] : 
                       (N1000)? mem[7815] : 
                       (N1002)? mem[7831] : 
                       (N1004)? mem[7847] : 
                       (N1006)? mem[7863] : 
                       (N1008)? mem[7879] : 
                       (N1010)? mem[7895] : 
                       (N1012)? mem[7911] : 
                       (N1014)? mem[7927] : 
                       (N1016)? mem[7943] : 
                       (N1018)? mem[7959] : 
                       (N1020)? mem[7975] : 
                       (N1022)? mem[7991] : 
                       (N1024)? mem[8007] : 
                       (N1026)? mem[8023] : 
                       (N1028)? mem[8039] : 
                       (N1030)? mem[8055] : 
                       (N1032)? mem[8071] : 
                       (N1034)? mem[8087] : 
                       (N1036)? mem[8103] : 
                       (N1038)? mem[8119] : 
                       (N1040)? mem[8135] : 
                       (N1042)? mem[8151] : 
                       (N1044)? mem[8167] : 
                       (N1046)? mem[8183] : 1'b0;
  assign r_data_o[6] = (N535)? mem[6] : 
                       (N537)? mem[22] : 
                       (N539)? mem[38] : 
                       (N541)? mem[54] : 
                       (N543)? mem[70] : 
                       (N545)? mem[86] : 
                       (N547)? mem[102] : 
                       (N549)? mem[118] : 
                       (N551)? mem[134] : 
                       (N553)? mem[150] : 
                       (N555)? mem[166] : 
                       (N557)? mem[182] : 
                       (N559)? mem[198] : 
                       (N561)? mem[214] : 
                       (N563)? mem[230] : 
                       (N565)? mem[246] : 
                       (N567)? mem[262] : 
                       (N569)? mem[278] : 
                       (N571)? mem[294] : 
                       (N573)? mem[310] : 
                       (N575)? mem[326] : 
                       (N577)? mem[342] : 
                       (N579)? mem[358] : 
                       (N581)? mem[374] : 
                       (N583)? mem[390] : 
                       (N585)? mem[406] : 
                       (N587)? mem[422] : 
                       (N589)? mem[438] : 
                       (N591)? mem[454] : 
                       (N593)? mem[470] : 
                       (N595)? mem[486] : 
                       (N597)? mem[502] : 
                       (N599)? mem[518] : 
                       (N601)? mem[534] : 
                       (N603)? mem[550] : 
                       (N605)? mem[566] : 
                       (N607)? mem[582] : 
                       (N609)? mem[598] : 
                       (N611)? mem[614] : 
                       (N613)? mem[630] : 
                       (N615)? mem[646] : 
                       (N617)? mem[662] : 
                       (N619)? mem[678] : 
                       (N621)? mem[694] : 
                       (N623)? mem[710] : 
                       (N625)? mem[726] : 
                       (N627)? mem[742] : 
                       (N629)? mem[758] : 
                       (N631)? mem[774] : 
                       (N633)? mem[790] : 
                       (N635)? mem[806] : 
                       (N637)? mem[822] : 
                       (N639)? mem[838] : 
                       (N641)? mem[854] : 
                       (N643)? mem[870] : 
                       (N645)? mem[886] : 
                       (N647)? mem[902] : 
                       (N649)? mem[918] : 
                       (N651)? mem[934] : 
                       (N653)? mem[950] : 
                       (N655)? mem[966] : 
                       (N657)? mem[982] : 
                       (N659)? mem[998] : 
                       (N661)? mem[1014] : 
                       (N663)? mem[1030] : 
                       (N665)? mem[1046] : 
                       (N667)? mem[1062] : 
                       (N669)? mem[1078] : 
                       (N671)? mem[1094] : 
                       (N673)? mem[1110] : 
                       (N675)? mem[1126] : 
                       (N677)? mem[1142] : 
                       (N679)? mem[1158] : 
                       (N681)? mem[1174] : 
                       (N683)? mem[1190] : 
                       (N685)? mem[1206] : 
                       (N687)? mem[1222] : 
                       (N689)? mem[1238] : 
                       (N691)? mem[1254] : 
                       (N693)? mem[1270] : 
                       (N695)? mem[1286] : 
                       (N697)? mem[1302] : 
                       (N699)? mem[1318] : 
                       (N701)? mem[1334] : 
                       (N703)? mem[1350] : 
                       (N705)? mem[1366] : 
                       (N707)? mem[1382] : 
                       (N709)? mem[1398] : 
                       (N711)? mem[1414] : 
                       (N713)? mem[1430] : 
                       (N715)? mem[1446] : 
                       (N717)? mem[1462] : 
                       (N719)? mem[1478] : 
                       (N721)? mem[1494] : 
                       (N723)? mem[1510] : 
                       (N725)? mem[1526] : 
                       (N727)? mem[1542] : 
                       (N729)? mem[1558] : 
                       (N731)? mem[1574] : 
                       (N733)? mem[1590] : 
                       (N735)? mem[1606] : 
                       (N737)? mem[1622] : 
                       (N739)? mem[1638] : 
                       (N741)? mem[1654] : 
                       (N743)? mem[1670] : 
                       (N745)? mem[1686] : 
                       (N747)? mem[1702] : 
                       (N749)? mem[1718] : 
                       (N751)? mem[1734] : 
                       (N753)? mem[1750] : 
                       (N755)? mem[1766] : 
                       (N757)? mem[1782] : 
                       (N759)? mem[1798] : 
                       (N761)? mem[1814] : 
                       (N763)? mem[1830] : 
                       (N765)? mem[1846] : 
                       (N767)? mem[1862] : 
                       (N769)? mem[1878] : 
                       (N771)? mem[1894] : 
                       (N773)? mem[1910] : 
                       (N775)? mem[1926] : 
                       (N777)? mem[1942] : 
                       (N779)? mem[1958] : 
                       (N781)? mem[1974] : 
                       (N783)? mem[1990] : 
                       (N785)? mem[2006] : 
                       (N787)? mem[2022] : 
                       (N789)? mem[2038] : 
                       (N791)? mem[2054] : 
                       (N793)? mem[2070] : 
                       (N795)? mem[2086] : 
                       (N797)? mem[2102] : 
                       (N799)? mem[2118] : 
                       (N801)? mem[2134] : 
                       (N803)? mem[2150] : 
                       (N805)? mem[2166] : 
                       (N807)? mem[2182] : 
                       (N809)? mem[2198] : 
                       (N811)? mem[2214] : 
                       (N813)? mem[2230] : 
                       (N815)? mem[2246] : 
                       (N817)? mem[2262] : 
                       (N819)? mem[2278] : 
                       (N821)? mem[2294] : 
                       (N823)? mem[2310] : 
                       (N825)? mem[2326] : 
                       (N827)? mem[2342] : 
                       (N829)? mem[2358] : 
                       (N831)? mem[2374] : 
                       (N833)? mem[2390] : 
                       (N835)? mem[2406] : 
                       (N837)? mem[2422] : 
                       (N839)? mem[2438] : 
                       (N841)? mem[2454] : 
                       (N843)? mem[2470] : 
                       (N845)? mem[2486] : 
                       (N847)? mem[2502] : 
                       (N849)? mem[2518] : 
                       (N851)? mem[2534] : 
                       (N853)? mem[2550] : 
                       (N855)? mem[2566] : 
                       (N857)? mem[2582] : 
                       (N859)? mem[2598] : 
                       (N861)? mem[2614] : 
                       (N863)? mem[2630] : 
                       (N865)? mem[2646] : 
                       (N867)? mem[2662] : 
                       (N869)? mem[2678] : 
                       (N871)? mem[2694] : 
                       (N873)? mem[2710] : 
                       (N875)? mem[2726] : 
                       (N877)? mem[2742] : 
                       (N879)? mem[2758] : 
                       (N881)? mem[2774] : 
                       (N883)? mem[2790] : 
                       (N885)? mem[2806] : 
                       (N887)? mem[2822] : 
                       (N889)? mem[2838] : 
                       (N891)? mem[2854] : 
                       (N893)? mem[2870] : 
                       (N895)? mem[2886] : 
                       (N897)? mem[2902] : 
                       (N899)? mem[2918] : 
                       (N901)? mem[2934] : 
                       (N903)? mem[2950] : 
                       (N905)? mem[2966] : 
                       (N907)? mem[2982] : 
                       (N909)? mem[2998] : 
                       (N911)? mem[3014] : 
                       (N913)? mem[3030] : 
                       (N915)? mem[3046] : 
                       (N917)? mem[3062] : 
                       (N919)? mem[3078] : 
                       (N921)? mem[3094] : 
                       (N923)? mem[3110] : 
                       (N925)? mem[3126] : 
                       (N927)? mem[3142] : 
                       (N929)? mem[3158] : 
                       (N931)? mem[3174] : 
                       (N933)? mem[3190] : 
                       (N935)? mem[3206] : 
                       (N937)? mem[3222] : 
                       (N939)? mem[3238] : 
                       (N941)? mem[3254] : 
                       (N943)? mem[3270] : 
                       (N945)? mem[3286] : 
                       (N947)? mem[3302] : 
                       (N949)? mem[3318] : 
                       (N951)? mem[3334] : 
                       (N953)? mem[3350] : 
                       (N955)? mem[3366] : 
                       (N957)? mem[3382] : 
                       (N959)? mem[3398] : 
                       (N961)? mem[3414] : 
                       (N963)? mem[3430] : 
                       (N965)? mem[3446] : 
                       (N967)? mem[3462] : 
                       (N969)? mem[3478] : 
                       (N971)? mem[3494] : 
                       (N973)? mem[3510] : 
                       (N975)? mem[3526] : 
                       (N977)? mem[3542] : 
                       (N979)? mem[3558] : 
                       (N981)? mem[3574] : 
                       (N983)? mem[3590] : 
                       (N985)? mem[3606] : 
                       (N987)? mem[3622] : 
                       (N989)? mem[3638] : 
                       (N991)? mem[3654] : 
                       (N993)? mem[3670] : 
                       (N995)? mem[3686] : 
                       (N997)? mem[3702] : 
                       (N999)? mem[3718] : 
                       (N1001)? mem[3734] : 
                       (N1003)? mem[3750] : 
                       (N1005)? mem[3766] : 
                       (N1007)? mem[3782] : 
                       (N1009)? mem[3798] : 
                       (N1011)? mem[3814] : 
                       (N1013)? mem[3830] : 
                       (N1015)? mem[3846] : 
                       (N1017)? mem[3862] : 
                       (N1019)? mem[3878] : 
                       (N1021)? mem[3894] : 
                       (N1023)? mem[3910] : 
                       (N1025)? mem[3926] : 
                       (N1027)? mem[3942] : 
                       (N1029)? mem[3958] : 
                       (N1031)? mem[3974] : 
                       (N1033)? mem[3990] : 
                       (N1035)? mem[4006] : 
                       (N1037)? mem[4022] : 
                       (N1039)? mem[4038] : 
                       (N1041)? mem[4054] : 
                       (N1043)? mem[4070] : 
                       (N1045)? mem[4086] : 
                       (N536)? mem[4102] : 
                       (N538)? mem[4118] : 
                       (N540)? mem[4134] : 
                       (N542)? mem[4150] : 
                       (N544)? mem[4166] : 
                       (N546)? mem[4182] : 
                       (N548)? mem[4198] : 
                       (N550)? mem[4214] : 
                       (N552)? mem[4230] : 
                       (N554)? mem[4246] : 
                       (N556)? mem[4262] : 
                       (N558)? mem[4278] : 
                       (N560)? mem[4294] : 
                       (N562)? mem[4310] : 
                       (N564)? mem[4326] : 
                       (N566)? mem[4342] : 
                       (N568)? mem[4358] : 
                       (N570)? mem[4374] : 
                       (N572)? mem[4390] : 
                       (N574)? mem[4406] : 
                       (N576)? mem[4422] : 
                       (N578)? mem[4438] : 
                       (N580)? mem[4454] : 
                       (N582)? mem[4470] : 
                       (N584)? mem[4486] : 
                       (N586)? mem[4502] : 
                       (N588)? mem[4518] : 
                       (N590)? mem[4534] : 
                       (N592)? mem[4550] : 
                       (N594)? mem[4566] : 
                       (N596)? mem[4582] : 
                       (N598)? mem[4598] : 
                       (N600)? mem[4614] : 
                       (N602)? mem[4630] : 
                       (N604)? mem[4646] : 
                       (N606)? mem[4662] : 
                       (N608)? mem[4678] : 
                       (N610)? mem[4694] : 
                       (N612)? mem[4710] : 
                       (N614)? mem[4726] : 
                       (N616)? mem[4742] : 
                       (N618)? mem[4758] : 
                       (N620)? mem[4774] : 
                       (N622)? mem[4790] : 
                       (N624)? mem[4806] : 
                       (N626)? mem[4822] : 
                       (N628)? mem[4838] : 
                       (N630)? mem[4854] : 
                       (N632)? mem[4870] : 
                       (N634)? mem[4886] : 
                       (N636)? mem[4902] : 
                       (N638)? mem[4918] : 
                       (N640)? mem[4934] : 
                       (N642)? mem[4950] : 
                       (N644)? mem[4966] : 
                       (N646)? mem[4982] : 
                       (N648)? mem[4998] : 
                       (N650)? mem[5014] : 
                       (N652)? mem[5030] : 
                       (N654)? mem[5046] : 
                       (N656)? mem[5062] : 
                       (N658)? mem[5078] : 
                       (N660)? mem[5094] : 
                       (N662)? mem[5110] : 
                       (N664)? mem[5126] : 
                       (N666)? mem[5142] : 
                       (N668)? mem[5158] : 
                       (N670)? mem[5174] : 
                       (N672)? mem[5190] : 
                       (N674)? mem[5206] : 
                       (N676)? mem[5222] : 
                       (N678)? mem[5238] : 
                       (N680)? mem[5254] : 
                       (N682)? mem[5270] : 
                       (N684)? mem[5286] : 
                       (N686)? mem[5302] : 
                       (N688)? mem[5318] : 
                       (N690)? mem[5334] : 
                       (N692)? mem[5350] : 
                       (N694)? mem[5366] : 
                       (N696)? mem[5382] : 
                       (N698)? mem[5398] : 
                       (N700)? mem[5414] : 
                       (N702)? mem[5430] : 
                       (N704)? mem[5446] : 
                       (N706)? mem[5462] : 
                       (N708)? mem[5478] : 
                       (N710)? mem[5494] : 
                       (N712)? mem[5510] : 
                       (N714)? mem[5526] : 
                       (N716)? mem[5542] : 
                       (N718)? mem[5558] : 
                       (N720)? mem[5574] : 
                       (N722)? mem[5590] : 
                       (N724)? mem[5606] : 
                       (N726)? mem[5622] : 
                       (N728)? mem[5638] : 
                       (N730)? mem[5654] : 
                       (N732)? mem[5670] : 
                       (N734)? mem[5686] : 
                       (N736)? mem[5702] : 
                       (N738)? mem[5718] : 
                       (N740)? mem[5734] : 
                       (N742)? mem[5750] : 
                       (N744)? mem[5766] : 
                       (N746)? mem[5782] : 
                       (N748)? mem[5798] : 
                       (N750)? mem[5814] : 
                       (N752)? mem[5830] : 
                       (N754)? mem[5846] : 
                       (N756)? mem[5862] : 
                       (N758)? mem[5878] : 
                       (N760)? mem[5894] : 
                       (N762)? mem[5910] : 
                       (N764)? mem[5926] : 
                       (N766)? mem[5942] : 
                       (N768)? mem[5958] : 
                       (N770)? mem[5974] : 
                       (N772)? mem[5990] : 
                       (N774)? mem[6006] : 
                       (N776)? mem[6022] : 
                       (N778)? mem[6038] : 
                       (N780)? mem[6054] : 
                       (N782)? mem[6070] : 
                       (N784)? mem[6086] : 
                       (N786)? mem[6102] : 
                       (N788)? mem[6118] : 
                       (N790)? mem[6134] : 
                       (N792)? mem[6150] : 
                       (N794)? mem[6166] : 
                       (N796)? mem[6182] : 
                       (N798)? mem[6198] : 
                       (N800)? mem[6214] : 
                       (N802)? mem[6230] : 
                       (N804)? mem[6246] : 
                       (N806)? mem[6262] : 
                       (N808)? mem[6278] : 
                       (N810)? mem[6294] : 
                       (N812)? mem[6310] : 
                       (N814)? mem[6326] : 
                       (N816)? mem[6342] : 
                       (N818)? mem[6358] : 
                       (N820)? mem[6374] : 
                       (N822)? mem[6390] : 
                       (N824)? mem[6406] : 
                       (N826)? mem[6422] : 
                       (N828)? mem[6438] : 
                       (N830)? mem[6454] : 
                       (N832)? mem[6470] : 
                       (N834)? mem[6486] : 
                       (N836)? mem[6502] : 
                       (N838)? mem[6518] : 
                       (N840)? mem[6534] : 
                       (N842)? mem[6550] : 
                       (N844)? mem[6566] : 
                       (N846)? mem[6582] : 
                       (N848)? mem[6598] : 
                       (N850)? mem[6614] : 
                       (N852)? mem[6630] : 
                       (N854)? mem[6646] : 
                       (N856)? mem[6662] : 
                       (N858)? mem[6678] : 
                       (N860)? mem[6694] : 
                       (N862)? mem[6710] : 
                       (N864)? mem[6726] : 
                       (N866)? mem[6742] : 
                       (N868)? mem[6758] : 
                       (N870)? mem[6774] : 
                       (N872)? mem[6790] : 
                       (N874)? mem[6806] : 
                       (N876)? mem[6822] : 
                       (N878)? mem[6838] : 
                       (N880)? mem[6854] : 
                       (N882)? mem[6870] : 
                       (N884)? mem[6886] : 
                       (N886)? mem[6902] : 
                       (N888)? mem[6918] : 
                       (N890)? mem[6934] : 
                       (N892)? mem[6950] : 
                       (N894)? mem[6966] : 
                       (N896)? mem[6982] : 
                       (N898)? mem[6998] : 
                       (N900)? mem[7014] : 
                       (N902)? mem[7030] : 
                       (N904)? mem[7046] : 
                       (N906)? mem[7062] : 
                       (N908)? mem[7078] : 
                       (N910)? mem[7094] : 
                       (N912)? mem[7110] : 
                       (N914)? mem[7126] : 
                       (N916)? mem[7142] : 
                       (N918)? mem[7158] : 
                       (N920)? mem[7174] : 
                       (N922)? mem[7190] : 
                       (N924)? mem[7206] : 
                       (N926)? mem[7222] : 
                       (N928)? mem[7238] : 
                       (N930)? mem[7254] : 
                       (N932)? mem[7270] : 
                       (N934)? mem[7286] : 
                       (N936)? mem[7302] : 
                       (N938)? mem[7318] : 
                       (N940)? mem[7334] : 
                       (N942)? mem[7350] : 
                       (N944)? mem[7366] : 
                       (N946)? mem[7382] : 
                       (N948)? mem[7398] : 
                       (N950)? mem[7414] : 
                       (N952)? mem[7430] : 
                       (N954)? mem[7446] : 
                       (N956)? mem[7462] : 
                       (N958)? mem[7478] : 
                       (N960)? mem[7494] : 
                       (N962)? mem[7510] : 
                       (N964)? mem[7526] : 
                       (N966)? mem[7542] : 
                       (N968)? mem[7558] : 
                       (N970)? mem[7574] : 
                       (N972)? mem[7590] : 
                       (N974)? mem[7606] : 
                       (N976)? mem[7622] : 
                       (N978)? mem[7638] : 
                       (N980)? mem[7654] : 
                       (N982)? mem[7670] : 
                       (N984)? mem[7686] : 
                       (N986)? mem[7702] : 
                       (N988)? mem[7718] : 
                       (N990)? mem[7734] : 
                       (N992)? mem[7750] : 
                       (N994)? mem[7766] : 
                       (N996)? mem[7782] : 
                       (N998)? mem[7798] : 
                       (N1000)? mem[7814] : 
                       (N1002)? mem[7830] : 
                       (N1004)? mem[7846] : 
                       (N1006)? mem[7862] : 
                       (N1008)? mem[7878] : 
                       (N1010)? mem[7894] : 
                       (N1012)? mem[7910] : 
                       (N1014)? mem[7926] : 
                       (N1016)? mem[7942] : 
                       (N1018)? mem[7958] : 
                       (N1020)? mem[7974] : 
                       (N1022)? mem[7990] : 
                       (N1024)? mem[8006] : 
                       (N1026)? mem[8022] : 
                       (N1028)? mem[8038] : 
                       (N1030)? mem[8054] : 
                       (N1032)? mem[8070] : 
                       (N1034)? mem[8086] : 
                       (N1036)? mem[8102] : 
                       (N1038)? mem[8118] : 
                       (N1040)? mem[8134] : 
                       (N1042)? mem[8150] : 
                       (N1044)? mem[8166] : 
                       (N1046)? mem[8182] : 1'b0;
  assign r_data_o[5] = (N535)? mem[5] : 
                       (N537)? mem[21] : 
                       (N539)? mem[37] : 
                       (N541)? mem[53] : 
                       (N543)? mem[69] : 
                       (N545)? mem[85] : 
                       (N547)? mem[101] : 
                       (N549)? mem[117] : 
                       (N551)? mem[133] : 
                       (N553)? mem[149] : 
                       (N555)? mem[165] : 
                       (N557)? mem[181] : 
                       (N559)? mem[197] : 
                       (N561)? mem[213] : 
                       (N563)? mem[229] : 
                       (N565)? mem[245] : 
                       (N567)? mem[261] : 
                       (N569)? mem[277] : 
                       (N571)? mem[293] : 
                       (N573)? mem[309] : 
                       (N575)? mem[325] : 
                       (N577)? mem[341] : 
                       (N579)? mem[357] : 
                       (N581)? mem[373] : 
                       (N583)? mem[389] : 
                       (N585)? mem[405] : 
                       (N587)? mem[421] : 
                       (N589)? mem[437] : 
                       (N591)? mem[453] : 
                       (N593)? mem[469] : 
                       (N595)? mem[485] : 
                       (N597)? mem[501] : 
                       (N599)? mem[517] : 
                       (N601)? mem[533] : 
                       (N603)? mem[549] : 
                       (N605)? mem[565] : 
                       (N607)? mem[581] : 
                       (N609)? mem[597] : 
                       (N611)? mem[613] : 
                       (N613)? mem[629] : 
                       (N615)? mem[645] : 
                       (N617)? mem[661] : 
                       (N619)? mem[677] : 
                       (N621)? mem[693] : 
                       (N623)? mem[709] : 
                       (N625)? mem[725] : 
                       (N627)? mem[741] : 
                       (N629)? mem[757] : 
                       (N631)? mem[773] : 
                       (N633)? mem[789] : 
                       (N635)? mem[805] : 
                       (N637)? mem[821] : 
                       (N639)? mem[837] : 
                       (N641)? mem[853] : 
                       (N643)? mem[869] : 
                       (N645)? mem[885] : 
                       (N647)? mem[901] : 
                       (N649)? mem[917] : 
                       (N651)? mem[933] : 
                       (N653)? mem[949] : 
                       (N655)? mem[965] : 
                       (N657)? mem[981] : 
                       (N659)? mem[997] : 
                       (N661)? mem[1013] : 
                       (N663)? mem[1029] : 
                       (N665)? mem[1045] : 
                       (N667)? mem[1061] : 
                       (N669)? mem[1077] : 
                       (N671)? mem[1093] : 
                       (N673)? mem[1109] : 
                       (N675)? mem[1125] : 
                       (N677)? mem[1141] : 
                       (N679)? mem[1157] : 
                       (N681)? mem[1173] : 
                       (N683)? mem[1189] : 
                       (N685)? mem[1205] : 
                       (N687)? mem[1221] : 
                       (N689)? mem[1237] : 
                       (N691)? mem[1253] : 
                       (N693)? mem[1269] : 
                       (N695)? mem[1285] : 
                       (N697)? mem[1301] : 
                       (N699)? mem[1317] : 
                       (N701)? mem[1333] : 
                       (N703)? mem[1349] : 
                       (N705)? mem[1365] : 
                       (N707)? mem[1381] : 
                       (N709)? mem[1397] : 
                       (N711)? mem[1413] : 
                       (N713)? mem[1429] : 
                       (N715)? mem[1445] : 
                       (N717)? mem[1461] : 
                       (N719)? mem[1477] : 
                       (N721)? mem[1493] : 
                       (N723)? mem[1509] : 
                       (N725)? mem[1525] : 
                       (N727)? mem[1541] : 
                       (N729)? mem[1557] : 
                       (N731)? mem[1573] : 
                       (N733)? mem[1589] : 
                       (N735)? mem[1605] : 
                       (N737)? mem[1621] : 
                       (N739)? mem[1637] : 
                       (N741)? mem[1653] : 
                       (N743)? mem[1669] : 
                       (N745)? mem[1685] : 
                       (N747)? mem[1701] : 
                       (N749)? mem[1717] : 
                       (N751)? mem[1733] : 
                       (N753)? mem[1749] : 
                       (N755)? mem[1765] : 
                       (N757)? mem[1781] : 
                       (N759)? mem[1797] : 
                       (N761)? mem[1813] : 
                       (N763)? mem[1829] : 
                       (N765)? mem[1845] : 
                       (N767)? mem[1861] : 
                       (N769)? mem[1877] : 
                       (N771)? mem[1893] : 
                       (N773)? mem[1909] : 
                       (N775)? mem[1925] : 
                       (N777)? mem[1941] : 
                       (N779)? mem[1957] : 
                       (N781)? mem[1973] : 
                       (N783)? mem[1989] : 
                       (N785)? mem[2005] : 
                       (N787)? mem[2021] : 
                       (N789)? mem[2037] : 
                       (N791)? mem[2053] : 
                       (N793)? mem[2069] : 
                       (N795)? mem[2085] : 
                       (N797)? mem[2101] : 
                       (N799)? mem[2117] : 
                       (N801)? mem[2133] : 
                       (N803)? mem[2149] : 
                       (N805)? mem[2165] : 
                       (N807)? mem[2181] : 
                       (N809)? mem[2197] : 
                       (N811)? mem[2213] : 
                       (N813)? mem[2229] : 
                       (N815)? mem[2245] : 
                       (N817)? mem[2261] : 
                       (N819)? mem[2277] : 
                       (N821)? mem[2293] : 
                       (N823)? mem[2309] : 
                       (N825)? mem[2325] : 
                       (N827)? mem[2341] : 
                       (N829)? mem[2357] : 
                       (N831)? mem[2373] : 
                       (N833)? mem[2389] : 
                       (N835)? mem[2405] : 
                       (N837)? mem[2421] : 
                       (N839)? mem[2437] : 
                       (N841)? mem[2453] : 
                       (N843)? mem[2469] : 
                       (N845)? mem[2485] : 
                       (N847)? mem[2501] : 
                       (N849)? mem[2517] : 
                       (N851)? mem[2533] : 
                       (N853)? mem[2549] : 
                       (N855)? mem[2565] : 
                       (N857)? mem[2581] : 
                       (N859)? mem[2597] : 
                       (N861)? mem[2613] : 
                       (N863)? mem[2629] : 
                       (N865)? mem[2645] : 
                       (N867)? mem[2661] : 
                       (N869)? mem[2677] : 
                       (N871)? mem[2693] : 
                       (N873)? mem[2709] : 
                       (N875)? mem[2725] : 
                       (N877)? mem[2741] : 
                       (N879)? mem[2757] : 
                       (N881)? mem[2773] : 
                       (N883)? mem[2789] : 
                       (N885)? mem[2805] : 
                       (N887)? mem[2821] : 
                       (N889)? mem[2837] : 
                       (N891)? mem[2853] : 
                       (N893)? mem[2869] : 
                       (N895)? mem[2885] : 
                       (N897)? mem[2901] : 
                       (N899)? mem[2917] : 
                       (N901)? mem[2933] : 
                       (N903)? mem[2949] : 
                       (N905)? mem[2965] : 
                       (N907)? mem[2981] : 
                       (N909)? mem[2997] : 
                       (N911)? mem[3013] : 
                       (N913)? mem[3029] : 
                       (N915)? mem[3045] : 
                       (N917)? mem[3061] : 
                       (N919)? mem[3077] : 
                       (N921)? mem[3093] : 
                       (N923)? mem[3109] : 
                       (N925)? mem[3125] : 
                       (N927)? mem[3141] : 
                       (N929)? mem[3157] : 
                       (N931)? mem[3173] : 
                       (N933)? mem[3189] : 
                       (N935)? mem[3205] : 
                       (N937)? mem[3221] : 
                       (N939)? mem[3237] : 
                       (N941)? mem[3253] : 
                       (N943)? mem[3269] : 
                       (N945)? mem[3285] : 
                       (N947)? mem[3301] : 
                       (N949)? mem[3317] : 
                       (N951)? mem[3333] : 
                       (N953)? mem[3349] : 
                       (N955)? mem[3365] : 
                       (N957)? mem[3381] : 
                       (N959)? mem[3397] : 
                       (N961)? mem[3413] : 
                       (N963)? mem[3429] : 
                       (N965)? mem[3445] : 
                       (N967)? mem[3461] : 
                       (N969)? mem[3477] : 
                       (N971)? mem[3493] : 
                       (N973)? mem[3509] : 
                       (N975)? mem[3525] : 
                       (N977)? mem[3541] : 
                       (N979)? mem[3557] : 
                       (N981)? mem[3573] : 
                       (N983)? mem[3589] : 
                       (N985)? mem[3605] : 
                       (N987)? mem[3621] : 
                       (N989)? mem[3637] : 
                       (N991)? mem[3653] : 
                       (N993)? mem[3669] : 
                       (N995)? mem[3685] : 
                       (N997)? mem[3701] : 
                       (N999)? mem[3717] : 
                       (N1001)? mem[3733] : 
                       (N1003)? mem[3749] : 
                       (N1005)? mem[3765] : 
                       (N1007)? mem[3781] : 
                       (N1009)? mem[3797] : 
                       (N1011)? mem[3813] : 
                       (N1013)? mem[3829] : 
                       (N1015)? mem[3845] : 
                       (N1017)? mem[3861] : 
                       (N1019)? mem[3877] : 
                       (N1021)? mem[3893] : 
                       (N1023)? mem[3909] : 
                       (N1025)? mem[3925] : 
                       (N1027)? mem[3941] : 
                       (N1029)? mem[3957] : 
                       (N1031)? mem[3973] : 
                       (N1033)? mem[3989] : 
                       (N1035)? mem[4005] : 
                       (N1037)? mem[4021] : 
                       (N1039)? mem[4037] : 
                       (N1041)? mem[4053] : 
                       (N1043)? mem[4069] : 
                       (N1045)? mem[4085] : 
                       (N536)? mem[4101] : 
                       (N538)? mem[4117] : 
                       (N540)? mem[4133] : 
                       (N542)? mem[4149] : 
                       (N544)? mem[4165] : 
                       (N546)? mem[4181] : 
                       (N548)? mem[4197] : 
                       (N550)? mem[4213] : 
                       (N552)? mem[4229] : 
                       (N554)? mem[4245] : 
                       (N556)? mem[4261] : 
                       (N558)? mem[4277] : 
                       (N560)? mem[4293] : 
                       (N562)? mem[4309] : 
                       (N564)? mem[4325] : 
                       (N566)? mem[4341] : 
                       (N568)? mem[4357] : 
                       (N570)? mem[4373] : 
                       (N572)? mem[4389] : 
                       (N574)? mem[4405] : 
                       (N576)? mem[4421] : 
                       (N578)? mem[4437] : 
                       (N580)? mem[4453] : 
                       (N582)? mem[4469] : 
                       (N584)? mem[4485] : 
                       (N586)? mem[4501] : 
                       (N588)? mem[4517] : 
                       (N590)? mem[4533] : 
                       (N592)? mem[4549] : 
                       (N594)? mem[4565] : 
                       (N596)? mem[4581] : 
                       (N598)? mem[4597] : 
                       (N600)? mem[4613] : 
                       (N602)? mem[4629] : 
                       (N604)? mem[4645] : 
                       (N606)? mem[4661] : 
                       (N608)? mem[4677] : 
                       (N610)? mem[4693] : 
                       (N612)? mem[4709] : 
                       (N614)? mem[4725] : 
                       (N616)? mem[4741] : 
                       (N618)? mem[4757] : 
                       (N620)? mem[4773] : 
                       (N622)? mem[4789] : 
                       (N624)? mem[4805] : 
                       (N626)? mem[4821] : 
                       (N628)? mem[4837] : 
                       (N630)? mem[4853] : 
                       (N632)? mem[4869] : 
                       (N634)? mem[4885] : 
                       (N636)? mem[4901] : 
                       (N638)? mem[4917] : 
                       (N640)? mem[4933] : 
                       (N642)? mem[4949] : 
                       (N644)? mem[4965] : 
                       (N646)? mem[4981] : 
                       (N648)? mem[4997] : 
                       (N650)? mem[5013] : 
                       (N652)? mem[5029] : 
                       (N654)? mem[5045] : 
                       (N656)? mem[5061] : 
                       (N658)? mem[5077] : 
                       (N660)? mem[5093] : 
                       (N662)? mem[5109] : 
                       (N664)? mem[5125] : 
                       (N666)? mem[5141] : 
                       (N668)? mem[5157] : 
                       (N670)? mem[5173] : 
                       (N672)? mem[5189] : 
                       (N674)? mem[5205] : 
                       (N676)? mem[5221] : 
                       (N678)? mem[5237] : 
                       (N680)? mem[5253] : 
                       (N682)? mem[5269] : 
                       (N684)? mem[5285] : 
                       (N686)? mem[5301] : 
                       (N688)? mem[5317] : 
                       (N690)? mem[5333] : 
                       (N692)? mem[5349] : 
                       (N694)? mem[5365] : 
                       (N696)? mem[5381] : 
                       (N698)? mem[5397] : 
                       (N700)? mem[5413] : 
                       (N702)? mem[5429] : 
                       (N704)? mem[5445] : 
                       (N706)? mem[5461] : 
                       (N708)? mem[5477] : 
                       (N710)? mem[5493] : 
                       (N712)? mem[5509] : 
                       (N714)? mem[5525] : 
                       (N716)? mem[5541] : 
                       (N718)? mem[5557] : 
                       (N720)? mem[5573] : 
                       (N722)? mem[5589] : 
                       (N724)? mem[5605] : 
                       (N726)? mem[5621] : 
                       (N728)? mem[5637] : 
                       (N730)? mem[5653] : 
                       (N732)? mem[5669] : 
                       (N734)? mem[5685] : 
                       (N736)? mem[5701] : 
                       (N738)? mem[5717] : 
                       (N740)? mem[5733] : 
                       (N742)? mem[5749] : 
                       (N744)? mem[5765] : 
                       (N746)? mem[5781] : 
                       (N748)? mem[5797] : 
                       (N750)? mem[5813] : 
                       (N752)? mem[5829] : 
                       (N754)? mem[5845] : 
                       (N756)? mem[5861] : 
                       (N758)? mem[5877] : 
                       (N760)? mem[5893] : 
                       (N762)? mem[5909] : 
                       (N764)? mem[5925] : 
                       (N766)? mem[5941] : 
                       (N768)? mem[5957] : 
                       (N770)? mem[5973] : 
                       (N772)? mem[5989] : 
                       (N774)? mem[6005] : 
                       (N776)? mem[6021] : 
                       (N778)? mem[6037] : 
                       (N780)? mem[6053] : 
                       (N782)? mem[6069] : 
                       (N784)? mem[6085] : 
                       (N786)? mem[6101] : 
                       (N788)? mem[6117] : 
                       (N790)? mem[6133] : 
                       (N792)? mem[6149] : 
                       (N794)? mem[6165] : 
                       (N796)? mem[6181] : 
                       (N798)? mem[6197] : 
                       (N800)? mem[6213] : 
                       (N802)? mem[6229] : 
                       (N804)? mem[6245] : 
                       (N806)? mem[6261] : 
                       (N808)? mem[6277] : 
                       (N810)? mem[6293] : 
                       (N812)? mem[6309] : 
                       (N814)? mem[6325] : 
                       (N816)? mem[6341] : 
                       (N818)? mem[6357] : 
                       (N820)? mem[6373] : 
                       (N822)? mem[6389] : 
                       (N824)? mem[6405] : 
                       (N826)? mem[6421] : 
                       (N828)? mem[6437] : 
                       (N830)? mem[6453] : 
                       (N832)? mem[6469] : 
                       (N834)? mem[6485] : 
                       (N836)? mem[6501] : 
                       (N838)? mem[6517] : 
                       (N840)? mem[6533] : 
                       (N842)? mem[6549] : 
                       (N844)? mem[6565] : 
                       (N846)? mem[6581] : 
                       (N848)? mem[6597] : 
                       (N850)? mem[6613] : 
                       (N852)? mem[6629] : 
                       (N854)? mem[6645] : 
                       (N856)? mem[6661] : 
                       (N858)? mem[6677] : 
                       (N860)? mem[6693] : 
                       (N862)? mem[6709] : 
                       (N864)? mem[6725] : 
                       (N866)? mem[6741] : 
                       (N868)? mem[6757] : 
                       (N870)? mem[6773] : 
                       (N872)? mem[6789] : 
                       (N874)? mem[6805] : 
                       (N876)? mem[6821] : 
                       (N878)? mem[6837] : 
                       (N880)? mem[6853] : 
                       (N882)? mem[6869] : 
                       (N884)? mem[6885] : 
                       (N886)? mem[6901] : 
                       (N888)? mem[6917] : 
                       (N890)? mem[6933] : 
                       (N892)? mem[6949] : 
                       (N894)? mem[6965] : 
                       (N896)? mem[6981] : 
                       (N898)? mem[6997] : 
                       (N900)? mem[7013] : 
                       (N902)? mem[7029] : 
                       (N904)? mem[7045] : 
                       (N906)? mem[7061] : 
                       (N908)? mem[7077] : 
                       (N910)? mem[7093] : 
                       (N912)? mem[7109] : 
                       (N914)? mem[7125] : 
                       (N916)? mem[7141] : 
                       (N918)? mem[7157] : 
                       (N920)? mem[7173] : 
                       (N922)? mem[7189] : 
                       (N924)? mem[7205] : 
                       (N926)? mem[7221] : 
                       (N928)? mem[7237] : 
                       (N930)? mem[7253] : 
                       (N932)? mem[7269] : 
                       (N934)? mem[7285] : 
                       (N936)? mem[7301] : 
                       (N938)? mem[7317] : 
                       (N940)? mem[7333] : 
                       (N942)? mem[7349] : 
                       (N944)? mem[7365] : 
                       (N946)? mem[7381] : 
                       (N948)? mem[7397] : 
                       (N950)? mem[7413] : 
                       (N952)? mem[7429] : 
                       (N954)? mem[7445] : 
                       (N956)? mem[7461] : 
                       (N958)? mem[7477] : 
                       (N960)? mem[7493] : 
                       (N962)? mem[7509] : 
                       (N964)? mem[7525] : 
                       (N966)? mem[7541] : 
                       (N968)? mem[7557] : 
                       (N970)? mem[7573] : 
                       (N972)? mem[7589] : 
                       (N974)? mem[7605] : 
                       (N976)? mem[7621] : 
                       (N978)? mem[7637] : 
                       (N980)? mem[7653] : 
                       (N982)? mem[7669] : 
                       (N984)? mem[7685] : 
                       (N986)? mem[7701] : 
                       (N988)? mem[7717] : 
                       (N990)? mem[7733] : 
                       (N992)? mem[7749] : 
                       (N994)? mem[7765] : 
                       (N996)? mem[7781] : 
                       (N998)? mem[7797] : 
                       (N1000)? mem[7813] : 
                       (N1002)? mem[7829] : 
                       (N1004)? mem[7845] : 
                       (N1006)? mem[7861] : 
                       (N1008)? mem[7877] : 
                       (N1010)? mem[7893] : 
                       (N1012)? mem[7909] : 
                       (N1014)? mem[7925] : 
                       (N1016)? mem[7941] : 
                       (N1018)? mem[7957] : 
                       (N1020)? mem[7973] : 
                       (N1022)? mem[7989] : 
                       (N1024)? mem[8005] : 
                       (N1026)? mem[8021] : 
                       (N1028)? mem[8037] : 
                       (N1030)? mem[8053] : 
                       (N1032)? mem[8069] : 
                       (N1034)? mem[8085] : 
                       (N1036)? mem[8101] : 
                       (N1038)? mem[8117] : 
                       (N1040)? mem[8133] : 
                       (N1042)? mem[8149] : 
                       (N1044)? mem[8165] : 
                       (N1046)? mem[8181] : 1'b0;
  assign r_data_o[4] = (N535)? mem[4] : 
                       (N537)? mem[20] : 
                       (N539)? mem[36] : 
                       (N541)? mem[52] : 
                       (N543)? mem[68] : 
                       (N545)? mem[84] : 
                       (N547)? mem[100] : 
                       (N549)? mem[116] : 
                       (N551)? mem[132] : 
                       (N553)? mem[148] : 
                       (N555)? mem[164] : 
                       (N557)? mem[180] : 
                       (N559)? mem[196] : 
                       (N561)? mem[212] : 
                       (N563)? mem[228] : 
                       (N565)? mem[244] : 
                       (N567)? mem[260] : 
                       (N569)? mem[276] : 
                       (N571)? mem[292] : 
                       (N573)? mem[308] : 
                       (N575)? mem[324] : 
                       (N577)? mem[340] : 
                       (N579)? mem[356] : 
                       (N581)? mem[372] : 
                       (N583)? mem[388] : 
                       (N585)? mem[404] : 
                       (N587)? mem[420] : 
                       (N589)? mem[436] : 
                       (N591)? mem[452] : 
                       (N593)? mem[468] : 
                       (N595)? mem[484] : 
                       (N597)? mem[500] : 
                       (N599)? mem[516] : 
                       (N601)? mem[532] : 
                       (N603)? mem[548] : 
                       (N605)? mem[564] : 
                       (N607)? mem[580] : 
                       (N609)? mem[596] : 
                       (N611)? mem[612] : 
                       (N613)? mem[628] : 
                       (N615)? mem[644] : 
                       (N617)? mem[660] : 
                       (N619)? mem[676] : 
                       (N621)? mem[692] : 
                       (N623)? mem[708] : 
                       (N625)? mem[724] : 
                       (N627)? mem[740] : 
                       (N629)? mem[756] : 
                       (N631)? mem[772] : 
                       (N633)? mem[788] : 
                       (N635)? mem[804] : 
                       (N637)? mem[820] : 
                       (N639)? mem[836] : 
                       (N641)? mem[852] : 
                       (N643)? mem[868] : 
                       (N645)? mem[884] : 
                       (N647)? mem[900] : 
                       (N649)? mem[916] : 
                       (N651)? mem[932] : 
                       (N653)? mem[948] : 
                       (N655)? mem[964] : 
                       (N657)? mem[980] : 
                       (N659)? mem[996] : 
                       (N661)? mem[1012] : 
                       (N663)? mem[1028] : 
                       (N665)? mem[1044] : 
                       (N667)? mem[1060] : 
                       (N669)? mem[1076] : 
                       (N671)? mem[1092] : 
                       (N673)? mem[1108] : 
                       (N675)? mem[1124] : 
                       (N677)? mem[1140] : 
                       (N679)? mem[1156] : 
                       (N681)? mem[1172] : 
                       (N683)? mem[1188] : 
                       (N685)? mem[1204] : 
                       (N687)? mem[1220] : 
                       (N689)? mem[1236] : 
                       (N691)? mem[1252] : 
                       (N693)? mem[1268] : 
                       (N695)? mem[1284] : 
                       (N697)? mem[1300] : 
                       (N699)? mem[1316] : 
                       (N701)? mem[1332] : 
                       (N703)? mem[1348] : 
                       (N705)? mem[1364] : 
                       (N707)? mem[1380] : 
                       (N709)? mem[1396] : 
                       (N711)? mem[1412] : 
                       (N713)? mem[1428] : 
                       (N715)? mem[1444] : 
                       (N717)? mem[1460] : 
                       (N719)? mem[1476] : 
                       (N721)? mem[1492] : 
                       (N723)? mem[1508] : 
                       (N725)? mem[1524] : 
                       (N727)? mem[1540] : 
                       (N729)? mem[1556] : 
                       (N731)? mem[1572] : 
                       (N733)? mem[1588] : 
                       (N735)? mem[1604] : 
                       (N737)? mem[1620] : 
                       (N739)? mem[1636] : 
                       (N741)? mem[1652] : 
                       (N743)? mem[1668] : 
                       (N745)? mem[1684] : 
                       (N747)? mem[1700] : 
                       (N749)? mem[1716] : 
                       (N751)? mem[1732] : 
                       (N753)? mem[1748] : 
                       (N755)? mem[1764] : 
                       (N757)? mem[1780] : 
                       (N759)? mem[1796] : 
                       (N761)? mem[1812] : 
                       (N763)? mem[1828] : 
                       (N765)? mem[1844] : 
                       (N767)? mem[1860] : 
                       (N769)? mem[1876] : 
                       (N771)? mem[1892] : 
                       (N773)? mem[1908] : 
                       (N775)? mem[1924] : 
                       (N777)? mem[1940] : 
                       (N779)? mem[1956] : 
                       (N781)? mem[1972] : 
                       (N783)? mem[1988] : 
                       (N785)? mem[2004] : 
                       (N787)? mem[2020] : 
                       (N789)? mem[2036] : 
                       (N791)? mem[2052] : 
                       (N793)? mem[2068] : 
                       (N795)? mem[2084] : 
                       (N797)? mem[2100] : 
                       (N799)? mem[2116] : 
                       (N801)? mem[2132] : 
                       (N803)? mem[2148] : 
                       (N805)? mem[2164] : 
                       (N807)? mem[2180] : 
                       (N809)? mem[2196] : 
                       (N811)? mem[2212] : 
                       (N813)? mem[2228] : 
                       (N815)? mem[2244] : 
                       (N817)? mem[2260] : 
                       (N819)? mem[2276] : 
                       (N821)? mem[2292] : 
                       (N823)? mem[2308] : 
                       (N825)? mem[2324] : 
                       (N827)? mem[2340] : 
                       (N829)? mem[2356] : 
                       (N831)? mem[2372] : 
                       (N833)? mem[2388] : 
                       (N835)? mem[2404] : 
                       (N837)? mem[2420] : 
                       (N839)? mem[2436] : 
                       (N841)? mem[2452] : 
                       (N843)? mem[2468] : 
                       (N845)? mem[2484] : 
                       (N847)? mem[2500] : 
                       (N849)? mem[2516] : 
                       (N851)? mem[2532] : 
                       (N853)? mem[2548] : 
                       (N855)? mem[2564] : 
                       (N857)? mem[2580] : 
                       (N859)? mem[2596] : 
                       (N861)? mem[2612] : 
                       (N863)? mem[2628] : 
                       (N865)? mem[2644] : 
                       (N867)? mem[2660] : 
                       (N869)? mem[2676] : 
                       (N871)? mem[2692] : 
                       (N873)? mem[2708] : 
                       (N875)? mem[2724] : 
                       (N877)? mem[2740] : 
                       (N879)? mem[2756] : 
                       (N881)? mem[2772] : 
                       (N883)? mem[2788] : 
                       (N885)? mem[2804] : 
                       (N887)? mem[2820] : 
                       (N889)? mem[2836] : 
                       (N891)? mem[2852] : 
                       (N893)? mem[2868] : 
                       (N895)? mem[2884] : 
                       (N897)? mem[2900] : 
                       (N899)? mem[2916] : 
                       (N901)? mem[2932] : 
                       (N903)? mem[2948] : 
                       (N905)? mem[2964] : 
                       (N907)? mem[2980] : 
                       (N909)? mem[2996] : 
                       (N911)? mem[3012] : 
                       (N913)? mem[3028] : 
                       (N915)? mem[3044] : 
                       (N917)? mem[3060] : 
                       (N919)? mem[3076] : 
                       (N921)? mem[3092] : 
                       (N923)? mem[3108] : 
                       (N925)? mem[3124] : 
                       (N927)? mem[3140] : 
                       (N929)? mem[3156] : 
                       (N931)? mem[3172] : 
                       (N933)? mem[3188] : 
                       (N935)? mem[3204] : 
                       (N937)? mem[3220] : 
                       (N939)? mem[3236] : 
                       (N941)? mem[3252] : 
                       (N943)? mem[3268] : 
                       (N945)? mem[3284] : 
                       (N947)? mem[3300] : 
                       (N949)? mem[3316] : 
                       (N951)? mem[3332] : 
                       (N953)? mem[3348] : 
                       (N955)? mem[3364] : 
                       (N957)? mem[3380] : 
                       (N959)? mem[3396] : 
                       (N961)? mem[3412] : 
                       (N963)? mem[3428] : 
                       (N965)? mem[3444] : 
                       (N967)? mem[3460] : 
                       (N969)? mem[3476] : 
                       (N971)? mem[3492] : 
                       (N973)? mem[3508] : 
                       (N975)? mem[3524] : 
                       (N977)? mem[3540] : 
                       (N979)? mem[3556] : 
                       (N981)? mem[3572] : 
                       (N983)? mem[3588] : 
                       (N985)? mem[3604] : 
                       (N987)? mem[3620] : 
                       (N989)? mem[3636] : 
                       (N991)? mem[3652] : 
                       (N993)? mem[3668] : 
                       (N995)? mem[3684] : 
                       (N997)? mem[3700] : 
                       (N999)? mem[3716] : 
                       (N1001)? mem[3732] : 
                       (N1003)? mem[3748] : 
                       (N1005)? mem[3764] : 
                       (N1007)? mem[3780] : 
                       (N1009)? mem[3796] : 
                       (N1011)? mem[3812] : 
                       (N1013)? mem[3828] : 
                       (N1015)? mem[3844] : 
                       (N1017)? mem[3860] : 
                       (N1019)? mem[3876] : 
                       (N1021)? mem[3892] : 
                       (N1023)? mem[3908] : 
                       (N1025)? mem[3924] : 
                       (N1027)? mem[3940] : 
                       (N1029)? mem[3956] : 
                       (N1031)? mem[3972] : 
                       (N1033)? mem[3988] : 
                       (N1035)? mem[4004] : 
                       (N1037)? mem[4020] : 
                       (N1039)? mem[4036] : 
                       (N1041)? mem[4052] : 
                       (N1043)? mem[4068] : 
                       (N1045)? mem[4084] : 
                       (N536)? mem[4100] : 
                       (N538)? mem[4116] : 
                       (N540)? mem[4132] : 
                       (N542)? mem[4148] : 
                       (N544)? mem[4164] : 
                       (N546)? mem[4180] : 
                       (N548)? mem[4196] : 
                       (N550)? mem[4212] : 
                       (N552)? mem[4228] : 
                       (N554)? mem[4244] : 
                       (N556)? mem[4260] : 
                       (N558)? mem[4276] : 
                       (N560)? mem[4292] : 
                       (N562)? mem[4308] : 
                       (N564)? mem[4324] : 
                       (N566)? mem[4340] : 
                       (N568)? mem[4356] : 
                       (N570)? mem[4372] : 
                       (N572)? mem[4388] : 
                       (N574)? mem[4404] : 
                       (N576)? mem[4420] : 
                       (N578)? mem[4436] : 
                       (N580)? mem[4452] : 
                       (N582)? mem[4468] : 
                       (N584)? mem[4484] : 
                       (N586)? mem[4500] : 
                       (N588)? mem[4516] : 
                       (N590)? mem[4532] : 
                       (N592)? mem[4548] : 
                       (N594)? mem[4564] : 
                       (N596)? mem[4580] : 
                       (N598)? mem[4596] : 
                       (N600)? mem[4612] : 
                       (N602)? mem[4628] : 
                       (N604)? mem[4644] : 
                       (N606)? mem[4660] : 
                       (N608)? mem[4676] : 
                       (N610)? mem[4692] : 
                       (N612)? mem[4708] : 
                       (N614)? mem[4724] : 
                       (N616)? mem[4740] : 
                       (N618)? mem[4756] : 
                       (N620)? mem[4772] : 
                       (N622)? mem[4788] : 
                       (N624)? mem[4804] : 
                       (N626)? mem[4820] : 
                       (N628)? mem[4836] : 
                       (N630)? mem[4852] : 
                       (N632)? mem[4868] : 
                       (N634)? mem[4884] : 
                       (N636)? mem[4900] : 
                       (N638)? mem[4916] : 
                       (N640)? mem[4932] : 
                       (N642)? mem[4948] : 
                       (N644)? mem[4964] : 
                       (N646)? mem[4980] : 
                       (N648)? mem[4996] : 
                       (N650)? mem[5012] : 
                       (N652)? mem[5028] : 
                       (N654)? mem[5044] : 
                       (N656)? mem[5060] : 
                       (N658)? mem[5076] : 
                       (N660)? mem[5092] : 
                       (N662)? mem[5108] : 
                       (N664)? mem[5124] : 
                       (N666)? mem[5140] : 
                       (N668)? mem[5156] : 
                       (N670)? mem[5172] : 
                       (N672)? mem[5188] : 
                       (N674)? mem[5204] : 
                       (N676)? mem[5220] : 
                       (N678)? mem[5236] : 
                       (N680)? mem[5252] : 
                       (N682)? mem[5268] : 
                       (N684)? mem[5284] : 
                       (N686)? mem[5300] : 
                       (N688)? mem[5316] : 
                       (N690)? mem[5332] : 
                       (N692)? mem[5348] : 
                       (N694)? mem[5364] : 
                       (N696)? mem[5380] : 
                       (N698)? mem[5396] : 
                       (N700)? mem[5412] : 
                       (N702)? mem[5428] : 
                       (N704)? mem[5444] : 
                       (N706)? mem[5460] : 
                       (N708)? mem[5476] : 
                       (N710)? mem[5492] : 
                       (N712)? mem[5508] : 
                       (N714)? mem[5524] : 
                       (N716)? mem[5540] : 
                       (N718)? mem[5556] : 
                       (N720)? mem[5572] : 
                       (N722)? mem[5588] : 
                       (N724)? mem[5604] : 
                       (N726)? mem[5620] : 
                       (N728)? mem[5636] : 
                       (N730)? mem[5652] : 
                       (N732)? mem[5668] : 
                       (N734)? mem[5684] : 
                       (N736)? mem[5700] : 
                       (N738)? mem[5716] : 
                       (N740)? mem[5732] : 
                       (N742)? mem[5748] : 
                       (N744)? mem[5764] : 
                       (N746)? mem[5780] : 
                       (N748)? mem[5796] : 
                       (N750)? mem[5812] : 
                       (N752)? mem[5828] : 
                       (N754)? mem[5844] : 
                       (N756)? mem[5860] : 
                       (N758)? mem[5876] : 
                       (N760)? mem[5892] : 
                       (N762)? mem[5908] : 
                       (N764)? mem[5924] : 
                       (N766)? mem[5940] : 
                       (N768)? mem[5956] : 
                       (N770)? mem[5972] : 
                       (N772)? mem[5988] : 
                       (N774)? mem[6004] : 
                       (N776)? mem[6020] : 
                       (N778)? mem[6036] : 
                       (N780)? mem[6052] : 
                       (N782)? mem[6068] : 
                       (N784)? mem[6084] : 
                       (N786)? mem[6100] : 
                       (N788)? mem[6116] : 
                       (N790)? mem[6132] : 
                       (N792)? mem[6148] : 
                       (N794)? mem[6164] : 
                       (N796)? mem[6180] : 
                       (N798)? mem[6196] : 
                       (N800)? mem[6212] : 
                       (N802)? mem[6228] : 
                       (N804)? mem[6244] : 
                       (N806)? mem[6260] : 
                       (N808)? mem[6276] : 
                       (N810)? mem[6292] : 
                       (N812)? mem[6308] : 
                       (N814)? mem[6324] : 
                       (N816)? mem[6340] : 
                       (N818)? mem[6356] : 
                       (N820)? mem[6372] : 
                       (N822)? mem[6388] : 
                       (N824)? mem[6404] : 
                       (N826)? mem[6420] : 
                       (N828)? mem[6436] : 
                       (N830)? mem[6452] : 
                       (N832)? mem[6468] : 
                       (N834)? mem[6484] : 
                       (N836)? mem[6500] : 
                       (N838)? mem[6516] : 
                       (N840)? mem[6532] : 
                       (N842)? mem[6548] : 
                       (N844)? mem[6564] : 
                       (N846)? mem[6580] : 
                       (N848)? mem[6596] : 
                       (N850)? mem[6612] : 
                       (N852)? mem[6628] : 
                       (N854)? mem[6644] : 
                       (N856)? mem[6660] : 
                       (N858)? mem[6676] : 
                       (N860)? mem[6692] : 
                       (N862)? mem[6708] : 
                       (N864)? mem[6724] : 
                       (N866)? mem[6740] : 
                       (N868)? mem[6756] : 
                       (N870)? mem[6772] : 
                       (N872)? mem[6788] : 
                       (N874)? mem[6804] : 
                       (N876)? mem[6820] : 
                       (N878)? mem[6836] : 
                       (N880)? mem[6852] : 
                       (N882)? mem[6868] : 
                       (N884)? mem[6884] : 
                       (N886)? mem[6900] : 
                       (N888)? mem[6916] : 
                       (N890)? mem[6932] : 
                       (N892)? mem[6948] : 
                       (N894)? mem[6964] : 
                       (N896)? mem[6980] : 
                       (N898)? mem[6996] : 
                       (N900)? mem[7012] : 
                       (N902)? mem[7028] : 
                       (N904)? mem[7044] : 
                       (N906)? mem[7060] : 
                       (N908)? mem[7076] : 
                       (N910)? mem[7092] : 
                       (N912)? mem[7108] : 
                       (N914)? mem[7124] : 
                       (N916)? mem[7140] : 
                       (N918)? mem[7156] : 
                       (N920)? mem[7172] : 
                       (N922)? mem[7188] : 
                       (N924)? mem[7204] : 
                       (N926)? mem[7220] : 
                       (N928)? mem[7236] : 
                       (N930)? mem[7252] : 
                       (N932)? mem[7268] : 
                       (N934)? mem[7284] : 
                       (N936)? mem[7300] : 
                       (N938)? mem[7316] : 
                       (N940)? mem[7332] : 
                       (N942)? mem[7348] : 
                       (N944)? mem[7364] : 
                       (N946)? mem[7380] : 
                       (N948)? mem[7396] : 
                       (N950)? mem[7412] : 
                       (N952)? mem[7428] : 
                       (N954)? mem[7444] : 
                       (N956)? mem[7460] : 
                       (N958)? mem[7476] : 
                       (N960)? mem[7492] : 
                       (N962)? mem[7508] : 
                       (N964)? mem[7524] : 
                       (N966)? mem[7540] : 
                       (N968)? mem[7556] : 
                       (N970)? mem[7572] : 
                       (N972)? mem[7588] : 
                       (N974)? mem[7604] : 
                       (N976)? mem[7620] : 
                       (N978)? mem[7636] : 
                       (N980)? mem[7652] : 
                       (N982)? mem[7668] : 
                       (N984)? mem[7684] : 
                       (N986)? mem[7700] : 
                       (N988)? mem[7716] : 
                       (N990)? mem[7732] : 
                       (N992)? mem[7748] : 
                       (N994)? mem[7764] : 
                       (N996)? mem[7780] : 
                       (N998)? mem[7796] : 
                       (N1000)? mem[7812] : 
                       (N1002)? mem[7828] : 
                       (N1004)? mem[7844] : 
                       (N1006)? mem[7860] : 
                       (N1008)? mem[7876] : 
                       (N1010)? mem[7892] : 
                       (N1012)? mem[7908] : 
                       (N1014)? mem[7924] : 
                       (N1016)? mem[7940] : 
                       (N1018)? mem[7956] : 
                       (N1020)? mem[7972] : 
                       (N1022)? mem[7988] : 
                       (N1024)? mem[8004] : 
                       (N1026)? mem[8020] : 
                       (N1028)? mem[8036] : 
                       (N1030)? mem[8052] : 
                       (N1032)? mem[8068] : 
                       (N1034)? mem[8084] : 
                       (N1036)? mem[8100] : 
                       (N1038)? mem[8116] : 
                       (N1040)? mem[8132] : 
                       (N1042)? mem[8148] : 
                       (N1044)? mem[8164] : 
                       (N1046)? mem[8180] : 1'b0;
  assign r_data_o[3] = (N535)? mem[3] : 
                       (N537)? mem[19] : 
                       (N539)? mem[35] : 
                       (N541)? mem[51] : 
                       (N543)? mem[67] : 
                       (N545)? mem[83] : 
                       (N547)? mem[99] : 
                       (N549)? mem[115] : 
                       (N551)? mem[131] : 
                       (N553)? mem[147] : 
                       (N555)? mem[163] : 
                       (N557)? mem[179] : 
                       (N559)? mem[195] : 
                       (N561)? mem[211] : 
                       (N563)? mem[227] : 
                       (N565)? mem[243] : 
                       (N567)? mem[259] : 
                       (N569)? mem[275] : 
                       (N571)? mem[291] : 
                       (N573)? mem[307] : 
                       (N575)? mem[323] : 
                       (N577)? mem[339] : 
                       (N579)? mem[355] : 
                       (N581)? mem[371] : 
                       (N583)? mem[387] : 
                       (N585)? mem[403] : 
                       (N587)? mem[419] : 
                       (N589)? mem[435] : 
                       (N591)? mem[451] : 
                       (N593)? mem[467] : 
                       (N595)? mem[483] : 
                       (N597)? mem[499] : 
                       (N599)? mem[515] : 
                       (N601)? mem[531] : 
                       (N603)? mem[547] : 
                       (N605)? mem[563] : 
                       (N607)? mem[579] : 
                       (N609)? mem[595] : 
                       (N611)? mem[611] : 
                       (N613)? mem[627] : 
                       (N615)? mem[643] : 
                       (N617)? mem[659] : 
                       (N619)? mem[675] : 
                       (N621)? mem[691] : 
                       (N623)? mem[707] : 
                       (N625)? mem[723] : 
                       (N627)? mem[739] : 
                       (N629)? mem[755] : 
                       (N631)? mem[771] : 
                       (N633)? mem[787] : 
                       (N635)? mem[803] : 
                       (N637)? mem[819] : 
                       (N639)? mem[835] : 
                       (N641)? mem[851] : 
                       (N643)? mem[867] : 
                       (N645)? mem[883] : 
                       (N647)? mem[899] : 
                       (N649)? mem[915] : 
                       (N651)? mem[931] : 
                       (N653)? mem[947] : 
                       (N655)? mem[963] : 
                       (N657)? mem[979] : 
                       (N659)? mem[995] : 
                       (N661)? mem[1011] : 
                       (N663)? mem[1027] : 
                       (N665)? mem[1043] : 
                       (N667)? mem[1059] : 
                       (N669)? mem[1075] : 
                       (N671)? mem[1091] : 
                       (N673)? mem[1107] : 
                       (N675)? mem[1123] : 
                       (N677)? mem[1139] : 
                       (N679)? mem[1155] : 
                       (N681)? mem[1171] : 
                       (N683)? mem[1187] : 
                       (N685)? mem[1203] : 
                       (N687)? mem[1219] : 
                       (N689)? mem[1235] : 
                       (N691)? mem[1251] : 
                       (N693)? mem[1267] : 
                       (N695)? mem[1283] : 
                       (N697)? mem[1299] : 
                       (N699)? mem[1315] : 
                       (N701)? mem[1331] : 
                       (N703)? mem[1347] : 
                       (N705)? mem[1363] : 
                       (N707)? mem[1379] : 
                       (N709)? mem[1395] : 
                       (N711)? mem[1411] : 
                       (N713)? mem[1427] : 
                       (N715)? mem[1443] : 
                       (N717)? mem[1459] : 
                       (N719)? mem[1475] : 
                       (N721)? mem[1491] : 
                       (N723)? mem[1507] : 
                       (N725)? mem[1523] : 
                       (N727)? mem[1539] : 
                       (N729)? mem[1555] : 
                       (N731)? mem[1571] : 
                       (N733)? mem[1587] : 
                       (N735)? mem[1603] : 
                       (N737)? mem[1619] : 
                       (N739)? mem[1635] : 
                       (N741)? mem[1651] : 
                       (N743)? mem[1667] : 
                       (N745)? mem[1683] : 
                       (N747)? mem[1699] : 
                       (N749)? mem[1715] : 
                       (N751)? mem[1731] : 
                       (N753)? mem[1747] : 
                       (N755)? mem[1763] : 
                       (N757)? mem[1779] : 
                       (N759)? mem[1795] : 
                       (N761)? mem[1811] : 
                       (N763)? mem[1827] : 
                       (N765)? mem[1843] : 
                       (N767)? mem[1859] : 
                       (N769)? mem[1875] : 
                       (N771)? mem[1891] : 
                       (N773)? mem[1907] : 
                       (N775)? mem[1923] : 
                       (N777)? mem[1939] : 
                       (N779)? mem[1955] : 
                       (N781)? mem[1971] : 
                       (N783)? mem[1987] : 
                       (N785)? mem[2003] : 
                       (N787)? mem[2019] : 
                       (N789)? mem[2035] : 
                       (N791)? mem[2051] : 
                       (N793)? mem[2067] : 
                       (N795)? mem[2083] : 
                       (N797)? mem[2099] : 
                       (N799)? mem[2115] : 
                       (N801)? mem[2131] : 
                       (N803)? mem[2147] : 
                       (N805)? mem[2163] : 
                       (N807)? mem[2179] : 
                       (N809)? mem[2195] : 
                       (N811)? mem[2211] : 
                       (N813)? mem[2227] : 
                       (N815)? mem[2243] : 
                       (N817)? mem[2259] : 
                       (N819)? mem[2275] : 
                       (N821)? mem[2291] : 
                       (N823)? mem[2307] : 
                       (N825)? mem[2323] : 
                       (N827)? mem[2339] : 
                       (N829)? mem[2355] : 
                       (N831)? mem[2371] : 
                       (N833)? mem[2387] : 
                       (N835)? mem[2403] : 
                       (N837)? mem[2419] : 
                       (N839)? mem[2435] : 
                       (N841)? mem[2451] : 
                       (N843)? mem[2467] : 
                       (N845)? mem[2483] : 
                       (N847)? mem[2499] : 
                       (N849)? mem[2515] : 
                       (N851)? mem[2531] : 
                       (N853)? mem[2547] : 
                       (N855)? mem[2563] : 
                       (N857)? mem[2579] : 
                       (N859)? mem[2595] : 
                       (N861)? mem[2611] : 
                       (N863)? mem[2627] : 
                       (N865)? mem[2643] : 
                       (N867)? mem[2659] : 
                       (N869)? mem[2675] : 
                       (N871)? mem[2691] : 
                       (N873)? mem[2707] : 
                       (N875)? mem[2723] : 
                       (N877)? mem[2739] : 
                       (N879)? mem[2755] : 
                       (N881)? mem[2771] : 
                       (N883)? mem[2787] : 
                       (N885)? mem[2803] : 
                       (N887)? mem[2819] : 
                       (N889)? mem[2835] : 
                       (N891)? mem[2851] : 
                       (N893)? mem[2867] : 
                       (N895)? mem[2883] : 
                       (N897)? mem[2899] : 
                       (N899)? mem[2915] : 
                       (N901)? mem[2931] : 
                       (N903)? mem[2947] : 
                       (N905)? mem[2963] : 
                       (N907)? mem[2979] : 
                       (N909)? mem[2995] : 
                       (N911)? mem[3011] : 
                       (N913)? mem[3027] : 
                       (N915)? mem[3043] : 
                       (N917)? mem[3059] : 
                       (N919)? mem[3075] : 
                       (N921)? mem[3091] : 
                       (N923)? mem[3107] : 
                       (N925)? mem[3123] : 
                       (N927)? mem[3139] : 
                       (N929)? mem[3155] : 
                       (N931)? mem[3171] : 
                       (N933)? mem[3187] : 
                       (N935)? mem[3203] : 
                       (N937)? mem[3219] : 
                       (N939)? mem[3235] : 
                       (N941)? mem[3251] : 
                       (N943)? mem[3267] : 
                       (N945)? mem[3283] : 
                       (N947)? mem[3299] : 
                       (N949)? mem[3315] : 
                       (N951)? mem[3331] : 
                       (N953)? mem[3347] : 
                       (N955)? mem[3363] : 
                       (N957)? mem[3379] : 
                       (N959)? mem[3395] : 
                       (N961)? mem[3411] : 
                       (N963)? mem[3427] : 
                       (N965)? mem[3443] : 
                       (N967)? mem[3459] : 
                       (N969)? mem[3475] : 
                       (N971)? mem[3491] : 
                       (N973)? mem[3507] : 
                       (N975)? mem[3523] : 
                       (N977)? mem[3539] : 
                       (N979)? mem[3555] : 
                       (N981)? mem[3571] : 
                       (N983)? mem[3587] : 
                       (N985)? mem[3603] : 
                       (N987)? mem[3619] : 
                       (N989)? mem[3635] : 
                       (N991)? mem[3651] : 
                       (N993)? mem[3667] : 
                       (N995)? mem[3683] : 
                       (N997)? mem[3699] : 
                       (N999)? mem[3715] : 
                       (N1001)? mem[3731] : 
                       (N1003)? mem[3747] : 
                       (N1005)? mem[3763] : 
                       (N1007)? mem[3779] : 
                       (N1009)? mem[3795] : 
                       (N1011)? mem[3811] : 
                       (N1013)? mem[3827] : 
                       (N1015)? mem[3843] : 
                       (N1017)? mem[3859] : 
                       (N1019)? mem[3875] : 
                       (N1021)? mem[3891] : 
                       (N1023)? mem[3907] : 
                       (N1025)? mem[3923] : 
                       (N1027)? mem[3939] : 
                       (N1029)? mem[3955] : 
                       (N1031)? mem[3971] : 
                       (N1033)? mem[3987] : 
                       (N1035)? mem[4003] : 
                       (N1037)? mem[4019] : 
                       (N1039)? mem[4035] : 
                       (N1041)? mem[4051] : 
                       (N1043)? mem[4067] : 
                       (N1045)? mem[4083] : 
                       (N536)? mem[4099] : 
                       (N538)? mem[4115] : 
                       (N540)? mem[4131] : 
                       (N542)? mem[4147] : 
                       (N544)? mem[4163] : 
                       (N546)? mem[4179] : 
                       (N548)? mem[4195] : 
                       (N550)? mem[4211] : 
                       (N552)? mem[4227] : 
                       (N554)? mem[4243] : 
                       (N556)? mem[4259] : 
                       (N558)? mem[4275] : 
                       (N560)? mem[4291] : 
                       (N562)? mem[4307] : 
                       (N564)? mem[4323] : 
                       (N566)? mem[4339] : 
                       (N568)? mem[4355] : 
                       (N570)? mem[4371] : 
                       (N572)? mem[4387] : 
                       (N574)? mem[4403] : 
                       (N576)? mem[4419] : 
                       (N578)? mem[4435] : 
                       (N580)? mem[4451] : 
                       (N582)? mem[4467] : 
                       (N584)? mem[4483] : 
                       (N586)? mem[4499] : 
                       (N588)? mem[4515] : 
                       (N590)? mem[4531] : 
                       (N592)? mem[4547] : 
                       (N594)? mem[4563] : 
                       (N596)? mem[4579] : 
                       (N598)? mem[4595] : 
                       (N600)? mem[4611] : 
                       (N602)? mem[4627] : 
                       (N604)? mem[4643] : 
                       (N606)? mem[4659] : 
                       (N608)? mem[4675] : 
                       (N610)? mem[4691] : 
                       (N612)? mem[4707] : 
                       (N614)? mem[4723] : 
                       (N616)? mem[4739] : 
                       (N618)? mem[4755] : 
                       (N620)? mem[4771] : 
                       (N622)? mem[4787] : 
                       (N624)? mem[4803] : 
                       (N626)? mem[4819] : 
                       (N628)? mem[4835] : 
                       (N630)? mem[4851] : 
                       (N632)? mem[4867] : 
                       (N634)? mem[4883] : 
                       (N636)? mem[4899] : 
                       (N638)? mem[4915] : 
                       (N640)? mem[4931] : 
                       (N642)? mem[4947] : 
                       (N644)? mem[4963] : 
                       (N646)? mem[4979] : 
                       (N648)? mem[4995] : 
                       (N650)? mem[5011] : 
                       (N652)? mem[5027] : 
                       (N654)? mem[5043] : 
                       (N656)? mem[5059] : 
                       (N658)? mem[5075] : 
                       (N660)? mem[5091] : 
                       (N662)? mem[5107] : 
                       (N664)? mem[5123] : 
                       (N666)? mem[5139] : 
                       (N668)? mem[5155] : 
                       (N670)? mem[5171] : 
                       (N672)? mem[5187] : 
                       (N674)? mem[5203] : 
                       (N676)? mem[5219] : 
                       (N678)? mem[5235] : 
                       (N680)? mem[5251] : 
                       (N682)? mem[5267] : 
                       (N684)? mem[5283] : 
                       (N686)? mem[5299] : 
                       (N688)? mem[5315] : 
                       (N690)? mem[5331] : 
                       (N692)? mem[5347] : 
                       (N694)? mem[5363] : 
                       (N696)? mem[5379] : 
                       (N698)? mem[5395] : 
                       (N700)? mem[5411] : 
                       (N702)? mem[5427] : 
                       (N704)? mem[5443] : 
                       (N706)? mem[5459] : 
                       (N708)? mem[5475] : 
                       (N710)? mem[5491] : 
                       (N712)? mem[5507] : 
                       (N714)? mem[5523] : 
                       (N716)? mem[5539] : 
                       (N718)? mem[5555] : 
                       (N720)? mem[5571] : 
                       (N722)? mem[5587] : 
                       (N724)? mem[5603] : 
                       (N726)? mem[5619] : 
                       (N728)? mem[5635] : 
                       (N730)? mem[5651] : 
                       (N732)? mem[5667] : 
                       (N734)? mem[5683] : 
                       (N736)? mem[5699] : 
                       (N738)? mem[5715] : 
                       (N740)? mem[5731] : 
                       (N742)? mem[5747] : 
                       (N744)? mem[5763] : 
                       (N746)? mem[5779] : 
                       (N748)? mem[5795] : 
                       (N750)? mem[5811] : 
                       (N752)? mem[5827] : 
                       (N754)? mem[5843] : 
                       (N756)? mem[5859] : 
                       (N758)? mem[5875] : 
                       (N760)? mem[5891] : 
                       (N762)? mem[5907] : 
                       (N764)? mem[5923] : 
                       (N766)? mem[5939] : 
                       (N768)? mem[5955] : 
                       (N770)? mem[5971] : 
                       (N772)? mem[5987] : 
                       (N774)? mem[6003] : 
                       (N776)? mem[6019] : 
                       (N778)? mem[6035] : 
                       (N780)? mem[6051] : 
                       (N782)? mem[6067] : 
                       (N784)? mem[6083] : 
                       (N786)? mem[6099] : 
                       (N788)? mem[6115] : 
                       (N790)? mem[6131] : 
                       (N792)? mem[6147] : 
                       (N794)? mem[6163] : 
                       (N796)? mem[6179] : 
                       (N798)? mem[6195] : 
                       (N800)? mem[6211] : 
                       (N802)? mem[6227] : 
                       (N804)? mem[6243] : 
                       (N806)? mem[6259] : 
                       (N808)? mem[6275] : 
                       (N810)? mem[6291] : 
                       (N812)? mem[6307] : 
                       (N814)? mem[6323] : 
                       (N816)? mem[6339] : 
                       (N818)? mem[6355] : 
                       (N820)? mem[6371] : 
                       (N822)? mem[6387] : 
                       (N824)? mem[6403] : 
                       (N826)? mem[6419] : 
                       (N828)? mem[6435] : 
                       (N830)? mem[6451] : 
                       (N832)? mem[6467] : 
                       (N834)? mem[6483] : 
                       (N836)? mem[6499] : 
                       (N838)? mem[6515] : 
                       (N840)? mem[6531] : 
                       (N842)? mem[6547] : 
                       (N844)? mem[6563] : 
                       (N846)? mem[6579] : 
                       (N848)? mem[6595] : 
                       (N850)? mem[6611] : 
                       (N852)? mem[6627] : 
                       (N854)? mem[6643] : 
                       (N856)? mem[6659] : 
                       (N858)? mem[6675] : 
                       (N860)? mem[6691] : 
                       (N862)? mem[6707] : 
                       (N864)? mem[6723] : 
                       (N866)? mem[6739] : 
                       (N868)? mem[6755] : 
                       (N870)? mem[6771] : 
                       (N872)? mem[6787] : 
                       (N874)? mem[6803] : 
                       (N876)? mem[6819] : 
                       (N878)? mem[6835] : 
                       (N880)? mem[6851] : 
                       (N882)? mem[6867] : 
                       (N884)? mem[6883] : 
                       (N886)? mem[6899] : 
                       (N888)? mem[6915] : 
                       (N890)? mem[6931] : 
                       (N892)? mem[6947] : 
                       (N894)? mem[6963] : 
                       (N896)? mem[6979] : 
                       (N898)? mem[6995] : 
                       (N900)? mem[7011] : 
                       (N902)? mem[7027] : 
                       (N904)? mem[7043] : 
                       (N906)? mem[7059] : 
                       (N908)? mem[7075] : 
                       (N910)? mem[7091] : 
                       (N912)? mem[7107] : 
                       (N914)? mem[7123] : 
                       (N916)? mem[7139] : 
                       (N918)? mem[7155] : 
                       (N920)? mem[7171] : 
                       (N922)? mem[7187] : 
                       (N924)? mem[7203] : 
                       (N926)? mem[7219] : 
                       (N928)? mem[7235] : 
                       (N930)? mem[7251] : 
                       (N932)? mem[7267] : 
                       (N934)? mem[7283] : 
                       (N936)? mem[7299] : 
                       (N938)? mem[7315] : 
                       (N940)? mem[7331] : 
                       (N942)? mem[7347] : 
                       (N944)? mem[7363] : 
                       (N946)? mem[7379] : 
                       (N948)? mem[7395] : 
                       (N950)? mem[7411] : 
                       (N952)? mem[7427] : 
                       (N954)? mem[7443] : 
                       (N956)? mem[7459] : 
                       (N958)? mem[7475] : 
                       (N960)? mem[7491] : 
                       (N962)? mem[7507] : 
                       (N964)? mem[7523] : 
                       (N966)? mem[7539] : 
                       (N968)? mem[7555] : 
                       (N970)? mem[7571] : 
                       (N972)? mem[7587] : 
                       (N974)? mem[7603] : 
                       (N976)? mem[7619] : 
                       (N978)? mem[7635] : 
                       (N980)? mem[7651] : 
                       (N982)? mem[7667] : 
                       (N984)? mem[7683] : 
                       (N986)? mem[7699] : 
                       (N988)? mem[7715] : 
                       (N990)? mem[7731] : 
                       (N992)? mem[7747] : 
                       (N994)? mem[7763] : 
                       (N996)? mem[7779] : 
                       (N998)? mem[7795] : 
                       (N1000)? mem[7811] : 
                       (N1002)? mem[7827] : 
                       (N1004)? mem[7843] : 
                       (N1006)? mem[7859] : 
                       (N1008)? mem[7875] : 
                       (N1010)? mem[7891] : 
                       (N1012)? mem[7907] : 
                       (N1014)? mem[7923] : 
                       (N1016)? mem[7939] : 
                       (N1018)? mem[7955] : 
                       (N1020)? mem[7971] : 
                       (N1022)? mem[7987] : 
                       (N1024)? mem[8003] : 
                       (N1026)? mem[8019] : 
                       (N1028)? mem[8035] : 
                       (N1030)? mem[8051] : 
                       (N1032)? mem[8067] : 
                       (N1034)? mem[8083] : 
                       (N1036)? mem[8099] : 
                       (N1038)? mem[8115] : 
                       (N1040)? mem[8131] : 
                       (N1042)? mem[8147] : 
                       (N1044)? mem[8163] : 
                       (N1046)? mem[8179] : 1'b0;
  assign r_data_o[2] = (N535)? mem[2] : 
                       (N537)? mem[18] : 
                       (N539)? mem[34] : 
                       (N541)? mem[50] : 
                       (N543)? mem[66] : 
                       (N545)? mem[82] : 
                       (N547)? mem[98] : 
                       (N549)? mem[114] : 
                       (N551)? mem[130] : 
                       (N553)? mem[146] : 
                       (N555)? mem[162] : 
                       (N557)? mem[178] : 
                       (N559)? mem[194] : 
                       (N561)? mem[210] : 
                       (N563)? mem[226] : 
                       (N565)? mem[242] : 
                       (N567)? mem[258] : 
                       (N569)? mem[274] : 
                       (N571)? mem[290] : 
                       (N573)? mem[306] : 
                       (N575)? mem[322] : 
                       (N577)? mem[338] : 
                       (N579)? mem[354] : 
                       (N581)? mem[370] : 
                       (N583)? mem[386] : 
                       (N585)? mem[402] : 
                       (N587)? mem[418] : 
                       (N589)? mem[434] : 
                       (N591)? mem[450] : 
                       (N593)? mem[466] : 
                       (N595)? mem[482] : 
                       (N597)? mem[498] : 
                       (N599)? mem[514] : 
                       (N601)? mem[530] : 
                       (N603)? mem[546] : 
                       (N605)? mem[562] : 
                       (N607)? mem[578] : 
                       (N609)? mem[594] : 
                       (N611)? mem[610] : 
                       (N613)? mem[626] : 
                       (N615)? mem[642] : 
                       (N617)? mem[658] : 
                       (N619)? mem[674] : 
                       (N621)? mem[690] : 
                       (N623)? mem[706] : 
                       (N625)? mem[722] : 
                       (N627)? mem[738] : 
                       (N629)? mem[754] : 
                       (N631)? mem[770] : 
                       (N633)? mem[786] : 
                       (N635)? mem[802] : 
                       (N637)? mem[818] : 
                       (N639)? mem[834] : 
                       (N641)? mem[850] : 
                       (N643)? mem[866] : 
                       (N645)? mem[882] : 
                       (N647)? mem[898] : 
                       (N649)? mem[914] : 
                       (N651)? mem[930] : 
                       (N653)? mem[946] : 
                       (N655)? mem[962] : 
                       (N657)? mem[978] : 
                       (N659)? mem[994] : 
                       (N661)? mem[1010] : 
                       (N663)? mem[1026] : 
                       (N665)? mem[1042] : 
                       (N667)? mem[1058] : 
                       (N669)? mem[1074] : 
                       (N671)? mem[1090] : 
                       (N673)? mem[1106] : 
                       (N675)? mem[1122] : 
                       (N677)? mem[1138] : 
                       (N679)? mem[1154] : 
                       (N681)? mem[1170] : 
                       (N683)? mem[1186] : 
                       (N685)? mem[1202] : 
                       (N687)? mem[1218] : 
                       (N689)? mem[1234] : 
                       (N691)? mem[1250] : 
                       (N693)? mem[1266] : 
                       (N695)? mem[1282] : 
                       (N697)? mem[1298] : 
                       (N699)? mem[1314] : 
                       (N701)? mem[1330] : 
                       (N703)? mem[1346] : 
                       (N705)? mem[1362] : 
                       (N707)? mem[1378] : 
                       (N709)? mem[1394] : 
                       (N711)? mem[1410] : 
                       (N713)? mem[1426] : 
                       (N715)? mem[1442] : 
                       (N717)? mem[1458] : 
                       (N719)? mem[1474] : 
                       (N721)? mem[1490] : 
                       (N723)? mem[1506] : 
                       (N725)? mem[1522] : 
                       (N727)? mem[1538] : 
                       (N729)? mem[1554] : 
                       (N731)? mem[1570] : 
                       (N733)? mem[1586] : 
                       (N735)? mem[1602] : 
                       (N737)? mem[1618] : 
                       (N739)? mem[1634] : 
                       (N741)? mem[1650] : 
                       (N743)? mem[1666] : 
                       (N745)? mem[1682] : 
                       (N747)? mem[1698] : 
                       (N749)? mem[1714] : 
                       (N751)? mem[1730] : 
                       (N753)? mem[1746] : 
                       (N755)? mem[1762] : 
                       (N757)? mem[1778] : 
                       (N759)? mem[1794] : 
                       (N761)? mem[1810] : 
                       (N763)? mem[1826] : 
                       (N765)? mem[1842] : 
                       (N767)? mem[1858] : 
                       (N769)? mem[1874] : 
                       (N771)? mem[1890] : 
                       (N773)? mem[1906] : 
                       (N775)? mem[1922] : 
                       (N777)? mem[1938] : 
                       (N779)? mem[1954] : 
                       (N781)? mem[1970] : 
                       (N783)? mem[1986] : 
                       (N785)? mem[2002] : 
                       (N787)? mem[2018] : 
                       (N789)? mem[2034] : 
                       (N791)? mem[2050] : 
                       (N793)? mem[2066] : 
                       (N795)? mem[2082] : 
                       (N797)? mem[2098] : 
                       (N799)? mem[2114] : 
                       (N801)? mem[2130] : 
                       (N803)? mem[2146] : 
                       (N805)? mem[2162] : 
                       (N807)? mem[2178] : 
                       (N809)? mem[2194] : 
                       (N811)? mem[2210] : 
                       (N813)? mem[2226] : 
                       (N815)? mem[2242] : 
                       (N817)? mem[2258] : 
                       (N819)? mem[2274] : 
                       (N821)? mem[2290] : 
                       (N823)? mem[2306] : 
                       (N825)? mem[2322] : 
                       (N827)? mem[2338] : 
                       (N829)? mem[2354] : 
                       (N831)? mem[2370] : 
                       (N833)? mem[2386] : 
                       (N835)? mem[2402] : 
                       (N837)? mem[2418] : 
                       (N839)? mem[2434] : 
                       (N841)? mem[2450] : 
                       (N843)? mem[2466] : 
                       (N845)? mem[2482] : 
                       (N847)? mem[2498] : 
                       (N849)? mem[2514] : 
                       (N851)? mem[2530] : 
                       (N853)? mem[2546] : 
                       (N855)? mem[2562] : 
                       (N857)? mem[2578] : 
                       (N859)? mem[2594] : 
                       (N861)? mem[2610] : 
                       (N863)? mem[2626] : 
                       (N865)? mem[2642] : 
                       (N867)? mem[2658] : 
                       (N869)? mem[2674] : 
                       (N871)? mem[2690] : 
                       (N873)? mem[2706] : 
                       (N875)? mem[2722] : 
                       (N877)? mem[2738] : 
                       (N879)? mem[2754] : 
                       (N881)? mem[2770] : 
                       (N883)? mem[2786] : 
                       (N885)? mem[2802] : 
                       (N887)? mem[2818] : 
                       (N889)? mem[2834] : 
                       (N891)? mem[2850] : 
                       (N893)? mem[2866] : 
                       (N895)? mem[2882] : 
                       (N897)? mem[2898] : 
                       (N899)? mem[2914] : 
                       (N901)? mem[2930] : 
                       (N903)? mem[2946] : 
                       (N905)? mem[2962] : 
                       (N907)? mem[2978] : 
                       (N909)? mem[2994] : 
                       (N911)? mem[3010] : 
                       (N913)? mem[3026] : 
                       (N915)? mem[3042] : 
                       (N917)? mem[3058] : 
                       (N919)? mem[3074] : 
                       (N921)? mem[3090] : 
                       (N923)? mem[3106] : 
                       (N925)? mem[3122] : 
                       (N927)? mem[3138] : 
                       (N929)? mem[3154] : 
                       (N931)? mem[3170] : 
                       (N933)? mem[3186] : 
                       (N935)? mem[3202] : 
                       (N937)? mem[3218] : 
                       (N939)? mem[3234] : 
                       (N941)? mem[3250] : 
                       (N943)? mem[3266] : 
                       (N945)? mem[3282] : 
                       (N947)? mem[3298] : 
                       (N949)? mem[3314] : 
                       (N951)? mem[3330] : 
                       (N953)? mem[3346] : 
                       (N955)? mem[3362] : 
                       (N957)? mem[3378] : 
                       (N959)? mem[3394] : 
                       (N961)? mem[3410] : 
                       (N963)? mem[3426] : 
                       (N965)? mem[3442] : 
                       (N967)? mem[3458] : 
                       (N969)? mem[3474] : 
                       (N971)? mem[3490] : 
                       (N973)? mem[3506] : 
                       (N975)? mem[3522] : 
                       (N977)? mem[3538] : 
                       (N979)? mem[3554] : 
                       (N981)? mem[3570] : 
                       (N983)? mem[3586] : 
                       (N985)? mem[3602] : 
                       (N987)? mem[3618] : 
                       (N989)? mem[3634] : 
                       (N991)? mem[3650] : 
                       (N993)? mem[3666] : 
                       (N995)? mem[3682] : 
                       (N997)? mem[3698] : 
                       (N999)? mem[3714] : 
                       (N1001)? mem[3730] : 
                       (N1003)? mem[3746] : 
                       (N1005)? mem[3762] : 
                       (N1007)? mem[3778] : 
                       (N1009)? mem[3794] : 
                       (N1011)? mem[3810] : 
                       (N1013)? mem[3826] : 
                       (N1015)? mem[3842] : 
                       (N1017)? mem[3858] : 
                       (N1019)? mem[3874] : 
                       (N1021)? mem[3890] : 
                       (N1023)? mem[3906] : 
                       (N1025)? mem[3922] : 
                       (N1027)? mem[3938] : 
                       (N1029)? mem[3954] : 
                       (N1031)? mem[3970] : 
                       (N1033)? mem[3986] : 
                       (N1035)? mem[4002] : 
                       (N1037)? mem[4018] : 
                       (N1039)? mem[4034] : 
                       (N1041)? mem[4050] : 
                       (N1043)? mem[4066] : 
                       (N1045)? mem[4082] : 
                       (N536)? mem[4098] : 
                       (N538)? mem[4114] : 
                       (N540)? mem[4130] : 
                       (N542)? mem[4146] : 
                       (N544)? mem[4162] : 
                       (N546)? mem[4178] : 
                       (N548)? mem[4194] : 
                       (N550)? mem[4210] : 
                       (N552)? mem[4226] : 
                       (N554)? mem[4242] : 
                       (N556)? mem[4258] : 
                       (N558)? mem[4274] : 
                       (N560)? mem[4290] : 
                       (N562)? mem[4306] : 
                       (N564)? mem[4322] : 
                       (N566)? mem[4338] : 
                       (N568)? mem[4354] : 
                       (N570)? mem[4370] : 
                       (N572)? mem[4386] : 
                       (N574)? mem[4402] : 
                       (N576)? mem[4418] : 
                       (N578)? mem[4434] : 
                       (N580)? mem[4450] : 
                       (N582)? mem[4466] : 
                       (N584)? mem[4482] : 
                       (N586)? mem[4498] : 
                       (N588)? mem[4514] : 
                       (N590)? mem[4530] : 
                       (N592)? mem[4546] : 
                       (N594)? mem[4562] : 
                       (N596)? mem[4578] : 
                       (N598)? mem[4594] : 
                       (N600)? mem[4610] : 
                       (N602)? mem[4626] : 
                       (N604)? mem[4642] : 
                       (N606)? mem[4658] : 
                       (N608)? mem[4674] : 
                       (N610)? mem[4690] : 
                       (N612)? mem[4706] : 
                       (N614)? mem[4722] : 
                       (N616)? mem[4738] : 
                       (N618)? mem[4754] : 
                       (N620)? mem[4770] : 
                       (N622)? mem[4786] : 
                       (N624)? mem[4802] : 
                       (N626)? mem[4818] : 
                       (N628)? mem[4834] : 
                       (N630)? mem[4850] : 
                       (N632)? mem[4866] : 
                       (N634)? mem[4882] : 
                       (N636)? mem[4898] : 
                       (N638)? mem[4914] : 
                       (N640)? mem[4930] : 
                       (N642)? mem[4946] : 
                       (N644)? mem[4962] : 
                       (N646)? mem[4978] : 
                       (N648)? mem[4994] : 
                       (N650)? mem[5010] : 
                       (N652)? mem[5026] : 
                       (N654)? mem[5042] : 
                       (N656)? mem[5058] : 
                       (N658)? mem[5074] : 
                       (N660)? mem[5090] : 
                       (N662)? mem[5106] : 
                       (N664)? mem[5122] : 
                       (N666)? mem[5138] : 
                       (N668)? mem[5154] : 
                       (N670)? mem[5170] : 
                       (N672)? mem[5186] : 
                       (N674)? mem[5202] : 
                       (N676)? mem[5218] : 
                       (N678)? mem[5234] : 
                       (N680)? mem[5250] : 
                       (N682)? mem[5266] : 
                       (N684)? mem[5282] : 
                       (N686)? mem[5298] : 
                       (N688)? mem[5314] : 
                       (N690)? mem[5330] : 
                       (N692)? mem[5346] : 
                       (N694)? mem[5362] : 
                       (N696)? mem[5378] : 
                       (N698)? mem[5394] : 
                       (N700)? mem[5410] : 
                       (N702)? mem[5426] : 
                       (N704)? mem[5442] : 
                       (N706)? mem[5458] : 
                       (N708)? mem[5474] : 
                       (N710)? mem[5490] : 
                       (N712)? mem[5506] : 
                       (N714)? mem[5522] : 
                       (N716)? mem[5538] : 
                       (N718)? mem[5554] : 
                       (N720)? mem[5570] : 
                       (N722)? mem[5586] : 
                       (N724)? mem[5602] : 
                       (N726)? mem[5618] : 
                       (N728)? mem[5634] : 
                       (N730)? mem[5650] : 
                       (N732)? mem[5666] : 
                       (N734)? mem[5682] : 
                       (N736)? mem[5698] : 
                       (N738)? mem[5714] : 
                       (N740)? mem[5730] : 
                       (N742)? mem[5746] : 
                       (N744)? mem[5762] : 
                       (N746)? mem[5778] : 
                       (N748)? mem[5794] : 
                       (N750)? mem[5810] : 
                       (N752)? mem[5826] : 
                       (N754)? mem[5842] : 
                       (N756)? mem[5858] : 
                       (N758)? mem[5874] : 
                       (N760)? mem[5890] : 
                       (N762)? mem[5906] : 
                       (N764)? mem[5922] : 
                       (N766)? mem[5938] : 
                       (N768)? mem[5954] : 
                       (N770)? mem[5970] : 
                       (N772)? mem[5986] : 
                       (N774)? mem[6002] : 
                       (N776)? mem[6018] : 
                       (N778)? mem[6034] : 
                       (N780)? mem[6050] : 
                       (N782)? mem[6066] : 
                       (N784)? mem[6082] : 
                       (N786)? mem[6098] : 
                       (N788)? mem[6114] : 
                       (N790)? mem[6130] : 
                       (N792)? mem[6146] : 
                       (N794)? mem[6162] : 
                       (N796)? mem[6178] : 
                       (N798)? mem[6194] : 
                       (N800)? mem[6210] : 
                       (N802)? mem[6226] : 
                       (N804)? mem[6242] : 
                       (N806)? mem[6258] : 
                       (N808)? mem[6274] : 
                       (N810)? mem[6290] : 
                       (N812)? mem[6306] : 
                       (N814)? mem[6322] : 
                       (N816)? mem[6338] : 
                       (N818)? mem[6354] : 
                       (N820)? mem[6370] : 
                       (N822)? mem[6386] : 
                       (N824)? mem[6402] : 
                       (N826)? mem[6418] : 
                       (N828)? mem[6434] : 
                       (N830)? mem[6450] : 
                       (N832)? mem[6466] : 
                       (N834)? mem[6482] : 
                       (N836)? mem[6498] : 
                       (N838)? mem[6514] : 
                       (N840)? mem[6530] : 
                       (N842)? mem[6546] : 
                       (N844)? mem[6562] : 
                       (N846)? mem[6578] : 
                       (N848)? mem[6594] : 
                       (N850)? mem[6610] : 
                       (N852)? mem[6626] : 
                       (N854)? mem[6642] : 
                       (N856)? mem[6658] : 
                       (N858)? mem[6674] : 
                       (N860)? mem[6690] : 
                       (N862)? mem[6706] : 
                       (N864)? mem[6722] : 
                       (N866)? mem[6738] : 
                       (N868)? mem[6754] : 
                       (N870)? mem[6770] : 
                       (N872)? mem[6786] : 
                       (N874)? mem[6802] : 
                       (N876)? mem[6818] : 
                       (N878)? mem[6834] : 
                       (N880)? mem[6850] : 
                       (N882)? mem[6866] : 
                       (N884)? mem[6882] : 
                       (N886)? mem[6898] : 
                       (N888)? mem[6914] : 
                       (N890)? mem[6930] : 
                       (N892)? mem[6946] : 
                       (N894)? mem[6962] : 
                       (N896)? mem[6978] : 
                       (N898)? mem[6994] : 
                       (N900)? mem[7010] : 
                       (N902)? mem[7026] : 
                       (N904)? mem[7042] : 
                       (N906)? mem[7058] : 
                       (N908)? mem[7074] : 
                       (N910)? mem[7090] : 
                       (N912)? mem[7106] : 
                       (N914)? mem[7122] : 
                       (N916)? mem[7138] : 
                       (N918)? mem[7154] : 
                       (N920)? mem[7170] : 
                       (N922)? mem[7186] : 
                       (N924)? mem[7202] : 
                       (N926)? mem[7218] : 
                       (N928)? mem[7234] : 
                       (N930)? mem[7250] : 
                       (N932)? mem[7266] : 
                       (N934)? mem[7282] : 
                       (N936)? mem[7298] : 
                       (N938)? mem[7314] : 
                       (N940)? mem[7330] : 
                       (N942)? mem[7346] : 
                       (N944)? mem[7362] : 
                       (N946)? mem[7378] : 
                       (N948)? mem[7394] : 
                       (N950)? mem[7410] : 
                       (N952)? mem[7426] : 
                       (N954)? mem[7442] : 
                       (N956)? mem[7458] : 
                       (N958)? mem[7474] : 
                       (N960)? mem[7490] : 
                       (N962)? mem[7506] : 
                       (N964)? mem[7522] : 
                       (N966)? mem[7538] : 
                       (N968)? mem[7554] : 
                       (N970)? mem[7570] : 
                       (N972)? mem[7586] : 
                       (N974)? mem[7602] : 
                       (N976)? mem[7618] : 
                       (N978)? mem[7634] : 
                       (N980)? mem[7650] : 
                       (N982)? mem[7666] : 
                       (N984)? mem[7682] : 
                       (N986)? mem[7698] : 
                       (N988)? mem[7714] : 
                       (N990)? mem[7730] : 
                       (N992)? mem[7746] : 
                       (N994)? mem[7762] : 
                       (N996)? mem[7778] : 
                       (N998)? mem[7794] : 
                       (N1000)? mem[7810] : 
                       (N1002)? mem[7826] : 
                       (N1004)? mem[7842] : 
                       (N1006)? mem[7858] : 
                       (N1008)? mem[7874] : 
                       (N1010)? mem[7890] : 
                       (N1012)? mem[7906] : 
                       (N1014)? mem[7922] : 
                       (N1016)? mem[7938] : 
                       (N1018)? mem[7954] : 
                       (N1020)? mem[7970] : 
                       (N1022)? mem[7986] : 
                       (N1024)? mem[8002] : 
                       (N1026)? mem[8018] : 
                       (N1028)? mem[8034] : 
                       (N1030)? mem[8050] : 
                       (N1032)? mem[8066] : 
                       (N1034)? mem[8082] : 
                       (N1036)? mem[8098] : 
                       (N1038)? mem[8114] : 
                       (N1040)? mem[8130] : 
                       (N1042)? mem[8146] : 
                       (N1044)? mem[8162] : 
                       (N1046)? mem[8178] : 1'b0;
  assign r_data_o[1] = (N535)? mem[1] : 
                       (N537)? mem[17] : 
                       (N539)? mem[33] : 
                       (N541)? mem[49] : 
                       (N543)? mem[65] : 
                       (N545)? mem[81] : 
                       (N547)? mem[97] : 
                       (N549)? mem[113] : 
                       (N551)? mem[129] : 
                       (N553)? mem[145] : 
                       (N555)? mem[161] : 
                       (N557)? mem[177] : 
                       (N559)? mem[193] : 
                       (N561)? mem[209] : 
                       (N563)? mem[225] : 
                       (N565)? mem[241] : 
                       (N567)? mem[257] : 
                       (N569)? mem[273] : 
                       (N571)? mem[289] : 
                       (N573)? mem[305] : 
                       (N575)? mem[321] : 
                       (N577)? mem[337] : 
                       (N579)? mem[353] : 
                       (N581)? mem[369] : 
                       (N583)? mem[385] : 
                       (N585)? mem[401] : 
                       (N587)? mem[417] : 
                       (N589)? mem[433] : 
                       (N591)? mem[449] : 
                       (N593)? mem[465] : 
                       (N595)? mem[481] : 
                       (N597)? mem[497] : 
                       (N599)? mem[513] : 
                       (N601)? mem[529] : 
                       (N603)? mem[545] : 
                       (N605)? mem[561] : 
                       (N607)? mem[577] : 
                       (N609)? mem[593] : 
                       (N611)? mem[609] : 
                       (N613)? mem[625] : 
                       (N615)? mem[641] : 
                       (N617)? mem[657] : 
                       (N619)? mem[673] : 
                       (N621)? mem[689] : 
                       (N623)? mem[705] : 
                       (N625)? mem[721] : 
                       (N627)? mem[737] : 
                       (N629)? mem[753] : 
                       (N631)? mem[769] : 
                       (N633)? mem[785] : 
                       (N635)? mem[801] : 
                       (N637)? mem[817] : 
                       (N639)? mem[833] : 
                       (N641)? mem[849] : 
                       (N643)? mem[865] : 
                       (N645)? mem[881] : 
                       (N647)? mem[897] : 
                       (N649)? mem[913] : 
                       (N651)? mem[929] : 
                       (N653)? mem[945] : 
                       (N655)? mem[961] : 
                       (N657)? mem[977] : 
                       (N659)? mem[993] : 
                       (N661)? mem[1009] : 
                       (N663)? mem[1025] : 
                       (N665)? mem[1041] : 
                       (N667)? mem[1057] : 
                       (N669)? mem[1073] : 
                       (N671)? mem[1089] : 
                       (N673)? mem[1105] : 
                       (N675)? mem[1121] : 
                       (N677)? mem[1137] : 
                       (N679)? mem[1153] : 
                       (N681)? mem[1169] : 
                       (N683)? mem[1185] : 
                       (N685)? mem[1201] : 
                       (N687)? mem[1217] : 
                       (N689)? mem[1233] : 
                       (N691)? mem[1249] : 
                       (N693)? mem[1265] : 
                       (N695)? mem[1281] : 
                       (N697)? mem[1297] : 
                       (N699)? mem[1313] : 
                       (N701)? mem[1329] : 
                       (N703)? mem[1345] : 
                       (N705)? mem[1361] : 
                       (N707)? mem[1377] : 
                       (N709)? mem[1393] : 
                       (N711)? mem[1409] : 
                       (N713)? mem[1425] : 
                       (N715)? mem[1441] : 
                       (N717)? mem[1457] : 
                       (N719)? mem[1473] : 
                       (N721)? mem[1489] : 
                       (N723)? mem[1505] : 
                       (N725)? mem[1521] : 
                       (N727)? mem[1537] : 
                       (N729)? mem[1553] : 
                       (N731)? mem[1569] : 
                       (N733)? mem[1585] : 
                       (N735)? mem[1601] : 
                       (N737)? mem[1617] : 
                       (N739)? mem[1633] : 
                       (N741)? mem[1649] : 
                       (N743)? mem[1665] : 
                       (N745)? mem[1681] : 
                       (N747)? mem[1697] : 
                       (N749)? mem[1713] : 
                       (N751)? mem[1729] : 
                       (N753)? mem[1745] : 
                       (N755)? mem[1761] : 
                       (N757)? mem[1777] : 
                       (N759)? mem[1793] : 
                       (N761)? mem[1809] : 
                       (N763)? mem[1825] : 
                       (N765)? mem[1841] : 
                       (N767)? mem[1857] : 
                       (N769)? mem[1873] : 
                       (N771)? mem[1889] : 
                       (N773)? mem[1905] : 
                       (N775)? mem[1921] : 
                       (N777)? mem[1937] : 
                       (N779)? mem[1953] : 
                       (N781)? mem[1969] : 
                       (N783)? mem[1985] : 
                       (N785)? mem[2001] : 
                       (N787)? mem[2017] : 
                       (N789)? mem[2033] : 
                       (N791)? mem[2049] : 
                       (N793)? mem[2065] : 
                       (N795)? mem[2081] : 
                       (N797)? mem[2097] : 
                       (N799)? mem[2113] : 
                       (N801)? mem[2129] : 
                       (N803)? mem[2145] : 
                       (N805)? mem[2161] : 
                       (N807)? mem[2177] : 
                       (N809)? mem[2193] : 
                       (N811)? mem[2209] : 
                       (N813)? mem[2225] : 
                       (N815)? mem[2241] : 
                       (N817)? mem[2257] : 
                       (N819)? mem[2273] : 
                       (N821)? mem[2289] : 
                       (N823)? mem[2305] : 
                       (N825)? mem[2321] : 
                       (N827)? mem[2337] : 
                       (N829)? mem[2353] : 
                       (N831)? mem[2369] : 
                       (N833)? mem[2385] : 
                       (N835)? mem[2401] : 
                       (N837)? mem[2417] : 
                       (N839)? mem[2433] : 
                       (N841)? mem[2449] : 
                       (N843)? mem[2465] : 
                       (N845)? mem[2481] : 
                       (N847)? mem[2497] : 
                       (N849)? mem[2513] : 
                       (N851)? mem[2529] : 
                       (N853)? mem[2545] : 
                       (N855)? mem[2561] : 
                       (N857)? mem[2577] : 
                       (N859)? mem[2593] : 
                       (N861)? mem[2609] : 
                       (N863)? mem[2625] : 
                       (N865)? mem[2641] : 
                       (N867)? mem[2657] : 
                       (N869)? mem[2673] : 
                       (N871)? mem[2689] : 
                       (N873)? mem[2705] : 
                       (N875)? mem[2721] : 
                       (N877)? mem[2737] : 
                       (N879)? mem[2753] : 
                       (N881)? mem[2769] : 
                       (N883)? mem[2785] : 
                       (N885)? mem[2801] : 
                       (N887)? mem[2817] : 
                       (N889)? mem[2833] : 
                       (N891)? mem[2849] : 
                       (N893)? mem[2865] : 
                       (N895)? mem[2881] : 
                       (N897)? mem[2897] : 
                       (N899)? mem[2913] : 
                       (N901)? mem[2929] : 
                       (N903)? mem[2945] : 
                       (N905)? mem[2961] : 
                       (N907)? mem[2977] : 
                       (N909)? mem[2993] : 
                       (N911)? mem[3009] : 
                       (N913)? mem[3025] : 
                       (N915)? mem[3041] : 
                       (N917)? mem[3057] : 
                       (N919)? mem[3073] : 
                       (N921)? mem[3089] : 
                       (N923)? mem[3105] : 
                       (N925)? mem[3121] : 
                       (N927)? mem[3137] : 
                       (N929)? mem[3153] : 
                       (N931)? mem[3169] : 
                       (N933)? mem[3185] : 
                       (N935)? mem[3201] : 
                       (N937)? mem[3217] : 
                       (N939)? mem[3233] : 
                       (N941)? mem[3249] : 
                       (N943)? mem[3265] : 
                       (N945)? mem[3281] : 
                       (N947)? mem[3297] : 
                       (N949)? mem[3313] : 
                       (N951)? mem[3329] : 
                       (N953)? mem[3345] : 
                       (N955)? mem[3361] : 
                       (N957)? mem[3377] : 
                       (N959)? mem[3393] : 
                       (N961)? mem[3409] : 
                       (N963)? mem[3425] : 
                       (N965)? mem[3441] : 
                       (N967)? mem[3457] : 
                       (N969)? mem[3473] : 
                       (N971)? mem[3489] : 
                       (N973)? mem[3505] : 
                       (N975)? mem[3521] : 
                       (N977)? mem[3537] : 
                       (N979)? mem[3553] : 
                       (N981)? mem[3569] : 
                       (N983)? mem[3585] : 
                       (N985)? mem[3601] : 
                       (N987)? mem[3617] : 
                       (N989)? mem[3633] : 
                       (N991)? mem[3649] : 
                       (N993)? mem[3665] : 
                       (N995)? mem[3681] : 
                       (N997)? mem[3697] : 
                       (N999)? mem[3713] : 
                       (N1001)? mem[3729] : 
                       (N1003)? mem[3745] : 
                       (N1005)? mem[3761] : 
                       (N1007)? mem[3777] : 
                       (N1009)? mem[3793] : 
                       (N1011)? mem[3809] : 
                       (N1013)? mem[3825] : 
                       (N1015)? mem[3841] : 
                       (N1017)? mem[3857] : 
                       (N1019)? mem[3873] : 
                       (N1021)? mem[3889] : 
                       (N1023)? mem[3905] : 
                       (N1025)? mem[3921] : 
                       (N1027)? mem[3937] : 
                       (N1029)? mem[3953] : 
                       (N1031)? mem[3969] : 
                       (N1033)? mem[3985] : 
                       (N1035)? mem[4001] : 
                       (N1037)? mem[4017] : 
                       (N1039)? mem[4033] : 
                       (N1041)? mem[4049] : 
                       (N1043)? mem[4065] : 
                       (N1045)? mem[4081] : 
                       (N536)? mem[4097] : 
                       (N538)? mem[4113] : 
                       (N540)? mem[4129] : 
                       (N542)? mem[4145] : 
                       (N544)? mem[4161] : 
                       (N546)? mem[4177] : 
                       (N548)? mem[4193] : 
                       (N550)? mem[4209] : 
                       (N552)? mem[4225] : 
                       (N554)? mem[4241] : 
                       (N556)? mem[4257] : 
                       (N558)? mem[4273] : 
                       (N560)? mem[4289] : 
                       (N562)? mem[4305] : 
                       (N564)? mem[4321] : 
                       (N566)? mem[4337] : 
                       (N568)? mem[4353] : 
                       (N570)? mem[4369] : 
                       (N572)? mem[4385] : 
                       (N574)? mem[4401] : 
                       (N576)? mem[4417] : 
                       (N578)? mem[4433] : 
                       (N580)? mem[4449] : 
                       (N582)? mem[4465] : 
                       (N584)? mem[4481] : 
                       (N586)? mem[4497] : 
                       (N588)? mem[4513] : 
                       (N590)? mem[4529] : 
                       (N592)? mem[4545] : 
                       (N594)? mem[4561] : 
                       (N596)? mem[4577] : 
                       (N598)? mem[4593] : 
                       (N600)? mem[4609] : 
                       (N602)? mem[4625] : 
                       (N604)? mem[4641] : 
                       (N606)? mem[4657] : 
                       (N608)? mem[4673] : 
                       (N610)? mem[4689] : 
                       (N612)? mem[4705] : 
                       (N614)? mem[4721] : 
                       (N616)? mem[4737] : 
                       (N618)? mem[4753] : 
                       (N620)? mem[4769] : 
                       (N622)? mem[4785] : 
                       (N624)? mem[4801] : 
                       (N626)? mem[4817] : 
                       (N628)? mem[4833] : 
                       (N630)? mem[4849] : 
                       (N632)? mem[4865] : 
                       (N634)? mem[4881] : 
                       (N636)? mem[4897] : 
                       (N638)? mem[4913] : 
                       (N640)? mem[4929] : 
                       (N642)? mem[4945] : 
                       (N644)? mem[4961] : 
                       (N646)? mem[4977] : 
                       (N648)? mem[4993] : 
                       (N650)? mem[5009] : 
                       (N652)? mem[5025] : 
                       (N654)? mem[5041] : 
                       (N656)? mem[5057] : 
                       (N658)? mem[5073] : 
                       (N660)? mem[5089] : 
                       (N662)? mem[5105] : 
                       (N664)? mem[5121] : 
                       (N666)? mem[5137] : 
                       (N668)? mem[5153] : 
                       (N670)? mem[5169] : 
                       (N672)? mem[5185] : 
                       (N674)? mem[5201] : 
                       (N676)? mem[5217] : 
                       (N678)? mem[5233] : 
                       (N680)? mem[5249] : 
                       (N682)? mem[5265] : 
                       (N684)? mem[5281] : 
                       (N686)? mem[5297] : 
                       (N688)? mem[5313] : 
                       (N690)? mem[5329] : 
                       (N692)? mem[5345] : 
                       (N694)? mem[5361] : 
                       (N696)? mem[5377] : 
                       (N698)? mem[5393] : 
                       (N700)? mem[5409] : 
                       (N702)? mem[5425] : 
                       (N704)? mem[5441] : 
                       (N706)? mem[5457] : 
                       (N708)? mem[5473] : 
                       (N710)? mem[5489] : 
                       (N712)? mem[5505] : 
                       (N714)? mem[5521] : 
                       (N716)? mem[5537] : 
                       (N718)? mem[5553] : 
                       (N720)? mem[5569] : 
                       (N722)? mem[5585] : 
                       (N724)? mem[5601] : 
                       (N726)? mem[5617] : 
                       (N728)? mem[5633] : 
                       (N730)? mem[5649] : 
                       (N732)? mem[5665] : 
                       (N734)? mem[5681] : 
                       (N736)? mem[5697] : 
                       (N738)? mem[5713] : 
                       (N740)? mem[5729] : 
                       (N742)? mem[5745] : 
                       (N744)? mem[5761] : 
                       (N746)? mem[5777] : 
                       (N748)? mem[5793] : 
                       (N750)? mem[5809] : 
                       (N752)? mem[5825] : 
                       (N754)? mem[5841] : 
                       (N756)? mem[5857] : 
                       (N758)? mem[5873] : 
                       (N760)? mem[5889] : 
                       (N762)? mem[5905] : 
                       (N764)? mem[5921] : 
                       (N766)? mem[5937] : 
                       (N768)? mem[5953] : 
                       (N770)? mem[5969] : 
                       (N772)? mem[5985] : 
                       (N774)? mem[6001] : 
                       (N776)? mem[6017] : 
                       (N778)? mem[6033] : 
                       (N780)? mem[6049] : 
                       (N782)? mem[6065] : 
                       (N784)? mem[6081] : 
                       (N786)? mem[6097] : 
                       (N788)? mem[6113] : 
                       (N790)? mem[6129] : 
                       (N792)? mem[6145] : 
                       (N794)? mem[6161] : 
                       (N796)? mem[6177] : 
                       (N798)? mem[6193] : 
                       (N800)? mem[6209] : 
                       (N802)? mem[6225] : 
                       (N804)? mem[6241] : 
                       (N806)? mem[6257] : 
                       (N808)? mem[6273] : 
                       (N810)? mem[6289] : 
                       (N812)? mem[6305] : 
                       (N814)? mem[6321] : 
                       (N816)? mem[6337] : 
                       (N818)? mem[6353] : 
                       (N820)? mem[6369] : 
                       (N822)? mem[6385] : 
                       (N824)? mem[6401] : 
                       (N826)? mem[6417] : 
                       (N828)? mem[6433] : 
                       (N830)? mem[6449] : 
                       (N832)? mem[6465] : 
                       (N834)? mem[6481] : 
                       (N836)? mem[6497] : 
                       (N838)? mem[6513] : 
                       (N840)? mem[6529] : 
                       (N842)? mem[6545] : 
                       (N844)? mem[6561] : 
                       (N846)? mem[6577] : 
                       (N848)? mem[6593] : 
                       (N850)? mem[6609] : 
                       (N852)? mem[6625] : 
                       (N854)? mem[6641] : 
                       (N856)? mem[6657] : 
                       (N858)? mem[6673] : 
                       (N860)? mem[6689] : 
                       (N862)? mem[6705] : 
                       (N864)? mem[6721] : 
                       (N866)? mem[6737] : 
                       (N868)? mem[6753] : 
                       (N870)? mem[6769] : 
                       (N872)? mem[6785] : 
                       (N874)? mem[6801] : 
                       (N876)? mem[6817] : 
                       (N878)? mem[6833] : 
                       (N880)? mem[6849] : 
                       (N882)? mem[6865] : 
                       (N884)? mem[6881] : 
                       (N886)? mem[6897] : 
                       (N888)? mem[6913] : 
                       (N890)? mem[6929] : 
                       (N892)? mem[6945] : 
                       (N894)? mem[6961] : 
                       (N896)? mem[6977] : 
                       (N898)? mem[6993] : 
                       (N900)? mem[7009] : 
                       (N902)? mem[7025] : 
                       (N904)? mem[7041] : 
                       (N906)? mem[7057] : 
                       (N908)? mem[7073] : 
                       (N910)? mem[7089] : 
                       (N912)? mem[7105] : 
                       (N914)? mem[7121] : 
                       (N916)? mem[7137] : 
                       (N918)? mem[7153] : 
                       (N920)? mem[7169] : 
                       (N922)? mem[7185] : 
                       (N924)? mem[7201] : 
                       (N926)? mem[7217] : 
                       (N928)? mem[7233] : 
                       (N930)? mem[7249] : 
                       (N932)? mem[7265] : 
                       (N934)? mem[7281] : 
                       (N936)? mem[7297] : 
                       (N938)? mem[7313] : 
                       (N940)? mem[7329] : 
                       (N942)? mem[7345] : 
                       (N944)? mem[7361] : 
                       (N946)? mem[7377] : 
                       (N948)? mem[7393] : 
                       (N950)? mem[7409] : 
                       (N952)? mem[7425] : 
                       (N954)? mem[7441] : 
                       (N956)? mem[7457] : 
                       (N958)? mem[7473] : 
                       (N960)? mem[7489] : 
                       (N962)? mem[7505] : 
                       (N964)? mem[7521] : 
                       (N966)? mem[7537] : 
                       (N968)? mem[7553] : 
                       (N970)? mem[7569] : 
                       (N972)? mem[7585] : 
                       (N974)? mem[7601] : 
                       (N976)? mem[7617] : 
                       (N978)? mem[7633] : 
                       (N980)? mem[7649] : 
                       (N982)? mem[7665] : 
                       (N984)? mem[7681] : 
                       (N986)? mem[7697] : 
                       (N988)? mem[7713] : 
                       (N990)? mem[7729] : 
                       (N992)? mem[7745] : 
                       (N994)? mem[7761] : 
                       (N996)? mem[7777] : 
                       (N998)? mem[7793] : 
                       (N1000)? mem[7809] : 
                       (N1002)? mem[7825] : 
                       (N1004)? mem[7841] : 
                       (N1006)? mem[7857] : 
                       (N1008)? mem[7873] : 
                       (N1010)? mem[7889] : 
                       (N1012)? mem[7905] : 
                       (N1014)? mem[7921] : 
                       (N1016)? mem[7937] : 
                       (N1018)? mem[7953] : 
                       (N1020)? mem[7969] : 
                       (N1022)? mem[7985] : 
                       (N1024)? mem[8001] : 
                       (N1026)? mem[8017] : 
                       (N1028)? mem[8033] : 
                       (N1030)? mem[8049] : 
                       (N1032)? mem[8065] : 
                       (N1034)? mem[8081] : 
                       (N1036)? mem[8097] : 
                       (N1038)? mem[8113] : 
                       (N1040)? mem[8129] : 
                       (N1042)? mem[8145] : 
                       (N1044)? mem[8161] : 
                       (N1046)? mem[8177] : 1'b0;
  assign r_data_o[0] = (N535)? mem[0] : 
                       (N537)? mem[16] : 
                       (N539)? mem[32] : 
                       (N541)? mem[48] : 
                       (N543)? mem[64] : 
                       (N545)? mem[80] : 
                       (N547)? mem[96] : 
                       (N549)? mem[112] : 
                       (N551)? mem[128] : 
                       (N553)? mem[144] : 
                       (N555)? mem[160] : 
                       (N557)? mem[176] : 
                       (N559)? mem[192] : 
                       (N561)? mem[208] : 
                       (N563)? mem[224] : 
                       (N565)? mem[240] : 
                       (N567)? mem[256] : 
                       (N569)? mem[272] : 
                       (N571)? mem[288] : 
                       (N573)? mem[304] : 
                       (N575)? mem[320] : 
                       (N577)? mem[336] : 
                       (N579)? mem[352] : 
                       (N581)? mem[368] : 
                       (N583)? mem[384] : 
                       (N585)? mem[400] : 
                       (N587)? mem[416] : 
                       (N589)? mem[432] : 
                       (N591)? mem[448] : 
                       (N593)? mem[464] : 
                       (N595)? mem[480] : 
                       (N597)? mem[496] : 
                       (N599)? mem[512] : 
                       (N601)? mem[528] : 
                       (N603)? mem[544] : 
                       (N605)? mem[560] : 
                       (N607)? mem[576] : 
                       (N609)? mem[592] : 
                       (N611)? mem[608] : 
                       (N613)? mem[624] : 
                       (N615)? mem[640] : 
                       (N617)? mem[656] : 
                       (N619)? mem[672] : 
                       (N621)? mem[688] : 
                       (N623)? mem[704] : 
                       (N625)? mem[720] : 
                       (N627)? mem[736] : 
                       (N629)? mem[752] : 
                       (N631)? mem[768] : 
                       (N633)? mem[784] : 
                       (N635)? mem[800] : 
                       (N637)? mem[816] : 
                       (N639)? mem[832] : 
                       (N641)? mem[848] : 
                       (N643)? mem[864] : 
                       (N645)? mem[880] : 
                       (N647)? mem[896] : 
                       (N649)? mem[912] : 
                       (N651)? mem[928] : 
                       (N653)? mem[944] : 
                       (N655)? mem[960] : 
                       (N657)? mem[976] : 
                       (N659)? mem[992] : 
                       (N661)? mem[1008] : 
                       (N663)? mem[1024] : 
                       (N665)? mem[1040] : 
                       (N667)? mem[1056] : 
                       (N669)? mem[1072] : 
                       (N671)? mem[1088] : 
                       (N673)? mem[1104] : 
                       (N675)? mem[1120] : 
                       (N677)? mem[1136] : 
                       (N679)? mem[1152] : 
                       (N681)? mem[1168] : 
                       (N683)? mem[1184] : 
                       (N685)? mem[1200] : 
                       (N687)? mem[1216] : 
                       (N689)? mem[1232] : 
                       (N691)? mem[1248] : 
                       (N693)? mem[1264] : 
                       (N695)? mem[1280] : 
                       (N697)? mem[1296] : 
                       (N699)? mem[1312] : 
                       (N701)? mem[1328] : 
                       (N703)? mem[1344] : 
                       (N705)? mem[1360] : 
                       (N707)? mem[1376] : 
                       (N709)? mem[1392] : 
                       (N711)? mem[1408] : 
                       (N713)? mem[1424] : 
                       (N715)? mem[1440] : 
                       (N717)? mem[1456] : 
                       (N719)? mem[1472] : 
                       (N721)? mem[1488] : 
                       (N723)? mem[1504] : 
                       (N725)? mem[1520] : 
                       (N727)? mem[1536] : 
                       (N729)? mem[1552] : 
                       (N731)? mem[1568] : 
                       (N733)? mem[1584] : 
                       (N735)? mem[1600] : 
                       (N737)? mem[1616] : 
                       (N739)? mem[1632] : 
                       (N741)? mem[1648] : 
                       (N743)? mem[1664] : 
                       (N745)? mem[1680] : 
                       (N747)? mem[1696] : 
                       (N749)? mem[1712] : 
                       (N751)? mem[1728] : 
                       (N753)? mem[1744] : 
                       (N755)? mem[1760] : 
                       (N757)? mem[1776] : 
                       (N759)? mem[1792] : 
                       (N761)? mem[1808] : 
                       (N763)? mem[1824] : 
                       (N765)? mem[1840] : 
                       (N767)? mem[1856] : 
                       (N769)? mem[1872] : 
                       (N771)? mem[1888] : 
                       (N773)? mem[1904] : 
                       (N775)? mem[1920] : 
                       (N777)? mem[1936] : 
                       (N779)? mem[1952] : 
                       (N781)? mem[1968] : 
                       (N783)? mem[1984] : 
                       (N785)? mem[2000] : 
                       (N787)? mem[2016] : 
                       (N789)? mem[2032] : 
                       (N791)? mem[2048] : 
                       (N793)? mem[2064] : 
                       (N795)? mem[2080] : 
                       (N797)? mem[2096] : 
                       (N799)? mem[2112] : 
                       (N801)? mem[2128] : 
                       (N803)? mem[2144] : 
                       (N805)? mem[2160] : 
                       (N807)? mem[2176] : 
                       (N809)? mem[2192] : 
                       (N811)? mem[2208] : 
                       (N813)? mem[2224] : 
                       (N815)? mem[2240] : 
                       (N817)? mem[2256] : 
                       (N819)? mem[2272] : 
                       (N821)? mem[2288] : 
                       (N823)? mem[2304] : 
                       (N825)? mem[2320] : 
                       (N827)? mem[2336] : 
                       (N829)? mem[2352] : 
                       (N831)? mem[2368] : 
                       (N833)? mem[2384] : 
                       (N835)? mem[2400] : 
                       (N837)? mem[2416] : 
                       (N839)? mem[2432] : 
                       (N841)? mem[2448] : 
                       (N843)? mem[2464] : 
                       (N845)? mem[2480] : 
                       (N847)? mem[2496] : 
                       (N849)? mem[2512] : 
                       (N851)? mem[2528] : 
                       (N853)? mem[2544] : 
                       (N855)? mem[2560] : 
                       (N857)? mem[2576] : 
                       (N859)? mem[2592] : 
                       (N861)? mem[2608] : 
                       (N863)? mem[2624] : 
                       (N865)? mem[2640] : 
                       (N867)? mem[2656] : 
                       (N869)? mem[2672] : 
                       (N871)? mem[2688] : 
                       (N873)? mem[2704] : 
                       (N875)? mem[2720] : 
                       (N877)? mem[2736] : 
                       (N879)? mem[2752] : 
                       (N881)? mem[2768] : 
                       (N883)? mem[2784] : 
                       (N885)? mem[2800] : 
                       (N887)? mem[2816] : 
                       (N889)? mem[2832] : 
                       (N891)? mem[2848] : 
                       (N893)? mem[2864] : 
                       (N895)? mem[2880] : 
                       (N897)? mem[2896] : 
                       (N899)? mem[2912] : 
                       (N901)? mem[2928] : 
                       (N903)? mem[2944] : 
                       (N905)? mem[2960] : 
                       (N907)? mem[2976] : 
                       (N909)? mem[2992] : 
                       (N911)? mem[3008] : 
                       (N913)? mem[3024] : 
                       (N915)? mem[3040] : 
                       (N917)? mem[3056] : 
                       (N919)? mem[3072] : 
                       (N921)? mem[3088] : 
                       (N923)? mem[3104] : 
                       (N925)? mem[3120] : 
                       (N927)? mem[3136] : 
                       (N929)? mem[3152] : 
                       (N931)? mem[3168] : 
                       (N933)? mem[3184] : 
                       (N935)? mem[3200] : 
                       (N937)? mem[3216] : 
                       (N939)? mem[3232] : 
                       (N941)? mem[3248] : 
                       (N943)? mem[3264] : 
                       (N945)? mem[3280] : 
                       (N947)? mem[3296] : 
                       (N949)? mem[3312] : 
                       (N951)? mem[3328] : 
                       (N953)? mem[3344] : 
                       (N955)? mem[3360] : 
                       (N957)? mem[3376] : 
                       (N959)? mem[3392] : 
                       (N961)? mem[3408] : 
                       (N963)? mem[3424] : 
                       (N965)? mem[3440] : 
                       (N967)? mem[3456] : 
                       (N969)? mem[3472] : 
                       (N971)? mem[3488] : 
                       (N973)? mem[3504] : 
                       (N975)? mem[3520] : 
                       (N977)? mem[3536] : 
                       (N979)? mem[3552] : 
                       (N981)? mem[3568] : 
                       (N983)? mem[3584] : 
                       (N985)? mem[3600] : 
                       (N987)? mem[3616] : 
                       (N989)? mem[3632] : 
                       (N991)? mem[3648] : 
                       (N993)? mem[3664] : 
                       (N995)? mem[3680] : 
                       (N997)? mem[3696] : 
                       (N999)? mem[3712] : 
                       (N1001)? mem[3728] : 
                       (N1003)? mem[3744] : 
                       (N1005)? mem[3760] : 
                       (N1007)? mem[3776] : 
                       (N1009)? mem[3792] : 
                       (N1011)? mem[3808] : 
                       (N1013)? mem[3824] : 
                       (N1015)? mem[3840] : 
                       (N1017)? mem[3856] : 
                       (N1019)? mem[3872] : 
                       (N1021)? mem[3888] : 
                       (N1023)? mem[3904] : 
                       (N1025)? mem[3920] : 
                       (N1027)? mem[3936] : 
                       (N1029)? mem[3952] : 
                       (N1031)? mem[3968] : 
                       (N1033)? mem[3984] : 
                       (N1035)? mem[4000] : 
                       (N1037)? mem[4016] : 
                       (N1039)? mem[4032] : 
                       (N1041)? mem[4048] : 
                       (N1043)? mem[4064] : 
                       (N1045)? mem[4080] : 
                       (N536)? mem[4096] : 
                       (N538)? mem[4112] : 
                       (N540)? mem[4128] : 
                       (N542)? mem[4144] : 
                       (N544)? mem[4160] : 
                       (N546)? mem[4176] : 
                       (N548)? mem[4192] : 
                       (N550)? mem[4208] : 
                       (N552)? mem[4224] : 
                       (N554)? mem[4240] : 
                       (N556)? mem[4256] : 
                       (N558)? mem[4272] : 
                       (N560)? mem[4288] : 
                       (N562)? mem[4304] : 
                       (N564)? mem[4320] : 
                       (N566)? mem[4336] : 
                       (N568)? mem[4352] : 
                       (N570)? mem[4368] : 
                       (N572)? mem[4384] : 
                       (N574)? mem[4400] : 
                       (N576)? mem[4416] : 
                       (N578)? mem[4432] : 
                       (N580)? mem[4448] : 
                       (N582)? mem[4464] : 
                       (N584)? mem[4480] : 
                       (N586)? mem[4496] : 
                       (N588)? mem[4512] : 
                       (N590)? mem[4528] : 
                       (N592)? mem[4544] : 
                       (N594)? mem[4560] : 
                       (N596)? mem[4576] : 
                       (N598)? mem[4592] : 
                       (N600)? mem[4608] : 
                       (N602)? mem[4624] : 
                       (N604)? mem[4640] : 
                       (N606)? mem[4656] : 
                       (N608)? mem[4672] : 
                       (N610)? mem[4688] : 
                       (N612)? mem[4704] : 
                       (N614)? mem[4720] : 
                       (N616)? mem[4736] : 
                       (N618)? mem[4752] : 
                       (N620)? mem[4768] : 
                       (N622)? mem[4784] : 
                       (N624)? mem[4800] : 
                       (N626)? mem[4816] : 
                       (N628)? mem[4832] : 
                       (N630)? mem[4848] : 
                       (N632)? mem[4864] : 
                       (N634)? mem[4880] : 
                       (N636)? mem[4896] : 
                       (N638)? mem[4912] : 
                       (N640)? mem[4928] : 
                       (N642)? mem[4944] : 
                       (N644)? mem[4960] : 
                       (N646)? mem[4976] : 
                       (N648)? mem[4992] : 
                       (N650)? mem[5008] : 
                       (N652)? mem[5024] : 
                       (N654)? mem[5040] : 
                       (N656)? mem[5056] : 
                       (N658)? mem[5072] : 
                       (N660)? mem[5088] : 
                       (N662)? mem[5104] : 
                       (N664)? mem[5120] : 
                       (N666)? mem[5136] : 
                       (N668)? mem[5152] : 
                       (N670)? mem[5168] : 
                       (N672)? mem[5184] : 
                       (N674)? mem[5200] : 
                       (N676)? mem[5216] : 
                       (N678)? mem[5232] : 
                       (N680)? mem[5248] : 
                       (N682)? mem[5264] : 
                       (N684)? mem[5280] : 
                       (N686)? mem[5296] : 
                       (N688)? mem[5312] : 
                       (N690)? mem[5328] : 
                       (N692)? mem[5344] : 
                       (N694)? mem[5360] : 
                       (N696)? mem[5376] : 
                       (N698)? mem[5392] : 
                       (N700)? mem[5408] : 
                       (N702)? mem[5424] : 
                       (N704)? mem[5440] : 
                       (N706)? mem[5456] : 
                       (N708)? mem[5472] : 
                       (N710)? mem[5488] : 
                       (N712)? mem[5504] : 
                       (N714)? mem[5520] : 
                       (N716)? mem[5536] : 
                       (N718)? mem[5552] : 
                       (N720)? mem[5568] : 
                       (N722)? mem[5584] : 
                       (N724)? mem[5600] : 
                       (N726)? mem[5616] : 
                       (N728)? mem[5632] : 
                       (N730)? mem[5648] : 
                       (N732)? mem[5664] : 
                       (N734)? mem[5680] : 
                       (N736)? mem[5696] : 
                       (N738)? mem[5712] : 
                       (N740)? mem[5728] : 
                       (N742)? mem[5744] : 
                       (N744)? mem[5760] : 
                       (N746)? mem[5776] : 
                       (N748)? mem[5792] : 
                       (N750)? mem[5808] : 
                       (N752)? mem[5824] : 
                       (N754)? mem[5840] : 
                       (N756)? mem[5856] : 
                       (N758)? mem[5872] : 
                       (N760)? mem[5888] : 
                       (N762)? mem[5904] : 
                       (N764)? mem[5920] : 
                       (N766)? mem[5936] : 
                       (N768)? mem[5952] : 
                       (N770)? mem[5968] : 
                       (N772)? mem[5984] : 
                       (N774)? mem[6000] : 
                       (N776)? mem[6016] : 
                       (N778)? mem[6032] : 
                       (N780)? mem[6048] : 
                       (N782)? mem[6064] : 
                       (N784)? mem[6080] : 
                       (N786)? mem[6096] : 
                       (N788)? mem[6112] : 
                       (N790)? mem[6128] : 
                       (N792)? mem[6144] : 
                       (N794)? mem[6160] : 
                       (N796)? mem[6176] : 
                       (N798)? mem[6192] : 
                       (N800)? mem[6208] : 
                       (N802)? mem[6224] : 
                       (N804)? mem[6240] : 
                       (N806)? mem[6256] : 
                       (N808)? mem[6272] : 
                       (N810)? mem[6288] : 
                       (N812)? mem[6304] : 
                       (N814)? mem[6320] : 
                       (N816)? mem[6336] : 
                       (N818)? mem[6352] : 
                       (N820)? mem[6368] : 
                       (N822)? mem[6384] : 
                       (N824)? mem[6400] : 
                       (N826)? mem[6416] : 
                       (N828)? mem[6432] : 
                       (N830)? mem[6448] : 
                       (N832)? mem[6464] : 
                       (N834)? mem[6480] : 
                       (N836)? mem[6496] : 
                       (N838)? mem[6512] : 
                       (N840)? mem[6528] : 
                       (N842)? mem[6544] : 
                       (N844)? mem[6560] : 
                       (N846)? mem[6576] : 
                       (N848)? mem[6592] : 
                       (N850)? mem[6608] : 
                       (N852)? mem[6624] : 
                       (N854)? mem[6640] : 
                       (N856)? mem[6656] : 
                       (N858)? mem[6672] : 
                       (N860)? mem[6688] : 
                       (N862)? mem[6704] : 
                       (N864)? mem[6720] : 
                       (N866)? mem[6736] : 
                       (N868)? mem[6752] : 
                       (N870)? mem[6768] : 
                       (N872)? mem[6784] : 
                       (N874)? mem[6800] : 
                       (N876)? mem[6816] : 
                       (N878)? mem[6832] : 
                       (N880)? mem[6848] : 
                       (N882)? mem[6864] : 
                       (N884)? mem[6880] : 
                       (N886)? mem[6896] : 
                       (N888)? mem[6912] : 
                       (N890)? mem[6928] : 
                       (N892)? mem[6944] : 
                       (N894)? mem[6960] : 
                       (N896)? mem[6976] : 
                       (N898)? mem[6992] : 
                       (N900)? mem[7008] : 
                       (N902)? mem[7024] : 
                       (N904)? mem[7040] : 
                       (N906)? mem[7056] : 
                       (N908)? mem[7072] : 
                       (N910)? mem[7088] : 
                       (N912)? mem[7104] : 
                       (N914)? mem[7120] : 
                       (N916)? mem[7136] : 
                       (N918)? mem[7152] : 
                       (N920)? mem[7168] : 
                       (N922)? mem[7184] : 
                       (N924)? mem[7200] : 
                       (N926)? mem[7216] : 
                       (N928)? mem[7232] : 
                       (N930)? mem[7248] : 
                       (N932)? mem[7264] : 
                       (N934)? mem[7280] : 
                       (N936)? mem[7296] : 
                       (N938)? mem[7312] : 
                       (N940)? mem[7328] : 
                       (N942)? mem[7344] : 
                       (N944)? mem[7360] : 
                       (N946)? mem[7376] : 
                       (N948)? mem[7392] : 
                       (N950)? mem[7408] : 
                       (N952)? mem[7424] : 
                       (N954)? mem[7440] : 
                       (N956)? mem[7456] : 
                       (N958)? mem[7472] : 
                       (N960)? mem[7488] : 
                       (N962)? mem[7504] : 
                       (N964)? mem[7520] : 
                       (N966)? mem[7536] : 
                       (N968)? mem[7552] : 
                       (N970)? mem[7568] : 
                       (N972)? mem[7584] : 
                       (N974)? mem[7600] : 
                       (N976)? mem[7616] : 
                       (N978)? mem[7632] : 
                       (N980)? mem[7648] : 
                       (N982)? mem[7664] : 
                       (N984)? mem[7680] : 
                       (N986)? mem[7696] : 
                       (N988)? mem[7712] : 
                       (N990)? mem[7728] : 
                       (N992)? mem[7744] : 
                       (N994)? mem[7760] : 
                       (N996)? mem[7776] : 
                       (N998)? mem[7792] : 
                       (N1000)? mem[7808] : 
                       (N1002)? mem[7824] : 
                       (N1004)? mem[7840] : 
                       (N1006)? mem[7856] : 
                       (N1008)? mem[7872] : 
                       (N1010)? mem[7888] : 
                       (N1012)? mem[7904] : 
                       (N1014)? mem[7920] : 
                       (N1016)? mem[7936] : 
                       (N1018)? mem[7952] : 
                       (N1020)? mem[7968] : 
                       (N1022)? mem[7984] : 
                       (N1024)? mem[8000] : 
                       (N1026)? mem[8016] : 
                       (N1028)? mem[8032] : 
                       (N1030)? mem[8048] : 
                       (N1032)? mem[8064] : 
                       (N1034)? mem[8080] : 
                       (N1036)? mem[8096] : 
                       (N1038)? mem[8112] : 
                       (N1040)? mem[8128] : 
                       (N1042)? mem[8144] : 
                       (N1044)? mem[8160] : 
                       (N1046)? mem[8176] : 1'b0;
  assign N2072 = w_addr_i[7] & w_addr_i[8];
  assign N2073 = N0 & w_addr_i[8];
  assign N0 = ~w_addr_i[7];
  assign N2074 = w_addr_i[7] & N1;
  assign N1 = ~w_addr_i[8];
  assign N2075 = N2 & N3;
  assign N2 = ~w_addr_i[7];
  assign N3 = ~w_addr_i[8];
  assign N2076 = w_addr_i[5] & w_addr_i[6];
  assign N2077 = N4 & w_addr_i[6];
  assign N4 = ~w_addr_i[5];
  assign N2078 = w_addr_i[5] & N5;
  assign N5 = ~w_addr_i[6];
  assign N2079 = N6 & N7;
  assign N6 = ~w_addr_i[5];
  assign N7 = ~w_addr_i[6];
  assign N2080 = N2072 & N2076;
  assign N2081 = N2072 & N2077;
  assign N2082 = N2072 & N2078;
  assign N2083 = N2072 & N2079;
  assign N2084 = N2073 & N2076;
  assign N2085 = N2073 & N2077;
  assign N2086 = N2073 & N2078;
  assign N2087 = N2073 & N2079;
  assign N2088 = N2074 & N2076;
  assign N2089 = N2074 & N2077;
  assign N2090 = N2074 & N2078;
  assign N2091 = N2074 & N2079;
  assign N2092 = N2075 & N2076;
  assign N2093 = N2075 & N2077;
  assign N2094 = N2075 & N2078;
  assign N2095 = N2075 & N2079;
  assign N2096 = w_addr_i[3] & w_addr_i[4];
  assign N2097 = N8 & w_addr_i[4];
  assign N8 = ~w_addr_i[3];
  assign N2098 = w_addr_i[3] & N9;
  assign N9 = ~w_addr_i[4];
  assign N2099 = N10 & N11;
  assign N10 = ~w_addr_i[3];
  assign N11 = ~w_addr_i[4];
  assign N2100 = ~w_addr_i[2];
  assign N2101 = w_addr_i[0] & w_addr_i[1];
  assign N2102 = N12 & w_addr_i[1];
  assign N12 = ~w_addr_i[0];
  assign N2103 = w_addr_i[0] & N13;
  assign N13 = ~w_addr_i[1];
  assign N2104 = N14 & N15;
  assign N14 = ~w_addr_i[0];
  assign N15 = ~w_addr_i[1];
  assign N2105 = w_addr_i[2] & N2101;
  assign N2106 = w_addr_i[2] & N2102;
  assign N2107 = w_addr_i[2] & N2103;
  assign N2108 = w_addr_i[2] & N2104;
  assign N2109 = N2100 & N2101;
  assign N2110 = N2100 & N2102;
  assign N2111 = N2100 & N2103;
  assign N2112 = N2100 & N2104;
  assign N2113 = N2096 & N2105;
  assign N2114 = N2096 & N2106;
  assign N2115 = N2096 & N2107;
  assign N2116 = N2096 & N2108;
  assign N2117 = N2096 & N2109;
  assign N2118 = N2096 & N2110;
  assign N2119 = N2096 & N2111;
  assign N2120 = N2096 & N2112;
  assign N2121 = N2097 & N2105;
  assign N2122 = N2097 & N2106;
  assign N2123 = N2097 & N2107;
  assign N2124 = N2097 & N2108;
  assign N2125 = N2097 & N2109;
  assign N2126 = N2097 & N2110;
  assign N2127 = N2097 & N2111;
  assign N2128 = N2097 & N2112;
  assign N2129 = N2098 & N2105;
  assign N2130 = N2098 & N2106;
  assign N2131 = N2098 & N2107;
  assign N2132 = N2098 & N2108;
  assign N2133 = N2098 & N2109;
  assign N2134 = N2098 & N2110;
  assign N2135 = N2098 & N2111;
  assign N2136 = N2098 & N2112;
  assign N2137 = N2099 & N2105;
  assign N2138 = N2099 & N2106;
  assign N2139 = N2099 & N2107;
  assign N2140 = N2099 & N2108;
  assign N2141 = N2099 & N2109;
  assign N2142 = N2099 & N2110;
  assign N2143 = N2099 & N2111;
  assign N2144 = N2099 & N2112;
  assign N1559 = N2080 & N2113;
  assign N1558 = N2080 & N2114;
  assign N1557 = N2080 & N2115;
  assign N1556 = N2080 & N2116;
  assign N1555 = N2080 & N2117;
  assign N1554 = N2080 & N2118;
  assign N1553 = N2080 & N2119;
  assign N1552 = N2080 & N2120;
  assign N1551 = N2080 & N2121;
  assign N1550 = N2080 & N2122;
  assign N1549 = N2080 & N2123;
  assign N1548 = N2080 & N2124;
  assign N1547 = N2080 & N2125;
  assign N1546 = N2080 & N2126;
  assign N1545 = N2080 & N2127;
  assign N1544 = N2080 & N2128;
  assign N1543 = N2080 & N2129;
  assign N1542 = N2080 & N2130;
  assign N1541 = N2080 & N2131;
  assign N1540 = N2080 & N2132;
  assign N1539 = N2080 & N2133;
  assign N1538 = N2080 & N2134;
  assign N1537 = N2080 & N2135;
  assign N1536 = N2080 & N2136;
  assign N1535 = N2080 & N2137;
  assign N1534 = N2080 & N2138;
  assign N1533 = N2080 & N2139;
  assign N1532 = N2080 & N2140;
  assign N1531 = N2080 & N2141;
  assign N1530 = N2080 & N2142;
  assign N1529 = N2080 & N2143;
  assign N1528 = N2080 & N2144;
  assign N1527 = N2081 & N2113;
  assign N1526 = N2081 & N2114;
  assign N1525 = N2081 & N2115;
  assign N1524 = N2081 & N2116;
  assign N1523 = N2081 & N2117;
  assign N1522 = N2081 & N2118;
  assign N1521 = N2081 & N2119;
  assign N1520 = N2081 & N2120;
  assign N1519 = N2081 & N2121;
  assign N1518 = N2081 & N2122;
  assign N1517 = N2081 & N2123;
  assign N1516 = N2081 & N2124;
  assign N1515 = N2081 & N2125;
  assign N1514 = N2081 & N2126;
  assign N1513 = N2081 & N2127;
  assign N1512 = N2081 & N2128;
  assign N1511 = N2081 & N2129;
  assign N1510 = N2081 & N2130;
  assign N1509 = N2081 & N2131;
  assign N1508 = N2081 & N2132;
  assign N1507 = N2081 & N2133;
  assign N1506 = N2081 & N2134;
  assign N1505 = N2081 & N2135;
  assign N1504 = N2081 & N2136;
  assign N1503 = N2081 & N2137;
  assign N1502 = N2081 & N2138;
  assign N1501 = N2081 & N2139;
  assign N1500 = N2081 & N2140;
  assign N1499 = N2081 & N2141;
  assign N1498 = N2081 & N2142;
  assign N1497 = N2081 & N2143;
  assign N1496 = N2081 & N2144;
  assign N1495 = N2082 & N2113;
  assign N1494 = N2082 & N2114;
  assign N1493 = N2082 & N2115;
  assign N1492 = N2082 & N2116;
  assign N1491 = N2082 & N2117;
  assign N1490 = N2082 & N2118;
  assign N1489 = N2082 & N2119;
  assign N1488 = N2082 & N2120;
  assign N1487 = N2082 & N2121;
  assign N1486 = N2082 & N2122;
  assign N1485 = N2082 & N2123;
  assign N1484 = N2082 & N2124;
  assign N1483 = N2082 & N2125;
  assign N1482 = N2082 & N2126;
  assign N1481 = N2082 & N2127;
  assign N1480 = N2082 & N2128;
  assign N1479 = N2082 & N2129;
  assign N1478 = N2082 & N2130;
  assign N1477 = N2082 & N2131;
  assign N1476 = N2082 & N2132;
  assign N1475 = N2082 & N2133;
  assign N1474 = N2082 & N2134;
  assign N1473 = N2082 & N2135;
  assign N1472 = N2082 & N2136;
  assign N1471 = N2082 & N2137;
  assign N1470 = N2082 & N2138;
  assign N1469 = N2082 & N2139;
  assign N1468 = N2082 & N2140;
  assign N1467 = N2082 & N2141;
  assign N1466 = N2082 & N2142;
  assign N1465 = N2082 & N2143;
  assign N1464 = N2082 & N2144;
  assign N1463 = N2083 & N2113;
  assign N1462 = N2083 & N2114;
  assign N1461 = N2083 & N2115;
  assign N1460 = N2083 & N2116;
  assign N1459 = N2083 & N2117;
  assign N1458 = N2083 & N2118;
  assign N1457 = N2083 & N2119;
  assign N1456 = N2083 & N2120;
  assign N1455 = N2083 & N2121;
  assign N1454 = N2083 & N2122;
  assign N1453 = N2083 & N2123;
  assign N1452 = N2083 & N2124;
  assign N1451 = N2083 & N2125;
  assign N1450 = N2083 & N2126;
  assign N1449 = N2083 & N2127;
  assign N1448 = N2083 & N2128;
  assign N1447 = N2083 & N2129;
  assign N1446 = N2083 & N2130;
  assign N1445 = N2083 & N2131;
  assign N1444 = N2083 & N2132;
  assign N1443 = N2083 & N2133;
  assign N1442 = N2083 & N2134;
  assign N1441 = N2083 & N2135;
  assign N1440 = N2083 & N2136;
  assign N1439 = N2083 & N2137;
  assign N1438 = N2083 & N2138;
  assign N1437 = N2083 & N2139;
  assign N1436 = N2083 & N2140;
  assign N1435 = N2083 & N2141;
  assign N1434 = N2083 & N2142;
  assign N1433 = N2083 & N2143;
  assign N1432 = N2083 & N2144;
  assign N1431 = N2084 & N2113;
  assign N1430 = N2084 & N2114;
  assign N1429 = N2084 & N2115;
  assign N1428 = N2084 & N2116;
  assign N1427 = N2084 & N2117;
  assign N1426 = N2084 & N2118;
  assign N1425 = N2084 & N2119;
  assign N1424 = N2084 & N2120;
  assign N1423 = N2084 & N2121;
  assign N1422 = N2084 & N2122;
  assign N1421 = N2084 & N2123;
  assign N1420 = N2084 & N2124;
  assign N1419 = N2084 & N2125;
  assign N1418 = N2084 & N2126;
  assign N1417 = N2084 & N2127;
  assign N1416 = N2084 & N2128;
  assign N1415 = N2084 & N2129;
  assign N1414 = N2084 & N2130;
  assign N1413 = N2084 & N2131;
  assign N1412 = N2084 & N2132;
  assign N1411 = N2084 & N2133;
  assign N1410 = N2084 & N2134;
  assign N1409 = N2084 & N2135;
  assign N1408 = N2084 & N2136;
  assign N1407 = N2084 & N2137;
  assign N1406 = N2084 & N2138;
  assign N1405 = N2084 & N2139;
  assign N1404 = N2084 & N2140;
  assign N1403 = N2084 & N2141;
  assign N1402 = N2084 & N2142;
  assign N1401 = N2084 & N2143;
  assign N1400 = N2084 & N2144;
  assign N1399 = N2085 & N2113;
  assign N1398 = N2085 & N2114;
  assign N1397 = N2085 & N2115;
  assign N1396 = N2085 & N2116;
  assign N1395 = N2085 & N2117;
  assign N1394 = N2085 & N2118;
  assign N1393 = N2085 & N2119;
  assign N1392 = N2085 & N2120;
  assign N1391 = N2085 & N2121;
  assign N1390 = N2085 & N2122;
  assign N1389 = N2085 & N2123;
  assign N1388 = N2085 & N2124;
  assign N1387 = N2085 & N2125;
  assign N1386 = N2085 & N2126;
  assign N1385 = N2085 & N2127;
  assign N1384 = N2085 & N2128;
  assign N1383 = N2085 & N2129;
  assign N1382 = N2085 & N2130;
  assign N1381 = N2085 & N2131;
  assign N1380 = N2085 & N2132;
  assign N1379 = N2085 & N2133;
  assign N1378 = N2085 & N2134;
  assign N1377 = N2085 & N2135;
  assign N1376 = N2085 & N2136;
  assign N1375 = N2085 & N2137;
  assign N1374 = N2085 & N2138;
  assign N1373 = N2085 & N2139;
  assign N1372 = N2085 & N2140;
  assign N1371 = N2085 & N2141;
  assign N1370 = N2085 & N2142;
  assign N1369 = N2085 & N2143;
  assign N1368 = N2085 & N2144;
  assign N1367 = N2086 & N2113;
  assign N1366 = N2086 & N2114;
  assign N1365 = N2086 & N2115;
  assign N1364 = N2086 & N2116;
  assign N1363 = N2086 & N2117;
  assign N1362 = N2086 & N2118;
  assign N1361 = N2086 & N2119;
  assign N1360 = N2086 & N2120;
  assign N1359 = N2086 & N2121;
  assign N1358 = N2086 & N2122;
  assign N1357 = N2086 & N2123;
  assign N1356 = N2086 & N2124;
  assign N1355 = N2086 & N2125;
  assign N1354 = N2086 & N2126;
  assign N1353 = N2086 & N2127;
  assign N1352 = N2086 & N2128;
  assign N1351 = N2086 & N2129;
  assign N1350 = N2086 & N2130;
  assign N1349 = N2086 & N2131;
  assign N1348 = N2086 & N2132;
  assign N1347 = N2086 & N2133;
  assign N1346 = N2086 & N2134;
  assign N1345 = N2086 & N2135;
  assign N1344 = N2086 & N2136;
  assign N1343 = N2086 & N2137;
  assign N1342 = N2086 & N2138;
  assign N1341 = N2086 & N2139;
  assign N1340 = N2086 & N2140;
  assign N1339 = N2086 & N2141;
  assign N1338 = N2086 & N2142;
  assign N1337 = N2086 & N2143;
  assign N1336 = N2086 & N2144;
  assign N1335 = N2087 & N2113;
  assign N1334 = N2087 & N2114;
  assign N1333 = N2087 & N2115;
  assign N1332 = N2087 & N2116;
  assign N1331 = N2087 & N2117;
  assign N1330 = N2087 & N2118;
  assign N1329 = N2087 & N2119;
  assign N1328 = N2087 & N2120;
  assign N1327 = N2087 & N2121;
  assign N1326 = N2087 & N2122;
  assign N1325 = N2087 & N2123;
  assign N1324 = N2087 & N2124;
  assign N1323 = N2087 & N2125;
  assign N1322 = N2087 & N2126;
  assign N1321 = N2087 & N2127;
  assign N1320 = N2087 & N2128;
  assign N1319 = N2087 & N2129;
  assign N1318 = N2087 & N2130;
  assign N1317 = N2087 & N2131;
  assign N1316 = N2087 & N2132;
  assign N1315 = N2087 & N2133;
  assign N1314 = N2087 & N2134;
  assign N1313 = N2087 & N2135;
  assign N1312 = N2087 & N2136;
  assign N1311 = N2087 & N2137;
  assign N1310 = N2087 & N2138;
  assign N1309 = N2087 & N2139;
  assign N1308 = N2087 & N2140;
  assign N1307 = N2087 & N2141;
  assign N1306 = N2087 & N2142;
  assign N1305 = N2087 & N2143;
  assign N1304 = N2087 & N2144;
  assign N1303 = N2088 & N2113;
  assign N1302 = N2088 & N2114;
  assign N1301 = N2088 & N2115;
  assign N1300 = N2088 & N2116;
  assign N1299 = N2088 & N2117;
  assign N1298 = N2088 & N2118;
  assign N1297 = N2088 & N2119;
  assign N1296 = N2088 & N2120;
  assign N1295 = N2088 & N2121;
  assign N1294 = N2088 & N2122;
  assign N1293 = N2088 & N2123;
  assign N1292 = N2088 & N2124;
  assign N1291 = N2088 & N2125;
  assign N1290 = N2088 & N2126;
  assign N1289 = N2088 & N2127;
  assign N1288 = N2088 & N2128;
  assign N1287 = N2088 & N2129;
  assign N1286 = N2088 & N2130;
  assign N1285 = N2088 & N2131;
  assign N1284 = N2088 & N2132;
  assign N1283 = N2088 & N2133;
  assign N1282 = N2088 & N2134;
  assign N1281 = N2088 & N2135;
  assign N1280 = N2088 & N2136;
  assign N1279 = N2088 & N2137;
  assign N1278 = N2088 & N2138;
  assign N1277 = N2088 & N2139;
  assign N1276 = N2088 & N2140;
  assign N1275 = N2088 & N2141;
  assign N1274 = N2088 & N2142;
  assign N1273 = N2088 & N2143;
  assign N1272 = N2088 & N2144;
  assign N1271 = N2089 & N2113;
  assign N1270 = N2089 & N2114;
  assign N1269 = N2089 & N2115;
  assign N1268 = N2089 & N2116;
  assign N1267 = N2089 & N2117;
  assign N1266 = N2089 & N2118;
  assign N1265 = N2089 & N2119;
  assign N1264 = N2089 & N2120;
  assign N1263 = N2089 & N2121;
  assign N1262 = N2089 & N2122;
  assign N1261 = N2089 & N2123;
  assign N1260 = N2089 & N2124;
  assign N1259 = N2089 & N2125;
  assign N1258 = N2089 & N2126;
  assign N1257 = N2089 & N2127;
  assign N1256 = N2089 & N2128;
  assign N1255 = N2089 & N2129;
  assign N1254 = N2089 & N2130;
  assign N1253 = N2089 & N2131;
  assign N1252 = N2089 & N2132;
  assign N1251 = N2089 & N2133;
  assign N1250 = N2089 & N2134;
  assign N1249 = N2089 & N2135;
  assign N1248 = N2089 & N2136;
  assign N1247 = N2089 & N2137;
  assign N1246 = N2089 & N2138;
  assign N1245 = N2089 & N2139;
  assign N1244 = N2089 & N2140;
  assign N1243 = N2089 & N2141;
  assign N1242 = N2089 & N2142;
  assign N1241 = N2089 & N2143;
  assign N1240 = N2089 & N2144;
  assign N1239 = N2090 & N2113;
  assign N1238 = N2090 & N2114;
  assign N1237 = N2090 & N2115;
  assign N1236 = N2090 & N2116;
  assign N1235 = N2090 & N2117;
  assign N1234 = N2090 & N2118;
  assign N1233 = N2090 & N2119;
  assign N1232 = N2090 & N2120;
  assign N1231 = N2090 & N2121;
  assign N1230 = N2090 & N2122;
  assign N1229 = N2090 & N2123;
  assign N1228 = N2090 & N2124;
  assign N1227 = N2090 & N2125;
  assign N1226 = N2090 & N2126;
  assign N1225 = N2090 & N2127;
  assign N1224 = N2090 & N2128;
  assign N1223 = N2090 & N2129;
  assign N1222 = N2090 & N2130;
  assign N1221 = N2090 & N2131;
  assign N1220 = N2090 & N2132;
  assign N1219 = N2090 & N2133;
  assign N1218 = N2090 & N2134;
  assign N1217 = N2090 & N2135;
  assign N1216 = N2090 & N2136;
  assign N1215 = N2090 & N2137;
  assign N1214 = N2090 & N2138;
  assign N1213 = N2090 & N2139;
  assign N1212 = N2090 & N2140;
  assign N1211 = N2090 & N2141;
  assign N1210 = N2090 & N2142;
  assign N1209 = N2090 & N2143;
  assign N1208 = N2090 & N2144;
  assign N1207 = N2091 & N2113;
  assign N1206 = N2091 & N2114;
  assign N1205 = N2091 & N2115;
  assign N1204 = N2091 & N2116;
  assign N1203 = N2091 & N2117;
  assign N1202 = N2091 & N2118;
  assign N1201 = N2091 & N2119;
  assign N1200 = N2091 & N2120;
  assign N1199 = N2091 & N2121;
  assign N1198 = N2091 & N2122;
  assign N1197 = N2091 & N2123;
  assign N1196 = N2091 & N2124;
  assign N1195 = N2091 & N2125;
  assign N1194 = N2091 & N2126;
  assign N1193 = N2091 & N2127;
  assign N1192 = N2091 & N2128;
  assign N1191 = N2091 & N2129;
  assign N1190 = N2091 & N2130;
  assign N1189 = N2091 & N2131;
  assign N1188 = N2091 & N2132;
  assign N1187 = N2091 & N2133;
  assign N1186 = N2091 & N2134;
  assign N1185 = N2091 & N2135;
  assign N1184 = N2091 & N2136;
  assign N1183 = N2091 & N2137;
  assign N1182 = N2091 & N2138;
  assign N1181 = N2091 & N2139;
  assign N1180 = N2091 & N2140;
  assign N1179 = N2091 & N2141;
  assign N1178 = N2091 & N2142;
  assign N1177 = N2091 & N2143;
  assign N1176 = N2091 & N2144;
  assign N1175 = N2092 & N2113;
  assign N1174 = N2092 & N2114;
  assign N1173 = N2092 & N2115;
  assign N1172 = N2092 & N2116;
  assign N1171 = N2092 & N2117;
  assign N1170 = N2092 & N2118;
  assign N1169 = N2092 & N2119;
  assign N1168 = N2092 & N2120;
  assign N1167 = N2092 & N2121;
  assign N1166 = N2092 & N2122;
  assign N1165 = N2092 & N2123;
  assign N1164 = N2092 & N2124;
  assign N1163 = N2092 & N2125;
  assign N1162 = N2092 & N2126;
  assign N1161 = N2092 & N2127;
  assign N1160 = N2092 & N2128;
  assign N1159 = N2092 & N2129;
  assign N1158 = N2092 & N2130;
  assign N1157 = N2092 & N2131;
  assign N1156 = N2092 & N2132;
  assign N1155 = N2092 & N2133;
  assign N1154 = N2092 & N2134;
  assign N1153 = N2092 & N2135;
  assign N1152 = N2092 & N2136;
  assign N1151 = N2092 & N2137;
  assign N1150 = N2092 & N2138;
  assign N1149 = N2092 & N2139;
  assign N1148 = N2092 & N2140;
  assign N1147 = N2092 & N2141;
  assign N1146 = N2092 & N2142;
  assign N1145 = N2092 & N2143;
  assign N1144 = N2092 & N2144;
  assign N1143 = N2093 & N2113;
  assign N1142 = N2093 & N2114;
  assign N1141 = N2093 & N2115;
  assign N1140 = N2093 & N2116;
  assign N1139 = N2093 & N2117;
  assign N1138 = N2093 & N2118;
  assign N1137 = N2093 & N2119;
  assign N1136 = N2093 & N2120;
  assign N1135 = N2093 & N2121;
  assign N1134 = N2093 & N2122;
  assign N1133 = N2093 & N2123;
  assign N1132 = N2093 & N2124;
  assign N1131 = N2093 & N2125;
  assign N1130 = N2093 & N2126;
  assign N1129 = N2093 & N2127;
  assign N1128 = N2093 & N2128;
  assign N1127 = N2093 & N2129;
  assign N1126 = N2093 & N2130;
  assign N1125 = N2093 & N2131;
  assign N1124 = N2093 & N2132;
  assign N1123 = N2093 & N2133;
  assign N1122 = N2093 & N2134;
  assign N1121 = N2093 & N2135;
  assign N1120 = N2093 & N2136;
  assign N1119 = N2093 & N2137;
  assign N1118 = N2093 & N2138;
  assign N1117 = N2093 & N2139;
  assign N1116 = N2093 & N2140;
  assign N1115 = N2093 & N2141;
  assign N1114 = N2093 & N2142;
  assign N1113 = N2093 & N2143;
  assign N1112 = N2093 & N2144;
  assign N1111 = N2094 & N2113;
  assign N1110 = N2094 & N2114;
  assign N1109 = N2094 & N2115;
  assign N1108 = N2094 & N2116;
  assign N1107 = N2094 & N2117;
  assign N1106 = N2094 & N2118;
  assign N1105 = N2094 & N2119;
  assign N1104 = N2094 & N2120;
  assign N1103 = N2094 & N2121;
  assign N1102 = N2094 & N2122;
  assign N1101 = N2094 & N2123;
  assign N1100 = N2094 & N2124;
  assign N1099 = N2094 & N2125;
  assign N1098 = N2094 & N2126;
  assign N1097 = N2094 & N2127;
  assign N1096 = N2094 & N2128;
  assign N1095 = N2094 & N2129;
  assign N1094 = N2094 & N2130;
  assign N1093 = N2094 & N2131;
  assign N1092 = N2094 & N2132;
  assign N1091 = N2094 & N2133;
  assign N1090 = N2094 & N2134;
  assign N1089 = N2094 & N2135;
  assign N1088 = N2094 & N2136;
  assign N1087 = N2094 & N2137;
  assign N1086 = N2094 & N2138;
  assign N1085 = N2094 & N2139;
  assign N1084 = N2094 & N2140;
  assign N1083 = N2094 & N2141;
  assign N1082 = N2094 & N2142;
  assign N1081 = N2094 & N2143;
  assign N1080 = N2094 & N2144;
  assign N1079 = N2095 & N2113;
  assign N1078 = N2095 & N2114;
  assign N1077 = N2095 & N2115;
  assign N1076 = N2095 & N2116;
  assign N1075 = N2095 & N2117;
  assign N1074 = N2095 & N2118;
  assign N1073 = N2095 & N2119;
  assign N1072 = N2095 & N2120;
  assign N1071 = N2095 & N2121;
  assign N1070 = N2095 & N2122;
  assign N1069 = N2095 & N2123;
  assign N1068 = N2095 & N2124;
  assign N1067 = N2095 & N2125;
  assign N1066 = N2095 & N2126;
  assign N1065 = N2095 & N2127;
  assign N1064 = N2095 & N2128;
  assign N1063 = N2095 & N2129;
  assign N1062 = N2095 & N2130;
  assign N1061 = N2095 & N2131;
  assign N1060 = N2095 & N2132;
  assign N1059 = N2095 & N2133;
  assign N1058 = N2095 & N2134;
  assign N1057 = N2095 & N2135;
  assign N1056 = N2095 & N2136;
  assign N1055 = N2095 & N2137;
  assign N1054 = N2095 & N2138;
  assign N1053 = N2095 & N2139;
  assign N1052 = N2095 & N2140;
  assign N1051 = N2095 & N2141;
  assign N1050 = N2095 & N2142;
  assign N1049 = N2095 & N2143;
  assign N1048 = N2095 & N2144;
  assign { N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560 } = (N16)? { N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050, N1049, N1048 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N17)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = w_v_i;
  assign N17 = N1047;
  assign N18 = ~r_addr_r[0];
  assign N19 = ~r_addr_r[1];
  assign N20 = N18 & N19;
  assign N21 = N18 & r_addr_r[1];
  assign N22 = r_addr_r[0] & N19;
  assign N23 = r_addr_r[0] & r_addr_r[1];
  assign N24 = ~r_addr_r[2];
  assign N25 = N20 & N24;
  assign N26 = N20 & r_addr_r[2];
  assign N27 = N22 & N24;
  assign N28 = N22 & r_addr_r[2];
  assign N29 = N21 & N24;
  assign N30 = N21 & r_addr_r[2];
  assign N31 = N23 & N24;
  assign N32 = N23 & r_addr_r[2];
  assign N33 = ~r_addr_r[3];
  assign N34 = N25 & N33;
  assign N35 = N25 & r_addr_r[3];
  assign N36 = N27 & N33;
  assign N37 = N27 & r_addr_r[3];
  assign N38 = N29 & N33;
  assign N39 = N29 & r_addr_r[3];
  assign N40 = N31 & N33;
  assign N41 = N31 & r_addr_r[3];
  assign N42 = N26 & N33;
  assign N43 = N26 & r_addr_r[3];
  assign N44 = N28 & N33;
  assign N45 = N28 & r_addr_r[3];
  assign N46 = N30 & N33;
  assign N47 = N30 & r_addr_r[3];
  assign N48 = N32 & N33;
  assign N49 = N32 & r_addr_r[3];
  assign N50 = ~r_addr_r[4];
  assign N51 = N34 & N50;
  assign N52 = N34 & r_addr_r[4];
  assign N53 = N36 & N50;
  assign N54 = N36 & r_addr_r[4];
  assign N55 = N38 & N50;
  assign N56 = N38 & r_addr_r[4];
  assign N57 = N40 & N50;
  assign N58 = N40 & r_addr_r[4];
  assign N59 = N42 & N50;
  assign N60 = N42 & r_addr_r[4];
  assign N61 = N44 & N50;
  assign N62 = N44 & r_addr_r[4];
  assign N63 = N46 & N50;
  assign N64 = N46 & r_addr_r[4];
  assign N65 = N48 & N50;
  assign N66 = N48 & r_addr_r[4];
  assign N67 = N35 & N50;
  assign N68 = N35 & r_addr_r[4];
  assign N69 = N37 & N50;
  assign N70 = N37 & r_addr_r[4];
  assign N71 = N39 & N50;
  assign N72 = N39 & r_addr_r[4];
  assign N73 = N41 & N50;
  assign N74 = N41 & r_addr_r[4];
  assign N75 = N43 & N50;
  assign N76 = N43 & r_addr_r[4];
  assign N77 = N45 & N50;
  assign N78 = N45 & r_addr_r[4];
  assign N79 = N47 & N50;
  assign N80 = N47 & r_addr_r[4];
  assign N81 = N49 & N50;
  assign N82 = N49 & r_addr_r[4];
  assign N83 = ~r_addr_r[5];
  assign N84 = N51 & N83;
  assign N85 = N51 & r_addr_r[5];
  assign N86 = N53 & N83;
  assign N87 = N53 & r_addr_r[5];
  assign N88 = N55 & N83;
  assign N89 = N55 & r_addr_r[5];
  assign N90 = N57 & N83;
  assign N91 = N57 & r_addr_r[5];
  assign N92 = N59 & N83;
  assign N93 = N59 & r_addr_r[5];
  assign N94 = N61 & N83;
  assign N95 = N61 & r_addr_r[5];
  assign N96 = N63 & N83;
  assign N97 = N63 & r_addr_r[5];
  assign N98 = N65 & N83;
  assign N99 = N65 & r_addr_r[5];
  assign N100 = N67 & N83;
  assign N101 = N67 & r_addr_r[5];
  assign N102 = N69 & N83;
  assign N103 = N69 & r_addr_r[5];
  assign N104 = N71 & N83;
  assign N105 = N71 & r_addr_r[5];
  assign N106 = N73 & N83;
  assign N107 = N73 & r_addr_r[5];
  assign N108 = N75 & N83;
  assign N109 = N75 & r_addr_r[5];
  assign N110 = N77 & N83;
  assign N111 = N77 & r_addr_r[5];
  assign N112 = N79 & N83;
  assign N113 = N79 & r_addr_r[5];
  assign N114 = N81 & N83;
  assign N115 = N81 & r_addr_r[5];
  assign N116 = N52 & N83;
  assign N117 = N52 & r_addr_r[5];
  assign N118 = N54 & N83;
  assign N119 = N54 & r_addr_r[5];
  assign N120 = N56 & N83;
  assign N121 = N56 & r_addr_r[5];
  assign N122 = N58 & N83;
  assign N123 = N58 & r_addr_r[5];
  assign N124 = N60 & N83;
  assign N125 = N60 & r_addr_r[5];
  assign N126 = N62 & N83;
  assign N127 = N62 & r_addr_r[5];
  assign N128 = N64 & N83;
  assign N129 = N64 & r_addr_r[5];
  assign N130 = N66 & N83;
  assign N131 = N66 & r_addr_r[5];
  assign N132 = N68 & N83;
  assign N133 = N68 & r_addr_r[5];
  assign N134 = N70 & N83;
  assign N135 = N70 & r_addr_r[5];
  assign N136 = N72 & N83;
  assign N137 = N72 & r_addr_r[5];
  assign N138 = N74 & N83;
  assign N139 = N74 & r_addr_r[5];
  assign N140 = N76 & N83;
  assign N141 = N76 & r_addr_r[5];
  assign N142 = N78 & N83;
  assign N143 = N78 & r_addr_r[5];
  assign N144 = N80 & N83;
  assign N145 = N80 & r_addr_r[5];
  assign N146 = N82 & N83;
  assign N147 = N82 & r_addr_r[5];
  assign N148 = ~r_addr_r[6];
  assign N149 = N84 & N148;
  assign N150 = N84 & r_addr_r[6];
  assign N151 = N86 & N148;
  assign N152 = N86 & r_addr_r[6];
  assign N153 = N88 & N148;
  assign N154 = N88 & r_addr_r[6];
  assign N155 = N90 & N148;
  assign N156 = N90 & r_addr_r[6];
  assign N157 = N92 & N148;
  assign N158 = N92 & r_addr_r[6];
  assign N159 = N94 & N148;
  assign N160 = N94 & r_addr_r[6];
  assign N161 = N96 & N148;
  assign N162 = N96 & r_addr_r[6];
  assign N163 = N98 & N148;
  assign N164 = N98 & r_addr_r[6];
  assign N165 = N100 & N148;
  assign N166 = N100 & r_addr_r[6];
  assign N167 = N102 & N148;
  assign N168 = N102 & r_addr_r[6];
  assign N169 = N104 & N148;
  assign N170 = N104 & r_addr_r[6];
  assign N171 = N106 & N148;
  assign N172 = N106 & r_addr_r[6];
  assign N173 = N108 & N148;
  assign N174 = N108 & r_addr_r[6];
  assign N175 = N110 & N148;
  assign N176 = N110 & r_addr_r[6];
  assign N177 = N112 & N148;
  assign N178 = N112 & r_addr_r[6];
  assign N179 = N114 & N148;
  assign N180 = N114 & r_addr_r[6];
  assign N181 = N116 & N148;
  assign N182 = N116 & r_addr_r[6];
  assign N183 = N118 & N148;
  assign N184 = N118 & r_addr_r[6];
  assign N185 = N120 & N148;
  assign N186 = N120 & r_addr_r[6];
  assign N187 = N122 & N148;
  assign N188 = N122 & r_addr_r[6];
  assign N189 = N124 & N148;
  assign N190 = N124 & r_addr_r[6];
  assign N191 = N126 & N148;
  assign N192 = N126 & r_addr_r[6];
  assign N193 = N128 & N148;
  assign N194 = N128 & r_addr_r[6];
  assign N195 = N130 & N148;
  assign N196 = N130 & r_addr_r[6];
  assign N197 = N132 & N148;
  assign N198 = N132 & r_addr_r[6];
  assign N199 = N134 & N148;
  assign N200 = N134 & r_addr_r[6];
  assign N201 = N136 & N148;
  assign N202 = N136 & r_addr_r[6];
  assign N203 = N138 & N148;
  assign N204 = N138 & r_addr_r[6];
  assign N205 = N140 & N148;
  assign N206 = N140 & r_addr_r[6];
  assign N207 = N142 & N148;
  assign N208 = N142 & r_addr_r[6];
  assign N209 = N144 & N148;
  assign N210 = N144 & r_addr_r[6];
  assign N211 = N146 & N148;
  assign N212 = N146 & r_addr_r[6];
  assign N213 = N85 & N148;
  assign N214 = N85 & r_addr_r[6];
  assign N215 = N87 & N148;
  assign N216 = N87 & r_addr_r[6];
  assign N217 = N89 & N148;
  assign N218 = N89 & r_addr_r[6];
  assign N219 = N91 & N148;
  assign N220 = N91 & r_addr_r[6];
  assign N221 = N93 & N148;
  assign N222 = N93 & r_addr_r[6];
  assign N223 = N95 & N148;
  assign N224 = N95 & r_addr_r[6];
  assign N225 = N97 & N148;
  assign N226 = N97 & r_addr_r[6];
  assign N227 = N99 & N148;
  assign N228 = N99 & r_addr_r[6];
  assign N229 = N101 & N148;
  assign N230 = N101 & r_addr_r[6];
  assign N231 = N103 & N148;
  assign N232 = N103 & r_addr_r[6];
  assign N233 = N105 & N148;
  assign N234 = N105 & r_addr_r[6];
  assign N235 = N107 & N148;
  assign N236 = N107 & r_addr_r[6];
  assign N237 = N109 & N148;
  assign N238 = N109 & r_addr_r[6];
  assign N239 = N111 & N148;
  assign N240 = N111 & r_addr_r[6];
  assign N241 = N113 & N148;
  assign N242 = N113 & r_addr_r[6];
  assign N243 = N115 & N148;
  assign N244 = N115 & r_addr_r[6];
  assign N245 = N117 & N148;
  assign N246 = N117 & r_addr_r[6];
  assign N247 = N119 & N148;
  assign N248 = N119 & r_addr_r[6];
  assign N249 = N121 & N148;
  assign N250 = N121 & r_addr_r[6];
  assign N251 = N123 & N148;
  assign N252 = N123 & r_addr_r[6];
  assign N253 = N125 & N148;
  assign N254 = N125 & r_addr_r[6];
  assign N255 = N127 & N148;
  assign N256 = N127 & r_addr_r[6];
  assign N257 = N129 & N148;
  assign N258 = N129 & r_addr_r[6];
  assign N259 = N131 & N148;
  assign N260 = N131 & r_addr_r[6];
  assign N261 = N133 & N148;
  assign N262 = N133 & r_addr_r[6];
  assign N263 = N135 & N148;
  assign N264 = N135 & r_addr_r[6];
  assign N265 = N137 & N148;
  assign N266 = N137 & r_addr_r[6];
  assign N267 = N139 & N148;
  assign N268 = N139 & r_addr_r[6];
  assign N269 = N141 & N148;
  assign N270 = N141 & r_addr_r[6];
  assign N271 = N143 & N148;
  assign N272 = N143 & r_addr_r[6];
  assign N273 = N145 & N148;
  assign N274 = N145 & r_addr_r[6];
  assign N275 = N147 & N148;
  assign N276 = N147 & r_addr_r[6];
  assign N277 = ~r_addr_r[7];
  assign N278 = N149 & N277;
  assign N279 = N149 & r_addr_r[7];
  assign N280 = N151 & N277;
  assign N281 = N151 & r_addr_r[7];
  assign N282 = N153 & N277;
  assign N283 = N153 & r_addr_r[7];
  assign N284 = N155 & N277;
  assign N285 = N155 & r_addr_r[7];
  assign N286 = N157 & N277;
  assign N287 = N157 & r_addr_r[7];
  assign N288 = N159 & N277;
  assign N289 = N159 & r_addr_r[7];
  assign N290 = N161 & N277;
  assign N291 = N161 & r_addr_r[7];
  assign N292 = N163 & N277;
  assign N293 = N163 & r_addr_r[7];
  assign N294 = N165 & N277;
  assign N295 = N165 & r_addr_r[7];
  assign N296 = N167 & N277;
  assign N297 = N167 & r_addr_r[7];
  assign N298 = N169 & N277;
  assign N299 = N169 & r_addr_r[7];
  assign N300 = N171 & N277;
  assign N301 = N171 & r_addr_r[7];
  assign N302 = N173 & N277;
  assign N303 = N173 & r_addr_r[7];
  assign N304 = N175 & N277;
  assign N305 = N175 & r_addr_r[7];
  assign N306 = N177 & N277;
  assign N307 = N177 & r_addr_r[7];
  assign N308 = N179 & N277;
  assign N309 = N179 & r_addr_r[7];
  assign N310 = N181 & N277;
  assign N311 = N181 & r_addr_r[7];
  assign N312 = N183 & N277;
  assign N313 = N183 & r_addr_r[7];
  assign N314 = N185 & N277;
  assign N315 = N185 & r_addr_r[7];
  assign N316 = N187 & N277;
  assign N317 = N187 & r_addr_r[7];
  assign N318 = N189 & N277;
  assign N319 = N189 & r_addr_r[7];
  assign N320 = N191 & N277;
  assign N321 = N191 & r_addr_r[7];
  assign N322 = N193 & N277;
  assign N323 = N193 & r_addr_r[7];
  assign N324 = N195 & N277;
  assign N325 = N195 & r_addr_r[7];
  assign N326 = N197 & N277;
  assign N327 = N197 & r_addr_r[7];
  assign N328 = N199 & N277;
  assign N329 = N199 & r_addr_r[7];
  assign N330 = N201 & N277;
  assign N331 = N201 & r_addr_r[7];
  assign N332 = N203 & N277;
  assign N333 = N203 & r_addr_r[7];
  assign N334 = N205 & N277;
  assign N335 = N205 & r_addr_r[7];
  assign N336 = N207 & N277;
  assign N337 = N207 & r_addr_r[7];
  assign N338 = N209 & N277;
  assign N339 = N209 & r_addr_r[7];
  assign N340 = N211 & N277;
  assign N341 = N211 & r_addr_r[7];
  assign N342 = N213 & N277;
  assign N343 = N213 & r_addr_r[7];
  assign N344 = N215 & N277;
  assign N345 = N215 & r_addr_r[7];
  assign N346 = N217 & N277;
  assign N347 = N217 & r_addr_r[7];
  assign N348 = N219 & N277;
  assign N349 = N219 & r_addr_r[7];
  assign N350 = N221 & N277;
  assign N351 = N221 & r_addr_r[7];
  assign N352 = N223 & N277;
  assign N353 = N223 & r_addr_r[7];
  assign N354 = N225 & N277;
  assign N355 = N225 & r_addr_r[7];
  assign N356 = N227 & N277;
  assign N357 = N227 & r_addr_r[7];
  assign N358 = N229 & N277;
  assign N359 = N229 & r_addr_r[7];
  assign N360 = N231 & N277;
  assign N361 = N231 & r_addr_r[7];
  assign N362 = N233 & N277;
  assign N363 = N233 & r_addr_r[7];
  assign N364 = N235 & N277;
  assign N365 = N235 & r_addr_r[7];
  assign N366 = N237 & N277;
  assign N367 = N237 & r_addr_r[7];
  assign N368 = N239 & N277;
  assign N369 = N239 & r_addr_r[7];
  assign N370 = N241 & N277;
  assign N371 = N241 & r_addr_r[7];
  assign N372 = N243 & N277;
  assign N373 = N243 & r_addr_r[7];
  assign N374 = N245 & N277;
  assign N375 = N245 & r_addr_r[7];
  assign N376 = N247 & N277;
  assign N377 = N247 & r_addr_r[7];
  assign N378 = N249 & N277;
  assign N379 = N249 & r_addr_r[7];
  assign N380 = N251 & N277;
  assign N381 = N251 & r_addr_r[7];
  assign N382 = N253 & N277;
  assign N383 = N253 & r_addr_r[7];
  assign N384 = N255 & N277;
  assign N385 = N255 & r_addr_r[7];
  assign N386 = N257 & N277;
  assign N387 = N257 & r_addr_r[7];
  assign N388 = N259 & N277;
  assign N389 = N259 & r_addr_r[7];
  assign N390 = N261 & N277;
  assign N391 = N261 & r_addr_r[7];
  assign N392 = N263 & N277;
  assign N393 = N263 & r_addr_r[7];
  assign N394 = N265 & N277;
  assign N395 = N265 & r_addr_r[7];
  assign N396 = N267 & N277;
  assign N397 = N267 & r_addr_r[7];
  assign N398 = N269 & N277;
  assign N399 = N269 & r_addr_r[7];
  assign N400 = N271 & N277;
  assign N401 = N271 & r_addr_r[7];
  assign N402 = N273 & N277;
  assign N403 = N273 & r_addr_r[7];
  assign N404 = N275 & N277;
  assign N405 = N275 & r_addr_r[7];
  assign N406 = N150 & N277;
  assign N407 = N150 & r_addr_r[7];
  assign N408 = N152 & N277;
  assign N409 = N152 & r_addr_r[7];
  assign N410 = N154 & N277;
  assign N411 = N154 & r_addr_r[7];
  assign N412 = N156 & N277;
  assign N413 = N156 & r_addr_r[7];
  assign N414 = N158 & N277;
  assign N415 = N158 & r_addr_r[7];
  assign N416 = N160 & N277;
  assign N417 = N160 & r_addr_r[7];
  assign N418 = N162 & N277;
  assign N419 = N162 & r_addr_r[7];
  assign N420 = N164 & N277;
  assign N421 = N164 & r_addr_r[7];
  assign N422 = N166 & N277;
  assign N423 = N166 & r_addr_r[7];
  assign N424 = N168 & N277;
  assign N425 = N168 & r_addr_r[7];
  assign N426 = N170 & N277;
  assign N427 = N170 & r_addr_r[7];
  assign N428 = N172 & N277;
  assign N429 = N172 & r_addr_r[7];
  assign N430 = N174 & N277;
  assign N431 = N174 & r_addr_r[7];
  assign N432 = N176 & N277;
  assign N433 = N176 & r_addr_r[7];
  assign N434 = N178 & N277;
  assign N435 = N178 & r_addr_r[7];
  assign N436 = N180 & N277;
  assign N437 = N180 & r_addr_r[7];
  assign N438 = N182 & N277;
  assign N439 = N182 & r_addr_r[7];
  assign N440 = N184 & N277;
  assign N441 = N184 & r_addr_r[7];
  assign N442 = N186 & N277;
  assign N443 = N186 & r_addr_r[7];
  assign N444 = N188 & N277;
  assign N445 = N188 & r_addr_r[7];
  assign N446 = N190 & N277;
  assign N447 = N190 & r_addr_r[7];
  assign N448 = N192 & N277;
  assign N449 = N192 & r_addr_r[7];
  assign N450 = N194 & N277;
  assign N451 = N194 & r_addr_r[7];
  assign N452 = N196 & N277;
  assign N453 = N196 & r_addr_r[7];
  assign N454 = N198 & N277;
  assign N455 = N198 & r_addr_r[7];
  assign N456 = N200 & N277;
  assign N457 = N200 & r_addr_r[7];
  assign N458 = N202 & N277;
  assign N459 = N202 & r_addr_r[7];
  assign N460 = N204 & N277;
  assign N461 = N204 & r_addr_r[7];
  assign N462 = N206 & N277;
  assign N463 = N206 & r_addr_r[7];
  assign N464 = N208 & N277;
  assign N465 = N208 & r_addr_r[7];
  assign N466 = N210 & N277;
  assign N467 = N210 & r_addr_r[7];
  assign N468 = N212 & N277;
  assign N469 = N212 & r_addr_r[7];
  assign N470 = N214 & N277;
  assign N471 = N214 & r_addr_r[7];
  assign N472 = N216 & N277;
  assign N473 = N216 & r_addr_r[7];
  assign N474 = N218 & N277;
  assign N475 = N218 & r_addr_r[7];
  assign N476 = N220 & N277;
  assign N477 = N220 & r_addr_r[7];
  assign N478 = N222 & N277;
  assign N479 = N222 & r_addr_r[7];
  assign N480 = N224 & N277;
  assign N481 = N224 & r_addr_r[7];
  assign N482 = N226 & N277;
  assign N483 = N226 & r_addr_r[7];
  assign N484 = N228 & N277;
  assign N485 = N228 & r_addr_r[7];
  assign N486 = N230 & N277;
  assign N487 = N230 & r_addr_r[7];
  assign N488 = N232 & N277;
  assign N489 = N232 & r_addr_r[7];
  assign N490 = N234 & N277;
  assign N491 = N234 & r_addr_r[7];
  assign N492 = N236 & N277;
  assign N493 = N236 & r_addr_r[7];
  assign N494 = N238 & N277;
  assign N495 = N238 & r_addr_r[7];
  assign N496 = N240 & N277;
  assign N497 = N240 & r_addr_r[7];
  assign N498 = N242 & N277;
  assign N499 = N242 & r_addr_r[7];
  assign N500 = N244 & N277;
  assign N501 = N244 & r_addr_r[7];
  assign N502 = N246 & N277;
  assign N503 = N246 & r_addr_r[7];
  assign N504 = N248 & N277;
  assign N505 = N248 & r_addr_r[7];
  assign N506 = N250 & N277;
  assign N507 = N250 & r_addr_r[7];
  assign N508 = N252 & N277;
  assign N509 = N252 & r_addr_r[7];
  assign N510 = N254 & N277;
  assign N511 = N254 & r_addr_r[7];
  assign N512 = N256 & N277;
  assign N513 = N256 & r_addr_r[7];
  assign N514 = N258 & N277;
  assign N515 = N258 & r_addr_r[7];
  assign N516 = N260 & N277;
  assign N517 = N260 & r_addr_r[7];
  assign N518 = N262 & N277;
  assign N519 = N262 & r_addr_r[7];
  assign N520 = N264 & N277;
  assign N521 = N264 & r_addr_r[7];
  assign N522 = N266 & N277;
  assign N523 = N266 & r_addr_r[7];
  assign N524 = N268 & N277;
  assign N525 = N268 & r_addr_r[7];
  assign N526 = N270 & N277;
  assign N527 = N270 & r_addr_r[7];
  assign N528 = N272 & N277;
  assign N529 = N272 & r_addr_r[7];
  assign N530 = N274 & N277;
  assign N531 = N274 & r_addr_r[7];
  assign N532 = N276 & N277;
  assign N533 = N276 & r_addr_r[7];
  assign N534 = ~r_addr_r[8];
  assign N535 = N278 & N534;
  assign N536 = N278 & r_addr_r[8];
  assign N537 = N280 & N534;
  assign N538 = N280 & r_addr_r[8];
  assign N539 = N282 & N534;
  assign N540 = N282 & r_addr_r[8];
  assign N541 = N284 & N534;
  assign N542 = N284 & r_addr_r[8];
  assign N543 = N286 & N534;
  assign N544 = N286 & r_addr_r[8];
  assign N545 = N288 & N534;
  assign N546 = N288 & r_addr_r[8];
  assign N547 = N290 & N534;
  assign N548 = N290 & r_addr_r[8];
  assign N549 = N292 & N534;
  assign N550 = N292 & r_addr_r[8];
  assign N551 = N294 & N534;
  assign N552 = N294 & r_addr_r[8];
  assign N553 = N296 & N534;
  assign N554 = N296 & r_addr_r[8];
  assign N555 = N298 & N534;
  assign N556 = N298 & r_addr_r[8];
  assign N557 = N300 & N534;
  assign N558 = N300 & r_addr_r[8];
  assign N559 = N302 & N534;
  assign N560 = N302 & r_addr_r[8];
  assign N561 = N304 & N534;
  assign N562 = N304 & r_addr_r[8];
  assign N563 = N306 & N534;
  assign N564 = N306 & r_addr_r[8];
  assign N565 = N308 & N534;
  assign N566 = N308 & r_addr_r[8];
  assign N567 = N310 & N534;
  assign N568 = N310 & r_addr_r[8];
  assign N569 = N312 & N534;
  assign N570 = N312 & r_addr_r[8];
  assign N571 = N314 & N534;
  assign N572 = N314 & r_addr_r[8];
  assign N573 = N316 & N534;
  assign N574 = N316 & r_addr_r[8];
  assign N575 = N318 & N534;
  assign N576 = N318 & r_addr_r[8];
  assign N577 = N320 & N534;
  assign N578 = N320 & r_addr_r[8];
  assign N579 = N322 & N534;
  assign N580 = N322 & r_addr_r[8];
  assign N581 = N324 & N534;
  assign N582 = N324 & r_addr_r[8];
  assign N583 = N326 & N534;
  assign N584 = N326 & r_addr_r[8];
  assign N585 = N328 & N534;
  assign N586 = N328 & r_addr_r[8];
  assign N587 = N330 & N534;
  assign N588 = N330 & r_addr_r[8];
  assign N589 = N332 & N534;
  assign N590 = N332 & r_addr_r[8];
  assign N591 = N334 & N534;
  assign N592 = N334 & r_addr_r[8];
  assign N593 = N336 & N534;
  assign N594 = N336 & r_addr_r[8];
  assign N595 = N338 & N534;
  assign N596 = N338 & r_addr_r[8];
  assign N597 = N340 & N534;
  assign N598 = N340 & r_addr_r[8];
  assign N599 = N342 & N534;
  assign N600 = N342 & r_addr_r[8];
  assign N601 = N344 & N534;
  assign N602 = N344 & r_addr_r[8];
  assign N603 = N346 & N534;
  assign N604 = N346 & r_addr_r[8];
  assign N605 = N348 & N534;
  assign N606 = N348 & r_addr_r[8];
  assign N607 = N350 & N534;
  assign N608 = N350 & r_addr_r[8];
  assign N609 = N352 & N534;
  assign N610 = N352 & r_addr_r[8];
  assign N611 = N354 & N534;
  assign N612 = N354 & r_addr_r[8];
  assign N613 = N356 & N534;
  assign N614 = N356 & r_addr_r[8];
  assign N615 = N358 & N534;
  assign N616 = N358 & r_addr_r[8];
  assign N617 = N360 & N534;
  assign N618 = N360 & r_addr_r[8];
  assign N619 = N362 & N534;
  assign N620 = N362 & r_addr_r[8];
  assign N621 = N364 & N534;
  assign N622 = N364 & r_addr_r[8];
  assign N623 = N366 & N534;
  assign N624 = N366 & r_addr_r[8];
  assign N625 = N368 & N534;
  assign N626 = N368 & r_addr_r[8];
  assign N627 = N370 & N534;
  assign N628 = N370 & r_addr_r[8];
  assign N629 = N372 & N534;
  assign N630 = N372 & r_addr_r[8];
  assign N631 = N374 & N534;
  assign N632 = N374 & r_addr_r[8];
  assign N633 = N376 & N534;
  assign N634 = N376 & r_addr_r[8];
  assign N635 = N378 & N534;
  assign N636 = N378 & r_addr_r[8];
  assign N637 = N380 & N534;
  assign N638 = N380 & r_addr_r[8];
  assign N639 = N382 & N534;
  assign N640 = N382 & r_addr_r[8];
  assign N641 = N384 & N534;
  assign N642 = N384 & r_addr_r[8];
  assign N643 = N386 & N534;
  assign N644 = N386 & r_addr_r[8];
  assign N645 = N388 & N534;
  assign N646 = N388 & r_addr_r[8];
  assign N647 = N390 & N534;
  assign N648 = N390 & r_addr_r[8];
  assign N649 = N392 & N534;
  assign N650 = N392 & r_addr_r[8];
  assign N651 = N394 & N534;
  assign N652 = N394 & r_addr_r[8];
  assign N653 = N396 & N534;
  assign N654 = N396 & r_addr_r[8];
  assign N655 = N398 & N534;
  assign N656 = N398 & r_addr_r[8];
  assign N657 = N400 & N534;
  assign N658 = N400 & r_addr_r[8];
  assign N659 = N402 & N534;
  assign N660 = N402 & r_addr_r[8];
  assign N661 = N404 & N534;
  assign N662 = N404 & r_addr_r[8];
  assign N663 = N406 & N534;
  assign N664 = N406 & r_addr_r[8];
  assign N665 = N408 & N534;
  assign N666 = N408 & r_addr_r[8];
  assign N667 = N410 & N534;
  assign N668 = N410 & r_addr_r[8];
  assign N669 = N412 & N534;
  assign N670 = N412 & r_addr_r[8];
  assign N671 = N414 & N534;
  assign N672 = N414 & r_addr_r[8];
  assign N673 = N416 & N534;
  assign N674 = N416 & r_addr_r[8];
  assign N675 = N418 & N534;
  assign N676 = N418 & r_addr_r[8];
  assign N677 = N420 & N534;
  assign N678 = N420 & r_addr_r[8];
  assign N679 = N422 & N534;
  assign N680 = N422 & r_addr_r[8];
  assign N681 = N424 & N534;
  assign N682 = N424 & r_addr_r[8];
  assign N683 = N426 & N534;
  assign N684 = N426 & r_addr_r[8];
  assign N685 = N428 & N534;
  assign N686 = N428 & r_addr_r[8];
  assign N687 = N430 & N534;
  assign N688 = N430 & r_addr_r[8];
  assign N689 = N432 & N534;
  assign N690 = N432 & r_addr_r[8];
  assign N691 = N434 & N534;
  assign N692 = N434 & r_addr_r[8];
  assign N693 = N436 & N534;
  assign N694 = N436 & r_addr_r[8];
  assign N695 = N438 & N534;
  assign N696 = N438 & r_addr_r[8];
  assign N697 = N440 & N534;
  assign N698 = N440 & r_addr_r[8];
  assign N699 = N442 & N534;
  assign N700 = N442 & r_addr_r[8];
  assign N701 = N444 & N534;
  assign N702 = N444 & r_addr_r[8];
  assign N703 = N446 & N534;
  assign N704 = N446 & r_addr_r[8];
  assign N705 = N448 & N534;
  assign N706 = N448 & r_addr_r[8];
  assign N707 = N450 & N534;
  assign N708 = N450 & r_addr_r[8];
  assign N709 = N452 & N534;
  assign N710 = N452 & r_addr_r[8];
  assign N711 = N454 & N534;
  assign N712 = N454 & r_addr_r[8];
  assign N713 = N456 & N534;
  assign N714 = N456 & r_addr_r[8];
  assign N715 = N458 & N534;
  assign N716 = N458 & r_addr_r[8];
  assign N717 = N460 & N534;
  assign N718 = N460 & r_addr_r[8];
  assign N719 = N462 & N534;
  assign N720 = N462 & r_addr_r[8];
  assign N721 = N464 & N534;
  assign N722 = N464 & r_addr_r[8];
  assign N723 = N466 & N534;
  assign N724 = N466 & r_addr_r[8];
  assign N725 = N468 & N534;
  assign N726 = N468 & r_addr_r[8];
  assign N727 = N470 & N534;
  assign N728 = N470 & r_addr_r[8];
  assign N729 = N472 & N534;
  assign N730 = N472 & r_addr_r[8];
  assign N731 = N474 & N534;
  assign N732 = N474 & r_addr_r[8];
  assign N733 = N476 & N534;
  assign N734 = N476 & r_addr_r[8];
  assign N735 = N478 & N534;
  assign N736 = N478 & r_addr_r[8];
  assign N737 = N480 & N534;
  assign N738 = N480 & r_addr_r[8];
  assign N739 = N482 & N534;
  assign N740 = N482 & r_addr_r[8];
  assign N741 = N484 & N534;
  assign N742 = N484 & r_addr_r[8];
  assign N743 = N486 & N534;
  assign N744 = N486 & r_addr_r[8];
  assign N745 = N488 & N534;
  assign N746 = N488 & r_addr_r[8];
  assign N747 = N490 & N534;
  assign N748 = N490 & r_addr_r[8];
  assign N749 = N492 & N534;
  assign N750 = N492 & r_addr_r[8];
  assign N751 = N494 & N534;
  assign N752 = N494 & r_addr_r[8];
  assign N753 = N496 & N534;
  assign N754 = N496 & r_addr_r[8];
  assign N755 = N498 & N534;
  assign N756 = N498 & r_addr_r[8];
  assign N757 = N500 & N534;
  assign N758 = N500 & r_addr_r[8];
  assign N759 = N502 & N534;
  assign N760 = N502 & r_addr_r[8];
  assign N761 = N504 & N534;
  assign N762 = N504 & r_addr_r[8];
  assign N763 = N506 & N534;
  assign N764 = N506 & r_addr_r[8];
  assign N765 = N508 & N534;
  assign N766 = N508 & r_addr_r[8];
  assign N767 = N510 & N534;
  assign N768 = N510 & r_addr_r[8];
  assign N769 = N512 & N534;
  assign N770 = N512 & r_addr_r[8];
  assign N771 = N514 & N534;
  assign N772 = N514 & r_addr_r[8];
  assign N773 = N516 & N534;
  assign N774 = N516 & r_addr_r[8];
  assign N775 = N518 & N534;
  assign N776 = N518 & r_addr_r[8];
  assign N777 = N520 & N534;
  assign N778 = N520 & r_addr_r[8];
  assign N779 = N522 & N534;
  assign N780 = N522 & r_addr_r[8];
  assign N781 = N524 & N534;
  assign N782 = N524 & r_addr_r[8];
  assign N783 = N526 & N534;
  assign N784 = N526 & r_addr_r[8];
  assign N785 = N528 & N534;
  assign N786 = N528 & r_addr_r[8];
  assign N787 = N530 & N534;
  assign N788 = N530 & r_addr_r[8];
  assign N789 = N532 & N534;
  assign N790 = N532 & r_addr_r[8];
  assign N791 = N279 & N534;
  assign N792 = N279 & r_addr_r[8];
  assign N793 = N281 & N534;
  assign N794 = N281 & r_addr_r[8];
  assign N795 = N283 & N534;
  assign N796 = N283 & r_addr_r[8];
  assign N797 = N285 & N534;
  assign N798 = N285 & r_addr_r[8];
  assign N799 = N287 & N534;
  assign N800 = N287 & r_addr_r[8];
  assign N801 = N289 & N534;
  assign N802 = N289 & r_addr_r[8];
  assign N803 = N291 & N534;
  assign N804 = N291 & r_addr_r[8];
  assign N805 = N293 & N534;
  assign N806 = N293 & r_addr_r[8];
  assign N807 = N295 & N534;
  assign N808 = N295 & r_addr_r[8];
  assign N809 = N297 & N534;
  assign N810 = N297 & r_addr_r[8];
  assign N811 = N299 & N534;
  assign N812 = N299 & r_addr_r[8];
  assign N813 = N301 & N534;
  assign N814 = N301 & r_addr_r[8];
  assign N815 = N303 & N534;
  assign N816 = N303 & r_addr_r[8];
  assign N817 = N305 & N534;
  assign N818 = N305 & r_addr_r[8];
  assign N819 = N307 & N534;
  assign N820 = N307 & r_addr_r[8];
  assign N821 = N309 & N534;
  assign N822 = N309 & r_addr_r[8];
  assign N823 = N311 & N534;
  assign N824 = N311 & r_addr_r[8];
  assign N825 = N313 & N534;
  assign N826 = N313 & r_addr_r[8];
  assign N827 = N315 & N534;
  assign N828 = N315 & r_addr_r[8];
  assign N829 = N317 & N534;
  assign N830 = N317 & r_addr_r[8];
  assign N831 = N319 & N534;
  assign N832 = N319 & r_addr_r[8];
  assign N833 = N321 & N534;
  assign N834 = N321 & r_addr_r[8];
  assign N835 = N323 & N534;
  assign N836 = N323 & r_addr_r[8];
  assign N837 = N325 & N534;
  assign N838 = N325 & r_addr_r[8];
  assign N839 = N327 & N534;
  assign N840 = N327 & r_addr_r[8];
  assign N841 = N329 & N534;
  assign N842 = N329 & r_addr_r[8];
  assign N843 = N331 & N534;
  assign N844 = N331 & r_addr_r[8];
  assign N845 = N333 & N534;
  assign N846 = N333 & r_addr_r[8];
  assign N847 = N335 & N534;
  assign N848 = N335 & r_addr_r[8];
  assign N849 = N337 & N534;
  assign N850 = N337 & r_addr_r[8];
  assign N851 = N339 & N534;
  assign N852 = N339 & r_addr_r[8];
  assign N853 = N341 & N534;
  assign N854 = N341 & r_addr_r[8];
  assign N855 = N343 & N534;
  assign N856 = N343 & r_addr_r[8];
  assign N857 = N345 & N534;
  assign N858 = N345 & r_addr_r[8];
  assign N859 = N347 & N534;
  assign N860 = N347 & r_addr_r[8];
  assign N861 = N349 & N534;
  assign N862 = N349 & r_addr_r[8];
  assign N863 = N351 & N534;
  assign N864 = N351 & r_addr_r[8];
  assign N865 = N353 & N534;
  assign N866 = N353 & r_addr_r[8];
  assign N867 = N355 & N534;
  assign N868 = N355 & r_addr_r[8];
  assign N869 = N357 & N534;
  assign N870 = N357 & r_addr_r[8];
  assign N871 = N359 & N534;
  assign N872 = N359 & r_addr_r[8];
  assign N873 = N361 & N534;
  assign N874 = N361 & r_addr_r[8];
  assign N875 = N363 & N534;
  assign N876 = N363 & r_addr_r[8];
  assign N877 = N365 & N534;
  assign N878 = N365 & r_addr_r[8];
  assign N879 = N367 & N534;
  assign N880 = N367 & r_addr_r[8];
  assign N881 = N369 & N534;
  assign N882 = N369 & r_addr_r[8];
  assign N883 = N371 & N534;
  assign N884 = N371 & r_addr_r[8];
  assign N885 = N373 & N534;
  assign N886 = N373 & r_addr_r[8];
  assign N887 = N375 & N534;
  assign N888 = N375 & r_addr_r[8];
  assign N889 = N377 & N534;
  assign N890 = N377 & r_addr_r[8];
  assign N891 = N379 & N534;
  assign N892 = N379 & r_addr_r[8];
  assign N893 = N381 & N534;
  assign N894 = N381 & r_addr_r[8];
  assign N895 = N383 & N534;
  assign N896 = N383 & r_addr_r[8];
  assign N897 = N385 & N534;
  assign N898 = N385 & r_addr_r[8];
  assign N899 = N387 & N534;
  assign N900 = N387 & r_addr_r[8];
  assign N901 = N389 & N534;
  assign N902 = N389 & r_addr_r[8];
  assign N903 = N391 & N534;
  assign N904 = N391 & r_addr_r[8];
  assign N905 = N393 & N534;
  assign N906 = N393 & r_addr_r[8];
  assign N907 = N395 & N534;
  assign N908 = N395 & r_addr_r[8];
  assign N909 = N397 & N534;
  assign N910 = N397 & r_addr_r[8];
  assign N911 = N399 & N534;
  assign N912 = N399 & r_addr_r[8];
  assign N913 = N401 & N534;
  assign N914 = N401 & r_addr_r[8];
  assign N915 = N403 & N534;
  assign N916 = N403 & r_addr_r[8];
  assign N917 = N405 & N534;
  assign N918 = N405 & r_addr_r[8];
  assign N919 = N407 & N534;
  assign N920 = N407 & r_addr_r[8];
  assign N921 = N409 & N534;
  assign N922 = N409 & r_addr_r[8];
  assign N923 = N411 & N534;
  assign N924 = N411 & r_addr_r[8];
  assign N925 = N413 & N534;
  assign N926 = N413 & r_addr_r[8];
  assign N927 = N415 & N534;
  assign N928 = N415 & r_addr_r[8];
  assign N929 = N417 & N534;
  assign N930 = N417 & r_addr_r[8];
  assign N931 = N419 & N534;
  assign N932 = N419 & r_addr_r[8];
  assign N933 = N421 & N534;
  assign N934 = N421 & r_addr_r[8];
  assign N935 = N423 & N534;
  assign N936 = N423 & r_addr_r[8];
  assign N937 = N425 & N534;
  assign N938 = N425 & r_addr_r[8];
  assign N939 = N427 & N534;
  assign N940 = N427 & r_addr_r[8];
  assign N941 = N429 & N534;
  assign N942 = N429 & r_addr_r[8];
  assign N943 = N431 & N534;
  assign N944 = N431 & r_addr_r[8];
  assign N945 = N433 & N534;
  assign N946 = N433 & r_addr_r[8];
  assign N947 = N435 & N534;
  assign N948 = N435 & r_addr_r[8];
  assign N949 = N437 & N534;
  assign N950 = N437 & r_addr_r[8];
  assign N951 = N439 & N534;
  assign N952 = N439 & r_addr_r[8];
  assign N953 = N441 & N534;
  assign N954 = N441 & r_addr_r[8];
  assign N955 = N443 & N534;
  assign N956 = N443 & r_addr_r[8];
  assign N957 = N445 & N534;
  assign N958 = N445 & r_addr_r[8];
  assign N959 = N447 & N534;
  assign N960 = N447 & r_addr_r[8];
  assign N961 = N449 & N534;
  assign N962 = N449 & r_addr_r[8];
  assign N963 = N451 & N534;
  assign N964 = N451 & r_addr_r[8];
  assign N965 = N453 & N534;
  assign N966 = N453 & r_addr_r[8];
  assign N967 = N455 & N534;
  assign N968 = N455 & r_addr_r[8];
  assign N969 = N457 & N534;
  assign N970 = N457 & r_addr_r[8];
  assign N971 = N459 & N534;
  assign N972 = N459 & r_addr_r[8];
  assign N973 = N461 & N534;
  assign N974 = N461 & r_addr_r[8];
  assign N975 = N463 & N534;
  assign N976 = N463 & r_addr_r[8];
  assign N977 = N465 & N534;
  assign N978 = N465 & r_addr_r[8];
  assign N979 = N467 & N534;
  assign N980 = N467 & r_addr_r[8];
  assign N981 = N469 & N534;
  assign N982 = N469 & r_addr_r[8];
  assign N983 = N471 & N534;
  assign N984 = N471 & r_addr_r[8];
  assign N985 = N473 & N534;
  assign N986 = N473 & r_addr_r[8];
  assign N987 = N475 & N534;
  assign N988 = N475 & r_addr_r[8];
  assign N989 = N477 & N534;
  assign N990 = N477 & r_addr_r[8];
  assign N991 = N479 & N534;
  assign N992 = N479 & r_addr_r[8];
  assign N993 = N481 & N534;
  assign N994 = N481 & r_addr_r[8];
  assign N995 = N483 & N534;
  assign N996 = N483 & r_addr_r[8];
  assign N997 = N485 & N534;
  assign N998 = N485 & r_addr_r[8];
  assign N999 = N487 & N534;
  assign N1000 = N487 & r_addr_r[8];
  assign N1001 = N489 & N534;
  assign N1002 = N489 & r_addr_r[8];
  assign N1003 = N491 & N534;
  assign N1004 = N491 & r_addr_r[8];
  assign N1005 = N493 & N534;
  assign N1006 = N493 & r_addr_r[8];
  assign N1007 = N495 & N534;
  assign N1008 = N495 & r_addr_r[8];
  assign N1009 = N497 & N534;
  assign N1010 = N497 & r_addr_r[8];
  assign N1011 = N499 & N534;
  assign N1012 = N499 & r_addr_r[8];
  assign N1013 = N501 & N534;
  assign N1014 = N501 & r_addr_r[8];
  assign N1015 = N503 & N534;
  assign N1016 = N503 & r_addr_r[8];
  assign N1017 = N505 & N534;
  assign N1018 = N505 & r_addr_r[8];
  assign N1019 = N507 & N534;
  assign N1020 = N507 & r_addr_r[8];
  assign N1021 = N509 & N534;
  assign N1022 = N509 & r_addr_r[8];
  assign N1023 = N511 & N534;
  assign N1024 = N511 & r_addr_r[8];
  assign N1025 = N513 & N534;
  assign N1026 = N513 & r_addr_r[8];
  assign N1027 = N515 & N534;
  assign N1028 = N515 & r_addr_r[8];
  assign N1029 = N517 & N534;
  assign N1030 = N517 & r_addr_r[8];
  assign N1031 = N519 & N534;
  assign N1032 = N519 & r_addr_r[8];
  assign N1033 = N521 & N534;
  assign N1034 = N521 & r_addr_r[8];
  assign N1035 = N523 & N534;
  assign N1036 = N523 & r_addr_r[8];
  assign N1037 = N525 & N534;
  assign N1038 = N525 & r_addr_r[8];
  assign N1039 = N527 & N534;
  assign N1040 = N527 & r_addr_r[8];
  assign N1041 = N529 & N534;
  assign N1042 = N529 & r_addr_r[8];
  assign N1043 = N531 & N534;
  assign N1044 = N531 & r_addr_r[8];
  assign N1045 = N533 & N534;
  assign N1046 = N533 & r_addr_r[8];
  assign N1047 = ~w_v_i;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { r_addr_r[8:0] } <= { r_addr_i[8:0] };
    end 
    if(N2071) begin
      { mem[8191:8176] } <= { w_data_i[15:0] };
    end 
    if(N2070) begin
      { mem[8175:8160] } <= { w_data_i[15:0] };
    end 
    if(N2069) begin
      { mem[8159:8144] } <= { w_data_i[15:0] };
    end 
    if(N2068) begin
      { mem[8143:8128] } <= { w_data_i[15:0] };
    end 
    if(N2067) begin
      { mem[8127:8112] } <= { w_data_i[15:0] };
    end 
    if(N2066) begin
      { mem[8111:8096] } <= { w_data_i[15:0] };
    end 
    if(N2065) begin
      { mem[8095:8080] } <= { w_data_i[15:0] };
    end 
    if(N2064) begin
      { mem[8079:8064] } <= { w_data_i[15:0] };
    end 
    if(N2063) begin
      { mem[8063:8048] } <= { w_data_i[15:0] };
    end 
    if(N2062) begin
      { mem[8047:8032] } <= { w_data_i[15:0] };
    end 
    if(N2061) begin
      { mem[8031:8016] } <= { w_data_i[15:0] };
    end 
    if(N2060) begin
      { mem[8015:8000] } <= { w_data_i[15:0] };
    end 
    if(N2059) begin
      { mem[7999:7984] } <= { w_data_i[15:0] };
    end 
    if(N2058) begin
      { mem[7983:7968] } <= { w_data_i[15:0] };
    end 
    if(N2057) begin
      { mem[7967:7952] } <= { w_data_i[15:0] };
    end 
    if(N2056) begin
      { mem[7951:7936] } <= { w_data_i[15:0] };
    end 
    if(N2055) begin
      { mem[7935:7920] } <= { w_data_i[15:0] };
    end 
    if(N2054) begin
      { mem[7919:7904] } <= { w_data_i[15:0] };
    end 
    if(N2053) begin
      { mem[7903:7888] } <= { w_data_i[15:0] };
    end 
    if(N2052) begin
      { mem[7887:7872] } <= { w_data_i[15:0] };
    end 
    if(N2051) begin
      { mem[7871:7856] } <= { w_data_i[15:0] };
    end 
    if(N2050) begin
      { mem[7855:7840] } <= { w_data_i[15:0] };
    end 
    if(N2049) begin
      { mem[7839:7824] } <= { w_data_i[15:0] };
    end 
    if(N2048) begin
      { mem[7823:7808] } <= { w_data_i[15:0] };
    end 
    if(N2047) begin
      { mem[7807:7792] } <= { w_data_i[15:0] };
    end 
    if(N2046) begin
      { mem[7791:7776] } <= { w_data_i[15:0] };
    end 
    if(N2045) begin
      { mem[7775:7760] } <= { w_data_i[15:0] };
    end 
    if(N2044) begin
      { mem[7759:7744] } <= { w_data_i[15:0] };
    end 
    if(N2043) begin
      { mem[7743:7728] } <= { w_data_i[15:0] };
    end 
    if(N2042) begin
      { mem[7727:7712] } <= { w_data_i[15:0] };
    end 
    if(N2041) begin
      { mem[7711:7696] } <= { w_data_i[15:0] };
    end 
    if(N2040) begin
      { mem[7695:7680] } <= { w_data_i[15:0] };
    end 
    if(N2039) begin
      { mem[7679:7664] } <= { w_data_i[15:0] };
    end 
    if(N2038) begin
      { mem[7663:7648] } <= { w_data_i[15:0] };
    end 
    if(N2037) begin
      { mem[7647:7632] } <= { w_data_i[15:0] };
    end 
    if(N2036) begin
      { mem[7631:7616] } <= { w_data_i[15:0] };
    end 
    if(N2035) begin
      { mem[7615:7600] } <= { w_data_i[15:0] };
    end 
    if(N2034) begin
      { mem[7599:7584] } <= { w_data_i[15:0] };
    end 
    if(N2033) begin
      { mem[7583:7568] } <= { w_data_i[15:0] };
    end 
    if(N2032) begin
      { mem[7567:7552] } <= { w_data_i[15:0] };
    end 
    if(N2031) begin
      { mem[7551:7536] } <= { w_data_i[15:0] };
    end 
    if(N2030) begin
      { mem[7535:7520] } <= { w_data_i[15:0] };
    end 
    if(N2029) begin
      { mem[7519:7504] } <= { w_data_i[15:0] };
    end 
    if(N2028) begin
      { mem[7503:7488] } <= { w_data_i[15:0] };
    end 
    if(N2027) begin
      { mem[7487:7472] } <= { w_data_i[15:0] };
    end 
    if(N2026) begin
      { mem[7471:7456] } <= { w_data_i[15:0] };
    end 
    if(N2025) begin
      { mem[7455:7440] } <= { w_data_i[15:0] };
    end 
    if(N2024) begin
      { mem[7439:7424] } <= { w_data_i[15:0] };
    end 
    if(N2023) begin
      { mem[7423:7408] } <= { w_data_i[15:0] };
    end 
    if(N2022) begin
      { mem[7407:7392] } <= { w_data_i[15:0] };
    end 
    if(N2021) begin
      { mem[7391:7376] } <= { w_data_i[15:0] };
    end 
    if(N2020) begin
      { mem[7375:7360] } <= { w_data_i[15:0] };
    end 
    if(N2019) begin
      { mem[7359:7344] } <= { w_data_i[15:0] };
    end 
    if(N2018) begin
      { mem[7343:7328] } <= { w_data_i[15:0] };
    end 
    if(N2017) begin
      { mem[7327:7312] } <= { w_data_i[15:0] };
    end 
    if(N2016) begin
      { mem[7311:7296] } <= { w_data_i[15:0] };
    end 
    if(N2015) begin
      { mem[7295:7280] } <= { w_data_i[15:0] };
    end 
    if(N2014) begin
      { mem[7279:7264] } <= { w_data_i[15:0] };
    end 
    if(N2013) begin
      { mem[7263:7248] } <= { w_data_i[15:0] };
    end 
    if(N2012) begin
      { mem[7247:7232] } <= { w_data_i[15:0] };
    end 
    if(N2011) begin
      { mem[7231:7216] } <= { w_data_i[15:0] };
    end 
    if(N2010) begin
      { mem[7215:7200] } <= { w_data_i[15:0] };
    end 
    if(N2009) begin
      { mem[7199:7184] } <= { w_data_i[15:0] };
    end 
    if(N2008) begin
      { mem[7183:7168] } <= { w_data_i[15:0] };
    end 
    if(N2007) begin
      { mem[7167:7152] } <= { w_data_i[15:0] };
    end 
    if(N2006) begin
      { mem[7151:7136] } <= { w_data_i[15:0] };
    end 
    if(N2005) begin
      { mem[7135:7120] } <= { w_data_i[15:0] };
    end 
    if(N2004) begin
      { mem[7119:7104] } <= { w_data_i[15:0] };
    end 
    if(N2003) begin
      { mem[7103:7088] } <= { w_data_i[15:0] };
    end 
    if(N2002) begin
      { mem[7087:7072] } <= { w_data_i[15:0] };
    end 
    if(N2001) begin
      { mem[7071:7056] } <= { w_data_i[15:0] };
    end 
    if(N2000) begin
      { mem[7055:7040] } <= { w_data_i[15:0] };
    end 
    if(N1999) begin
      { mem[7039:7024] } <= { w_data_i[15:0] };
    end 
    if(N1998) begin
      { mem[7023:7008] } <= { w_data_i[15:0] };
    end 
    if(N1997) begin
      { mem[7007:6992] } <= { w_data_i[15:0] };
    end 
    if(N1996) begin
      { mem[6991:6976] } <= { w_data_i[15:0] };
    end 
    if(N1995) begin
      { mem[6975:6960] } <= { w_data_i[15:0] };
    end 
    if(N1994) begin
      { mem[6959:6944] } <= { w_data_i[15:0] };
    end 
    if(N1993) begin
      { mem[6943:6928] } <= { w_data_i[15:0] };
    end 
    if(N1992) begin
      { mem[6927:6912] } <= { w_data_i[15:0] };
    end 
    if(N1991) begin
      { mem[6911:6896] } <= { w_data_i[15:0] };
    end 
    if(N1990) begin
      { mem[6895:6880] } <= { w_data_i[15:0] };
    end 
    if(N1989) begin
      { mem[6879:6864] } <= { w_data_i[15:0] };
    end 
    if(N1988) begin
      { mem[6863:6848] } <= { w_data_i[15:0] };
    end 
    if(N1987) begin
      { mem[6847:6832] } <= { w_data_i[15:0] };
    end 
    if(N1986) begin
      { mem[6831:6816] } <= { w_data_i[15:0] };
    end 
    if(N1985) begin
      { mem[6815:6800] } <= { w_data_i[15:0] };
    end 
    if(N1984) begin
      { mem[6799:6784] } <= { w_data_i[15:0] };
    end 
    if(N1983) begin
      { mem[6783:6768] } <= { w_data_i[15:0] };
    end 
    if(N1982) begin
      { mem[6767:6752] } <= { w_data_i[15:0] };
    end 
    if(N1981) begin
      { mem[6751:6736] } <= { w_data_i[15:0] };
    end 
    if(N1980) begin
      { mem[6735:6720] } <= { w_data_i[15:0] };
    end 
    if(N1979) begin
      { mem[6719:6704] } <= { w_data_i[15:0] };
    end 
    if(N1978) begin
      { mem[6703:6688] } <= { w_data_i[15:0] };
    end 
    if(N1977) begin
      { mem[6687:6672] } <= { w_data_i[15:0] };
    end 
    if(N1976) begin
      { mem[6671:6656] } <= { w_data_i[15:0] };
    end 
    if(N1975) begin
      { mem[6655:6640] } <= { w_data_i[15:0] };
    end 
    if(N1974) begin
      { mem[6639:6624] } <= { w_data_i[15:0] };
    end 
    if(N1973) begin
      { mem[6623:6608] } <= { w_data_i[15:0] };
    end 
    if(N1972) begin
      { mem[6607:6592] } <= { w_data_i[15:0] };
    end 
    if(N1971) begin
      { mem[6591:6576] } <= { w_data_i[15:0] };
    end 
    if(N1970) begin
      { mem[6575:6560] } <= { w_data_i[15:0] };
    end 
    if(N1969) begin
      { mem[6559:6544] } <= { w_data_i[15:0] };
    end 
    if(N1968) begin
      { mem[6543:6528] } <= { w_data_i[15:0] };
    end 
    if(N1967) begin
      { mem[6527:6512] } <= { w_data_i[15:0] };
    end 
    if(N1966) begin
      { mem[6511:6496] } <= { w_data_i[15:0] };
    end 
    if(N1965) begin
      { mem[6495:6480] } <= { w_data_i[15:0] };
    end 
    if(N1964) begin
      { mem[6479:6464] } <= { w_data_i[15:0] };
    end 
    if(N1963) begin
      { mem[6463:6448] } <= { w_data_i[15:0] };
    end 
    if(N1962) begin
      { mem[6447:6432] } <= { w_data_i[15:0] };
    end 
    if(N1961) begin
      { mem[6431:6416] } <= { w_data_i[15:0] };
    end 
    if(N1960) begin
      { mem[6415:6400] } <= { w_data_i[15:0] };
    end 
    if(N1959) begin
      { mem[6399:6384] } <= { w_data_i[15:0] };
    end 
    if(N1958) begin
      { mem[6383:6368] } <= { w_data_i[15:0] };
    end 
    if(N1957) begin
      { mem[6367:6352] } <= { w_data_i[15:0] };
    end 
    if(N1956) begin
      { mem[6351:6336] } <= { w_data_i[15:0] };
    end 
    if(N1955) begin
      { mem[6335:6320] } <= { w_data_i[15:0] };
    end 
    if(N1954) begin
      { mem[6319:6304] } <= { w_data_i[15:0] };
    end 
    if(N1953) begin
      { mem[6303:6288] } <= { w_data_i[15:0] };
    end 
    if(N1952) begin
      { mem[6287:6272] } <= { w_data_i[15:0] };
    end 
    if(N1951) begin
      { mem[6271:6256] } <= { w_data_i[15:0] };
    end 
    if(N1950) begin
      { mem[6255:6240] } <= { w_data_i[15:0] };
    end 
    if(N1949) begin
      { mem[6239:6224] } <= { w_data_i[15:0] };
    end 
    if(N1948) begin
      { mem[6223:6208] } <= { w_data_i[15:0] };
    end 
    if(N1947) begin
      { mem[6207:6192] } <= { w_data_i[15:0] };
    end 
    if(N1946) begin
      { mem[6191:6176] } <= { w_data_i[15:0] };
    end 
    if(N1945) begin
      { mem[6175:6160] } <= { w_data_i[15:0] };
    end 
    if(N1944) begin
      { mem[6159:6144] } <= { w_data_i[15:0] };
    end 
    if(N1943) begin
      { mem[6143:6128] } <= { w_data_i[15:0] };
    end 
    if(N1942) begin
      { mem[6127:6112] } <= { w_data_i[15:0] };
    end 
    if(N1941) begin
      { mem[6111:6096] } <= { w_data_i[15:0] };
    end 
    if(N1940) begin
      { mem[6095:6080] } <= { w_data_i[15:0] };
    end 
    if(N1939) begin
      { mem[6079:6064] } <= { w_data_i[15:0] };
    end 
    if(N1938) begin
      { mem[6063:6048] } <= { w_data_i[15:0] };
    end 
    if(N1937) begin
      { mem[6047:6032] } <= { w_data_i[15:0] };
    end 
    if(N1936) begin
      { mem[6031:6016] } <= { w_data_i[15:0] };
    end 
    if(N1935) begin
      { mem[6015:6000] } <= { w_data_i[15:0] };
    end 
    if(N1934) begin
      { mem[5999:5984] } <= { w_data_i[15:0] };
    end 
    if(N1933) begin
      { mem[5983:5968] } <= { w_data_i[15:0] };
    end 
    if(N1932) begin
      { mem[5967:5952] } <= { w_data_i[15:0] };
    end 
    if(N1931) begin
      { mem[5951:5936] } <= { w_data_i[15:0] };
    end 
    if(N1930) begin
      { mem[5935:5920] } <= { w_data_i[15:0] };
    end 
    if(N1929) begin
      { mem[5919:5904] } <= { w_data_i[15:0] };
    end 
    if(N1928) begin
      { mem[5903:5888] } <= { w_data_i[15:0] };
    end 
    if(N1927) begin
      { mem[5887:5872] } <= { w_data_i[15:0] };
    end 
    if(N1926) begin
      { mem[5871:5856] } <= { w_data_i[15:0] };
    end 
    if(N1925) begin
      { mem[5855:5840] } <= { w_data_i[15:0] };
    end 
    if(N1924) begin
      { mem[5839:5824] } <= { w_data_i[15:0] };
    end 
    if(N1923) begin
      { mem[5823:5808] } <= { w_data_i[15:0] };
    end 
    if(N1922) begin
      { mem[5807:5792] } <= { w_data_i[15:0] };
    end 
    if(N1921) begin
      { mem[5791:5776] } <= { w_data_i[15:0] };
    end 
    if(N1920) begin
      { mem[5775:5760] } <= { w_data_i[15:0] };
    end 
    if(N1919) begin
      { mem[5759:5744] } <= { w_data_i[15:0] };
    end 
    if(N1918) begin
      { mem[5743:5728] } <= { w_data_i[15:0] };
    end 
    if(N1917) begin
      { mem[5727:5712] } <= { w_data_i[15:0] };
    end 
    if(N1916) begin
      { mem[5711:5696] } <= { w_data_i[15:0] };
    end 
    if(N1915) begin
      { mem[5695:5680] } <= { w_data_i[15:0] };
    end 
    if(N1914) begin
      { mem[5679:5664] } <= { w_data_i[15:0] };
    end 
    if(N1913) begin
      { mem[5663:5648] } <= { w_data_i[15:0] };
    end 
    if(N1912) begin
      { mem[5647:5632] } <= { w_data_i[15:0] };
    end 
    if(N1911) begin
      { mem[5631:5616] } <= { w_data_i[15:0] };
    end 
    if(N1910) begin
      { mem[5615:5600] } <= { w_data_i[15:0] };
    end 
    if(N1909) begin
      { mem[5599:5584] } <= { w_data_i[15:0] };
    end 
    if(N1908) begin
      { mem[5583:5568] } <= { w_data_i[15:0] };
    end 
    if(N1907) begin
      { mem[5567:5552] } <= { w_data_i[15:0] };
    end 
    if(N1906) begin
      { mem[5551:5536] } <= { w_data_i[15:0] };
    end 
    if(N1905) begin
      { mem[5535:5520] } <= { w_data_i[15:0] };
    end 
    if(N1904) begin
      { mem[5519:5504] } <= { w_data_i[15:0] };
    end 
    if(N1903) begin
      { mem[5503:5488] } <= { w_data_i[15:0] };
    end 
    if(N1902) begin
      { mem[5487:5472] } <= { w_data_i[15:0] };
    end 
    if(N1901) begin
      { mem[5471:5456] } <= { w_data_i[15:0] };
    end 
    if(N1900) begin
      { mem[5455:5440] } <= { w_data_i[15:0] };
    end 
    if(N1899) begin
      { mem[5439:5424] } <= { w_data_i[15:0] };
    end 
    if(N1898) begin
      { mem[5423:5408] } <= { w_data_i[15:0] };
    end 
    if(N1897) begin
      { mem[5407:5392] } <= { w_data_i[15:0] };
    end 
    if(N1896) begin
      { mem[5391:5376] } <= { w_data_i[15:0] };
    end 
    if(N1895) begin
      { mem[5375:5360] } <= { w_data_i[15:0] };
    end 
    if(N1894) begin
      { mem[5359:5344] } <= { w_data_i[15:0] };
    end 
    if(N1893) begin
      { mem[5343:5328] } <= { w_data_i[15:0] };
    end 
    if(N1892) begin
      { mem[5327:5312] } <= { w_data_i[15:0] };
    end 
    if(N1891) begin
      { mem[5311:5296] } <= { w_data_i[15:0] };
    end 
    if(N1890) begin
      { mem[5295:5280] } <= { w_data_i[15:0] };
    end 
    if(N1889) begin
      { mem[5279:5264] } <= { w_data_i[15:0] };
    end 
    if(N1888) begin
      { mem[5263:5248] } <= { w_data_i[15:0] };
    end 
    if(N1887) begin
      { mem[5247:5232] } <= { w_data_i[15:0] };
    end 
    if(N1886) begin
      { mem[5231:5216] } <= { w_data_i[15:0] };
    end 
    if(N1885) begin
      { mem[5215:5200] } <= { w_data_i[15:0] };
    end 
    if(N1884) begin
      { mem[5199:5184] } <= { w_data_i[15:0] };
    end 
    if(N1883) begin
      { mem[5183:5168] } <= { w_data_i[15:0] };
    end 
    if(N1882) begin
      { mem[5167:5152] } <= { w_data_i[15:0] };
    end 
    if(N1881) begin
      { mem[5151:5136] } <= { w_data_i[15:0] };
    end 
    if(N1880) begin
      { mem[5135:5120] } <= { w_data_i[15:0] };
    end 
    if(N1879) begin
      { mem[5119:5104] } <= { w_data_i[15:0] };
    end 
    if(N1878) begin
      { mem[5103:5088] } <= { w_data_i[15:0] };
    end 
    if(N1877) begin
      { mem[5087:5072] } <= { w_data_i[15:0] };
    end 
    if(N1876) begin
      { mem[5071:5056] } <= { w_data_i[15:0] };
    end 
    if(N1875) begin
      { mem[5055:5040] } <= { w_data_i[15:0] };
    end 
    if(N1874) begin
      { mem[5039:5024] } <= { w_data_i[15:0] };
    end 
    if(N1873) begin
      { mem[5023:5008] } <= { w_data_i[15:0] };
    end 
    if(N1872) begin
      { mem[5007:4992] } <= { w_data_i[15:0] };
    end 
    if(N1871) begin
      { mem[4991:4976] } <= { w_data_i[15:0] };
    end 
    if(N1870) begin
      { mem[4975:4960] } <= { w_data_i[15:0] };
    end 
    if(N1869) begin
      { mem[4959:4944] } <= { w_data_i[15:0] };
    end 
    if(N1868) begin
      { mem[4943:4928] } <= { w_data_i[15:0] };
    end 
    if(N1867) begin
      { mem[4927:4912] } <= { w_data_i[15:0] };
    end 
    if(N1866) begin
      { mem[4911:4896] } <= { w_data_i[15:0] };
    end 
    if(N1865) begin
      { mem[4895:4880] } <= { w_data_i[15:0] };
    end 
    if(N1864) begin
      { mem[4879:4864] } <= { w_data_i[15:0] };
    end 
    if(N1863) begin
      { mem[4863:4848] } <= { w_data_i[15:0] };
    end 
    if(N1862) begin
      { mem[4847:4832] } <= { w_data_i[15:0] };
    end 
    if(N1861) begin
      { mem[4831:4816] } <= { w_data_i[15:0] };
    end 
    if(N1860) begin
      { mem[4815:4800] } <= { w_data_i[15:0] };
    end 
    if(N1859) begin
      { mem[4799:4784] } <= { w_data_i[15:0] };
    end 
    if(N1858) begin
      { mem[4783:4768] } <= { w_data_i[15:0] };
    end 
    if(N1857) begin
      { mem[4767:4752] } <= { w_data_i[15:0] };
    end 
    if(N1856) begin
      { mem[4751:4736] } <= { w_data_i[15:0] };
    end 
    if(N1855) begin
      { mem[4735:4720] } <= { w_data_i[15:0] };
    end 
    if(N1854) begin
      { mem[4719:4704] } <= { w_data_i[15:0] };
    end 
    if(N1853) begin
      { mem[4703:4688] } <= { w_data_i[15:0] };
    end 
    if(N1852) begin
      { mem[4687:4672] } <= { w_data_i[15:0] };
    end 
    if(N1851) begin
      { mem[4671:4656] } <= { w_data_i[15:0] };
    end 
    if(N1850) begin
      { mem[4655:4640] } <= { w_data_i[15:0] };
    end 
    if(N1849) begin
      { mem[4639:4624] } <= { w_data_i[15:0] };
    end 
    if(N1848) begin
      { mem[4623:4608] } <= { w_data_i[15:0] };
    end 
    if(N1847) begin
      { mem[4607:4592] } <= { w_data_i[15:0] };
    end 
    if(N1846) begin
      { mem[4591:4576] } <= { w_data_i[15:0] };
    end 
    if(N1845) begin
      { mem[4575:4560] } <= { w_data_i[15:0] };
    end 
    if(N1844) begin
      { mem[4559:4544] } <= { w_data_i[15:0] };
    end 
    if(N1843) begin
      { mem[4543:4528] } <= { w_data_i[15:0] };
    end 
    if(N1842) begin
      { mem[4527:4512] } <= { w_data_i[15:0] };
    end 
    if(N1841) begin
      { mem[4511:4496] } <= { w_data_i[15:0] };
    end 
    if(N1840) begin
      { mem[4495:4480] } <= { w_data_i[15:0] };
    end 
    if(N1839) begin
      { mem[4479:4464] } <= { w_data_i[15:0] };
    end 
    if(N1838) begin
      { mem[4463:4448] } <= { w_data_i[15:0] };
    end 
    if(N1837) begin
      { mem[4447:4432] } <= { w_data_i[15:0] };
    end 
    if(N1836) begin
      { mem[4431:4416] } <= { w_data_i[15:0] };
    end 
    if(N1835) begin
      { mem[4415:4400] } <= { w_data_i[15:0] };
    end 
    if(N1834) begin
      { mem[4399:4384] } <= { w_data_i[15:0] };
    end 
    if(N1833) begin
      { mem[4383:4368] } <= { w_data_i[15:0] };
    end 
    if(N1832) begin
      { mem[4367:4352] } <= { w_data_i[15:0] };
    end 
    if(N1831) begin
      { mem[4351:4336] } <= { w_data_i[15:0] };
    end 
    if(N1830) begin
      { mem[4335:4320] } <= { w_data_i[15:0] };
    end 
    if(N1829) begin
      { mem[4319:4304] } <= { w_data_i[15:0] };
    end 
    if(N1828) begin
      { mem[4303:4288] } <= { w_data_i[15:0] };
    end 
    if(N1827) begin
      { mem[4287:4272] } <= { w_data_i[15:0] };
    end 
    if(N1826) begin
      { mem[4271:4256] } <= { w_data_i[15:0] };
    end 
    if(N1825) begin
      { mem[4255:4240] } <= { w_data_i[15:0] };
    end 
    if(N1824) begin
      { mem[4239:4224] } <= { w_data_i[15:0] };
    end 
    if(N1823) begin
      { mem[4223:4208] } <= { w_data_i[15:0] };
    end 
    if(N1822) begin
      { mem[4207:4192] } <= { w_data_i[15:0] };
    end 
    if(N1821) begin
      { mem[4191:4176] } <= { w_data_i[15:0] };
    end 
    if(N1820) begin
      { mem[4175:4160] } <= { w_data_i[15:0] };
    end 
    if(N1819) begin
      { mem[4159:4144] } <= { w_data_i[15:0] };
    end 
    if(N1818) begin
      { mem[4143:4128] } <= { w_data_i[15:0] };
    end 
    if(N1817) begin
      { mem[4127:4112] } <= { w_data_i[15:0] };
    end 
    if(N1816) begin
      { mem[4111:4096] } <= { w_data_i[15:0] };
    end 
    if(N1815) begin
      { mem[4095:4080] } <= { w_data_i[15:0] };
    end 
    if(N1814) begin
      { mem[4079:4064] } <= { w_data_i[15:0] };
    end 
    if(N1813) begin
      { mem[4063:4048] } <= { w_data_i[15:0] };
    end 
    if(N1812) begin
      { mem[4047:4032] } <= { w_data_i[15:0] };
    end 
    if(N1811) begin
      { mem[4031:4016] } <= { w_data_i[15:0] };
    end 
    if(N1810) begin
      { mem[4015:4000] } <= { w_data_i[15:0] };
    end 
    if(N1809) begin
      { mem[3999:3984] } <= { w_data_i[15:0] };
    end 
    if(N1808) begin
      { mem[3983:3968] } <= { w_data_i[15:0] };
    end 
    if(N1807) begin
      { mem[3967:3952] } <= { w_data_i[15:0] };
    end 
    if(N1806) begin
      { mem[3951:3936] } <= { w_data_i[15:0] };
    end 
    if(N1805) begin
      { mem[3935:3920] } <= { w_data_i[15:0] };
    end 
    if(N1804) begin
      { mem[3919:3904] } <= { w_data_i[15:0] };
    end 
    if(N1803) begin
      { mem[3903:3888] } <= { w_data_i[15:0] };
    end 
    if(N1802) begin
      { mem[3887:3872] } <= { w_data_i[15:0] };
    end 
    if(N1801) begin
      { mem[3871:3856] } <= { w_data_i[15:0] };
    end 
    if(N1800) begin
      { mem[3855:3840] } <= { w_data_i[15:0] };
    end 
    if(N1799) begin
      { mem[3839:3824] } <= { w_data_i[15:0] };
    end 
    if(N1798) begin
      { mem[3823:3808] } <= { w_data_i[15:0] };
    end 
    if(N1797) begin
      { mem[3807:3792] } <= { w_data_i[15:0] };
    end 
    if(N1796) begin
      { mem[3791:3776] } <= { w_data_i[15:0] };
    end 
    if(N1795) begin
      { mem[3775:3760] } <= { w_data_i[15:0] };
    end 
    if(N1794) begin
      { mem[3759:3744] } <= { w_data_i[15:0] };
    end 
    if(N1793) begin
      { mem[3743:3728] } <= { w_data_i[15:0] };
    end 
    if(N1792) begin
      { mem[3727:3712] } <= { w_data_i[15:0] };
    end 
    if(N1791) begin
      { mem[3711:3696] } <= { w_data_i[15:0] };
    end 
    if(N1790) begin
      { mem[3695:3680] } <= { w_data_i[15:0] };
    end 
    if(N1789) begin
      { mem[3679:3664] } <= { w_data_i[15:0] };
    end 
    if(N1788) begin
      { mem[3663:3648] } <= { w_data_i[15:0] };
    end 
    if(N1787) begin
      { mem[3647:3632] } <= { w_data_i[15:0] };
    end 
    if(N1786) begin
      { mem[3631:3616] } <= { w_data_i[15:0] };
    end 
    if(N1785) begin
      { mem[3615:3600] } <= { w_data_i[15:0] };
    end 
    if(N1784) begin
      { mem[3599:3584] } <= { w_data_i[15:0] };
    end 
    if(N1783) begin
      { mem[3583:3568] } <= { w_data_i[15:0] };
    end 
    if(N1782) begin
      { mem[3567:3552] } <= { w_data_i[15:0] };
    end 
    if(N1781) begin
      { mem[3551:3536] } <= { w_data_i[15:0] };
    end 
    if(N1780) begin
      { mem[3535:3520] } <= { w_data_i[15:0] };
    end 
    if(N1779) begin
      { mem[3519:3504] } <= { w_data_i[15:0] };
    end 
    if(N1778) begin
      { mem[3503:3488] } <= { w_data_i[15:0] };
    end 
    if(N1777) begin
      { mem[3487:3472] } <= { w_data_i[15:0] };
    end 
    if(N1776) begin
      { mem[3471:3456] } <= { w_data_i[15:0] };
    end 
    if(N1775) begin
      { mem[3455:3440] } <= { w_data_i[15:0] };
    end 
    if(N1774) begin
      { mem[3439:3424] } <= { w_data_i[15:0] };
    end 
    if(N1773) begin
      { mem[3423:3408] } <= { w_data_i[15:0] };
    end 
    if(N1772) begin
      { mem[3407:3392] } <= { w_data_i[15:0] };
    end 
    if(N1771) begin
      { mem[3391:3376] } <= { w_data_i[15:0] };
    end 
    if(N1770) begin
      { mem[3375:3360] } <= { w_data_i[15:0] };
    end 
    if(N1769) begin
      { mem[3359:3344] } <= { w_data_i[15:0] };
    end 
    if(N1768) begin
      { mem[3343:3328] } <= { w_data_i[15:0] };
    end 
    if(N1767) begin
      { mem[3327:3312] } <= { w_data_i[15:0] };
    end 
    if(N1766) begin
      { mem[3311:3296] } <= { w_data_i[15:0] };
    end 
    if(N1765) begin
      { mem[3295:3280] } <= { w_data_i[15:0] };
    end 
    if(N1764) begin
      { mem[3279:3264] } <= { w_data_i[15:0] };
    end 
    if(N1763) begin
      { mem[3263:3248] } <= { w_data_i[15:0] };
    end 
    if(N1762) begin
      { mem[3247:3232] } <= { w_data_i[15:0] };
    end 
    if(N1761) begin
      { mem[3231:3216] } <= { w_data_i[15:0] };
    end 
    if(N1760) begin
      { mem[3215:3200] } <= { w_data_i[15:0] };
    end 
    if(N1759) begin
      { mem[3199:3184] } <= { w_data_i[15:0] };
    end 
    if(N1758) begin
      { mem[3183:3168] } <= { w_data_i[15:0] };
    end 
    if(N1757) begin
      { mem[3167:3152] } <= { w_data_i[15:0] };
    end 
    if(N1756) begin
      { mem[3151:3136] } <= { w_data_i[15:0] };
    end 
    if(N1755) begin
      { mem[3135:3120] } <= { w_data_i[15:0] };
    end 
    if(N1754) begin
      { mem[3119:3104] } <= { w_data_i[15:0] };
    end 
    if(N1753) begin
      { mem[3103:3088] } <= { w_data_i[15:0] };
    end 
    if(N1752) begin
      { mem[3087:3072] } <= { w_data_i[15:0] };
    end 
    if(N1751) begin
      { mem[3071:3056] } <= { w_data_i[15:0] };
    end 
    if(N1750) begin
      { mem[3055:3040] } <= { w_data_i[15:0] };
    end 
    if(N1749) begin
      { mem[3039:3024] } <= { w_data_i[15:0] };
    end 
    if(N1748) begin
      { mem[3023:3008] } <= { w_data_i[15:0] };
    end 
    if(N1747) begin
      { mem[3007:2992] } <= { w_data_i[15:0] };
    end 
    if(N1746) begin
      { mem[2991:2976] } <= { w_data_i[15:0] };
    end 
    if(N1745) begin
      { mem[2975:2960] } <= { w_data_i[15:0] };
    end 
    if(N1744) begin
      { mem[2959:2944] } <= { w_data_i[15:0] };
    end 
    if(N1743) begin
      { mem[2943:2928] } <= { w_data_i[15:0] };
    end 
    if(N1742) begin
      { mem[2927:2912] } <= { w_data_i[15:0] };
    end 
    if(N1741) begin
      { mem[2911:2896] } <= { w_data_i[15:0] };
    end 
    if(N1740) begin
      { mem[2895:2880] } <= { w_data_i[15:0] };
    end 
    if(N1739) begin
      { mem[2879:2864] } <= { w_data_i[15:0] };
    end 
    if(N1738) begin
      { mem[2863:2848] } <= { w_data_i[15:0] };
    end 
    if(N1737) begin
      { mem[2847:2832] } <= { w_data_i[15:0] };
    end 
    if(N1736) begin
      { mem[2831:2816] } <= { w_data_i[15:0] };
    end 
    if(N1735) begin
      { mem[2815:2800] } <= { w_data_i[15:0] };
    end 
    if(N1734) begin
      { mem[2799:2784] } <= { w_data_i[15:0] };
    end 
    if(N1733) begin
      { mem[2783:2768] } <= { w_data_i[15:0] };
    end 
    if(N1732) begin
      { mem[2767:2752] } <= { w_data_i[15:0] };
    end 
    if(N1731) begin
      { mem[2751:2736] } <= { w_data_i[15:0] };
    end 
    if(N1730) begin
      { mem[2735:2720] } <= { w_data_i[15:0] };
    end 
    if(N1729) begin
      { mem[2719:2704] } <= { w_data_i[15:0] };
    end 
    if(N1728) begin
      { mem[2703:2688] } <= { w_data_i[15:0] };
    end 
    if(N1727) begin
      { mem[2687:2672] } <= { w_data_i[15:0] };
    end 
    if(N1726) begin
      { mem[2671:2656] } <= { w_data_i[15:0] };
    end 
    if(N1725) begin
      { mem[2655:2640] } <= { w_data_i[15:0] };
    end 
    if(N1724) begin
      { mem[2639:2624] } <= { w_data_i[15:0] };
    end 
    if(N1723) begin
      { mem[2623:2608] } <= { w_data_i[15:0] };
    end 
    if(N1722) begin
      { mem[2607:2592] } <= { w_data_i[15:0] };
    end 
    if(N1721) begin
      { mem[2591:2576] } <= { w_data_i[15:0] };
    end 
    if(N1720) begin
      { mem[2575:2560] } <= { w_data_i[15:0] };
    end 
    if(N1719) begin
      { mem[2559:2544] } <= { w_data_i[15:0] };
    end 
    if(N1718) begin
      { mem[2543:2528] } <= { w_data_i[15:0] };
    end 
    if(N1717) begin
      { mem[2527:2512] } <= { w_data_i[15:0] };
    end 
    if(N1716) begin
      { mem[2511:2496] } <= { w_data_i[15:0] };
    end 
    if(N1715) begin
      { mem[2495:2480] } <= { w_data_i[15:0] };
    end 
    if(N1714) begin
      { mem[2479:2464] } <= { w_data_i[15:0] };
    end 
    if(N1713) begin
      { mem[2463:2448] } <= { w_data_i[15:0] };
    end 
    if(N1712) begin
      { mem[2447:2432] } <= { w_data_i[15:0] };
    end 
    if(N1711) begin
      { mem[2431:2416] } <= { w_data_i[15:0] };
    end 
    if(N1710) begin
      { mem[2415:2400] } <= { w_data_i[15:0] };
    end 
    if(N1709) begin
      { mem[2399:2384] } <= { w_data_i[15:0] };
    end 
    if(N1708) begin
      { mem[2383:2368] } <= { w_data_i[15:0] };
    end 
    if(N1707) begin
      { mem[2367:2352] } <= { w_data_i[15:0] };
    end 
    if(N1706) begin
      { mem[2351:2336] } <= { w_data_i[15:0] };
    end 
    if(N1705) begin
      { mem[2335:2320] } <= { w_data_i[15:0] };
    end 
    if(N1704) begin
      { mem[2319:2304] } <= { w_data_i[15:0] };
    end 
    if(N1703) begin
      { mem[2303:2288] } <= { w_data_i[15:0] };
    end 
    if(N1702) begin
      { mem[2287:2272] } <= { w_data_i[15:0] };
    end 
    if(N1701) begin
      { mem[2271:2256] } <= { w_data_i[15:0] };
    end 
    if(N1700) begin
      { mem[2255:2240] } <= { w_data_i[15:0] };
    end 
    if(N1699) begin
      { mem[2239:2224] } <= { w_data_i[15:0] };
    end 
    if(N1698) begin
      { mem[2223:2208] } <= { w_data_i[15:0] };
    end 
    if(N1697) begin
      { mem[2207:2192] } <= { w_data_i[15:0] };
    end 
    if(N1696) begin
      { mem[2191:2176] } <= { w_data_i[15:0] };
    end 
    if(N1695) begin
      { mem[2175:2160] } <= { w_data_i[15:0] };
    end 
    if(N1694) begin
      { mem[2159:2144] } <= { w_data_i[15:0] };
    end 
    if(N1693) begin
      { mem[2143:2128] } <= { w_data_i[15:0] };
    end 
    if(N1692) begin
      { mem[2127:2112] } <= { w_data_i[15:0] };
    end 
    if(N1691) begin
      { mem[2111:2096] } <= { w_data_i[15:0] };
    end 
    if(N1690) begin
      { mem[2095:2080] } <= { w_data_i[15:0] };
    end 
    if(N1689) begin
      { mem[2079:2064] } <= { w_data_i[15:0] };
    end 
    if(N1688) begin
      { mem[2063:2048] } <= { w_data_i[15:0] };
    end 
    if(N1687) begin
      { mem[2047:2032] } <= { w_data_i[15:0] };
    end 
    if(N1686) begin
      { mem[2031:2016] } <= { w_data_i[15:0] };
    end 
    if(N1685) begin
      { mem[2015:2000] } <= { w_data_i[15:0] };
    end 
    if(N1684) begin
      { mem[1999:1984] } <= { w_data_i[15:0] };
    end 
    if(N1683) begin
      { mem[1983:1968] } <= { w_data_i[15:0] };
    end 
    if(N1682) begin
      { mem[1967:1952] } <= { w_data_i[15:0] };
    end 
    if(N1681) begin
      { mem[1951:1936] } <= { w_data_i[15:0] };
    end 
    if(N1680) begin
      { mem[1935:1920] } <= { w_data_i[15:0] };
    end 
    if(N1679) begin
      { mem[1919:1904] } <= { w_data_i[15:0] };
    end 
    if(N1678) begin
      { mem[1903:1888] } <= { w_data_i[15:0] };
    end 
    if(N1677) begin
      { mem[1887:1872] } <= { w_data_i[15:0] };
    end 
    if(N1676) begin
      { mem[1871:1856] } <= { w_data_i[15:0] };
    end 
    if(N1675) begin
      { mem[1855:1840] } <= { w_data_i[15:0] };
    end 
    if(N1674) begin
      { mem[1839:1824] } <= { w_data_i[15:0] };
    end 
    if(N1673) begin
      { mem[1823:1808] } <= { w_data_i[15:0] };
    end 
    if(N1672) begin
      { mem[1807:1792] } <= { w_data_i[15:0] };
    end 
    if(N1671) begin
      { mem[1791:1776] } <= { w_data_i[15:0] };
    end 
    if(N1670) begin
      { mem[1775:1760] } <= { w_data_i[15:0] };
    end 
    if(N1669) begin
      { mem[1759:1744] } <= { w_data_i[15:0] };
    end 
    if(N1668) begin
      { mem[1743:1728] } <= { w_data_i[15:0] };
    end 
    if(N1667) begin
      { mem[1727:1712] } <= { w_data_i[15:0] };
    end 
    if(N1666) begin
      { mem[1711:1696] } <= { w_data_i[15:0] };
    end 
    if(N1665) begin
      { mem[1695:1680] } <= { w_data_i[15:0] };
    end 
    if(N1664) begin
      { mem[1679:1664] } <= { w_data_i[15:0] };
    end 
    if(N1663) begin
      { mem[1663:1648] } <= { w_data_i[15:0] };
    end 
    if(N1662) begin
      { mem[1647:1632] } <= { w_data_i[15:0] };
    end 
    if(N1661) begin
      { mem[1631:1616] } <= { w_data_i[15:0] };
    end 
    if(N1660) begin
      { mem[1615:1600] } <= { w_data_i[15:0] };
    end 
    if(N1659) begin
      { mem[1599:1584] } <= { w_data_i[15:0] };
    end 
    if(N1658) begin
      { mem[1583:1568] } <= { w_data_i[15:0] };
    end 
    if(N1657) begin
      { mem[1567:1552] } <= { w_data_i[15:0] };
    end 
    if(N1656) begin
      { mem[1551:1536] } <= { w_data_i[15:0] };
    end 
    if(N1655) begin
      { mem[1535:1520] } <= { w_data_i[15:0] };
    end 
    if(N1654) begin
      { mem[1519:1504] } <= { w_data_i[15:0] };
    end 
    if(N1653) begin
      { mem[1503:1488] } <= { w_data_i[15:0] };
    end 
    if(N1652) begin
      { mem[1487:1472] } <= { w_data_i[15:0] };
    end 
    if(N1651) begin
      { mem[1471:1456] } <= { w_data_i[15:0] };
    end 
    if(N1650) begin
      { mem[1455:1440] } <= { w_data_i[15:0] };
    end 
    if(N1649) begin
      { mem[1439:1424] } <= { w_data_i[15:0] };
    end 
    if(N1648) begin
      { mem[1423:1408] } <= { w_data_i[15:0] };
    end 
    if(N1647) begin
      { mem[1407:1392] } <= { w_data_i[15:0] };
    end 
    if(N1646) begin
      { mem[1391:1376] } <= { w_data_i[15:0] };
    end 
    if(N1645) begin
      { mem[1375:1360] } <= { w_data_i[15:0] };
    end 
    if(N1644) begin
      { mem[1359:1344] } <= { w_data_i[15:0] };
    end 
    if(N1643) begin
      { mem[1343:1328] } <= { w_data_i[15:0] };
    end 
    if(N1642) begin
      { mem[1327:1312] } <= { w_data_i[15:0] };
    end 
    if(N1641) begin
      { mem[1311:1296] } <= { w_data_i[15:0] };
    end 
    if(N1640) begin
      { mem[1295:1280] } <= { w_data_i[15:0] };
    end 
    if(N1639) begin
      { mem[1279:1264] } <= { w_data_i[15:0] };
    end 
    if(N1638) begin
      { mem[1263:1248] } <= { w_data_i[15:0] };
    end 
    if(N1637) begin
      { mem[1247:1232] } <= { w_data_i[15:0] };
    end 
    if(N1636) begin
      { mem[1231:1216] } <= { w_data_i[15:0] };
    end 
    if(N1635) begin
      { mem[1215:1200] } <= { w_data_i[15:0] };
    end 
    if(N1634) begin
      { mem[1199:1184] } <= { w_data_i[15:0] };
    end 
    if(N1633) begin
      { mem[1183:1168] } <= { w_data_i[15:0] };
    end 
    if(N1632) begin
      { mem[1167:1152] } <= { w_data_i[15:0] };
    end 
    if(N1631) begin
      { mem[1151:1136] } <= { w_data_i[15:0] };
    end 
    if(N1630) begin
      { mem[1135:1120] } <= { w_data_i[15:0] };
    end 
    if(N1629) begin
      { mem[1119:1104] } <= { w_data_i[15:0] };
    end 
    if(N1628) begin
      { mem[1103:1088] } <= { w_data_i[15:0] };
    end 
    if(N1627) begin
      { mem[1087:1072] } <= { w_data_i[15:0] };
    end 
    if(N1626) begin
      { mem[1071:1056] } <= { w_data_i[15:0] };
    end 
    if(N1625) begin
      { mem[1055:1040] } <= { w_data_i[15:0] };
    end 
    if(N1624) begin
      { mem[1039:1024] } <= { w_data_i[15:0] };
    end 
    if(N1623) begin
      { mem[1023:1008] } <= { w_data_i[15:0] };
    end 
    if(N1622) begin
      { mem[1007:992] } <= { w_data_i[15:0] };
    end 
    if(N1621) begin
      { mem[991:976] } <= { w_data_i[15:0] };
    end 
    if(N1620) begin
      { mem[975:960] } <= { w_data_i[15:0] };
    end 
    if(N1619) begin
      { mem[959:944] } <= { w_data_i[15:0] };
    end 
    if(N1618) begin
      { mem[943:928] } <= { w_data_i[15:0] };
    end 
    if(N1617) begin
      { mem[927:912] } <= { w_data_i[15:0] };
    end 
    if(N1616) begin
      { mem[911:896] } <= { w_data_i[15:0] };
    end 
    if(N1615) begin
      { mem[895:880] } <= { w_data_i[15:0] };
    end 
    if(N1614) begin
      { mem[879:864] } <= { w_data_i[15:0] };
    end 
    if(N1613) begin
      { mem[863:848] } <= { w_data_i[15:0] };
    end 
    if(N1612) begin
      { mem[847:832] } <= { w_data_i[15:0] };
    end 
    if(N1611) begin
      { mem[831:816] } <= { w_data_i[15:0] };
    end 
    if(N1610) begin
      { mem[815:800] } <= { w_data_i[15:0] };
    end 
    if(N1609) begin
      { mem[799:784] } <= { w_data_i[15:0] };
    end 
    if(N1608) begin
      { mem[783:768] } <= { w_data_i[15:0] };
    end 
    if(N1607) begin
      { mem[767:752] } <= { w_data_i[15:0] };
    end 
    if(N1606) begin
      { mem[751:736] } <= { w_data_i[15:0] };
    end 
    if(N1605) begin
      { mem[735:720] } <= { w_data_i[15:0] };
    end 
    if(N1604) begin
      { mem[719:704] } <= { w_data_i[15:0] };
    end 
    if(N1603) begin
      { mem[703:688] } <= { w_data_i[15:0] };
    end 
    if(N1602) begin
      { mem[687:672] } <= { w_data_i[15:0] };
    end 
    if(N1601) begin
      { mem[671:656] } <= { w_data_i[15:0] };
    end 
    if(N1600) begin
      { mem[655:640] } <= { w_data_i[15:0] };
    end 
    if(N1599) begin
      { mem[639:624] } <= { w_data_i[15:0] };
    end 
    if(N1598) begin
      { mem[623:608] } <= { w_data_i[15:0] };
    end 
    if(N1597) begin
      { mem[607:592] } <= { w_data_i[15:0] };
    end 
    if(N1596) begin
      { mem[591:576] } <= { w_data_i[15:0] };
    end 
    if(N1595) begin
      { mem[575:560] } <= { w_data_i[15:0] };
    end 
    if(N1594) begin
      { mem[559:544] } <= { w_data_i[15:0] };
    end 
    if(N1593) begin
      { mem[543:528] } <= { w_data_i[15:0] };
    end 
    if(N1592) begin
      { mem[527:512] } <= { w_data_i[15:0] };
    end 
    if(N1591) begin
      { mem[511:496] } <= { w_data_i[15:0] };
    end 
    if(N1590) begin
      { mem[495:480] } <= { w_data_i[15:0] };
    end 
    if(N1589) begin
      { mem[479:464] } <= { w_data_i[15:0] };
    end 
    if(N1588) begin
      { mem[463:448] } <= { w_data_i[15:0] };
    end 
    if(N1587) begin
      { mem[447:432] } <= { w_data_i[15:0] };
    end 
    if(N1586) begin
      { mem[431:416] } <= { w_data_i[15:0] };
    end 
    if(N1585) begin
      { mem[415:400] } <= { w_data_i[15:0] };
    end 
    if(N1584) begin
      { mem[399:384] } <= { w_data_i[15:0] };
    end 
    if(N1583) begin
      { mem[383:368] } <= { w_data_i[15:0] };
    end 
    if(N1582) begin
      { mem[367:352] } <= { w_data_i[15:0] };
    end 
    if(N1581) begin
      { mem[351:336] } <= { w_data_i[15:0] };
    end 
    if(N1580) begin
      { mem[335:320] } <= { w_data_i[15:0] };
    end 
    if(N1579) begin
      { mem[319:304] } <= { w_data_i[15:0] };
    end 
    if(N1578) begin
      { mem[303:288] } <= { w_data_i[15:0] };
    end 
    if(N1577) begin
      { mem[287:272] } <= { w_data_i[15:0] };
    end 
    if(N1576) begin
      { mem[271:256] } <= { w_data_i[15:0] };
    end 
    if(N1575) begin
      { mem[255:240] } <= { w_data_i[15:0] };
    end 
    if(N1574) begin
      { mem[239:224] } <= { w_data_i[15:0] };
    end 
    if(N1573) begin
      { mem[223:208] } <= { w_data_i[15:0] };
    end 
    if(N1572) begin
      { mem[207:192] } <= { w_data_i[15:0] };
    end 
    if(N1571) begin
      { mem[191:176] } <= { w_data_i[15:0] };
    end 
    if(N1570) begin
      { mem[175:160] } <= { w_data_i[15:0] };
    end 
    if(N1569) begin
      { mem[159:144] } <= { w_data_i[15:0] };
    end 
    if(N1568) begin
      { mem[143:128] } <= { w_data_i[15:0] };
    end 
    if(N1567) begin
      { mem[127:112] } <= { w_data_i[15:0] };
    end 
    if(N1566) begin
      { mem[111:96] } <= { w_data_i[15:0] };
    end 
    if(N1565) begin
      { mem[95:80] } <= { w_data_i[15:0] };
    end 
    if(N1564) begin
      { mem[79:64] } <= { w_data_i[15:0] };
    end 
    if(N1563) begin
      { mem[63:48] } <= { w_data_i[15:0] };
    end 
    if(N1562) begin
      { mem[47:32] } <= { w_data_i[15:0] };
    end 
    if(N1561) begin
      { mem[31:16] } <= { w_data_i[15:0] };
    end 
    if(N1560) begin
      { mem[15:0] } <= { w_data_i[15:0] };
    end 
  end


endmodule



module bsg_mem_1r1w_sync_width_p16_els_p512_read_write_same_addr_p0
(
  clk_i,
  reset_i,
  w_v_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_addr_i,
  r_data_o
);

  input [8:0] w_addr_i;
  input [15:0] w_data_i;
  input [8:0] r_addr_i;
  output [15:0] r_data_o;
  input clk_i;
  input reset_i;
  input w_v_i;
  input r_v_i;
  wire [15:0] r_data_o;

  bsg_mem_1r1w_sync_synth_width_p16_els_p512_read_write_same_addr_p0_harden_p0
  synth
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .w_v_i(w_v_i),
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_v_i(r_v_i),
    .r_addr_i(r_addr_i),
    .r_data_o(r_data_o)
  );


endmodule

