

module top
(
  ready_i,
  reqs_i,
  grants_o
);

  input [127:0] reqs_i;
  output [127:0] grants_o;
  input ready_i;

  bsg_arb_fixed
  wrapper
  (
    .reqs_i(reqs_i),
    .grants_o(grants_o),
    .ready_i(ready_i)
  );


endmodule



module bsg_scan_width_p128_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [127:0] i;
  output [127:0] o;
  wire [127:0] o;
  wire t_3__127_,t_3__126_,t_3__125_,t_3__124_,t_3__123_,t_3__122_,t_3__121_,t_3__120_,
  t_3__119_,t_3__118_,t_3__117_,t_3__116_,t_3__115_,t_3__114_,t_3__113_,t_3__112_,
  t_3__111_,t_3__110_,t_3__109_,t_3__108_,t_3__107_,t_3__106_,t_3__105_,t_3__104_,
  t_3__103_,t_3__102_,t_3__101_,t_3__100_,t_3__99_,t_3__98_,t_3__97_,t_3__96_,
  t_3__95_,t_3__94_,t_3__93_,t_3__92_,t_3__91_,t_3__90_,t_3__89_,t_3__88_,t_3__87_,
  t_3__86_,t_3__85_,t_3__84_,t_3__83_,t_3__82_,t_3__81_,t_3__80_,t_3__79_,t_3__78_,
  t_3__77_,t_3__76_,t_3__75_,t_3__74_,t_3__73_,t_3__72_,t_3__71_,t_3__70_,t_3__69_,
  t_3__68_,t_3__67_,t_3__66_,t_3__65_,t_3__64_,t_3__63_,t_3__62_,t_3__61_,t_3__60_,
  t_3__59_,t_3__58_,t_3__57_,t_3__56_,t_3__55_,t_3__54_,t_3__53_,t_3__52_,
  t_3__51_,t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,t_3__45_,t_3__44_,t_3__43_,
  t_3__42_,t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,t_3__36_,t_3__35_,t_3__34_,
  t_3__33_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,t_3__26_,t_3__25_,
  t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,t_3__17_,t_3__16_,
  t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,
  t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_2__127_,t_2__126_,t_2__125_,
  t_2__124_,t_2__123_,t_2__122_,t_2__121_,t_2__120_,t_2__119_,t_2__118_,t_2__117_,
  t_2__116_,t_2__115_,t_2__114_,t_2__113_,t_2__112_,t_2__111_,t_2__110_,t_2__109_,
  t_2__108_,t_2__107_,t_2__106_,t_2__105_,t_2__104_,t_2__103_,t_2__102_,t_2__101_,
  t_2__100_,t_2__99_,t_2__98_,t_2__97_,t_2__96_,t_2__95_,t_2__94_,t_2__93_,
  t_2__92_,t_2__91_,t_2__90_,t_2__89_,t_2__88_,t_2__87_,t_2__86_,t_2__85_,t_2__84_,
  t_2__83_,t_2__82_,t_2__81_,t_2__80_,t_2__79_,t_2__78_,t_2__77_,t_2__76_,t_2__75_,
  t_2__74_,t_2__73_,t_2__72_,t_2__71_,t_2__70_,t_2__69_,t_2__68_,t_2__67_,t_2__66_,
  t_2__65_,t_2__64_,t_2__63_,t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,t_2__57_,
  t_2__56_,t_2__55_,t_2__54_,t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,t_2__48_,
  t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,t_2__39_,
  t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,t_2__30_,
  t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,
  t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,
  t_2__2_,t_2__1_,t_2__0_,t_1__127_,t_1__126_,t_1__125_,t_1__124_,t_1__123_,t_1__122_,
  t_1__121_,t_1__120_,t_1__119_,t_1__118_,t_1__117_,t_1__116_,t_1__115_,t_1__114_,
  t_1__113_,t_1__112_,t_1__111_,t_1__110_,t_1__109_,t_1__108_,t_1__107_,t_1__106_,
  t_1__105_,t_1__104_,t_1__103_,t_1__102_,t_1__101_,t_1__100_,t_1__99_,t_1__98_,
  t_1__97_,t_1__96_,t_1__95_,t_1__94_,t_1__93_,t_1__92_,t_1__91_,t_1__90_,t_1__89_,
  t_1__88_,t_1__87_,t_1__86_,t_1__85_,t_1__84_,t_1__83_,t_1__82_,t_1__81_,t_1__80_,
  t_1__79_,t_1__78_,t_1__77_,t_1__76_,t_1__75_,t_1__74_,t_1__73_,t_1__72_,
  t_1__71_,t_1__70_,t_1__69_,t_1__68_,t_1__67_,t_1__66_,t_1__65_,t_1__64_,t_1__63_,
  t_1__62_,t_1__61_,t_1__60_,t_1__59_,t_1__58_,t_1__57_,t_1__56_,t_1__55_,t_1__54_,
  t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,t_1__48_,t_1__47_,t_1__46_,t_1__45_,
  t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,t_1__39_,t_1__38_,t_1__37_,t_1__36_,
  t_1__35_,t_1__34_,t_1__33_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,t_1__27_,
  t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,t_1__18_,
  t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,t_1__9_,
  t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_,t_6__127_,
  t_6__126_,t_6__125_,t_6__124_,t_6__123_,t_6__122_,t_6__121_,t_6__120_,t_6__119_,
  t_6__118_,t_6__117_,t_6__116_,t_6__115_,t_6__114_,t_6__113_,t_6__112_,t_6__111_,
  t_6__110_,t_6__109_,t_6__108_,t_6__107_,t_6__106_,t_6__105_,t_6__104_,t_6__103_,
  t_6__102_,t_6__101_,t_6__100_,t_6__99_,t_6__98_,t_6__97_,t_6__96_,t_6__95_,
  t_6__94_,t_6__93_,t_6__92_,t_6__91_,t_6__90_,t_6__89_,t_6__88_,t_6__87_,t_6__86_,
  t_6__85_,t_6__84_,t_6__83_,t_6__82_,t_6__81_,t_6__80_,t_6__79_,t_6__78_,t_6__77_,
  t_6__76_,t_6__75_,t_6__74_,t_6__73_,t_6__72_,t_6__71_,t_6__70_,t_6__69_,t_6__68_,
  t_6__67_,t_6__66_,t_6__65_,t_6__64_,t_6__63_,t_6__62_,t_6__61_,t_6__60_,t_6__59_,
  t_6__58_,t_6__57_,t_6__56_,t_6__55_,t_6__54_,t_6__53_,t_6__52_,t_6__51_,t_6__50_,
  t_6__49_,t_6__48_,t_6__47_,t_6__46_,t_6__45_,t_6__44_,t_6__43_,t_6__42_,
  t_6__41_,t_6__40_,t_6__39_,t_6__38_,t_6__37_,t_6__36_,t_6__35_,t_6__34_,t_6__33_,
  t_6__32_,t_6__31_,t_6__30_,t_6__29_,t_6__28_,t_6__27_,t_6__26_,t_6__25_,t_6__24_,
  t_6__23_,t_6__22_,t_6__21_,t_6__20_,t_6__19_,t_6__18_,t_6__17_,t_6__16_,t_6__15_,
  t_6__14_,t_6__13_,t_6__12_,t_6__11_,t_6__10_,t_6__9_,t_6__8_,t_6__7_,t_6__6_,t_6__5_,
  t_6__4_,t_6__3_,t_6__2_,t_6__1_,t_6__0_,t_5__127_,t_5__126_,t_5__125_,t_5__124_,
  t_5__123_,t_5__122_,t_5__121_,t_5__120_,t_5__119_,t_5__118_,t_5__117_,t_5__116_,
  t_5__115_,t_5__114_,t_5__113_,t_5__112_,t_5__111_,t_5__110_,t_5__109_,t_5__108_,
  t_5__107_,t_5__106_,t_5__105_,t_5__104_,t_5__103_,t_5__102_,t_5__101_,t_5__100_,
  t_5__99_,t_5__98_,t_5__97_,t_5__96_,t_5__95_,t_5__94_,t_5__93_,t_5__92_,
  t_5__91_,t_5__90_,t_5__89_,t_5__88_,t_5__87_,t_5__86_,t_5__85_,t_5__84_,t_5__83_,
  t_5__82_,t_5__81_,t_5__80_,t_5__79_,t_5__78_,t_5__77_,t_5__76_,t_5__75_,t_5__74_,
  t_5__73_,t_5__72_,t_5__71_,t_5__70_,t_5__69_,t_5__68_,t_5__67_,t_5__66_,t_5__65_,
  t_5__64_,t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,t_5__58_,t_5__57_,t_5__56_,
  t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,
  t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,
  t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,
  t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,
  t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,
  t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,
  t_5__1_,t_5__0_,t_4__127_,t_4__126_,t_4__125_,t_4__124_,t_4__123_,t_4__122_,t_4__121_,
  t_4__120_,t_4__119_,t_4__118_,t_4__117_,t_4__116_,t_4__115_,t_4__114_,t_4__113_,
  t_4__112_,t_4__111_,t_4__110_,t_4__109_,t_4__108_,t_4__107_,t_4__106_,t_4__105_,
  t_4__104_,t_4__103_,t_4__102_,t_4__101_,t_4__100_,t_4__99_,t_4__98_,t_4__97_,
  t_4__96_,t_4__95_,t_4__94_,t_4__93_,t_4__92_,t_4__91_,t_4__90_,t_4__89_,t_4__88_,
  t_4__87_,t_4__86_,t_4__85_,t_4__84_,t_4__83_,t_4__82_,t_4__81_,t_4__80_,t_4__79_,
  t_4__78_,t_4__77_,t_4__76_,t_4__75_,t_4__74_,t_4__73_,t_4__72_,t_4__71_,t_4__70_,
  t_4__69_,t_4__68_,t_4__67_,t_4__66_,t_4__65_,t_4__64_,t_4__63_,t_4__62_,
  t_4__61_,t_4__60_,t_4__59_,t_4__58_,t_4__57_,t_4__56_,t_4__55_,t_4__54_,t_4__53_,
  t_4__52_,t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,
  t_4__43_,t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,
  t_4__34_,t_4__33_,t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,
  t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,
  t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,
  t_4__7_,t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_;
  assign t_1__127_ = i[0] | 1'b0;
  assign t_1__126_ = i[1] | i[0];
  assign t_1__125_ = i[2] | i[1];
  assign t_1__124_ = i[3] | i[2];
  assign t_1__123_ = i[4] | i[3];
  assign t_1__122_ = i[5] | i[4];
  assign t_1__121_ = i[6] | i[5];
  assign t_1__120_ = i[7] | i[6];
  assign t_1__119_ = i[8] | i[7];
  assign t_1__118_ = i[9] | i[8];
  assign t_1__117_ = i[10] | i[9];
  assign t_1__116_ = i[11] | i[10];
  assign t_1__115_ = i[12] | i[11];
  assign t_1__114_ = i[13] | i[12];
  assign t_1__113_ = i[14] | i[13];
  assign t_1__112_ = i[15] | i[14];
  assign t_1__111_ = i[16] | i[15];
  assign t_1__110_ = i[17] | i[16];
  assign t_1__109_ = i[18] | i[17];
  assign t_1__108_ = i[19] | i[18];
  assign t_1__107_ = i[20] | i[19];
  assign t_1__106_ = i[21] | i[20];
  assign t_1__105_ = i[22] | i[21];
  assign t_1__104_ = i[23] | i[22];
  assign t_1__103_ = i[24] | i[23];
  assign t_1__102_ = i[25] | i[24];
  assign t_1__101_ = i[26] | i[25];
  assign t_1__100_ = i[27] | i[26];
  assign t_1__99_ = i[28] | i[27];
  assign t_1__98_ = i[29] | i[28];
  assign t_1__97_ = i[30] | i[29];
  assign t_1__96_ = i[31] | i[30];
  assign t_1__95_ = i[32] | i[31];
  assign t_1__94_ = i[33] | i[32];
  assign t_1__93_ = i[34] | i[33];
  assign t_1__92_ = i[35] | i[34];
  assign t_1__91_ = i[36] | i[35];
  assign t_1__90_ = i[37] | i[36];
  assign t_1__89_ = i[38] | i[37];
  assign t_1__88_ = i[39] | i[38];
  assign t_1__87_ = i[40] | i[39];
  assign t_1__86_ = i[41] | i[40];
  assign t_1__85_ = i[42] | i[41];
  assign t_1__84_ = i[43] | i[42];
  assign t_1__83_ = i[44] | i[43];
  assign t_1__82_ = i[45] | i[44];
  assign t_1__81_ = i[46] | i[45];
  assign t_1__80_ = i[47] | i[46];
  assign t_1__79_ = i[48] | i[47];
  assign t_1__78_ = i[49] | i[48];
  assign t_1__77_ = i[50] | i[49];
  assign t_1__76_ = i[51] | i[50];
  assign t_1__75_ = i[52] | i[51];
  assign t_1__74_ = i[53] | i[52];
  assign t_1__73_ = i[54] | i[53];
  assign t_1__72_ = i[55] | i[54];
  assign t_1__71_ = i[56] | i[55];
  assign t_1__70_ = i[57] | i[56];
  assign t_1__69_ = i[58] | i[57];
  assign t_1__68_ = i[59] | i[58];
  assign t_1__67_ = i[60] | i[59];
  assign t_1__66_ = i[61] | i[60];
  assign t_1__65_ = i[62] | i[61];
  assign t_1__64_ = i[63] | i[62];
  assign t_1__63_ = i[64] | i[63];
  assign t_1__62_ = i[65] | i[64];
  assign t_1__61_ = i[66] | i[65];
  assign t_1__60_ = i[67] | i[66];
  assign t_1__59_ = i[68] | i[67];
  assign t_1__58_ = i[69] | i[68];
  assign t_1__57_ = i[70] | i[69];
  assign t_1__56_ = i[71] | i[70];
  assign t_1__55_ = i[72] | i[71];
  assign t_1__54_ = i[73] | i[72];
  assign t_1__53_ = i[74] | i[73];
  assign t_1__52_ = i[75] | i[74];
  assign t_1__51_ = i[76] | i[75];
  assign t_1__50_ = i[77] | i[76];
  assign t_1__49_ = i[78] | i[77];
  assign t_1__48_ = i[79] | i[78];
  assign t_1__47_ = i[80] | i[79];
  assign t_1__46_ = i[81] | i[80];
  assign t_1__45_ = i[82] | i[81];
  assign t_1__44_ = i[83] | i[82];
  assign t_1__43_ = i[84] | i[83];
  assign t_1__42_ = i[85] | i[84];
  assign t_1__41_ = i[86] | i[85];
  assign t_1__40_ = i[87] | i[86];
  assign t_1__39_ = i[88] | i[87];
  assign t_1__38_ = i[89] | i[88];
  assign t_1__37_ = i[90] | i[89];
  assign t_1__36_ = i[91] | i[90];
  assign t_1__35_ = i[92] | i[91];
  assign t_1__34_ = i[93] | i[92];
  assign t_1__33_ = i[94] | i[93];
  assign t_1__32_ = i[95] | i[94];
  assign t_1__31_ = i[96] | i[95];
  assign t_1__30_ = i[97] | i[96];
  assign t_1__29_ = i[98] | i[97];
  assign t_1__28_ = i[99] | i[98];
  assign t_1__27_ = i[100] | i[99];
  assign t_1__26_ = i[101] | i[100];
  assign t_1__25_ = i[102] | i[101];
  assign t_1__24_ = i[103] | i[102];
  assign t_1__23_ = i[104] | i[103];
  assign t_1__22_ = i[105] | i[104];
  assign t_1__21_ = i[106] | i[105];
  assign t_1__20_ = i[107] | i[106];
  assign t_1__19_ = i[108] | i[107];
  assign t_1__18_ = i[109] | i[108];
  assign t_1__17_ = i[110] | i[109];
  assign t_1__16_ = i[111] | i[110];
  assign t_1__15_ = i[112] | i[111];
  assign t_1__14_ = i[113] | i[112];
  assign t_1__13_ = i[114] | i[113];
  assign t_1__12_ = i[115] | i[114];
  assign t_1__11_ = i[116] | i[115];
  assign t_1__10_ = i[117] | i[116];
  assign t_1__9_ = i[118] | i[117];
  assign t_1__8_ = i[119] | i[118];
  assign t_1__7_ = i[120] | i[119];
  assign t_1__6_ = i[121] | i[120];
  assign t_1__5_ = i[122] | i[121];
  assign t_1__4_ = i[123] | i[122];
  assign t_1__3_ = i[124] | i[123];
  assign t_1__2_ = i[125] | i[124];
  assign t_1__1_ = i[126] | i[125];
  assign t_1__0_ = i[127] | i[126];
  assign t_2__127_ = t_1__127_ | 1'b0;
  assign t_2__126_ = t_1__126_ | 1'b0;
  assign t_2__125_ = t_1__125_ | t_1__127_;
  assign t_2__124_ = t_1__124_ | t_1__126_;
  assign t_2__123_ = t_1__123_ | t_1__125_;
  assign t_2__122_ = t_1__122_ | t_1__124_;
  assign t_2__121_ = t_1__121_ | t_1__123_;
  assign t_2__120_ = t_1__120_ | t_1__122_;
  assign t_2__119_ = t_1__119_ | t_1__121_;
  assign t_2__118_ = t_1__118_ | t_1__120_;
  assign t_2__117_ = t_1__117_ | t_1__119_;
  assign t_2__116_ = t_1__116_ | t_1__118_;
  assign t_2__115_ = t_1__115_ | t_1__117_;
  assign t_2__114_ = t_1__114_ | t_1__116_;
  assign t_2__113_ = t_1__113_ | t_1__115_;
  assign t_2__112_ = t_1__112_ | t_1__114_;
  assign t_2__111_ = t_1__111_ | t_1__113_;
  assign t_2__110_ = t_1__110_ | t_1__112_;
  assign t_2__109_ = t_1__109_ | t_1__111_;
  assign t_2__108_ = t_1__108_ | t_1__110_;
  assign t_2__107_ = t_1__107_ | t_1__109_;
  assign t_2__106_ = t_1__106_ | t_1__108_;
  assign t_2__105_ = t_1__105_ | t_1__107_;
  assign t_2__104_ = t_1__104_ | t_1__106_;
  assign t_2__103_ = t_1__103_ | t_1__105_;
  assign t_2__102_ = t_1__102_ | t_1__104_;
  assign t_2__101_ = t_1__101_ | t_1__103_;
  assign t_2__100_ = t_1__100_ | t_1__102_;
  assign t_2__99_ = t_1__99_ | t_1__101_;
  assign t_2__98_ = t_1__98_ | t_1__100_;
  assign t_2__97_ = t_1__97_ | t_1__99_;
  assign t_2__96_ = t_1__96_ | t_1__98_;
  assign t_2__95_ = t_1__95_ | t_1__97_;
  assign t_2__94_ = t_1__94_ | t_1__96_;
  assign t_2__93_ = t_1__93_ | t_1__95_;
  assign t_2__92_ = t_1__92_ | t_1__94_;
  assign t_2__91_ = t_1__91_ | t_1__93_;
  assign t_2__90_ = t_1__90_ | t_1__92_;
  assign t_2__89_ = t_1__89_ | t_1__91_;
  assign t_2__88_ = t_1__88_ | t_1__90_;
  assign t_2__87_ = t_1__87_ | t_1__89_;
  assign t_2__86_ = t_1__86_ | t_1__88_;
  assign t_2__85_ = t_1__85_ | t_1__87_;
  assign t_2__84_ = t_1__84_ | t_1__86_;
  assign t_2__83_ = t_1__83_ | t_1__85_;
  assign t_2__82_ = t_1__82_ | t_1__84_;
  assign t_2__81_ = t_1__81_ | t_1__83_;
  assign t_2__80_ = t_1__80_ | t_1__82_;
  assign t_2__79_ = t_1__79_ | t_1__81_;
  assign t_2__78_ = t_1__78_ | t_1__80_;
  assign t_2__77_ = t_1__77_ | t_1__79_;
  assign t_2__76_ = t_1__76_ | t_1__78_;
  assign t_2__75_ = t_1__75_ | t_1__77_;
  assign t_2__74_ = t_1__74_ | t_1__76_;
  assign t_2__73_ = t_1__73_ | t_1__75_;
  assign t_2__72_ = t_1__72_ | t_1__74_;
  assign t_2__71_ = t_1__71_ | t_1__73_;
  assign t_2__70_ = t_1__70_ | t_1__72_;
  assign t_2__69_ = t_1__69_ | t_1__71_;
  assign t_2__68_ = t_1__68_ | t_1__70_;
  assign t_2__67_ = t_1__67_ | t_1__69_;
  assign t_2__66_ = t_1__66_ | t_1__68_;
  assign t_2__65_ = t_1__65_ | t_1__67_;
  assign t_2__64_ = t_1__64_ | t_1__66_;
  assign t_2__63_ = t_1__63_ | t_1__65_;
  assign t_2__62_ = t_1__62_ | t_1__64_;
  assign t_2__61_ = t_1__61_ | t_1__63_;
  assign t_2__60_ = t_1__60_ | t_1__62_;
  assign t_2__59_ = t_1__59_ | t_1__61_;
  assign t_2__58_ = t_1__58_ | t_1__60_;
  assign t_2__57_ = t_1__57_ | t_1__59_;
  assign t_2__56_ = t_1__56_ | t_1__58_;
  assign t_2__55_ = t_1__55_ | t_1__57_;
  assign t_2__54_ = t_1__54_ | t_1__56_;
  assign t_2__53_ = t_1__53_ | t_1__55_;
  assign t_2__52_ = t_1__52_ | t_1__54_;
  assign t_2__51_ = t_1__51_ | t_1__53_;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__127_ = t_2__127_ | 1'b0;
  assign t_3__126_ = t_2__126_ | 1'b0;
  assign t_3__125_ = t_2__125_ | 1'b0;
  assign t_3__124_ = t_2__124_ | 1'b0;
  assign t_3__123_ = t_2__123_ | t_2__127_;
  assign t_3__122_ = t_2__122_ | t_2__126_;
  assign t_3__121_ = t_2__121_ | t_2__125_;
  assign t_3__120_ = t_2__120_ | t_2__124_;
  assign t_3__119_ = t_2__119_ | t_2__123_;
  assign t_3__118_ = t_2__118_ | t_2__122_;
  assign t_3__117_ = t_2__117_ | t_2__121_;
  assign t_3__116_ = t_2__116_ | t_2__120_;
  assign t_3__115_ = t_2__115_ | t_2__119_;
  assign t_3__114_ = t_2__114_ | t_2__118_;
  assign t_3__113_ = t_2__113_ | t_2__117_;
  assign t_3__112_ = t_2__112_ | t_2__116_;
  assign t_3__111_ = t_2__111_ | t_2__115_;
  assign t_3__110_ = t_2__110_ | t_2__114_;
  assign t_3__109_ = t_2__109_ | t_2__113_;
  assign t_3__108_ = t_2__108_ | t_2__112_;
  assign t_3__107_ = t_2__107_ | t_2__111_;
  assign t_3__106_ = t_2__106_ | t_2__110_;
  assign t_3__105_ = t_2__105_ | t_2__109_;
  assign t_3__104_ = t_2__104_ | t_2__108_;
  assign t_3__103_ = t_2__103_ | t_2__107_;
  assign t_3__102_ = t_2__102_ | t_2__106_;
  assign t_3__101_ = t_2__101_ | t_2__105_;
  assign t_3__100_ = t_2__100_ | t_2__104_;
  assign t_3__99_ = t_2__99_ | t_2__103_;
  assign t_3__98_ = t_2__98_ | t_2__102_;
  assign t_3__97_ = t_2__97_ | t_2__101_;
  assign t_3__96_ = t_2__96_ | t_2__100_;
  assign t_3__95_ = t_2__95_ | t_2__99_;
  assign t_3__94_ = t_2__94_ | t_2__98_;
  assign t_3__93_ = t_2__93_ | t_2__97_;
  assign t_3__92_ = t_2__92_ | t_2__96_;
  assign t_3__91_ = t_2__91_ | t_2__95_;
  assign t_3__90_ = t_2__90_ | t_2__94_;
  assign t_3__89_ = t_2__89_ | t_2__93_;
  assign t_3__88_ = t_2__88_ | t_2__92_;
  assign t_3__87_ = t_2__87_ | t_2__91_;
  assign t_3__86_ = t_2__86_ | t_2__90_;
  assign t_3__85_ = t_2__85_ | t_2__89_;
  assign t_3__84_ = t_2__84_ | t_2__88_;
  assign t_3__83_ = t_2__83_ | t_2__87_;
  assign t_3__82_ = t_2__82_ | t_2__86_;
  assign t_3__81_ = t_2__81_ | t_2__85_;
  assign t_3__80_ = t_2__80_ | t_2__84_;
  assign t_3__79_ = t_2__79_ | t_2__83_;
  assign t_3__78_ = t_2__78_ | t_2__82_;
  assign t_3__77_ = t_2__77_ | t_2__81_;
  assign t_3__76_ = t_2__76_ | t_2__80_;
  assign t_3__75_ = t_2__75_ | t_2__79_;
  assign t_3__74_ = t_2__74_ | t_2__78_;
  assign t_3__73_ = t_2__73_ | t_2__77_;
  assign t_3__72_ = t_2__72_ | t_2__76_;
  assign t_3__71_ = t_2__71_ | t_2__75_;
  assign t_3__70_ = t_2__70_ | t_2__74_;
  assign t_3__69_ = t_2__69_ | t_2__73_;
  assign t_3__68_ = t_2__68_ | t_2__72_;
  assign t_3__67_ = t_2__67_ | t_2__71_;
  assign t_3__66_ = t_2__66_ | t_2__70_;
  assign t_3__65_ = t_2__65_ | t_2__69_;
  assign t_3__64_ = t_2__64_ | t_2__68_;
  assign t_3__63_ = t_2__63_ | t_2__67_;
  assign t_3__62_ = t_2__62_ | t_2__66_;
  assign t_3__61_ = t_2__61_ | t_2__65_;
  assign t_3__60_ = t_2__60_ | t_2__64_;
  assign t_3__59_ = t_2__59_ | t_2__63_;
  assign t_3__58_ = t_2__58_ | t_2__62_;
  assign t_3__57_ = t_2__57_ | t_2__61_;
  assign t_3__56_ = t_2__56_ | t_2__60_;
  assign t_3__55_ = t_2__55_ | t_2__59_;
  assign t_3__54_ = t_2__54_ | t_2__58_;
  assign t_3__53_ = t_2__53_ | t_2__57_;
  assign t_3__52_ = t_2__52_ | t_2__56_;
  assign t_3__51_ = t_2__51_ | t_2__55_;
  assign t_3__50_ = t_2__50_ | t_2__54_;
  assign t_3__49_ = t_2__49_ | t_2__53_;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__127_ = t_3__127_ | 1'b0;
  assign t_4__126_ = t_3__126_ | 1'b0;
  assign t_4__125_ = t_3__125_ | 1'b0;
  assign t_4__124_ = t_3__124_ | 1'b0;
  assign t_4__123_ = t_3__123_ | 1'b0;
  assign t_4__122_ = t_3__122_ | 1'b0;
  assign t_4__121_ = t_3__121_ | 1'b0;
  assign t_4__120_ = t_3__120_ | 1'b0;
  assign t_4__119_ = t_3__119_ | t_3__127_;
  assign t_4__118_ = t_3__118_ | t_3__126_;
  assign t_4__117_ = t_3__117_ | t_3__125_;
  assign t_4__116_ = t_3__116_ | t_3__124_;
  assign t_4__115_ = t_3__115_ | t_3__123_;
  assign t_4__114_ = t_3__114_ | t_3__122_;
  assign t_4__113_ = t_3__113_ | t_3__121_;
  assign t_4__112_ = t_3__112_ | t_3__120_;
  assign t_4__111_ = t_3__111_ | t_3__119_;
  assign t_4__110_ = t_3__110_ | t_3__118_;
  assign t_4__109_ = t_3__109_ | t_3__117_;
  assign t_4__108_ = t_3__108_ | t_3__116_;
  assign t_4__107_ = t_3__107_ | t_3__115_;
  assign t_4__106_ = t_3__106_ | t_3__114_;
  assign t_4__105_ = t_3__105_ | t_3__113_;
  assign t_4__104_ = t_3__104_ | t_3__112_;
  assign t_4__103_ = t_3__103_ | t_3__111_;
  assign t_4__102_ = t_3__102_ | t_3__110_;
  assign t_4__101_ = t_3__101_ | t_3__109_;
  assign t_4__100_ = t_3__100_ | t_3__108_;
  assign t_4__99_ = t_3__99_ | t_3__107_;
  assign t_4__98_ = t_3__98_ | t_3__106_;
  assign t_4__97_ = t_3__97_ | t_3__105_;
  assign t_4__96_ = t_3__96_ | t_3__104_;
  assign t_4__95_ = t_3__95_ | t_3__103_;
  assign t_4__94_ = t_3__94_ | t_3__102_;
  assign t_4__93_ = t_3__93_ | t_3__101_;
  assign t_4__92_ = t_3__92_ | t_3__100_;
  assign t_4__91_ = t_3__91_ | t_3__99_;
  assign t_4__90_ = t_3__90_ | t_3__98_;
  assign t_4__89_ = t_3__89_ | t_3__97_;
  assign t_4__88_ = t_3__88_ | t_3__96_;
  assign t_4__87_ = t_3__87_ | t_3__95_;
  assign t_4__86_ = t_3__86_ | t_3__94_;
  assign t_4__85_ = t_3__85_ | t_3__93_;
  assign t_4__84_ = t_3__84_ | t_3__92_;
  assign t_4__83_ = t_3__83_ | t_3__91_;
  assign t_4__82_ = t_3__82_ | t_3__90_;
  assign t_4__81_ = t_3__81_ | t_3__89_;
  assign t_4__80_ = t_3__80_ | t_3__88_;
  assign t_4__79_ = t_3__79_ | t_3__87_;
  assign t_4__78_ = t_3__78_ | t_3__86_;
  assign t_4__77_ = t_3__77_ | t_3__85_;
  assign t_4__76_ = t_3__76_ | t_3__84_;
  assign t_4__75_ = t_3__75_ | t_3__83_;
  assign t_4__74_ = t_3__74_ | t_3__82_;
  assign t_4__73_ = t_3__73_ | t_3__81_;
  assign t_4__72_ = t_3__72_ | t_3__80_;
  assign t_4__71_ = t_3__71_ | t_3__79_;
  assign t_4__70_ = t_3__70_ | t_3__78_;
  assign t_4__69_ = t_3__69_ | t_3__77_;
  assign t_4__68_ = t_3__68_ | t_3__76_;
  assign t_4__67_ = t_3__67_ | t_3__75_;
  assign t_4__66_ = t_3__66_ | t_3__74_;
  assign t_4__65_ = t_3__65_ | t_3__73_;
  assign t_4__64_ = t_3__64_ | t_3__72_;
  assign t_4__63_ = t_3__63_ | t_3__71_;
  assign t_4__62_ = t_3__62_ | t_3__70_;
  assign t_4__61_ = t_3__61_ | t_3__69_;
  assign t_4__60_ = t_3__60_ | t_3__68_;
  assign t_4__59_ = t_3__59_ | t_3__67_;
  assign t_4__58_ = t_3__58_ | t_3__66_;
  assign t_4__57_ = t_3__57_ | t_3__65_;
  assign t_4__56_ = t_3__56_ | t_3__64_;
  assign t_4__55_ = t_3__55_ | t_3__63_;
  assign t_4__54_ = t_3__54_ | t_3__62_;
  assign t_4__53_ = t_3__53_ | t_3__61_;
  assign t_4__52_ = t_3__52_ | t_3__60_;
  assign t_4__51_ = t_3__51_ | t_3__59_;
  assign t_4__50_ = t_3__50_ | t_3__58_;
  assign t_4__49_ = t_3__49_ | t_3__57_;
  assign t_4__48_ = t_3__48_ | t_3__56_;
  assign t_4__47_ = t_3__47_ | t_3__55_;
  assign t_4__46_ = t_3__46_ | t_3__54_;
  assign t_4__45_ = t_3__45_ | t_3__53_;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__127_ = t_4__127_ | 1'b0;
  assign t_5__126_ = t_4__126_ | 1'b0;
  assign t_5__125_ = t_4__125_ | 1'b0;
  assign t_5__124_ = t_4__124_ | 1'b0;
  assign t_5__123_ = t_4__123_ | 1'b0;
  assign t_5__122_ = t_4__122_ | 1'b0;
  assign t_5__121_ = t_4__121_ | 1'b0;
  assign t_5__120_ = t_4__120_ | 1'b0;
  assign t_5__119_ = t_4__119_ | 1'b0;
  assign t_5__118_ = t_4__118_ | 1'b0;
  assign t_5__117_ = t_4__117_ | 1'b0;
  assign t_5__116_ = t_4__116_ | 1'b0;
  assign t_5__115_ = t_4__115_ | 1'b0;
  assign t_5__114_ = t_4__114_ | 1'b0;
  assign t_5__113_ = t_4__113_ | 1'b0;
  assign t_5__112_ = t_4__112_ | 1'b0;
  assign t_5__111_ = t_4__111_ | t_4__127_;
  assign t_5__110_ = t_4__110_ | t_4__126_;
  assign t_5__109_ = t_4__109_ | t_4__125_;
  assign t_5__108_ = t_4__108_ | t_4__124_;
  assign t_5__107_ = t_4__107_ | t_4__123_;
  assign t_5__106_ = t_4__106_ | t_4__122_;
  assign t_5__105_ = t_4__105_ | t_4__121_;
  assign t_5__104_ = t_4__104_ | t_4__120_;
  assign t_5__103_ = t_4__103_ | t_4__119_;
  assign t_5__102_ = t_4__102_ | t_4__118_;
  assign t_5__101_ = t_4__101_ | t_4__117_;
  assign t_5__100_ = t_4__100_ | t_4__116_;
  assign t_5__99_ = t_4__99_ | t_4__115_;
  assign t_5__98_ = t_4__98_ | t_4__114_;
  assign t_5__97_ = t_4__97_ | t_4__113_;
  assign t_5__96_ = t_4__96_ | t_4__112_;
  assign t_5__95_ = t_4__95_ | t_4__111_;
  assign t_5__94_ = t_4__94_ | t_4__110_;
  assign t_5__93_ = t_4__93_ | t_4__109_;
  assign t_5__92_ = t_4__92_ | t_4__108_;
  assign t_5__91_ = t_4__91_ | t_4__107_;
  assign t_5__90_ = t_4__90_ | t_4__106_;
  assign t_5__89_ = t_4__89_ | t_4__105_;
  assign t_5__88_ = t_4__88_ | t_4__104_;
  assign t_5__87_ = t_4__87_ | t_4__103_;
  assign t_5__86_ = t_4__86_ | t_4__102_;
  assign t_5__85_ = t_4__85_ | t_4__101_;
  assign t_5__84_ = t_4__84_ | t_4__100_;
  assign t_5__83_ = t_4__83_ | t_4__99_;
  assign t_5__82_ = t_4__82_ | t_4__98_;
  assign t_5__81_ = t_4__81_ | t_4__97_;
  assign t_5__80_ = t_4__80_ | t_4__96_;
  assign t_5__79_ = t_4__79_ | t_4__95_;
  assign t_5__78_ = t_4__78_ | t_4__94_;
  assign t_5__77_ = t_4__77_ | t_4__93_;
  assign t_5__76_ = t_4__76_ | t_4__92_;
  assign t_5__75_ = t_4__75_ | t_4__91_;
  assign t_5__74_ = t_4__74_ | t_4__90_;
  assign t_5__73_ = t_4__73_ | t_4__89_;
  assign t_5__72_ = t_4__72_ | t_4__88_;
  assign t_5__71_ = t_4__71_ | t_4__87_;
  assign t_5__70_ = t_4__70_ | t_4__86_;
  assign t_5__69_ = t_4__69_ | t_4__85_;
  assign t_5__68_ = t_4__68_ | t_4__84_;
  assign t_5__67_ = t_4__67_ | t_4__83_;
  assign t_5__66_ = t_4__66_ | t_4__82_;
  assign t_5__65_ = t_4__65_ | t_4__81_;
  assign t_5__64_ = t_4__64_ | t_4__80_;
  assign t_5__63_ = t_4__63_ | t_4__79_;
  assign t_5__62_ = t_4__62_ | t_4__78_;
  assign t_5__61_ = t_4__61_ | t_4__77_;
  assign t_5__60_ = t_4__60_ | t_4__76_;
  assign t_5__59_ = t_4__59_ | t_4__75_;
  assign t_5__58_ = t_4__58_ | t_4__74_;
  assign t_5__57_ = t_4__57_ | t_4__73_;
  assign t_5__56_ = t_4__56_ | t_4__72_;
  assign t_5__55_ = t_4__55_ | t_4__71_;
  assign t_5__54_ = t_4__54_ | t_4__70_;
  assign t_5__53_ = t_4__53_ | t_4__69_;
  assign t_5__52_ = t_4__52_ | t_4__68_;
  assign t_5__51_ = t_4__51_ | t_4__67_;
  assign t_5__50_ = t_4__50_ | t_4__66_;
  assign t_5__49_ = t_4__49_ | t_4__65_;
  assign t_5__48_ = t_4__48_ | t_4__64_;
  assign t_5__47_ = t_4__47_ | t_4__63_;
  assign t_5__46_ = t_4__46_ | t_4__62_;
  assign t_5__45_ = t_4__45_ | t_4__61_;
  assign t_5__44_ = t_4__44_ | t_4__60_;
  assign t_5__43_ = t_4__43_ | t_4__59_;
  assign t_5__42_ = t_4__42_ | t_4__58_;
  assign t_5__41_ = t_4__41_ | t_4__57_;
  assign t_5__40_ = t_4__40_ | t_4__56_;
  assign t_5__39_ = t_4__39_ | t_4__55_;
  assign t_5__38_ = t_4__38_ | t_4__54_;
  assign t_5__37_ = t_4__37_ | t_4__53_;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign t_6__127_ = t_5__127_ | 1'b0;
  assign t_6__126_ = t_5__126_ | 1'b0;
  assign t_6__125_ = t_5__125_ | 1'b0;
  assign t_6__124_ = t_5__124_ | 1'b0;
  assign t_6__123_ = t_5__123_ | 1'b0;
  assign t_6__122_ = t_5__122_ | 1'b0;
  assign t_6__121_ = t_5__121_ | 1'b0;
  assign t_6__120_ = t_5__120_ | 1'b0;
  assign t_6__119_ = t_5__119_ | 1'b0;
  assign t_6__118_ = t_5__118_ | 1'b0;
  assign t_6__117_ = t_5__117_ | 1'b0;
  assign t_6__116_ = t_5__116_ | 1'b0;
  assign t_6__115_ = t_5__115_ | 1'b0;
  assign t_6__114_ = t_5__114_ | 1'b0;
  assign t_6__113_ = t_5__113_ | 1'b0;
  assign t_6__112_ = t_5__112_ | 1'b0;
  assign t_6__111_ = t_5__111_ | 1'b0;
  assign t_6__110_ = t_5__110_ | 1'b0;
  assign t_6__109_ = t_5__109_ | 1'b0;
  assign t_6__108_ = t_5__108_ | 1'b0;
  assign t_6__107_ = t_5__107_ | 1'b0;
  assign t_6__106_ = t_5__106_ | 1'b0;
  assign t_6__105_ = t_5__105_ | 1'b0;
  assign t_6__104_ = t_5__104_ | 1'b0;
  assign t_6__103_ = t_5__103_ | 1'b0;
  assign t_6__102_ = t_5__102_ | 1'b0;
  assign t_6__101_ = t_5__101_ | 1'b0;
  assign t_6__100_ = t_5__100_ | 1'b0;
  assign t_6__99_ = t_5__99_ | 1'b0;
  assign t_6__98_ = t_5__98_ | 1'b0;
  assign t_6__97_ = t_5__97_ | 1'b0;
  assign t_6__96_ = t_5__96_ | 1'b0;
  assign t_6__95_ = t_5__95_ | t_5__127_;
  assign t_6__94_ = t_5__94_ | t_5__126_;
  assign t_6__93_ = t_5__93_ | t_5__125_;
  assign t_6__92_ = t_5__92_ | t_5__124_;
  assign t_6__91_ = t_5__91_ | t_5__123_;
  assign t_6__90_ = t_5__90_ | t_5__122_;
  assign t_6__89_ = t_5__89_ | t_5__121_;
  assign t_6__88_ = t_5__88_ | t_5__120_;
  assign t_6__87_ = t_5__87_ | t_5__119_;
  assign t_6__86_ = t_5__86_ | t_5__118_;
  assign t_6__85_ = t_5__85_ | t_5__117_;
  assign t_6__84_ = t_5__84_ | t_5__116_;
  assign t_6__83_ = t_5__83_ | t_5__115_;
  assign t_6__82_ = t_5__82_ | t_5__114_;
  assign t_6__81_ = t_5__81_ | t_5__113_;
  assign t_6__80_ = t_5__80_ | t_5__112_;
  assign t_6__79_ = t_5__79_ | t_5__111_;
  assign t_6__78_ = t_5__78_ | t_5__110_;
  assign t_6__77_ = t_5__77_ | t_5__109_;
  assign t_6__76_ = t_5__76_ | t_5__108_;
  assign t_6__75_ = t_5__75_ | t_5__107_;
  assign t_6__74_ = t_5__74_ | t_5__106_;
  assign t_6__73_ = t_5__73_ | t_5__105_;
  assign t_6__72_ = t_5__72_ | t_5__104_;
  assign t_6__71_ = t_5__71_ | t_5__103_;
  assign t_6__70_ = t_5__70_ | t_5__102_;
  assign t_6__69_ = t_5__69_ | t_5__101_;
  assign t_6__68_ = t_5__68_ | t_5__100_;
  assign t_6__67_ = t_5__67_ | t_5__99_;
  assign t_6__66_ = t_5__66_ | t_5__98_;
  assign t_6__65_ = t_5__65_ | t_5__97_;
  assign t_6__64_ = t_5__64_ | t_5__96_;
  assign t_6__63_ = t_5__63_ | t_5__95_;
  assign t_6__62_ = t_5__62_ | t_5__94_;
  assign t_6__61_ = t_5__61_ | t_5__93_;
  assign t_6__60_ = t_5__60_ | t_5__92_;
  assign t_6__59_ = t_5__59_ | t_5__91_;
  assign t_6__58_ = t_5__58_ | t_5__90_;
  assign t_6__57_ = t_5__57_ | t_5__89_;
  assign t_6__56_ = t_5__56_ | t_5__88_;
  assign t_6__55_ = t_5__55_ | t_5__87_;
  assign t_6__54_ = t_5__54_ | t_5__86_;
  assign t_6__53_ = t_5__53_ | t_5__85_;
  assign t_6__52_ = t_5__52_ | t_5__84_;
  assign t_6__51_ = t_5__51_ | t_5__83_;
  assign t_6__50_ = t_5__50_ | t_5__82_;
  assign t_6__49_ = t_5__49_ | t_5__81_;
  assign t_6__48_ = t_5__48_ | t_5__80_;
  assign t_6__47_ = t_5__47_ | t_5__79_;
  assign t_6__46_ = t_5__46_ | t_5__78_;
  assign t_6__45_ = t_5__45_ | t_5__77_;
  assign t_6__44_ = t_5__44_ | t_5__76_;
  assign t_6__43_ = t_5__43_ | t_5__75_;
  assign t_6__42_ = t_5__42_ | t_5__74_;
  assign t_6__41_ = t_5__41_ | t_5__73_;
  assign t_6__40_ = t_5__40_ | t_5__72_;
  assign t_6__39_ = t_5__39_ | t_5__71_;
  assign t_6__38_ = t_5__38_ | t_5__70_;
  assign t_6__37_ = t_5__37_ | t_5__69_;
  assign t_6__36_ = t_5__36_ | t_5__68_;
  assign t_6__35_ = t_5__35_ | t_5__67_;
  assign t_6__34_ = t_5__34_ | t_5__66_;
  assign t_6__33_ = t_5__33_ | t_5__65_;
  assign t_6__32_ = t_5__32_ | t_5__64_;
  assign t_6__31_ = t_5__31_ | t_5__63_;
  assign t_6__30_ = t_5__30_ | t_5__62_;
  assign t_6__29_ = t_5__29_ | t_5__61_;
  assign t_6__28_ = t_5__28_ | t_5__60_;
  assign t_6__27_ = t_5__27_ | t_5__59_;
  assign t_6__26_ = t_5__26_ | t_5__58_;
  assign t_6__25_ = t_5__25_ | t_5__57_;
  assign t_6__24_ = t_5__24_ | t_5__56_;
  assign t_6__23_ = t_5__23_ | t_5__55_;
  assign t_6__22_ = t_5__22_ | t_5__54_;
  assign t_6__21_ = t_5__21_ | t_5__53_;
  assign t_6__20_ = t_5__20_ | t_5__52_;
  assign t_6__19_ = t_5__19_ | t_5__51_;
  assign t_6__18_ = t_5__18_ | t_5__50_;
  assign t_6__17_ = t_5__17_ | t_5__49_;
  assign t_6__16_ = t_5__16_ | t_5__48_;
  assign t_6__15_ = t_5__15_ | t_5__47_;
  assign t_6__14_ = t_5__14_ | t_5__46_;
  assign t_6__13_ = t_5__13_ | t_5__45_;
  assign t_6__12_ = t_5__12_ | t_5__44_;
  assign t_6__11_ = t_5__11_ | t_5__43_;
  assign t_6__10_ = t_5__10_ | t_5__42_;
  assign t_6__9_ = t_5__9_ | t_5__41_;
  assign t_6__8_ = t_5__8_ | t_5__40_;
  assign t_6__7_ = t_5__7_ | t_5__39_;
  assign t_6__6_ = t_5__6_ | t_5__38_;
  assign t_6__5_ = t_5__5_ | t_5__37_;
  assign t_6__4_ = t_5__4_ | t_5__36_;
  assign t_6__3_ = t_5__3_ | t_5__35_;
  assign t_6__2_ = t_5__2_ | t_5__34_;
  assign t_6__1_ = t_5__1_ | t_5__33_;
  assign t_6__0_ = t_5__0_ | t_5__32_;
  assign o[0] = t_6__127_ | 1'b0;
  assign o[1] = t_6__126_ | 1'b0;
  assign o[2] = t_6__125_ | 1'b0;
  assign o[3] = t_6__124_ | 1'b0;
  assign o[4] = t_6__123_ | 1'b0;
  assign o[5] = t_6__122_ | 1'b0;
  assign o[6] = t_6__121_ | 1'b0;
  assign o[7] = t_6__120_ | 1'b0;
  assign o[8] = t_6__119_ | 1'b0;
  assign o[9] = t_6__118_ | 1'b0;
  assign o[10] = t_6__117_ | 1'b0;
  assign o[11] = t_6__116_ | 1'b0;
  assign o[12] = t_6__115_ | 1'b0;
  assign o[13] = t_6__114_ | 1'b0;
  assign o[14] = t_6__113_ | 1'b0;
  assign o[15] = t_6__112_ | 1'b0;
  assign o[16] = t_6__111_ | 1'b0;
  assign o[17] = t_6__110_ | 1'b0;
  assign o[18] = t_6__109_ | 1'b0;
  assign o[19] = t_6__108_ | 1'b0;
  assign o[20] = t_6__107_ | 1'b0;
  assign o[21] = t_6__106_ | 1'b0;
  assign o[22] = t_6__105_ | 1'b0;
  assign o[23] = t_6__104_ | 1'b0;
  assign o[24] = t_6__103_ | 1'b0;
  assign o[25] = t_6__102_ | 1'b0;
  assign o[26] = t_6__101_ | 1'b0;
  assign o[27] = t_6__100_ | 1'b0;
  assign o[28] = t_6__99_ | 1'b0;
  assign o[29] = t_6__98_ | 1'b0;
  assign o[30] = t_6__97_ | 1'b0;
  assign o[31] = t_6__96_ | 1'b0;
  assign o[32] = t_6__95_ | 1'b0;
  assign o[33] = t_6__94_ | 1'b0;
  assign o[34] = t_6__93_ | 1'b0;
  assign o[35] = t_6__92_ | 1'b0;
  assign o[36] = t_6__91_ | 1'b0;
  assign o[37] = t_6__90_ | 1'b0;
  assign o[38] = t_6__89_ | 1'b0;
  assign o[39] = t_6__88_ | 1'b0;
  assign o[40] = t_6__87_ | 1'b0;
  assign o[41] = t_6__86_ | 1'b0;
  assign o[42] = t_6__85_ | 1'b0;
  assign o[43] = t_6__84_ | 1'b0;
  assign o[44] = t_6__83_ | 1'b0;
  assign o[45] = t_6__82_ | 1'b0;
  assign o[46] = t_6__81_ | 1'b0;
  assign o[47] = t_6__80_ | 1'b0;
  assign o[48] = t_6__79_ | 1'b0;
  assign o[49] = t_6__78_ | 1'b0;
  assign o[50] = t_6__77_ | 1'b0;
  assign o[51] = t_6__76_ | 1'b0;
  assign o[52] = t_6__75_ | 1'b0;
  assign o[53] = t_6__74_ | 1'b0;
  assign o[54] = t_6__73_ | 1'b0;
  assign o[55] = t_6__72_ | 1'b0;
  assign o[56] = t_6__71_ | 1'b0;
  assign o[57] = t_6__70_ | 1'b0;
  assign o[58] = t_6__69_ | 1'b0;
  assign o[59] = t_6__68_ | 1'b0;
  assign o[60] = t_6__67_ | 1'b0;
  assign o[61] = t_6__66_ | 1'b0;
  assign o[62] = t_6__65_ | 1'b0;
  assign o[63] = t_6__64_ | 1'b0;
  assign o[64] = t_6__63_ | t_6__127_;
  assign o[65] = t_6__62_ | t_6__126_;
  assign o[66] = t_6__61_ | t_6__125_;
  assign o[67] = t_6__60_ | t_6__124_;
  assign o[68] = t_6__59_ | t_6__123_;
  assign o[69] = t_6__58_ | t_6__122_;
  assign o[70] = t_6__57_ | t_6__121_;
  assign o[71] = t_6__56_ | t_6__120_;
  assign o[72] = t_6__55_ | t_6__119_;
  assign o[73] = t_6__54_ | t_6__118_;
  assign o[74] = t_6__53_ | t_6__117_;
  assign o[75] = t_6__52_ | t_6__116_;
  assign o[76] = t_6__51_ | t_6__115_;
  assign o[77] = t_6__50_ | t_6__114_;
  assign o[78] = t_6__49_ | t_6__113_;
  assign o[79] = t_6__48_ | t_6__112_;
  assign o[80] = t_6__47_ | t_6__111_;
  assign o[81] = t_6__46_ | t_6__110_;
  assign o[82] = t_6__45_ | t_6__109_;
  assign o[83] = t_6__44_ | t_6__108_;
  assign o[84] = t_6__43_ | t_6__107_;
  assign o[85] = t_6__42_ | t_6__106_;
  assign o[86] = t_6__41_ | t_6__105_;
  assign o[87] = t_6__40_ | t_6__104_;
  assign o[88] = t_6__39_ | t_6__103_;
  assign o[89] = t_6__38_ | t_6__102_;
  assign o[90] = t_6__37_ | t_6__101_;
  assign o[91] = t_6__36_ | t_6__100_;
  assign o[92] = t_6__35_ | t_6__99_;
  assign o[93] = t_6__34_ | t_6__98_;
  assign o[94] = t_6__33_ | t_6__97_;
  assign o[95] = t_6__32_ | t_6__96_;
  assign o[96] = t_6__31_ | t_6__95_;
  assign o[97] = t_6__30_ | t_6__94_;
  assign o[98] = t_6__29_ | t_6__93_;
  assign o[99] = t_6__28_ | t_6__92_;
  assign o[100] = t_6__27_ | t_6__91_;
  assign o[101] = t_6__26_ | t_6__90_;
  assign o[102] = t_6__25_ | t_6__89_;
  assign o[103] = t_6__24_ | t_6__88_;
  assign o[104] = t_6__23_ | t_6__87_;
  assign o[105] = t_6__22_ | t_6__86_;
  assign o[106] = t_6__21_ | t_6__85_;
  assign o[107] = t_6__20_ | t_6__84_;
  assign o[108] = t_6__19_ | t_6__83_;
  assign o[109] = t_6__18_ | t_6__82_;
  assign o[110] = t_6__17_ | t_6__81_;
  assign o[111] = t_6__16_ | t_6__80_;
  assign o[112] = t_6__15_ | t_6__79_;
  assign o[113] = t_6__14_ | t_6__78_;
  assign o[114] = t_6__13_ | t_6__77_;
  assign o[115] = t_6__12_ | t_6__76_;
  assign o[116] = t_6__11_ | t_6__75_;
  assign o[117] = t_6__10_ | t_6__74_;
  assign o[118] = t_6__9_ | t_6__73_;
  assign o[119] = t_6__8_ | t_6__72_;
  assign o[120] = t_6__7_ | t_6__71_;
  assign o[121] = t_6__6_ | t_6__70_;
  assign o[122] = t_6__5_ | t_6__69_;
  assign o[123] = t_6__4_ | t_6__68_;
  assign o[124] = t_6__3_ | t_6__67_;
  assign o[125] = t_6__2_ | t_6__66_;
  assign o[126] = t_6__1_ | t_6__65_;
  assign o[127] = t_6__0_ | t_6__64_;

endmodule



module bsg_priority_encode_one_hot_out_width_p128_lo_to_hi_p1
(
  i,
  o
);

  input [127:0] i;
  output [127:0] o;
  wire [127:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126;
  wire [127:1] scan_lo;

  bsg_scan_width_p128_or_p1_lo_to_hi_p1
  genblk1_scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[127] = scan_lo[127] & N0;
  assign N0 = ~scan_lo[126];
  assign o[126] = scan_lo[126] & N1;
  assign N1 = ~scan_lo[125];
  assign o[125] = scan_lo[125] & N2;
  assign N2 = ~scan_lo[124];
  assign o[124] = scan_lo[124] & N3;
  assign N3 = ~scan_lo[123];
  assign o[123] = scan_lo[123] & N4;
  assign N4 = ~scan_lo[122];
  assign o[122] = scan_lo[122] & N5;
  assign N5 = ~scan_lo[121];
  assign o[121] = scan_lo[121] & N6;
  assign N6 = ~scan_lo[120];
  assign o[120] = scan_lo[120] & N7;
  assign N7 = ~scan_lo[119];
  assign o[119] = scan_lo[119] & N8;
  assign N8 = ~scan_lo[118];
  assign o[118] = scan_lo[118] & N9;
  assign N9 = ~scan_lo[117];
  assign o[117] = scan_lo[117] & N10;
  assign N10 = ~scan_lo[116];
  assign o[116] = scan_lo[116] & N11;
  assign N11 = ~scan_lo[115];
  assign o[115] = scan_lo[115] & N12;
  assign N12 = ~scan_lo[114];
  assign o[114] = scan_lo[114] & N13;
  assign N13 = ~scan_lo[113];
  assign o[113] = scan_lo[113] & N14;
  assign N14 = ~scan_lo[112];
  assign o[112] = scan_lo[112] & N15;
  assign N15 = ~scan_lo[111];
  assign o[111] = scan_lo[111] & N16;
  assign N16 = ~scan_lo[110];
  assign o[110] = scan_lo[110] & N17;
  assign N17 = ~scan_lo[109];
  assign o[109] = scan_lo[109] & N18;
  assign N18 = ~scan_lo[108];
  assign o[108] = scan_lo[108] & N19;
  assign N19 = ~scan_lo[107];
  assign o[107] = scan_lo[107] & N20;
  assign N20 = ~scan_lo[106];
  assign o[106] = scan_lo[106] & N21;
  assign N21 = ~scan_lo[105];
  assign o[105] = scan_lo[105] & N22;
  assign N22 = ~scan_lo[104];
  assign o[104] = scan_lo[104] & N23;
  assign N23 = ~scan_lo[103];
  assign o[103] = scan_lo[103] & N24;
  assign N24 = ~scan_lo[102];
  assign o[102] = scan_lo[102] & N25;
  assign N25 = ~scan_lo[101];
  assign o[101] = scan_lo[101] & N26;
  assign N26 = ~scan_lo[100];
  assign o[100] = scan_lo[100] & N27;
  assign N27 = ~scan_lo[99];
  assign o[99] = scan_lo[99] & N28;
  assign N28 = ~scan_lo[98];
  assign o[98] = scan_lo[98] & N29;
  assign N29 = ~scan_lo[97];
  assign o[97] = scan_lo[97] & N30;
  assign N30 = ~scan_lo[96];
  assign o[96] = scan_lo[96] & N31;
  assign N31 = ~scan_lo[95];
  assign o[95] = scan_lo[95] & N32;
  assign N32 = ~scan_lo[94];
  assign o[94] = scan_lo[94] & N33;
  assign N33 = ~scan_lo[93];
  assign o[93] = scan_lo[93] & N34;
  assign N34 = ~scan_lo[92];
  assign o[92] = scan_lo[92] & N35;
  assign N35 = ~scan_lo[91];
  assign o[91] = scan_lo[91] & N36;
  assign N36 = ~scan_lo[90];
  assign o[90] = scan_lo[90] & N37;
  assign N37 = ~scan_lo[89];
  assign o[89] = scan_lo[89] & N38;
  assign N38 = ~scan_lo[88];
  assign o[88] = scan_lo[88] & N39;
  assign N39 = ~scan_lo[87];
  assign o[87] = scan_lo[87] & N40;
  assign N40 = ~scan_lo[86];
  assign o[86] = scan_lo[86] & N41;
  assign N41 = ~scan_lo[85];
  assign o[85] = scan_lo[85] & N42;
  assign N42 = ~scan_lo[84];
  assign o[84] = scan_lo[84] & N43;
  assign N43 = ~scan_lo[83];
  assign o[83] = scan_lo[83] & N44;
  assign N44 = ~scan_lo[82];
  assign o[82] = scan_lo[82] & N45;
  assign N45 = ~scan_lo[81];
  assign o[81] = scan_lo[81] & N46;
  assign N46 = ~scan_lo[80];
  assign o[80] = scan_lo[80] & N47;
  assign N47 = ~scan_lo[79];
  assign o[79] = scan_lo[79] & N48;
  assign N48 = ~scan_lo[78];
  assign o[78] = scan_lo[78] & N49;
  assign N49 = ~scan_lo[77];
  assign o[77] = scan_lo[77] & N50;
  assign N50 = ~scan_lo[76];
  assign o[76] = scan_lo[76] & N51;
  assign N51 = ~scan_lo[75];
  assign o[75] = scan_lo[75] & N52;
  assign N52 = ~scan_lo[74];
  assign o[74] = scan_lo[74] & N53;
  assign N53 = ~scan_lo[73];
  assign o[73] = scan_lo[73] & N54;
  assign N54 = ~scan_lo[72];
  assign o[72] = scan_lo[72] & N55;
  assign N55 = ~scan_lo[71];
  assign o[71] = scan_lo[71] & N56;
  assign N56 = ~scan_lo[70];
  assign o[70] = scan_lo[70] & N57;
  assign N57 = ~scan_lo[69];
  assign o[69] = scan_lo[69] & N58;
  assign N58 = ~scan_lo[68];
  assign o[68] = scan_lo[68] & N59;
  assign N59 = ~scan_lo[67];
  assign o[67] = scan_lo[67] & N60;
  assign N60 = ~scan_lo[66];
  assign o[66] = scan_lo[66] & N61;
  assign N61 = ~scan_lo[65];
  assign o[65] = scan_lo[65] & N62;
  assign N62 = ~scan_lo[64];
  assign o[64] = scan_lo[64] & N63;
  assign N63 = ~scan_lo[63];
  assign o[63] = scan_lo[63] & N64;
  assign N64 = ~scan_lo[62];
  assign o[62] = scan_lo[62] & N65;
  assign N65 = ~scan_lo[61];
  assign o[61] = scan_lo[61] & N66;
  assign N66 = ~scan_lo[60];
  assign o[60] = scan_lo[60] & N67;
  assign N67 = ~scan_lo[59];
  assign o[59] = scan_lo[59] & N68;
  assign N68 = ~scan_lo[58];
  assign o[58] = scan_lo[58] & N69;
  assign N69 = ~scan_lo[57];
  assign o[57] = scan_lo[57] & N70;
  assign N70 = ~scan_lo[56];
  assign o[56] = scan_lo[56] & N71;
  assign N71 = ~scan_lo[55];
  assign o[55] = scan_lo[55] & N72;
  assign N72 = ~scan_lo[54];
  assign o[54] = scan_lo[54] & N73;
  assign N73 = ~scan_lo[53];
  assign o[53] = scan_lo[53] & N74;
  assign N74 = ~scan_lo[52];
  assign o[52] = scan_lo[52] & N75;
  assign N75 = ~scan_lo[51];
  assign o[51] = scan_lo[51] & N76;
  assign N76 = ~scan_lo[50];
  assign o[50] = scan_lo[50] & N77;
  assign N77 = ~scan_lo[49];
  assign o[49] = scan_lo[49] & N78;
  assign N78 = ~scan_lo[48];
  assign o[48] = scan_lo[48] & N79;
  assign N79 = ~scan_lo[47];
  assign o[47] = scan_lo[47] & N80;
  assign N80 = ~scan_lo[46];
  assign o[46] = scan_lo[46] & N81;
  assign N81 = ~scan_lo[45];
  assign o[45] = scan_lo[45] & N82;
  assign N82 = ~scan_lo[44];
  assign o[44] = scan_lo[44] & N83;
  assign N83 = ~scan_lo[43];
  assign o[43] = scan_lo[43] & N84;
  assign N84 = ~scan_lo[42];
  assign o[42] = scan_lo[42] & N85;
  assign N85 = ~scan_lo[41];
  assign o[41] = scan_lo[41] & N86;
  assign N86 = ~scan_lo[40];
  assign o[40] = scan_lo[40] & N87;
  assign N87 = ~scan_lo[39];
  assign o[39] = scan_lo[39] & N88;
  assign N88 = ~scan_lo[38];
  assign o[38] = scan_lo[38] & N89;
  assign N89 = ~scan_lo[37];
  assign o[37] = scan_lo[37] & N90;
  assign N90 = ~scan_lo[36];
  assign o[36] = scan_lo[36] & N91;
  assign N91 = ~scan_lo[35];
  assign o[35] = scan_lo[35] & N92;
  assign N92 = ~scan_lo[34];
  assign o[34] = scan_lo[34] & N93;
  assign N93 = ~scan_lo[33];
  assign o[33] = scan_lo[33] & N94;
  assign N94 = ~scan_lo[32];
  assign o[32] = scan_lo[32] & N95;
  assign N95 = ~scan_lo[31];
  assign o[31] = scan_lo[31] & N96;
  assign N96 = ~scan_lo[30];
  assign o[30] = scan_lo[30] & N97;
  assign N97 = ~scan_lo[29];
  assign o[29] = scan_lo[29] & N98;
  assign N98 = ~scan_lo[28];
  assign o[28] = scan_lo[28] & N99;
  assign N99 = ~scan_lo[27];
  assign o[27] = scan_lo[27] & N100;
  assign N100 = ~scan_lo[26];
  assign o[26] = scan_lo[26] & N101;
  assign N101 = ~scan_lo[25];
  assign o[25] = scan_lo[25] & N102;
  assign N102 = ~scan_lo[24];
  assign o[24] = scan_lo[24] & N103;
  assign N103 = ~scan_lo[23];
  assign o[23] = scan_lo[23] & N104;
  assign N104 = ~scan_lo[22];
  assign o[22] = scan_lo[22] & N105;
  assign N105 = ~scan_lo[21];
  assign o[21] = scan_lo[21] & N106;
  assign N106 = ~scan_lo[20];
  assign o[20] = scan_lo[20] & N107;
  assign N107 = ~scan_lo[19];
  assign o[19] = scan_lo[19] & N108;
  assign N108 = ~scan_lo[18];
  assign o[18] = scan_lo[18] & N109;
  assign N109 = ~scan_lo[17];
  assign o[17] = scan_lo[17] & N110;
  assign N110 = ~scan_lo[16];
  assign o[16] = scan_lo[16] & N111;
  assign N111 = ~scan_lo[15];
  assign o[15] = scan_lo[15] & N112;
  assign N112 = ~scan_lo[14];
  assign o[14] = scan_lo[14] & N113;
  assign N113 = ~scan_lo[13];
  assign o[13] = scan_lo[13] & N114;
  assign N114 = ~scan_lo[12];
  assign o[12] = scan_lo[12] & N115;
  assign N115 = ~scan_lo[11];
  assign o[11] = scan_lo[11] & N116;
  assign N116 = ~scan_lo[10];
  assign o[10] = scan_lo[10] & N117;
  assign N117 = ~scan_lo[9];
  assign o[9] = scan_lo[9] & N118;
  assign N118 = ~scan_lo[8];
  assign o[8] = scan_lo[8] & N119;
  assign N119 = ~scan_lo[7];
  assign o[7] = scan_lo[7] & N120;
  assign N120 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N121;
  assign N121 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N122;
  assign N122 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N123;
  assign N123 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N124;
  assign N124 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N125;
  assign N125 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N126;
  assign N126 = ~o[0];

endmodule



module bsg_arb_fixed
(
  ready_i,
  reqs_i,
  grants_o
);

  input [127:0] reqs_i;
  output [127:0] grants_o;
  input ready_i;
  wire [127:0] grants_o,grants_unmasked_lo;

  bsg_priority_encode_one_hot_out_width_p128_lo_to_hi_p1
  enc
  (
    .i(reqs_i),
    .o(grants_unmasked_lo)
  );

  assign grants_o[127] = grants_unmasked_lo[127] & ready_i;
  assign grants_o[126] = grants_unmasked_lo[126] & ready_i;
  assign grants_o[125] = grants_unmasked_lo[125] & ready_i;
  assign grants_o[124] = grants_unmasked_lo[124] & ready_i;
  assign grants_o[123] = grants_unmasked_lo[123] & ready_i;
  assign grants_o[122] = grants_unmasked_lo[122] & ready_i;
  assign grants_o[121] = grants_unmasked_lo[121] & ready_i;
  assign grants_o[120] = grants_unmasked_lo[120] & ready_i;
  assign grants_o[119] = grants_unmasked_lo[119] & ready_i;
  assign grants_o[118] = grants_unmasked_lo[118] & ready_i;
  assign grants_o[117] = grants_unmasked_lo[117] & ready_i;
  assign grants_o[116] = grants_unmasked_lo[116] & ready_i;
  assign grants_o[115] = grants_unmasked_lo[115] & ready_i;
  assign grants_o[114] = grants_unmasked_lo[114] & ready_i;
  assign grants_o[113] = grants_unmasked_lo[113] & ready_i;
  assign grants_o[112] = grants_unmasked_lo[112] & ready_i;
  assign grants_o[111] = grants_unmasked_lo[111] & ready_i;
  assign grants_o[110] = grants_unmasked_lo[110] & ready_i;
  assign grants_o[109] = grants_unmasked_lo[109] & ready_i;
  assign grants_o[108] = grants_unmasked_lo[108] & ready_i;
  assign grants_o[107] = grants_unmasked_lo[107] & ready_i;
  assign grants_o[106] = grants_unmasked_lo[106] & ready_i;
  assign grants_o[105] = grants_unmasked_lo[105] & ready_i;
  assign grants_o[104] = grants_unmasked_lo[104] & ready_i;
  assign grants_o[103] = grants_unmasked_lo[103] & ready_i;
  assign grants_o[102] = grants_unmasked_lo[102] & ready_i;
  assign grants_o[101] = grants_unmasked_lo[101] & ready_i;
  assign grants_o[100] = grants_unmasked_lo[100] & ready_i;
  assign grants_o[99] = grants_unmasked_lo[99] & ready_i;
  assign grants_o[98] = grants_unmasked_lo[98] & ready_i;
  assign grants_o[97] = grants_unmasked_lo[97] & ready_i;
  assign grants_o[96] = grants_unmasked_lo[96] & ready_i;
  assign grants_o[95] = grants_unmasked_lo[95] & ready_i;
  assign grants_o[94] = grants_unmasked_lo[94] & ready_i;
  assign grants_o[93] = grants_unmasked_lo[93] & ready_i;
  assign grants_o[92] = grants_unmasked_lo[92] & ready_i;
  assign grants_o[91] = grants_unmasked_lo[91] & ready_i;
  assign grants_o[90] = grants_unmasked_lo[90] & ready_i;
  assign grants_o[89] = grants_unmasked_lo[89] & ready_i;
  assign grants_o[88] = grants_unmasked_lo[88] & ready_i;
  assign grants_o[87] = grants_unmasked_lo[87] & ready_i;
  assign grants_o[86] = grants_unmasked_lo[86] & ready_i;
  assign grants_o[85] = grants_unmasked_lo[85] & ready_i;
  assign grants_o[84] = grants_unmasked_lo[84] & ready_i;
  assign grants_o[83] = grants_unmasked_lo[83] & ready_i;
  assign grants_o[82] = grants_unmasked_lo[82] & ready_i;
  assign grants_o[81] = grants_unmasked_lo[81] & ready_i;
  assign grants_o[80] = grants_unmasked_lo[80] & ready_i;
  assign grants_o[79] = grants_unmasked_lo[79] & ready_i;
  assign grants_o[78] = grants_unmasked_lo[78] & ready_i;
  assign grants_o[77] = grants_unmasked_lo[77] & ready_i;
  assign grants_o[76] = grants_unmasked_lo[76] & ready_i;
  assign grants_o[75] = grants_unmasked_lo[75] & ready_i;
  assign grants_o[74] = grants_unmasked_lo[74] & ready_i;
  assign grants_o[73] = grants_unmasked_lo[73] & ready_i;
  assign grants_o[72] = grants_unmasked_lo[72] & ready_i;
  assign grants_o[71] = grants_unmasked_lo[71] & ready_i;
  assign grants_o[70] = grants_unmasked_lo[70] & ready_i;
  assign grants_o[69] = grants_unmasked_lo[69] & ready_i;
  assign grants_o[68] = grants_unmasked_lo[68] & ready_i;
  assign grants_o[67] = grants_unmasked_lo[67] & ready_i;
  assign grants_o[66] = grants_unmasked_lo[66] & ready_i;
  assign grants_o[65] = grants_unmasked_lo[65] & ready_i;
  assign grants_o[64] = grants_unmasked_lo[64] & ready_i;
  assign grants_o[63] = grants_unmasked_lo[63] & ready_i;
  assign grants_o[62] = grants_unmasked_lo[62] & ready_i;
  assign grants_o[61] = grants_unmasked_lo[61] & ready_i;
  assign grants_o[60] = grants_unmasked_lo[60] & ready_i;
  assign grants_o[59] = grants_unmasked_lo[59] & ready_i;
  assign grants_o[58] = grants_unmasked_lo[58] & ready_i;
  assign grants_o[57] = grants_unmasked_lo[57] & ready_i;
  assign grants_o[56] = grants_unmasked_lo[56] & ready_i;
  assign grants_o[55] = grants_unmasked_lo[55] & ready_i;
  assign grants_o[54] = grants_unmasked_lo[54] & ready_i;
  assign grants_o[53] = grants_unmasked_lo[53] & ready_i;
  assign grants_o[52] = grants_unmasked_lo[52] & ready_i;
  assign grants_o[51] = grants_unmasked_lo[51] & ready_i;
  assign grants_o[50] = grants_unmasked_lo[50] & ready_i;
  assign grants_o[49] = grants_unmasked_lo[49] & ready_i;
  assign grants_o[48] = grants_unmasked_lo[48] & ready_i;
  assign grants_o[47] = grants_unmasked_lo[47] & ready_i;
  assign grants_o[46] = grants_unmasked_lo[46] & ready_i;
  assign grants_o[45] = grants_unmasked_lo[45] & ready_i;
  assign grants_o[44] = grants_unmasked_lo[44] & ready_i;
  assign grants_o[43] = grants_unmasked_lo[43] & ready_i;
  assign grants_o[42] = grants_unmasked_lo[42] & ready_i;
  assign grants_o[41] = grants_unmasked_lo[41] & ready_i;
  assign grants_o[40] = grants_unmasked_lo[40] & ready_i;
  assign grants_o[39] = grants_unmasked_lo[39] & ready_i;
  assign grants_o[38] = grants_unmasked_lo[38] & ready_i;
  assign grants_o[37] = grants_unmasked_lo[37] & ready_i;
  assign grants_o[36] = grants_unmasked_lo[36] & ready_i;
  assign grants_o[35] = grants_unmasked_lo[35] & ready_i;
  assign grants_o[34] = grants_unmasked_lo[34] & ready_i;
  assign grants_o[33] = grants_unmasked_lo[33] & ready_i;
  assign grants_o[32] = grants_unmasked_lo[32] & ready_i;
  assign grants_o[31] = grants_unmasked_lo[31] & ready_i;
  assign grants_o[30] = grants_unmasked_lo[30] & ready_i;
  assign grants_o[29] = grants_unmasked_lo[29] & ready_i;
  assign grants_o[28] = grants_unmasked_lo[28] & ready_i;
  assign grants_o[27] = grants_unmasked_lo[27] & ready_i;
  assign grants_o[26] = grants_unmasked_lo[26] & ready_i;
  assign grants_o[25] = grants_unmasked_lo[25] & ready_i;
  assign grants_o[24] = grants_unmasked_lo[24] & ready_i;
  assign grants_o[23] = grants_unmasked_lo[23] & ready_i;
  assign grants_o[22] = grants_unmasked_lo[22] & ready_i;
  assign grants_o[21] = grants_unmasked_lo[21] & ready_i;
  assign grants_o[20] = grants_unmasked_lo[20] & ready_i;
  assign grants_o[19] = grants_unmasked_lo[19] & ready_i;
  assign grants_o[18] = grants_unmasked_lo[18] & ready_i;
  assign grants_o[17] = grants_unmasked_lo[17] & ready_i;
  assign grants_o[16] = grants_unmasked_lo[16] & ready_i;
  assign grants_o[15] = grants_unmasked_lo[15] & ready_i;
  assign grants_o[14] = grants_unmasked_lo[14] & ready_i;
  assign grants_o[13] = grants_unmasked_lo[13] & ready_i;
  assign grants_o[12] = grants_unmasked_lo[12] & ready_i;
  assign grants_o[11] = grants_unmasked_lo[11] & ready_i;
  assign grants_o[10] = grants_unmasked_lo[10] & ready_i;
  assign grants_o[9] = grants_unmasked_lo[9] & ready_i;
  assign grants_o[8] = grants_unmasked_lo[8] & ready_i;
  assign grants_o[7] = grants_unmasked_lo[7] & ready_i;
  assign grants_o[6] = grants_unmasked_lo[6] & ready_i;
  assign grants_o[5] = grants_unmasked_lo[5] & ready_i;
  assign grants_o[4] = grants_unmasked_lo[4] & ready_i;
  assign grants_o[3] = grants_unmasked_lo[3] & ready_i;
  assign grants_o[2] = grants_unmasked_lo[2] & ready_i;
  assign grants_o[1] = grants_unmasked_lo[1] & ready_i;
  assign grants_o[0] = grants_unmasked_lo[0] & ready_i;

endmodule

