

module top
(
  clk_i,
  reset_i,
  v_i,
  tag_i,
  data_i,
  yumi_o,
  v_o,
  yumi_i,
  data_o
);

  input [5:0] tag_i;
  input [7:0] data_i;
  output [63:0] v_o;
  input [63:0] yumi_i;
  output [511:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  output yumi_o;

  bsg_1_to_n_tagged_fifo
  wrapper
  (
    .tag_i(tag_i),
    .data_i(data_i),
    .v_o(v_o),
    .yumi_i(yumi_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_o(yumi_o)
  );


endmodule



module bsg_decode_num_out_p64
(
  i,
  o
);

  input [5:0] i;
  output [63:0] o;
  wire [63:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_decode_with_v_num_out_p64
(
  i,
  v_i,
  o
);

  input [5:0] i;
  output [63:0] o;
  input v_i;
  wire [63:0] o,lo;

  bsg_decode_num_out_p64
  bd
  (
    .i(i),
    .o(lo)
  );

  assign o[63] = v_i & lo[63];
  assign o[62] = v_i & lo[62];
  assign o[61] = v_i & lo[61];
  assign o[60] = v_i & lo[60];
  assign o[59] = v_i & lo[59];
  assign o[58] = v_i & lo[58];
  assign o[57] = v_i & lo[57];
  assign o[56] = v_i & lo[56];
  assign o[55] = v_i & lo[55];
  assign o[54] = v_i & lo[54];
  assign o[53] = v_i & lo[53];
  assign o[52] = v_i & lo[52];
  assign o[51] = v_i & lo[51];
  assign o[50] = v_i & lo[50];
  assign o[49] = v_i & lo[49];
  assign o[48] = v_i & lo[48];
  assign o[47] = v_i & lo[47];
  assign o[46] = v_i & lo[46];
  assign o[45] = v_i & lo[45];
  assign o[44] = v_i & lo[44];
  assign o[43] = v_i & lo[43];
  assign o[42] = v_i & lo[42];
  assign o[41] = v_i & lo[41];
  assign o[40] = v_i & lo[40];
  assign o[39] = v_i & lo[39];
  assign o[38] = v_i & lo[38];
  assign o[37] = v_i & lo[37];
  assign o[36] = v_i & lo[36];
  assign o[35] = v_i & lo[35];
  assign o[34] = v_i & lo[34];
  assign o[33] = v_i & lo[33];
  assign o[32] = v_i & lo[32];
  assign o[31] = v_i & lo[31];
  assign o[30] = v_i & lo[30];
  assign o[29] = v_i & lo[29];
  assign o[28] = v_i & lo[28];
  assign o[27] = v_i & lo[27];
  assign o[26] = v_i & lo[26];
  assign o[25] = v_i & lo[25];
  assign o[24] = v_i & lo[24];
  assign o[23] = v_i & lo[23];
  assign o[22] = v_i & lo[22];
  assign o[21] = v_i & lo[21];
  assign o[20] = v_i & lo[20];
  assign o[19] = v_i & lo[19];
  assign o[18] = v_i & lo[18];
  assign o[17] = v_i & lo[17];
  assign o[16] = v_i & lo[16];
  assign o[15] = v_i & lo[15];
  assign o[14] = v_i & lo[14];
  assign o[13] = v_i & lo[13];
  assign o[12] = v_i & lo[12];
  assign o[11] = v_i & lo[11];
  assign o[10] = v_i & lo[10];
  assign o[9] = v_i & lo[9];
  assign o[8] = v_i & lo[8];
  assign o[7] = v_i & lo[7];
  assign o[6] = v_i & lo[6];
  assign o[5] = v_i & lo[5];
  assign o[4] = v_i & lo[4];
  assign o[3] = v_i & lo[3];
  assign o[2] = v_i & lo[2];
  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bsg_1_to_n_tagged_num_out_p64
(
  clk_i,
  reset_i,
  v_i,
  tag_i,
  yumi_o,
  v_o,
  ready_i
);

  input [5:0] tag_i;
  output [63:0] v_o;
  input [63:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output yumi_o;
  wire [63:0] v_o;
  wire yumi_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130;

  bsg_decode_with_v_num_out_p64
  many_bdv
  (
    .i(tag_i),
    .v_i(v_i),
    .o(v_o)
  );

  assign N130 = (N66)? ready_i[0] : 
                (N68)? ready_i[1] : 
                (N70)? ready_i[2] : 
                (N72)? ready_i[3] : 
                (N74)? ready_i[4] : 
                (N76)? ready_i[5] : 
                (N78)? ready_i[6] : 
                (N80)? ready_i[7] : 
                (N82)? ready_i[8] : 
                (N84)? ready_i[9] : 
                (N86)? ready_i[10] : 
                (N88)? ready_i[11] : 
                (N90)? ready_i[12] : 
                (N92)? ready_i[13] : 
                (N94)? ready_i[14] : 
                (N96)? ready_i[15] : 
                (N98)? ready_i[16] : 
                (N100)? ready_i[17] : 
                (N102)? ready_i[18] : 
                (N104)? ready_i[19] : 
                (N106)? ready_i[20] : 
                (N108)? ready_i[21] : 
                (N110)? ready_i[22] : 
                (N112)? ready_i[23] : 
                (N114)? ready_i[24] : 
                (N116)? ready_i[25] : 
                (N118)? ready_i[26] : 
                (N120)? ready_i[27] : 
                (N122)? ready_i[28] : 
                (N124)? ready_i[29] : 
                (N126)? ready_i[30] : 
                (N128)? ready_i[31] : 
                (N67)? ready_i[32] : 
                (N69)? ready_i[33] : 
                (N71)? ready_i[34] : 
                (N73)? ready_i[35] : 
                (N75)? ready_i[36] : 
                (N77)? ready_i[37] : 
                (N79)? ready_i[38] : 
                (N81)? ready_i[39] : 
                (N83)? ready_i[40] : 
                (N85)? ready_i[41] : 
                (N87)? ready_i[42] : 
                (N89)? ready_i[43] : 
                (N91)? ready_i[44] : 
                (N93)? ready_i[45] : 
                (N95)? ready_i[46] : 
                (N97)? ready_i[47] : 
                (N99)? ready_i[48] : 
                (N101)? ready_i[49] : 
                (N103)? ready_i[50] : 
                (N105)? ready_i[51] : 
                (N107)? ready_i[52] : 
                (N109)? ready_i[53] : 
                (N111)? ready_i[54] : 
                (N113)? ready_i[55] : 
                (N115)? ready_i[56] : 
                (N117)? ready_i[57] : 
                (N119)? ready_i[58] : 
                (N121)? ready_i[59] : 
                (N123)? ready_i[60] : 
                (N125)? ready_i[61] : 
                (N127)? ready_i[62] : 
                (N129)? ready_i[63] : 1'b0;
  assign N0 = ~tag_i[0];
  assign N1 = ~tag_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & tag_i[1];
  assign N4 = tag_i[0] & N1;
  assign N5 = tag_i[0] & tag_i[1];
  assign N6 = ~tag_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & tag_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & tag_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & tag_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & tag_i[2];
  assign N15 = ~tag_i[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & tag_i[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & tag_i[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & tag_i[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & tag_i[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & tag_i[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & tag_i[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & tag_i[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & tag_i[3];
  assign N32 = ~tag_i[4];
  assign N33 = N16 & N32;
  assign N34 = N16 & tag_i[4];
  assign N35 = N18 & N32;
  assign N36 = N18 & tag_i[4];
  assign N37 = N20 & N32;
  assign N38 = N20 & tag_i[4];
  assign N39 = N22 & N32;
  assign N40 = N22 & tag_i[4];
  assign N41 = N24 & N32;
  assign N42 = N24 & tag_i[4];
  assign N43 = N26 & N32;
  assign N44 = N26 & tag_i[4];
  assign N45 = N28 & N32;
  assign N46 = N28 & tag_i[4];
  assign N47 = N30 & N32;
  assign N48 = N30 & tag_i[4];
  assign N49 = N17 & N32;
  assign N50 = N17 & tag_i[4];
  assign N51 = N19 & N32;
  assign N52 = N19 & tag_i[4];
  assign N53 = N21 & N32;
  assign N54 = N21 & tag_i[4];
  assign N55 = N23 & N32;
  assign N56 = N23 & tag_i[4];
  assign N57 = N25 & N32;
  assign N58 = N25 & tag_i[4];
  assign N59 = N27 & N32;
  assign N60 = N27 & tag_i[4];
  assign N61 = N29 & N32;
  assign N62 = N29 & tag_i[4];
  assign N63 = N31 & N32;
  assign N64 = N31 & tag_i[4];
  assign N65 = ~tag_i[5];
  assign N66 = N33 & N65;
  assign N67 = N33 & tag_i[5];
  assign N68 = N35 & N65;
  assign N69 = N35 & tag_i[5];
  assign N70 = N37 & N65;
  assign N71 = N37 & tag_i[5];
  assign N72 = N39 & N65;
  assign N73 = N39 & tag_i[5];
  assign N74 = N41 & N65;
  assign N75 = N41 & tag_i[5];
  assign N76 = N43 & N65;
  assign N77 = N43 & tag_i[5];
  assign N78 = N45 & N65;
  assign N79 = N45 & tag_i[5];
  assign N80 = N47 & N65;
  assign N81 = N47 & tag_i[5];
  assign N82 = N49 & N65;
  assign N83 = N49 & tag_i[5];
  assign N84 = N51 & N65;
  assign N85 = N51 & tag_i[5];
  assign N86 = N53 & N65;
  assign N87 = N53 & tag_i[5];
  assign N88 = N55 & N65;
  assign N89 = N55 & tag_i[5];
  assign N90 = N57 & N65;
  assign N91 = N57 & tag_i[5];
  assign N92 = N59 & N65;
  assign N93 = N59 & tag_i[5];
  assign N94 = N61 & N65;
  assign N95 = N61 & tag_i[5];
  assign N96 = N63 & N65;
  assign N97 = N63 & tag_i[5];
  assign N98 = N34 & N65;
  assign N99 = N34 & tag_i[5];
  assign N100 = N36 & N65;
  assign N101 = N36 & tag_i[5];
  assign N102 = N38 & N65;
  assign N103 = N38 & tag_i[5];
  assign N104 = N40 & N65;
  assign N105 = N40 & tag_i[5];
  assign N106 = N42 & N65;
  assign N107 = N42 & tag_i[5];
  assign N108 = N44 & N65;
  assign N109 = N44 & tag_i[5];
  assign N110 = N46 & N65;
  assign N111 = N46 & tag_i[5];
  assign N112 = N48 & N65;
  assign N113 = N48 & tag_i[5];
  assign N114 = N50 & N65;
  assign N115 = N50 & tag_i[5];
  assign N116 = N52 & N65;
  assign N117 = N52 & tag_i[5];
  assign N118 = N54 & N65;
  assign N119 = N54 & tag_i[5];
  assign N120 = N56 & N65;
  assign N121 = N56 & tag_i[5];
  assign N122 = N58 & N65;
  assign N123 = N58 & tag_i[5];
  assign N124 = N60 & N65;
  assign N125 = N60 & tag_i[5];
  assign N126 = N62 & N65;
  assign N127 = N62 & tag_i[5];
  assign N128 = N64 & N65;
  assign N129 = N64 & tag_i[5];
  assign yumi_o = N130 & v_i;

endmodule



module bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  ready_o,
  v_o,
  data_o,
  yumi_i
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [7:0] data_o,little_data,big_data_lo;
  wire ready_o,v_o,N0,N1,N2,N3,little_ready_lo,little_will_have_space,N4,N5,big_deq,N6,
  big_full_lo,big_empty_lo,N7,N8,little_valid,big_enq,N9,N10,N11,N12,N13,
  big_valid,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;
  reg big_deq_r;

  bsg_fifo_1rw_large
  big1p
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(big_valid),
    .enq_not_deq_i(big_enq),
    .full_o(big_full_lo),
    .empty_o(big_empty_lo),
    .data_o(big_data_lo)
  );


  bsg_two_fifo
  little2p
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(little_ready_lo),
    .data_i(little_data),
    .v_i(little_valid),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );

  assign N6 = (N0)? 1'b0 : 
              (N1)? big_deq : 1'b0;
  assign N0 = N5;
  assign N1 = N4;
  assign little_valid = (N2)? 1'b1 : 
                        (N15)? N10 : 
                        (N8)? 1'b0 : 1'b0;
  assign N2 = big_deq_r;
  assign big_enq = (N2)? v_i : 
                   (N15)? N11 : 
                   (N8)? N12 : 1'b0;
  assign big_deq = (N2)? N9 : 
                   (N15)? 1'b0 : 
                   (N8)? N13 : 1'b0;
  assign little_data = (N2)? big_data_lo : 
                       (N3)? data_i : 1'b0;
  assign N3 = N16;
  assign little_will_have_space = little_ready_lo | yumi_i;
  assign N4 = ~reset_i;
  assign N5 = reset_i;
  assign ready_o = ~big_full_lo;
  assign N7 = big_empty_lo | big_deq_r;
  assign N8 = ~N7;
  assign N9 = N19 & N20;
  assign N19 = N17 & N18;
  assign N17 = ~big_empty_lo;
  assign N18 = ~v_i;
  assign N20 = ~v_o;
  assign N10 = v_i & little_will_have_space;
  assign N11 = v_i & N21;
  assign N21 = ~little_will_have_space;
  assign N12 = v_i & N22;
  assign N22 = ~big_full_lo;
  assign N13 = N23 & little_will_have_space;
  assign N23 = ~N12;
  assign big_valid = big_enq | big_deq;
  assign N14 = ~big_deq_r;
  assign N15 = big_empty_lo & N14;
  assign N16 = ~big_deq_r;

  always @(posedge clk_i) begin
    if(1'b1) begin
      big_deq_r <= N6;
    end 
  end


endmodule



module bsg_1_to_n_tagged_fifo
(
  clk_i,
  reset_i,
  v_i,
  tag_i,
  data_i,
  yumi_o,
  v_o,
  yumi_i,
  data_o
);

  input [5:0] tag_i;
  input [7:0] data_i;
  output [63:0] v_o;
  input [63:0] yumi_i;
  output [511:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  output yumi_o;
  wire [63:0] v_o,valid_lo,ready_li;
  wire [511:0] data_o;
  wire yumi_o;

  bsg_1_to_n_tagged_num_out_p64
  u_1_to_n
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .tag_i(tag_i),
    .yumi_o(yumi_o),
    .v_o(valid_lo),
    .ready_i(ready_li)
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_0__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[0]),
    .ready_o(ready_li[0]),
    .v_o(v_o[0]),
    .data_o(data_o[7:0]),
    .yumi_i(yumi_i[0])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_1__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[1]),
    .ready_o(ready_li[1]),
    .v_o(v_o[1]),
    .data_o(data_o[15:8]),
    .yumi_i(yumi_i[1])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_2__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[2]),
    .ready_o(ready_li[2]),
    .v_o(v_o[2]),
    .data_o(data_o[23:16]),
    .yumi_i(yumi_i[2])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_3__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[3]),
    .ready_o(ready_li[3]),
    .v_o(v_o[3]),
    .data_o(data_o[31:24]),
    .yumi_i(yumi_i[3])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_4__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[4]),
    .ready_o(ready_li[4]),
    .v_o(v_o[4]),
    .data_o(data_o[39:32]),
    .yumi_i(yumi_i[4])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_5__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[5]),
    .ready_o(ready_li[5]),
    .v_o(v_o[5]),
    .data_o(data_o[47:40]),
    .yumi_i(yumi_i[5])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_6__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[6]),
    .ready_o(ready_li[6]),
    .v_o(v_o[6]),
    .data_o(data_o[55:48]),
    .yumi_i(yumi_i[6])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_7__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[7]),
    .ready_o(ready_li[7]),
    .v_o(v_o[7]),
    .data_o(data_o[63:56]),
    .yumi_i(yumi_i[7])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_8__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[8]),
    .ready_o(ready_li[8]),
    .v_o(v_o[8]),
    .data_o(data_o[71:64]),
    .yumi_i(yumi_i[8])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_9__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[9]),
    .ready_o(ready_li[9]),
    .v_o(v_o[9]),
    .data_o(data_o[79:72]),
    .yumi_i(yumi_i[9])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_10__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[10]),
    .ready_o(ready_li[10]),
    .v_o(v_o[10]),
    .data_o(data_o[87:80]),
    .yumi_i(yumi_i[10])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_11__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[11]),
    .ready_o(ready_li[11]),
    .v_o(v_o[11]),
    .data_o(data_o[95:88]),
    .yumi_i(yumi_i[11])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_12__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[12]),
    .ready_o(ready_li[12]),
    .v_o(v_o[12]),
    .data_o(data_o[103:96]),
    .yumi_i(yumi_i[12])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_13__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[13]),
    .ready_o(ready_li[13]),
    .v_o(v_o[13]),
    .data_o(data_o[111:104]),
    .yumi_i(yumi_i[13])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_14__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[14]),
    .ready_o(ready_li[14]),
    .v_o(v_o[14]),
    .data_o(data_o[119:112]),
    .yumi_i(yumi_i[14])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_15__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[15]),
    .ready_o(ready_li[15]),
    .v_o(v_o[15]),
    .data_o(data_o[127:120]),
    .yumi_i(yumi_i[15])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_16__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[16]),
    .ready_o(ready_li[16]),
    .v_o(v_o[16]),
    .data_o(data_o[135:128]),
    .yumi_i(yumi_i[16])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_17__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[17]),
    .ready_o(ready_li[17]),
    .v_o(v_o[17]),
    .data_o(data_o[143:136]),
    .yumi_i(yumi_i[17])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_18__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[18]),
    .ready_o(ready_li[18]),
    .v_o(v_o[18]),
    .data_o(data_o[151:144]),
    .yumi_i(yumi_i[18])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_19__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[19]),
    .ready_o(ready_li[19]),
    .v_o(v_o[19]),
    .data_o(data_o[159:152]),
    .yumi_i(yumi_i[19])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_20__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[20]),
    .ready_o(ready_li[20]),
    .v_o(v_o[20]),
    .data_o(data_o[167:160]),
    .yumi_i(yumi_i[20])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_21__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[21]),
    .ready_o(ready_li[21]),
    .v_o(v_o[21]),
    .data_o(data_o[175:168]),
    .yumi_i(yumi_i[21])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_22__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[22]),
    .ready_o(ready_li[22]),
    .v_o(v_o[22]),
    .data_o(data_o[183:176]),
    .yumi_i(yumi_i[22])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_23__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[23]),
    .ready_o(ready_li[23]),
    .v_o(v_o[23]),
    .data_o(data_o[191:184]),
    .yumi_i(yumi_i[23])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_24__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[24]),
    .ready_o(ready_li[24]),
    .v_o(v_o[24]),
    .data_o(data_o[199:192]),
    .yumi_i(yumi_i[24])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_25__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[25]),
    .ready_o(ready_li[25]),
    .v_o(v_o[25]),
    .data_o(data_o[207:200]),
    .yumi_i(yumi_i[25])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_26__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[26]),
    .ready_o(ready_li[26]),
    .v_o(v_o[26]),
    .data_o(data_o[215:208]),
    .yumi_i(yumi_i[26])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_27__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[27]),
    .ready_o(ready_li[27]),
    .v_o(v_o[27]),
    .data_o(data_o[223:216]),
    .yumi_i(yumi_i[27])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_28__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[28]),
    .ready_o(ready_li[28]),
    .v_o(v_o[28]),
    .data_o(data_o[231:224]),
    .yumi_i(yumi_i[28])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_29__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[29]),
    .ready_o(ready_li[29]),
    .v_o(v_o[29]),
    .data_o(data_o[239:232]),
    .yumi_i(yumi_i[29])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_30__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[30]),
    .ready_o(ready_li[30]),
    .v_o(v_o[30]),
    .data_o(data_o[247:240]),
    .yumi_i(yumi_i[30])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_31__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[31]),
    .ready_o(ready_li[31]),
    .v_o(v_o[31]),
    .data_o(data_o[255:248]),
    .yumi_i(yumi_i[31])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_32__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[32]),
    .ready_o(ready_li[32]),
    .v_o(v_o[32]),
    .data_o(data_o[263:256]),
    .yumi_i(yumi_i[32])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_33__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[33]),
    .ready_o(ready_li[33]),
    .v_o(v_o[33]),
    .data_o(data_o[271:264]),
    .yumi_i(yumi_i[33])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_34__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[34]),
    .ready_o(ready_li[34]),
    .v_o(v_o[34]),
    .data_o(data_o[279:272]),
    .yumi_i(yumi_i[34])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_35__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[35]),
    .ready_o(ready_li[35]),
    .v_o(v_o[35]),
    .data_o(data_o[287:280]),
    .yumi_i(yumi_i[35])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_36__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[36]),
    .ready_o(ready_li[36]),
    .v_o(v_o[36]),
    .data_o(data_o[295:288]),
    .yumi_i(yumi_i[36])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_37__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[37]),
    .ready_o(ready_li[37]),
    .v_o(v_o[37]),
    .data_o(data_o[303:296]),
    .yumi_i(yumi_i[37])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_38__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[38]),
    .ready_o(ready_li[38]),
    .v_o(v_o[38]),
    .data_o(data_o[311:304]),
    .yumi_i(yumi_i[38])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_39__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[39]),
    .ready_o(ready_li[39]),
    .v_o(v_o[39]),
    .data_o(data_o[319:312]),
    .yumi_i(yumi_i[39])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_40__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[40]),
    .ready_o(ready_li[40]),
    .v_o(v_o[40]),
    .data_o(data_o[327:320]),
    .yumi_i(yumi_i[40])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_41__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[41]),
    .ready_o(ready_li[41]),
    .v_o(v_o[41]),
    .data_o(data_o[335:328]),
    .yumi_i(yumi_i[41])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_42__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[42]),
    .ready_o(ready_li[42]),
    .v_o(v_o[42]),
    .data_o(data_o[343:336]),
    .yumi_i(yumi_i[42])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_43__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[43]),
    .ready_o(ready_li[43]),
    .v_o(v_o[43]),
    .data_o(data_o[351:344]),
    .yumi_i(yumi_i[43])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_44__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[44]),
    .ready_o(ready_li[44]),
    .v_o(v_o[44]),
    .data_o(data_o[359:352]),
    .yumi_i(yumi_i[44])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_45__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[45]),
    .ready_o(ready_li[45]),
    .v_o(v_o[45]),
    .data_o(data_o[367:360]),
    .yumi_i(yumi_i[45])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_46__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[46]),
    .ready_o(ready_li[46]),
    .v_o(v_o[46]),
    .data_o(data_o[375:368]),
    .yumi_i(yumi_i[46])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_47__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[47]),
    .ready_o(ready_li[47]),
    .v_o(v_o[47]),
    .data_o(data_o[383:376]),
    .yumi_i(yumi_i[47])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_48__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[48]),
    .ready_o(ready_li[48]),
    .v_o(v_o[48]),
    .data_o(data_o[391:384]),
    .yumi_i(yumi_i[48])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_49__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[49]),
    .ready_o(ready_li[49]),
    .v_o(v_o[49]),
    .data_o(data_o[399:392]),
    .yumi_i(yumi_i[49])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_50__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[50]),
    .ready_o(ready_li[50]),
    .v_o(v_o[50]),
    .data_o(data_o[407:400]),
    .yumi_i(yumi_i[50])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_51__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[51]),
    .ready_o(ready_li[51]),
    .v_o(v_o[51]),
    .data_o(data_o[415:408]),
    .yumi_i(yumi_i[51])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_52__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[52]),
    .ready_o(ready_li[52]),
    .v_o(v_o[52]),
    .data_o(data_o[423:416]),
    .yumi_i(yumi_i[52])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_53__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[53]),
    .ready_o(ready_li[53]),
    .v_o(v_o[53]),
    .data_o(data_o[431:424]),
    .yumi_i(yumi_i[53])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_54__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[54]),
    .ready_o(ready_li[54]),
    .v_o(v_o[54]),
    .data_o(data_o[439:432]),
    .yumi_i(yumi_i[54])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_55__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[55]),
    .ready_o(ready_li[55]),
    .v_o(v_o[55]),
    .data_o(data_o[447:440]),
    .yumi_i(yumi_i[55])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_56__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[56]),
    .ready_o(ready_li[56]),
    .v_o(v_o[56]),
    .data_o(data_o[455:448]),
    .yumi_i(yumi_i[56])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_57__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[57]),
    .ready_o(ready_li[57]),
    .v_o(v_o[57]),
    .data_o(data_o[463:456]),
    .yumi_i(yumi_i[57])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_58__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[58]),
    .ready_o(ready_li[58]),
    .v_o(v_o[58]),
    .data_o(data_o[471:464]),
    .yumi_i(yumi_i[58])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_59__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[59]),
    .ready_o(ready_li[59]),
    .v_o(v_o[59]),
    .data_o(data_o[479:472]),
    .yumi_i(yumi_i[59])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_60__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[60]),
    .ready_o(ready_li[60]),
    .v_o(v_o[60]),
    .data_o(data_o[487:480]),
    .yumi_i(yumi_i[60])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_61__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[61]),
    .ready_o(ready_li[61]),
    .v_o(v_o[61]),
    .data_o(data_o[495:488]),
    .yumi_i(yumi_i[61])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_62__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[62]),
    .ready_o(ready_li[62]),
    .v_o(v_o[62]),
    .data_o(data_o[503:496]),
    .yumi_i(yumi_i[62])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_63__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[63]),
    .ready_o(ready_li[63]),
    .v_o(v_o[63]),
    .data_o(data_o[511:504]),
    .yumi_i(yumi_i[63])
  );


endmodule

