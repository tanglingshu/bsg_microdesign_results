

module top
(
  o
);

  output [127:0] o;

  bsg_tielo
  wrapper
  (
    .o(o)
  );


endmodule



module bsg_tielo
(
  o
);

  output [127:0] o;
  wire [127:0] o;
  assign o[0] = 1'b0;
  assign o[1] = 1'b0;
  assign o[2] = 1'b0;
  assign o[3] = 1'b0;
  assign o[4] = 1'b0;
  assign o[5] = 1'b0;
  assign o[6] = 1'b0;
  assign o[7] = 1'b0;
  assign o[8] = 1'b0;
  assign o[9] = 1'b0;
  assign o[10] = 1'b0;
  assign o[11] = 1'b0;
  assign o[12] = 1'b0;
  assign o[13] = 1'b0;
  assign o[14] = 1'b0;
  assign o[15] = 1'b0;
  assign o[16] = 1'b0;
  assign o[17] = 1'b0;
  assign o[18] = 1'b0;
  assign o[19] = 1'b0;
  assign o[20] = 1'b0;
  assign o[21] = 1'b0;
  assign o[22] = 1'b0;
  assign o[23] = 1'b0;
  assign o[24] = 1'b0;
  assign o[25] = 1'b0;
  assign o[26] = 1'b0;
  assign o[27] = 1'b0;
  assign o[28] = 1'b0;
  assign o[29] = 1'b0;
  assign o[30] = 1'b0;
  assign o[31] = 1'b0;
  assign o[32] = 1'b0;
  assign o[33] = 1'b0;
  assign o[34] = 1'b0;
  assign o[35] = 1'b0;
  assign o[36] = 1'b0;
  assign o[37] = 1'b0;
  assign o[38] = 1'b0;
  assign o[39] = 1'b0;
  assign o[40] = 1'b0;
  assign o[41] = 1'b0;
  assign o[42] = 1'b0;
  assign o[43] = 1'b0;
  assign o[44] = 1'b0;
  assign o[45] = 1'b0;
  assign o[46] = 1'b0;
  assign o[47] = 1'b0;
  assign o[48] = 1'b0;
  assign o[49] = 1'b0;
  assign o[50] = 1'b0;
  assign o[51] = 1'b0;
  assign o[52] = 1'b0;
  assign o[53] = 1'b0;
  assign o[54] = 1'b0;
  assign o[55] = 1'b0;
  assign o[56] = 1'b0;
  assign o[57] = 1'b0;
  assign o[58] = 1'b0;
  assign o[59] = 1'b0;
  assign o[60] = 1'b0;
  assign o[61] = 1'b0;
  assign o[62] = 1'b0;
  assign o[63] = 1'b0;
  assign o[64] = 1'b0;
  assign o[65] = 1'b0;
  assign o[66] = 1'b0;
  assign o[67] = 1'b0;
  assign o[68] = 1'b0;
  assign o[69] = 1'b0;
  assign o[70] = 1'b0;
  assign o[71] = 1'b0;
  assign o[72] = 1'b0;
  assign o[73] = 1'b0;
  assign o[74] = 1'b0;
  assign o[75] = 1'b0;
  assign o[76] = 1'b0;
  assign o[77] = 1'b0;
  assign o[78] = 1'b0;
  assign o[79] = 1'b0;
  assign o[80] = 1'b0;
  assign o[81] = 1'b0;
  assign o[82] = 1'b0;
  assign o[83] = 1'b0;
  assign o[84] = 1'b0;
  assign o[85] = 1'b0;
  assign o[86] = 1'b0;
  assign o[87] = 1'b0;
  assign o[88] = 1'b0;
  assign o[89] = 1'b0;
  assign o[90] = 1'b0;
  assign o[91] = 1'b0;
  assign o[92] = 1'b0;
  assign o[93] = 1'b0;
  assign o[94] = 1'b0;
  assign o[95] = 1'b0;
  assign o[96] = 1'b0;
  assign o[97] = 1'b0;
  assign o[98] = 1'b0;
  assign o[99] = 1'b0;
  assign o[100] = 1'b0;
  assign o[101] = 1'b0;
  assign o[102] = 1'b0;
  assign o[103] = 1'b0;
  assign o[104] = 1'b0;
  assign o[105] = 1'b0;
  assign o[106] = 1'b0;
  assign o[107] = 1'b0;
  assign o[108] = 1'b0;
  assign o[109] = 1'b0;
  assign o[110] = 1'b0;
  assign o[111] = 1'b0;
  assign o[112] = 1'b0;
  assign o[113] = 1'b0;
  assign o[114] = 1'b0;
  assign o[115] = 1'b0;
  assign o[116] = 1'b0;
  assign o[117] = 1'b0;
  assign o[118] = 1'b0;
  assign o[119] = 1'b0;
  assign o[120] = 1'b0;
  assign o[121] = 1'b0;
  assign o[122] = 1'b0;
  assign o[123] = 1'b0;
  assign o[124] = 1'b0;
  assign o[125] = 1'b0;
  assign o[126] = 1'b0;
  assign o[127] = 1'b0;

endmodule

