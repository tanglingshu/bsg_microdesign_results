

module top
(
  clk_i,
  data_i,
  data_o
);

  input [127:0] data_i;
  output [127:0] data_o;
  input clk_i;

  bsg_dff_chain
  wrapper
  (
    .data_i(data_i),
    .data_o(data_o),
    .clk_i(clk_i)
  );


endmodule



module bsg_dff_width_p128
(
  clk_i,
  data_i,
  data_o
);

  input [127:0] data_i;
  output [127:0] data_o;
  input clk_i;
  reg [127:0] data_o;

  always @(posedge clk_i) begin
    if(1'b1) begin
      { data_o[127:0] } <= { data_i[127:0] };
    end 
  end


endmodule



module bsg_dff_chain
(
  clk_i,
  data_i,
  data_o
);

  input [127:0] data_i;
  output [127:0] data_o;
  input clk_i;
  wire [127:0] data_o;
  wire chained_data_delayed_127__127_,chained_data_delayed_127__126_,
  chained_data_delayed_127__125_,chained_data_delayed_127__124_,chained_data_delayed_127__123_,
  chained_data_delayed_127__122_,chained_data_delayed_127__121_,
  chained_data_delayed_127__120_,chained_data_delayed_127__119_,chained_data_delayed_127__118_,
  chained_data_delayed_127__117_,chained_data_delayed_127__116_,
  chained_data_delayed_127__115_,chained_data_delayed_127__114_,chained_data_delayed_127__113_,
  chained_data_delayed_127__112_,chained_data_delayed_127__111_,chained_data_delayed_127__110_,
  chained_data_delayed_127__109_,chained_data_delayed_127__108_,
  chained_data_delayed_127__107_,chained_data_delayed_127__106_,chained_data_delayed_127__105_,
  chained_data_delayed_127__104_,chained_data_delayed_127__103_,
  chained_data_delayed_127__102_,chained_data_delayed_127__101_,chained_data_delayed_127__100_,
  chained_data_delayed_127__99_,chained_data_delayed_127__98_,chained_data_delayed_127__97_,
  chained_data_delayed_127__96_,chained_data_delayed_127__95_,
  chained_data_delayed_127__94_,chained_data_delayed_127__93_,chained_data_delayed_127__92_,
  chained_data_delayed_127__91_,chained_data_delayed_127__90_,chained_data_delayed_127__89_,
  chained_data_delayed_127__88_,chained_data_delayed_127__87_,
  chained_data_delayed_127__86_,chained_data_delayed_127__85_,chained_data_delayed_127__84_,
  chained_data_delayed_127__83_,chained_data_delayed_127__82_,chained_data_delayed_127__81_,
  chained_data_delayed_127__80_,chained_data_delayed_127__79_,
  chained_data_delayed_127__78_,chained_data_delayed_127__77_,chained_data_delayed_127__76_,
  chained_data_delayed_127__75_,chained_data_delayed_127__74_,chained_data_delayed_127__73_,
  chained_data_delayed_127__72_,chained_data_delayed_127__71_,
  chained_data_delayed_127__70_,chained_data_delayed_127__69_,chained_data_delayed_127__68_,
  chained_data_delayed_127__67_,chained_data_delayed_127__66_,chained_data_delayed_127__65_,
  chained_data_delayed_127__64_,chained_data_delayed_127__63_,
  chained_data_delayed_127__62_,chained_data_delayed_127__61_,chained_data_delayed_127__60_,
  chained_data_delayed_127__59_,chained_data_delayed_127__58_,chained_data_delayed_127__57_,
  chained_data_delayed_127__56_,chained_data_delayed_127__55_,
  chained_data_delayed_127__54_,chained_data_delayed_127__53_,chained_data_delayed_127__52_,
  chained_data_delayed_127__51_,chained_data_delayed_127__50_,chained_data_delayed_127__49_,
  chained_data_delayed_127__48_,chained_data_delayed_127__47_,
  chained_data_delayed_127__46_,chained_data_delayed_127__45_,chained_data_delayed_127__44_,
  chained_data_delayed_127__43_,chained_data_delayed_127__42_,chained_data_delayed_127__41_,
  chained_data_delayed_127__40_,chained_data_delayed_127__39_,
  chained_data_delayed_127__38_,chained_data_delayed_127__37_,chained_data_delayed_127__36_,
  chained_data_delayed_127__35_,chained_data_delayed_127__34_,chained_data_delayed_127__33_,
  chained_data_delayed_127__32_,chained_data_delayed_127__31_,
  chained_data_delayed_127__30_,chained_data_delayed_127__29_,chained_data_delayed_127__28_,
  chained_data_delayed_127__27_,chained_data_delayed_127__26_,chained_data_delayed_127__25_,
  chained_data_delayed_127__24_,chained_data_delayed_127__23_,
  chained_data_delayed_127__22_,chained_data_delayed_127__21_,chained_data_delayed_127__20_,
  chained_data_delayed_127__19_,chained_data_delayed_127__18_,chained_data_delayed_127__17_,
  chained_data_delayed_127__16_,chained_data_delayed_127__15_,
  chained_data_delayed_127__14_,chained_data_delayed_127__13_,chained_data_delayed_127__12_,
  chained_data_delayed_127__11_,chained_data_delayed_127__10_,chained_data_delayed_127__9_,
  chained_data_delayed_127__8_,chained_data_delayed_127__7_,
  chained_data_delayed_127__6_,chained_data_delayed_127__5_,chained_data_delayed_127__4_,
  chained_data_delayed_127__3_,chained_data_delayed_127__2_,chained_data_delayed_127__1_,
  chained_data_delayed_127__0_,chained_data_delayed_126__127_,chained_data_delayed_126__126_,
  chained_data_delayed_126__125_,chained_data_delayed_126__124_,
  chained_data_delayed_126__123_,chained_data_delayed_126__122_,chained_data_delayed_126__121_,
  chained_data_delayed_126__120_,chained_data_delayed_126__119_,
  chained_data_delayed_126__118_,chained_data_delayed_126__117_,chained_data_delayed_126__116_,
  chained_data_delayed_126__115_,chained_data_delayed_126__114_,
  chained_data_delayed_126__113_,chained_data_delayed_126__112_,chained_data_delayed_126__111_,
  chained_data_delayed_126__110_,chained_data_delayed_126__109_,chained_data_delayed_126__108_,
  chained_data_delayed_126__107_,chained_data_delayed_126__106_,
  chained_data_delayed_126__105_,chained_data_delayed_126__104_,chained_data_delayed_126__103_,
  chained_data_delayed_126__102_,chained_data_delayed_126__101_,
  chained_data_delayed_126__100_,chained_data_delayed_126__99_,chained_data_delayed_126__98_,
  chained_data_delayed_126__97_,chained_data_delayed_126__96_,chained_data_delayed_126__95_,
  chained_data_delayed_126__94_,chained_data_delayed_126__93_,
  chained_data_delayed_126__92_,chained_data_delayed_126__91_,chained_data_delayed_126__90_,
  chained_data_delayed_126__89_,chained_data_delayed_126__88_,chained_data_delayed_126__87_,
  chained_data_delayed_126__86_,chained_data_delayed_126__85_,
  chained_data_delayed_126__84_,chained_data_delayed_126__83_,chained_data_delayed_126__82_,
  chained_data_delayed_126__81_,chained_data_delayed_126__80_,chained_data_delayed_126__79_,
  chained_data_delayed_126__78_,chained_data_delayed_126__77_,
  chained_data_delayed_126__76_,chained_data_delayed_126__75_,chained_data_delayed_126__74_,
  chained_data_delayed_126__73_,chained_data_delayed_126__72_,chained_data_delayed_126__71_,
  chained_data_delayed_126__70_,chained_data_delayed_126__69_,
  chained_data_delayed_126__68_,chained_data_delayed_126__67_,chained_data_delayed_126__66_,
  chained_data_delayed_126__65_,chained_data_delayed_126__64_,chained_data_delayed_126__63_,
  chained_data_delayed_126__62_,chained_data_delayed_126__61_,
  chained_data_delayed_126__60_,chained_data_delayed_126__59_,chained_data_delayed_126__58_,
  chained_data_delayed_126__57_,chained_data_delayed_126__56_,chained_data_delayed_126__55_,
  chained_data_delayed_126__54_,chained_data_delayed_126__53_,
  chained_data_delayed_126__52_,chained_data_delayed_126__51_,chained_data_delayed_126__50_,
  chained_data_delayed_126__49_,chained_data_delayed_126__48_,chained_data_delayed_126__47_,
  chained_data_delayed_126__46_,chained_data_delayed_126__45_,
  chained_data_delayed_126__44_,chained_data_delayed_126__43_,chained_data_delayed_126__42_,
  chained_data_delayed_126__41_,chained_data_delayed_126__40_,chained_data_delayed_126__39_,
  chained_data_delayed_126__38_,chained_data_delayed_126__37_,
  chained_data_delayed_126__36_,chained_data_delayed_126__35_,chained_data_delayed_126__34_,
  chained_data_delayed_126__33_,chained_data_delayed_126__32_,chained_data_delayed_126__31_,
  chained_data_delayed_126__30_,chained_data_delayed_126__29_,
  chained_data_delayed_126__28_,chained_data_delayed_126__27_,chained_data_delayed_126__26_,
  chained_data_delayed_126__25_,chained_data_delayed_126__24_,chained_data_delayed_126__23_,
  chained_data_delayed_126__22_,chained_data_delayed_126__21_,
  chained_data_delayed_126__20_,chained_data_delayed_126__19_,chained_data_delayed_126__18_,
  chained_data_delayed_126__17_,chained_data_delayed_126__16_,chained_data_delayed_126__15_,
  chained_data_delayed_126__14_,chained_data_delayed_126__13_,
  chained_data_delayed_126__12_,chained_data_delayed_126__11_,chained_data_delayed_126__10_,
  chained_data_delayed_126__9_,chained_data_delayed_126__8_,chained_data_delayed_126__7_,
  chained_data_delayed_126__6_,chained_data_delayed_126__5_,chained_data_delayed_126__4_,
  chained_data_delayed_126__3_,chained_data_delayed_126__2_,
  chained_data_delayed_126__1_,chained_data_delayed_126__0_,chained_data_delayed_125__127_,
  chained_data_delayed_125__126_,chained_data_delayed_125__125_,chained_data_delayed_125__124_,
  chained_data_delayed_125__123_,chained_data_delayed_125__122_,
  chained_data_delayed_125__121_,chained_data_delayed_125__120_,chained_data_delayed_125__119_,
  chained_data_delayed_125__118_,chained_data_delayed_125__117_,
  chained_data_delayed_125__116_,chained_data_delayed_125__115_,chained_data_delayed_125__114_,
  chained_data_delayed_125__113_,chained_data_delayed_125__112_,
  chained_data_delayed_125__111_,chained_data_delayed_125__110_,chained_data_delayed_125__109_,
  chained_data_delayed_125__108_,chained_data_delayed_125__107_,chained_data_delayed_125__106_,
  chained_data_delayed_125__105_,chained_data_delayed_125__104_,
  chained_data_delayed_125__103_,chained_data_delayed_125__102_,chained_data_delayed_125__101_,
  chained_data_delayed_125__100_,chained_data_delayed_125__99_,
  chained_data_delayed_125__98_,chained_data_delayed_125__97_,chained_data_delayed_125__96_,
  chained_data_delayed_125__95_,chained_data_delayed_125__94_,chained_data_delayed_125__93_,
  chained_data_delayed_125__92_,chained_data_delayed_125__91_,
  chained_data_delayed_125__90_,chained_data_delayed_125__89_,chained_data_delayed_125__88_,
  chained_data_delayed_125__87_,chained_data_delayed_125__86_,chained_data_delayed_125__85_,
  chained_data_delayed_125__84_,chained_data_delayed_125__83_,
  chained_data_delayed_125__82_,chained_data_delayed_125__81_,chained_data_delayed_125__80_,
  chained_data_delayed_125__79_,chained_data_delayed_125__78_,chained_data_delayed_125__77_,
  chained_data_delayed_125__76_,chained_data_delayed_125__75_,
  chained_data_delayed_125__74_,chained_data_delayed_125__73_,chained_data_delayed_125__72_,
  chained_data_delayed_125__71_,chained_data_delayed_125__70_,chained_data_delayed_125__69_,
  chained_data_delayed_125__68_,chained_data_delayed_125__67_,
  chained_data_delayed_125__66_,chained_data_delayed_125__65_,chained_data_delayed_125__64_,
  chained_data_delayed_125__63_,chained_data_delayed_125__62_,chained_data_delayed_125__61_,
  chained_data_delayed_125__60_,chained_data_delayed_125__59_,
  chained_data_delayed_125__58_,chained_data_delayed_125__57_,chained_data_delayed_125__56_,
  chained_data_delayed_125__55_,chained_data_delayed_125__54_,chained_data_delayed_125__53_,
  chained_data_delayed_125__52_,chained_data_delayed_125__51_,
  chained_data_delayed_125__50_,chained_data_delayed_125__49_,chained_data_delayed_125__48_,
  chained_data_delayed_125__47_,chained_data_delayed_125__46_,chained_data_delayed_125__45_,
  chained_data_delayed_125__44_,chained_data_delayed_125__43_,
  chained_data_delayed_125__42_,chained_data_delayed_125__41_,chained_data_delayed_125__40_,
  chained_data_delayed_125__39_,chained_data_delayed_125__38_,chained_data_delayed_125__37_,
  chained_data_delayed_125__36_,chained_data_delayed_125__35_,
  chained_data_delayed_125__34_,chained_data_delayed_125__33_,chained_data_delayed_125__32_,
  chained_data_delayed_125__31_,chained_data_delayed_125__30_,chained_data_delayed_125__29_,
  chained_data_delayed_125__28_,chained_data_delayed_125__27_,
  chained_data_delayed_125__26_,chained_data_delayed_125__25_,chained_data_delayed_125__24_,
  chained_data_delayed_125__23_,chained_data_delayed_125__22_,chained_data_delayed_125__21_,
  chained_data_delayed_125__20_,chained_data_delayed_125__19_,
  chained_data_delayed_125__18_,chained_data_delayed_125__17_,chained_data_delayed_125__16_,
  chained_data_delayed_125__15_,chained_data_delayed_125__14_,chained_data_delayed_125__13_,
  chained_data_delayed_125__12_,chained_data_delayed_125__11_,
  chained_data_delayed_125__10_,chained_data_delayed_125__9_,chained_data_delayed_125__8_,
  chained_data_delayed_125__7_,chained_data_delayed_125__6_,chained_data_delayed_125__5_,
  chained_data_delayed_125__4_,chained_data_delayed_125__3_,chained_data_delayed_125__2_,
  chained_data_delayed_125__1_,chained_data_delayed_125__0_,
  chained_data_delayed_4__127_,chained_data_delayed_4__126_,chained_data_delayed_4__125_,
  chained_data_delayed_4__124_,chained_data_delayed_4__123_,chained_data_delayed_4__122_,
  chained_data_delayed_4__121_,chained_data_delayed_4__120_,chained_data_delayed_4__119_,
  chained_data_delayed_4__118_,chained_data_delayed_4__117_,
  chained_data_delayed_4__116_,chained_data_delayed_4__115_,chained_data_delayed_4__114_,
  chained_data_delayed_4__113_,chained_data_delayed_4__112_,chained_data_delayed_4__111_,
  chained_data_delayed_4__110_,chained_data_delayed_4__109_,chained_data_delayed_4__108_,
  chained_data_delayed_4__107_,chained_data_delayed_4__106_,
  chained_data_delayed_4__105_,chained_data_delayed_4__104_,chained_data_delayed_4__103_,
  chained_data_delayed_4__102_,chained_data_delayed_4__101_,chained_data_delayed_4__100_,
  chained_data_delayed_4__99_,chained_data_delayed_4__98_,chained_data_delayed_4__97_,
  chained_data_delayed_4__96_,chained_data_delayed_4__95_,chained_data_delayed_4__94_,
  chained_data_delayed_4__93_,chained_data_delayed_4__92_,chained_data_delayed_4__91_,
  chained_data_delayed_4__90_,chained_data_delayed_4__89_,
  chained_data_delayed_4__88_,chained_data_delayed_4__87_,chained_data_delayed_4__86_,
  chained_data_delayed_4__85_,chained_data_delayed_4__84_,chained_data_delayed_4__83_,
  chained_data_delayed_4__82_,chained_data_delayed_4__81_,chained_data_delayed_4__80_,
  chained_data_delayed_4__79_,chained_data_delayed_4__78_,chained_data_delayed_4__77_,
  chained_data_delayed_4__76_,chained_data_delayed_4__75_,chained_data_delayed_4__74_,
  chained_data_delayed_4__73_,chained_data_delayed_4__72_,chained_data_delayed_4__71_,
  chained_data_delayed_4__70_,chained_data_delayed_4__69_,
  chained_data_delayed_4__68_,chained_data_delayed_4__67_,chained_data_delayed_4__66_,
  chained_data_delayed_4__65_,chained_data_delayed_4__64_,chained_data_delayed_4__63_,
  chained_data_delayed_4__62_,chained_data_delayed_4__61_,chained_data_delayed_4__60_,
  chained_data_delayed_4__59_,chained_data_delayed_4__58_,chained_data_delayed_4__57_,
  chained_data_delayed_4__56_,chained_data_delayed_4__55_,chained_data_delayed_4__54_,
  chained_data_delayed_4__53_,chained_data_delayed_4__52_,chained_data_delayed_4__51_,
  chained_data_delayed_4__50_,chained_data_delayed_4__49_,
  chained_data_delayed_4__48_,chained_data_delayed_4__47_,chained_data_delayed_4__46_,
  chained_data_delayed_4__45_,chained_data_delayed_4__44_,chained_data_delayed_4__43_,
  chained_data_delayed_4__42_,chained_data_delayed_4__41_,chained_data_delayed_4__40_,
  chained_data_delayed_4__39_,chained_data_delayed_4__38_,chained_data_delayed_4__37_,
  chained_data_delayed_4__36_,chained_data_delayed_4__35_,chained_data_delayed_4__34_,
  chained_data_delayed_4__33_,chained_data_delayed_4__32_,chained_data_delayed_4__31_,
  chained_data_delayed_4__30_,chained_data_delayed_4__29_,
  chained_data_delayed_4__28_,chained_data_delayed_4__27_,chained_data_delayed_4__26_,
  chained_data_delayed_4__25_,chained_data_delayed_4__24_,chained_data_delayed_4__23_,
  chained_data_delayed_4__22_,chained_data_delayed_4__21_,chained_data_delayed_4__20_,
  chained_data_delayed_4__19_,chained_data_delayed_4__18_,chained_data_delayed_4__17_,
  chained_data_delayed_4__16_,chained_data_delayed_4__15_,chained_data_delayed_4__14_,
  chained_data_delayed_4__13_,chained_data_delayed_4__12_,chained_data_delayed_4__11_,
  chained_data_delayed_4__10_,chained_data_delayed_4__9_,chained_data_delayed_4__8_,
  chained_data_delayed_4__7_,chained_data_delayed_4__6_,
  chained_data_delayed_4__5_,chained_data_delayed_4__4_,chained_data_delayed_4__3_,
  chained_data_delayed_4__2_,chained_data_delayed_4__1_,chained_data_delayed_4__0_,
  chained_data_delayed_3__127_,chained_data_delayed_3__126_,chained_data_delayed_3__125_,
  chained_data_delayed_3__124_,chained_data_delayed_3__123_,chained_data_delayed_3__122_,
  chained_data_delayed_3__121_,chained_data_delayed_3__120_,chained_data_delayed_3__119_,
  chained_data_delayed_3__118_,chained_data_delayed_3__117_,
  chained_data_delayed_3__116_,chained_data_delayed_3__115_,chained_data_delayed_3__114_,
  chained_data_delayed_3__113_,chained_data_delayed_3__112_,chained_data_delayed_3__111_,
  chained_data_delayed_3__110_,chained_data_delayed_3__109_,chained_data_delayed_3__108_,
  chained_data_delayed_3__107_,chained_data_delayed_3__106_,
  chained_data_delayed_3__105_,chained_data_delayed_3__104_,chained_data_delayed_3__103_,
  chained_data_delayed_3__102_,chained_data_delayed_3__101_,chained_data_delayed_3__100_,
  chained_data_delayed_3__99_,chained_data_delayed_3__98_,chained_data_delayed_3__97_,
  chained_data_delayed_3__96_,chained_data_delayed_3__95_,chained_data_delayed_3__94_,
  chained_data_delayed_3__93_,chained_data_delayed_3__92_,chained_data_delayed_3__91_,
  chained_data_delayed_3__90_,chained_data_delayed_3__89_,
  chained_data_delayed_3__88_,chained_data_delayed_3__87_,chained_data_delayed_3__86_,
  chained_data_delayed_3__85_,chained_data_delayed_3__84_,chained_data_delayed_3__83_,
  chained_data_delayed_3__82_,chained_data_delayed_3__81_,chained_data_delayed_3__80_,
  chained_data_delayed_3__79_,chained_data_delayed_3__78_,chained_data_delayed_3__77_,
  chained_data_delayed_3__76_,chained_data_delayed_3__75_,chained_data_delayed_3__74_,
  chained_data_delayed_3__73_,chained_data_delayed_3__72_,chained_data_delayed_3__71_,
  chained_data_delayed_3__70_,chained_data_delayed_3__69_,
  chained_data_delayed_3__68_,chained_data_delayed_3__67_,chained_data_delayed_3__66_,
  chained_data_delayed_3__65_,chained_data_delayed_3__64_,chained_data_delayed_3__63_,
  chained_data_delayed_3__62_,chained_data_delayed_3__61_,chained_data_delayed_3__60_,
  chained_data_delayed_3__59_,chained_data_delayed_3__58_,chained_data_delayed_3__57_,
  chained_data_delayed_3__56_,chained_data_delayed_3__55_,chained_data_delayed_3__54_,
  chained_data_delayed_3__53_,chained_data_delayed_3__52_,chained_data_delayed_3__51_,
  chained_data_delayed_3__50_,chained_data_delayed_3__49_,
  chained_data_delayed_3__48_,chained_data_delayed_3__47_,chained_data_delayed_3__46_,
  chained_data_delayed_3__45_,chained_data_delayed_3__44_,chained_data_delayed_3__43_,
  chained_data_delayed_3__42_,chained_data_delayed_3__41_,chained_data_delayed_3__40_,
  chained_data_delayed_3__39_,chained_data_delayed_3__38_,chained_data_delayed_3__37_,
  chained_data_delayed_3__36_,chained_data_delayed_3__35_,chained_data_delayed_3__34_,
  chained_data_delayed_3__33_,chained_data_delayed_3__32_,chained_data_delayed_3__31_,
  chained_data_delayed_3__30_,chained_data_delayed_3__29_,
  chained_data_delayed_3__28_,chained_data_delayed_3__27_,chained_data_delayed_3__26_,
  chained_data_delayed_3__25_,chained_data_delayed_3__24_,chained_data_delayed_3__23_,
  chained_data_delayed_3__22_,chained_data_delayed_3__21_,chained_data_delayed_3__20_,
  chained_data_delayed_3__19_,chained_data_delayed_3__18_,chained_data_delayed_3__17_,
  chained_data_delayed_3__16_,chained_data_delayed_3__15_,chained_data_delayed_3__14_,
  chained_data_delayed_3__13_,chained_data_delayed_3__12_,chained_data_delayed_3__11_,
  chained_data_delayed_3__10_,chained_data_delayed_3__9_,
  chained_data_delayed_3__8_,chained_data_delayed_3__7_,chained_data_delayed_3__6_,
  chained_data_delayed_3__5_,chained_data_delayed_3__4_,chained_data_delayed_3__3_,
  chained_data_delayed_3__2_,chained_data_delayed_3__1_,chained_data_delayed_3__0_,
  chained_data_delayed_2__127_,chained_data_delayed_2__126_,chained_data_delayed_2__125_,
  chained_data_delayed_2__124_,chained_data_delayed_2__123_,chained_data_delayed_2__122_,
  chained_data_delayed_2__121_,chained_data_delayed_2__120_,chained_data_delayed_2__119_,
  chained_data_delayed_2__118_,chained_data_delayed_2__117_,
  chained_data_delayed_2__116_,chained_data_delayed_2__115_,chained_data_delayed_2__114_,
  chained_data_delayed_2__113_,chained_data_delayed_2__112_,chained_data_delayed_2__111_,
  chained_data_delayed_2__110_,chained_data_delayed_2__109_,chained_data_delayed_2__108_,
  chained_data_delayed_2__107_,chained_data_delayed_2__106_,
  chained_data_delayed_2__105_,chained_data_delayed_2__104_,chained_data_delayed_2__103_,
  chained_data_delayed_2__102_,chained_data_delayed_2__101_,chained_data_delayed_2__100_,
  chained_data_delayed_2__99_,chained_data_delayed_2__98_,chained_data_delayed_2__97_,
  chained_data_delayed_2__96_,chained_data_delayed_2__95_,chained_data_delayed_2__94_,
  chained_data_delayed_2__93_,chained_data_delayed_2__92_,
  chained_data_delayed_2__91_,chained_data_delayed_2__90_,chained_data_delayed_2__89_,
  chained_data_delayed_2__88_,chained_data_delayed_2__87_,chained_data_delayed_2__86_,
  chained_data_delayed_2__85_,chained_data_delayed_2__84_,chained_data_delayed_2__83_,
  chained_data_delayed_2__82_,chained_data_delayed_2__81_,chained_data_delayed_2__80_,
  chained_data_delayed_2__79_,chained_data_delayed_2__78_,chained_data_delayed_2__77_,
  chained_data_delayed_2__76_,chained_data_delayed_2__75_,chained_data_delayed_2__74_,
  chained_data_delayed_2__73_,chained_data_delayed_2__72_,
  chained_data_delayed_2__71_,chained_data_delayed_2__70_,chained_data_delayed_2__69_,
  chained_data_delayed_2__68_,chained_data_delayed_2__67_,chained_data_delayed_2__66_,
  chained_data_delayed_2__65_,chained_data_delayed_2__64_,chained_data_delayed_2__63_,
  chained_data_delayed_2__62_,chained_data_delayed_2__61_,chained_data_delayed_2__60_,
  chained_data_delayed_2__59_,chained_data_delayed_2__58_,chained_data_delayed_2__57_,
  chained_data_delayed_2__56_,chained_data_delayed_2__55_,chained_data_delayed_2__54_,
  chained_data_delayed_2__53_,chained_data_delayed_2__52_,
  chained_data_delayed_2__51_,chained_data_delayed_2__50_,chained_data_delayed_2__49_,
  chained_data_delayed_2__48_,chained_data_delayed_2__47_,chained_data_delayed_2__46_,
  chained_data_delayed_2__45_,chained_data_delayed_2__44_,chained_data_delayed_2__43_,
  chained_data_delayed_2__42_,chained_data_delayed_2__41_,chained_data_delayed_2__40_,
  chained_data_delayed_2__39_,chained_data_delayed_2__38_,chained_data_delayed_2__37_,
  chained_data_delayed_2__36_,chained_data_delayed_2__35_,chained_data_delayed_2__34_,
  chained_data_delayed_2__33_,chained_data_delayed_2__32_,
  chained_data_delayed_2__31_,chained_data_delayed_2__30_,chained_data_delayed_2__29_,
  chained_data_delayed_2__28_,chained_data_delayed_2__27_,chained_data_delayed_2__26_,
  chained_data_delayed_2__25_,chained_data_delayed_2__24_,chained_data_delayed_2__23_,
  chained_data_delayed_2__22_,chained_data_delayed_2__21_,chained_data_delayed_2__20_,
  chained_data_delayed_2__19_,chained_data_delayed_2__18_,chained_data_delayed_2__17_,
  chained_data_delayed_2__16_,chained_data_delayed_2__15_,chained_data_delayed_2__14_,
  chained_data_delayed_2__13_,chained_data_delayed_2__12_,
  chained_data_delayed_2__11_,chained_data_delayed_2__10_,chained_data_delayed_2__9_,
  chained_data_delayed_2__8_,chained_data_delayed_2__7_,chained_data_delayed_2__6_,
  chained_data_delayed_2__5_,chained_data_delayed_2__4_,chained_data_delayed_2__3_,
  chained_data_delayed_2__2_,chained_data_delayed_2__1_,chained_data_delayed_2__0_,
  chained_data_delayed_1__127_,chained_data_delayed_1__126_,chained_data_delayed_1__125_,
  chained_data_delayed_1__124_,chained_data_delayed_1__123_,chained_data_delayed_1__122_,
  chained_data_delayed_1__121_,chained_data_delayed_1__120_,
  chained_data_delayed_1__119_,chained_data_delayed_1__118_,chained_data_delayed_1__117_,
  chained_data_delayed_1__116_,chained_data_delayed_1__115_,chained_data_delayed_1__114_,
  chained_data_delayed_1__113_,chained_data_delayed_1__112_,chained_data_delayed_1__111_,
  chained_data_delayed_1__110_,chained_data_delayed_1__109_,chained_data_delayed_1__108_,
  chained_data_delayed_1__107_,chained_data_delayed_1__106_,
  chained_data_delayed_1__105_,chained_data_delayed_1__104_,chained_data_delayed_1__103_,
  chained_data_delayed_1__102_,chained_data_delayed_1__101_,chained_data_delayed_1__100_,
  chained_data_delayed_1__99_,chained_data_delayed_1__98_,chained_data_delayed_1__97_,
  chained_data_delayed_1__96_,chained_data_delayed_1__95_,chained_data_delayed_1__94_,
  chained_data_delayed_1__93_,chained_data_delayed_1__92_,
  chained_data_delayed_1__91_,chained_data_delayed_1__90_,chained_data_delayed_1__89_,
  chained_data_delayed_1__88_,chained_data_delayed_1__87_,chained_data_delayed_1__86_,
  chained_data_delayed_1__85_,chained_data_delayed_1__84_,chained_data_delayed_1__83_,
  chained_data_delayed_1__82_,chained_data_delayed_1__81_,chained_data_delayed_1__80_,
  chained_data_delayed_1__79_,chained_data_delayed_1__78_,chained_data_delayed_1__77_,
  chained_data_delayed_1__76_,chained_data_delayed_1__75_,chained_data_delayed_1__74_,
  chained_data_delayed_1__73_,chained_data_delayed_1__72_,
  chained_data_delayed_1__71_,chained_data_delayed_1__70_,chained_data_delayed_1__69_,
  chained_data_delayed_1__68_,chained_data_delayed_1__67_,chained_data_delayed_1__66_,
  chained_data_delayed_1__65_,chained_data_delayed_1__64_,chained_data_delayed_1__63_,
  chained_data_delayed_1__62_,chained_data_delayed_1__61_,chained_data_delayed_1__60_,
  chained_data_delayed_1__59_,chained_data_delayed_1__58_,chained_data_delayed_1__57_,
  chained_data_delayed_1__56_,chained_data_delayed_1__55_,chained_data_delayed_1__54_,
  chained_data_delayed_1__53_,chained_data_delayed_1__52_,
  chained_data_delayed_1__51_,chained_data_delayed_1__50_,chained_data_delayed_1__49_,
  chained_data_delayed_1__48_,chained_data_delayed_1__47_,chained_data_delayed_1__46_,
  chained_data_delayed_1__45_,chained_data_delayed_1__44_,chained_data_delayed_1__43_,
  chained_data_delayed_1__42_,chained_data_delayed_1__41_,chained_data_delayed_1__40_,
  chained_data_delayed_1__39_,chained_data_delayed_1__38_,chained_data_delayed_1__37_,
  chained_data_delayed_1__36_,chained_data_delayed_1__35_,chained_data_delayed_1__34_,
  chained_data_delayed_1__33_,chained_data_delayed_1__32_,
  chained_data_delayed_1__31_,chained_data_delayed_1__30_,chained_data_delayed_1__29_,
  chained_data_delayed_1__28_,chained_data_delayed_1__27_,chained_data_delayed_1__26_,
  chained_data_delayed_1__25_,chained_data_delayed_1__24_,chained_data_delayed_1__23_,
  chained_data_delayed_1__22_,chained_data_delayed_1__21_,chained_data_delayed_1__20_,
  chained_data_delayed_1__19_,chained_data_delayed_1__18_,chained_data_delayed_1__17_,
  chained_data_delayed_1__16_,chained_data_delayed_1__15_,chained_data_delayed_1__14_,
  chained_data_delayed_1__13_,chained_data_delayed_1__12_,
  chained_data_delayed_1__11_,chained_data_delayed_1__10_,chained_data_delayed_1__9_,
  chained_data_delayed_1__8_,chained_data_delayed_1__7_,chained_data_delayed_1__6_,
  chained_data_delayed_1__5_,chained_data_delayed_1__4_,chained_data_delayed_1__3_,
  chained_data_delayed_1__2_,chained_data_delayed_1__1_,chained_data_delayed_1__0_,
  chained_data_delayed_8__127_,chained_data_delayed_8__126_,chained_data_delayed_8__125_,
  chained_data_delayed_8__124_,chained_data_delayed_8__123_,chained_data_delayed_8__122_,
  chained_data_delayed_8__121_,chained_data_delayed_8__120_,
  chained_data_delayed_8__119_,chained_data_delayed_8__118_,chained_data_delayed_8__117_,
  chained_data_delayed_8__116_,chained_data_delayed_8__115_,chained_data_delayed_8__114_,
  chained_data_delayed_8__113_,chained_data_delayed_8__112_,chained_data_delayed_8__111_,
  chained_data_delayed_8__110_,chained_data_delayed_8__109_,
  chained_data_delayed_8__108_,chained_data_delayed_8__107_,chained_data_delayed_8__106_,
  chained_data_delayed_8__105_,chained_data_delayed_8__104_,chained_data_delayed_8__103_,
  chained_data_delayed_8__102_,chained_data_delayed_8__101_,chained_data_delayed_8__100_,
  chained_data_delayed_8__99_,chained_data_delayed_8__98_,chained_data_delayed_8__97_,
  chained_data_delayed_8__96_,chained_data_delayed_8__95_,
  chained_data_delayed_8__94_,chained_data_delayed_8__93_,chained_data_delayed_8__92_,
  chained_data_delayed_8__91_,chained_data_delayed_8__90_,chained_data_delayed_8__89_,
  chained_data_delayed_8__88_,chained_data_delayed_8__87_,chained_data_delayed_8__86_,
  chained_data_delayed_8__85_,chained_data_delayed_8__84_,chained_data_delayed_8__83_,
  chained_data_delayed_8__82_,chained_data_delayed_8__81_,chained_data_delayed_8__80_,
  chained_data_delayed_8__79_,chained_data_delayed_8__78_,chained_data_delayed_8__77_,
  chained_data_delayed_8__76_,chained_data_delayed_8__75_,
  chained_data_delayed_8__74_,chained_data_delayed_8__73_,chained_data_delayed_8__72_,
  chained_data_delayed_8__71_,chained_data_delayed_8__70_,chained_data_delayed_8__69_,
  chained_data_delayed_8__68_,chained_data_delayed_8__67_,chained_data_delayed_8__66_,
  chained_data_delayed_8__65_,chained_data_delayed_8__64_,chained_data_delayed_8__63_,
  chained_data_delayed_8__62_,chained_data_delayed_8__61_,chained_data_delayed_8__60_,
  chained_data_delayed_8__59_,chained_data_delayed_8__58_,chained_data_delayed_8__57_,
  chained_data_delayed_8__56_,chained_data_delayed_8__55_,
  chained_data_delayed_8__54_,chained_data_delayed_8__53_,chained_data_delayed_8__52_,
  chained_data_delayed_8__51_,chained_data_delayed_8__50_,chained_data_delayed_8__49_,
  chained_data_delayed_8__48_,chained_data_delayed_8__47_,chained_data_delayed_8__46_,
  chained_data_delayed_8__45_,chained_data_delayed_8__44_,chained_data_delayed_8__43_,
  chained_data_delayed_8__42_,chained_data_delayed_8__41_,chained_data_delayed_8__40_,
  chained_data_delayed_8__39_,chained_data_delayed_8__38_,chained_data_delayed_8__37_,
  chained_data_delayed_8__36_,chained_data_delayed_8__35_,
  chained_data_delayed_8__34_,chained_data_delayed_8__33_,chained_data_delayed_8__32_,
  chained_data_delayed_8__31_,chained_data_delayed_8__30_,chained_data_delayed_8__29_,
  chained_data_delayed_8__28_,chained_data_delayed_8__27_,chained_data_delayed_8__26_,
  chained_data_delayed_8__25_,chained_data_delayed_8__24_,chained_data_delayed_8__23_,
  chained_data_delayed_8__22_,chained_data_delayed_8__21_,chained_data_delayed_8__20_,
  chained_data_delayed_8__19_,chained_data_delayed_8__18_,chained_data_delayed_8__17_,
  chained_data_delayed_8__16_,chained_data_delayed_8__15_,
  chained_data_delayed_8__14_,chained_data_delayed_8__13_,chained_data_delayed_8__12_,
  chained_data_delayed_8__11_,chained_data_delayed_8__10_,chained_data_delayed_8__9_,
  chained_data_delayed_8__8_,chained_data_delayed_8__7_,chained_data_delayed_8__6_,
  chained_data_delayed_8__5_,chained_data_delayed_8__4_,chained_data_delayed_8__3_,
  chained_data_delayed_8__2_,chained_data_delayed_8__1_,chained_data_delayed_8__0_,
  chained_data_delayed_7__127_,chained_data_delayed_7__126_,chained_data_delayed_7__125_,
  chained_data_delayed_7__124_,chained_data_delayed_7__123_,chained_data_delayed_7__122_,
  chained_data_delayed_7__121_,chained_data_delayed_7__120_,
  chained_data_delayed_7__119_,chained_data_delayed_7__118_,chained_data_delayed_7__117_,
  chained_data_delayed_7__116_,chained_data_delayed_7__115_,chained_data_delayed_7__114_,
  chained_data_delayed_7__113_,chained_data_delayed_7__112_,chained_data_delayed_7__111_,
  chained_data_delayed_7__110_,chained_data_delayed_7__109_,
  chained_data_delayed_7__108_,chained_data_delayed_7__107_,chained_data_delayed_7__106_,
  chained_data_delayed_7__105_,chained_data_delayed_7__104_,chained_data_delayed_7__103_,
  chained_data_delayed_7__102_,chained_data_delayed_7__101_,chained_data_delayed_7__100_,
  chained_data_delayed_7__99_,chained_data_delayed_7__98_,chained_data_delayed_7__97_,
  chained_data_delayed_7__96_,chained_data_delayed_7__95_,
  chained_data_delayed_7__94_,chained_data_delayed_7__93_,chained_data_delayed_7__92_,
  chained_data_delayed_7__91_,chained_data_delayed_7__90_,chained_data_delayed_7__89_,
  chained_data_delayed_7__88_,chained_data_delayed_7__87_,chained_data_delayed_7__86_,
  chained_data_delayed_7__85_,chained_data_delayed_7__84_,chained_data_delayed_7__83_,
  chained_data_delayed_7__82_,chained_data_delayed_7__81_,chained_data_delayed_7__80_,
  chained_data_delayed_7__79_,chained_data_delayed_7__78_,chained_data_delayed_7__77_,
  chained_data_delayed_7__76_,chained_data_delayed_7__75_,
  chained_data_delayed_7__74_,chained_data_delayed_7__73_,chained_data_delayed_7__72_,
  chained_data_delayed_7__71_,chained_data_delayed_7__70_,chained_data_delayed_7__69_,
  chained_data_delayed_7__68_,chained_data_delayed_7__67_,chained_data_delayed_7__66_,
  chained_data_delayed_7__65_,chained_data_delayed_7__64_,chained_data_delayed_7__63_,
  chained_data_delayed_7__62_,chained_data_delayed_7__61_,chained_data_delayed_7__60_,
  chained_data_delayed_7__59_,chained_data_delayed_7__58_,chained_data_delayed_7__57_,
  chained_data_delayed_7__56_,chained_data_delayed_7__55_,
  chained_data_delayed_7__54_,chained_data_delayed_7__53_,chained_data_delayed_7__52_,
  chained_data_delayed_7__51_,chained_data_delayed_7__50_,chained_data_delayed_7__49_,
  chained_data_delayed_7__48_,chained_data_delayed_7__47_,chained_data_delayed_7__46_,
  chained_data_delayed_7__45_,chained_data_delayed_7__44_,chained_data_delayed_7__43_,
  chained_data_delayed_7__42_,chained_data_delayed_7__41_,chained_data_delayed_7__40_,
  chained_data_delayed_7__39_,chained_data_delayed_7__38_,chained_data_delayed_7__37_,
  chained_data_delayed_7__36_,chained_data_delayed_7__35_,
  chained_data_delayed_7__34_,chained_data_delayed_7__33_,chained_data_delayed_7__32_,
  chained_data_delayed_7__31_,chained_data_delayed_7__30_,chained_data_delayed_7__29_,
  chained_data_delayed_7__28_,chained_data_delayed_7__27_,chained_data_delayed_7__26_,
  chained_data_delayed_7__25_,chained_data_delayed_7__24_,chained_data_delayed_7__23_,
  chained_data_delayed_7__22_,chained_data_delayed_7__21_,chained_data_delayed_7__20_,
  chained_data_delayed_7__19_,chained_data_delayed_7__18_,chained_data_delayed_7__17_,
  chained_data_delayed_7__16_,chained_data_delayed_7__15_,
  chained_data_delayed_7__14_,chained_data_delayed_7__13_,chained_data_delayed_7__12_,
  chained_data_delayed_7__11_,chained_data_delayed_7__10_,chained_data_delayed_7__9_,
  chained_data_delayed_7__8_,chained_data_delayed_7__7_,chained_data_delayed_7__6_,
  chained_data_delayed_7__5_,chained_data_delayed_7__4_,chained_data_delayed_7__3_,
  chained_data_delayed_7__2_,chained_data_delayed_7__1_,chained_data_delayed_7__0_,
  chained_data_delayed_6__127_,chained_data_delayed_6__126_,chained_data_delayed_6__125_,
  chained_data_delayed_6__124_,chained_data_delayed_6__123_,chained_data_delayed_6__122_,
  chained_data_delayed_6__121_,chained_data_delayed_6__120_,
  chained_data_delayed_6__119_,chained_data_delayed_6__118_,chained_data_delayed_6__117_,
  chained_data_delayed_6__116_,chained_data_delayed_6__115_,chained_data_delayed_6__114_,
  chained_data_delayed_6__113_,chained_data_delayed_6__112_,chained_data_delayed_6__111_,
  chained_data_delayed_6__110_,chained_data_delayed_6__109_,
  chained_data_delayed_6__108_,chained_data_delayed_6__107_,chained_data_delayed_6__106_,
  chained_data_delayed_6__105_,chained_data_delayed_6__104_,chained_data_delayed_6__103_,
  chained_data_delayed_6__102_,chained_data_delayed_6__101_,chained_data_delayed_6__100_,
  chained_data_delayed_6__99_,chained_data_delayed_6__98_,
  chained_data_delayed_6__97_,chained_data_delayed_6__96_,chained_data_delayed_6__95_,
  chained_data_delayed_6__94_,chained_data_delayed_6__93_,chained_data_delayed_6__92_,
  chained_data_delayed_6__91_,chained_data_delayed_6__90_,chained_data_delayed_6__89_,
  chained_data_delayed_6__88_,chained_data_delayed_6__87_,chained_data_delayed_6__86_,
  chained_data_delayed_6__85_,chained_data_delayed_6__84_,chained_data_delayed_6__83_,
  chained_data_delayed_6__82_,chained_data_delayed_6__81_,chained_data_delayed_6__80_,
  chained_data_delayed_6__79_,chained_data_delayed_6__78_,
  chained_data_delayed_6__77_,chained_data_delayed_6__76_,chained_data_delayed_6__75_,
  chained_data_delayed_6__74_,chained_data_delayed_6__73_,chained_data_delayed_6__72_,
  chained_data_delayed_6__71_,chained_data_delayed_6__70_,chained_data_delayed_6__69_,
  chained_data_delayed_6__68_,chained_data_delayed_6__67_,chained_data_delayed_6__66_,
  chained_data_delayed_6__65_,chained_data_delayed_6__64_,chained_data_delayed_6__63_,
  chained_data_delayed_6__62_,chained_data_delayed_6__61_,chained_data_delayed_6__60_,
  chained_data_delayed_6__59_,chained_data_delayed_6__58_,
  chained_data_delayed_6__57_,chained_data_delayed_6__56_,chained_data_delayed_6__55_,
  chained_data_delayed_6__54_,chained_data_delayed_6__53_,chained_data_delayed_6__52_,
  chained_data_delayed_6__51_,chained_data_delayed_6__50_,chained_data_delayed_6__49_,
  chained_data_delayed_6__48_,chained_data_delayed_6__47_,chained_data_delayed_6__46_,
  chained_data_delayed_6__45_,chained_data_delayed_6__44_,chained_data_delayed_6__43_,
  chained_data_delayed_6__42_,chained_data_delayed_6__41_,chained_data_delayed_6__40_,
  chained_data_delayed_6__39_,chained_data_delayed_6__38_,
  chained_data_delayed_6__37_,chained_data_delayed_6__36_,chained_data_delayed_6__35_,
  chained_data_delayed_6__34_,chained_data_delayed_6__33_,chained_data_delayed_6__32_,
  chained_data_delayed_6__31_,chained_data_delayed_6__30_,chained_data_delayed_6__29_,
  chained_data_delayed_6__28_,chained_data_delayed_6__27_,chained_data_delayed_6__26_,
  chained_data_delayed_6__25_,chained_data_delayed_6__24_,chained_data_delayed_6__23_,
  chained_data_delayed_6__22_,chained_data_delayed_6__21_,chained_data_delayed_6__20_,
  chained_data_delayed_6__19_,chained_data_delayed_6__18_,
  chained_data_delayed_6__17_,chained_data_delayed_6__16_,chained_data_delayed_6__15_,
  chained_data_delayed_6__14_,chained_data_delayed_6__13_,chained_data_delayed_6__12_,
  chained_data_delayed_6__11_,chained_data_delayed_6__10_,chained_data_delayed_6__9_,
  chained_data_delayed_6__8_,chained_data_delayed_6__7_,chained_data_delayed_6__6_,
  chained_data_delayed_6__5_,chained_data_delayed_6__4_,chained_data_delayed_6__3_,
  chained_data_delayed_6__2_,chained_data_delayed_6__1_,chained_data_delayed_6__0_,
  chained_data_delayed_5__127_,chained_data_delayed_5__126_,chained_data_delayed_5__125_,
  chained_data_delayed_5__124_,chained_data_delayed_5__123_,
  chained_data_delayed_5__122_,chained_data_delayed_5__121_,chained_data_delayed_5__120_,
  chained_data_delayed_5__119_,chained_data_delayed_5__118_,chained_data_delayed_5__117_,
  chained_data_delayed_5__116_,chained_data_delayed_5__115_,chained_data_delayed_5__114_,
  chained_data_delayed_5__113_,chained_data_delayed_5__112_,
  chained_data_delayed_5__111_,chained_data_delayed_5__110_,chained_data_delayed_5__109_,
  chained_data_delayed_5__108_,chained_data_delayed_5__107_,chained_data_delayed_5__106_,
  chained_data_delayed_5__105_,chained_data_delayed_5__104_,chained_data_delayed_5__103_,
  chained_data_delayed_5__102_,chained_data_delayed_5__101_,chained_data_delayed_5__100_,
  chained_data_delayed_5__99_,chained_data_delayed_5__98_,
  chained_data_delayed_5__97_,chained_data_delayed_5__96_,chained_data_delayed_5__95_,
  chained_data_delayed_5__94_,chained_data_delayed_5__93_,chained_data_delayed_5__92_,
  chained_data_delayed_5__91_,chained_data_delayed_5__90_,chained_data_delayed_5__89_,
  chained_data_delayed_5__88_,chained_data_delayed_5__87_,chained_data_delayed_5__86_,
  chained_data_delayed_5__85_,chained_data_delayed_5__84_,chained_data_delayed_5__83_,
  chained_data_delayed_5__82_,chained_data_delayed_5__81_,chained_data_delayed_5__80_,
  chained_data_delayed_5__79_,chained_data_delayed_5__78_,
  chained_data_delayed_5__77_,chained_data_delayed_5__76_,chained_data_delayed_5__75_,
  chained_data_delayed_5__74_,chained_data_delayed_5__73_,chained_data_delayed_5__72_,
  chained_data_delayed_5__71_,chained_data_delayed_5__70_,chained_data_delayed_5__69_,
  chained_data_delayed_5__68_,chained_data_delayed_5__67_,chained_data_delayed_5__66_,
  chained_data_delayed_5__65_,chained_data_delayed_5__64_,chained_data_delayed_5__63_,
  chained_data_delayed_5__62_,chained_data_delayed_5__61_,chained_data_delayed_5__60_,
  chained_data_delayed_5__59_,chained_data_delayed_5__58_,
  chained_data_delayed_5__57_,chained_data_delayed_5__56_,chained_data_delayed_5__55_,
  chained_data_delayed_5__54_,chained_data_delayed_5__53_,chained_data_delayed_5__52_,
  chained_data_delayed_5__51_,chained_data_delayed_5__50_,chained_data_delayed_5__49_,
  chained_data_delayed_5__48_,chained_data_delayed_5__47_,chained_data_delayed_5__46_,
  chained_data_delayed_5__45_,chained_data_delayed_5__44_,chained_data_delayed_5__43_,
  chained_data_delayed_5__42_,chained_data_delayed_5__41_,chained_data_delayed_5__40_,
  chained_data_delayed_5__39_,chained_data_delayed_5__38_,
  chained_data_delayed_5__37_,chained_data_delayed_5__36_,chained_data_delayed_5__35_,
  chained_data_delayed_5__34_,chained_data_delayed_5__33_,chained_data_delayed_5__32_,
  chained_data_delayed_5__31_,chained_data_delayed_5__30_,chained_data_delayed_5__29_,
  chained_data_delayed_5__28_,chained_data_delayed_5__27_,chained_data_delayed_5__26_,
  chained_data_delayed_5__25_,chained_data_delayed_5__24_,chained_data_delayed_5__23_,
  chained_data_delayed_5__22_,chained_data_delayed_5__21_,chained_data_delayed_5__20_,
  chained_data_delayed_5__19_,chained_data_delayed_5__18_,
  chained_data_delayed_5__17_,chained_data_delayed_5__16_,chained_data_delayed_5__15_,
  chained_data_delayed_5__14_,chained_data_delayed_5__13_,chained_data_delayed_5__12_,
  chained_data_delayed_5__11_,chained_data_delayed_5__10_,chained_data_delayed_5__9_,
  chained_data_delayed_5__8_,chained_data_delayed_5__7_,chained_data_delayed_5__6_,
  chained_data_delayed_5__5_,chained_data_delayed_5__4_,chained_data_delayed_5__3_,
  chained_data_delayed_5__2_,chained_data_delayed_5__1_,chained_data_delayed_5__0_,
  chained_data_delayed_12__127_,chained_data_delayed_12__126_,chained_data_delayed_12__125_,
  chained_data_delayed_12__124_,chained_data_delayed_12__123_,
  chained_data_delayed_12__122_,chained_data_delayed_12__121_,chained_data_delayed_12__120_,
  chained_data_delayed_12__119_,chained_data_delayed_12__118_,chained_data_delayed_12__117_,
  chained_data_delayed_12__116_,chained_data_delayed_12__115_,
  chained_data_delayed_12__114_,chained_data_delayed_12__113_,chained_data_delayed_12__112_,
  chained_data_delayed_12__111_,chained_data_delayed_12__110_,chained_data_delayed_12__109_,
  chained_data_delayed_12__108_,chained_data_delayed_12__107_,
  chained_data_delayed_12__106_,chained_data_delayed_12__105_,chained_data_delayed_12__104_,
  chained_data_delayed_12__103_,chained_data_delayed_12__102_,chained_data_delayed_12__101_,
  chained_data_delayed_12__100_,chained_data_delayed_12__99_,
  chained_data_delayed_12__98_,chained_data_delayed_12__97_,chained_data_delayed_12__96_,
  chained_data_delayed_12__95_,chained_data_delayed_12__94_,chained_data_delayed_12__93_,
  chained_data_delayed_12__92_,chained_data_delayed_12__91_,chained_data_delayed_12__90_,
  chained_data_delayed_12__89_,chained_data_delayed_12__88_,
  chained_data_delayed_12__87_,chained_data_delayed_12__86_,chained_data_delayed_12__85_,
  chained_data_delayed_12__84_,chained_data_delayed_12__83_,chained_data_delayed_12__82_,
  chained_data_delayed_12__81_,chained_data_delayed_12__80_,chained_data_delayed_12__79_,
  chained_data_delayed_12__78_,chained_data_delayed_12__77_,
  chained_data_delayed_12__76_,chained_data_delayed_12__75_,chained_data_delayed_12__74_,
  chained_data_delayed_12__73_,chained_data_delayed_12__72_,chained_data_delayed_12__71_,
  chained_data_delayed_12__70_,chained_data_delayed_12__69_,chained_data_delayed_12__68_,
  chained_data_delayed_12__67_,chained_data_delayed_12__66_,
  chained_data_delayed_12__65_,chained_data_delayed_12__64_,chained_data_delayed_12__63_,
  chained_data_delayed_12__62_,chained_data_delayed_12__61_,chained_data_delayed_12__60_,
  chained_data_delayed_12__59_,chained_data_delayed_12__58_,chained_data_delayed_12__57_,
  chained_data_delayed_12__56_,chained_data_delayed_12__55_,
  chained_data_delayed_12__54_,chained_data_delayed_12__53_,chained_data_delayed_12__52_,
  chained_data_delayed_12__51_,chained_data_delayed_12__50_,chained_data_delayed_12__49_,
  chained_data_delayed_12__48_,chained_data_delayed_12__47_,chained_data_delayed_12__46_,
  chained_data_delayed_12__45_,chained_data_delayed_12__44_,
  chained_data_delayed_12__43_,chained_data_delayed_12__42_,chained_data_delayed_12__41_,
  chained_data_delayed_12__40_,chained_data_delayed_12__39_,chained_data_delayed_12__38_,
  chained_data_delayed_12__37_,chained_data_delayed_12__36_,chained_data_delayed_12__35_,
  chained_data_delayed_12__34_,chained_data_delayed_12__33_,
  chained_data_delayed_12__32_,chained_data_delayed_12__31_,chained_data_delayed_12__30_,
  chained_data_delayed_12__29_,chained_data_delayed_12__28_,chained_data_delayed_12__27_,
  chained_data_delayed_12__26_,chained_data_delayed_12__25_,chained_data_delayed_12__24_,
  chained_data_delayed_12__23_,chained_data_delayed_12__22_,
  chained_data_delayed_12__21_,chained_data_delayed_12__20_,chained_data_delayed_12__19_,
  chained_data_delayed_12__18_,chained_data_delayed_12__17_,chained_data_delayed_12__16_,
  chained_data_delayed_12__15_,chained_data_delayed_12__14_,chained_data_delayed_12__13_,
  chained_data_delayed_12__12_,chained_data_delayed_12__11_,chained_data_delayed_12__10_,
  chained_data_delayed_12__9_,chained_data_delayed_12__8_,
  chained_data_delayed_12__7_,chained_data_delayed_12__6_,chained_data_delayed_12__5_,
  chained_data_delayed_12__4_,chained_data_delayed_12__3_,chained_data_delayed_12__2_,
  chained_data_delayed_12__1_,chained_data_delayed_12__0_,chained_data_delayed_11__127_,
  chained_data_delayed_11__126_,chained_data_delayed_11__125_,chained_data_delayed_11__124_,
  chained_data_delayed_11__123_,chained_data_delayed_11__122_,
  chained_data_delayed_11__121_,chained_data_delayed_11__120_,chained_data_delayed_11__119_,
  chained_data_delayed_11__118_,chained_data_delayed_11__117_,chained_data_delayed_11__116_,
  chained_data_delayed_11__115_,chained_data_delayed_11__114_,
  chained_data_delayed_11__113_,chained_data_delayed_11__112_,chained_data_delayed_11__111_,
  chained_data_delayed_11__110_,chained_data_delayed_11__109_,chained_data_delayed_11__108_,
  chained_data_delayed_11__107_,chained_data_delayed_11__106_,
  chained_data_delayed_11__105_,chained_data_delayed_11__104_,chained_data_delayed_11__103_,
  chained_data_delayed_11__102_,chained_data_delayed_11__101_,chained_data_delayed_11__100_,
  chained_data_delayed_11__99_,chained_data_delayed_11__98_,
  chained_data_delayed_11__97_,chained_data_delayed_11__96_,chained_data_delayed_11__95_,
  chained_data_delayed_11__94_,chained_data_delayed_11__93_,chained_data_delayed_11__92_,
  chained_data_delayed_11__91_,chained_data_delayed_11__90_,chained_data_delayed_11__89_,
  chained_data_delayed_11__88_,chained_data_delayed_11__87_,
  chained_data_delayed_11__86_,chained_data_delayed_11__85_,chained_data_delayed_11__84_,
  chained_data_delayed_11__83_,chained_data_delayed_11__82_,chained_data_delayed_11__81_,
  chained_data_delayed_11__80_,chained_data_delayed_11__79_,chained_data_delayed_11__78_,
  chained_data_delayed_11__77_,chained_data_delayed_11__76_,
  chained_data_delayed_11__75_,chained_data_delayed_11__74_,chained_data_delayed_11__73_,
  chained_data_delayed_11__72_,chained_data_delayed_11__71_,chained_data_delayed_11__70_,
  chained_data_delayed_11__69_,chained_data_delayed_11__68_,chained_data_delayed_11__67_,
  chained_data_delayed_11__66_,chained_data_delayed_11__65_,
  chained_data_delayed_11__64_,chained_data_delayed_11__63_,chained_data_delayed_11__62_,
  chained_data_delayed_11__61_,chained_data_delayed_11__60_,chained_data_delayed_11__59_,
  chained_data_delayed_11__58_,chained_data_delayed_11__57_,chained_data_delayed_11__56_,
  chained_data_delayed_11__55_,chained_data_delayed_11__54_,
  chained_data_delayed_11__53_,chained_data_delayed_11__52_,chained_data_delayed_11__51_,
  chained_data_delayed_11__50_,chained_data_delayed_11__49_,chained_data_delayed_11__48_,
  chained_data_delayed_11__47_,chained_data_delayed_11__46_,chained_data_delayed_11__45_,
  chained_data_delayed_11__44_,chained_data_delayed_11__43_,
  chained_data_delayed_11__42_,chained_data_delayed_11__41_,chained_data_delayed_11__40_,
  chained_data_delayed_11__39_,chained_data_delayed_11__38_,chained_data_delayed_11__37_,
  chained_data_delayed_11__36_,chained_data_delayed_11__35_,chained_data_delayed_11__34_,
  chained_data_delayed_11__33_,chained_data_delayed_11__32_,
  chained_data_delayed_11__31_,chained_data_delayed_11__30_,chained_data_delayed_11__29_,
  chained_data_delayed_11__28_,chained_data_delayed_11__27_,chained_data_delayed_11__26_,
  chained_data_delayed_11__25_,chained_data_delayed_11__24_,chained_data_delayed_11__23_,
  chained_data_delayed_11__22_,chained_data_delayed_11__21_,chained_data_delayed_11__20_,
  chained_data_delayed_11__19_,chained_data_delayed_11__18_,
  chained_data_delayed_11__17_,chained_data_delayed_11__16_,chained_data_delayed_11__15_,
  chained_data_delayed_11__14_,chained_data_delayed_11__13_,chained_data_delayed_11__12_,
  chained_data_delayed_11__11_,chained_data_delayed_11__10_,chained_data_delayed_11__9_,
  chained_data_delayed_11__8_,chained_data_delayed_11__7_,
  chained_data_delayed_11__6_,chained_data_delayed_11__5_,chained_data_delayed_11__4_,
  chained_data_delayed_11__3_,chained_data_delayed_11__2_,chained_data_delayed_11__1_,
  chained_data_delayed_11__0_,chained_data_delayed_10__127_,chained_data_delayed_10__126_,
  chained_data_delayed_10__125_,chained_data_delayed_10__124_,chained_data_delayed_10__123_,
  chained_data_delayed_10__122_,chained_data_delayed_10__121_,
  chained_data_delayed_10__120_,chained_data_delayed_10__119_,chained_data_delayed_10__118_,
  chained_data_delayed_10__117_,chained_data_delayed_10__116_,chained_data_delayed_10__115_,
  chained_data_delayed_10__114_,chained_data_delayed_10__113_,
  chained_data_delayed_10__112_,chained_data_delayed_10__111_,chained_data_delayed_10__110_,
  chained_data_delayed_10__109_,chained_data_delayed_10__108_,chained_data_delayed_10__107_,
  chained_data_delayed_10__106_,chained_data_delayed_10__105_,
  chained_data_delayed_10__104_,chained_data_delayed_10__103_,chained_data_delayed_10__102_,
  chained_data_delayed_10__101_,chained_data_delayed_10__100_,chained_data_delayed_10__99_,
  chained_data_delayed_10__98_,chained_data_delayed_10__97_,
  chained_data_delayed_10__96_,chained_data_delayed_10__95_,chained_data_delayed_10__94_,
  chained_data_delayed_10__93_,chained_data_delayed_10__92_,chained_data_delayed_10__91_,
  chained_data_delayed_10__90_,chained_data_delayed_10__89_,chained_data_delayed_10__88_,
  chained_data_delayed_10__87_,chained_data_delayed_10__86_,
  chained_data_delayed_10__85_,chained_data_delayed_10__84_,chained_data_delayed_10__83_,
  chained_data_delayed_10__82_,chained_data_delayed_10__81_,chained_data_delayed_10__80_,
  chained_data_delayed_10__79_,chained_data_delayed_10__78_,chained_data_delayed_10__77_,
  chained_data_delayed_10__76_,chained_data_delayed_10__75_,
  chained_data_delayed_10__74_,chained_data_delayed_10__73_,chained_data_delayed_10__72_,
  chained_data_delayed_10__71_,chained_data_delayed_10__70_,chained_data_delayed_10__69_,
  chained_data_delayed_10__68_,chained_data_delayed_10__67_,chained_data_delayed_10__66_,
  chained_data_delayed_10__65_,chained_data_delayed_10__64_,
  chained_data_delayed_10__63_,chained_data_delayed_10__62_,chained_data_delayed_10__61_,
  chained_data_delayed_10__60_,chained_data_delayed_10__59_,chained_data_delayed_10__58_,
  chained_data_delayed_10__57_,chained_data_delayed_10__56_,chained_data_delayed_10__55_,
  chained_data_delayed_10__54_,chained_data_delayed_10__53_,
  chained_data_delayed_10__52_,chained_data_delayed_10__51_,chained_data_delayed_10__50_,
  chained_data_delayed_10__49_,chained_data_delayed_10__48_,chained_data_delayed_10__47_,
  chained_data_delayed_10__46_,chained_data_delayed_10__45_,chained_data_delayed_10__44_,
  chained_data_delayed_10__43_,chained_data_delayed_10__42_,
  chained_data_delayed_10__41_,chained_data_delayed_10__40_,chained_data_delayed_10__39_,
  chained_data_delayed_10__38_,chained_data_delayed_10__37_,chained_data_delayed_10__36_,
  chained_data_delayed_10__35_,chained_data_delayed_10__34_,chained_data_delayed_10__33_,
  chained_data_delayed_10__32_,chained_data_delayed_10__31_,chained_data_delayed_10__30_,
  chained_data_delayed_10__29_,chained_data_delayed_10__28_,
  chained_data_delayed_10__27_,chained_data_delayed_10__26_,chained_data_delayed_10__25_,
  chained_data_delayed_10__24_,chained_data_delayed_10__23_,chained_data_delayed_10__22_,
  chained_data_delayed_10__21_,chained_data_delayed_10__20_,chained_data_delayed_10__19_,
  chained_data_delayed_10__18_,chained_data_delayed_10__17_,
  chained_data_delayed_10__16_,chained_data_delayed_10__15_,chained_data_delayed_10__14_,
  chained_data_delayed_10__13_,chained_data_delayed_10__12_,chained_data_delayed_10__11_,
  chained_data_delayed_10__10_,chained_data_delayed_10__9_,chained_data_delayed_10__8_,
  chained_data_delayed_10__7_,chained_data_delayed_10__6_,chained_data_delayed_10__5_,
  chained_data_delayed_10__4_,chained_data_delayed_10__3_,
  chained_data_delayed_10__2_,chained_data_delayed_10__1_,chained_data_delayed_10__0_,
  chained_data_delayed_9__127_,chained_data_delayed_9__126_,chained_data_delayed_9__125_,
  chained_data_delayed_9__124_,chained_data_delayed_9__123_,chained_data_delayed_9__122_,
  chained_data_delayed_9__121_,chained_data_delayed_9__120_,
  chained_data_delayed_9__119_,chained_data_delayed_9__118_,chained_data_delayed_9__117_,
  chained_data_delayed_9__116_,chained_data_delayed_9__115_,chained_data_delayed_9__114_,
  chained_data_delayed_9__113_,chained_data_delayed_9__112_,chained_data_delayed_9__111_,
  chained_data_delayed_9__110_,chained_data_delayed_9__109_,chained_data_delayed_9__108_,
  chained_data_delayed_9__107_,chained_data_delayed_9__106_,
  chained_data_delayed_9__105_,chained_data_delayed_9__104_,chained_data_delayed_9__103_,
  chained_data_delayed_9__102_,chained_data_delayed_9__101_,chained_data_delayed_9__100_,
  chained_data_delayed_9__99_,chained_data_delayed_9__98_,chained_data_delayed_9__97_,
  chained_data_delayed_9__96_,chained_data_delayed_9__95_,chained_data_delayed_9__94_,
  chained_data_delayed_9__93_,chained_data_delayed_9__92_,
  chained_data_delayed_9__91_,chained_data_delayed_9__90_,chained_data_delayed_9__89_,
  chained_data_delayed_9__88_,chained_data_delayed_9__87_,chained_data_delayed_9__86_,
  chained_data_delayed_9__85_,chained_data_delayed_9__84_,chained_data_delayed_9__83_,
  chained_data_delayed_9__82_,chained_data_delayed_9__81_,chained_data_delayed_9__80_,
  chained_data_delayed_9__79_,chained_data_delayed_9__78_,chained_data_delayed_9__77_,
  chained_data_delayed_9__76_,chained_data_delayed_9__75_,chained_data_delayed_9__74_,
  chained_data_delayed_9__73_,chained_data_delayed_9__72_,
  chained_data_delayed_9__71_,chained_data_delayed_9__70_,chained_data_delayed_9__69_,
  chained_data_delayed_9__68_,chained_data_delayed_9__67_,chained_data_delayed_9__66_,
  chained_data_delayed_9__65_,chained_data_delayed_9__64_,chained_data_delayed_9__63_,
  chained_data_delayed_9__62_,chained_data_delayed_9__61_,chained_data_delayed_9__60_,
  chained_data_delayed_9__59_,chained_data_delayed_9__58_,chained_data_delayed_9__57_,
  chained_data_delayed_9__56_,chained_data_delayed_9__55_,chained_data_delayed_9__54_,
  chained_data_delayed_9__53_,chained_data_delayed_9__52_,
  chained_data_delayed_9__51_,chained_data_delayed_9__50_,chained_data_delayed_9__49_,
  chained_data_delayed_9__48_,chained_data_delayed_9__47_,chained_data_delayed_9__46_,
  chained_data_delayed_9__45_,chained_data_delayed_9__44_,chained_data_delayed_9__43_,
  chained_data_delayed_9__42_,chained_data_delayed_9__41_,chained_data_delayed_9__40_,
  chained_data_delayed_9__39_,chained_data_delayed_9__38_,chained_data_delayed_9__37_,
  chained_data_delayed_9__36_,chained_data_delayed_9__35_,chained_data_delayed_9__34_,
  chained_data_delayed_9__33_,chained_data_delayed_9__32_,
  chained_data_delayed_9__31_,chained_data_delayed_9__30_,chained_data_delayed_9__29_,
  chained_data_delayed_9__28_,chained_data_delayed_9__27_,chained_data_delayed_9__26_,
  chained_data_delayed_9__25_,chained_data_delayed_9__24_,chained_data_delayed_9__23_,
  chained_data_delayed_9__22_,chained_data_delayed_9__21_,chained_data_delayed_9__20_,
  chained_data_delayed_9__19_,chained_data_delayed_9__18_,chained_data_delayed_9__17_,
  chained_data_delayed_9__16_,chained_data_delayed_9__15_,chained_data_delayed_9__14_,
  chained_data_delayed_9__13_,chained_data_delayed_9__12_,
  chained_data_delayed_9__11_,chained_data_delayed_9__10_,chained_data_delayed_9__9_,
  chained_data_delayed_9__8_,chained_data_delayed_9__7_,chained_data_delayed_9__6_,
  chained_data_delayed_9__5_,chained_data_delayed_9__4_,chained_data_delayed_9__3_,
  chained_data_delayed_9__2_,chained_data_delayed_9__1_,chained_data_delayed_9__0_,
  chained_data_delayed_16__127_,chained_data_delayed_16__126_,chained_data_delayed_16__125_,
  chained_data_delayed_16__124_,chained_data_delayed_16__123_,
  chained_data_delayed_16__122_,chained_data_delayed_16__121_,chained_data_delayed_16__120_,
  chained_data_delayed_16__119_,chained_data_delayed_16__118_,chained_data_delayed_16__117_,
  chained_data_delayed_16__116_,chained_data_delayed_16__115_,
  chained_data_delayed_16__114_,chained_data_delayed_16__113_,chained_data_delayed_16__112_,
  chained_data_delayed_16__111_,chained_data_delayed_16__110_,chained_data_delayed_16__109_,
  chained_data_delayed_16__108_,chained_data_delayed_16__107_,
  chained_data_delayed_16__106_,chained_data_delayed_16__105_,chained_data_delayed_16__104_,
  chained_data_delayed_16__103_,chained_data_delayed_16__102_,chained_data_delayed_16__101_,
  chained_data_delayed_16__100_,chained_data_delayed_16__99_,chained_data_delayed_16__98_,
  chained_data_delayed_16__97_,chained_data_delayed_16__96_,
  chained_data_delayed_16__95_,chained_data_delayed_16__94_,chained_data_delayed_16__93_,
  chained_data_delayed_16__92_,chained_data_delayed_16__91_,chained_data_delayed_16__90_,
  chained_data_delayed_16__89_,chained_data_delayed_16__88_,chained_data_delayed_16__87_,
  chained_data_delayed_16__86_,chained_data_delayed_16__85_,
  chained_data_delayed_16__84_,chained_data_delayed_16__83_,chained_data_delayed_16__82_,
  chained_data_delayed_16__81_,chained_data_delayed_16__80_,chained_data_delayed_16__79_,
  chained_data_delayed_16__78_,chained_data_delayed_16__77_,chained_data_delayed_16__76_,
  chained_data_delayed_16__75_,chained_data_delayed_16__74_,
  chained_data_delayed_16__73_,chained_data_delayed_16__72_,chained_data_delayed_16__71_,
  chained_data_delayed_16__70_,chained_data_delayed_16__69_,chained_data_delayed_16__68_,
  chained_data_delayed_16__67_,chained_data_delayed_16__66_,chained_data_delayed_16__65_,
  chained_data_delayed_16__64_,chained_data_delayed_16__63_,
  chained_data_delayed_16__62_,chained_data_delayed_16__61_,chained_data_delayed_16__60_,
  chained_data_delayed_16__59_,chained_data_delayed_16__58_,chained_data_delayed_16__57_,
  chained_data_delayed_16__56_,chained_data_delayed_16__55_,chained_data_delayed_16__54_,
  chained_data_delayed_16__53_,chained_data_delayed_16__52_,
  chained_data_delayed_16__51_,chained_data_delayed_16__50_,chained_data_delayed_16__49_,
  chained_data_delayed_16__48_,chained_data_delayed_16__47_,chained_data_delayed_16__46_,
  chained_data_delayed_16__45_,chained_data_delayed_16__44_,chained_data_delayed_16__43_,
  chained_data_delayed_16__42_,chained_data_delayed_16__41_,
  chained_data_delayed_16__40_,chained_data_delayed_16__39_,chained_data_delayed_16__38_,
  chained_data_delayed_16__37_,chained_data_delayed_16__36_,chained_data_delayed_16__35_,
  chained_data_delayed_16__34_,chained_data_delayed_16__33_,chained_data_delayed_16__32_,
  chained_data_delayed_16__31_,chained_data_delayed_16__30_,
  chained_data_delayed_16__29_,chained_data_delayed_16__28_,chained_data_delayed_16__27_,
  chained_data_delayed_16__26_,chained_data_delayed_16__25_,chained_data_delayed_16__24_,
  chained_data_delayed_16__23_,chained_data_delayed_16__22_,chained_data_delayed_16__21_,
  chained_data_delayed_16__20_,chained_data_delayed_16__19_,chained_data_delayed_16__18_,
  chained_data_delayed_16__17_,chained_data_delayed_16__16_,
  chained_data_delayed_16__15_,chained_data_delayed_16__14_,chained_data_delayed_16__13_,
  chained_data_delayed_16__12_,chained_data_delayed_16__11_,chained_data_delayed_16__10_,
  chained_data_delayed_16__9_,chained_data_delayed_16__8_,chained_data_delayed_16__7_,
  chained_data_delayed_16__6_,chained_data_delayed_16__5_,chained_data_delayed_16__4_,
  chained_data_delayed_16__3_,chained_data_delayed_16__2_,
  chained_data_delayed_16__1_,chained_data_delayed_16__0_,chained_data_delayed_15__127_,
  chained_data_delayed_15__126_,chained_data_delayed_15__125_,chained_data_delayed_15__124_,
  chained_data_delayed_15__123_,chained_data_delayed_15__122_,
  chained_data_delayed_15__121_,chained_data_delayed_15__120_,chained_data_delayed_15__119_,
  chained_data_delayed_15__118_,chained_data_delayed_15__117_,chained_data_delayed_15__116_,
  chained_data_delayed_15__115_,chained_data_delayed_15__114_,
  chained_data_delayed_15__113_,chained_data_delayed_15__112_,chained_data_delayed_15__111_,
  chained_data_delayed_15__110_,chained_data_delayed_15__109_,chained_data_delayed_15__108_,
  chained_data_delayed_15__107_,chained_data_delayed_15__106_,
  chained_data_delayed_15__105_,chained_data_delayed_15__104_,chained_data_delayed_15__103_,
  chained_data_delayed_15__102_,chained_data_delayed_15__101_,chained_data_delayed_15__100_,
  chained_data_delayed_15__99_,chained_data_delayed_15__98_,chained_data_delayed_15__97_,
  chained_data_delayed_15__96_,chained_data_delayed_15__95_,
  chained_data_delayed_15__94_,chained_data_delayed_15__93_,chained_data_delayed_15__92_,
  chained_data_delayed_15__91_,chained_data_delayed_15__90_,chained_data_delayed_15__89_,
  chained_data_delayed_15__88_,chained_data_delayed_15__87_,chained_data_delayed_15__86_,
  chained_data_delayed_15__85_,chained_data_delayed_15__84_,
  chained_data_delayed_15__83_,chained_data_delayed_15__82_,chained_data_delayed_15__81_,
  chained_data_delayed_15__80_,chained_data_delayed_15__79_,chained_data_delayed_15__78_,
  chained_data_delayed_15__77_,chained_data_delayed_15__76_,chained_data_delayed_15__75_,
  chained_data_delayed_15__74_,chained_data_delayed_15__73_,
  chained_data_delayed_15__72_,chained_data_delayed_15__71_,chained_data_delayed_15__70_,
  chained_data_delayed_15__69_,chained_data_delayed_15__68_,chained_data_delayed_15__67_,
  chained_data_delayed_15__66_,chained_data_delayed_15__65_,chained_data_delayed_15__64_,
  chained_data_delayed_15__63_,chained_data_delayed_15__62_,
  chained_data_delayed_15__61_,chained_data_delayed_15__60_,chained_data_delayed_15__59_,
  chained_data_delayed_15__58_,chained_data_delayed_15__57_,chained_data_delayed_15__56_,
  chained_data_delayed_15__55_,chained_data_delayed_15__54_,chained_data_delayed_15__53_,
  chained_data_delayed_15__52_,chained_data_delayed_15__51_,
  chained_data_delayed_15__50_,chained_data_delayed_15__49_,chained_data_delayed_15__48_,
  chained_data_delayed_15__47_,chained_data_delayed_15__46_,chained_data_delayed_15__45_,
  chained_data_delayed_15__44_,chained_data_delayed_15__43_,chained_data_delayed_15__42_,
  chained_data_delayed_15__41_,chained_data_delayed_15__40_,
  chained_data_delayed_15__39_,chained_data_delayed_15__38_,chained_data_delayed_15__37_,
  chained_data_delayed_15__36_,chained_data_delayed_15__35_,chained_data_delayed_15__34_,
  chained_data_delayed_15__33_,chained_data_delayed_15__32_,chained_data_delayed_15__31_,
  chained_data_delayed_15__30_,chained_data_delayed_15__29_,chained_data_delayed_15__28_,
  chained_data_delayed_15__27_,chained_data_delayed_15__26_,
  chained_data_delayed_15__25_,chained_data_delayed_15__24_,chained_data_delayed_15__23_,
  chained_data_delayed_15__22_,chained_data_delayed_15__21_,chained_data_delayed_15__20_,
  chained_data_delayed_15__19_,chained_data_delayed_15__18_,chained_data_delayed_15__17_,
  chained_data_delayed_15__16_,chained_data_delayed_15__15_,
  chained_data_delayed_15__14_,chained_data_delayed_15__13_,chained_data_delayed_15__12_,
  chained_data_delayed_15__11_,chained_data_delayed_15__10_,chained_data_delayed_15__9_,
  chained_data_delayed_15__8_,chained_data_delayed_15__7_,chained_data_delayed_15__6_,
  chained_data_delayed_15__5_,chained_data_delayed_15__4_,chained_data_delayed_15__3_,
  chained_data_delayed_15__2_,chained_data_delayed_15__1_,
  chained_data_delayed_15__0_,chained_data_delayed_14__127_,chained_data_delayed_14__126_,
  chained_data_delayed_14__125_,chained_data_delayed_14__124_,chained_data_delayed_14__123_,
  chained_data_delayed_14__122_,chained_data_delayed_14__121_,
  chained_data_delayed_14__120_,chained_data_delayed_14__119_,chained_data_delayed_14__118_,
  chained_data_delayed_14__117_,chained_data_delayed_14__116_,chained_data_delayed_14__115_,
  chained_data_delayed_14__114_,chained_data_delayed_14__113_,
  chained_data_delayed_14__112_,chained_data_delayed_14__111_,chained_data_delayed_14__110_,
  chained_data_delayed_14__109_,chained_data_delayed_14__108_,chained_data_delayed_14__107_,
  chained_data_delayed_14__106_,chained_data_delayed_14__105_,
  chained_data_delayed_14__104_,chained_data_delayed_14__103_,chained_data_delayed_14__102_,
  chained_data_delayed_14__101_,chained_data_delayed_14__100_,chained_data_delayed_14__99_,
  chained_data_delayed_14__98_,chained_data_delayed_14__97_,chained_data_delayed_14__96_,
  chained_data_delayed_14__95_,chained_data_delayed_14__94_,
  chained_data_delayed_14__93_,chained_data_delayed_14__92_,chained_data_delayed_14__91_,
  chained_data_delayed_14__90_,chained_data_delayed_14__89_,chained_data_delayed_14__88_,
  chained_data_delayed_14__87_,chained_data_delayed_14__86_,chained_data_delayed_14__85_,
  chained_data_delayed_14__84_,chained_data_delayed_14__83_,
  chained_data_delayed_14__82_,chained_data_delayed_14__81_,chained_data_delayed_14__80_,
  chained_data_delayed_14__79_,chained_data_delayed_14__78_,chained_data_delayed_14__77_,
  chained_data_delayed_14__76_,chained_data_delayed_14__75_,chained_data_delayed_14__74_,
  chained_data_delayed_14__73_,chained_data_delayed_14__72_,
  chained_data_delayed_14__71_,chained_data_delayed_14__70_,chained_data_delayed_14__69_,
  chained_data_delayed_14__68_,chained_data_delayed_14__67_,chained_data_delayed_14__66_,
  chained_data_delayed_14__65_,chained_data_delayed_14__64_,chained_data_delayed_14__63_,
  chained_data_delayed_14__62_,chained_data_delayed_14__61_,
  chained_data_delayed_14__60_,chained_data_delayed_14__59_,chained_data_delayed_14__58_,
  chained_data_delayed_14__57_,chained_data_delayed_14__56_,chained_data_delayed_14__55_,
  chained_data_delayed_14__54_,chained_data_delayed_14__53_,chained_data_delayed_14__52_,
  chained_data_delayed_14__51_,chained_data_delayed_14__50_,
  chained_data_delayed_14__49_,chained_data_delayed_14__48_,chained_data_delayed_14__47_,
  chained_data_delayed_14__46_,chained_data_delayed_14__45_,chained_data_delayed_14__44_,
  chained_data_delayed_14__43_,chained_data_delayed_14__42_,chained_data_delayed_14__41_,
  chained_data_delayed_14__40_,chained_data_delayed_14__39_,chained_data_delayed_14__38_,
  chained_data_delayed_14__37_,chained_data_delayed_14__36_,
  chained_data_delayed_14__35_,chained_data_delayed_14__34_,chained_data_delayed_14__33_,
  chained_data_delayed_14__32_,chained_data_delayed_14__31_,chained_data_delayed_14__30_,
  chained_data_delayed_14__29_,chained_data_delayed_14__28_,chained_data_delayed_14__27_,
  chained_data_delayed_14__26_,chained_data_delayed_14__25_,
  chained_data_delayed_14__24_,chained_data_delayed_14__23_,chained_data_delayed_14__22_,
  chained_data_delayed_14__21_,chained_data_delayed_14__20_,chained_data_delayed_14__19_,
  chained_data_delayed_14__18_,chained_data_delayed_14__17_,chained_data_delayed_14__16_,
  chained_data_delayed_14__15_,chained_data_delayed_14__14_,
  chained_data_delayed_14__13_,chained_data_delayed_14__12_,chained_data_delayed_14__11_,
  chained_data_delayed_14__10_,chained_data_delayed_14__9_,chained_data_delayed_14__8_,
  chained_data_delayed_14__7_,chained_data_delayed_14__6_,chained_data_delayed_14__5_,
  chained_data_delayed_14__4_,chained_data_delayed_14__3_,chained_data_delayed_14__2_,
  chained_data_delayed_14__1_,chained_data_delayed_14__0_,
  chained_data_delayed_13__127_,chained_data_delayed_13__126_,chained_data_delayed_13__125_,
  chained_data_delayed_13__124_,chained_data_delayed_13__123_,chained_data_delayed_13__122_,
  chained_data_delayed_13__121_,chained_data_delayed_13__120_,
  chained_data_delayed_13__119_,chained_data_delayed_13__118_,chained_data_delayed_13__117_,
  chained_data_delayed_13__116_,chained_data_delayed_13__115_,chained_data_delayed_13__114_,
  chained_data_delayed_13__113_,chained_data_delayed_13__112_,
  chained_data_delayed_13__111_,chained_data_delayed_13__110_,chained_data_delayed_13__109_,
  chained_data_delayed_13__108_,chained_data_delayed_13__107_,chained_data_delayed_13__106_,
  chained_data_delayed_13__105_,chained_data_delayed_13__104_,
  chained_data_delayed_13__103_,chained_data_delayed_13__102_,chained_data_delayed_13__101_,
  chained_data_delayed_13__100_,chained_data_delayed_13__99_,chained_data_delayed_13__98_,
  chained_data_delayed_13__97_,chained_data_delayed_13__96_,chained_data_delayed_13__95_,
  chained_data_delayed_13__94_,chained_data_delayed_13__93_,
  chained_data_delayed_13__92_,chained_data_delayed_13__91_,chained_data_delayed_13__90_,
  chained_data_delayed_13__89_,chained_data_delayed_13__88_,chained_data_delayed_13__87_,
  chained_data_delayed_13__86_,chained_data_delayed_13__85_,chained_data_delayed_13__84_,
  chained_data_delayed_13__83_,chained_data_delayed_13__82_,
  chained_data_delayed_13__81_,chained_data_delayed_13__80_,chained_data_delayed_13__79_,
  chained_data_delayed_13__78_,chained_data_delayed_13__77_,chained_data_delayed_13__76_,
  chained_data_delayed_13__75_,chained_data_delayed_13__74_,chained_data_delayed_13__73_,
  chained_data_delayed_13__72_,chained_data_delayed_13__71_,
  chained_data_delayed_13__70_,chained_data_delayed_13__69_,chained_data_delayed_13__68_,
  chained_data_delayed_13__67_,chained_data_delayed_13__66_,chained_data_delayed_13__65_,
  chained_data_delayed_13__64_,chained_data_delayed_13__63_,chained_data_delayed_13__62_,
  chained_data_delayed_13__61_,chained_data_delayed_13__60_,
  chained_data_delayed_13__59_,chained_data_delayed_13__58_,chained_data_delayed_13__57_,
  chained_data_delayed_13__56_,chained_data_delayed_13__55_,chained_data_delayed_13__54_,
  chained_data_delayed_13__53_,chained_data_delayed_13__52_,chained_data_delayed_13__51_,
  chained_data_delayed_13__50_,chained_data_delayed_13__49_,chained_data_delayed_13__48_,
  chained_data_delayed_13__47_,chained_data_delayed_13__46_,
  chained_data_delayed_13__45_,chained_data_delayed_13__44_,chained_data_delayed_13__43_,
  chained_data_delayed_13__42_,chained_data_delayed_13__41_,chained_data_delayed_13__40_,
  chained_data_delayed_13__39_,chained_data_delayed_13__38_,chained_data_delayed_13__37_,
  chained_data_delayed_13__36_,chained_data_delayed_13__35_,
  chained_data_delayed_13__34_,chained_data_delayed_13__33_,chained_data_delayed_13__32_,
  chained_data_delayed_13__31_,chained_data_delayed_13__30_,chained_data_delayed_13__29_,
  chained_data_delayed_13__28_,chained_data_delayed_13__27_,chained_data_delayed_13__26_,
  chained_data_delayed_13__25_,chained_data_delayed_13__24_,
  chained_data_delayed_13__23_,chained_data_delayed_13__22_,chained_data_delayed_13__21_,
  chained_data_delayed_13__20_,chained_data_delayed_13__19_,chained_data_delayed_13__18_,
  chained_data_delayed_13__17_,chained_data_delayed_13__16_,chained_data_delayed_13__15_,
  chained_data_delayed_13__14_,chained_data_delayed_13__13_,
  chained_data_delayed_13__12_,chained_data_delayed_13__11_,chained_data_delayed_13__10_,
  chained_data_delayed_13__9_,chained_data_delayed_13__8_,chained_data_delayed_13__7_,
  chained_data_delayed_13__6_,chained_data_delayed_13__5_,chained_data_delayed_13__4_,
  chained_data_delayed_13__3_,chained_data_delayed_13__2_,chained_data_delayed_13__1_,
  chained_data_delayed_13__0_,chained_data_delayed_20__127_,
  chained_data_delayed_20__126_,chained_data_delayed_20__125_,chained_data_delayed_20__124_,
  chained_data_delayed_20__123_,chained_data_delayed_20__122_,chained_data_delayed_20__121_,
  chained_data_delayed_20__120_,chained_data_delayed_20__119_,
  chained_data_delayed_20__118_,chained_data_delayed_20__117_,chained_data_delayed_20__116_,
  chained_data_delayed_20__115_,chained_data_delayed_20__114_,chained_data_delayed_20__113_,
  chained_data_delayed_20__112_,chained_data_delayed_20__111_,
  chained_data_delayed_20__110_,chained_data_delayed_20__109_,chained_data_delayed_20__108_,
  chained_data_delayed_20__107_,chained_data_delayed_20__106_,chained_data_delayed_20__105_,
  chained_data_delayed_20__104_,chained_data_delayed_20__103_,
  chained_data_delayed_20__102_,chained_data_delayed_20__101_,chained_data_delayed_20__100_,
  chained_data_delayed_20__99_,chained_data_delayed_20__98_,chained_data_delayed_20__97_,
  chained_data_delayed_20__96_,chained_data_delayed_20__95_,chained_data_delayed_20__94_,
  chained_data_delayed_20__93_,chained_data_delayed_20__92_,
  chained_data_delayed_20__91_,chained_data_delayed_20__90_,chained_data_delayed_20__89_,
  chained_data_delayed_20__88_,chained_data_delayed_20__87_,chained_data_delayed_20__86_,
  chained_data_delayed_20__85_,chained_data_delayed_20__84_,chained_data_delayed_20__83_,
  chained_data_delayed_20__82_,chained_data_delayed_20__81_,
  chained_data_delayed_20__80_,chained_data_delayed_20__79_,chained_data_delayed_20__78_,
  chained_data_delayed_20__77_,chained_data_delayed_20__76_,chained_data_delayed_20__75_,
  chained_data_delayed_20__74_,chained_data_delayed_20__73_,chained_data_delayed_20__72_,
  chained_data_delayed_20__71_,chained_data_delayed_20__70_,
  chained_data_delayed_20__69_,chained_data_delayed_20__68_,chained_data_delayed_20__67_,
  chained_data_delayed_20__66_,chained_data_delayed_20__65_,chained_data_delayed_20__64_,
  chained_data_delayed_20__63_,chained_data_delayed_20__62_,chained_data_delayed_20__61_,
  chained_data_delayed_20__60_,chained_data_delayed_20__59_,chained_data_delayed_20__58_,
  chained_data_delayed_20__57_,chained_data_delayed_20__56_,
  chained_data_delayed_20__55_,chained_data_delayed_20__54_,chained_data_delayed_20__53_,
  chained_data_delayed_20__52_,chained_data_delayed_20__51_,chained_data_delayed_20__50_,
  chained_data_delayed_20__49_,chained_data_delayed_20__48_,chained_data_delayed_20__47_,
  chained_data_delayed_20__46_,chained_data_delayed_20__45_,
  chained_data_delayed_20__44_,chained_data_delayed_20__43_,chained_data_delayed_20__42_,
  chained_data_delayed_20__41_,chained_data_delayed_20__40_,chained_data_delayed_20__39_,
  chained_data_delayed_20__38_,chained_data_delayed_20__37_,chained_data_delayed_20__36_,
  chained_data_delayed_20__35_,chained_data_delayed_20__34_,
  chained_data_delayed_20__33_,chained_data_delayed_20__32_,chained_data_delayed_20__31_,
  chained_data_delayed_20__30_,chained_data_delayed_20__29_,chained_data_delayed_20__28_,
  chained_data_delayed_20__27_,chained_data_delayed_20__26_,chained_data_delayed_20__25_,
  chained_data_delayed_20__24_,chained_data_delayed_20__23_,
  chained_data_delayed_20__22_,chained_data_delayed_20__21_,chained_data_delayed_20__20_,
  chained_data_delayed_20__19_,chained_data_delayed_20__18_,chained_data_delayed_20__17_,
  chained_data_delayed_20__16_,chained_data_delayed_20__15_,chained_data_delayed_20__14_,
  chained_data_delayed_20__13_,chained_data_delayed_20__12_,
  chained_data_delayed_20__11_,chained_data_delayed_20__10_,chained_data_delayed_20__9_,
  chained_data_delayed_20__8_,chained_data_delayed_20__7_,chained_data_delayed_20__6_,
  chained_data_delayed_20__5_,chained_data_delayed_20__4_,chained_data_delayed_20__3_,
  chained_data_delayed_20__2_,chained_data_delayed_20__1_,chained_data_delayed_20__0_,
  chained_data_delayed_19__127_,chained_data_delayed_19__126_,
  chained_data_delayed_19__125_,chained_data_delayed_19__124_,chained_data_delayed_19__123_,
  chained_data_delayed_19__122_,chained_data_delayed_19__121_,chained_data_delayed_19__120_,
  chained_data_delayed_19__119_,chained_data_delayed_19__118_,
  chained_data_delayed_19__117_,chained_data_delayed_19__116_,chained_data_delayed_19__115_,
  chained_data_delayed_19__114_,chained_data_delayed_19__113_,chained_data_delayed_19__112_,
  chained_data_delayed_19__111_,chained_data_delayed_19__110_,
  chained_data_delayed_19__109_,chained_data_delayed_19__108_,chained_data_delayed_19__107_,
  chained_data_delayed_19__106_,chained_data_delayed_19__105_,chained_data_delayed_19__104_,
  chained_data_delayed_19__103_,chained_data_delayed_19__102_,
  chained_data_delayed_19__101_,chained_data_delayed_19__100_,chained_data_delayed_19__99_,
  chained_data_delayed_19__98_,chained_data_delayed_19__97_,chained_data_delayed_19__96_,
  chained_data_delayed_19__95_,chained_data_delayed_19__94_,chained_data_delayed_19__93_,
  chained_data_delayed_19__92_,chained_data_delayed_19__91_,
  chained_data_delayed_19__90_,chained_data_delayed_19__89_,chained_data_delayed_19__88_,
  chained_data_delayed_19__87_,chained_data_delayed_19__86_,chained_data_delayed_19__85_,
  chained_data_delayed_19__84_,chained_data_delayed_19__83_,chained_data_delayed_19__82_,
  chained_data_delayed_19__81_,chained_data_delayed_19__80_,
  chained_data_delayed_19__79_,chained_data_delayed_19__78_,chained_data_delayed_19__77_,
  chained_data_delayed_19__76_,chained_data_delayed_19__75_,chained_data_delayed_19__74_,
  chained_data_delayed_19__73_,chained_data_delayed_19__72_,chained_data_delayed_19__71_,
  chained_data_delayed_19__70_,chained_data_delayed_19__69_,chained_data_delayed_19__68_,
  chained_data_delayed_19__67_,chained_data_delayed_19__66_,
  chained_data_delayed_19__65_,chained_data_delayed_19__64_,chained_data_delayed_19__63_,
  chained_data_delayed_19__62_,chained_data_delayed_19__61_,chained_data_delayed_19__60_,
  chained_data_delayed_19__59_,chained_data_delayed_19__58_,chained_data_delayed_19__57_,
  chained_data_delayed_19__56_,chained_data_delayed_19__55_,
  chained_data_delayed_19__54_,chained_data_delayed_19__53_,chained_data_delayed_19__52_,
  chained_data_delayed_19__51_,chained_data_delayed_19__50_,chained_data_delayed_19__49_,
  chained_data_delayed_19__48_,chained_data_delayed_19__47_,chained_data_delayed_19__46_,
  chained_data_delayed_19__45_,chained_data_delayed_19__44_,
  chained_data_delayed_19__43_,chained_data_delayed_19__42_,chained_data_delayed_19__41_,
  chained_data_delayed_19__40_,chained_data_delayed_19__39_,chained_data_delayed_19__38_,
  chained_data_delayed_19__37_,chained_data_delayed_19__36_,chained_data_delayed_19__35_,
  chained_data_delayed_19__34_,chained_data_delayed_19__33_,
  chained_data_delayed_19__32_,chained_data_delayed_19__31_,chained_data_delayed_19__30_,
  chained_data_delayed_19__29_,chained_data_delayed_19__28_,chained_data_delayed_19__27_,
  chained_data_delayed_19__26_,chained_data_delayed_19__25_,chained_data_delayed_19__24_,
  chained_data_delayed_19__23_,chained_data_delayed_19__22_,
  chained_data_delayed_19__21_,chained_data_delayed_19__20_,chained_data_delayed_19__19_,
  chained_data_delayed_19__18_,chained_data_delayed_19__17_,chained_data_delayed_19__16_,
  chained_data_delayed_19__15_,chained_data_delayed_19__14_,chained_data_delayed_19__13_,
  chained_data_delayed_19__12_,chained_data_delayed_19__11_,
  chained_data_delayed_19__10_,chained_data_delayed_19__9_,chained_data_delayed_19__8_,
  chained_data_delayed_19__7_,chained_data_delayed_19__6_,chained_data_delayed_19__5_,
  chained_data_delayed_19__4_,chained_data_delayed_19__3_,chained_data_delayed_19__2_,
  chained_data_delayed_19__1_,chained_data_delayed_19__0_,chained_data_delayed_18__127_,
  chained_data_delayed_18__126_,chained_data_delayed_18__125_,
  chained_data_delayed_18__124_,chained_data_delayed_18__123_,chained_data_delayed_18__122_,
  chained_data_delayed_18__121_,chained_data_delayed_18__120_,chained_data_delayed_18__119_,
  chained_data_delayed_18__118_,chained_data_delayed_18__117_,
  chained_data_delayed_18__116_,chained_data_delayed_18__115_,chained_data_delayed_18__114_,
  chained_data_delayed_18__113_,chained_data_delayed_18__112_,chained_data_delayed_18__111_,
  chained_data_delayed_18__110_,chained_data_delayed_18__109_,
  chained_data_delayed_18__108_,chained_data_delayed_18__107_,chained_data_delayed_18__106_,
  chained_data_delayed_18__105_,chained_data_delayed_18__104_,chained_data_delayed_18__103_,
  chained_data_delayed_18__102_,chained_data_delayed_18__101_,
  chained_data_delayed_18__100_,chained_data_delayed_18__99_,chained_data_delayed_18__98_,
  chained_data_delayed_18__97_,chained_data_delayed_18__96_,chained_data_delayed_18__95_,
  chained_data_delayed_18__94_,chained_data_delayed_18__93_,chained_data_delayed_18__92_,
  chained_data_delayed_18__91_,chained_data_delayed_18__90_,
  chained_data_delayed_18__89_,chained_data_delayed_18__88_,chained_data_delayed_18__87_,
  chained_data_delayed_18__86_,chained_data_delayed_18__85_,chained_data_delayed_18__84_,
  chained_data_delayed_18__83_,chained_data_delayed_18__82_,chained_data_delayed_18__81_,
  chained_data_delayed_18__80_,chained_data_delayed_18__79_,chained_data_delayed_18__78_,
  chained_data_delayed_18__77_,chained_data_delayed_18__76_,
  chained_data_delayed_18__75_,chained_data_delayed_18__74_,chained_data_delayed_18__73_,
  chained_data_delayed_18__72_,chained_data_delayed_18__71_,chained_data_delayed_18__70_,
  chained_data_delayed_18__69_,chained_data_delayed_18__68_,chained_data_delayed_18__67_,
  chained_data_delayed_18__66_,chained_data_delayed_18__65_,
  chained_data_delayed_18__64_,chained_data_delayed_18__63_,chained_data_delayed_18__62_,
  chained_data_delayed_18__61_,chained_data_delayed_18__60_,chained_data_delayed_18__59_,
  chained_data_delayed_18__58_,chained_data_delayed_18__57_,chained_data_delayed_18__56_,
  chained_data_delayed_18__55_,chained_data_delayed_18__54_,
  chained_data_delayed_18__53_,chained_data_delayed_18__52_,chained_data_delayed_18__51_,
  chained_data_delayed_18__50_,chained_data_delayed_18__49_,chained_data_delayed_18__48_,
  chained_data_delayed_18__47_,chained_data_delayed_18__46_,chained_data_delayed_18__45_,
  chained_data_delayed_18__44_,chained_data_delayed_18__43_,
  chained_data_delayed_18__42_,chained_data_delayed_18__41_,chained_data_delayed_18__40_,
  chained_data_delayed_18__39_,chained_data_delayed_18__38_,chained_data_delayed_18__37_,
  chained_data_delayed_18__36_,chained_data_delayed_18__35_,chained_data_delayed_18__34_,
  chained_data_delayed_18__33_,chained_data_delayed_18__32_,
  chained_data_delayed_18__31_,chained_data_delayed_18__30_,chained_data_delayed_18__29_,
  chained_data_delayed_18__28_,chained_data_delayed_18__27_,chained_data_delayed_18__26_,
  chained_data_delayed_18__25_,chained_data_delayed_18__24_,chained_data_delayed_18__23_,
  chained_data_delayed_18__22_,chained_data_delayed_18__21_,
  chained_data_delayed_18__20_,chained_data_delayed_18__19_,chained_data_delayed_18__18_,
  chained_data_delayed_18__17_,chained_data_delayed_18__16_,chained_data_delayed_18__15_,
  chained_data_delayed_18__14_,chained_data_delayed_18__13_,chained_data_delayed_18__12_,
  chained_data_delayed_18__11_,chained_data_delayed_18__10_,chained_data_delayed_18__9_,
  chained_data_delayed_18__8_,chained_data_delayed_18__7_,
  chained_data_delayed_18__6_,chained_data_delayed_18__5_,chained_data_delayed_18__4_,
  chained_data_delayed_18__3_,chained_data_delayed_18__2_,chained_data_delayed_18__1_,
  chained_data_delayed_18__0_,chained_data_delayed_17__127_,chained_data_delayed_17__126_,
  chained_data_delayed_17__125_,chained_data_delayed_17__124_,
  chained_data_delayed_17__123_,chained_data_delayed_17__122_,chained_data_delayed_17__121_,
  chained_data_delayed_17__120_,chained_data_delayed_17__119_,chained_data_delayed_17__118_,
  chained_data_delayed_17__117_,chained_data_delayed_17__116_,
  chained_data_delayed_17__115_,chained_data_delayed_17__114_,chained_data_delayed_17__113_,
  chained_data_delayed_17__112_,chained_data_delayed_17__111_,chained_data_delayed_17__110_,
  chained_data_delayed_17__109_,chained_data_delayed_17__108_,
  chained_data_delayed_17__107_,chained_data_delayed_17__106_,chained_data_delayed_17__105_,
  chained_data_delayed_17__104_,chained_data_delayed_17__103_,chained_data_delayed_17__102_,
  chained_data_delayed_17__101_,chained_data_delayed_17__100_,
  chained_data_delayed_17__99_,chained_data_delayed_17__98_,chained_data_delayed_17__97_,
  chained_data_delayed_17__96_,chained_data_delayed_17__95_,chained_data_delayed_17__94_,
  chained_data_delayed_17__93_,chained_data_delayed_17__92_,chained_data_delayed_17__91_,
  chained_data_delayed_17__90_,chained_data_delayed_17__89_,chained_data_delayed_17__88_,
  chained_data_delayed_17__87_,chained_data_delayed_17__86_,
  chained_data_delayed_17__85_,chained_data_delayed_17__84_,chained_data_delayed_17__83_,
  chained_data_delayed_17__82_,chained_data_delayed_17__81_,chained_data_delayed_17__80_,
  chained_data_delayed_17__79_,chained_data_delayed_17__78_,chained_data_delayed_17__77_,
  chained_data_delayed_17__76_,chained_data_delayed_17__75_,
  chained_data_delayed_17__74_,chained_data_delayed_17__73_,chained_data_delayed_17__72_,
  chained_data_delayed_17__71_,chained_data_delayed_17__70_,chained_data_delayed_17__69_,
  chained_data_delayed_17__68_,chained_data_delayed_17__67_,chained_data_delayed_17__66_,
  chained_data_delayed_17__65_,chained_data_delayed_17__64_,
  chained_data_delayed_17__63_,chained_data_delayed_17__62_,chained_data_delayed_17__61_,
  chained_data_delayed_17__60_,chained_data_delayed_17__59_,chained_data_delayed_17__58_,
  chained_data_delayed_17__57_,chained_data_delayed_17__56_,chained_data_delayed_17__55_,
  chained_data_delayed_17__54_,chained_data_delayed_17__53_,
  chained_data_delayed_17__52_,chained_data_delayed_17__51_,chained_data_delayed_17__50_,
  chained_data_delayed_17__49_,chained_data_delayed_17__48_,chained_data_delayed_17__47_,
  chained_data_delayed_17__46_,chained_data_delayed_17__45_,chained_data_delayed_17__44_,
  chained_data_delayed_17__43_,chained_data_delayed_17__42_,
  chained_data_delayed_17__41_,chained_data_delayed_17__40_,chained_data_delayed_17__39_,
  chained_data_delayed_17__38_,chained_data_delayed_17__37_,chained_data_delayed_17__36_,
  chained_data_delayed_17__35_,chained_data_delayed_17__34_,chained_data_delayed_17__33_,
  chained_data_delayed_17__32_,chained_data_delayed_17__31_,
  chained_data_delayed_17__30_,chained_data_delayed_17__29_,chained_data_delayed_17__28_,
  chained_data_delayed_17__27_,chained_data_delayed_17__26_,chained_data_delayed_17__25_,
  chained_data_delayed_17__24_,chained_data_delayed_17__23_,chained_data_delayed_17__22_,
  chained_data_delayed_17__21_,chained_data_delayed_17__20_,
  chained_data_delayed_17__19_,chained_data_delayed_17__18_,chained_data_delayed_17__17_,
  chained_data_delayed_17__16_,chained_data_delayed_17__15_,chained_data_delayed_17__14_,
  chained_data_delayed_17__13_,chained_data_delayed_17__12_,chained_data_delayed_17__11_,
  chained_data_delayed_17__10_,chained_data_delayed_17__9_,chained_data_delayed_17__8_,
  chained_data_delayed_17__7_,chained_data_delayed_17__6_,
  chained_data_delayed_17__5_,chained_data_delayed_17__4_,chained_data_delayed_17__3_,
  chained_data_delayed_17__2_,chained_data_delayed_17__1_,chained_data_delayed_17__0_,
  chained_data_delayed_24__127_,chained_data_delayed_24__126_,chained_data_delayed_24__125_,
  chained_data_delayed_24__124_,chained_data_delayed_24__123_,
  chained_data_delayed_24__122_,chained_data_delayed_24__121_,chained_data_delayed_24__120_,
  chained_data_delayed_24__119_,chained_data_delayed_24__118_,chained_data_delayed_24__117_,
  chained_data_delayed_24__116_,chained_data_delayed_24__115_,
  chained_data_delayed_24__114_,chained_data_delayed_24__113_,chained_data_delayed_24__112_,
  chained_data_delayed_24__111_,chained_data_delayed_24__110_,chained_data_delayed_24__109_,
  chained_data_delayed_24__108_,chained_data_delayed_24__107_,
  chained_data_delayed_24__106_,chained_data_delayed_24__105_,chained_data_delayed_24__104_,
  chained_data_delayed_24__103_,chained_data_delayed_24__102_,chained_data_delayed_24__101_,
  chained_data_delayed_24__100_,chained_data_delayed_24__99_,chained_data_delayed_24__98_,
  chained_data_delayed_24__97_,chained_data_delayed_24__96_,
  chained_data_delayed_24__95_,chained_data_delayed_24__94_,chained_data_delayed_24__93_,
  chained_data_delayed_24__92_,chained_data_delayed_24__91_,chained_data_delayed_24__90_,
  chained_data_delayed_24__89_,chained_data_delayed_24__88_,chained_data_delayed_24__87_,
  chained_data_delayed_24__86_,chained_data_delayed_24__85_,
  chained_data_delayed_24__84_,chained_data_delayed_24__83_,chained_data_delayed_24__82_,
  chained_data_delayed_24__81_,chained_data_delayed_24__80_,chained_data_delayed_24__79_,
  chained_data_delayed_24__78_,chained_data_delayed_24__77_,chained_data_delayed_24__76_,
  chained_data_delayed_24__75_,chained_data_delayed_24__74_,
  chained_data_delayed_24__73_,chained_data_delayed_24__72_,chained_data_delayed_24__71_,
  chained_data_delayed_24__70_,chained_data_delayed_24__69_,chained_data_delayed_24__68_,
  chained_data_delayed_24__67_,chained_data_delayed_24__66_,chained_data_delayed_24__65_,
  chained_data_delayed_24__64_,chained_data_delayed_24__63_,
  chained_data_delayed_24__62_,chained_data_delayed_24__61_,chained_data_delayed_24__60_,
  chained_data_delayed_24__59_,chained_data_delayed_24__58_,chained_data_delayed_24__57_,
  chained_data_delayed_24__56_,chained_data_delayed_24__55_,chained_data_delayed_24__54_,
  chained_data_delayed_24__53_,chained_data_delayed_24__52_,
  chained_data_delayed_24__51_,chained_data_delayed_24__50_,chained_data_delayed_24__49_,
  chained_data_delayed_24__48_,chained_data_delayed_24__47_,chained_data_delayed_24__46_,
  chained_data_delayed_24__45_,chained_data_delayed_24__44_,chained_data_delayed_24__43_,
  chained_data_delayed_24__42_,chained_data_delayed_24__41_,
  chained_data_delayed_24__40_,chained_data_delayed_24__39_,chained_data_delayed_24__38_,
  chained_data_delayed_24__37_,chained_data_delayed_24__36_,chained_data_delayed_24__35_,
  chained_data_delayed_24__34_,chained_data_delayed_24__33_,chained_data_delayed_24__32_,
  chained_data_delayed_24__31_,chained_data_delayed_24__30_,
  chained_data_delayed_24__29_,chained_data_delayed_24__28_,chained_data_delayed_24__27_,
  chained_data_delayed_24__26_,chained_data_delayed_24__25_,chained_data_delayed_24__24_,
  chained_data_delayed_24__23_,chained_data_delayed_24__22_,chained_data_delayed_24__21_,
  chained_data_delayed_24__20_,chained_data_delayed_24__19_,chained_data_delayed_24__18_,
  chained_data_delayed_24__17_,chained_data_delayed_24__16_,
  chained_data_delayed_24__15_,chained_data_delayed_24__14_,chained_data_delayed_24__13_,
  chained_data_delayed_24__12_,chained_data_delayed_24__11_,chained_data_delayed_24__10_,
  chained_data_delayed_24__9_,chained_data_delayed_24__8_,chained_data_delayed_24__7_,
  chained_data_delayed_24__6_,chained_data_delayed_24__5_,chained_data_delayed_24__4_,
  chained_data_delayed_24__3_,chained_data_delayed_24__2_,
  chained_data_delayed_24__1_,chained_data_delayed_24__0_,chained_data_delayed_23__127_,
  chained_data_delayed_23__126_,chained_data_delayed_23__125_,chained_data_delayed_23__124_,
  chained_data_delayed_23__123_,chained_data_delayed_23__122_,
  chained_data_delayed_23__121_,chained_data_delayed_23__120_,chained_data_delayed_23__119_,
  chained_data_delayed_23__118_,chained_data_delayed_23__117_,chained_data_delayed_23__116_,
  chained_data_delayed_23__115_,chained_data_delayed_23__114_,
  chained_data_delayed_23__113_,chained_data_delayed_23__112_,chained_data_delayed_23__111_,
  chained_data_delayed_23__110_,chained_data_delayed_23__109_,chained_data_delayed_23__108_,
  chained_data_delayed_23__107_,chained_data_delayed_23__106_,
  chained_data_delayed_23__105_,chained_data_delayed_23__104_,chained_data_delayed_23__103_,
  chained_data_delayed_23__102_,chained_data_delayed_23__101_,chained_data_delayed_23__100_,
  chained_data_delayed_23__99_,chained_data_delayed_23__98_,chained_data_delayed_23__97_,
  chained_data_delayed_23__96_,chained_data_delayed_23__95_,
  chained_data_delayed_23__94_,chained_data_delayed_23__93_,chained_data_delayed_23__92_,
  chained_data_delayed_23__91_,chained_data_delayed_23__90_,chained_data_delayed_23__89_,
  chained_data_delayed_23__88_,chained_data_delayed_23__87_,chained_data_delayed_23__86_,
  chained_data_delayed_23__85_,chained_data_delayed_23__84_,
  chained_data_delayed_23__83_,chained_data_delayed_23__82_,chained_data_delayed_23__81_,
  chained_data_delayed_23__80_,chained_data_delayed_23__79_,chained_data_delayed_23__78_,
  chained_data_delayed_23__77_,chained_data_delayed_23__76_,chained_data_delayed_23__75_,
  chained_data_delayed_23__74_,chained_data_delayed_23__73_,
  chained_data_delayed_23__72_,chained_data_delayed_23__71_,chained_data_delayed_23__70_,
  chained_data_delayed_23__69_,chained_data_delayed_23__68_,chained_data_delayed_23__67_,
  chained_data_delayed_23__66_,chained_data_delayed_23__65_,chained_data_delayed_23__64_,
  chained_data_delayed_23__63_,chained_data_delayed_23__62_,
  chained_data_delayed_23__61_,chained_data_delayed_23__60_,chained_data_delayed_23__59_,
  chained_data_delayed_23__58_,chained_data_delayed_23__57_,chained_data_delayed_23__56_,
  chained_data_delayed_23__55_,chained_data_delayed_23__54_,chained_data_delayed_23__53_,
  chained_data_delayed_23__52_,chained_data_delayed_23__51_,
  chained_data_delayed_23__50_,chained_data_delayed_23__49_,chained_data_delayed_23__48_,
  chained_data_delayed_23__47_,chained_data_delayed_23__46_,chained_data_delayed_23__45_,
  chained_data_delayed_23__44_,chained_data_delayed_23__43_,chained_data_delayed_23__42_,
  chained_data_delayed_23__41_,chained_data_delayed_23__40_,
  chained_data_delayed_23__39_,chained_data_delayed_23__38_,chained_data_delayed_23__37_,
  chained_data_delayed_23__36_,chained_data_delayed_23__35_,chained_data_delayed_23__34_,
  chained_data_delayed_23__33_,chained_data_delayed_23__32_,chained_data_delayed_23__31_,
  chained_data_delayed_23__30_,chained_data_delayed_23__29_,chained_data_delayed_23__28_,
  chained_data_delayed_23__27_,chained_data_delayed_23__26_,
  chained_data_delayed_23__25_,chained_data_delayed_23__24_,chained_data_delayed_23__23_,
  chained_data_delayed_23__22_,chained_data_delayed_23__21_,chained_data_delayed_23__20_,
  chained_data_delayed_23__19_,chained_data_delayed_23__18_,chained_data_delayed_23__17_,
  chained_data_delayed_23__16_,chained_data_delayed_23__15_,
  chained_data_delayed_23__14_,chained_data_delayed_23__13_,chained_data_delayed_23__12_,
  chained_data_delayed_23__11_,chained_data_delayed_23__10_,chained_data_delayed_23__9_,
  chained_data_delayed_23__8_,chained_data_delayed_23__7_,chained_data_delayed_23__6_,
  chained_data_delayed_23__5_,chained_data_delayed_23__4_,chained_data_delayed_23__3_,
  chained_data_delayed_23__2_,chained_data_delayed_23__1_,
  chained_data_delayed_23__0_,chained_data_delayed_22__127_,chained_data_delayed_22__126_,
  chained_data_delayed_22__125_,chained_data_delayed_22__124_,chained_data_delayed_22__123_,
  chained_data_delayed_22__122_,chained_data_delayed_22__121_,
  chained_data_delayed_22__120_,chained_data_delayed_22__119_,chained_data_delayed_22__118_,
  chained_data_delayed_22__117_,chained_data_delayed_22__116_,chained_data_delayed_22__115_,
  chained_data_delayed_22__114_,chained_data_delayed_22__113_,
  chained_data_delayed_22__112_,chained_data_delayed_22__111_,chained_data_delayed_22__110_,
  chained_data_delayed_22__109_,chained_data_delayed_22__108_,chained_data_delayed_22__107_,
  chained_data_delayed_22__106_,chained_data_delayed_22__105_,
  chained_data_delayed_22__104_,chained_data_delayed_22__103_,chained_data_delayed_22__102_,
  chained_data_delayed_22__101_,chained_data_delayed_22__100_,chained_data_delayed_22__99_,
  chained_data_delayed_22__98_,chained_data_delayed_22__97_,chained_data_delayed_22__96_,
  chained_data_delayed_22__95_,chained_data_delayed_22__94_,
  chained_data_delayed_22__93_,chained_data_delayed_22__92_,chained_data_delayed_22__91_,
  chained_data_delayed_22__90_,chained_data_delayed_22__89_,chained_data_delayed_22__88_,
  chained_data_delayed_22__87_,chained_data_delayed_22__86_,chained_data_delayed_22__85_,
  chained_data_delayed_22__84_,chained_data_delayed_22__83_,
  chained_data_delayed_22__82_,chained_data_delayed_22__81_,chained_data_delayed_22__80_,
  chained_data_delayed_22__79_,chained_data_delayed_22__78_,chained_data_delayed_22__77_,
  chained_data_delayed_22__76_,chained_data_delayed_22__75_,chained_data_delayed_22__74_,
  chained_data_delayed_22__73_,chained_data_delayed_22__72_,
  chained_data_delayed_22__71_,chained_data_delayed_22__70_,chained_data_delayed_22__69_,
  chained_data_delayed_22__68_,chained_data_delayed_22__67_,chained_data_delayed_22__66_,
  chained_data_delayed_22__65_,chained_data_delayed_22__64_,chained_data_delayed_22__63_,
  chained_data_delayed_22__62_,chained_data_delayed_22__61_,
  chained_data_delayed_22__60_,chained_data_delayed_22__59_,chained_data_delayed_22__58_,
  chained_data_delayed_22__57_,chained_data_delayed_22__56_,chained_data_delayed_22__55_,
  chained_data_delayed_22__54_,chained_data_delayed_22__53_,chained_data_delayed_22__52_,
  chained_data_delayed_22__51_,chained_data_delayed_22__50_,
  chained_data_delayed_22__49_,chained_data_delayed_22__48_,chained_data_delayed_22__47_,
  chained_data_delayed_22__46_,chained_data_delayed_22__45_,chained_data_delayed_22__44_,
  chained_data_delayed_22__43_,chained_data_delayed_22__42_,chained_data_delayed_22__41_,
  chained_data_delayed_22__40_,chained_data_delayed_22__39_,chained_data_delayed_22__38_,
  chained_data_delayed_22__37_,chained_data_delayed_22__36_,
  chained_data_delayed_22__35_,chained_data_delayed_22__34_,chained_data_delayed_22__33_,
  chained_data_delayed_22__32_,chained_data_delayed_22__31_,chained_data_delayed_22__30_,
  chained_data_delayed_22__29_,chained_data_delayed_22__28_,chained_data_delayed_22__27_,
  chained_data_delayed_22__26_,chained_data_delayed_22__25_,
  chained_data_delayed_22__24_,chained_data_delayed_22__23_,chained_data_delayed_22__22_,
  chained_data_delayed_22__21_,chained_data_delayed_22__20_,chained_data_delayed_22__19_,
  chained_data_delayed_22__18_,chained_data_delayed_22__17_,chained_data_delayed_22__16_,
  chained_data_delayed_22__15_,chained_data_delayed_22__14_,
  chained_data_delayed_22__13_,chained_data_delayed_22__12_,chained_data_delayed_22__11_,
  chained_data_delayed_22__10_,chained_data_delayed_22__9_,chained_data_delayed_22__8_,
  chained_data_delayed_22__7_,chained_data_delayed_22__6_,chained_data_delayed_22__5_,
  chained_data_delayed_22__4_,chained_data_delayed_22__3_,chained_data_delayed_22__2_,
  chained_data_delayed_22__1_,chained_data_delayed_22__0_,
  chained_data_delayed_21__127_,chained_data_delayed_21__126_,chained_data_delayed_21__125_,
  chained_data_delayed_21__124_,chained_data_delayed_21__123_,chained_data_delayed_21__122_,
  chained_data_delayed_21__121_,chained_data_delayed_21__120_,
  chained_data_delayed_21__119_,chained_data_delayed_21__118_,chained_data_delayed_21__117_,
  chained_data_delayed_21__116_,chained_data_delayed_21__115_,chained_data_delayed_21__114_,
  chained_data_delayed_21__113_,chained_data_delayed_21__112_,
  chained_data_delayed_21__111_,chained_data_delayed_21__110_,chained_data_delayed_21__109_,
  chained_data_delayed_21__108_,chained_data_delayed_21__107_,chained_data_delayed_21__106_,
  chained_data_delayed_21__105_,chained_data_delayed_21__104_,
  chained_data_delayed_21__103_,chained_data_delayed_21__102_,chained_data_delayed_21__101_,
  chained_data_delayed_21__100_,chained_data_delayed_21__99_,chained_data_delayed_21__98_,
  chained_data_delayed_21__97_,chained_data_delayed_21__96_,chained_data_delayed_21__95_,
  chained_data_delayed_21__94_,chained_data_delayed_21__93_,
  chained_data_delayed_21__92_,chained_data_delayed_21__91_,chained_data_delayed_21__90_,
  chained_data_delayed_21__89_,chained_data_delayed_21__88_,chained_data_delayed_21__87_,
  chained_data_delayed_21__86_,chained_data_delayed_21__85_,chained_data_delayed_21__84_,
  chained_data_delayed_21__83_,chained_data_delayed_21__82_,
  chained_data_delayed_21__81_,chained_data_delayed_21__80_,chained_data_delayed_21__79_,
  chained_data_delayed_21__78_,chained_data_delayed_21__77_,chained_data_delayed_21__76_,
  chained_data_delayed_21__75_,chained_data_delayed_21__74_,chained_data_delayed_21__73_,
  chained_data_delayed_21__72_,chained_data_delayed_21__71_,
  chained_data_delayed_21__70_,chained_data_delayed_21__69_,chained_data_delayed_21__68_,
  chained_data_delayed_21__67_,chained_data_delayed_21__66_,chained_data_delayed_21__65_,
  chained_data_delayed_21__64_,chained_data_delayed_21__63_,chained_data_delayed_21__62_,
  chained_data_delayed_21__61_,chained_data_delayed_21__60_,
  chained_data_delayed_21__59_,chained_data_delayed_21__58_,chained_data_delayed_21__57_,
  chained_data_delayed_21__56_,chained_data_delayed_21__55_,chained_data_delayed_21__54_,
  chained_data_delayed_21__53_,chained_data_delayed_21__52_,chained_data_delayed_21__51_,
  chained_data_delayed_21__50_,chained_data_delayed_21__49_,chained_data_delayed_21__48_,
  chained_data_delayed_21__47_,chained_data_delayed_21__46_,
  chained_data_delayed_21__45_,chained_data_delayed_21__44_,chained_data_delayed_21__43_,
  chained_data_delayed_21__42_,chained_data_delayed_21__41_,chained_data_delayed_21__40_,
  chained_data_delayed_21__39_,chained_data_delayed_21__38_,chained_data_delayed_21__37_,
  chained_data_delayed_21__36_,chained_data_delayed_21__35_,
  chained_data_delayed_21__34_,chained_data_delayed_21__33_,chained_data_delayed_21__32_,
  chained_data_delayed_21__31_,chained_data_delayed_21__30_,chained_data_delayed_21__29_,
  chained_data_delayed_21__28_,chained_data_delayed_21__27_,chained_data_delayed_21__26_,
  chained_data_delayed_21__25_,chained_data_delayed_21__24_,
  chained_data_delayed_21__23_,chained_data_delayed_21__22_,chained_data_delayed_21__21_,
  chained_data_delayed_21__20_,chained_data_delayed_21__19_,chained_data_delayed_21__18_,
  chained_data_delayed_21__17_,chained_data_delayed_21__16_,chained_data_delayed_21__15_,
  chained_data_delayed_21__14_,chained_data_delayed_21__13_,
  chained_data_delayed_21__12_,chained_data_delayed_21__11_,chained_data_delayed_21__10_,
  chained_data_delayed_21__9_,chained_data_delayed_21__8_,chained_data_delayed_21__7_,
  chained_data_delayed_21__6_,chained_data_delayed_21__5_,chained_data_delayed_21__4_,
  chained_data_delayed_21__3_,chained_data_delayed_21__2_,chained_data_delayed_21__1_,
  chained_data_delayed_21__0_,chained_data_delayed_28__127_,
  chained_data_delayed_28__126_,chained_data_delayed_28__125_,chained_data_delayed_28__124_,
  chained_data_delayed_28__123_,chained_data_delayed_28__122_,chained_data_delayed_28__121_,
  chained_data_delayed_28__120_,chained_data_delayed_28__119_,
  chained_data_delayed_28__118_,chained_data_delayed_28__117_,chained_data_delayed_28__116_,
  chained_data_delayed_28__115_,chained_data_delayed_28__114_,chained_data_delayed_28__113_,
  chained_data_delayed_28__112_,chained_data_delayed_28__111_,
  chained_data_delayed_28__110_,chained_data_delayed_28__109_,chained_data_delayed_28__108_,
  chained_data_delayed_28__107_,chained_data_delayed_28__106_,chained_data_delayed_28__105_,
  chained_data_delayed_28__104_,chained_data_delayed_28__103_,
  chained_data_delayed_28__102_,chained_data_delayed_28__101_,chained_data_delayed_28__100_,
  chained_data_delayed_28__99_,chained_data_delayed_28__98_,chained_data_delayed_28__97_,
  chained_data_delayed_28__96_,chained_data_delayed_28__95_,chained_data_delayed_28__94_,
  chained_data_delayed_28__93_,chained_data_delayed_28__92_,
  chained_data_delayed_28__91_,chained_data_delayed_28__90_,chained_data_delayed_28__89_,
  chained_data_delayed_28__88_,chained_data_delayed_28__87_,chained_data_delayed_28__86_,
  chained_data_delayed_28__85_,chained_data_delayed_28__84_,chained_data_delayed_28__83_,
  chained_data_delayed_28__82_,chained_data_delayed_28__81_,
  chained_data_delayed_28__80_,chained_data_delayed_28__79_,chained_data_delayed_28__78_,
  chained_data_delayed_28__77_,chained_data_delayed_28__76_,chained_data_delayed_28__75_,
  chained_data_delayed_28__74_,chained_data_delayed_28__73_,chained_data_delayed_28__72_,
  chained_data_delayed_28__71_,chained_data_delayed_28__70_,
  chained_data_delayed_28__69_,chained_data_delayed_28__68_,chained_data_delayed_28__67_,
  chained_data_delayed_28__66_,chained_data_delayed_28__65_,chained_data_delayed_28__64_,
  chained_data_delayed_28__63_,chained_data_delayed_28__62_,chained_data_delayed_28__61_,
  chained_data_delayed_28__60_,chained_data_delayed_28__59_,chained_data_delayed_28__58_,
  chained_data_delayed_28__57_,chained_data_delayed_28__56_,
  chained_data_delayed_28__55_,chained_data_delayed_28__54_,chained_data_delayed_28__53_,
  chained_data_delayed_28__52_,chained_data_delayed_28__51_,chained_data_delayed_28__50_,
  chained_data_delayed_28__49_,chained_data_delayed_28__48_,chained_data_delayed_28__47_,
  chained_data_delayed_28__46_,chained_data_delayed_28__45_,
  chained_data_delayed_28__44_,chained_data_delayed_28__43_,chained_data_delayed_28__42_,
  chained_data_delayed_28__41_,chained_data_delayed_28__40_,chained_data_delayed_28__39_,
  chained_data_delayed_28__38_,chained_data_delayed_28__37_,chained_data_delayed_28__36_,
  chained_data_delayed_28__35_,chained_data_delayed_28__34_,
  chained_data_delayed_28__33_,chained_data_delayed_28__32_,chained_data_delayed_28__31_,
  chained_data_delayed_28__30_,chained_data_delayed_28__29_,chained_data_delayed_28__28_,
  chained_data_delayed_28__27_,chained_data_delayed_28__26_,chained_data_delayed_28__25_,
  chained_data_delayed_28__24_,chained_data_delayed_28__23_,
  chained_data_delayed_28__22_,chained_data_delayed_28__21_,chained_data_delayed_28__20_,
  chained_data_delayed_28__19_,chained_data_delayed_28__18_,chained_data_delayed_28__17_,
  chained_data_delayed_28__16_,chained_data_delayed_28__15_,chained_data_delayed_28__14_,
  chained_data_delayed_28__13_,chained_data_delayed_28__12_,
  chained_data_delayed_28__11_,chained_data_delayed_28__10_,chained_data_delayed_28__9_,
  chained_data_delayed_28__8_,chained_data_delayed_28__7_,chained_data_delayed_28__6_,
  chained_data_delayed_28__5_,chained_data_delayed_28__4_,chained_data_delayed_28__3_,
  chained_data_delayed_28__2_,chained_data_delayed_28__1_,chained_data_delayed_28__0_,
  chained_data_delayed_27__127_,chained_data_delayed_27__126_,
  chained_data_delayed_27__125_,chained_data_delayed_27__124_,chained_data_delayed_27__123_,
  chained_data_delayed_27__122_,chained_data_delayed_27__121_,chained_data_delayed_27__120_,
  chained_data_delayed_27__119_,chained_data_delayed_27__118_,
  chained_data_delayed_27__117_,chained_data_delayed_27__116_,chained_data_delayed_27__115_,
  chained_data_delayed_27__114_,chained_data_delayed_27__113_,chained_data_delayed_27__112_,
  chained_data_delayed_27__111_,chained_data_delayed_27__110_,
  chained_data_delayed_27__109_,chained_data_delayed_27__108_,chained_data_delayed_27__107_,
  chained_data_delayed_27__106_,chained_data_delayed_27__105_,chained_data_delayed_27__104_,
  chained_data_delayed_27__103_,chained_data_delayed_27__102_,
  chained_data_delayed_27__101_,chained_data_delayed_27__100_,chained_data_delayed_27__99_,
  chained_data_delayed_27__98_,chained_data_delayed_27__97_,chained_data_delayed_27__96_,
  chained_data_delayed_27__95_,chained_data_delayed_27__94_,chained_data_delayed_27__93_,
  chained_data_delayed_27__92_,chained_data_delayed_27__91_,
  chained_data_delayed_27__90_,chained_data_delayed_27__89_,chained_data_delayed_27__88_,
  chained_data_delayed_27__87_,chained_data_delayed_27__86_,chained_data_delayed_27__85_,
  chained_data_delayed_27__84_,chained_data_delayed_27__83_,chained_data_delayed_27__82_,
  chained_data_delayed_27__81_,chained_data_delayed_27__80_,
  chained_data_delayed_27__79_,chained_data_delayed_27__78_,chained_data_delayed_27__77_,
  chained_data_delayed_27__76_,chained_data_delayed_27__75_,chained_data_delayed_27__74_,
  chained_data_delayed_27__73_,chained_data_delayed_27__72_,chained_data_delayed_27__71_,
  chained_data_delayed_27__70_,chained_data_delayed_27__69_,chained_data_delayed_27__68_,
  chained_data_delayed_27__67_,chained_data_delayed_27__66_,
  chained_data_delayed_27__65_,chained_data_delayed_27__64_,chained_data_delayed_27__63_,
  chained_data_delayed_27__62_,chained_data_delayed_27__61_,chained_data_delayed_27__60_,
  chained_data_delayed_27__59_,chained_data_delayed_27__58_,chained_data_delayed_27__57_,
  chained_data_delayed_27__56_,chained_data_delayed_27__55_,
  chained_data_delayed_27__54_,chained_data_delayed_27__53_,chained_data_delayed_27__52_,
  chained_data_delayed_27__51_,chained_data_delayed_27__50_,chained_data_delayed_27__49_,
  chained_data_delayed_27__48_,chained_data_delayed_27__47_,chained_data_delayed_27__46_,
  chained_data_delayed_27__45_,chained_data_delayed_27__44_,
  chained_data_delayed_27__43_,chained_data_delayed_27__42_,chained_data_delayed_27__41_,
  chained_data_delayed_27__40_,chained_data_delayed_27__39_,chained_data_delayed_27__38_,
  chained_data_delayed_27__37_,chained_data_delayed_27__36_,chained_data_delayed_27__35_,
  chained_data_delayed_27__34_,chained_data_delayed_27__33_,
  chained_data_delayed_27__32_,chained_data_delayed_27__31_,chained_data_delayed_27__30_,
  chained_data_delayed_27__29_,chained_data_delayed_27__28_,chained_data_delayed_27__27_,
  chained_data_delayed_27__26_,chained_data_delayed_27__25_,chained_data_delayed_27__24_,
  chained_data_delayed_27__23_,chained_data_delayed_27__22_,
  chained_data_delayed_27__21_,chained_data_delayed_27__20_,chained_data_delayed_27__19_,
  chained_data_delayed_27__18_,chained_data_delayed_27__17_,chained_data_delayed_27__16_,
  chained_data_delayed_27__15_,chained_data_delayed_27__14_,chained_data_delayed_27__13_,
  chained_data_delayed_27__12_,chained_data_delayed_27__11_,
  chained_data_delayed_27__10_,chained_data_delayed_27__9_,chained_data_delayed_27__8_,
  chained_data_delayed_27__7_,chained_data_delayed_27__6_,chained_data_delayed_27__5_,
  chained_data_delayed_27__4_,chained_data_delayed_27__3_,chained_data_delayed_27__2_,
  chained_data_delayed_27__1_,chained_data_delayed_27__0_,chained_data_delayed_26__127_,
  chained_data_delayed_26__126_,chained_data_delayed_26__125_,
  chained_data_delayed_26__124_,chained_data_delayed_26__123_,chained_data_delayed_26__122_,
  chained_data_delayed_26__121_,chained_data_delayed_26__120_,chained_data_delayed_26__119_,
  chained_data_delayed_26__118_,chained_data_delayed_26__117_,
  chained_data_delayed_26__116_,chained_data_delayed_26__115_,chained_data_delayed_26__114_,
  chained_data_delayed_26__113_,chained_data_delayed_26__112_,chained_data_delayed_26__111_,
  chained_data_delayed_26__110_,chained_data_delayed_26__109_,
  chained_data_delayed_26__108_,chained_data_delayed_26__107_,chained_data_delayed_26__106_,
  chained_data_delayed_26__105_,chained_data_delayed_26__104_,chained_data_delayed_26__103_,
  chained_data_delayed_26__102_,chained_data_delayed_26__101_,
  chained_data_delayed_26__100_,chained_data_delayed_26__99_,chained_data_delayed_26__98_,
  chained_data_delayed_26__97_,chained_data_delayed_26__96_,chained_data_delayed_26__95_,
  chained_data_delayed_26__94_,chained_data_delayed_26__93_,chained_data_delayed_26__92_,
  chained_data_delayed_26__91_,chained_data_delayed_26__90_,
  chained_data_delayed_26__89_,chained_data_delayed_26__88_,chained_data_delayed_26__87_,
  chained_data_delayed_26__86_,chained_data_delayed_26__85_,chained_data_delayed_26__84_,
  chained_data_delayed_26__83_,chained_data_delayed_26__82_,chained_data_delayed_26__81_,
  chained_data_delayed_26__80_,chained_data_delayed_26__79_,chained_data_delayed_26__78_,
  chained_data_delayed_26__77_,chained_data_delayed_26__76_,
  chained_data_delayed_26__75_,chained_data_delayed_26__74_,chained_data_delayed_26__73_,
  chained_data_delayed_26__72_,chained_data_delayed_26__71_,chained_data_delayed_26__70_,
  chained_data_delayed_26__69_,chained_data_delayed_26__68_,chained_data_delayed_26__67_,
  chained_data_delayed_26__66_,chained_data_delayed_26__65_,
  chained_data_delayed_26__64_,chained_data_delayed_26__63_,chained_data_delayed_26__62_,
  chained_data_delayed_26__61_,chained_data_delayed_26__60_,chained_data_delayed_26__59_,
  chained_data_delayed_26__58_,chained_data_delayed_26__57_,chained_data_delayed_26__56_,
  chained_data_delayed_26__55_,chained_data_delayed_26__54_,
  chained_data_delayed_26__53_,chained_data_delayed_26__52_,chained_data_delayed_26__51_,
  chained_data_delayed_26__50_,chained_data_delayed_26__49_,chained_data_delayed_26__48_,
  chained_data_delayed_26__47_,chained_data_delayed_26__46_,chained_data_delayed_26__45_,
  chained_data_delayed_26__44_,chained_data_delayed_26__43_,
  chained_data_delayed_26__42_,chained_data_delayed_26__41_,chained_data_delayed_26__40_,
  chained_data_delayed_26__39_,chained_data_delayed_26__38_,chained_data_delayed_26__37_,
  chained_data_delayed_26__36_,chained_data_delayed_26__35_,chained_data_delayed_26__34_,
  chained_data_delayed_26__33_,chained_data_delayed_26__32_,
  chained_data_delayed_26__31_,chained_data_delayed_26__30_,chained_data_delayed_26__29_,
  chained_data_delayed_26__28_,chained_data_delayed_26__27_,chained_data_delayed_26__26_,
  chained_data_delayed_26__25_,chained_data_delayed_26__24_,chained_data_delayed_26__23_,
  chained_data_delayed_26__22_,chained_data_delayed_26__21_,
  chained_data_delayed_26__20_,chained_data_delayed_26__19_,chained_data_delayed_26__18_,
  chained_data_delayed_26__17_,chained_data_delayed_26__16_,chained_data_delayed_26__15_,
  chained_data_delayed_26__14_,chained_data_delayed_26__13_,chained_data_delayed_26__12_,
  chained_data_delayed_26__11_,chained_data_delayed_26__10_,chained_data_delayed_26__9_,
  chained_data_delayed_26__8_,chained_data_delayed_26__7_,
  chained_data_delayed_26__6_,chained_data_delayed_26__5_,chained_data_delayed_26__4_,
  chained_data_delayed_26__3_,chained_data_delayed_26__2_,chained_data_delayed_26__1_,
  chained_data_delayed_26__0_,chained_data_delayed_25__127_,chained_data_delayed_25__126_,
  chained_data_delayed_25__125_,chained_data_delayed_25__124_,
  chained_data_delayed_25__123_,chained_data_delayed_25__122_,chained_data_delayed_25__121_,
  chained_data_delayed_25__120_,chained_data_delayed_25__119_,chained_data_delayed_25__118_,
  chained_data_delayed_25__117_,chained_data_delayed_25__116_,
  chained_data_delayed_25__115_,chained_data_delayed_25__114_,chained_data_delayed_25__113_,
  chained_data_delayed_25__112_,chained_data_delayed_25__111_,chained_data_delayed_25__110_,
  chained_data_delayed_25__109_,chained_data_delayed_25__108_,
  chained_data_delayed_25__107_,chained_data_delayed_25__106_,chained_data_delayed_25__105_,
  chained_data_delayed_25__104_,chained_data_delayed_25__103_,chained_data_delayed_25__102_,
  chained_data_delayed_25__101_,chained_data_delayed_25__100_,
  chained_data_delayed_25__99_,chained_data_delayed_25__98_,chained_data_delayed_25__97_,
  chained_data_delayed_25__96_,chained_data_delayed_25__95_,chained_data_delayed_25__94_,
  chained_data_delayed_25__93_,chained_data_delayed_25__92_,chained_data_delayed_25__91_,
  chained_data_delayed_25__90_,chained_data_delayed_25__89_,chained_data_delayed_25__88_,
  chained_data_delayed_25__87_,chained_data_delayed_25__86_,
  chained_data_delayed_25__85_,chained_data_delayed_25__84_,chained_data_delayed_25__83_,
  chained_data_delayed_25__82_,chained_data_delayed_25__81_,chained_data_delayed_25__80_,
  chained_data_delayed_25__79_,chained_data_delayed_25__78_,chained_data_delayed_25__77_,
  chained_data_delayed_25__76_,chained_data_delayed_25__75_,
  chained_data_delayed_25__74_,chained_data_delayed_25__73_,chained_data_delayed_25__72_,
  chained_data_delayed_25__71_,chained_data_delayed_25__70_,chained_data_delayed_25__69_,
  chained_data_delayed_25__68_,chained_data_delayed_25__67_,chained_data_delayed_25__66_,
  chained_data_delayed_25__65_,chained_data_delayed_25__64_,
  chained_data_delayed_25__63_,chained_data_delayed_25__62_,chained_data_delayed_25__61_,
  chained_data_delayed_25__60_,chained_data_delayed_25__59_,chained_data_delayed_25__58_,
  chained_data_delayed_25__57_,chained_data_delayed_25__56_,chained_data_delayed_25__55_,
  chained_data_delayed_25__54_,chained_data_delayed_25__53_,
  chained_data_delayed_25__52_,chained_data_delayed_25__51_,chained_data_delayed_25__50_,
  chained_data_delayed_25__49_,chained_data_delayed_25__48_,chained_data_delayed_25__47_,
  chained_data_delayed_25__46_,chained_data_delayed_25__45_,chained_data_delayed_25__44_,
  chained_data_delayed_25__43_,chained_data_delayed_25__42_,
  chained_data_delayed_25__41_,chained_data_delayed_25__40_,chained_data_delayed_25__39_,
  chained_data_delayed_25__38_,chained_data_delayed_25__37_,chained_data_delayed_25__36_,
  chained_data_delayed_25__35_,chained_data_delayed_25__34_,chained_data_delayed_25__33_,
  chained_data_delayed_25__32_,chained_data_delayed_25__31_,
  chained_data_delayed_25__30_,chained_data_delayed_25__29_,chained_data_delayed_25__28_,
  chained_data_delayed_25__27_,chained_data_delayed_25__26_,chained_data_delayed_25__25_,
  chained_data_delayed_25__24_,chained_data_delayed_25__23_,chained_data_delayed_25__22_,
  chained_data_delayed_25__21_,chained_data_delayed_25__20_,
  chained_data_delayed_25__19_,chained_data_delayed_25__18_,chained_data_delayed_25__17_,
  chained_data_delayed_25__16_,chained_data_delayed_25__15_,chained_data_delayed_25__14_,
  chained_data_delayed_25__13_,chained_data_delayed_25__12_,chained_data_delayed_25__11_,
  chained_data_delayed_25__10_,chained_data_delayed_25__9_,chained_data_delayed_25__8_,
  chained_data_delayed_25__7_,chained_data_delayed_25__6_,
  chained_data_delayed_25__5_,chained_data_delayed_25__4_,chained_data_delayed_25__3_,
  chained_data_delayed_25__2_,chained_data_delayed_25__1_,chained_data_delayed_25__0_,
  chained_data_delayed_32__127_,chained_data_delayed_32__126_,chained_data_delayed_32__125_,
  chained_data_delayed_32__124_,chained_data_delayed_32__123_,
  chained_data_delayed_32__122_,chained_data_delayed_32__121_,chained_data_delayed_32__120_,
  chained_data_delayed_32__119_,chained_data_delayed_32__118_,chained_data_delayed_32__117_,
  chained_data_delayed_32__116_,chained_data_delayed_32__115_,
  chained_data_delayed_32__114_,chained_data_delayed_32__113_,chained_data_delayed_32__112_,
  chained_data_delayed_32__111_,chained_data_delayed_32__110_,chained_data_delayed_32__109_,
  chained_data_delayed_32__108_,chained_data_delayed_32__107_,
  chained_data_delayed_32__106_,chained_data_delayed_32__105_,chained_data_delayed_32__104_,
  chained_data_delayed_32__103_,chained_data_delayed_32__102_,chained_data_delayed_32__101_,
  chained_data_delayed_32__100_,chained_data_delayed_32__99_,chained_data_delayed_32__98_,
  chained_data_delayed_32__97_,chained_data_delayed_32__96_,
  chained_data_delayed_32__95_,chained_data_delayed_32__94_,chained_data_delayed_32__93_,
  chained_data_delayed_32__92_,chained_data_delayed_32__91_,chained_data_delayed_32__90_,
  chained_data_delayed_32__89_,chained_data_delayed_32__88_,chained_data_delayed_32__87_,
  chained_data_delayed_32__86_,chained_data_delayed_32__85_,
  chained_data_delayed_32__84_,chained_data_delayed_32__83_,chained_data_delayed_32__82_,
  chained_data_delayed_32__81_,chained_data_delayed_32__80_,chained_data_delayed_32__79_,
  chained_data_delayed_32__78_,chained_data_delayed_32__77_,chained_data_delayed_32__76_,
  chained_data_delayed_32__75_,chained_data_delayed_32__74_,
  chained_data_delayed_32__73_,chained_data_delayed_32__72_,chained_data_delayed_32__71_,
  chained_data_delayed_32__70_,chained_data_delayed_32__69_,chained_data_delayed_32__68_,
  chained_data_delayed_32__67_,chained_data_delayed_32__66_,chained_data_delayed_32__65_,
  chained_data_delayed_32__64_,chained_data_delayed_32__63_,
  chained_data_delayed_32__62_,chained_data_delayed_32__61_,chained_data_delayed_32__60_,
  chained_data_delayed_32__59_,chained_data_delayed_32__58_,chained_data_delayed_32__57_,
  chained_data_delayed_32__56_,chained_data_delayed_32__55_,chained_data_delayed_32__54_,
  chained_data_delayed_32__53_,chained_data_delayed_32__52_,
  chained_data_delayed_32__51_,chained_data_delayed_32__50_,chained_data_delayed_32__49_,
  chained_data_delayed_32__48_,chained_data_delayed_32__47_,chained_data_delayed_32__46_,
  chained_data_delayed_32__45_,chained_data_delayed_32__44_,chained_data_delayed_32__43_,
  chained_data_delayed_32__42_,chained_data_delayed_32__41_,
  chained_data_delayed_32__40_,chained_data_delayed_32__39_,chained_data_delayed_32__38_,
  chained_data_delayed_32__37_,chained_data_delayed_32__36_,chained_data_delayed_32__35_,
  chained_data_delayed_32__34_,chained_data_delayed_32__33_,chained_data_delayed_32__32_,
  chained_data_delayed_32__31_,chained_data_delayed_32__30_,
  chained_data_delayed_32__29_,chained_data_delayed_32__28_,chained_data_delayed_32__27_,
  chained_data_delayed_32__26_,chained_data_delayed_32__25_,chained_data_delayed_32__24_,
  chained_data_delayed_32__23_,chained_data_delayed_32__22_,chained_data_delayed_32__21_,
  chained_data_delayed_32__20_,chained_data_delayed_32__19_,chained_data_delayed_32__18_,
  chained_data_delayed_32__17_,chained_data_delayed_32__16_,
  chained_data_delayed_32__15_,chained_data_delayed_32__14_,chained_data_delayed_32__13_,
  chained_data_delayed_32__12_,chained_data_delayed_32__11_,chained_data_delayed_32__10_,
  chained_data_delayed_32__9_,chained_data_delayed_32__8_,chained_data_delayed_32__7_,
  chained_data_delayed_32__6_,chained_data_delayed_32__5_,chained_data_delayed_32__4_,
  chained_data_delayed_32__3_,chained_data_delayed_32__2_,
  chained_data_delayed_32__1_,chained_data_delayed_32__0_,chained_data_delayed_31__127_,
  chained_data_delayed_31__126_,chained_data_delayed_31__125_,chained_data_delayed_31__124_,
  chained_data_delayed_31__123_,chained_data_delayed_31__122_,
  chained_data_delayed_31__121_,chained_data_delayed_31__120_,chained_data_delayed_31__119_,
  chained_data_delayed_31__118_,chained_data_delayed_31__117_,chained_data_delayed_31__116_,
  chained_data_delayed_31__115_,chained_data_delayed_31__114_,
  chained_data_delayed_31__113_,chained_data_delayed_31__112_,chained_data_delayed_31__111_,
  chained_data_delayed_31__110_,chained_data_delayed_31__109_,chained_data_delayed_31__108_,
  chained_data_delayed_31__107_,chained_data_delayed_31__106_,
  chained_data_delayed_31__105_,chained_data_delayed_31__104_,chained_data_delayed_31__103_,
  chained_data_delayed_31__102_,chained_data_delayed_31__101_,chained_data_delayed_31__100_,
  chained_data_delayed_31__99_,chained_data_delayed_31__98_,chained_data_delayed_31__97_,
  chained_data_delayed_31__96_,chained_data_delayed_31__95_,
  chained_data_delayed_31__94_,chained_data_delayed_31__93_,chained_data_delayed_31__92_,
  chained_data_delayed_31__91_,chained_data_delayed_31__90_,chained_data_delayed_31__89_,
  chained_data_delayed_31__88_,chained_data_delayed_31__87_,chained_data_delayed_31__86_,
  chained_data_delayed_31__85_,chained_data_delayed_31__84_,
  chained_data_delayed_31__83_,chained_data_delayed_31__82_,chained_data_delayed_31__81_,
  chained_data_delayed_31__80_,chained_data_delayed_31__79_,chained_data_delayed_31__78_,
  chained_data_delayed_31__77_,chained_data_delayed_31__76_,chained_data_delayed_31__75_,
  chained_data_delayed_31__74_,chained_data_delayed_31__73_,
  chained_data_delayed_31__72_,chained_data_delayed_31__71_,chained_data_delayed_31__70_,
  chained_data_delayed_31__69_,chained_data_delayed_31__68_,chained_data_delayed_31__67_,
  chained_data_delayed_31__66_,chained_data_delayed_31__65_,chained_data_delayed_31__64_,
  chained_data_delayed_31__63_,chained_data_delayed_31__62_,
  chained_data_delayed_31__61_,chained_data_delayed_31__60_,chained_data_delayed_31__59_,
  chained_data_delayed_31__58_,chained_data_delayed_31__57_,chained_data_delayed_31__56_,
  chained_data_delayed_31__55_,chained_data_delayed_31__54_,chained_data_delayed_31__53_,
  chained_data_delayed_31__52_,chained_data_delayed_31__51_,
  chained_data_delayed_31__50_,chained_data_delayed_31__49_,chained_data_delayed_31__48_,
  chained_data_delayed_31__47_,chained_data_delayed_31__46_,chained_data_delayed_31__45_,
  chained_data_delayed_31__44_,chained_data_delayed_31__43_,chained_data_delayed_31__42_,
  chained_data_delayed_31__41_,chained_data_delayed_31__40_,
  chained_data_delayed_31__39_,chained_data_delayed_31__38_,chained_data_delayed_31__37_,
  chained_data_delayed_31__36_,chained_data_delayed_31__35_,chained_data_delayed_31__34_,
  chained_data_delayed_31__33_,chained_data_delayed_31__32_,chained_data_delayed_31__31_,
  chained_data_delayed_31__30_,chained_data_delayed_31__29_,chained_data_delayed_31__28_,
  chained_data_delayed_31__27_,chained_data_delayed_31__26_,
  chained_data_delayed_31__25_,chained_data_delayed_31__24_,chained_data_delayed_31__23_,
  chained_data_delayed_31__22_,chained_data_delayed_31__21_,chained_data_delayed_31__20_,
  chained_data_delayed_31__19_,chained_data_delayed_31__18_,chained_data_delayed_31__17_,
  chained_data_delayed_31__16_,chained_data_delayed_31__15_,
  chained_data_delayed_31__14_,chained_data_delayed_31__13_,chained_data_delayed_31__12_,
  chained_data_delayed_31__11_,chained_data_delayed_31__10_,chained_data_delayed_31__9_,
  chained_data_delayed_31__8_,chained_data_delayed_31__7_,chained_data_delayed_31__6_,
  chained_data_delayed_31__5_,chained_data_delayed_31__4_,chained_data_delayed_31__3_,
  chained_data_delayed_31__2_,chained_data_delayed_31__1_,
  chained_data_delayed_31__0_,chained_data_delayed_30__127_,chained_data_delayed_30__126_,
  chained_data_delayed_30__125_,chained_data_delayed_30__124_,chained_data_delayed_30__123_,
  chained_data_delayed_30__122_,chained_data_delayed_30__121_,
  chained_data_delayed_30__120_,chained_data_delayed_30__119_,chained_data_delayed_30__118_,
  chained_data_delayed_30__117_,chained_data_delayed_30__116_,chained_data_delayed_30__115_,
  chained_data_delayed_30__114_,chained_data_delayed_30__113_,
  chained_data_delayed_30__112_,chained_data_delayed_30__111_,chained_data_delayed_30__110_,
  chained_data_delayed_30__109_,chained_data_delayed_30__108_,chained_data_delayed_30__107_,
  chained_data_delayed_30__106_,chained_data_delayed_30__105_,
  chained_data_delayed_30__104_,chained_data_delayed_30__103_,chained_data_delayed_30__102_,
  chained_data_delayed_30__101_,chained_data_delayed_30__100_,chained_data_delayed_30__99_,
  chained_data_delayed_30__98_,chained_data_delayed_30__97_,chained_data_delayed_30__96_,
  chained_data_delayed_30__95_,chained_data_delayed_30__94_,
  chained_data_delayed_30__93_,chained_data_delayed_30__92_,chained_data_delayed_30__91_,
  chained_data_delayed_30__90_,chained_data_delayed_30__89_,chained_data_delayed_30__88_,
  chained_data_delayed_30__87_,chained_data_delayed_30__86_,chained_data_delayed_30__85_,
  chained_data_delayed_30__84_,chained_data_delayed_30__83_,
  chained_data_delayed_30__82_,chained_data_delayed_30__81_,chained_data_delayed_30__80_,
  chained_data_delayed_30__79_,chained_data_delayed_30__78_,chained_data_delayed_30__77_,
  chained_data_delayed_30__76_,chained_data_delayed_30__75_,chained_data_delayed_30__74_,
  chained_data_delayed_30__73_,chained_data_delayed_30__72_,
  chained_data_delayed_30__71_,chained_data_delayed_30__70_,chained_data_delayed_30__69_,
  chained_data_delayed_30__68_,chained_data_delayed_30__67_,chained_data_delayed_30__66_,
  chained_data_delayed_30__65_,chained_data_delayed_30__64_,chained_data_delayed_30__63_,
  chained_data_delayed_30__62_,chained_data_delayed_30__61_,
  chained_data_delayed_30__60_,chained_data_delayed_30__59_,chained_data_delayed_30__58_,
  chained_data_delayed_30__57_,chained_data_delayed_30__56_,chained_data_delayed_30__55_,
  chained_data_delayed_30__54_,chained_data_delayed_30__53_,chained_data_delayed_30__52_,
  chained_data_delayed_30__51_,chained_data_delayed_30__50_,
  chained_data_delayed_30__49_,chained_data_delayed_30__48_,chained_data_delayed_30__47_,
  chained_data_delayed_30__46_,chained_data_delayed_30__45_,chained_data_delayed_30__44_,
  chained_data_delayed_30__43_,chained_data_delayed_30__42_,chained_data_delayed_30__41_,
  chained_data_delayed_30__40_,chained_data_delayed_30__39_,chained_data_delayed_30__38_,
  chained_data_delayed_30__37_,chained_data_delayed_30__36_,
  chained_data_delayed_30__35_,chained_data_delayed_30__34_,chained_data_delayed_30__33_,
  chained_data_delayed_30__32_,chained_data_delayed_30__31_,chained_data_delayed_30__30_,
  chained_data_delayed_30__29_,chained_data_delayed_30__28_,chained_data_delayed_30__27_,
  chained_data_delayed_30__26_,chained_data_delayed_30__25_,
  chained_data_delayed_30__24_,chained_data_delayed_30__23_,chained_data_delayed_30__22_,
  chained_data_delayed_30__21_,chained_data_delayed_30__20_,chained_data_delayed_30__19_,
  chained_data_delayed_30__18_,chained_data_delayed_30__17_,chained_data_delayed_30__16_,
  chained_data_delayed_30__15_,chained_data_delayed_30__14_,
  chained_data_delayed_30__13_,chained_data_delayed_30__12_,chained_data_delayed_30__11_,
  chained_data_delayed_30__10_,chained_data_delayed_30__9_,chained_data_delayed_30__8_,
  chained_data_delayed_30__7_,chained_data_delayed_30__6_,chained_data_delayed_30__5_,
  chained_data_delayed_30__4_,chained_data_delayed_30__3_,chained_data_delayed_30__2_,
  chained_data_delayed_30__1_,chained_data_delayed_30__0_,
  chained_data_delayed_29__127_,chained_data_delayed_29__126_,chained_data_delayed_29__125_,
  chained_data_delayed_29__124_,chained_data_delayed_29__123_,chained_data_delayed_29__122_,
  chained_data_delayed_29__121_,chained_data_delayed_29__120_,
  chained_data_delayed_29__119_,chained_data_delayed_29__118_,chained_data_delayed_29__117_,
  chained_data_delayed_29__116_,chained_data_delayed_29__115_,chained_data_delayed_29__114_,
  chained_data_delayed_29__113_,chained_data_delayed_29__112_,
  chained_data_delayed_29__111_,chained_data_delayed_29__110_,chained_data_delayed_29__109_,
  chained_data_delayed_29__108_,chained_data_delayed_29__107_,chained_data_delayed_29__106_,
  chained_data_delayed_29__105_,chained_data_delayed_29__104_,
  chained_data_delayed_29__103_,chained_data_delayed_29__102_,chained_data_delayed_29__101_,
  chained_data_delayed_29__100_,chained_data_delayed_29__99_,chained_data_delayed_29__98_,
  chained_data_delayed_29__97_,chained_data_delayed_29__96_,chained_data_delayed_29__95_,
  chained_data_delayed_29__94_,chained_data_delayed_29__93_,
  chained_data_delayed_29__92_,chained_data_delayed_29__91_,chained_data_delayed_29__90_,
  chained_data_delayed_29__89_,chained_data_delayed_29__88_,chained_data_delayed_29__87_,
  chained_data_delayed_29__86_,chained_data_delayed_29__85_,chained_data_delayed_29__84_,
  chained_data_delayed_29__83_,chained_data_delayed_29__82_,
  chained_data_delayed_29__81_,chained_data_delayed_29__80_,chained_data_delayed_29__79_,
  chained_data_delayed_29__78_,chained_data_delayed_29__77_,chained_data_delayed_29__76_,
  chained_data_delayed_29__75_,chained_data_delayed_29__74_,chained_data_delayed_29__73_,
  chained_data_delayed_29__72_,chained_data_delayed_29__71_,
  chained_data_delayed_29__70_,chained_data_delayed_29__69_,chained_data_delayed_29__68_,
  chained_data_delayed_29__67_,chained_data_delayed_29__66_,chained_data_delayed_29__65_,
  chained_data_delayed_29__64_,chained_data_delayed_29__63_,chained_data_delayed_29__62_,
  chained_data_delayed_29__61_,chained_data_delayed_29__60_,
  chained_data_delayed_29__59_,chained_data_delayed_29__58_,chained_data_delayed_29__57_,
  chained_data_delayed_29__56_,chained_data_delayed_29__55_,chained_data_delayed_29__54_,
  chained_data_delayed_29__53_,chained_data_delayed_29__52_,chained_data_delayed_29__51_,
  chained_data_delayed_29__50_,chained_data_delayed_29__49_,chained_data_delayed_29__48_,
  chained_data_delayed_29__47_,chained_data_delayed_29__46_,
  chained_data_delayed_29__45_,chained_data_delayed_29__44_,chained_data_delayed_29__43_,
  chained_data_delayed_29__42_,chained_data_delayed_29__41_,chained_data_delayed_29__40_,
  chained_data_delayed_29__39_,chained_data_delayed_29__38_,chained_data_delayed_29__37_,
  chained_data_delayed_29__36_,chained_data_delayed_29__35_,
  chained_data_delayed_29__34_,chained_data_delayed_29__33_,chained_data_delayed_29__32_,
  chained_data_delayed_29__31_,chained_data_delayed_29__30_,chained_data_delayed_29__29_,
  chained_data_delayed_29__28_,chained_data_delayed_29__27_,chained_data_delayed_29__26_,
  chained_data_delayed_29__25_,chained_data_delayed_29__24_,
  chained_data_delayed_29__23_,chained_data_delayed_29__22_,chained_data_delayed_29__21_,
  chained_data_delayed_29__20_,chained_data_delayed_29__19_,chained_data_delayed_29__18_,
  chained_data_delayed_29__17_,chained_data_delayed_29__16_,chained_data_delayed_29__15_,
  chained_data_delayed_29__14_,chained_data_delayed_29__13_,
  chained_data_delayed_29__12_,chained_data_delayed_29__11_,chained_data_delayed_29__10_,
  chained_data_delayed_29__9_,chained_data_delayed_29__8_,chained_data_delayed_29__7_,
  chained_data_delayed_29__6_,chained_data_delayed_29__5_,chained_data_delayed_29__4_,
  chained_data_delayed_29__3_,chained_data_delayed_29__2_,chained_data_delayed_29__1_,
  chained_data_delayed_29__0_,chained_data_delayed_36__127_,
  chained_data_delayed_36__126_,chained_data_delayed_36__125_,chained_data_delayed_36__124_,
  chained_data_delayed_36__123_,chained_data_delayed_36__122_,chained_data_delayed_36__121_,
  chained_data_delayed_36__120_,chained_data_delayed_36__119_,
  chained_data_delayed_36__118_,chained_data_delayed_36__117_,chained_data_delayed_36__116_,
  chained_data_delayed_36__115_,chained_data_delayed_36__114_,chained_data_delayed_36__113_,
  chained_data_delayed_36__112_,chained_data_delayed_36__111_,
  chained_data_delayed_36__110_,chained_data_delayed_36__109_,chained_data_delayed_36__108_,
  chained_data_delayed_36__107_,chained_data_delayed_36__106_,chained_data_delayed_36__105_,
  chained_data_delayed_36__104_,chained_data_delayed_36__103_,
  chained_data_delayed_36__102_,chained_data_delayed_36__101_,chained_data_delayed_36__100_,
  chained_data_delayed_36__99_,chained_data_delayed_36__98_,chained_data_delayed_36__97_,
  chained_data_delayed_36__96_,chained_data_delayed_36__95_,chained_data_delayed_36__94_,
  chained_data_delayed_36__93_,chained_data_delayed_36__92_,
  chained_data_delayed_36__91_,chained_data_delayed_36__90_,chained_data_delayed_36__89_,
  chained_data_delayed_36__88_,chained_data_delayed_36__87_,chained_data_delayed_36__86_,
  chained_data_delayed_36__85_,chained_data_delayed_36__84_,chained_data_delayed_36__83_,
  chained_data_delayed_36__82_,chained_data_delayed_36__81_,
  chained_data_delayed_36__80_,chained_data_delayed_36__79_,chained_data_delayed_36__78_,
  chained_data_delayed_36__77_,chained_data_delayed_36__76_,chained_data_delayed_36__75_,
  chained_data_delayed_36__74_,chained_data_delayed_36__73_,chained_data_delayed_36__72_,
  chained_data_delayed_36__71_,chained_data_delayed_36__70_,
  chained_data_delayed_36__69_,chained_data_delayed_36__68_,chained_data_delayed_36__67_,
  chained_data_delayed_36__66_,chained_data_delayed_36__65_,chained_data_delayed_36__64_,
  chained_data_delayed_36__63_,chained_data_delayed_36__62_,chained_data_delayed_36__61_,
  chained_data_delayed_36__60_,chained_data_delayed_36__59_,chained_data_delayed_36__58_,
  chained_data_delayed_36__57_,chained_data_delayed_36__56_,
  chained_data_delayed_36__55_,chained_data_delayed_36__54_,chained_data_delayed_36__53_,
  chained_data_delayed_36__52_,chained_data_delayed_36__51_,chained_data_delayed_36__50_,
  chained_data_delayed_36__49_,chained_data_delayed_36__48_,chained_data_delayed_36__47_,
  chained_data_delayed_36__46_,chained_data_delayed_36__45_,
  chained_data_delayed_36__44_,chained_data_delayed_36__43_,chained_data_delayed_36__42_,
  chained_data_delayed_36__41_,chained_data_delayed_36__40_,chained_data_delayed_36__39_,
  chained_data_delayed_36__38_,chained_data_delayed_36__37_,chained_data_delayed_36__36_,
  chained_data_delayed_36__35_,chained_data_delayed_36__34_,
  chained_data_delayed_36__33_,chained_data_delayed_36__32_,chained_data_delayed_36__31_,
  chained_data_delayed_36__30_,chained_data_delayed_36__29_,chained_data_delayed_36__28_,
  chained_data_delayed_36__27_,chained_data_delayed_36__26_,chained_data_delayed_36__25_,
  chained_data_delayed_36__24_,chained_data_delayed_36__23_,
  chained_data_delayed_36__22_,chained_data_delayed_36__21_,chained_data_delayed_36__20_,
  chained_data_delayed_36__19_,chained_data_delayed_36__18_,chained_data_delayed_36__17_,
  chained_data_delayed_36__16_,chained_data_delayed_36__15_,chained_data_delayed_36__14_,
  chained_data_delayed_36__13_,chained_data_delayed_36__12_,
  chained_data_delayed_36__11_,chained_data_delayed_36__10_,chained_data_delayed_36__9_,
  chained_data_delayed_36__8_,chained_data_delayed_36__7_,chained_data_delayed_36__6_,
  chained_data_delayed_36__5_,chained_data_delayed_36__4_,chained_data_delayed_36__3_,
  chained_data_delayed_36__2_,chained_data_delayed_36__1_,chained_data_delayed_36__0_,
  chained_data_delayed_35__127_,chained_data_delayed_35__126_,
  chained_data_delayed_35__125_,chained_data_delayed_35__124_,chained_data_delayed_35__123_,
  chained_data_delayed_35__122_,chained_data_delayed_35__121_,chained_data_delayed_35__120_,
  chained_data_delayed_35__119_,chained_data_delayed_35__118_,
  chained_data_delayed_35__117_,chained_data_delayed_35__116_,chained_data_delayed_35__115_,
  chained_data_delayed_35__114_,chained_data_delayed_35__113_,chained_data_delayed_35__112_,
  chained_data_delayed_35__111_,chained_data_delayed_35__110_,
  chained_data_delayed_35__109_,chained_data_delayed_35__108_,chained_data_delayed_35__107_,
  chained_data_delayed_35__106_,chained_data_delayed_35__105_,chained_data_delayed_35__104_,
  chained_data_delayed_35__103_,chained_data_delayed_35__102_,
  chained_data_delayed_35__101_,chained_data_delayed_35__100_,chained_data_delayed_35__99_,
  chained_data_delayed_35__98_,chained_data_delayed_35__97_,chained_data_delayed_35__96_,
  chained_data_delayed_35__95_,chained_data_delayed_35__94_,chained_data_delayed_35__93_,
  chained_data_delayed_35__92_,chained_data_delayed_35__91_,
  chained_data_delayed_35__90_,chained_data_delayed_35__89_,chained_data_delayed_35__88_,
  chained_data_delayed_35__87_,chained_data_delayed_35__86_,chained_data_delayed_35__85_,
  chained_data_delayed_35__84_,chained_data_delayed_35__83_,chained_data_delayed_35__82_,
  chained_data_delayed_35__81_,chained_data_delayed_35__80_,
  chained_data_delayed_35__79_,chained_data_delayed_35__78_,chained_data_delayed_35__77_,
  chained_data_delayed_35__76_,chained_data_delayed_35__75_,chained_data_delayed_35__74_,
  chained_data_delayed_35__73_,chained_data_delayed_35__72_,chained_data_delayed_35__71_,
  chained_data_delayed_35__70_,chained_data_delayed_35__69_,chained_data_delayed_35__68_,
  chained_data_delayed_35__67_,chained_data_delayed_35__66_,
  chained_data_delayed_35__65_,chained_data_delayed_35__64_,chained_data_delayed_35__63_,
  chained_data_delayed_35__62_,chained_data_delayed_35__61_,chained_data_delayed_35__60_,
  chained_data_delayed_35__59_,chained_data_delayed_35__58_,chained_data_delayed_35__57_,
  chained_data_delayed_35__56_,chained_data_delayed_35__55_,
  chained_data_delayed_35__54_,chained_data_delayed_35__53_,chained_data_delayed_35__52_,
  chained_data_delayed_35__51_,chained_data_delayed_35__50_,chained_data_delayed_35__49_,
  chained_data_delayed_35__48_,chained_data_delayed_35__47_,chained_data_delayed_35__46_,
  chained_data_delayed_35__45_,chained_data_delayed_35__44_,
  chained_data_delayed_35__43_,chained_data_delayed_35__42_,chained_data_delayed_35__41_,
  chained_data_delayed_35__40_,chained_data_delayed_35__39_,chained_data_delayed_35__38_,
  chained_data_delayed_35__37_,chained_data_delayed_35__36_,chained_data_delayed_35__35_,
  chained_data_delayed_35__34_,chained_data_delayed_35__33_,
  chained_data_delayed_35__32_,chained_data_delayed_35__31_,chained_data_delayed_35__30_,
  chained_data_delayed_35__29_,chained_data_delayed_35__28_,chained_data_delayed_35__27_,
  chained_data_delayed_35__26_,chained_data_delayed_35__25_,chained_data_delayed_35__24_,
  chained_data_delayed_35__23_,chained_data_delayed_35__22_,
  chained_data_delayed_35__21_,chained_data_delayed_35__20_,chained_data_delayed_35__19_,
  chained_data_delayed_35__18_,chained_data_delayed_35__17_,chained_data_delayed_35__16_,
  chained_data_delayed_35__15_,chained_data_delayed_35__14_,chained_data_delayed_35__13_,
  chained_data_delayed_35__12_,chained_data_delayed_35__11_,
  chained_data_delayed_35__10_,chained_data_delayed_35__9_,chained_data_delayed_35__8_,
  chained_data_delayed_35__7_,chained_data_delayed_35__6_,chained_data_delayed_35__5_,
  chained_data_delayed_35__4_,chained_data_delayed_35__3_,chained_data_delayed_35__2_,
  chained_data_delayed_35__1_,chained_data_delayed_35__0_,chained_data_delayed_34__127_,
  chained_data_delayed_34__126_,chained_data_delayed_34__125_,
  chained_data_delayed_34__124_,chained_data_delayed_34__123_,chained_data_delayed_34__122_,
  chained_data_delayed_34__121_,chained_data_delayed_34__120_,chained_data_delayed_34__119_,
  chained_data_delayed_34__118_,chained_data_delayed_34__117_,
  chained_data_delayed_34__116_,chained_data_delayed_34__115_,chained_data_delayed_34__114_,
  chained_data_delayed_34__113_,chained_data_delayed_34__112_,chained_data_delayed_34__111_,
  chained_data_delayed_34__110_,chained_data_delayed_34__109_,
  chained_data_delayed_34__108_,chained_data_delayed_34__107_,chained_data_delayed_34__106_,
  chained_data_delayed_34__105_,chained_data_delayed_34__104_,chained_data_delayed_34__103_,
  chained_data_delayed_34__102_,chained_data_delayed_34__101_,
  chained_data_delayed_34__100_,chained_data_delayed_34__99_,chained_data_delayed_34__98_,
  chained_data_delayed_34__97_,chained_data_delayed_34__96_,chained_data_delayed_34__95_,
  chained_data_delayed_34__94_,chained_data_delayed_34__93_,chained_data_delayed_34__92_,
  chained_data_delayed_34__91_,chained_data_delayed_34__90_,
  chained_data_delayed_34__89_,chained_data_delayed_34__88_,chained_data_delayed_34__87_,
  chained_data_delayed_34__86_,chained_data_delayed_34__85_,chained_data_delayed_34__84_,
  chained_data_delayed_34__83_,chained_data_delayed_34__82_,chained_data_delayed_34__81_,
  chained_data_delayed_34__80_,chained_data_delayed_34__79_,chained_data_delayed_34__78_,
  chained_data_delayed_34__77_,chained_data_delayed_34__76_,
  chained_data_delayed_34__75_,chained_data_delayed_34__74_,chained_data_delayed_34__73_,
  chained_data_delayed_34__72_,chained_data_delayed_34__71_,chained_data_delayed_34__70_,
  chained_data_delayed_34__69_,chained_data_delayed_34__68_,chained_data_delayed_34__67_,
  chained_data_delayed_34__66_,chained_data_delayed_34__65_,
  chained_data_delayed_34__64_,chained_data_delayed_34__63_,chained_data_delayed_34__62_,
  chained_data_delayed_34__61_,chained_data_delayed_34__60_,chained_data_delayed_34__59_,
  chained_data_delayed_34__58_,chained_data_delayed_34__57_,chained_data_delayed_34__56_,
  chained_data_delayed_34__55_,chained_data_delayed_34__54_,
  chained_data_delayed_34__53_,chained_data_delayed_34__52_,chained_data_delayed_34__51_,
  chained_data_delayed_34__50_,chained_data_delayed_34__49_,chained_data_delayed_34__48_,
  chained_data_delayed_34__47_,chained_data_delayed_34__46_,chained_data_delayed_34__45_,
  chained_data_delayed_34__44_,chained_data_delayed_34__43_,
  chained_data_delayed_34__42_,chained_data_delayed_34__41_,chained_data_delayed_34__40_,
  chained_data_delayed_34__39_,chained_data_delayed_34__38_,chained_data_delayed_34__37_,
  chained_data_delayed_34__36_,chained_data_delayed_34__35_,chained_data_delayed_34__34_,
  chained_data_delayed_34__33_,chained_data_delayed_34__32_,
  chained_data_delayed_34__31_,chained_data_delayed_34__30_,chained_data_delayed_34__29_,
  chained_data_delayed_34__28_,chained_data_delayed_34__27_,chained_data_delayed_34__26_,
  chained_data_delayed_34__25_,chained_data_delayed_34__24_,chained_data_delayed_34__23_,
  chained_data_delayed_34__22_,chained_data_delayed_34__21_,
  chained_data_delayed_34__20_,chained_data_delayed_34__19_,chained_data_delayed_34__18_,
  chained_data_delayed_34__17_,chained_data_delayed_34__16_,chained_data_delayed_34__15_,
  chained_data_delayed_34__14_,chained_data_delayed_34__13_,chained_data_delayed_34__12_,
  chained_data_delayed_34__11_,chained_data_delayed_34__10_,chained_data_delayed_34__9_,
  chained_data_delayed_34__8_,chained_data_delayed_34__7_,
  chained_data_delayed_34__6_,chained_data_delayed_34__5_,chained_data_delayed_34__4_,
  chained_data_delayed_34__3_,chained_data_delayed_34__2_,chained_data_delayed_34__1_,
  chained_data_delayed_34__0_,chained_data_delayed_33__127_,chained_data_delayed_33__126_,
  chained_data_delayed_33__125_,chained_data_delayed_33__124_,
  chained_data_delayed_33__123_,chained_data_delayed_33__122_,chained_data_delayed_33__121_,
  chained_data_delayed_33__120_,chained_data_delayed_33__119_,chained_data_delayed_33__118_,
  chained_data_delayed_33__117_,chained_data_delayed_33__116_,
  chained_data_delayed_33__115_,chained_data_delayed_33__114_,chained_data_delayed_33__113_,
  chained_data_delayed_33__112_,chained_data_delayed_33__111_,chained_data_delayed_33__110_,
  chained_data_delayed_33__109_,chained_data_delayed_33__108_,
  chained_data_delayed_33__107_,chained_data_delayed_33__106_,chained_data_delayed_33__105_,
  chained_data_delayed_33__104_,chained_data_delayed_33__103_,chained_data_delayed_33__102_,
  chained_data_delayed_33__101_,chained_data_delayed_33__100_,
  chained_data_delayed_33__99_,chained_data_delayed_33__98_,chained_data_delayed_33__97_,
  chained_data_delayed_33__96_,chained_data_delayed_33__95_,chained_data_delayed_33__94_,
  chained_data_delayed_33__93_,chained_data_delayed_33__92_,chained_data_delayed_33__91_,
  chained_data_delayed_33__90_,chained_data_delayed_33__89_,chained_data_delayed_33__88_,
  chained_data_delayed_33__87_,chained_data_delayed_33__86_,
  chained_data_delayed_33__85_,chained_data_delayed_33__84_,chained_data_delayed_33__83_,
  chained_data_delayed_33__82_,chained_data_delayed_33__81_,chained_data_delayed_33__80_,
  chained_data_delayed_33__79_,chained_data_delayed_33__78_,chained_data_delayed_33__77_,
  chained_data_delayed_33__76_,chained_data_delayed_33__75_,
  chained_data_delayed_33__74_,chained_data_delayed_33__73_,chained_data_delayed_33__72_,
  chained_data_delayed_33__71_,chained_data_delayed_33__70_,chained_data_delayed_33__69_,
  chained_data_delayed_33__68_,chained_data_delayed_33__67_,chained_data_delayed_33__66_,
  chained_data_delayed_33__65_,chained_data_delayed_33__64_,
  chained_data_delayed_33__63_,chained_data_delayed_33__62_,chained_data_delayed_33__61_,
  chained_data_delayed_33__60_,chained_data_delayed_33__59_,chained_data_delayed_33__58_,
  chained_data_delayed_33__57_,chained_data_delayed_33__56_,chained_data_delayed_33__55_,
  chained_data_delayed_33__54_,chained_data_delayed_33__53_,
  chained_data_delayed_33__52_,chained_data_delayed_33__51_,chained_data_delayed_33__50_,
  chained_data_delayed_33__49_,chained_data_delayed_33__48_,chained_data_delayed_33__47_,
  chained_data_delayed_33__46_,chained_data_delayed_33__45_,chained_data_delayed_33__44_,
  chained_data_delayed_33__43_,chained_data_delayed_33__42_,
  chained_data_delayed_33__41_,chained_data_delayed_33__40_,chained_data_delayed_33__39_,
  chained_data_delayed_33__38_,chained_data_delayed_33__37_,chained_data_delayed_33__36_,
  chained_data_delayed_33__35_,chained_data_delayed_33__34_,chained_data_delayed_33__33_,
  chained_data_delayed_33__32_,chained_data_delayed_33__31_,
  chained_data_delayed_33__30_,chained_data_delayed_33__29_,chained_data_delayed_33__28_,
  chained_data_delayed_33__27_,chained_data_delayed_33__26_,chained_data_delayed_33__25_,
  chained_data_delayed_33__24_,chained_data_delayed_33__23_,chained_data_delayed_33__22_,
  chained_data_delayed_33__21_,chained_data_delayed_33__20_,
  chained_data_delayed_33__19_,chained_data_delayed_33__18_,chained_data_delayed_33__17_,
  chained_data_delayed_33__16_,chained_data_delayed_33__15_,chained_data_delayed_33__14_,
  chained_data_delayed_33__13_,chained_data_delayed_33__12_,chained_data_delayed_33__11_,
  chained_data_delayed_33__10_,chained_data_delayed_33__9_,chained_data_delayed_33__8_,
  chained_data_delayed_33__7_,chained_data_delayed_33__6_,
  chained_data_delayed_33__5_,chained_data_delayed_33__4_,chained_data_delayed_33__3_,
  chained_data_delayed_33__2_,chained_data_delayed_33__1_,chained_data_delayed_33__0_,
  chained_data_delayed_40__127_,chained_data_delayed_40__126_,chained_data_delayed_40__125_,
  chained_data_delayed_40__124_,chained_data_delayed_40__123_,
  chained_data_delayed_40__122_,chained_data_delayed_40__121_,chained_data_delayed_40__120_,
  chained_data_delayed_40__119_,chained_data_delayed_40__118_,chained_data_delayed_40__117_,
  chained_data_delayed_40__116_,chained_data_delayed_40__115_,
  chained_data_delayed_40__114_,chained_data_delayed_40__113_,chained_data_delayed_40__112_,
  chained_data_delayed_40__111_,chained_data_delayed_40__110_,chained_data_delayed_40__109_,
  chained_data_delayed_40__108_,chained_data_delayed_40__107_,
  chained_data_delayed_40__106_,chained_data_delayed_40__105_,chained_data_delayed_40__104_,
  chained_data_delayed_40__103_,chained_data_delayed_40__102_,chained_data_delayed_40__101_,
  chained_data_delayed_40__100_,chained_data_delayed_40__99_,chained_data_delayed_40__98_,
  chained_data_delayed_40__97_,chained_data_delayed_40__96_,
  chained_data_delayed_40__95_,chained_data_delayed_40__94_,chained_data_delayed_40__93_,
  chained_data_delayed_40__92_,chained_data_delayed_40__91_,chained_data_delayed_40__90_,
  chained_data_delayed_40__89_,chained_data_delayed_40__88_,chained_data_delayed_40__87_,
  chained_data_delayed_40__86_,chained_data_delayed_40__85_,
  chained_data_delayed_40__84_,chained_data_delayed_40__83_,chained_data_delayed_40__82_,
  chained_data_delayed_40__81_,chained_data_delayed_40__80_,chained_data_delayed_40__79_,
  chained_data_delayed_40__78_,chained_data_delayed_40__77_,chained_data_delayed_40__76_,
  chained_data_delayed_40__75_,chained_data_delayed_40__74_,
  chained_data_delayed_40__73_,chained_data_delayed_40__72_,chained_data_delayed_40__71_,
  chained_data_delayed_40__70_,chained_data_delayed_40__69_,chained_data_delayed_40__68_,
  chained_data_delayed_40__67_,chained_data_delayed_40__66_,chained_data_delayed_40__65_,
  chained_data_delayed_40__64_,chained_data_delayed_40__63_,
  chained_data_delayed_40__62_,chained_data_delayed_40__61_,chained_data_delayed_40__60_,
  chained_data_delayed_40__59_,chained_data_delayed_40__58_,chained_data_delayed_40__57_,
  chained_data_delayed_40__56_,chained_data_delayed_40__55_,chained_data_delayed_40__54_,
  chained_data_delayed_40__53_,chained_data_delayed_40__52_,
  chained_data_delayed_40__51_,chained_data_delayed_40__50_,chained_data_delayed_40__49_,
  chained_data_delayed_40__48_,chained_data_delayed_40__47_,chained_data_delayed_40__46_,
  chained_data_delayed_40__45_,chained_data_delayed_40__44_,chained_data_delayed_40__43_,
  chained_data_delayed_40__42_,chained_data_delayed_40__41_,
  chained_data_delayed_40__40_,chained_data_delayed_40__39_,chained_data_delayed_40__38_,
  chained_data_delayed_40__37_,chained_data_delayed_40__36_,chained_data_delayed_40__35_,
  chained_data_delayed_40__34_,chained_data_delayed_40__33_,chained_data_delayed_40__32_,
  chained_data_delayed_40__31_,chained_data_delayed_40__30_,
  chained_data_delayed_40__29_,chained_data_delayed_40__28_,chained_data_delayed_40__27_,
  chained_data_delayed_40__26_,chained_data_delayed_40__25_,chained_data_delayed_40__24_,
  chained_data_delayed_40__23_,chained_data_delayed_40__22_,chained_data_delayed_40__21_,
  chained_data_delayed_40__20_,chained_data_delayed_40__19_,chained_data_delayed_40__18_,
  chained_data_delayed_40__17_,chained_data_delayed_40__16_,
  chained_data_delayed_40__15_,chained_data_delayed_40__14_,chained_data_delayed_40__13_,
  chained_data_delayed_40__12_,chained_data_delayed_40__11_,chained_data_delayed_40__10_,
  chained_data_delayed_40__9_,chained_data_delayed_40__8_,chained_data_delayed_40__7_,
  chained_data_delayed_40__6_,chained_data_delayed_40__5_,chained_data_delayed_40__4_,
  chained_data_delayed_40__3_,chained_data_delayed_40__2_,
  chained_data_delayed_40__1_,chained_data_delayed_40__0_,chained_data_delayed_39__127_,
  chained_data_delayed_39__126_,chained_data_delayed_39__125_,chained_data_delayed_39__124_,
  chained_data_delayed_39__123_,chained_data_delayed_39__122_,
  chained_data_delayed_39__121_,chained_data_delayed_39__120_,chained_data_delayed_39__119_,
  chained_data_delayed_39__118_,chained_data_delayed_39__117_,chained_data_delayed_39__116_,
  chained_data_delayed_39__115_,chained_data_delayed_39__114_,
  chained_data_delayed_39__113_,chained_data_delayed_39__112_,chained_data_delayed_39__111_,
  chained_data_delayed_39__110_,chained_data_delayed_39__109_,chained_data_delayed_39__108_,
  chained_data_delayed_39__107_,chained_data_delayed_39__106_,
  chained_data_delayed_39__105_,chained_data_delayed_39__104_,chained_data_delayed_39__103_,
  chained_data_delayed_39__102_,chained_data_delayed_39__101_,chained_data_delayed_39__100_,
  chained_data_delayed_39__99_,chained_data_delayed_39__98_,chained_data_delayed_39__97_,
  chained_data_delayed_39__96_,chained_data_delayed_39__95_,
  chained_data_delayed_39__94_,chained_data_delayed_39__93_,chained_data_delayed_39__92_,
  chained_data_delayed_39__91_,chained_data_delayed_39__90_,chained_data_delayed_39__89_,
  chained_data_delayed_39__88_,chained_data_delayed_39__87_,chained_data_delayed_39__86_,
  chained_data_delayed_39__85_,chained_data_delayed_39__84_,
  chained_data_delayed_39__83_,chained_data_delayed_39__82_,chained_data_delayed_39__81_,
  chained_data_delayed_39__80_,chained_data_delayed_39__79_,chained_data_delayed_39__78_,
  chained_data_delayed_39__77_,chained_data_delayed_39__76_,chained_data_delayed_39__75_,
  chained_data_delayed_39__74_,chained_data_delayed_39__73_,
  chained_data_delayed_39__72_,chained_data_delayed_39__71_,chained_data_delayed_39__70_,
  chained_data_delayed_39__69_,chained_data_delayed_39__68_,chained_data_delayed_39__67_,
  chained_data_delayed_39__66_,chained_data_delayed_39__65_,chained_data_delayed_39__64_,
  chained_data_delayed_39__63_,chained_data_delayed_39__62_,
  chained_data_delayed_39__61_,chained_data_delayed_39__60_,chained_data_delayed_39__59_,
  chained_data_delayed_39__58_,chained_data_delayed_39__57_,chained_data_delayed_39__56_,
  chained_data_delayed_39__55_,chained_data_delayed_39__54_,chained_data_delayed_39__53_,
  chained_data_delayed_39__52_,chained_data_delayed_39__51_,
  chained_data_delayed_39__50_,chained_data_delayed_39__49_,chained_data_delayed_39__48_,
  chained_data_delayed_39__47_,chained_data_delayed_39__46_,chained_data_delayed_39__45_,
  chained_data_delayed_39__44_,chained_data_delayed_39__43_,chained_data_delayed_39__42_,
  chained_data_delayed_39__41_,chained_data_delayed_39__40_,
  chained_data_delayed_39__39_,chained_data_delayed_39__38_,chained_data_delayed_39__37_,
  chained_data_delayed_39__36_,chained_data_delayed_39__35_,chained_data_delayed_39__34_,
  chained_data_delayed_39__33_,chained_data_delayed_39__32_,chained_data_delayed_39__31_,
  chained_data_delayed_39__30_,chained_data_delayed_39__29_,chained_data_delayed_39__28_,
  chained_data_delayed_39__27_,chained_data_delayed_39__26_,
  chained_data_delayed_39__25_,chained_data_delayed_39__24_,chained_data_delayed_39__23_,
  chained_data_delayed_39__22_,chained_data_delayed_39__21_,chained_data_delayed_39__20_,
  chained_data_delayed_39__19_,chained_data_delayed_39__18_,chained_data_delayed_39__17_,
  chained_data_delayed_39__16_,chained_data_delayed_39__15_,
  chained_data_delayed_39__14_,chained_data_delayed_39__13_,chained_data_delayed_39__12_,
  chained_data_delayed_39__11_,chained_data_delayed_39__10_,chained_data_delayed_39__9_,
  chained_data_delayed_39__8_,chained_data_delayed_39__7_,chained_data_delayed_39__6_,
  chained_data_delayed_39__5_,chained_data_delayed_39__4_,chained_data_delayed_39__3_,
  chained_data_delayed_39__2_,chained_data_delayed_39__1_,
  chained_data_delayed_39__0_,chained_data_delayed_38__127_,chained_data_delayed_38__126_,
  chained_data_delayed_38__125_,chained_data_delayed_38__124_,chained_data_delayed_38__123_,
  chained_data_delayed_38__122_,chained_data_delayed_38__121_,
  chained_data_delayed_38__120_,chained_data_delayed_38__119_,chained_data_delayed_38__118_,
  chained_data_delayed_38__117_,chained_data_delayed_38__116_,chained_data_delayed_38__115_,
  chained_data_delayed_38__114_,chained_data_delayed_38__113_,
  chained_data_delayed_38__112_,chained_data_delayed_38__111_,chained_data_delayed_38__110_,
  chained_data_delayed_38__109_,chained_data_delayed_38__108_,chained_data_delayed_38__107_,
  chained_data_delayed_38__106_,chained_data_delayed_38__105_,
  chained_data_delayed_38__104_,chained_data_delayed_38__103_,chained_data_delayed_38__102_,
  chained_data_delayed_38__101_,chained_data_delayed_38__100_,chained_data_delayed_38__99_,
  chained_data_delayed_38__98_,chained_data_delayed_38__97_,chained_data_delayed_38__96_,
  chained_data_delayed_38__95_,chained_data_delayed_38__94_,
  chained_data_delayed_38__93_,chained_data_delayed_38__92_,chained_data_delayed_38__91_,
  chained_data_delayed_38__90_,chained_data_delayed_38__89_,chained_data_delayed_38__88_,
  chained_data_delayed_38__87_,chained_data_delayed_38__86_,chained_data_delayed_38__85_,
  chained_data_delayed_38__84_,chained_data_delayed_38__83_,
  chained_data_delayed_38__82_,chained_data_delayed_38__81_,chained_data_delayed_38__80_,
  chained_data_delayed_38__79_,chained_data_delayed_38__78_,chained_data_delayed_38__77_,
  chained_data_delayed_38__76_,chained_data_delayed_38__75_,chained_data_delayed_38__74_,
  chained_data_delayed_38__73_,chained_data_delayed_38__72_,
  chained_data_delayed_38__71_,chained_data_delayed_38__70_,chained_data_delayed_38__69_,
  chained_data_delayed_38__68_,chained_data_delayed_38__67_,chained_data_delayed_38__66_,
  chained_data_delayed_38__65_,chained_data_delayed_38__64_,chained_data_delayed_38__63_,
  chained_data_delayed_38__62_,chained_data_delayed_38__61_,
  chained_data_delayed_38__60_,chained_data_delayed_38__59_,chained_data_delayed_38__58_,
  chained_data_delayed_38__57_,chained_data_delayed_38__56_,chained_data_delayed_38__55_,
  chained_data_delayed_38__54_,chained_data_delayed_38__53_,chained_data_delayed_38__52_,
  chained_data_delayed_38__51_,chained_data_delayed_38__50_,
  chained_data_delayed_38__49_,chained_data_delayed_38__48_,chained_data_delayed_38__47_,
  chained_data_delayed_38__46_,chained_data_delayed_38__45_,chained_data_delayed_38__44_,
  chained_data_delayed_38__43_,chained_data_delayed_38__42_,chained_data_delayed_38__41_,
  chained_data_delayed_38__40_,chained_data_delayed_38__39_,chained_data_delayed_38__38_,
  chained_data_delayed_38__37_,chained_data_delayed_38__36_,
  chained_data_delayed_38__35_,chained_data_delayed_38__34_,chained_data_delayed_38__33_,
  chained_data_delayed_38__32_,chained_data_delayed_38__31_,chained_data_delayed_38__30_,
  chained_data_delayed_38__29_,chained_data_delayed_38__28_,chained_data_delayed_38__27_,
  chained_data_delayed_38__26_,chained_data_delayed_38__25_,
  chained_data_delayed_38__24_,chained_data_delayed_38__23_,chained_data_delayed_38__22_,
  chained_data_delayed_38__21_,chained_data_delayed_38__20_,chained_data_delayed_38__19_,
  chained_data_delayed_38__18_,chained_data_delayed_38__17_,chained_data_delayed_38__16_,
  chained_data_delayed_38__15_,chained_data_delayed_38__14_,
  chained_data_delayed_38__13_,chained_data_delayed_38__12_,chained_data_delayed_38__11_,
  chained_data_delayed_38__10_,chained_data_delayed_38__9_,chained_data_delayed_38__8_,
  chained_data_delayed_38__7_,chained_data_delayed_38__6_,chained_data_delayed_38__5_,
  chained_data_delayed_38__4_,chained_data_delayed_38__3_,chained_data_delayed_38__2_,
  chained_data_delayed_38__1_,chained_data_delayed_38__0_,
  chained_data_delayed_37__127_,chained_data_delayed_37__126_,chained_data_delayed_37__125_,
  chained_data_delayed_37__124_,chained_data_delayed_37__123_,chained_data_delayed_37__122_,
  chained_data_delayed_37__121_,chained_data_delayed_37__120_,
  chained_data_delayed_37__119_,chained_data_delayed_37__118_,chained_data_delayed_37__117_,
  chained_data_delayed_37__116_,chained_data_delayed_37__115_,chained_data_delayed_37__114_,
  chained_data_delayed_37__113_,chained_data_delayed_37__112_,
  chained_data_delayed_37__111_,chained_data_delayed_37__110_,chained_data_delayed_37__109_,
  chained_data_delayed_37__108_,chained_data_delayed_37__107_,chained_data_delayed_37__106_,
  chained_data_delayed_37__105_,chained_data_delayed_37__104_,
  chained_data_delayed_37__103_,chained_data_delayed_37__102_,chained_data_delayed_37__101_,
  chained_data_delayed_37__100_,chained_data_delayed_37__99_,chained_data_delayed_37__98_,
  chained_data_delayed_37__97_,chained_data_delayed_37__96_,chained_data_delayed_37__95_,
  chained_data_delayed_37__94_,chained_data_delayed_37__93_,
  chained_data_delayed_37__92_,chained_data_delayed_37__91_,chained_data_delayed_37__90_,
  chained_data_delayed_37__89_,chained_data_delayed_37__88_,chained_data_delayed_37__87_,
  chained_data_delayed_37__86_,chained_data_delayed_37__85_,chained_data_delayed_37__84_,
  chained_data_delayed_37__83_,chained_data_delayed_37__82_,
  chained_data_delayed_37__81_,chained_data_delayed_37__80_,chained_data_delayed_37__79_,
  chained_data_delayed_37__78_,chained_data_delayed_37__77_,chained_data_delayed_37__76_,
  chained_data_delayed_37__75_,chained_data_delayed_37__74_,chained_data_delayed_37__73_,
  chained_data_delayed_37__72_,chained_data_delayed_37__71_,
  chained_data_delayed_37__70_,chained_data_delayed_37__69_,chained_data_delayed_37__68_,
  chained_data_delayed_37__67_,chained_data_delayed_37__66_,chained_data_delayed_37__65_,
  chained_data_delayed_37__64_,chained_data_delayed_37__63_,chained_data_delayed_37__62_,
  chained_data_delayed_37__61_,chained_data_delayed_37__60_,
  chained_data_delayed_37__59_,chained_data_delayed_37__58_,chained_data_delayed_37__57_,
  chained_data_delayed_37__56_,chained_data_delayed_37__55_,chained_data_delayed_37__54_,
  chained_data_delayed_37__53_,chained_data_delayed_37__52_,chained_data_delayed_37__51_,
  chained_data_delayed_37__50_,chained_data_delayed_37__49_,chained_data_delayed_37__48_,
  chained_data_delayed_37__47_,chained_data_delayed_37__46_,
  chained_data_delayed_37__45_,chained_data_delayed_37__44_,chained_data_delayed_37__43_,
  chained_data_delayed_37__42_,chained_data_delayed_37__41_,chained_data_delayed_37__40_,
  chained_data_delayed_37__39_,chained_data_delayed_37__38_,chained_data_delayed_37__37_,
  chained_data_delayed_37__36_,chained_data_delayed_37__35_,
  chained_data_delayed_37__34_,chained_data_delayed_37__33_,chained_data_delayed_37__32_,
  chained_data_delayed_37__31_,chained_data_delayed_37__30_,chained_data_delayed_37__29_,
  chained_data_delayed_37__28_,chained_data_delayed_37__27_,chained_data_delayed_37__26_,
  chained_data_delayed_37__25_,chained_data_delayed_37__24_,
  chained_data_delayed_37__23_,chained_data_delayed_37__22_,chained_data_delayed_37__21_,
  chained_data_delayed_37__20_,chained_data_delayed_37__19_,chained_data_delayed_37__18_,
  chained_data_delayed_37__17_,chained_data_delayed_37__16_,chained_data_delayed_37__15_,
  chained_data_delayed_37__14_,chained_data_delayed_37__13_,
  chained_data_delayed_37__12_,chained_data_delayed_37__11_,chained_data_delayed_37__10_,
  chained_data_delayed_37__9_,chained_data_delayed_37__8_,chained_data_delayed_37__7_,
  chained_data_delayed_37__6_,chained_data_delayed_37__5_,chained_data_delayed_37__4_,
  chained_data_delayed_37__3_,chained_data_delayed_37__2_,chained_data_delayed_37__1_,
  chained_data_delayed_37__0_,chained_data_delayed_44__127_,
  chained_data_delayed_44__126_,chained_data_delayed_44__125_,chained_data_delayed_44__124_,
  chained_data_delayed_44__123_,chained_data_delayed_44__122_,chained_data_delayed_44__121_,
  chained_data_delayed_44__120_,chained_data_delayed_44__119_,
  chained_data_delayed_44__118_,chained_data_delayed_44__117_,chained_data_delayed_44__116_,
  chained_data_delayed_44__115_,chained_data_delayed_44__114_,chained_data_delayed_44__113_,
  chained_data_delayed_44__112_,chained_data_delayed_44__111_,
  chained_data_delayed_44__110_,chained_data_delayed_44__109_,chained_data_delayed_44__108_,
  chained_data_delayed_44__107_,chained_data_delayed_44__106_,chained_data_delayed_44__105_,
  chained_data_delayed_44__104_,chained_data_delayed_44__103_,
  chained_data_delayed_44__102_,chained_data_delayed_44__101_,chained_data_delayed_44__100_,
  chained_data_delayed_44__99_,chained_data_delayed_44__98_,chained_data_delayed_44__97_,
  chained_data_delayed_44__96_,chained_data_delayed_44__95_,chained_data_delayed_44__94_,
  chained_data_delayed_44__93_,chained_data_delayed_44__92_,
  chained_data_delayed_44__91_,chained_data_delayed_44__90_,chained_data_delayed_44__89_,
  chained_data_delayed_44__88_,chained_data_delayed_44__87_,chained_data_delayed_44__86_,
  chained_data_delayed_44__85_,chained_data_delayed_44__84_,chained_data_delayed_44__83_,
  chained_data_delayed_44__82_,chained_data_delayed_44__81_,
  chained_data_delayed_44__80_,chained_data_delayed_44__79_,chained_data_delayed_44__78_,
  chained_data_delayed_44__77_,chained_data_delayed_44__76_,chained_data_delayed_44__75_,
  chained_data_delayed_44__74_,chained_data_delayed_44__73_,chained_data_delayed_44__72_,
  chained_data_delayed_44__71_,chained_data_delayed_44__70_,
  chained_data_delayed_44__69_,chained_data_delayed_44__68_,chained_data_delayed_44__67_,
  chained_data_delayed_44__66_,chained_data_delayed_44__65_,chained_data_delayed_44__64_,
  chained_data_delayed_44__63_,chained_data_delayed_44__62_,chained_data_delayed_44__61_,
  chained_data_delayed_44__60_,chained_data_delayed_44__59_,chained_data_delayed_44__58_,
  chained_data_delayed_44__57_,chained_data_delayed_44__56_,
  chained_data_delayed_44__55_,chained_data_delayed_44__54_,chained_data_delayed_44__53_,
  chained_data_delayed_44__52_,chained_data_delayed_44__51_,chained_data_delayed_44__50_,
  chained_data_delayed_44__49_,chained_data_delayed_44__48_,chained_data_delayed_44__47_,
  chained_data_delayed_44__46_,chained_data_delayed_44__45_,
  chained_data_delayed_44__44_,chained_data_delayed_44__43_,chained_data_delayed_44__42_,
  chained_data_delayed_44__41_,chained_data_delayed_44__40_,chained_data_delayed_44__39_,
  chained_data_delayed_44__38_,chained_data_delayed_44__37_,chained_data_delayed_44__36_,
  chained_data_delayed_44__35_,chained_data_delayed_44__34_,
  chained_data_delayed_44__33_,chained_data_delayed_44__32_,chained_data_delayed_44__31_,
  chained_data_delayed_44__30_,chained_data_delayed_44__29_,chained_data_delayed_44__28_,
  chained_data_delayed_44__27_,chained_data_delayed_44__26_,chained_data_delayed_44__25_,
  chained_data_delayed_44__24_,chained_data_delayed_44__23_,
  chained_data_delayed_44__22_,chained_data_delayed_44__21_,chained_data_delayed_44__20_,
  chained_data_delayed_44__19_,chained_data_delayed_44__18_,chained_data_delayed_44__17_,
  chained_data_delayed_44__16_,chained_data_delayed_44__15_,chained_data_delayed_44__14_,
  chained_data_delayed_44__13_,chained_data_delayed_44__12_,
  chained_data_delayed_44__11_,chained_data_delayed_44__10_,chained_data_delayed_44__9_,
  chained_data_delayed_44__8_,chained_data_delayed_44__7_,chained_data_delayed_44__6_,
  chained_data_delayed_44__5_,chained_data_delayed_44__4_,chained_data_delayed_44__3_,
  chained_data_delayed_44__2_,chained_data_delayed_44__1_,chained_data_delayed_44__0_,
  chained_data_delayed_43__127_,chained_data_delayed_43__126_,
  chained_data_delayed_43__125_,chained_data_delayed_43__124_,chained_data_delayed_43__123_,
  chained_data_delayed_43__122_,chained_data_delayed_43__121_,chained_data_delayed_43__120_,
  chained_data_delayed_43__119_,chained_data_delayed_43__118_,
  chained_data_delayed_43__117_,chained_data_delayed_43__116_,chained_data_delayed_43__115_,
  chained_data_delayed_43__114_,chained_data_delayed_43__113_,chained_data_delayed_43__112_,
  chained_data_delayed_43__111_,chained_data_delayed_43__110_,
  chained_data_delayed_43__109_,chained_data_delayed_43__108_,chained_data_delayed_43__107_,
  chained_data_delayed_43__106_,chained_data_delayed_43__105_,chained_data_delayed_43__104_,
  chained_data_delayed_43__103_,chained_data_delayed_43__102_,
  chained_data_delayed_43__101_,chained_data_delayed_43__100_,chained_data_delayed_43__99_,
  chained_data_delayed_43__98_,chained_data_delayed_43__97_,chained_data_delayed_43__96_,
  chained_data_delayed_43__95_,chained_data_delayed_43__94_,chained_data_delayed_43__93_,
  chained_data_delayed_43__92_,chained_data_delayed_43__91_,
  chained_data_delayed_43__90_,chained_data_delayed_43__89_,chained_data_delayed_43__88_,
  chained_data_delayed_43__87_,chained_data_delayed_43__86_,chained_data_delayed_43__85_,
  chained_data_delayed_43__84_,chained_data_delayed_43__83_,chained_data_delayed_43__82_,
  chained_data_delayed_43__81_,chained_data_delayed_43__80_,
  chained_data_delayed_43__79_,chained_data_delayed_43__78_,chained_data_delayed_43__77_,
  chained_data_delayed_43__76_,chained_data_delayed_43__75_,chained_data_delayed_43__74_,
  chained_data_delayed_43__73_,chained_data_delayed_43__72_,chained_data_delayed_43__71_,
  chained_data_delayed_43__70_,chained_data_delayed_43__69_,chained_data_delayed_43__68_,
  chained_data_delayed_43__67_,chained_data_delayed_43__66_,
  chained_data_delayed_43__65_,chained_data_delayed_43__64_,chained_data_delayed_43__63_,
  chained_data_delayed_43__62_,chained_data_delayed_43__61_,chained_data_delayed_43__60_,
  chained_data_delayed_43__59_,chained_data_delayed_43__58_,chained_data_delayed_43__57_,
  chained_data_delayed_43__56_,chained_data_delayed_43__55_,
  chained_data_delayed_43__54_,chained_data_delayed_43__53_,chained_data_delayed_43__52_,
  chained_data_delayed_43__51_,chained_data_delayed_43__50_,chained_data_delayed_43__49_,
  chained_data_delayed_43__48_,chained_data_delayed_43__47_,chained_data_delayed_43__46_,
  chained_data_delayed_43__45_,chained_data_delayed_43__44_,
  chained_data_delayed_43__43_,chained_data_delayed_43__42_,chained_data_delayed_43__41_,
  chained_data_delayed_43__40_,chained_data_delayed_43__39_,chained_data_delayed_43__38_,
  chained_data_delayed_43__37_,chained_data_delayed_43__36_,chained_data_delayed_43__35_,
  chained_data_delayed_43__34_,chained_data_delayed_43__33_,
  chained_data_delayed_43__32_,chained_data_delayed_43__31_,chained_data_delayed_43__30_,
  chained_data_delayed_43__29_,chained_data_delayed_43__28_,chained_data_delayed_43__27_,
  chained_data_delayed_43__26_,chained_data_delayed_43__25_,chained_data_delayed_43__24_,
  chained_data_delayed_43__23_,chained_data_delayed_43__22_,
  chained_data_delayed_43__21_,chained_data_delayed_43__20_,chained_data_delayed_43__19_,
  chained_data_delayed_43__18_,chained_data_delayed_43__17_,chained_data_delayed_43__16_,
  chained_data_delayed_43__15_,chained_data_delayed_43__14_,chained_data_delayed_43__13_,
  chained_data_delayed_43__12_,chained_data_delayed_43__11_,
  chained_data_delayed_43__10_,chained_data_delayed_43__9_,chained_data_delayed_43__8_,
  chained_data_delayed_43__7_,chained_data_delayed_43__6_,chained_data_delayed_43__5_,
  chained_data_delayed_43__4_,chained_data_delayed_43__3_,chained_data_delayed_43__2_,
  chained_data_delayed_43__1_,chained_data_delayed_43__0_,chained_data_delayed_42__127_,
  chained_data_delayed_42__126_,chained_data_delayed_42__125_,
  chained_data_delayed_42__124_,chained_data_delayed_42__123_,chained_data_delayed_42__122_,
  chained_data_delayed_42__121_,chained_data_delayed_42__120_,chained_data_delayed_42__119_,
  chained_data_delayed_42__118_,chained_data_delayed_42__117_,
  chained_data_delayed_42__116_,chained_data_delayed_42__115_,chained_data_delayed_42__114_,
  chained_data_delayed_42__113_,chained_data_delayed_42__112_,chained_data_delayed_42__111_,
  chained_data_delayed_42__110_,chained_data_delayed_42__109_,
  chained_data_delayed_42__108_,chained_data_delayed_42__107_,chained_data_delayed_42__106_,
  chained_data_delayed_42__105_,chained_data_delayed_42__104_,chained_data_delayed_42__103_,
  chained_data_delayed_42__102_,chained_data_delayed_42__101_,
  chained_data_delayed_42__100_,chained_data_delayed_42__99_,chained_data_delayed_42__98_,
  chained_data_delayed_42__97_,chained_data_delayed_42__96_,chained_data_delayed_42__95_,
  chained_data_delayed_42__94_,chained_data_delayed_42__93_,chained_data_delayed_42__92_,
  chained_data_delayed_42__91_,chained_data_delayed_42__90_,
  chained_data_delayed_42__89_,chained_data_delayed_42__88_,chained_data_delayed_42__87_,
  chained_data_delayed_42__86_,chained_data_delayed_42__85_,chained_data_delayed_42__84_,
  chained_data_delayed_42__83_,chained_data_delayed_42__82_,chained_data_delayed_42__81_,
  chained_data_delayed_42__80_,chained_data_delayed_42__79_,chained_data_delayed_42__78_,
  chained_data_delayed_42__77_,chained_data_delayed_42__76_,
  chained_data_delayed_42__75_,chained_data_delayed_42__74_,chained_data_delayed_42__73_,
  chained_data_delayed_42__72_,chained_data_delayed_42__71_,chained_data_delayed_42__70_,
  chained_data_delayed_42__69_,chained_data_delayed_42__68_,chained_data_delayed_42__67_,
  chained_data_delayed_42__66_,chained_data_delayed_42__65_,
  chained_data_delayed_42__64_,chained_data_delayed_42__63_,chained_data_delayed_42__62_,
  chained_data_delayed_42__61_,chained_data_delayed_42__60_,chained_data_delayed_42__59_,
  chained_data_delayed_42__58_,chained_data_delayed_42__57_,chained_data_delayed_42__56_,
  chained_data_delayed_42__55_,chained_data_delayed_42__54_,
  chained_data_delayed_42__53_,chained_data_delayed_42__52_,chained_data_delayed_42__51_,
  chained_data_delayed_42__50_,chained_data_delayed_42__49_,chained_data_delayed_42__48_,
  chained_data_delayed_42__47_,chained_data_delayed_42__46_,chained_data_delayed_42__45_,
  chained_data_delayed_42__44_,chained_data_delayed_42__43_,
  chained_data_delayed_42__42_,chained_data_delayed_42__41_,chained_data_delayed_42__40_,
  chained_data_delayed_42__39_,chained_data_delayed_42__38_,chained_data_delayed_42__37_,
  chained_data_delayed_42__36_,chained_data_delayed_42__35_,chained_data_delayed_42__34_,
  chained_data_delayed_42__33_,chained_data_delayed_42__32_,
  chained_data_delayed_42__31_,chained_data_delayed_42__30_,chained_data_delayed_42__29_,
  chained_data_delayed_42__28_,chained_data_delayed_42__27_,chained_data_delayed_42__26_,
  chained_data_delayed_42__25_,chained_data_delayed_42__24_,chained_data_delayed_42__23_,
  chained_data_delayed_42__22_,chained_data_delayed_42__21_,
  chained_data_delayed_42__20_,chained_data_delayed_42__19_,chained_data_delayed_42__18_,
  chained_data_delayed_42__17_,chained_data_delayed_42__16_,chained_data_delayed_42__15_,
  chained_data_delayed_42__14_,chained_data_delayed_42__13_,chained_data_delayed_42__12_,
  chained_data_delayed_42__11_,chained_data_delayed_42__10_,chained_data_delayed_42__9_,
  chained_data_delayed_42__8_,chained_data_delayed_42__7_,
  chained_data_delayed_42__6_,chained_data_delayed_42__5_,chained_data_delayed_42__4_,
  chained_data_delayed_42__3_,chained_data_delayed_42__2_,chained_data_delayed_42__1_,
  chained_data_delayed_42__0_,chained_data_delayed_41__127_,chained_data_delayed_41__126_,
  chained_data_delayed_41__125_,chained_data_delayed_41__124_,
  chained_data_delayed_41__123_,chained_data_delayed_41__122_,chained_data_delayed_41__121_,
  chained_data_delayed_41__120_,chained_data_delayed_41__119_,chained_data_delayed_41__118_,
  chained_data_delayed_41__117_,chained_data_delayed_41__116_,
  chained_data_delayed_41__115_,chained_data_delayed_41__114_,chained_data_delayed_41__113_,
  chained_data_delayed_41__112_,chained_data_delayed_41__111_,chained_data_delayed_41__110_,
  chained_data_delayed_41__109_,chained_data_delayed_41__108_,
  chained_data_delayed_41__107_,chained_data_delayed_41__106_,chained_data_delayed_41__105_,
  chained_data_delayed_41__104_,chained_data_delayed_41__103_,chained_data_delayed_41__102_,
  chained_data_delayed_41__101_,chained_data_delayed_41__100_,
  chained_data_delayed_41__99_,chained_data_delayed_41__98_,chained_data_delayed_41__97_,
  chained_data_delayed_41__96_,chained_data_delayed_41__95_,chained_data_delayed_41__94_,
  chained_data_delayed_41__93_,chained_data_delayed_41__92_,chained_data_delayed_41__91_,
  chained_data_delayed_41__90_,chained_data_delayed_41__89_,chained_data_delayed_41__88_,
  chained_data_delayed_41__87_,chained_data_delayed_41__86_,
  chained_data_delayed_41__85_,chained_data_delayed_41__84_,chained_data_delayed_41__83_,
  chained_data_delayed_41__82_,chained_data_delayed_41__81_,chained_data_delayed_41__80_,
  chained_data_delayed_41__79_,chained_data_delayed_41__78_,chained_data_delayed_41__77_,
  chained_data_delayed_41__76_,chained_data_delayed_41__75_,
  chained_data_delayed_41__74_,chained_data_delayed_41__73_,chained_data_delayed_41__72_,
  chained_data_delayed_41__71_,chained_data_delayed_41__70_,chained_data_delayed_41__69_,
  chained_data_delayed_41__68_,chained_data_delayed_41__67_,chained_data_delayed_41__66_,
  chained_data_delayed_41__65_,chained_data_delayed_41__64_,
  chained_data_delayed_41__63_,chained_data_delayed_41__62_,chained_data_delayed_41__61_,
  chained_data_delayed_41__60_,chained_data_delayed_41__59_,chained_data_delayed_41__58_,
  chained_data_delayed_41__57_,chained_data_delayed_41__56_,chained_data_delayed_41__55_,
  chained_data_delayed_41__54_,chained_data_delayed_41__53_,
  chained_data_delayed_41__52_,chained_data_delayed_41__51_,chained_data_delayed_41__50_,
  chained_data_delayed_41__49_,chained_data_delayed_41__48_,chained_data_delayed_41__47_,
  chained_data_delayed_41__46_,chained_data_delayed_41__45_,chained_data_delayed_41__44_,
  chained_data_delayed_41__43_,chained_data_delayed_41__42_,
  chained_data_delayed_41__41_,chained_data_delayed_41__40_,chained_data_delayed_41__39_,
  chained_data_delayed_41__38_,chained_data_delayed_41__37_,chained_data_delayed_41__36_,
  chained_data_delayed_41__35_,chained_data_delayed_41__34_,chained_data_delayed_41__33_,
  chained_data_delayed_41__32_,chained_data_delayed_41__31_,
  chained_data_delayed_41__30_,chained_data_delayed_41__29_,chained_data_delayed_41__28_,
  chained_data_delayed_41__27_,chained_data_delayed_41__26_,chained_data_delayed_41__25_,
  chained_data_delayed_41__24_,chained_data_delayed_41__23_,chained_data_delayed_41__22_,
  chained_data_delayed_41__21_,chained_data_delayed_41__20_,
  chained_data_delayed_41__19_,chained_data_delayed_41__18_,chained_data_delayed_41__17_,
  chained_data_delayed_41__16_,chained_data_delayed_41__15_,chained_data_delayed_41__14_,
  chained_data_delayed_41__13_,chained_data_delayed_41__12_,chained_data_delayed_41__11_,
  chained_data_delayed_41__10_,chained_data_delayed_41__9_,chained_data_delayed_41__8_,
  chained_data_delayed_41__7_,chained_data_delayed_41__6_,
  chained_data_delayed_41__5_,chained_data_delayed_41__4_,chained_data_delayed_41__3_,
  chained_data_delayed_41__2_,chained_data_delayed_41__1_,chained_data_delayed_41__0_,
  chained_data_delayed_48__127_,chained_data_delayed_48__126_,chained_data_delayed_48__125_,
  chained_data_delayed_48__124_,chained_data_delayed_48__123_,
  chained_data_delayed_48__122_,chained_data_delayed_48__121_,chained_data_delayed_48__120_,
  chained_data_delayed_48__119_,chained_data_delayed_48__118_,chained_data_delayed_48__117_,
  chained_data_delayed_48__116_,chained_data_delayed_48__115_,
  chained_data_delayed_48__114_,chained_data_delayed_48__113_,chained_data_delayed_48__112_,
  chained_data_delayed_48__111_,chained_data_delayed_48__110_,chained_data_delayed_48__109_,
  chained_data_delayed_48__108_,chained_data_delayed_48__107_,
  chained_data_delayed_48__106_,chained_data_delayed_48__105_,chained_data_delayed_48__104_,
  chained_data_delayed_48__103_,chained_data_delayed_48__102_,chained_data_delayed_48__101_,
  chained_data_delayed_48__100_,chained_data_delayed_48__99_,chained_data_delayed_48__98_,
  chained_data_delayed_48__97_,chained_data_delayed_48__96_,
  chained_data_delayed_48__95_,chained_data_delayed_48__94_,chained_data_delayed_48__93_,
  chained_data_delayed_48__92_,chained_data_delayed_48__91_,chained_data_delayed_48__90_,
  chained_data_delayed_48__89_,chained_data_delayed_48__88_,chained_data_delayed_48__87_,
  chained_data_delayed_48__86_,chained_data_delayed_48__85_,
  chained_data_delayed_48__84_,chained_data_delayed_48__83_,chained_data_delayed_48__82_,
  chained_data_delayed_48__81_,chained_data_delayed_48__80_,chained_data_delayed_48__79_,
  chained_data_delayed_48__78_,chained_data_delayed_48__77_,chained_data_delayed_48__76_,
  chained_data_delayed_48__75_,chained_data_delayed_48__74_,
  chained_data_delayed_48__73_,chained_data_delayed_48__72_,chained_data_delayed_48__71_,
  chained_data_delayed_48__70_,chained_data_delayed_48__69_,chained_data_delayed_48__68_,
  chained_data_delayed_48__67_,chained_data_delayed_48__66_,chained_data_delayed_48__65_,
  chained_data_delayed_48__64_,chained_data_delayed_48__63_,
  chained_data_delayed_48__62_,chained_data_delayed_48__61_,chained_data_delayed_48__60_,
  chained_data_delayed_48__59_,chained_data_delayed_48__58_,chained_data_delayed_48__57_,
  chained_data_delayed_48__56_,chained_data_delayed_48__55_,chained_data_delayed_48__54_,
  chained_data_delayed_48__53_,chained_data_delayed_48__52_,
  chained_data_delayed_48__51_,chained_data_delayed_48__50_,chained_data_delayed_48__49_,
  chained_data_delayed_48__48_,chained_data_delayed_48__47_,chained_data_delayed_48__46_,
  chained_data_delayed_48__45_,chained_data_delayed_48__44_,chained_data_delayed_48__43_,
  chained_data_delayed_48__42_,chained_data_delayed_48__41_,
  chained_data_delayed_48__40_,chained_data_delayed_48__39_,chained_data_delayed_48__38_,
  chained_data_delayed_48__37_,chained_data_delayed_48__36_,chained_data_delayed_48__35_,
  chained_data_delayed_48__34_,chained_data_delayed_48__33_,chained_data_delayed_48__32_,
  chained_data_delayed_48__31_,chained_data_delayed_48__30_,
  chained_data_delayed_48__29_,chained_data_delayed_48__28_,chained_data_delayed_48__27_,
  chained_data_delayed_48__26_,chained_data_delayed_48__25_,chained_data_delayed_48__24_,
  chained_data_delayed_48__23_,chained_data_delayed_48__22_,chained_data_delayed_48__21_,
  chained_data_delayed_48__20_,chained_data_delayed_48__19_,chained_data_delayed_48__18_,
  chained_data_delayed_48__17_,chained_data_delayed_48__16_,
  chained_data_delayed_48__15_,chained_data_delayed_48__14_,chained_data_delayed_48__13_,
  chained_data_delayed_48__12_,chained_data_delayed_48__11_,chained_data_delayed_48__10_,
  chained_data_delayed_48__9_,chained_data_delayed_48__8_,chained_data_delayed_48__7_,
  chained_data_delayed_48__6_,chained_data_delayed_48__5_,chained_data_delayed_48__4_,
  chained_data_delayed_48__3_,chained_data_delayed_48__2_,
  chained_data_delayed_48__1_,chained_data_delayed_48__0_,chained_data_delayed_47__127_,
  chained_data_delayed_47__126_,chained_data_delayed_47__125_,chained_data_delayed_47__124_,
  chained_data_delayed_47__123_,chained_data_delayed_47__122_,
  chained_data_delayed_47__121_,chained_data_delayed_47__120_,chained_data_delayed_47__119_,
  chained_data_delayed_47__118_,chained_data_delayed_47__117_,chained_data_delayed_47__116_,
  chained_data_delayed_47__115_,chained_data_delayed_47__114_,
  chained_data_delayed_47__113_,chained_data_delayed_47__112_,chained_data_delayed_47__111_,
  chained_data_delayed_47__110_,chained_data_delayed_47__109_,chained_data_delayed_47__108_,
  chained_data_delayed_47__107_,chained_data_delayed_47__106_,
  chained_data_delayed_47__105_,chained_data_delayed_47__104_,chained_data_delayed_47__103_,
  chained_data_delayed_47__102_,chained_data_delayed_47__101_,chained_data_delayed_47__100_,
  chained_data_delayed_47__99_,chained_data_delayed_47__98_,chained_data_delayed_47__97_,
  chained_data_delayed_47__96_,chained_data_delayed_47__95_,
  chained_data_delayed_47__94_,chained_data_delayed_47__93_,chained_data_delayed_47__92_,
  chained_data_delayed_47__91_,chained_data_delayed_47__90_,chained_data_delayed_47__89_,
  chained_data_delayed_47__88_,chained_data_delayed_47__87_,chained_data_delayed_47__86_,
  chained_data_delayed_47__85_,chained_data_delayed_47__84_,
  chained_data_delayed_47__83_,chained_data_delayed_47__82_,chained_data_delayed_47__81_,
  chained_data_delayed_47__80_,chained_data_delayed_47__79_,chained_data_delayed_47__78_,
  chained_data_delayed_47__77_,chained_data_delayed_47__76_,chained_data_delayed_47__75_,
  chained_data_delayed_47__74_,chained_data_delayed_47__73_,
  chained_data_delayed_47__72_,chained_data_delayed_47__71_,chained_data_delayed_47__70_,
  chained_data_delayed_47__69_,chained_data_delayed_47__68_,chained_data_delayed_47__67_,
  chained_data_delayed_47__66_,chained_data_delayed_47__65_,chained_data_delayed_47__64_,
  chained_data_delayed_47__63_,chained_data_delayed_47__62_,
  chained_data_delayed_47__61_,chained_data_delayed_47__60_,chained_data_delayed_47__59_,
  chained_data_delayed_47__58_,chained_data_delayed_47__57_,chained_data_delayed_47__56_,
  chained_data_delayed_47__55_,chained_data_delayed_47__54_,chained_data_delayed_47__53_,
  chained_data_delayed_47__52_,chained_data_delayed_47__51_,
  chained_data_delayed_47__50_,chained_data_delayed_47__49_,chained_data_delayed_47__48_,
  chained_data_delayed_47__47_,chained_data_delayed_47__46_,chained_data_delayed_47__45_,
  chained_data_delayed_47__44_,chained_data_delayed_47__43_,chained_data_delayed_47__42_,
  chained_data_delayed_47__41_,chained_data_delayed_47__40_,
  chained_data_delayed_47__39_,chained_data_delayed_47__38_,chained_data_delayed_47__37_,
  chained_data_delayed_47__36_,chained_data_delayed_47__35_,chained_data_delayed_47__34_,
  chained_data_delayed_47__33_,chained_data_delayed_47__32_,chained_data_delayed_47__31_,
  chained_data_delayed_47__30_,chained_data_delayed_47__29_,chained_data_delayed_47__28_,
  chained_data_delayed_47__27_,chained_data_delayed_47__26_,
  chained_data_delayed_47__25_,chained_data_delayed_47__24_,chained_data_delayed_47__23_,
  chained_data_delayed_47__22_,chained_data_delayed_47__21_,chained_data_delayed_47__20_,
  chained_data_delayed_47__19_,chained_data_delayed_47__18_,chained_data_delayed_47__17_,
  chained_data_delayed_47__16_,chained_data_delayed_47__15_,
  chained_data_delayed_47__14_,chained_data_delayed_47__13_,chained_data_delayed_47__12_,
  chained_data_delayed_47__11_,chained_data_delayed_47__10_,chained_data_delayed_47__9_,
  chained_data_delayed_47__8_,chained_data_delayed_47__7_,chained_data_delayed_47__6_,
  chained_data_delayed_47__5_,chained_data_delayed_47__4_,chained_data_delayed_47__3_,
  chained_data_delayed_47__2_,chained_data_delayed_47__1_,
  chained_data_delayed_47__0_,chained_data_delayed_46__127_,chained_data_delayed_46__126_,
  chained_data_delayed_46__125_,chained_data_delayed_46__124_,chained_data_delayed_46__123_,
  chained_data_delayed_46__122_,chained_data_delayed_46__121_,
  chained_data_delayed_46__120_,chained_data_delayed_46__119_,chained_data_delayed_46__118_,
  chained_data_delayed_46__117_,chained_data_delayed_46__116_,chained_data_delayed_46__115_,
  chained_data_delayed_46__114_,chained_data_delayed_46__113_,
  chained_data_delayed_46__112_,chained_data_delayed_46__111_,chained_data_delayed_46__110_,
  chained_data_delayed_46__109_,chained_data_delayed_46__108_,chained_data_delayed_46__107_,
  chained_data_delayed_46__106_,chained_data_delayed_46__105_,
  chained_data_delayed_46__104_,chained_data_delayed_46__103_,chained_data_delayed_46__102_,
  chained_data_delayed_46__101_,chained_data_delayed_46__100_,chained_data_delayed_46__99_,
  chained_data_delayed_46__98_,chained_data_delayed_46__97_,chained_data_delayed_46__96_,
  chained_data_delayed_46__95_,chained_data_delayed_46__94_,
  chained_data_delayed_46__93_,chained_data_delayed_46__92_,chained_data_delayed_46__91_,
  chained_data_delayed_46__90_,chained_data_delayed_46__89_,chained_data_delayed_46__88_,
  chained_data_delayed_46__87_,chained_data_delayed_46__86_,chained_data_delayed_46__85_,
  chained_data_delayed_46__84_,chained_data_delayed_46__83_,
  chained_data_delayed_46__82_,chained_data_delayed_46__81_,chained_data_delayed_46__80_,
  chained_data_delayed_46__79_,chained_data_delayed_46__78_,chained_data_delayed_46__77_,
  chained_data_delayed_46__76_,chained_data_delayed_46__75_,chained_data_delayed_46__74_,
  chained_data_delayed_46__73_,chained_data_delayed_46__72_,
  chained_data_delayed_46__71_,chained_data_delayed_46__70_,chained_data_delayed_46__69_,
  chained_data_delayed_46__68_,chained_data_delayed_46__67_,chained_data_delayed_46__66_,
  chained_data_delayed_46__65_,chained_data_delayed_46__64_,chained_data_delayed_46__63_,
  chained_data_delayed_46__62_,chained_data_delayed_46__61_,
  chained_data_delayed_46__60_,chained_data_delayed_46__59_,chained_data_delayed_46__58_,
  chained_data_delayed_46__57_,chained_data_delayed_46__56_,chained_data_delayed_46__55_,
  chained_data_delayed_46__54_,chained_data_delayed_46__53_,chained_data_delayed_46__52_,
  chained_data_delayed_46__51_,chained_data_delayed_46__50_,
  chained_data_delayed_46__49_,chained_data_delayed_46__48_,chained_data_delayed_46__47_,
  chained_data_delayed_46__46_,chained_data_delayed_46__45_,chained_data_delayed_46__44_,
  chained_data_delayed_46__43_,chained_data_delayed_46__42_,chained_data_delayed_46__41_,
  chained_data_delayed_46__40_,chained_data_delayed_46__39_,chained_data_delayed_46__38_,
  chained_data_delayed_46__37_,chained_data_delayed_46__36_,
  chained_data_delayed_46__35_,chained_data_delayed_46__34_,chained_data_delayed_46__33_,
  chained_data_delayed_46__32_,chained_data_delayed_46__31_,chained_data_delayed_46__30_,
  chained_data_delayed_46__29_,chained_data_delayed_46__28_,chained_data_delayed_46__27_,
  chained_data_delayed_46__26_,chained_data_delayed_46__25_,
  chained_data_delayed_46__24_,chained_data_delayed_46__23_,chained_data_delayed_46__22_,
  chained_data_delayed_46__21_,chained_data_delayed_46__20_,chained_data_delayed_46__19_,
  chained_data_delayed_46__18_,chained_data_delayed_46__17_,chained_data_delayed_46__16_,
  chained_data_delayed_46__15_,chained_data_delayed_46__14_,
  chained_data_delayed_46__13_,chained_data_delayed_46__12_,chained_data_delayed_46__11_,
  chained_data_delayed_46__10_,chained_data_delayed_46__9_,chained_data_delayed_46__8_,
  chained_data_delayed_46__7_,chained_data_delayed_46__6_,chained_data_delayed_46__5_,
  chained_data_delayed_46__4_,chained_data_delayed_46__3_,chained_data_delayed_46__2_,
  chained_data_delayed_46__1_,chained_data_delayed_46__0_,
  chained_data_delayed_45__127_,chained_data_delayed_45__126_,chained_data_delayed_45__125_,
  chained_data_delayed_45__124_,chained_data_delayed_45__123_,chained_data_delayed_45__122_,
  chained_data_delayed_45__121_,chained_data_delayed_45__120_,
  chained_data_delayed_45__119_,chained_data_delayed_45__118_,chained_data_delayed_45__117_,
  chained_data_delayed_45__116_,chained_data_delayed_45__115_,chained_data_delayed_45__114_,
  chained_data_delayed_45__113_,chained_data_delayed_45__112_,
  chained_data_delayed_45__111_,chained_data_delayed_45__110_,chained_data_delayed_45__109_,
  chained_data_delayed_45__108_,chained_data_delayed_45__107_,chained_data_delayed_45__106_,
  chained_data_delayed_45__105_,chained_data_delayed_45__104_,
  chained_data_delayed_45__103_,chained_data_delayed_45__102_,chained_data_delayed_45__101_,
  chained_data_delayed_45__100_,chained_data_delayed_45__99_,chained_data_delayed_45__98_,
  chained_data_delayed_45__97_,chained_data_delayed_45__96_,chained_data_delayed_45__95_,
  chained_data_delayed_45__94_,chained_data_delayed_45__93_,
  chained_data_delayed_45__92_,chained_data_delayed_45__91_,chained_data_delayed_45__90_,
  chained_data_delayed_45__89_,chained_data_delayed_45__88_,chained_data_delayed_45__87_,
  chained_data_delayed_45__86_,chained_data_delayed_45__85_,chained_data_delayed_45__84_,
  chained_data_delayed_45__83_,chained_data_delayed_45__82_,
  chained_data_delayed_45__81_,chained_data_delayed_45__80_,chained_data_delayed_45__79_,
  chained_data_delayed_45__78_,chained_data_delayed_45__77_,chained_data_delayed_45__76_,
  chained_data_delayed_45__75_,chained_data_delayed_45__74_,chained_data_delayed_45__73_,
  chained_data_delayed_45__72_,chained_data_delayed_45__71_,
  chained_data_delayed_45__70_,chained_data_delayed_45__69_,chained_data_delayed_45__68_,
  chained_data_delayed_45__67_,chained_data_delayed_45__66_,chained_data_delayed_45__65_,
  chained_data_delayed_45__64_,chained_data_delayed_45__63_,chained_data_delayed_45__62_,
  chained_data_delayed_45__61_,chained_data_delayed_45__60_,
  chained_data_delayed_45__59_,chained_data_delayed_45__58_,chained_data_delayed_45__57_,
  chained_data_delayed_45__56_,chained_data_delayed_45__55_,chained_data_delayed_45__54_,
  chained_data_delayed_45__53_,chained_data_delayed_45__52_,chained_data_delayed_45__51_,
  chained_data_delayed_45__50_,chained_data_delayed_45__49_,chained_data_delayed_45__48_,
  chained_data_delayed_45__47_,chained_data_delayed_45__46_,
  chained_data_delayed_45__45_,chained_data_delayed_45__44_,chained_data_delayed_45__43_,
  chained_data_delayed_45__42_,chained_data_delayed_45__41_,chained_data_delayed_45__40_,
  chained_data_delayed_45__39_,chained_data_delayed_45__38_,chained_data_delayed_45__37_,
  chained_data_delayed_45__36_,chained_data_delayed_45__35_,
  chained_data_delayed_45__34_,chained_data_delayed_45__33_,chained_data_delayed_45__32_,
  chained_data_delayed_45__31_,chained_data_delayed_45__30_,chained_data_delayed_45__29_,
  chained_data_delayed_45__28_,chained_data_delayed_45__27_,chained_data_delayed_45__26_,
  chained_data_delayed_45__25_,chained_data_delayed_45__24_,
  chained_data_delayed_45__23_,chained_data_delayed_45__22_,chained_data_delayed_45__21_,
  chained_data_delayed_45__20_,chained_data_delayed_45__19_,chained_data_delayed_45__18_,
  chained_data_delayed_45__17_,chained_data_delayed_45__16_,chained_data_delayed_45__15_,
  chained_data_delayed_45__14_,chained_data_delayed_45__13_,
  chained_data_delayed_45__12_,chained_data_delayed_45__11_,chained_data_delayed_45__10_,
  chained_data_delayed_45__9_,chained_data_delayed_45__8_,chained_data_delayed_45__7_,
  chained_data_delayed_45__6_,chained_data_delayed_45__5_,chained_data_delayed_45__4_,
  chained_data_delayed_45__3_,chained_data_delayed_45__2_,chained_data_delayed_45__1_,
  chained_data_delayed_45__0_,chained_data_delayed_52__127_,
  chained_data_delayed_52__126_,chained_data_delayed_52__125_,chained_data_delayed_52__124_,
  chained_data_delayed_52__123_,chained_data_delayed_52__122_,chained_data_delayed_52__121_,
  chained_data_delayed_52__120_,chained_data_delayed_52__119_,
  chained_data_delayed_52__118_,chained_data_delayed_52__117_,chained_data_delayed_52__116_,
  chained_data_delayed_52__115_,chained_data_delayed_52__114_,chained_data_delayed_52__113_,
  chained_data_delayed_52__112_,chained_data_delayed_52__111_,
  chained_data_delayed_52__110_,chained_data_delayed_52__109_,chained_data_delayed_52__108_,
  chained_data_delayed_52__107_,chained_data_delayed_52__106_,chained_data_delayed_52__105_,
  chained_data_delayed_52__104_,chained_data_delayed_52__103_,
  chained_data_delayed_52__102_,chained_data_delayed_52__101_,chained_data_delayed_52__100_,
  chained_data_delayed_52__99_,chained_data_delayed_52__98_,chained_data_delayed_52__97_,
  chained_data_delayed_52__96_,chained_data_delayed_52__95_,chained_data_delayed_52__94_,
  chained_data_delayed_52__93_,chained_data_delayed_52__92_,
  chained_data_delayed_52__91_,chained_data_delayed_52__90_,chained_data_delayed_52__89_,
  chained_data_delayed_52__88_,chained_data_delayed_52__87_,chained_data_delayed_52__86_,
  chained_data_delayed_52__85_,chained_data_delayed_52__84_,chained_data_delayed_52__83_,
  chained_data_delayed_52__82_,chained_data_delayed_52__81_,
  chained_data_delayed_52__80_,chained_data_delayed_52__79_,chained_data_delayed_52__78_,
  chained_data_delayed_52__77_,chained_data_delayed_52__76_,chained_data_delayed_52__75_,
  chained_data_delayed_52__74_,chained_data_delayed_52__73_,chained_data_delayed_52__72_,
  chained_data_delayed_52__71_,chained_data_delayed_52__70_,
  chained_data_delayed_52__69_,chained_data_delayed_52__68_,chained_data_delayed_52__67_,
  chained_data_delayed_52__66_,chained_data_delayed_52__65_,chained_data_delayed_52__64_,
  chained_data_delayed_52__63_,chained_data_delayed_52__62_,chained_data_delayed_52__61_,
  chained_data_delayed_52__60_,chained_data_delayed_52__59_,chained_data_delayed_52__58_,
  chained_data_delayed_52__57_,chained_data_delayed_52__56_,
  chained_data_delayed_52__55_,chained_data_delayed_52__54_,chained_data_delayed_52__53_,
  chained_data_delayed_52__52_,chained_data_delayed_52__51_,chained_data_delayed_52__50_,
  chained_data_delayed_52__49_,chained_data_delayed_52__48_,chained_data_delayed_52__47_,
  chained_data_delayed_52__46_,chained_data_delayed_52__45_,
  chained_data_delayed_52__44_,chained_data_delayed_52__43_,chained_data_delayed_52__42_,
  chained_data_delayed_52__41_,chained_data_delayed_52__40_,chained_data_delayed_52__39_,
  chained_data_delayed_52__38_,chained_data_delayed_52__37_,chained_data_delayed_52__36_,
  chained_data_delayed_52__35_,chained_data_delayed_52__34_,
  chained_data_delayed_52__33_,chained_data_delayed_52__32_,chained_data_delayed_52__31_,
  chained_data_delayed_52__30_,chained_data_delayed_52__29_,chained_data_delayed_52__28_,
  chained_data_delayed_52__27_,chained_data_delayed_52__26_,chained_data_delayed_52__25_,
  chained_data_delayed_52__24_,chained_data_delayed_52__23_,
  chained_data_delayed_52__22_,chained_data_delayed_52__21_,chained_data_delayed_52__20_,
  chained_data_delayed_52__19_,chained_data_delayed_52__18_,chained_data_delayed_52__17_,
  chained_data_delayed_52__16_,chained_data_delayed_52__15_,chained_data_delayed_52__14_,
  chained_data_delayed_52__13_,chained_data_delayed_52__12_,
  chained_data_delayed_52__11_,chained_data_delayed_52__10_,chained_data_delayed_52__9_,
  chained_data_delayed_52__8_,chained_data_delayed_52__7_,chained_data_delayed_52__6_,
  chained_data_delayed_52__5_,chained_data_delayed_52__4_,chained_data_delayed_52__3_,
  chained_data_delayed_52__2_,chained_data_delayed_52__1_,chained_data_delayed_52__0_,
  chained_data_delayed_51__127_,chained_data_delayed_51__126_,
  chained_data_delayed_51__125_,chained_data_delayed_51__124_,chained_data_delayed_51__123_,
  chained_data_delayed_51__122_,chained_data_delayed_51__121_,chained_data_delayed_51__120_,
  chained_data_delayed_51__119_,chained_data_delayed_51__118_,
  chained_data_delayed_51__117_,chained_data_delayed_51__116_,chained_data_delayed_51__115_,
  chained_data_delayed_51__114_,chained_data_delayed_51__113_,chained_data_delayed_51__112_,
  chained_data_delayed_51__111_,chained_data_delayed_51__110_,
  chained_data_delayed_51__109_,chained_data_delayed_51__108_,chained_data_delayed_51__107_,
  chained_data_delayed_51__106_,chained_data_delayed_51__105_,chained_data_delayed_51__104_,
  chained_data_delayed_51__103_,chained_data_delayed_51__102_,
  chained_data_delayed_51__101_,chained_data_delayed_51__100_,chained_data_delayed_51__99_,
  chained_data_delayed_51__98_,chained_data_delayed_51__97_,chained_data_delayed_51__96_,
  chained_data_delayed_51__95_,chained_data_delayed_51__94_,chained_data_delayed_51__93_,
  chained_data_delayed_51__92_,chained_data_delayed_51__91_,
  chained_data_delayed_51__90_,chained_data_delayed_51__89_,chained_data_delayed_51__88_,
  chained_data_delayed_51__87_,chained_data_delayed_51__86_,chained_data_delayed_51__85_,
  chained_data_delayed_51__84_,chained_data_delayed_51__83_,chained_data_delayed_51__82_,
  chained_data_delayed_51__81_,chained_data_delayed_51__80_,
  chained_data_delayed_51__79_,chained_data_delayed_51__78_,chained_data_delayed_51__77_,
  chained_data_delayed_51__76_,chained_data_delayed_51__75_,chained_data_delayed_51__74_,
  chained_data_delayed_51__73_,chained_data_delayed_51__72_,chained_data_delayed_51__71_,
  chained_data_delayed_51__70_,chained_data_delayed_51__69_,chained_data_delayed_51__68_,
  chained_data_delayed_51__67_,chained_data_delayed_51__66_,
  chained_data_delayed_51__65_,chained_data_delayed_51__64_,chained_data_delayed_51__63_,
  chained_data_delayed_51__62_,chained_data_delayed_51__61_,chained_data_delayed_51__60_,
  chained_data_delayed_51__59_,chained_data_delayed_51__58_,chained_data_delayed_51__57_,
  chained_data_delayed_51__56_,chained_data_delayed_51__55_,
  chained_data_delayed_51__54_,chained_data_delayed_51__53_,chained_data_delayed_51__52_,
  chained_data_delayed_51__51_,chained_data_delayed_51__50_,chained_data_delayed_51__49_,
  chained_data_delayed_51__48_,chained_data_delayed_51__47_,chained_data_delayed_51__46_,
  chained_data_delayed_51__45_,chained_data_delayed_51__44_,
  chained_data_delayed_51__43_,chained_data_delayed_51__42_,chained_data_delayed_51__41_,
  chained_data_delayed_51__40_,chained_data_delayed_51__39_,chained_data_delayed_51__38_,
  chained_data_delayed_51__37_,chained_data_delayed_51__36_,chained_data_delayed_51__35_,
  chained_data_delayed_51__34_,chained_data_delayed_51__33_,
  chained_data_delayed_51__32_,chained_data_delayed_51__31_,chained_data_delayed_51__30_,
  chained_data_delayed_51__29_,chained_data_delayed_51__28_,chained_data_delayed_51__27_,
  chained_data_delayed_51__26_,chained_data_delayed_51__25_,chained_data_delayed_51__24_,
  chained_data_delayed_51__23_,chained_data_delayed_51__22_,
  chained_data_delayed_51__21_,chained_data_delayed_51__20_,chained_data_delayed_51__19_,
  chained_data_delayed_51__18_,chained_data_delayed_51__17_,chained_data_delayed_51__16_,
  chained_data_delayed_51__15_,chained_data_delayed_51__14_,chained_data_delayed_51__13_,
  chained_data_delayed_51__12_,chained_data_delayed_51__11_,
  chained_data_delayed_51__10_,chained_data_delayed_51__9_,chained_data_delayed_51__8_,
  chained_data_delayed_51__7_,chained_data_delayed_51__6_,chained_data_delayed_51__5_,
  chained_data_delayed_51__4_,chained_data_delayed_51__3_,chained_data_delayed_51__2_,
  chained_data_delayed_51__1_,chained_data_delayed_51__0_,chained_data_delayed_50__127_,
  chained_data_delayed_50__126_,chained_data_delayed_50__125_,
  chained_data_delayed_50__124_,chained_data_delayed_50__123_,chained_data_delayed_50__122_,
  chained_data_delayed_50__121_,chained_data_delayed_50__120_,chained_data_delayed_50__119_,
  chained_data_delayed_50__118_,chained_data_delayed_50__117_,
  chained_data_delayed_50__116_,chained_data_delayed_50__115_,chained_data_delayed_50__114_,
  chained_data_delayed_50__113_,chained_data_delayed_50__112_,chained_data_delayed_50__111_,
  chained_data_delayed_50__110_,chained_data_delayed_50__109_,
  chained_data_delayed_50__108_,chained_data_delayed_50__107_,chained_data_delayed_50__106_,
  chained_data_delayed_50__105_,chained_data_delayed_50__104_,chained_data_delayed_50__103_,
  chained_data_delayed_50__102_,chained_data_delayed_50__101_,
  chained_data_delayed_50__100_,chained_data_delayed_50__99_,chained_data_delayed_50__98_,
  chained_data_delayed_50__97_,chained_data_delayed_50__96_,chained_data_delayed_50__95_,
  chained_data_delayed_50__94_,chained_data_delayed_50__93_,chained_data_delayed_50__92_,
  chained_data_delayed_50__91_,chained_data_delayed_50__90_,
  chained_data_delayed_50__89_,chained_data_delayed_50__88_,chained_data_delayed_50__87_,
  chained_data_delayed_50__86_,chained_data_delayed_50__85_,chained_data_delayed_50__84_,
  chained_data_delayed_50__83_,chained_data_delayed_50__82_,chained_data_delayed_50__81_,
  chained_data_delayed_50__80_,chained_data_delayed_50__79_,chained_data_delayed_50__78_,
  chained_data_delayed_50__77_,chained_data_delayed_50__76_,
  chained_data_delayed_50__75_,chained_data_delayed_50__74_,chained_data_delayed_50__73_,
  chained_data_delayed_50__72_,chained_data_delayed_50__71_,chained_data_delayed_50__70_,
  chained_data_delayed_50__69_,chained_data_delayed_50__68_,chained_data_delayed_50__67_,
  chained_data_delayed_50__66_,chained_data_delayed_50__65_,
  chained_data_delayed_50__64_,chained_data_delayed_50__63_,chained_data_delayed_50__62_,
  chained_data_delayed_50__61_,chained_data_delayed_50__60_,chained_data_delayed_50__59_,
  chained_data_delayed_50__58_,chained_data_delayed_50__57_,chained_data_delayed_50__56_,
  chained_data_delayed_50__55_,chained_data_delayed_50__54_,
  chained_data_delayed_50__53_,chained_data_delayed_50__52_,chained_data_delayed_50__51_,
  chained_data_delayed_50__50_,chained_data_delayed_50__49_,chained_data_delayed_50__48_,
  chained_data_delayed_50__47_,chained_data_delayed_50__46_,chained_data_delayed_50__45_,
  chained_data_delayed_50__44_,chained_data_delayed_50__43_,
  chained_data_delayed_50__42_,chained_data_delayed_50__41_,chained_data_delayed_50__40_,
  chained_data_delayed_50__39_,chained_data_delayed_50__38_,chained_data_delayed_50__37_,
  chained_data_delayed_50__36_,chained_data_delayed_50__35_,chained_data_delayed_50__34_,
  chained_data_delayed_50__33_,chained_data_delayed_50__32_,
  chained_data_delayed_50__31_,chained_data_delayed_50__30_,chained_data_delayed_50__29_,
  chained_data_delayed_50__28_,chained_data_delayed_50__27_,chained_data_delayed_50__26_,
  chained_data_delayed_50__25_,chained_data_delayed_50__24_,chained_data_delayed_50__23_,
  chained_data_delayed_50__22_,chained_data_delayed_50__21_,
  chained_data_delayed_50__20_,chained_data_delayed_50__19_,chained_data_delayed_50__18_,
  chained_data_delayed_50__17_,chained_data_delayed_50__16_,chained_data_delayed_50__15_,
  chained_data_delayed_50__14_,chained_data_delayed_50__13_,chained_data_delayed_50__12_,
  chained_data_delayed_50__11_,chained_data_delayed_50__10_,chained_data_delayed_50__9_,
  chained_data_delayed_50__8_,chained_data_delayed_50__7_,
  chained_data_delayed_50__6_,chained_data_delayed_50__5_,chained_data_delayed_50__4_,
  chained_data_delayed_50__3_,chained_data_delayed_50__2_,chained_data_delayed_50__1_,
  chained_data_delayed_50__0_,chained_data_delayed_49__127_,chained_data_delayed_49__126_,
  chained_data_delayed_49__125_,chained_data_delayed_49__124_,
  chained_data_delayed_49__123_,chained_data_delayed_49__122_,chained_data_delayed_49__121_,
  chained_data_delayed_49__120_,chained_data_delayed_49__119_,chained_data_delayed_49__118_,
  chained_data_delayed_49__117_,chained_data_delayed_49__116_,
  chained_data_delayed_49__115_,chained_data_delayed_49__114_,chained_data_delayed_49__113_,
  chained_data_delayed_49__112_,chained_data_delayed_49__111_,chained_data_delayed_49__110_,
  chained_data_delayed_49__109_,chained_data_delayed_49__108_,
  chained_data_delayed_49__107_,chained_data_delayed_49__106_,chained_data_delayed_49__105_,
  chained_data_delayed_49__104_,chained_data_delayed_49__103_,chained_data_delayed_49__102_,
  chained_data_delayed_49__101_,chained_data_delayed_49__100_,
  chained_data_delayed_49__99_,chained_data_delayed_49__98_,chained_data_delayed_49__97_,
  chained_data_delayed_49__96_,chained_data_delayed_49__95_,chained_data_delayed_49__94_,
  chained_data_delayed_49__93_,chained_data_delayed_49__92_,chained_data_delayed_49__91_,
  chained_data_delayed_49__90_,chained_data_delayed_49__89_,chained_data_delayed_49__88_,
  chained_data_delayed_49__87_,chained_data_delayed_49__86_,
  chained_data_delayed_49__85_,chained_data_delayed_49__84_,chained_data_delayed_49__83_,
  chained_data_delayed_49__82_,chained_data_delayed_49__81_,chained_data_delayed_49__80_,
  chained_data_delayed_49__79_,chained_data_delayed_49__78_,chained_data_delayed_49__77_,
  chained_data_delayed_49__76_,chained_data_delayed_49__75_,
  chained_data_delayed_49__74_,chained_data_delayed_49__73_,chained_data_delayed_49__72_,
  chained_data_delayed_49__71_,chained_data_delayed_49__70_,chained_data_delayed_49__69_,
  chained_data_delayed_49__68_,chained_data_delayed_49__67_,chained_data_delayed_49__66_,
  chained_data_delayed_49__65_,chained_data_delayed_49__64_,
  chained_data_delayed_49__63_,chained_data_delayed_49__62_,chained_data_delayed_49__61_,
  chained_data_delayed_49__60_,chained_data_delayed_49__59_,chained_data_delayed_49__58_,
  chained_data_delayed_49__57_,chained_data_delayed_49__56_,chained_data_delayed_49__55_,
  chained_data_delayed_49__54_,chained_data_delayed_49__53_,
  chained_data_delayed_49__52_,chained_data_delayed_49__51_,chained_data_delayed_49__50_,
  chained_data_delayed_49__49_,chained_data_delayed_49__48_,chained_data_delayed_49__47_,
  chained_data_delayed_49__46_,chained_data_delayed_49__45_,chained_data_delayed_49__44_,
  chained_data_delayed_49__43_,chained_data_delayed_49__42_,
  chained_data_delayed_49__41_,chained_data_delayed_49__40_,chained_data_delayed_49__39_,
  chained_data_delayed_49__38_,chained_data_delayed_49__37_,chained_data_delayed_49__36_,
  chained_data_delayed_49__35_,chained_data_delayed_49__34_,chained_data_delayed_49__33_,
  chained_data_delayed_49__32_,chained_data_delayed_49__31_,
  chained_data_delayed_49__30_,chained_data_delayed_49__29_,chained_data_delayed_49__28_,
  chained_data_delayed_49__27_,chained_data_delayed_49__26_,chained_data_delayed_49__25_,
  chained_data_delayed_49__24_,chained_data_delayed_49__23_,chained_data_delayed_49__22_,
  chained_data_delayed_49__21_,chained_data_delayed_49__20_,
  chained_data_delayed_49__19_,chained_data_delayed_49__18_,chained_data_delayed_49__17_,
  chained_data_delayed_49__16_,chained_data_delayed_49__15_,chained_data_delayed_49__14_,
  chained_data_delayed_49__13_,chained_data_delayed_49__12_,chained_data_delayed_49__11_,
  chained_data_delayed_49__10_,chained_data_delayed_49__9_,chained_data_delayed_49__8_,
  chained_data_delayed_49__7_,chained_data_delayed_49__6_,
  chained_data_delayed_49__5_,chained_data_delayed_49__4_,chained_data_delayed_49__3_,
  chained_data_delayed_49__2_,chained_data_delayed_49__1_,chained_data_delayed_49__0_,
  chained_data_delayed_56__127_,chained_data_delayed_56__126_,chained_data_delayed_56__125_,
  chained_data_delayed_56__124_,chained_data_delayed_56__123_,
  chained_data_delayed_56__122_,chained_data_delayed_56__121_,chained_data_delayed_56__120_,
  chained_data_delayed_56__119_,chained_data_delayed_56__118_,chained_data_delayed_56__117_,
  chained_data_delayed_56__116_,chained_data_delayed_56__115_,
  chained_data_delayed_56__114_,chained_data_delayed_56__113_,chained_data_delayed_56__112_,
  chained_data_delayed_56__111_,chained_data_delayed_56__110_,chained_data_delayed_56__109_,
  chained_data_delayed_56__108_,chained_data_delayed_56__107_,
  chained_data_delayed_56__106_,chained_data_delayed_56__105_,chained_data_delayed_56__104_,
  chained_data_delayed_56__103_,chained_data_delayed_56__102_,chained_data_delayed_56__101_,
  chained_data_delayed_56__100_,chained_data_delayed_56__99_,chained_data_delayed_56__98_,
  chained_data_delayed_56__97_,chained_data_delayed_56__96_,
  chained_data_delayed_56__95_,chained_data_delayed_56__94_,chained_data_delayed_56__93_,
  chained_data_delayed_56__92_,chained_data_delayed_56__91_,chained_data_delayed_56__90_,
  chained_data_delayed_56__89_,chained_data_delayed_56__88_,chained_data_delayed_56__87_,
  chained_data_delayed_56__86_,chained_data_delayed_56__85_,
  chained_data_delayed_56__84_,chained_data_delayed_56__83_,chained_data_delayed_56__82_,
  chained_data_delayed_56__81_,chained_data_delayed_56__80_,chained_data_delayed_56__79_,
  chained_data_delayed_56__78_,chained_data_delayed_56__77_,chained_data_delayed_56__76_,
  chained_data_delayed_56__75_,chained_data_delayed_56__74_,
  chained_data_delayed_56__73_,chained_data_delayed_56__72_,chained_data_delayed_56__71_,
  chained_data_delayed_56__70_,chained_data_delayed_56__69_,chained_data_delayed_56__68_,
  chained_data_delayed_56__67_,chained_data_delayed_56__66_,chained_data_delayed_56__65_,
  chained_data_delayed_56__64_,chained_data_delayed_56__63_,
  chained_data_delayed_56__62_,chained_data_delayed_56__61_,chained_data_delayed_56__60_,
  chained_data_delayed_56__59_,chained_data_delayed_56__58_,chained_data_delayed_56__57_,
  chained_data_delayed_56__56_,chained_data_delayed_56__55_,chained_data_delayed_56__54_,
  chained_data_delayed_56__53_,chained_data_delayed_56__52_,
  chained_data_delayed_56__51_,chained_data_delayed_56__50_,chained_data_delayed_56__49_,
  chained_data_delayed_56__48_,chained_data_delayed_56__47_,chained_data_delayed_56__46_,
  chained_data_delayed_56__45_,chained_data_delayed_56__44_,chained_data_delayed_56__43_,
  chained_data_delayed_56__42_,chained_data_delayed_56__41_,
  chained_data_delayed_56__40_,chained_data_delayed_56__39_,chained_data_delayed_56__38_,
  chained_data_delayed_56__37_,chained_data_delayed_56__36_,chained_data_delayed_56__35_,
  chained_data_delayed_56__34_,chained_data_delayed_56__33_,chained_data_delayed_56__32_,
  chained_data_delayed_56__31_,chained_data_delayed_56__30_,
  chained_data_delayed_56__29_,chained_data_delayed_56__28_,chained_data_delayed_56__27_,
  chained_data_delayed_56__26_,chained_data_delayed_56__25_,chained_data_delayed_56__24_,
  chained_data_delayed_56__23_,chained_data_delayed_56__22_,chained_data_delayed_56__21_,
  chained_data_delayed_56__20_,chained_data_delayed_56__19_,chained_data_delayed_56__18_,
  chained_data_delayed_56__17_,chained_data_delayed_56__16_,
  chained_data_delayed_56__15_,chained_data_delayed_56__14_,chained_data_delayed_56__13_,
  chained_data_delayed_56__12_,chained_data_delayed_56__11_,chained_data_delayed_56__10_,
  chained_data_delayed_56__9_,chained_data_delayed_56__8_,chained_data_delayed_56__7_,
  chained_data_delayed_56__6_,chained_data_delayed_56__5_,chained_data_delayed_56__4_,
  chained_data_delayed_56__3_,chained_data_delayed_56__2_,
  chained_data_delayed_56__1_,chained_data_delayed_56__0_,chained_data_delayed_55__127_,
  chained_data_delayed_55__126_,chained_data_delayed_55__125_,chained_data_delayed_55__124_,
  chained_data_delayed_55__123_,chained_data_delayed_55__122_,
  chained_data_delayed_55__121_,chained_data_delayed_55__120_,chained_data_delayed_55__119_,
  chained_data_delayed_55__118_,chained_data_delayed_55__117_,chained_data_delayed_55__116_,
  chained_data_delayed_55__115_,chained_data_delayed_55__114_,
  chained_data_delayed_55__113_,chained_data_delayed_55__112_,chained_data_delayed_55__111_,
  chained_data_delayed_55__110_,chained_data_delayed_55__109_,chained_data_delayed_55__108_,
  chained_data_delayed_55__107_,chained_data_delayed_55__106_,
  chained_data_delayed_55__105_,chained_data_delayed_55__104_,chained_data_delayed_55__103_,
  chained_data_delayed_55__102_,chained_data_delayed_55__101_,chained_data_delayed_55__100_,
  chained_data_delayed_55__99_,chained_data_delayed_55__98_,chained_data_delayed_55__97_,
  chained_data_delayed_55__96_,chained_data_delayed_55__95_,
  chained_data_delayed_55__94_,chained_data_delayed_55__93_,chained_data_delayed_55__92_,
  chained_data_delayed_55__91_,chained_data_delayed_55__90_,chained_data_delayed_55__89_,
  chained_data_delayed_55__88_,chained_data_delayed_55__87_,chained_data_delayed_55__86_,
  chained_data_delayed_55__85_,chained_data_delayed_55__84_,
  chained_data_delayed_55__83_,chained_data_delayed_55__82_,chained_data_delayed_55__81_,
  chained_data_delayed_55__80_,chained_data_delayed_55__79_,chained_data_delayed_55__78_,
  chained_data_delayed_55__77_,chained_data_delayed_55__76_,chained_data_delayed_55__75_,
  chained_data_delayed_55__74_,chained_data_delayed_55__73_,
  chained_data_delayed_55__72_,chained_data_delayed_55__71_,chained_data_delayed_55__70_,
  chained_data_delayed_55__69_,chained_data_delayed_55__68_,chained_data_delayed_55__67_,
  chained_data_delayed_55__66_,chained_data_delayed_55__65_,chained_data_delayed_55__64_,
  chained_data_delayed_55__63_,chained_data_delayed_55__62_,
  chained_data_delayed_55__61_,chained_data_delayed_55__60_,chained_data_delayed_55__59_,
  chained_data_delayed_55__58_,chained_data_delayed_55__57_,chained_data_delayed_55__56_,
  chained_data_delayed_55__55_,chained_data_delayed_55__54_,chained_data_delayed_55__53_,
  chained_data_delayed_55__52_,chained_data_delayed_55__51_,
  chained_data_delayed_55__50_,chained_data_delayed_55__49_,chained_data_delayed_55__48_,
  chained_data_delayed_55__47_,chained_data_delayed_55__46_,chained_data_delayed_55__45_,
  chained_data_delayed_55__44_,chained_data_delayed_55__43_,chained_data_delayed_55__42_,
  chained_data_delayed_55__41_,chained_data_delayed_55__40_,
  chained_data_delayed_55__39_,chained_data_delayed_55__38_,chained_data_delayed_55__37_,
  chained_data_delayed_55__36_,chained_data_delayed_55__35_,chained_data_delayed_55__34_,
  chained_data_delayed_55__33_,chained_data_delayed_55__32_,chained_data_delayed_55__31_,
  chained_data_delayed_55__30_,chained_data_delayed_55__29_,chained_data_delayed_55__28_,
  chained_data_delayed_55__27_,chained_data_delayed_55__26_,
  chained_data_delayed_55__25_,chained_data_delayed_55__24_,chained_data_delayed_55__23_,
  chained_data_delayed_55__22_,chained_data_delayed_55__21_,chained_data_delayed_55__20_,
  chained_data_delayed_55__19_,chained_data_delayed_55__18_,chained_data_delayed_55__17_,
  chained_data_delayed_55__16_,chained_data_delayed_55__15_,
  chained_data_delayed_55__14_,chained_data_delayed_55__13_,chained_data_delayed_55__12_,
  chained_data_delayed_55__11_,chained_data_delayed_55__10_,chained_data_delayed_55__9_,
  chained_data_delayed_55__8_,chained_data_delayed_55__7_,chained_data_delayed_55__6_,
  chained_data_delayed_55__5_,chained_data_delayed_55__4_,chained_data_delayed_55__3_,
  chained_data_delayed_55__2_,chained_data_delayed_55__1_,
  chained_data_delayed_55__0_,chained_data_delayed_54__127_,chained_data_delayed_54__126_,
  chained_data_delayed_54__125_,chained_data_delayed_54__124_,chained_data_delayed_54__123_,
  chained_data_delayed_54__122_,chained_data_delayed_54__121_,
  chained_data_delayed_54__120_,chained_data_delayed_54__119_,chained_data_delayed_54__118_,
  chained_data_delayed_54__117_,chained_data_delayed_54__116_,chained_data_delayed_54__115_,
  chained_data_delayed_54__114_,chained_data_delayed_54__113_,
  chained_data_delayed_54__112_,chained_data_delayed_54__111_,chained_data_delayed_54__110_,
  chained_data_delayed_54__109_,chained_data_delayed_54__108_,chained_data_delayed_54__107_,
  chained_data_delayed_54__106_,chained_data_delayed_54__105_,
  chained_data_delayed_54__104_,chained_data_delayed_54__103_,chained_data_delayed_54__102_,
  chained_data_delayed_54__101_,chained_data_delayed_54__100_,chained_data_delayed_54__99_,
  chained_data_delayed_54__98_,chained_data_delayed_54__97_,chained_data_delayed_54__96_,
  chained_data_delayed_54__95_,chained_data_delayed_54__94_,
  chained_data_delayed_54__93_,chained_data_delayed_54__92_,chained_data_delayed_54__91_,
  chained_data_delayed_54__90_,chained_data_delayed_54__89_,chained_data_delayed_54__88_,
  chained_data_delayed_54__87_,chained_data_delayed_54__86_,chained_data_delayed_54__85_,
  chained_data_delayed_54__84_,chained_data_delayed_54__83_,
  chained_data_delayed_54__82_,chained_data_delayed_54__81_,chained_data_delayed_54__80_,
  chained_data_delayed_54__79_,chained_data_delayed_54__78_,chained_data_delayed_54__77_,
  chained_data_delayed_54__76_,chained_data_delayed_54__75_,chained_data_delayed_54__74_,
  chained_data_delayed_54__73_,chained_data_delayed_54__72_,
  chained_data_delayed_54__71_,chained_data_delayed_54__70_,chained_data_delayed_54__69_,
  chained_data_delayed_54__68_,chained_data_delayed_54__67_,chained_data_delayed_54__66_,
  chained_data_delayed_54__65_,chained_data_delayed_54__64_,chained_data_delayed_54__63_,
  chained_data_delayed_54__62_,chained_data_delayed_54__61_,
  chained_data_delayed_54__60_,chained_data_delayed_54__59_,chained_data_delayed_54__58_,
  chained_data_delayed_54__57_,chained_data_delayed_54__56_,chained_data_delayed_54__55_,
  chained_data_delayed_54__54_,chained_data_delayed_54__53_,chained_data_delayed_54__52_,
  chained_data_delayed_54__51_,chained_data_delayed_54__50_,
  chained_data_delayed_54__49_,chained_data_delayed_54__48_,chained_data_delayed_54__47_,
  chained_data_delayed_54__46_,chained_data_delayed_54__45_,chained_data_delayed_54__44_,
  chained_data_delayed_54__43_,chained_data_delayed_54__42_,chained_data_delayed_54__41_,
  chained_data_delayed_54__40_,chained_data_delayed_54__39_,chained_data_delayed_54__38_,
  chained_data_delayed_54__37_,chained_data_delayed_54__36_,
  chained_data_delayed_54__35_,chained_data_delayed_54__34_,chained_data_delayed_54__33_,
  chained_data_delayed_54__32_,chained_data_delayed_54__31_,chained_data_delayed_54__30_,
  chained_data_delayed_54__29_,chained_data_delayed_54__28_,chained_data_delayed_54__27_,
  chained_data_delayed_54__26_,chained_data_delayed_54__25_,
  chained_data_delayed_54__24_,chained_data_delayed_54__23_,chained_data_delayed_54__22_,
  chained_data_delayed_54__21_,chained_data_delayed_54__20_,chained_data_delayed_54__19_,
  chained_data_delayed_54__18_,chained_data_delayed_54__17_,chained_data_delayed_54__16_,
  chained_data_delayed_54__15_,chained_data_delayed_54__14_,
  chained_data_delayed_54__13_,chained_data_delayed_54__12_,chained_data_delayed_54__11_,
  chained_data_delayed_54__10_,chained_data_delayed_54__9_,chained_data_delayed_54__8_,
  chained_data_delayed_54__7_,chained_data_delayed_54__6_,chained_data_delayed_54__5_,
  chained_data_delayed_54__4_,chained_data_delayed_54__3_,chained_data_delayed_54__2_,
  chained_data_delayed_54__1_,chained_data_delayed_54__0_,
  chained_data_delayed_53__127_,chained_data_delayed_53__126_,chained_data_delayed_53__125_,
  chained_data_delayed_53__124_,chained_data_delayed_53__123_,chained_data_delayed_53__122_,
  chained_data_delayed_53__121_,chained_data_delayed_53__120_,
  chained_data_delayed_53__119_,chained_data_delayed_53__118_,chained_data_delayed_53__117_,
  chained_data_delayed_53__116_,chained_data_delayed_53__115_,chained_data_delayed_53__114_,
  chained_data_delayed_53__113_,chained_data_delayed_53__112_,
  chained_data_delayed_53__111_,chained_data_delayed_53__110_,chained_data_delayed_53__109_,
  chained_data_delayed_53__108_,chained_data_delayed_53__107_,chained_data_delayed_53__106_,
  chained_data_delayed_53__105_,chained_data_delayed_53__104_,
  chained_data_delayed_53__103_,chained_data_delayed_53__102_,chained_data_delayed_53__101_,
  chained_data_delayed_53__100_,chained_data_delayed_53__99_,chained_data_delayed_53__98_,
  chained_data_delayed_53__97_,chained_data_delayed_53__96_,chained_data_delayed_53__95_,
  chained_data_delayed_53__94_,chained_data_delayed_53__93_,
  chained_data_delayed_53__92_,chained_data_delayed_53__91_,chained_data_delayed_53__90_,
  chained_data_delayed_53__89_,chained_data_delayed_53__88_,chained_data_delayed_53__87_,
  chained_data_delayed_53__86_,chained_data_delayed_53__85_,chained_data_delayed_53__84_,
  chained_data_delayed_53__83_,chained_data_delayed_53__82_,
  chained_data_delayed_53__81_,chained_data_delayed_53__80_,chained_data_delayed_53__79_,
  chained_data_delayed_53__78_,chained_data_delayed_53__77_,chained_data_delayed_53__76_,
  chained_data_delayed_53__75_,chained_data_delayed_53__74_,chained_data_delayed_53__73_,
  chained_data_delayed_53__72_,chained_data_delayed_53__71_,
  chained_data_delayed_53__70_,chained_data_delayed_53__69_,chained_data_delayed_53__68_,
  chained_data_delayed_53__67_,chained_data_delayed_53__66_,chained_data_delayed_53__65_,
  chained_data_delayed_53__64_,chained_data_delayed_53__63_,chained_data_delayed_53__62_,
  chained_data_delayed_53__61_,chained_data_delayed_53__60_,
  chained_data_delayed_53__59_,chained_data_delayed_53__58_,chained_data_delayed_53__57_,
  chained_data_delayed_53__56_,chained_data_delayed_53__55_,chained_data_delayed_53__54_,
  chained_data_delayed_53__53_,chained_data_delayed_53__52_,chained_data_delayed_53__51_,
  chained_data_delayed_53__50_,chained_data_delayed_53__49_,chained_data_delayed_53__48_,
  chained_data_delayed_53__47_,chained_data_delayed_53__46_,
  chained_data_delayed_53__45_,chained_data_delayed_53__44_,chained_data_delayed_53__43_,
  chained_data_delayed_53__42_,chained_data_delayed_53__41_,chained_data_delayed_53__40_,
  chained_data_delayed_53__39_,chained_data_delayed_53__38_,chained_data_delayed_53__37_,
  chained_data_delayed_53__36_,chained_data_delayed_53__35_,
  chained_data_delayed_53__34_,chained_data_delayed_53__33_,chained_data_delayed_53__32_,
  chained_data_delayed_53__31_,chained_data_delayed_53__30_,chained_data_delayed_53__29_,
  chained_data_delayed_53__28_,chained_data_delayed_53__27_,chained_data_delayed_53__26_,
  chained_data_delayed_53__25_,chained_data_delayed_53__24_,
  chained_data_delayed_53__23_,chained_data_delayed_53__22_,chained_data_delayed_53__21_,
  chained_data_delayed_53__20_,chained_data_delayed_53__19_,chained_data_delayed_53__18_,
  chained_data_delayed_53__17_,chained_data_delayed_53__16_,chained_data_delayed_53__15_,
  chained_data_delayed_53__14_,chained_data_delayed_53__13_,
  chained_data_delayed_53__12_,chained_data_delayed_53__11_,chained_data_delayed_53__10_,
  chained_data_delayed_53__9_,chained_data_delayed_53__8_,chained_data_delayed_53__7_,
  chained_data_delayed_53__6_,chained_data_delayed_53__5_,chained_data_delayed_53__4_,
  chained_data_delayed_53__3_,chained_data_delayed_53__2_,chained_data_delayed_53__1_,
  chained_data_delayed_53__0_,chained_data_delayed_60__127_,
  chained_data_delayed_60__126_,chained_data_delayed_60__125_,chained_data_delayed_60__124_,
  chained_data_delayed_60__123_,chained_data_delayed_60__122_,chained_data_delayed_60__121_,
  chained_data_delayed_60__120_,chained_data_delayed_60__119_,
  chained_data_delayed_60__118_,chained_data_delayed_60__117_,chained_data_delayed_60__116_,
  chained_data_delayed_60__115_,chained_data_delayed_60__114_,chained_data_delayed_60__113_,
  chained_data_delayed_60__112_,chained_data_delayed_60__111_,
  chained_data_delayed_60__110_,chained_data_delayed_60__109_,chained_data_delayed_60__108_,
  chained_data_delayed_60__107_,chained_data_delayed_60__106_,chained_data_delayed_60__105_,
  chained_data_delayed_60__104_,chained_data_delayed_60__103_,
  chained_data_delayed_60__102_,chained_data_delayed_60__101_,chained_data_delayed_60__100_,
  chained_data_delayed_60__99_,chained_data_delayed_60__98_,chained_data_delayed_60__97_,
  chained_data_delayed_60__96_,chained_data_delayed_60__95_,chained_data_delayed_60__94_,
  chained_data_delayed_60__93_,chained_data_delayed_60__92_,
  chained_data_delayed_60__91_,chained_data_delayed_60__90_,chained_data_delayed_60__89_,
  chained_data_delayed_60__88_,chained_data_delayed_60__87_,chained_data_delayed_60__86_,
  chained_data_delayed_60__85_,chained_data_delayed_60__84_,chained_data_delayed_60__83_,
  chained_data_delayed_60__82_,chained_data_delayed_60__81_,
  chained_data_delayed_60__80_,chained_data_delayed_60__79_,chained_data_delayed_60__78_,
  chained_data_delayed_60__77_,chained_data_delayed_60__76_,chained_data_delayed_60__75_,
  chained_data_delayed_60__74_,chained_data_delayed_60__73_,chained_data_delayed_60__72_,
  chained_data_delayed_60__71_,chained_data_delayed_60__70_,
  chained_data_delayed_60__69_,chained_data_delayed_60__68_,chained_data_delayed_60__67_,
  chained_data_delayed_60__66_,chained_data_delayed_60__65_,chained_data_delayed_60__64_,
  chained_data_delayed_60__63_,chained_data_delayed_60__62_,chained_data_delayed_60__61_,
  chained_data_delayed_60__60_,chained_data_delayed_60__59_,chained_data_delayed_60__58_,
  chained_data_delayed_60__57_,chained_data_delayed_60__56_,
  chained_data_delayed_60__55_,chained_data_delayed_60__54_,chained_data_delayed_60__53_,
  chained_data_delayed_60__52_,chained_data_delayed_60__51_,chained_data_delayed_60__50_,
  chained_data_delayed_60__49_,chained_data_delayed_60__48_,chained_data_delayed_60__47_,
  chained_data_delayed_60__46_,chained_data_delayed_60__45_,
  chained_data_delayed_60__44_,chained_data_delayed_60__43_,chained_data_delayed_60__42_,
  chained_data_delayed_60__41_,chained_data_delayed_60__40_,chained_data_delayed_60__39_,
  chained_data_delayed_60__38_,chained_data_delayed_60__37_,chained_data_delayed_60__36_,
  chained_data_delayed_60__35_,chained_data_delayed_60__34_,
  chained_data_delayed_60__33_,chained_data_delayed_60__32_,chained_data_delayed_60__31_,
  chained_data_delayed_60__30_,chained_data_delayed_60__29_,chained_data_delayed_60__28_,
  chained_data_delayed_60__27_,chained_data_delayed_60__26_,chained_data_delayed_60__25_,
  chained_data_delayed_60__24_,chained_data_delayed_60__23_,
  chained_data_delayed_60__22_,chained_data_delayed_60__21_,chained_data_delayed_60__20_,
  chained_data_delayed_60__19_,chained_data_delayed_60__18_,chained_data_delayed_60__17_,
  chained_data_delayed_60__16_,chained_data_delayed_60__15_,chained_data_delayed_60__14_,
  chained_data_delayed_60__13_,chained_data_delayed_60__12_,
  chained_data_delayed_60__11_,chained_data_delayed_60__10_,chained_data_delayed_60__9_,
  chained_data_delayed_60__8_,chained_data_delayed_60__7_,chained_data_delayed_60__6_,
  chained_data_delayed_60__5_,chained_data_delayed_60__4_,chained_data_delayed_60__3_,
  chained_data_delayed_60__2_,chained_data_delayed_60__1_,chained_data_delayed_60__0_,
  chained_data_delayed_59__127_,chained_data_delayed_59__126_,
  chained_data_delayed_59__125_,chained_data_delayed_59__124_,chained_data_delayed_59__123_,
  chained_data_delayed_59__122_,chained_data_delayed_59__121_,chained_data_delayed_59__120_,
  chained_data_delayed_59__119_,chained_data_delayed_59__118_,
  chained_data_delayed_59__117_,chained_data_delayed_59__116_,chained_data_delayed_59__115_,
  chained_data_delayed_59__114_,chained_data_delayed_59__113_,chained_data_delayed_59__112_,
  chained_data_delayed_59__111_,chained_data_delayed_59__110_,
  chained_data_delayed_59__109_,chained_data_delayed_59__108_,chained_data_delayed_59__107_,
  chained_data_delayed_59__106_,chained_data_delayed_59__105_,chained_data_delayed_59__104_,
  chained_data_delayed_59__103_,chained_data_delayed_59__102_,
  chained_data_delayed_59__101_,chained_data_delayed_59__100_,chained_data_delayed_59__99_,
  chained_data_delayed_59__98_,chained_data_delayed_59__97_,chained_data_delayed_59__96_,
  chained_data_delayed_59__95_,chained_data_delayed_59__94_,chained_data_delayed_59__93_,
  chained_data_delayed_59__92_,chained_data_delayed_59__91_,
  chained_data_delayed_59__90_,chained_data_delayed_59__89_,chained_data_delayed_59__88_,
  chained_data_delayed_59__87_,chained_data_delayed_59__86_,chained_data_delayed_59__85_,
  chained_data_delayed_59__84_,chained_data_delayed_59__83_,chained_data_delayed_59__82_,
  chained_data_delayed_59__81_,chained_data_delayed_59__80_,
  chained_data_delayed_59__79_,chained_data_delayed_59__78_,chained_data_delayed_59__77_,
  chained_data_delayed_59__76_,chained_data_delayed_59__75_,chained_data_delayed_59__74_,
  chained_data_delayed_59__73_,chained_data_delayed_59__72_,chained_data_delayed_59__71_,
  chained_data_delayed_59__70_,chained_data_delayed_59__69_,chained_data_delayed_59__68_,
  chained_data_delayed_59__67_,chained_data_delayed_59__66_,
  chained_data_delayed_59__65_,chained_data_delayed_59__64_,chained_data_delayed_59__63_,
  chained_data_delayed_59__62_,chained_data_delayed_59__61_,chained_data_delayed_59__60_,
  chained_data_delayed_59__59_,chained_data_delayed_59__58_,chained_data_delayed_59__57_,
  chained_data_delayed_59__56_,chained_data_delayed_59__55_,
  chained_data_delayed_59__54_,chained_data_delayed_59__53_,chained_data_delayed_59__52_,
  chained_data_delayed_59__51_,chained_data_delayed_59__50_,chained_data_delayed_59__49_,
  chained_data_delayed_59__48_,chained_data_delayed_59__47_,chained_data_delayed_59__46_,
  chained_data_delayed_59__45_,chained_data_delayed_59__44_,
  chained_data_delayed_59__43_,chained_data_delayed_59__42_,chained_data_delayed_59__41_,
  chained_data_delayed_59__40_,chained_data_delayed_59__39_,chained_data_delayed_59__38_,
  chained_data_delayed_59__37_,chained_data_delayed_59__36_,chained_data_delayed_59__35_,
  chained_data_delayed_59__34_,chained_data_delayed_59__33_,
  chained_data_delayed_59__32_,chained_data_delayed_59__31_,chained_data_delayed_59__30_,
  chained_data_delayed_59__29_,chained_data_delayed_59__28_,chained_data_delayed_59__27_,
  chained_data_delayed_59__26_,chained_data_delayed_59__25_,chained_data_delayed_59__24_,
  chained_data_delayed_59__23_,chained_data_delayed_59__22_,
  chained_data_delayed_59__21_,chained_data_delayed_59__20_,chained_data_delayed_59__19_,
  chained_data_delayed_59__18_,chained_data_delayed_59__17_,chained_data_delayed_59__16_,
  chained_data_delayed_59__15_,chained_data_delayed_59__14_,chained_data_delayed_59__13_,
  chained_data_delayed_59__12_,chained_data_delayed_59__11_,
  chained_data_delayed_59__10_,chained_data_delayed_59__9_,chained_data_delayed_59__8_,
  chained_data_delayed_59__7_,chained_data_delayed_59__6_,chained_data_delayed_59__5_,
  chained_data_delayed_59__4_,chained_data_delayed_59__3_,chained_data_delayed_59__2_,
  chained_data_delayed_59__1_,chained_data_delayed_59__0_,chained_data_delayed_58__127_,
  chained_data_delayed_58__126_,chained_data_delayed_58__125_,
  chained_data_delayed_58__124_,chained_data_delayed_58__123_,chained_data_delayed_58__122_,
  chained_data_delayed_58__121_,chained_data_delayed_58__120_,chained_data_delayed_58__119_,
  chained_data_delayed_58__118_,chained_data_delayed_58__117_,
  chained_data_delayed_58__116_,chained_data_delayed_58__115_,chained_data_delayed_58__114_,
  chained_data_delayed_58__113_,chained_data_delayed_58__112_,chained_data_delayed_58__111_,
  chained_data_delayed_58__110_,chained_data_delayed_58__109_,
  chained_data_delayed_58__108_,chained_data_delayed_58__107_,chained_data_delayed_58__106_,
  chained_data_delayed_58__105_,chained_data_delayed_58__104_,chained_data_delayed_58__103_,
  chained_data_delayed_58__102_,chained_data_delayed_58__101_,
  chained_data_delayed_58__100_,chained_data_delayed_58__99_,chained_data_delayed_58__98_,
  chained_data_delayed_58__97_,chained_data_delayed_58__96_,chained_data_delayed_58__95_,
  chained_data_delayed_58__94_,chained_data_delayed_58__93_,chained_data_delayed_58__92_,
  chained_data_delayed_58__91_,chained_data_delayed_58__90_,
  chained_data_delayed_58__89_,chained_data_delayed_58__88_,chained_data_delayed_58__87_,
  chained_data_delayed_58__86_,chained_data_delayed_58__85_,chained_data_delayed_58__84_,
  chained_data_delayed_58__83_,chained_data_delayed_58__82_,chained_data_delayed_58__81_,
  chained_data_delayed_58__80_,chained_data_delayed_58__79_,chained_data_delayed_58__78_,
  chained_data_delayed_58__77_,chained_data_delayed_58__76_,
  chained_data_delayed_58__75_,chained_data_delayed_58__74_,chained_data_delayed_58__73_,
  chained_data_delayed_58__72_,chained_data_delayed_58__71_,chained_data_delayed_58__70_,
  chained_data_delayed_58__69_,chained_data_delayed_58__68_,chained_data_delayed_58__67_,
  chained_data_delayed_58__66_,chained_data_delayed_58__65_,
  chained_data_delayed_58__64_,chained_data_delayed_58__63_,chained_data_delayed_58__62_,
  chained_data_delayed_58__61_,chained_data_delayed_58__60_,chained_data_delayed_58__59_,
  chained_data_delayed_58__58_,chained_data_delayed_58__57_,chained_data_delayed_58__56_,
  chained_data_delayed_58__55_,chained_data_delayed_58__54_,
  chained_data_delayed_58__53_,chained_data_delayed_58__52_,chained_data_delayed_58__51_,
  chained_data_delayed_58__50_,chained_data_delayed_58__49_,chained_data_delayed_58__48_,
  chained_data_delayed_58__47_,chained_data_delayed_58__46_,chained_data_delayed_58__45_,
  chained_data_delayed_58__44_,chained_data_delayed_58__43_,
  chained_data_delayed_58__42_,chained_data_delayed_58__41_,chained_data_delayed_58__40_,
  chained_data_delayed_58__39_,chained_data_delayed_58__38_,chained_data_delayed_58__37_,
  chained_data_delayed_58__36_,chained_data_delayed_58__35_,chained_data_delayed_58__34_,
  chained_data_delayed_58__33_,chained_data_delayed_58__32_,
  chained_data_delayed_58__31_,chained_data_delayed_58__30_,chained_data_delayed_58__29_,
  chained_data_delayed_58__28_,chained_data_delayed_58__27_,chained_data_delayed_58__26_,
  chained_data_delayed_58__25_,chained_data_delayed_58__24_,chained_data_delayed_58__23_,
  chained_data_delayed_58__22_,chained_data_delayed_58__21_,
  chained_data_delayed_58__20_,chained_data_delayed_58__19_,chained_data_delayed_58__18_,
  chained_data_delayed_58__17_,chained_data_delayed_58__16_,chained_data_delayed_58__15_,
  chained_data_delayed_58__14_,chained_data_delayed_58__13_,chained_data_delayed_58__12_,
  chained_data_delayed_58__11_,chained_data_delayed_58__10_,chained_data_delayed_58__9_,
  chained_data_delayed_58__8_,chained_data_delayed_58__7_,
  chained_data_delayed_58__6_,chained_data_delayed_58__5_,chained_data_delayed_58__4_,
  chained_data_delayed_58__3_,chained_data_delayed_58__2_,chained_data_delayed_58__1_,
  chained_data_delayed_58__0_,chained_data_delayed_57__127_,chained_data_delayed_57__126_,
  chained_data_delayed_57__125_,chained_data_delayed_57__124_,
  chained_data_delayed_57__123_,chained_data_delayed_57__122_,chained_data_delayed_57__121_,
  chained_data_delayed_57__120_,chained_data_delayed_57__119_,chained_data_delayed_57__118_,
  chained_data_delayed_57__117_,chained_data_delayed_57__116_,
  chained_data_delayed_57__115_,chained_data_delayed_57__114_,chained_data_delayed_57__113_,
  chained_data_delayed_57__112_,chained_data_delayed_57__111_,chained_data_delayed_57__110_,
  chained_data_delayed_57__109_,chained_data_delayed_57__108_,
  chained_data_delayed_57__107_,chained_data_delayed_57__106_,chained_data_delayed_57__105_,
  chained_data_delayed_57__104_,chained_data_delayed_57__103_,chained_data_delayed_57__102_,
  chained_data_delayed_57__101_,chained_data_delayed_57__100_,
  chained_data_delayed_57__99_,chained_data_delayed_57__98_,chained_data_delayed_57__97_,
  chained_data_delayed_57__96_,chained_data_delayed_57__95_,chained_data_delayed_57__94_,
  chained_data_delayed_57__93_,chained_data_delayed_57__92_,chained_data_delayed_57__91_,
  chained_data_delayed_57__90_,chained_data_delayed_57__89_,chained_data_delayed_57__88_,
  chained_data_delayed_57__87_,chained_data_delayed_57__86_,
  chained_data_delayed_57__85_,chained_data_delayed_57__84_,chained_data_delayed_57__83_,
  chained_data_delayed_57__82_,chained_data_delayed_57__81_,chained_data_delayed_57__80_,
  chained_data_delayed_57__79_,chained_data_delayed_57__78_,chained_data_delayed_57__77_,
  chained_data_delayed_57__76_,chained_data_delayed_57__75_,
  chained_data_delayed_57__74_,chained_data_delayed_57__73_,chained_data_delayed_57__72_,
  chained_data_delayed_57__71_,chained_data_delayed_57__70_,chained_data_delayed_57__69_,
  chained_data_delayed_57__68_,chained_data_delayed_57__67_,chained_data_delayed_57__66_,
  chained_data_delayed_57__65_,chained_data_delayed_57__64_,
  chained_data_delayed_57__63_,chained_data_delayed_57__62_,chained_data_delayed_57__61_,
  chained_data_delayed_57__60_,chained_data_delayed_57__59_,chained_data_delayed_57__58_,
  chained_data_delayed_57__57_,chained_data_delayed_57__56_,chained_data_delayed_57__55_,
  chained_data_delayed_57__54_,chained_data_delayed_57__53_,
  chained_data_delayed_57__52_,chained_data_delayed_57__51_,chained_data_delayed_57__50_,
  chained_data_delayed_57__49_,chained_data_delayed_57__48_,chained_data_delayed_57__47_,
  chained_data_delayed_57__46_,chained_data_delayed_57__45_,chained_data_delayed_57__44_,
  chained_data_delayed_57__43_,chained_data_delayed_57__42_,
  chained_data_delayed_57__41_,chained_data_delayed_57__40_,chained_data_delayed_57__39_,
  chained_data_delayed_57__38_,chained_data_delayed_57__37_,chained_data_delayed_57__36_,
  chained_data_delayed_57__35_,chained_data_delayed_57__34_,chained_data_delayed_57__33_,
  chained_data_delayed_57__32_,chained_data_delayed_57__31_,
  chained_data_delayed_57__30_,chained_data_delayed_57__29_,chained_data_delayed_57__28_,
  chained_data_delayed_57__27_,chained_data_delayed_57__26_,chained_data_delayed_57__25_,
  chained_data_delayed_57__24_,chained_data_delayed_57__23_,chained_data_delayed_57__22_,
  chained_data_delayed_57__21_,chained_data_delayed_57__20_,
  chained_data_delayed_57__19_,chained_data_delayed_57__18_,chained_data_delayed_57__17_,
  chained_data_delayed_57__16_,chained_data_delayed_57__15_,chained_data_delayed_57__14_,
  chained_data_delayed_57__13_,chained_data_delayed_57__12_,chained_data_delayed_57__11_,
  chained_data_delayed_57__10_,chained_data_delayed_57__9_,chained_data_delayed_57__8_,
  chained_data_delayed_57__7_,chained_data_delayed_57__6_,
  chained_data_delayed_57__5_,chained_data_delayed_57__4_,chained_data_delayed_57__3_,
  chained_data_delayed_57__2_,chained_data_delayed_57__1_,chained_data_delayed_57__0_,
  chained_data_delayed_64__127_,chained_data_delayed_64__126_,chained_data_delayed_64__125_,
  chained_data_delayed_64__124_,chained_data_delayed_64__123_,
  chained_data_delayed_64__122_,chained_data_delayed_64__121_,chained_data_delayed_64__120_,
  chained_data_delayed_64__119_,chained_data_delayed_64__118_,chained_data_delayed_64__117_,
  chained_data_delayed_64__116_,chained_data_delayed_64__115_,
  chained_data_delayed_64__114_,chained_data_delayed_64__113_,chained_data_delayed_64__112_,
  chained_data_delayed_64__111_,chained_data_delayed_64__110_,chained_data_delayed_64__109_,
  chained_data_delayed_64__108_,chained_data_delayed_64__107_,
  chained_data_delayed_64__106_,chained_data_delayed_64__105_,chained_data_delayed_64__104_,
  chained_data_delayed_64__103_,chained_data_delayed_64__102_,chained_data_delayed_64__101_,
  chained_data_delayed_64__100_,chained_data_delayed_64__99_,chained_data_delayed_64__98_,
  chained_data_delayed_64__97_,chained_data_delayed_64__96_,
  chained_data_delayed_64__95_,chained_data_delayed_64__94_,chained_data_delayed_64__93_,
  chained_data_delayed_64__92_,chained_data_delayed_64__91_,chained_data_delayed_64__90_,
  chained_data_delayed_64__89_,chained_data_delayed_64__88_,chained_data_delayed_64__87_,
  chained_data_delayed_64__86_,chained_data_delayed_64__85_,
  chained_data_delayed_64__84_,chained_data_delayed_64__83_,chained_data_delayed_64__82_,
  chained_data_delayed_64__81_,chained_data_delayed_64__80_,chained_data_delayed_64__79_,
  chained_data_delayed_64__78_,chained_data_delayed_64__77_,chained_data_delayed_64__76_,
  chained_data_delayed_64__75_,chained_data_delayed_64__74_,
  chained_data_delayed_64__73_,chained_data_delayed_64__72_,chained_data_delayed_64__71_,
  chained_data_delayed_64__70_,chained_data_delayed_64__69_,chained_data_delayed_64__68_,
  chained_data_delayed_64__67_,chained_data_delayed_64__66_,chained_data_delayed_64__65_,
  chained_data_delayed_64__64_,chained_data_delayed_64__63_,
  chained_data_delayed_64__62_,chained_data_delayed_64__61_,chained_data_delayed_64__60_,
  chained_data_delayed_64__59_,chained_data_delayed_64__58_,chained_data_delayed_64__57_,
  chained_data_delayed_64__56_,chained_data_delayed_64__55_,chained_data_delayed_64__54_,
  chained_data_delayed_64__53_,chained_data_delayed_64__52_,
  chained_data_delayed_64__51_,chained_data_delayed_64__50_,chained_data_delayed_64__49_,
  chained_data_delayed_64__48_,chained_data_delayed_64__47_,chained_data_delayed_64__46_,
  chained_data_delayed_64__45_,chained_data_delayed_64__44_,chained_data_delayed_64__43_,
  chained_data_delayed_64__42_,chained_data_delayed_64__41_,
  chained_data_delayed_64__40_,chained_data_delayed_64__39_,chained_data_delayed_64__38_,
  chained_data_delayed_64__37_,chained_data_delayed_64__36_,chained_data_delayed_64__35_,
  chained_data_delayed_64__34_,chained_data_delayed_64__33_,chained_data_delayed_64__32_,
  chained_data_delayed_64__31_,chained_data_delayed_64__30_,
  chained_data_delayed_64__29_,chained_data_delayed_64__28_,chained_data_delayed_64__27_,
  chained_data_delayed_64__26_,chained_data_delayed_64__25_,chained_data_delayed_64__24_,
  chained_data_delayed_64__23_,chained_data_delayed_64__22_,chained_data_delayed_64__21_,
  chained_data_delayed_64__20_,chained_data_delayed_64__19_,chained_data_delayed_64__18_,
  chained_data_delayed_64__17_,chained_data_delayed_64__16_,
  chained_data_delayed_64__15_,chained_data_delayed_64__14_,chained_data_delayed_64__13_,
  chained_data_delayed_64__12_,chained_data_delayed_64__11_,chained_data_delayed_64__10_,
  chained_data_delayed_64__9_,chained_data_delayed_64__8_,chained_data_delayed_64__7_,
  chained_data_delayed_64__6_,chained_data_delayed_64__5_,chained_data_delayed_64__4_,
  chained_data_delayed_64__3_,chained_data_delayed_64__2_,
  chained_data_delayed_64__1_,chained_data_delayed_64__0_,chained_data_delayed_63__127_,
  chained_data_delayed_63__126_,chained_data_delayed_63__125_,chained_data_delayed_63__124_,
  chained_data_delayed_63__123_,chained_data_delayed_63__122_,
  chained_data_delayed_63__121_,chained_data_delayed_63__120_,chained_data_delayed_63__119_,
  chained_data_delayed_63__118_,chained_data_delayed_63__117_,chained_data_delayed_63__116_,
  chained_data_delayed_63__115_,chained_data_delayed_63__114_,
  chained_data_delayed_63__113_,chained_data_delayed_63__112_,chained_data_delayed_63__111_,
  chained_data_delayed_63__110_,chained_data_delayed_63__109_,chained_data_delayed_63__108_,
  chained_data_delayed_63__107_,chained_data_delayed_63__106_,
  chained_data_delayed_63__105_,chained_data_delayed_63__104_,chained_data_delayed_63__103_,
  chained_data_delayed_63__102_,chained_data_delayed_63__101_,chained_data_delayed_63__100_,
  chained_data_delayed_63__99_,chained_data_delayed_63__98_,chained_data_delayed_63__97_,
  chained_data_delayed_63__96_,chained_data_delayed_63__95_,
  chained_data_delayed_63__94_,chained_data_delayed_63__93_,chained_data_delayed_63__92_,
  chained_data_delayed_63__91_,chained_data_delayed_63__90_,chained_data_delayed_63__89_,
  chained_data_delayed_63__88_,chained_data_delayed_63__87_,chained_data_delayed_63__86_,
  chained_data_delayed_63__85_,chained_data_delayed_63__84_,
  chained_data_delayed_63__83_,chained_data_delayed_63__82_,chained_data_delayed_63__81_,
  chained_data_delayed_63__80_,chained_data_delayed_63__79_,chained_data_delayed_63__78_,
  chained_data_delayed_63__77_,chained_data_delayed_63__76_,chained_data_delayed_63__75_,
  chained_data_delayed_63__74_,chained_data_delayed_63__73_,
  chained_data_delayed_63__72_,chained_data_delayed_63__71_,chained_data_delayed_63__70_,
  chained_data_delayed_63__69_,chained_data_delayed_63__68_,chained_data_delayed_63__67_,
  chained_data_delayed_63__66_,chained_data_delayed_63__65_,chained_data_delayed_63__64_,
  chained_data_delayed_63__63_,chained_data_delayed_63__62_,
  chained_data_delayed_63__61_,chained_data_delayed_63__60_,chained_data_delayed_63__59_,
  chained_data_delayed_63__58_,chained_data_delayed_63__57_,chained_data_delayed_63__56_,
  chained_data_delayed_63__55_,chained_data_delayed_63__54_,chained_data_delayed_63__53_,
  chained_data_delayed_63__52_,chained_data_delayed_63__51_,
  chained_data_delayed_63__50_,chained_data_delayed_63__49_,chained_data_delayed_63__48_,
  chained_data_delayed_63__47_,chained_data_delayed_63__46_,chained_data_delayed_63__45_,
  chained_data_delayed_63__44_,chained_data_delayed_63__43_,chained_data_delayed_63__42_,
  chained_data_delayed_63__41_,chained_data_delayed_63__40_,
  chained_data_delayed_63__39_,chained_data_delayed_63__38_,chained_data_delayed_63__37_,
  chained_data_delayed_63__36_,chained_data_delayed_63__35_,chained_data_delayed_63__34_,
  chained_data_delayed_63__33_,chained_data_delayed_63__32_,chained_data_delayed_63__31_,
  chained_data_delayed_63__30_,chained_data_delayed_63__29_,chained_data_delayed_63__28_,
  chained_data_delayed_63__27_,chained_data_delayed_63__26_,
  chained_data_delayed_63__25_,chained_data_delayed_63__24_,chained_data_delayed_63__23_,
  chained_data_delayed_63__22_,chained_data_delayed_63__21_,chained_data_delayed_63__20_,
  chained_data_delayed_63__19_,chained_data_delayed_63__18_,chained_data_delayed_63__17_,
  chained_data_delayed_63__16_,chained_data_delayed_63__15_,
  chained_data_delayed_63__14_,chained_data_delayed_63__13_,chained_data_delayed_63__12_,
  chained_data_delayed_63__11_,chained_data_delayed_63__10_,chained_data_delayed_63__9_,
  chained_data_delayed_63__8_,chained_data_delayed_63__7_,chained_data_delayed_63__6_,
  chained_data_delayed_63__5_,chained_data_delayed_63__4_,chained_data_delayed_63__3_,
  chained_data_delayed_63__2_,chained_data_delayed_63__1_,
  chained_data_delayed_63__0_,chained_data_delayed_62__127_,chained_data_delayed_62__126_,
  chained_data_delayed_62__125_,chained_data_delayed_62__124_,chained_data_delayed_62__123_,
  chained_data_delayed_62__122_,chained_data_delayed_62__121_,
  chained_data_delayed_62__120_,chained_data_delayed_62__119_,chained_data_delayed_62__118_,
  chained_data_delayed_62__117_,chained_data_delayed_62__116_,chained_data_delayed_62__115_,
  chained_data_delayed_62__114_,chained_data_delayed_62__113_,
  chained_data_delayed_62__112_,chained_data_delayed_62__111_,chained_data_delayed_62__110_,
  chained_data_delayed_62__109_,chained_data_delayed_62__108_,chained_data_delayed_62__107_,
  chained_data_delayed_62__106_,chained_data_delayed_62__105_,
  chained_data_delayed_62__104_,chained_data_delayed_62__103_,chained_data_delayed_62__102_,
  chained_data_delayed_62__101_,chained_data_delayed_62__100_,chained_data_delayed_62__99_,
  chained_data_delayed_62__98_,chained_data_delayed_62__97_,chained_data_delayed_62__96_,
  chained_data_delayed_62__95_,chained_data_delayed_62__94_,
  chained_data_delayed_62__93_,chained_data_delayed_62__92_,chained_data_delayed_62__91_,
  chained_data_delayed_62__90_,chained_data_delayed_62__89_,chained_data_delayed_62__88_,
  chained_data_delayed_62__87_,chained_data_delayed_62__86_,chained_data_delayed_62__85_,
  chained_data_delayed_62__84_,chained_data_delayed_62__83_,
  chained_data_delayed_62__82_,chained_data_delayed_62__81_,chained_data_delayed_62__80_,
  chained_data_delayed_62__79_,chained_data_delayed_62__78_,chained_data_delayed_62__77_,
  chained_data_delayed_62__76_,chained_data_delayed_62__75_,chained_data_delayed_62__74_,
  chained_data_delayed_62__73_,chained_data_delayed_62__72_,
  chained_data_delayed_62__71_,chained_data_delayed_62__70_,chained_data_delayed_62__69_,
  chained_data_delayed_62__68_,chained_data_delayed_62__67_,chained_data_delayed_62__66_,
  chained_data_delayed_62__65_,chained_data_delayed_62__64_,chained_data_delayed_62__63_,
  chained_data_delayed_62__62_,chained_data_delayed_62__61_,
  chained_data_delayed_62__60_,chained_data_delayed_62__59_,chained_data_delayed_62__58_,
  chained_data_delayed_62__57_,chained_data_delayed_62__56_,chained_data_delayed_62__55_,
  chained_data_delayed_62__54_,chained_data_delayed_62__53_,chained_data_delayed_62__52_,
  chained_data_delayed_62__51_,chained_data_delayed_62__50_,
  chained_data_delayed_62__49_,chained_data_delayed_62__48_,chained_data_delayed_62__47_,
  chained_data_delayed_62__46_,chained_data_delayed_62__45_,chained_data_delayed_62__44_,
  chained_data_delayed_62__43_,chained_data_delayed_62__42_,chained_data_delayed_62__41_,
  chained_data_delayed_62__40_,chained_data_delayed_62__39_,chained_data_delayed_62__38_,
  chained_data_delayed_62__37_,chained_data_delayed_62__36_,
  chained_data_delayed_62__35_,chained_data_delayed_62__34_,chained_data_delayed_62__33_,
  chained_data_delayed_62__32_,chained_data_delayed_62__31_,chained_data_delayed_62__30_,
  chained_data_delayed_62__29_,chained_data_delayed_62__28_,chained_data_delayed_62__27_,
  chained_data_delayed_62__26_,chained_data_delayed_62__25_,
  chained_data_delayed_62__24_,chained_data_delayed_62__23_,chained_data_delayed_62__22_,
  chained_data_delayed_62__21_,chained_data_delayed_62__20_,chained_data_delayed_62__19_,
  chained_data_delayed_62__18_,chained_data_delayed_62__17_,chained_data_delayed_62__16_,
  chained_data_delayed_62__15_,chained_data_delayed_62__14_,
  chained_data_delayed_62__13_,chained_data_delayed_62__12_,chained_data_delayed_62__11_,
  chained_data_delayed_62__10_,chained_data_delayed_62__9_,chained_data_delayed_62__8_,
  chained_data_delayed_62__7_,chained_data_delayed_62__6_,chained_data_delayed_62__5_,
  chained_data_delayed_62__4_,chained_data_delayed_62__3_,chained_data_delayed_62__2_,
  chained_data_delayed_62__1_,chained_data_delayed_62__0_,
  chained_data_delayed_61__127_,chained_data_delayed_61__126_,chained_data_delayed_61__125_,
  chained_data_delayed_61__124_,chained_data_delayed_61__123_,chained_data_delayed_61__122_,
  chained_data_delayed_61__121_,chained_data_delayed_61__120_,
  chained_data_delayed_61__119_,chained_data_delayed_61__118_,chained_data_delayed_61__117_,
  chained_data_delayed_61__116_,chained_data_delayed_61__115_,chained_data_delayed_61__114_,
  chained_data_delayed_61__113_,chained_data_delayed_61__112_,
  chained_data_delayed_61__111_,chained_data_delayed_61__110_,chained_data_delayed_61__109_,
  chained_data_delayed_61__108_,chained_data_delayed_61__107_,chained_data_delayed_61__106_,
  chained_data_delayed_61__105_,chained_data_delayed_61__104_,
  chained_data_delayed_61__103_,chained_data_delayed_61__102_,chained_data_delayed_61__101_,
  chained_data_delayed_61__100_,chained_data_delayed_61__99_,chained_data_delayed_61__98_,
  chained_data_delayed_61__97_,chained_data_delayed_61__96_,chained_data_delayed_61__95_,
  chained_data_delayed_61__94_,chained_data_delayed_61__93_,
  chained_data_delayed_61__92_,chained_data_delayed_61__91_,chained_data_delayed_61__90_,
  chained_data_delayed_61__89_,chained_data_delayed_61__88_,chained_data_delayed_61__87_,
  chained_data_delayed_61__86_,chained_data_delayed_61__85_,chained_data_delayed_61__84_,
  chained_data_delayed_61__83_,chained_data_delayed_61__82_,
  chained_data_delayed_61__81_,chained_data_delayed_61__80_,chained_data_delayed_61__79_,
  chained_data_delayed_61__78_,chained_data_delayed_61__77_,chained_data_delayed_61__76_,
  chained_data_delayed_61__75_,chained_data_delayed_61__74_,chained_data_delayed_61__73_,
  chained_data_delayed_61__72_,chained_data_delayed_61__71_,
  chained_data_delayed_61__70_,chained_data_delayed_61__69_,chained_data_delayed_61__68_,
  chained_data_delayed_61__67_,chained_data_delayed_61__66_,chained_data_delayed_61__65_,
  chained_data_delayed_61__64_,chained_data_delayed_61__63_,chained_data_delayed_61__62_,
  chained_data_delayed_61__61_,chained_data_delayed_61__60_,
  chained_data_delayed_61__59_,chained_data_delayed_61__58_,chained_data_delayed_61__57_,
  chained_data_delayed_61__56_,chained_data_delayed_61__55_,chained_data_delayed_61__54_,
  chained_data_delayed_61__53_,chained_data_delayed_61__52_,chained_data_delayed_61__51_,
  chained_data_delayed_61__50_,chained_data_delayed_61__49_,chained_data_delayed_61__48_,
  chained_data_delayed_61__47_,chained_data_delayed_61__46_,
  chained_data_delayed_61__45_,chained_data_delayed_61__44_,chained_data_delayed_61__43_,
  chained_data_delayed_61__42_,chained_data_delayed_61__41_,chained_data_delayed_61__40_,
  chained_data_delayed_61__39_,chained_data_delayed_61__38_,chained_data_delayed_61__37_,
  chained_data_delayed_61__36_,chained_data_delayed_61__35_,
  chained_data_delayed_61__34_,chained_data_delayed_61__33_,chained_data_delayed_61__32_,
  chained_data_delayed_61__31_,chained_data_delayed_61__30_,chained_data_delayed_61__29_,
  chained_data_delayed_61__28_,chained_data_delayed_61__27_,chained_data_delayed_61__26_,
  chained_data_delayed_61__25_,chained_data_delayed_61__24_,
  chained_data_delayed_61__23_,chained_data_delayed_61__22_,chained_data_delayed_61__21_,
  chained_data_delayed_61__20_,chained_data_delayed_61__19_,chained_data_delayed_61__18_,
  chained_data_delayed_61__17_,chained_data_delayed_61__16_,chained_data_delayed_61__15_,
  chained_data_delayed_61__14_,chained_data_delayed_61__13_,
  chained_data_delayed_61__12_,chained_data_delayed_61__11_,chained_data_delayed_61__10_,
  chained_data_delayed_61__9_,chained_data_delayed_61__8_,chained_data_delayed_61__7_,
  chained_data_delayed_61__6_,chained_data_delayed_61__5_,chained_data_delayed_61__4_,
  chained_data_delayed_61__3_,chained_data_delayed_61__2_,chained_data_delayed_61__1_,
  chained_data_delayed_61__0_,chained_data_delayed_68__127_,
  chained_data_delayed_68__126_,chained_data_delayed_68__125_,chained_data_delayed_68__124_,
  chained_data_delayed_68__123_,chained_data_delayed_68__122_,chained_data_delayed_68__121_,
  chained_data_delayed_68__120_,chained_data_delayed_68__119_,
  chained_data_delayed_68__118_,chained_data_delayed_68__117_,chained_data_delayed_68__116_,
  chained_data_delayed_68__115_,chained_data_delayed_68__114_,chained_data_delayed_68__113_,
  chained_data_delayed_68__112_,chained_data_delayed_68__111_,
  chained_data_delayed_68__110_,chained_data_delayed_68__109_,chained_data_delayed_68__108_,
  chained_data_delayed_68__107_,chained_data_delayed_68__106_,chained_data_delayed_68__105_,
  chained_data_delayed_68__104_,chained_data_delayed_68__103_,
  chained_data_delayed_68__102_,chained_data_delayed_68__101_,chained_data_delayed_68__100_,
  chained_data_delayed_68__99_,chained_data_delayed_68__98_,chained_data_delayed_68__97_,
  chained_data_delayed_68__96_,chained_data_delayed_68__95_,chained_data_delayed_68__94_,
  chained_data_delayed_68__93_,chained_data_delayed_68__92_,
  chained_data_delayed_68__91_,chained_data_delayed_68__90_,chained_data_delayed_68__89_,
  chained_data_delayed_68__88_,chained_data_delayed_68__87_,chained_data_delayed_68__86_,
  chained_data_delayed_68__85_,chained_data_delayed_68__84_,chained_data_delayed_68__83_,
  chained_data_delayed_68__82_,chained_data_delayed_68__81_,
  chained_data_delayed_68__80_,chained_data_delayed_68__79_,chained_data_delayed_68__78_,
  chained_data_delayed_68__77_,chained_data_delayed_68__76_,chained_data_delayed_68__75_,
  chained_data_delayed_68__74_,chained_data_delayed_68__73_,chained_data_delayed_68__72_,
  chained_data_delayed_68__71_,chained_data_delayed_68__70_,
  chained_data_delayed_68__69_,chained_data_delayed_68__68_,chained_data_delayed_68__67_,
  chained_data_delayed_68__66_,chained_data_delayed_68__65_,chained_data_delayed_68__64_,
  chained_data_delayed_68__63_,chained_data_delayed_68__62_,chained_data_delayed_68__61_,
  chained_data_delayed_68__60_,chained_data_delayed_68__59_,chained_data_delayed_68__58_,
  chained_data_delayed_68__57_,chained_data_delayed_68__56_,
  chained_data_delayed_68__55_,chained_data_delayed_68__54_,chained_data_delayed_68__53_,
  chained_data_delayed_68__52_,chained_data_delayed_68__51_,chained_data_delayed_68__50_,
  chained_data_delayed_68__49_,chained_data_delayed_68__48_,chained_data_delayed_68__47_,
  chained_data_delayed_68__46_,chained_data_delayed_68__45_,
  chained_data_delayed_68__44_,chained_data_delayed_68__43_,chained_data_delayed_68__42_,
  chained_data_delayed_68__41_,chained_data_delayed_68__40_,chained_data_delayed_68__39_,
  chained_data_delayed_68__38_,chained_data_delayed_68__37_,chained_data_delayed_68__36_,
  chained_data_delayed_68__35_,chained_data_delayed_68__34_,
  chained_data_delayed_68__33_,chained_data_delayed_68__32_,chained_data_delayed_68__31_,
  chained_data_delayed_68__30_,chained_data_delayed_68__29_,chained_data_delayed_68__28_,
  chained_data_delayed_68__27_,chained_data_delayed_68__26_,chained_data_delayed_68__25_,
  chained_data_delayed_68__24_,chained_data_delayed_68__23_,
  chained_data_delayed_68__22_,chained_data_delayed_68__21_,chained_data_delayed_68__20_,
  chained_data_delayed_68__19_,chained_data_delayed_68__18_,chained_data_delayed_68__17_,
  chained_data_delayed_68__16_,chained_data_delayed_68__15_,chained_data_delayed_68__14_,
  chained_data_delayed_68__13_,chained_data_delayed_68__12_,
  chained_data_delayed_68__11_,chained_data_delayed_68__10_,chained_data_delayed_68__9_,
  chained_data_delayed_68__8_,chained_data_delayed_68__7_,chained_data_delayed_68__6_,
  chained_data_delayed_68__5_,chained_data_delayed_68__4_,chained_data_delayed_68__3_,
  chained_data_delayed_68__2_,chained_data_delayed_68__1_,chained_data_delayed_68__0_,
  chained_data_delayed_67__127_,chained_data_delayed_67__126_,
  chained_data_delayed_67__125_,chained_data_delayed_67__124_,chained_data_delayed_67__123_,
  chained_data_delayed_67__122_,chained_data_delayed_67__121_,chained_data_delayed_67__120_,
  chained_data_delayed_67__119_,chained_data_delayed_67__118_,
  chained_data_delayed_67__117_,chained_data_delayed_67__116_,chained_data_delayed_67__115_,
  chained_data_delayed_67__114_,chained_data_delayed_67__113_,chained_data_delayed_67__112_,
  chained_data_delayed_67__111_,chained_data_delayed_67__110_,
  chained_data_delayed_67__109_,chained_data_delayed_67__108_,chained_data_delayed_67__107_,
  chained_data_delayed_67__106_,chained_data_delayed_67__105_,chained_data_delayed_67__104_,
  chained_data_delayed_67__103_,chained_data_delayed_67__102_,
  chained_data_delayed_67__101_,chained_data_delayed_67__100_,chained_data_delayed_67__99_,
  chained_data_delayed_67__98_,chained_data_delayed_67__97_,chained_data_delayed_67__96_,
  chained_data_delayed_67__95_,chained_data_delayed_67__94_,chained_data_delayed_67__93_,
  chained_data_delayed_67__92_,chained_data_delayed_67__91_,
  chained_data_delayed_67__90_,chained_data_delayed_67__89_,chained_data_delayed_67__88_,
  chained_data_delayed_67__87_,chained_data_delayed_67__86_,chained_data_delayed_67__85_,
  chained_data_delayed_67__84_,chained_data_delayed_67__83_,chained_data_delayed_67__82_,
  chained_data_delayed_67__81_,chained_data_delayed_67__80_,
  chained_data_delayed_67__79_,chained_data_delayed_67__78_,chained_data_delayed_67__77_,
  chained_data_delayed_67__76_,chained_data_delayed_67__75_,chained_data_delayed_67__74_,
  chained_data_delayed_67__73_,chained_data_delayed_67__72_,chained_data_delayed_67__71_,
  chained_data_delayed_67__70_,chained_data_delayed_67__69_,chained_data_delayed_67__68_,
  chained_data_delayed_67__67_,chained_data_delayed_67__66_,
  chained_data_delayed_67__65_,chained_data_delayed_67__64_,chained_data_delayed_67__63_,
  chained_data_delayed_67__62_,chained_data_delayed_67__61_,chained_data_delayed_67__60_,
  chained_data_delayed_67__59_,chained_data_delayed_67__58_,chained_data_delayed_67__57_,
  chained_data_delayed_67__56_,chained_data_delayed_67__55_,
  chained_data_delayed_67__54_,chained_data_delayed_67__53_,chained_data_delayed_67__52_,
  chained_data_delayed_67__51_,chained_data_delayed_67__50_,chained_data_delayed_67__49_,
  chained_data_delayed_67__48_,chained_data_delayed_67__47_,chained_data_delayed_67__46_,
  chained_data_delayed_67__45_,chained_data_delayed_67__44_,
  chained_data_delayed_67__43_,chained_data_delayed_67__42_,chained_data_delayed_67__41_,
  chained_data_delayed_67__40_,chained_data_delayed_67__39_,chained_data_delayed_67__38_,
  chained_data_delayed_67__37_,chained_data_delayed_67__36_,chained_data_delayed_67__35_,
  chained_data_delayed_67__34_,chained_data_delayed_67__33_,
  chained_data_delayed_67__32_,chained_data_delayed_67__31_,chained_data_delayed_67__30_,
  chained_data_delayed_67__29_,chained_data_delayed_67__28_,chained_data_delayed_67__27_,
  chained_data_delayed_67__26_,chained_data_delayed_67__25_,chained_data_delayed_67__24_,
  chained_data_delayed_67__23_,chained_data_delayed_67__22_,
  chained_data_delayed_67__21_,chained_data_delayed_67__20_,chained_data_delayed_67__19_,
  chained_data_delayed_67__18_,chained_data_delayed_67__17_,chained_data_delayed_67__16_,
  chained_data_delayed_67__15_,chained_data_delayed_67__14_,chained_data_delayed_67__13_,
  chained_data_delayed_67__12_,chained_data_delayed_67__11_,
  chained_data_delayed_67__10_,chained_data_delayed_67__9_,chained_data_delayed_67__8_,
  chained_data_delayed_67__7_,chained_data_delayed_67__6_,chained_data_delayed_67__5_,
  chained_data_delayed_67__4_,chained_data_delayed_67__3_,chained_data_delayed_67__2_,
  chained_data_delayed_67__1_,chained_data_delayed_67__0_,chained_data_delayed_66__127_,
  chained_data_delayed_66__126_,chained_data_delayed_66__125_,
  chained_data_delayed_66__124_,chained_data_delayed_66__123_,chained_data_delayed_66__122_,
  chained_data_delayed_66__121_,chained_data_delayed_66__120_,chained_data_delayed_66__119_,
  chained_data_delayed_66__118_,chained_data_delayed_66__117_,
  chained_data_delayed_66__116_,chained_data_delayed_66__115_,chained_data_delayed_66__114_,
  chained_data_delayed_66__113_,chained_data_delayed_66__112_,chained_data_delayed_66__111_,
  chained_data_delayed_66__110_,chained_data_delayed_66__109_,
  chained_data_delayed_66__108_,chained_data_delayed_66__107_,chained_data_delayed_66__106_,
  chained_data_delayed_66__105_,chained_data_delayed_66__104_,chained_data_delayed_66__103_,
  chained_data_delayed_66__102_,chained_data_delayed_66__101_,
  chained_data_delayed_66__100_,chained_data_delayed_66__99_,chained_data_delayed_66__98_,
  chained_data_delayed_66__97_,chained_data_delayed_66__96_,chained_data_delayed_66__95_,
  chained_data_delayed_66__94_,chained_data_delayed_66__93_,chained_data_delayed_66__92_,
  chained_data_delayed_66__91_,chained_data_delayed_66__90_,
  chained_data_delayed_66__89_,chained_data_delayed_66__88_,chained_data_delayed_66__87_,
  chained_data_delayed_66__86_,chained_data_delayed_66__85_,chained_data_delayed_66__84_,
  chained_data_delayed_66__83_,chained_data_delayed_66__82_,chained_data_delayed_66__81_,
  chained_data_delayed_66__80_,chained_data_delayed_66__79_,chained_data_delayed_66__78_,
  chained_data_delayed_66__77_,chained_data_delayed_66__76_,
  chained_data_delayed_66__75_,chained_data_delayed_66__74_,chained_data_delayed_66__73_,
  chained_data_delayed_66__72_,chained_data_delayed_66__71_,chained_data_delayed_66__70_,
  chained_data_delayed_66__69_,chained_data_delayed_66__68_,chained_data_delayed_66__67_,
  chained_data_delayed_66__66_,chained_data_delayed_66__65_,
  chained_data_delayed_66__64_,chained_data_delayed_66__63_,chained_data_delayed_66__62_,
  chained_data_delayed_66__61_,chained_data_delayed_66__60_,chained_data_delayed_66__59_,
  chained_data_delayed_66__58_,chained_data_delayed_66__57_,chained_data_delayed_66__56_,
  chained_data_delayed_66__55_,chained_data_delayed_66__54_,
  chained_data_delayed_66__53_,chained_data_delayed_66__52_,chained_data_delayed_66__51_,
  chained_data_delayed_66__50_,chained_data_delayed_66__49_,chained_data_delayed_66__48_,
  chained_data_delayed_66__47_,chained_data_delayed_66__46_,chained_data_delayed_66__45_,
  chained_data_delayed_66__44_,chained_data_delayed_66__43_,
  chained_data_delayed_66__42_,chained_data_delayed_66__41_,chained_data_delayed_66__40_,
  chained_data_delayed_66__39_,chained_data_delayed_66__38_,chained_data_delayed_66__37_,
  chained_data_delayed_66__36_,chained_data_delayed_66__35_,chained_data_delayed_66__34_,
  chained_data_delayed_66__33_,chained_data_delayed_66__32_,
  chained_data_delayed_66__31_,chained_data_delayed_66__30_,chained_data_delayed_66__29_,
  chained_data_delayed_66__28_,chained_data_delayed_66__27_,chained_data_delayed_66__26_,
  chained_data_delayed_66__25_,chained_data_delayed_66__24_,chained_data_delayed_66__23_,
  chained_data_delayed_66__22_,chained_data_delayed_66__21_,
  chained_data_delayed_66__20_,chained_data_delayed_66__19_,chained_data_delayed_66__18_,
  chained_data_delayed_66__17_,chained_data_delayed_66__16_,chained_data_delayed_66__15_,
  chained_data_delayed_66__14_,chained_data_delayed_66__13_,chained_data_delayed_66__12_,
  chained_data_delayed_66__11_,chained_data_delayed_66__10_,chained_data_delayed_66__9_,
  chained_data_delayed_66__8_,chained_data_delayed_66__7_,
  chained_data_delayed_66__6_,chained_data_delayed_66__5_,chained_data_delayed_66__4_,
  chained_data_delayed_66__3_,chained_data_delayed_66__2_,chained_data_delayed_66__1_,
  chained_data_delayed_66__0_,chained_data_delayed_65__127_,chained_data_delayed_65__126_,
  chained_data_delayed_65__125_,chained_data_delayed_65__124_,
  chained_data_delayed_65__123_,chained_data_delayed_65__122_,chained_data_delayed_65__121_,
  chained_data_delayed_65__120_,chained_data_delayed_65__119_,chained_data_delayed_65__118_,
  chained_data_delayed_65__117_,chained_data_delayed_65__116_,
  chained_data_delayed_65__115_,chained_data_delayed_65__114_,chained_data_delayed_65__113_,
  chained_data_delayed_65__112_,chained_data_delayed_65__111_,chained_data_delayed_65__110_,
  chained_data_delayed_65__109_,chained_data_delayed_65__108_,
  chained_data_delayed_65__107_,chained_data_delayed_65__106_,chained_data_delayed_65__105_,
  chained_data_delayed_65__104_,chained_data_delayed_65__103_,chained_data_delayed_65__102_,
  chained_data_delayed_65__101_,chained_data_delayed_65__100_,
  chained_data_delayed_65__99_,chained_data_delayed_65__98_,chained_data_delayed_65__97_,
  chained_data_delayed_65__96_,chained_data_delayed_65__95_,chained_data_delayed_65__94_,
  chained_data_delayed_65__93_,chained_data_delayed_65__92_,chained_data_delayed_65__91_,
  chained_data_delayed_65__90_,chained_data_delayed_65__89_,chained_data_delayed_65__88_,
  chained_data_delayed_65__87_,chained_data_delayed_65__86_,
  chained_data_delayed_65__85_,chained_data_delayed_65__84_,chained_data_delayed_65__83_,
  chained_data_delayed_65__82_,chained_data_delayed_65__81_,chained_data_delayed_65__80_,
  chained_data_delayed_65__79_,chained_data_delayed_65__78_,chained_data_delayed_65__77_,
  chained_data_delayed_65__76_,chained_data_delayed_65__75_,
  chained_data_delayed_65__74_,chained_data_delayed_65__73_,chained_data_delayed_65__72_,
  chained_data_delayed_65__71_,chained_data_delayed_65__70_,chained_data_delayed_65__69_,
  chained_data_delayed_65__68_,chained_data_delayed_65__67_,chained_data_delayed_65__66_,
  chained_data_delayed_65__65_,chained_data_delayed_65__64_,
  chained_data_delayed_65__63_,chained_data_delayed_65__62_,chained_data_delayed_65__61_,
  chained_data_delayed_65__60_,chained_data_delayed_65__59_,chained_data_delayed_65__58_,
  chained_data_delayed_65__57_,chained_data_delayed_65__56_,chained_data_delayed_65__55_,
  chained_data_delayed_65__54_,chained_data_delayed_65__53_,
  chained_data_delayed_65__52_,chained_data_delayed_65__51_,chained_data_delayed_65__50_,
  chained_data_delayed_65__49_,chained_data_delayed_65__48_,chained_data_delayed_65__47_,
  chained_data_delayed_65__46_,chained_data_delayed_65__45_,chained_data_delayed_65__44_,
  chained_data_delayed_65__43_,chained_data_delayed_65__42_,
  chained_data_delayed_65__41_,chained_data_delayed_65__40_,chained_data_delayed_65__39_,
  chained_data_delayed_65__38_,chained_data_delayed_65__37_,chained_data_delayed_65__36_,
  chained_data_delayed_65__35_,chained_data_delayed_65__34_,chained_data_delayed_65__33_,
  chained_data_delayed_65__32_,chained_data_delayed_65__31_,
  chained_data_delayed_65__30_,chained_data_delayed_65__29_,chained_data_delayed_65__28_,
  chained_data_delayed_65__27_,chained_data_delayed_65__26_,chained_data_delayed_65__25_,
  chained_data_delayed_65__24_,chained_data_delayed_65__23_,chained_data_delayed_65__22_,
  chained_data_delayed_65__21_,chained_data_delayed_65__20_,
  chained_data_delayed_65__19_,chained_data_delayed_65__18_,chained_data_delayed_65__17_,
  chained_data_delayed_65__16_,chained_data_delayed_65__15_,chained_data_delayed_65__14_,
  chained_data_delayed_65__13_,chained_data_delayed_65__12_,chained_data_delayed_65__11_,
  chained_data_delayed_65__10_,chained_data_delayed_65__9_,chained_data_delayed_65__8_,
  chained_data_delayed_65__7_,chained_data_delayed_65__6_,
  chained_data_delayed_65__5_,chained_data_delayed_65__4_,chained_data_delayed_65__3_,
  chained_data_delayed_65__2_,chained_data_delayed_65__1_,chained_data_delayed_65__0_,
  chained_data_delayed_72__127_,chained_data_delayed_72__126_,chained_data_delayed_72__125_,
  chained_data_delayed_72__124_,chained_data_delayed_72__123_,
  chained_data_delayed_72__122_,chained_data_delayed_72__121_,chained_data_delayed_72__120_,
  chained_data_delayed_72__119_,chained_data_delayed_72__118_,chained_data_delayed_72__117_,
  chained_data_delayed_72__116_,chained_data_delayed_72__115_,
  chained_data_delayed_72__114_,chained_data_delayed_72__113_,chained_data_delayed_72__112_,
  chained_data_delayed_72__111_,chained_data_delayed_72__110_,chained_data_delayed_72__109_,
  chained_data_delayed_72__108_,chained_data_delayed_72__107_,
  chained_data_delayed_72__106_,chained_data_delayed_72__105_,chained_data_delayed_72__104_,
  chained_data_delayed_72__103_,chained_data_delayed_72__102_,chained_data_delayed_72__101_,
  chained_data_delayed_72__100_,chained_data_delayed_72__99_,chained_data_delayed_72__98_,
  chained_data_delayed_72__97_,chained_data_delayed_72__96_,
  chained_data_delayed_72__95_,chained_data_delayed_72__94_,chained_data_delayed_72__93_,
  chained_data_delayed_72__92_,chained_data_delayed_72__91_,chained_data_delayed_72__90_,
  chained_data_delayed_72__89_,chained_data_delayed_72__88_,chained_data_delayed_72__87_,
  chained_data_delayed_72__86_,chained_data_delayed_72__85_,
  chained_data_delayed_72__84_,chained_data_delayed_72__83_,chained_data_delayed_72__82_,
  chained_data_delayed_72__81_,chained_data_delayed_72__80_,chained_data_delayed_72__79_,
  chained_data_delayed_72__78_,chained_data_delayed_72__77_,chained_data_delayed_72__76_,
  chained_data_delayed_72__75_,chained_data_delayed_72__74_,
  chained_data_delayed_72__73_,chained_data_delayed_72__72_,chained_data_delayed_72__71_,
  chained_data_delayed_72__70_,chained_data_delayed_72__69_,chained_data_delayed_72__68_,
  chained_data_delayed_72__67_,chained_data_delayed_72__66_,chained_data_delayed_72__65_,
  chained_data_delayed_72__64_,chained_data_delayed_72__63_,
  chained_data_delayed_72__62_,chained_data_delayed_72__61_,chained_data_delayed_72__60_,
  chained_data_delayed_72__59_,chained_data_delayed_72__58_,chained_data_delayed_72__57_,
  chained_data_delayed_72__56_,chained_data_delayed_72__55_,chained_data_delayed_72__54_,
  chained_data_delayed_72__53_,chained_data_delayed_72__52_,
  chained_data_delayed_72__51_,chained_data_delayed_72__50_,chained_data_delayed_72__49_,
  chained_data_delayed_72__48_,chained_data_delayed_72__47_,chained_data_delayed_72__46_,
  chained_data_delayed_72__45_,chained_data_delayed_72__44_,chained_data_delayed_72__43_,
  chained_data_delayed_72__42_,chained_data_delayed_72__41_,
  chained_data_delayed_72__40_,chained_data_delayed_72__39_,chained_data_delayed_72__38_,
  chained_data_delayed_72__37_,chained_data_delayed_72__36_,chained_data_delayed_72__35_,
  chained_data_delayed_72__34_,chained_data_delayed_72__33_,chained_data_delayed_72__32_,
  chained_data_delayed_72__31_,chained_data_delayed_72__30_,
  chained_data_delayed_72__29_,chained_data_delayed_72__28_,chained_data_delayed_72__27_,
  chained_data_delayed_72__26_,chained_data_delayed_72__25_,chained_data_delayed_72__24_,
  chained_data_delayed_72__23_,chained_data_delayed_72__22_,chained_data_delayed_72__21_,
  chained_data_delayed_72__20_,chained_data_delayed_72__19_,chained_data_delayed_72__18_,
  chained_data_delayed_72__17_,chained_data_delayed_72__16_,
  chained_data_delayed_72__15_,chained_data_delayed_72__14_,chained_data_delayed_72__13_,
  chained_data_delayed_72__12_,chained_data_delayed_72__11_,chained_data_delayed_72__10_,
  chained_data_delayed_72__9_,chained_data_delayed_72__8_,chained_data_delayed_72__7_,
  chained_data_delayed_72__6_,chained_data_delayed_72__5_,chained_data_delayed_72__4_,
  chained_data_delayed_72__3_,chained_data_delayed_72__2_,
  chained_data_delayed_72__1_,chained_data_delayed_72__0_,chained_data_delayed_71__127_,
  chained_data_delayed_71__126_,chained_data_delayed_71__125_,chained_data_delayed_71__124_,
  chained_data_delayed_71__123_,chained_data_delayed_71__122_,
  chained_data_delayed_71__121_,chained_data_delayed_71__120_,chained_data_delayed_71__119_,
  chained_data_delayed_71__118_,chained_data_delayed_71__117_,chained_data_delayed_71__116_,
  chained_data_delayed_71__115_,chained_data_delayed_71__114_,
  chained_data_delayed_71__113_,chained_data_delayed_71__112_,chained_data_delayed_71__111_,
  chained_data_delayed_71__110_,chained_data_delayed_71__109_,chained_data_delayed_71__108_,
  chained_data_delayed_71__107_,chained_data_delayed_71__106_,
  chained_data_delayed_71__105_,chained_data_delayed_71__104_,chained_data_delayed_71__103_,
  chained_data_delayed_71__102_,chained_data_delayed_71__101_,chained_data_delayed_71__100_,
  chained_data_delayed_71__99_,chained_data_delayed_71__98_,chained_data_delayed_71__97_,
  chained_data_delayed_71__96_,chained_data_delayed_71__95_,
  chained_data_delayed_71__94_,chained_data_delayed_71__93_,chained_data_delayed_71__92_,
  chained_data_delayed_71__91_,chained_data_delayed_71__90_,chained_data_delayed_71__89_,
  chained_data_delayed_71__88_,chained_data_delayed_71__87_,chained_data_delayed_71__86_,
  chained_data_delayed_71__85_,chained_data_delayed_71__84_,
  chained_data_delayed_71__83_,chained_data_delayed_71__82_,chained_data_delayed_71__81_,
  chained_data_delayed_71__80_,chained_data_delayed_71__79_,chained_data_delayed_71__78_,
  chained_data_delayed_71__77_,chained_data_delayed_71__76_,chained_data_delayed_71__75_,
  chained_data_delayed_71__74_,chained_data_delayed_71__73_,
  chained_data_delayed_71__72_,chained_data_delayed_71__71_,chained_data_delayed_71__70_,
  chained_data_delayed_71__69_,chained_data_delayed_71__68_,chained_data_delayed_71__67_,
  chained_data_delayed_71__66_,chained_data_delayed_71__65_,chained_data_delayed_71__64_,
  chained_data_delayed_71__63_,chained_data_delayed_71__62_,
  chained_data_delayed_71__61_,chained_data_delayed_71__60_,chained_data_delayed_71__59_,
  chained_data_delayed_71__58_,chained_data_delayed_71__57_,chained_data_delayed_71__56_,
  chained_data_delayed_71__55_,chained_data_delayed_71__54_,chained_data_delayed_71__53_,
  chained_data_delayed_71__52_,chained_data_delayed_71__51_,
  chained_data_delayed_71__50_,chained_data_delayed_71__49_,chained_data_delayed_71__48_,
  chained_data_delayed_71__47_,chained_data_delayed_71__46_,chained_data_delayed_71__45_,
  chained_data_delayed_71__44_,chained_data_delayed_71__43_,chained_data_delayed_71__42_,
  chained_data_delayed_71__41_,chained_data_delayed_71__40_,
  chained_data_delayed_71__39_,chained_data_delayed_71__38_,chained_data_delayed_71__37_,
  chained_data_delayed_71__36_,chained_data_delayed_71__35_,chained_data_delayed_71__34_,
  chained_data_delayed_71__33_,chained_data_delayed_71__32_,chained_data_delayed_71__31_,
  chained_data_delayed_71__30_,chained_data_delayed_71__29_,chained_data_delayed_71__28_,
  chained_data_delayed_71__27_,chained_data_delayed_71__26_,
  chained_data_delayed_71__25_,chained_data_delayed_71__24_,chained_data_delayed_71__23_,
  chained_data_delayed_71__22_,chained_data_delayed_71__21_,chained_data_delayed_71__20_,
  chained_data_delayed_71__19_,chained_data_delayed_71__18_,chained_data_delayed_71__17_,
  chained_data_delayed_71__16_,chained_data_delayed_71__15_,
  chained_data_delayed_71__14_,chained_data_delayed_71__13_,chained_data_delayed_71__12_,
  chained_data_delayed_71__11_,chained_data_delayed_71__10_,chained_data_delayed_71__9_,
  chained_data_delayed_71__8_,chained_data_delayed_71__7_,chained_data_delayed_71__6_,
  chained_data_delayed_71__5_,chained_data_delayed_71__4_,chained_data_delayed_71__3_,
  chained_data_delayed_71__2_,chained_data_delayed_71__1_,
  chained_data_delayed_71__0_,chained_data_delayed_70__127_,chained_data_delayed_70__126_,
  chained_data_delayed_70__125_,chained_data_delayed_70__124_,chained_data_delayed_70__123_,
  chained_data_delayed_70__122_,chained_data_delayed_70__121_,
  chained_data_delayed_70__120_,chained_data_delayed_70__119_,chained_data_delayed_70__118_,
  chained_data_delayed_70__117_,chained_data_delayed_70__116_,chained_data_delayed_70__115_,
  chained_data_delayed_70__114_,chained_data_delayed_70__113_,
  chained_data_delayed_70__112_,chained_data_delayed_70__111_,chained_data_delayed_70__110_,
  chained_data_delayed_70__109_,chained_data_delayed_70__108_,chained_data_delayed_70__107_,
  chained_data_delayed_70__106_,chained_data_delayed_70__105_,
  chained_data_delayed_70__104_,chained_data_delayed_70__103_,chained_data_delayed_70__102_,
  chained_data_delayed_70__101_,chained_data_delayed_70__100_,chained_data_delayed_70__99_,
  chained_data_delayed_70__98_,chained_data_delayed_70__97_,chained_data_delayed_70__96_,
  chained_data_delayed_70__95_,chained_data_delayed_70__94_,
  chained_data_delayed_70__93_,chained_data_delayed_70__92_,chained_data_delayed_70__91_,
  chained_data_delayed_70__90_,chained_data_delayed_70__89_,chained_data_delayed_70__88_,
  chained_data_delayed_70__87_,chained_data_delayed_70__86_,chained_data_delayed_70__85_,
  chained_data_delayed_70__84_,chained_data_delayed_70__83_,
  chained_data_delayed_70__82_,chained_data_delayed_70__81_,chained_data_delayed_70__80_,
  chained_data_delayed_70__79_,chained_data_delayed_70__78_,chained_data_delayed_70__77_,
  chained_data_delayed_70__76_,chained_data_delayed_70__75_,chained_data_delayed_70__74_,
  chained_data_delayed_70__73_,chained_data_delayed_70__72_,
  chained_data_delayed_70__71_,chained_data_delayed_70__70_,chained_data_delayed_70__69_,
  chained_data_delayed_70__68_,chained_data_delayed_70__67_,chained_data_delayed_70__66_,
  chained_data_delayed_70__65_,chained_data_delayed_70__64_,chained_data_delayed_70__63_,
  chained_data_delayed_70__62_,chained_data_delayed_70__61_,
  chained_data_delayed_70__60_,chained_data_delayed_70__59_,chained_data_delayed_70__58_,
  chained_data_delayed_70__57_,chained_data_delayed_70__56_,chained_data_delayed_70__55_,
  chained_data_delayed_70__54_,chained_data_delayed_70__53_,chained_data_delayed_70__52_,
  chained_data_delayed_70__51_,chained_data_delayed_70__50_,
  chained_data_delayed_70__49_,chained_data_delayed_70__48_,chained_data_delayed_70__47_,
  chained_data_delayed_70__46_,chained_data_delayed_70__45_,chained_data_delayed_70__44_,
  chained_data_delayed_70__43_,chained_data_delayed_70__42_,chained_data_delayed_70__41_,
  chained_data_delayed_70__40_,chained_data_delayed_70__39_,chained_data_delayed_70__38_,
  chained_data_delayed_70__37_,chained_data_delayed_70__36_,
  chained_data_delayed_70__35_,chained_data_delayed_70__34_,chained_data_delayed_70__33_,
  chained_data_delayed_70__32_,chained_data_delayed_70__31_,chained_data_delayed_70__30_,
  chained_data_delayed_70__29_,chained_data_delayed_70__28_,chained_data_delayed_70__27_,
  chained_data_delayed_70__26_,chained_data_delayed_70__25_,
  chained_data_delayed_70__24_,chained_data_delayed_70__23_,chained_data_delayed_70__22_,
  chained_data_delayed_70__21_,chained_data_delayed_70__20_,chained_data_delayed_70__19_,
  chained_data_delayed_70__18_,chained_data_delayed_70__17_,chained_data_delayed_70__16_,
  chained_data_delayed_70__15_,chained_data_delayed_70__14_,
  chained_data_delayed_70__13_,chained_data_delayed_70__12_,chained_data_delayed_70__11_,
  chained_data_delayed_70__10_,chained_data_delayed_70__9_,chained_data_delayed_70__8_,
  chained_data_delayed_70__7_,chained_data_delayed_70__6_,chained_data_delayed_70__5_,
  chained_data_delayed_70__4_,chained_data_delayed_70__3_,chained_data_delayed_70__2_,
  chained_data_delayed_70__1_,chained_data_delayed_70__0_,
  chained_data_delayed_69__127_,chained_data_delayed_69__126_,chained_data_delayed_69__125_,
  chained_data_delayed_69__124_,chained_data_delayed_69__123_,chained_data_delayed_69__122_,
  chained_data_delayed_69__121_,chained_data_delayed_69__120_,
  chained_data_delayed_69__119_,chained_data_delayed_69__118_,chained_data_delayed_69__117_,
  chained_data_delayed_69__116_,chained_data_delayed_69__115_,chained_data_delayed_69__114_,
  chained_data_delayed_69__113_,chained_data_delayed_69__112_,
  chained_data_delayed_69__111_,chained_data_delayed_69__110_,chained_data_delayed_69__109_,
  chained_data_delayed_69__108_,chained_data_delayed_69__107_,chained_data_delayed_69__106_,
  chained_data_delayed_69__105_,chained_data_delayed_69__104_,
  chained_data_delayed_69__103_,chained_data_delayed_69__102_,chained_data_delayed_69__101_,
  chained_data_delayed_69__100_,chained_data_delayed_69__99_,chained_data_delayed_69__98_,
  chained_data_delayed_69__97_,chained_data_delayed_69__96_,chained_data_delayed_69__95_,
  chained_data_delayed_69__94_,chained_data_delayed_69__93_,
  chained_data_delayed_69__92_,chained_data_delayed_69__91_,chained_data_delayed_69__90_,
  chained_data_delayed_69__89_,chained_data_delayed_69__88_,chained_data_delayed_69__87_,
  chained_data_delayed_69__86_,chained_data_delayed_69__85_,chained_data_delayed_69__84_,
  chained_data_delayed_69__83_,chained_data_delayed_69__82_,
  chained_data_delayed_69__81_,chained_data_delayed_69__80_,chained_data_delayed_69__79_,
  chained_data_delayed_69__78_,chained_data_delayed_69__77_,chained_data_delayed_69__76_,
  chained_data_delayed_69__75_,chained_data_delayed_69__74_,chained_data_delayed_69__73_,
  chained_data_delayed_69__72_,chained_data_delayed_69__71_,
  chained_data_delayed_69__70_,chained_data_delayed_69__69_,chained_data_delayed_69__68_,
  chained_data_delayed_69__67_,chained_data_delayed_69__66_,chained_data_delayed_69__65_,
  chained_data_delayed_69__64_,chained_data_delayed_69__63_,chained_data_delayed_69__62_,
  chained_data_delayed_69__61_,chained_data_delayed_69__60_,
  chained_data_delayed_69__59_,chained_data_delayed_69__58_,chained_data_delayed_69__57_,
  chained_data_delayed_69__56_,chained_data_delayed_69__55_,chained_data_delayed_69__54_,
  chained_data_delayed_69__53_,chained_data_delayed_69__52_,chained_data_delayed_69__51_,
  chained_data_delayed_69__50_,chained_data_delayed_69__49_,chained_data_delayed_69__48_,
  chained_data_delayed_69__47_,chained_data_delayed_69__46_,
  chained_data_delayed_69__45_,chained_data_delayed_69__44_,chained_data_delayed_69__43_,
  chained_data_delayed_69__42_,chained_data_delayed_69__41_,chained_data_delayed_69__40_,
  chained_data_delayed_69__39_,chained_data_delayed_69__38_,chained_data_delayed_69__37_,
  chained_data_delayed_69__36_,chained_data_delayed_69__35_,
  chained_data_delayed_69__34_,chained_data_delayed_69__33_,chained_data_delayed_69__32_,
  chained_data_delayed_69__31_,chained_data_delayed_69__30_,chained_data_delayed_69__29_,
  chained_data_delayed_69__28_,chained_data_delayed_69__27_,chained_data_delayed_69__26_,
  chained_data_delayed_69__25_,chained_data_delayed_69__24_,
  chained_data_delayed_69__23_,chained_data_delayed_69__22_,chained_data_delayed_69__21_,
  chained_data_delayed_69__20_,chained_data_delayed_69__19_,chained_data_delayed_69__18_,
  chained_data_delayed_69__17_,chained_data_delayed_69__16_,chained_data_delayed_69__15_,
  chained_data_delayed_69__14_,chained_data_delayed_69__13_,
  chained_data_delayed_69__12_,chained_data_delayed_69__11_,chained_data_delayed_69__10_,
  chained_data_delayed_69__9_,chained_data_delayed_69__8_,chained_data_delayed_69__7_,
  chained_data_delayed_69__6_,chained_data_delayed_69__5_,chained_data_delayed_69__4_,
  chained_data_delayed_69__3_,chained_data_delayed_69__2_,chained_data_delayed_69__1_,
  chained_data_delayed_69__0_,chained_data_delayed_76__127_,
  chained_data_delayed_76__126_,chained_data_delayed_76__125_,chained_data_delayed_76__124_,
  chained_data_delayed_76__123_,chained_data_delayed_76__122_,chained_data_delayed_76__121_,
  chained_data_delayed_76__120_,chained_data_delayed_76__119_,
  chained_data_delayed_76__118_,chained_data_delayed_76__117_,chained_data_delayed_76__116_,
  chained_data_delayed_76__115_,chained_data_delayed_76__114_,chained_data_delayed_76__113_,
  chained_data_delayed_76__112_,chained_data_delayed_76__111_,
  chained_data_delayed_76__110_,chained_data_delayed_76__109_,chained_data_delayed_76__108_,
  chained_data_delayed_76__107_,chained_data_delayed_76__106_,chained_data_delayed_76__105_,
  chained_data_delayed_76__104_,chained_data_delayed_76__103_,
  chained_data_delayed_76__102_,chained_data_delayed_76__101_,chained_data_delayed_76__100_,
  chained_data_delayed_76__99_,chained_data_delayed_76__98_,chained_data_delayed_76__97_,
  chained_data_delayed_76__96_,chained_data_delayed_76__95_,chained_data_delayed_76__94_,
  chained_data_delayed_76__93_,chained_data_delayed_76__92_,
  chained_data_delayed_76__91_,chained_data_delayed_76__90_,chained_data_delayed_76__89_,
  chained_data_delayed_76__88_,chained_data_delayed_76__87_,chained_data_delayed_76__86_,
  chained_data_delayed_76__85_,chained_data_delayed_76__84_,chained_data_delayed_76__83_,
  chained_data_delayed_76__82_,chained_data_delayed_76__81_,
  chained_data_delayed_76__80_,chained_data_delayed_76__79_,chained_data_delayed_76__78_,
  chained_data_delayed_76__77_,chained_data_delayed_76__76_,chained_data_delayed_76__75_,
  chained_data_delayed_76__74_,chained_data_delayed_76__73_,chained_data_delayed_76__72_,
  chained_data_delayed_76__71_,chained_data_delayed_76__70_,
  chained_data_delayed_76__69_,chained_data_delayed_76__68_,chained_data_delayed_76__67_,
  chained_data_delayed_76__66_,chained_data_delayed_76__65_,chained_data_delayed_76__64_,
  chained_data_delayed_76__63_,chained_data_delayed_76__62_,chained_data_delayed_76__61_,
  chained_data_delayed_76__60_,chained_data_delayed_76__59_,chained_data_delayed_76__58_,
  chained_data_delayed_76__57_,chained_data_delayed_76__56_,
  chained_data_delayed_76__55_,chained_data_delayed_76__54_,chained_data_delayed_76__53_,
  chained_data_delayed_76__52_,chained_data_delayed_76__51_,chained_data_delayed_76__50_,
  chained_data_delayed_76__49_,chained_data_delayed_76__48_,chained_data_delayed_76__47_,
  chained_data_delayed_76__46_,chained_data_delayed_76__45_,
  chained_data_delayed_76__44_,chained_data_delayed_76__43_,chained_data_delayed_76__42_,
  chained_data_delayed_76__41_,chained_data_delayed_76__40_,chained_data_delayed_76__39_,
  chained_data_delayed_76__38_,chained_data_delayed_76__37_,chained_data_delayed_76__36_,
  chained_data_delayed_76__35_,chained_data_delayed_76__34_,
  chained_data_delayed_76__33_,chained_data_delayed_76__32_,chained_data_delayed_76__31_,
  chained_data_delayed_76__30_,chained_data_delayed_76__29_,chained_data_delayed_76__28_,
  chained_data_delayed_76__27_,chained_data_delayed_76__26_,chained_data_delayed_76__25_,
  chained_data_delayed_76__24_,chained_data_delayed_76__23_,
  chained_data_delayed_76__22_,chained_data_delayed_76__21_,chained_data_delayed_76__20_,
  chained_data_delayed_76__19_,chained_data_delayed_76__18_,chained_data_delayed_76__17_,
  chained_data_delayed_76__16_,chained_data_delayed_76__15_,chained_data_delayed_76__14_,
  chained_data_delayed_76__13_,chained_data_delayed_76__12_,
  chained_data_delayed_76__11_,chained_data_delayed_76__10_,chained_data_delayed_76__9_,
  chained_data_delayed_76__8_,chained_data_delayed_76__7_,chained_data_delayed_76__6_,
  chained_data_delayed_76__5_,chained_data_delayed_76__4_,chained_data_delayed_76__3_,
  chained_data_delayed_76__2_,chained_data_delayed_76__1_,chained_data_delayed_76__0_,
  chained_data_delayed_75__127_,chained_data_delayed_75__126_,
  chained_data_delayed_75__125_,chained_data_delayed_75__124_,chained_data_delayed_75__123_,
  chained_data_delayed_75__122_,chained_data_delayed_75__121_,chained_data_delayed_75__120_,
  chained_data_delayed_75__119_,chained_data_delayed_75__118_,
  chained_data_delayed_75__117_,chained_data_delayed_75__116_,chained_data_delayed_75__115_,
  chained_data_delayed_75__114_,chained_data_delayed_75__113_,chained_data_delayed_75__112_,
  chained_data_delayed_75__111_,chained_data_delayed_75__110_,
  chained_data_delayed_75__109_,chained_data_delayed_75__108_,chained_data_delayed_75__107_,
  chained_data_delayed_75__106_,chained_data_delayed_75__105_,chained_data_delayed_75__104_,
  chained_data_delayed_75__103_,chained_data_delayed_75__102_,
  chained_data_delayed_75__101_,chained_data_delayed_75__100_,chained_data_delayed_75__99_,
  chained_data_delayed_75__98_,chained_data_delayed_75__97_,chained_data_delayed_75__96_,
  chained_data_delayed_75__95_,chained_data_delayed_75__94_,chained_data_delayed_75__93_,
  chained_data_delayed_75__92_,chained_data_delayed_75__91_,
  chained_data_delayed_75__90_,chained_data_delayed_75__89_,chained_data_delayed_75__88_,
  chained_data_delayed_75__87_,chained_data_delayed_75__86_,chained_data_delayed_75__85_,
  chained_data_delayed_75__84_,chained_data_delayed_75__83_,chained_data_delayed_75__82_,
  chained_data_delayed_75__81_,chained_data_delayed_75__80_,
  chained_data_delayed_75__79_,chained_data_delayed_75__78_,chained_data_delayed_75__77_,
  chained_data_delayed_75__76_,chained_data_delayed_75__75_,chained_data_delayed_75__74_,
  chained_data_delayed_75__73_,chained_data_delayed_75__72_,chained_data_delayed_75__71_,
  chained_data_delayed_75__70_,chained_data_delayed_75__69_,chained_data_delayed_75__68_,
  chained_data_delayed_75__67_,chained_data_delayed_75__66_,
  chained_data_delayed_75__65_,chained_data_delayed_75__64_,chained_data_delayed_75__63_,
  chained_data_delayed_75__62_,chained_data_delayed_75__61_,chained_data_delayed_75__60_,
  chained_data_delayed_75__59_,chained_data_delayed_75__58_,chained_data_delayed_75__57_,
  chained_data_delayed_75__56_,chained_data_delayed_75__55_,
  chained_data_delayed_75__54_,chained_data_delayed_75__53_,chained_data_delayed_75__52_,
  chained_data_delayed_75__51_,chained_data_delayed_75__50_,chained_data_delayed_75__49_,
  chained_data_delayed_75__48_,chained_data_delayed_75__47_,chained_data_delayed_75__46_,
  chained_data_delayed_75__45_,chained_data_delayed_75__44_,
  chained_data_delayed_75__43_,chained_data_delayed_75__42_,chained_data_delayed_75__41_,
  chained_data_delayed_75__40_,chained_data_delayed_75__39_,chained_data_delayed_75__38_,
  chained_data_delayed_75__37_,chained_data_delayed_75__36_,chained_data_delayed_75__35_,
  chained_data_delayed_75__34_,chained_data_delayed_75__33_,
  chained_data_delayed_75__32_,chained_data_delayed_75__31_,chained_data_delayed_75__30_,
  chained_data_delayed_75__29_,chained_data_delayed_75__28_,chained_data_delayed_75__27_,
  chained_data_delayed_75__26_,chained_data_delayed_75__25_,chained_data_delayed_75__24_,
  chained_data_delayed_75__23_,chained_data_delayed_75__22_,
  chained_data_delayed_75__21_,chained_data_delayed_75__20_,chained_data_delayed_75__19_,
  chained_data_delayed_75__18_,chained_data_delayed_75__17_,chained_data_delayed_75__16_,
  chained_data_delayed_75__15_,chained_data_delayed_75__14_,chained_data_delayed_75__13_,
  chained_data_delayed_75__12_,chained_data_delayed_75__11_,
  chained_data_delayed_75__10_,chained_data_delayed_75__9_,chained_data_delayed_75__8_,
  chained_data_delayed_75__7_,chained_data_delayed_75__6_,chained_data_delayed_75__5_,
  chained_data_delayed_75__4_,chained_data_delayed_75__3_,chained_data_delayed_75__2_,
  chained_data_delayed_75__1_,chained_data_delayed_75__0_,chained_data_delayed_74__127_,
  chained_data_delayed_74__126_,chained_data_delayed_74__125_,
  chained_data_delayed_74__124_,chained_data_delayed_74__123_,chained_data_delayed_74__122_,
  chained_data_delayed_74__121_,chained_data_delayed_74__120_,chained_data_delayed_74__119_,
  chained_data_delayed_74__118_,chained_data_delayed_74__117_,
  chained_data_delayed_74__116_,chained_data_delayed_74__115_,chained_data_delayed_74__114_,
  chained_data_delayed_74__113_,chained_data_delayed_74__112_,chained_data_delayed_74__111_,
  chained_data_delayed_74__110_,chained_data_delayed_74__109_,
  chained_data_delayed_74__108_,chained_data_delayed_74__107_,chained_data_delayed_74__106_,
  chained_data_delayed_74__105_,chained_data_delayed_74__104_,chained_data_delayed_74__103_,
  chained_data_delayed_74__102_,chained_data_delayed_74__101_,
  chained_data_delayed_74__100_,chained_data_delayed_74__99_,chained_data_delayed_74__98_,
  chained_data_delayed_74__97_,chained_data_delayed_74__96_,chained_data_delayed_74__95_,
  chained_data_delayed_74__94_,chained_data_delayed_74__93_,chained_data_delayed_74__92_,
  chained_data_delayed_74__91_,chained_data_delayed_74__90_,
  chained_data_delayed_74__89_,chained_data_delayed_74__88_,chained_data_delayed_74__87_,
  chained_data_delayed_74__86_,chained_data_delayed_74__85_,chained_data_delayed_74__84_,
  chained_data_delayed_74__83_,chained_data_delayed_74__82_,chained_data_delayed_74__81_,
  chained_data_delayed_74__80_,chained_data_delayed_74__79_,chained_data_delayed_74__78_,
  chained_data_delayed_74__77_,chained_data_delayed_74__76_,
  chained_data_delayed_74__75_,chained_data_delayed_74__74_,chained_data_delayed_74__73_,
  chained_data_delayed_74__72_,chained_data_delayed_74__71_,chained_data_delayed_74__70_,
  chained_data_delayed_74__69_,chained_data_delayed_74__68_,chained_data_delayed_74__67_,
  chained_data_delayed_74__66_,chained_data_delayed_74__65_,
  chained_data_delayed_74__64_,chained_data_delayed_74__63_,chained_data_delayed_74__62_,
  chained_data_delayed_74__61_,chained_data_delayed_74__60_,chained_data_delayed_74__59_,
  chained_data_delayed_74__58_,chained_data_delayed_74__57_,chained_data_delayed_74__56_,
  chained_data_delayed_74__55_,chained_data_delayed_74__54_,
  chained_data_delayed_74__53_,chained_data_delayed_74__52_,chained_data_delayed_74__51_,
  chained_data_delayed_74__50_,chained_data_delayed_74__49_,chained_data_delayed_74__48_,
  chained_data_delayed_74__47_,chained_data_delayed_74__46_,chained_data_delayed_74__45_,
  chained_data_delayed_74__44_,chained_data_delayed_74__43_,
  chained_data_delayed_74__42_,chained_data_delayed_74__41_,chained_data_delayed_74__40_,
  chained_data_delayed_74__39_,chained_data_delayed_74__38_,chained_data_delayed_74__37_,
  chained_data_delayed_74__36_,chained_data_delayed_74__35_,chained_data_delayed_74__34_,
  chained_data_delayed_74__33_,chained_data_delayed_74__32_,
  chained_data_delayed_74__31_,chained_data_delayed_74__30_,chained_data_delayed_74__29_,
  chained_data_delayed_74__28_,chained_data_delayed_74__27_,chained_data_delayed_74__26_,
  chained_data_delayed_74__25_,chained_data_delayed_74__24_,chained_data_delayed_74__23_,
  chained_data_delayed_74__22_,chained_data_delayed_74__21_,
  chained_data_delayed_74__20_,chained_data_delayed_74__19_,chained_data_delayed_74__18_,
  chained_data_delayed_74__17_,chained_data_delayed_74__16_,chained_data_delayed_74__15_,
  chained_data_delayed_74__14_,chained_data_delayed_74__13_,chained_data_delayed_74__12_,
  chained_data_delayed_74__11_,chained_data_delayed_74__10_,chained_data_delayed_74__9_,
  chained_data_delayed_74__8_,chained_data_delayed_74__7_,
  chained_data_delayed_74__6_,chained_data_delayed_74__5_,chained_data_delayed_74__4_,
  chained_data_delayed_74__3_,chained_data_delayed_74__2_,chained_data_delayed_74__1_,
  chained_data_delayed_74__0_,chained_data_delayed_73__127_,chained_data_delayed_73__126_,
  chained_data_delayed_73__125_,chained_data_delayed_73__124_,
  chained_data_delayed_73__123_,chained_data_delayed_73__122_,chained_data_delayed_73__121_,
  chained_data_delayed_73__120_,chained_data_delayed_73__119_,chained_data_delayed_73__118_,
  chained_data_delayed_73__117_,chained_data_delayed_73__116_,
  chained_data_delayed_73__115_,chained_data_delayed_73__114_,chained_data_delayed_73__113_,
  chained_data_delayed_73__112_,chained_data_delayed_73__111_,chained_data_delayed_73__110_,
  chained_data_delayed_73__109_,chained_data_delayed_73__108_,
  chained_data_delayed_73__107_,chained_data_delayed_73__106_,chained_data_delayed_73__105_,
  chained_data_delayed_73__104_,chained_data_delayed_73__103_,chained_data_delayed_73__102_,
  chained_data_delayed_73__101_,chained_data_delayed_73__100_,
  chained_data_delayed_73__99_,chained_data_delayed_73__98_,chained_data_delayed_73__97_,
  chained_data_delayed_73__96_,chained_data_delayed_73__95_,chained_data_delayed_73__94_,
  chained_data_delayed_73__93_,chained_data_delayed_73__92_,chained_data_delayed_73__91_,
  chained_data_delayed_73__90_,chained_data_delayed_73__89_,chained_data_delayed_73__88_,
  chained_data_delayed_73__87_,chained_data_delayed_73__86_,
  chained_data_delayed_73__85_,chained_data_delayed_73__84_,chained_data_delayed_73__83_,
  chained_data_delayed_73__82_,chained_data_delayed_73__81_,chained_data_delayed_73__80_,
  chained_data_delayed_73__79_,chained_data_delayed_73__78_,chained_data_delayed_73__77_,
  chained_data_delayed_73__76_,chained_data_delayed_73__75_,
  chained_data_delayed_73__74_,chained_data_delayed_73__73_,chained_data_delayed_73__72_,
  chained_data_delayed_73__71_,chained_data_delayed_73__70_,chained_data_delayed_73__69_,
  chained_data_delayed_73__68_,chained_data_delayed_73__67_,chained_data_delayed_73__66_,
  chained_data_delayed_73__65_,chained_data_delayed_73__64_,
  chained_data_delayed_73__63_,chained_data_delayed_73__62_,chained_data_delayed_73__61_,
  chained_data_delayed_73__60_,chained_data_delayed_73__59_,chained_data_delayed_73__58_,
  chained_data_delayed_73__57_,chained_data_delayed_73__56_,chained_data_delayed_73__55_,
  chained_data_delayed_73__54_,chained_data_delayed_73__53_,
  chained_data_delayed_73__52_,chained_data_delayed_73__51_,chained_data_delayed_73__50_,
  chained_data_delayed_73__49_,chained_data_delayed_73__48_,chained_data_delayed_73__47_,
  chained_data_delayed_73__46_,chained_data_delayed_73__45_,chained_data_delayed_73__44_,
  chained_data_delayed_73__43_,chained_data_delayed_73__42_,
  chained_data_delayed_73__41_,chained_data_delayed_73__40_,chained_data_delayed_73__39_,
  chained_data_delayed_73__38_,chained_data_delayed_73__37_,chained_data_delayed_73__36_,
  chained_data_delayed_73__35_,chained_data_delayed_73__34_,chained_data_delayed_73__33_,
  chained_data_delayed_73__32_,chained_data_delayed_73__31_,
  chained_data_delayed_73__30_,chained_data_delayed_73__29_,chained_data_delayed_73__28_,
  chained_data_delayed_73__27_,chained_data_delayed_73__26_,chained_data_delayed_73__25_,
  chained_data_delayed_73__24_,chained_data_delayed_73__23_,chained_data_delayed_73__22_,
  chained_data_delayed_73__21_,chained_data_delayed_73__20_,
  chained_data_delayed_73__19_,chained_data_delayed_73__18_,chained_data_delayed_73__17_,
  chained_data_delayed_73__16_,chained_data_delayed_73__15_,chained_data_delayed_73__14_,
  chained_data_delayed_73__13_,chained_data_delayed_73__12_,chained_data_delayed_73__11_,
  chained_data_delayed_73__10_,chained_data_delayed_73__9_,chained_data_delayed_73__8_,
  chained_data_delayed_73__7_,chained_data_delayed_73__6_,
  chained_data_delayed_73__5_,chained_data_delayed_73__4_,chained_data_delayed_73__3_,
  chained_data_delayed_73__2_,chained_data_delayed_73__1_,chained_data_delayed_73__0_,
  chained_data_delayed_80__127_,chained_data_delayed_80__126_,chained_data_delayed_80__125_,
  chained_data_delayed_80__124_,chained_data_delayed_80__123_,
  chained_data_delayed_80__122_,chained_data_delayed_80__121_,chained_data_delayed_80__120_,
  chained_data_delayed_80__119_,chained_data_delayed_80__118_,chained_data_delayed_80__117_,
  chained_data_delayed_80__116_,chained_data_delayed_80__115_,
  chained_data_delayed_80__114_,chained_data_delayed_80__113_,chained_data_delayed_80__112_,
  chained_data_delayed_80__111_,chained_data_delayed_80__110_,chained_data_delayed_80__109_,
  chained_data_delayed_80__108_,chained_data_delayed_80__107_,
  chained_data_delayed_80__106_,chained_data_delayed_80__105_,chained_data_delayed_80__104_,
  chained_data_delayed_80__103_,chained_data_delayed_80__102_,chained_data_delayed_80__101_,
  chained_data_delayed_80__100_,chained_data_delayed_80__99_,chained_data_delayed_80__98_,
  chained_data_delayed_80__97_,chained_data_delayed_80__96_,
  chained_data_delayed_80__95_,chained_data_delayed_80__94_,chained_data_delayed_80__93_,
  chained_data_delayed_80__92_,chained_data_delayed_80__91_,chained_data_delayed_80__90_,
  chained_data_delayed_80__89_,chained_data_delayed_80__88_,chained_data_delayed_80__87_,
  chained_data_delayed_80__86_,chained_data_delayed_80__85_,
  chained_data_delayed_80__84_,chained_data_delayed_80__83_,chained_data_delayed_80__82_,
  chained_data_delayed_80__81_,chained_data_delayed_80__80_,chained_data_delayed_80__79_,
  chained_data_delayed_80__78_,chained_data_delayed_80__77_,chained_data_delayed_80__76_,
  chained_data_delayed_80__75_,chained_data_delayed_80__74_,
  chained_data_delayed_80__73_,chained_data_delayed_80__72_,chained_data_delayed_80__71_,
  chained_data_delayed_80__70_,chained_data_delayed_80__69_,chained_data_delayed_80__68_,
  chained_data_delayed_80__67_,chained_data_delayed_80__66_,chained_data_delayed_80__65_,
  chained_data_delayed_80__64_,chained_data_delayed_80__63_,
  chained_data_delayed_80__62_,chained_data_delayed_80__61_,chained_data_delayed_80__60_,
  chained_data_delayed_80__59_,chained_data_delayed_80__58_,chained_data_delayed_80__57_,
  chained_data_delayed_80__56_,chained_data_delayed_80__55_,chained_data_delayed_80__54_,
  chained_data_delayed_80__53_,chained_data_delayed_80__52_,
  chained_data_delayed_80__51_,chained_data_delayed_80__50_,chained_data_delayed_80__49_,
  chained_data_delayed_80__48_,chained_data_delayed_80__47_,chained_data_delayed_80__46_,
  chained_data_delayed_80__45_,chained_data_delayed_80__44_,chained_data_delayed_80__43_,
  chained_data_delayed_80__42_,chained_data_delayed_80__41_,
  chained_data_delayed_80__40_,chained_data_delayed_80__39_,chained_data_delayed_80__38_,
  chained_data_delayed_80__37_,chained_data_delayed_80__36_,chained_data_delayed_80__35_,
  chained_data_delayed_80__34_,chained_data_delayed_80__33_,chained_data_delayed_80__32_,
  chained_data_delayed_80__31_,chained_data_delayed_80__30_,
  chained_data_delayed_80__29_,chained_data_delayed_80__28_,chained_data_delayed_80__27_,
  chained_data_delayed_80__26_,chained_data_delayed_80__25_,chained_data_delayed_80__24_,
  chained_data_delayed_80__23_,chained_data_delayed_80__22_,chained_data_delayed_80__21_,
  chained_data_delayed_80__20_,chained_data_delayed_80__19_,chained_data_delayed_80__18_,
  chained_data_delayed_80__17_,chained_data_delayed_80__16_,
  chained_data_delayed_80__15_,chained_data_delayed_80__14_,chained_data_delayed_80__13_,
  chained_data_delayed_80__12_,chained_data_delayed_80__11_,chained_data_delayed_80__10_,
  chained_data_delayed_80__9_,chained_data_delayed_80__8_,chained_data_delayed_80__7_,
  chained_data_delayed_80__6_,chained_data_delayed_80__5_,chained_data_delayed_80__4_,
  chained_data_delayed_80__3_,chained_data_delayed_80__2_,
  chained_data_delayed_80__1_,chained_data_delayed_80__0_,chained_data_delayed_79__127_,
  chained_data_delayed_79__126_,chained_data_delayed_79__125_,chained_data_delayed_79__124_,
  chained_data_delayed_79__123_,chained_data_delayed_79__122_,
  chained_data_delayed_79__121_,chained_data_delayed_79__120_,chained_data_delayed_79__119_,
  chained_data_delayed_79__118_,chained_data_delayed_79__117_,chained_data_delayed_79__116_,
  chained_data_delayed_79__115_,chained_data_delayed_79__114_,
  chained_data_delayed_79__113_,chained_data_delayed_79__112_,chained_data_delayed_79__111_,
  chained_data_delayed_79__110_,chained_data_delayed_79__109_,chained_data_delayed_79__108_,
  chained_data_delayed_79__107_,chained_data_delayed_79__106_,
  chained_data_delayed_79__105_,chained_data_delayed_79__104_,chained_data_delayed_79__103_,
  chained_data_delayed_79__102_,chained_data_delayed_79__101_,chained_data_delayed_79__100_,
  chained_data_delayed_79__99_,chained_data_delayed_79__98_,chained_data_delayed_79__97_,
  chained_data_delayed_79__96_,chained_data_delayed_79__95_,
  chained_data_delayed_79__94_,chained_data_delayed_79__93_,chained_data_delayed_79__92_,
  chained_data_delayed_79__91_,chained_data_delayed_79__90_,chained_data_delayed_79__89_,
  chained_data_delayed_79__88_,chained_data_delayed_79__87_,chained_data_delayed_79__86_,
  chained_data_delayed_79__85_,chained_data_delayed_79__84_,
  chained_data_delayed_79__83_,chained_data_delayed_79__82_,chained_data_delayed_79__81_,
  chained_data_delayed_79__80_,chained_data_delayed_79__79_,chained_data_delayed_79__78_,
  chained_data_delayed_79__77_,chained_data_delayed_79__76_,chained_data_delayed_79__75_,
  chained_data_delayed_79__74_,chained_data_delayed_79__73_,
  chained_data_delayed_79__72_,chained_data_delayed_79__71_,chained_data_delayed_79__70_,
  chained_data_delayed_79__69_,chained_data_delayed_79__68_,chained_data_delayed_79__67_,
  chained_data_delayed_79__66_,chained_data_delayed_79__65_,chained_data_delayed_79__64_,
  chained_data_delayed_79__63_,chained_data_delayed_79__62_,
  chained_data_delayed_79__61_,chained_data_delayed_79__60_,chained_data_delayed_79__59_,
  chained_data_delayed_79__58_,chained_data_delayed_79__57_,chained_data_delayed_79__56_,
  chained_data_delayed_79__55_,chained_data_delayed_79__54_,chained_data_delayed_79__53_,
  chained_data_delayed_79__52_,chained_data_delayed_79__51_,
  chained_data_delayed_79__50_,chained_data_delayed_79__49_,chained_data_delayed_79__48_,
  chained_data_delayed_79__47_,chained_data_delayed_79__46_,chained_data_delayed_79__45_,
  chained_data_delayed_79__44_,chained_data_delayed_79__43_,chained_data_delayed_79__42_,
  chained_data_delayed_79__41_,chained_data_delayed_79__40_,
  chained_data_delayed_79__39_,chained_data_delayed_79__38_,chained_data_delayed_79__37_,
  chained_data_delayed_79__36_,chained_data_delayed_79__35_,chained_data_delayed_79__34_,
  chained_data_delayed_79__33_,chained_data_delayed_79__32_,chained_data_delayed_79__31_,
  chained_data_delayed_79__30_,chained_data_delayed_79__29_,chained_data_delayed_79__28_,
  chained_data_delayed_79__27_,chained_data_delayed_79__26_,
  chained_data_delayed_79__25_,chained_data_delayed_79__24_,chained_data_delayed_79__23_,
  chained_data_delayed_79__22_,chained_data_delayed_79__21_,chained_data_delayed_79__20_,
  chained_data_delayed_79__19_,chained_data_delayed_79__18_,chained_data_delayed_79__17_,
  chained_data_delayed_79__16_,chained_data_delayed_79__15_,
  chained_data_delayed_79__14_,chained_data_delayed_79__13_,chained_data_delayed_79__12_,
  chained_data_delayed_79__11_,chained_data_delayed_79__10_,chained_data_delayed_79__9_,
  chained_data_delayed_79__8_,chained_data_delayed_79__7_,chained_data_delayed_79__6_,
  chained_data_delayed_79__5_,chained_data_delayed_79__4_,chained_data_delayed_79__3_,
  chained_data_delayed_79__2_,chained_data_delayed_79__1_,
  chained_data_delayed_79__0_,chained_data_delayed_78__127_,chained_data_delayed_78__126_,
  chained_data_delayed_78__125_,chained_data_delayed_78__124_,chained_data_delayed_78__123_,
  chained_data_delayed_78__122_,chained_data_delayed_78__121_,
  chained_data_delayed_78__120_,chained_data_delayed_78__119_,chained_data_delayed_78__118_,
  chained_data_delayed_78__117_,chained_data_delayed_78__116_,chained_data_delayed_78__115_,
  chained_data_delayed_78__114_,chained_data_delayed_78__113_,
  chained_data_delayed_78__112_,chained_data_delayed_78__111_,chained_data_delayed_78__110_,
  chained_data_delayed_78__109_,chained_data_delayed_78__108_,chained_data_delayed_78__107_,
  chained_data_delayed_78__106_,chained_data_delayed_78__105_,
  chained_data_delayed_78__104_,chained_data_delayed_78__103_,chained_data_delayed_78__102_,
  chained_data_delayed_78__101_,chained_data_delayed_78__100_,chained_data_delayed_78__99_,
  chained_data_delayed_78__98_,chained_data_delayed_78__97_,chained_data_delayed_78__96_,
  chained_data_delayed_78__95_,chained_data_delayed_78__94_,
  chained_data_delayed_78__93_,chained_data_delayed_78__92_,chained_data_delayed_78__91_,
  chained_data_delayed_78__90_,chained_data_delayed_78__89_,chained_data_delayed_78__88_,
  chained_data_delayed_78__87_,chained_data_delayed_78__86_,chained_data_delayed_78__85_,
  chained_data_delayed_78__84_,chained_data_delayed_78__83_,
  chained_data_delayed_78__82_,chained_data_delayed_78__81_,chained_data_delayed_78__80_,
  chained_data_delayed_78__79_,chained_data_delayed_78__78_,chained_data_delayed_78__77_,
  chained_data_delayed_78__76_,chained_data_delayed_78__75_,chained_data_delayed_78__74_,
  chained_data_delayed_78__73_,chained_data_delayed_78__72_,
  chained_data_delayed_78__71_,chained_data_delayed_78__70_,chained_data_delayed_78__69_,
  chained_data_delayed_78__68_,chained_data_delayed_78__67_,chained_data_delayed_78__66_,
  chained_data_delayed_78__65_,chained_data_delayed_78__64_,chained_data_delayed_78__63_,
  chained_data_delayed_78__62_,chained_data_delayed_78__61_,
  chained_data_delayed_78__60_,chained_data_delayed_78__59_,chained_data_delayed_78__58_,
  chained_data_delayed_78__57_,chained_data_delayed_78__56_,chained_data_delayed_78__55_,
  chained_data_delayed_78__54_,chained_data_delayed_78__53_,chained_data_delayed_78__52_,
  chained_data_delayed_78__51_,chained_data_delayed_78__50_,
  chained_data_delayed_78__49_,chained_data_delayed_78__48_,chained_data_delayed_78__47_,
  chained_data_delayed_78__46_,chained_data_delayed_78__45_,chained_data_delayed_78__44_,
  chained_data_delayed_78__43_,chained_data_delayed_78__42_,chained_data_delayed_78__41_,
  chained_data_delayed_78__40_,chained_data_delayed_78__39_,chained_data_delayed_78__38_,
  chained_data_delayed_78__37_,chained_data_delayed_78__36_,
  chained_data_delayed_78__35_,chained_data_delayed_78__34_,chained_data_delayed_78__33_,
  chained_data_delayed_78__32_,chained_data_delayed_78__31_,chained_data_delayed_78__30_,
  chained_data_delayed_78__29_,chained_data_delayed_78__28_,chained_data_delayed_78__27_,
  chained_data_delayed_78__26_,chained_data_delayed_78__25_,
  chained_data_delayed_78__24_,chained_data_delayed_78__23_,chained_data_delayed_78__22_,
  chained_data_delayed_78__21_,chained_data_delayed_78__20_,chained_data_delayed_78__19_,
  chained_data_delayed_78__18_,chained_data_delayed_78__17_,chained_data_delayed_78__16_,
  chained_data_delayed_78__15_,chained_data_delayed_78__14_,
  chained_data_delayed_78__13_,chained_data_delayed_78__12_,chained_data_delayed_78__11_,
  chained_data_delayed_78__10_,chained_data_delayed_78__9_,chained_data_delayed_78__8_,
  chained_data_delayed_78__7_,chained_data_delayed_78__6_,chained_data_delayed_78__5_,
  chained_data_delayed_78__4_,chained_data_delayed_78__3_,chained_data_delayed_78__2_,
  chained_data_delayed_78__1_,chained_data_delayed_78__0_,
  chained_data_delayed_77__127_,chained_data_delayed_77__126_,chained_data_delayed_77__125_,
  chained_data_delayed_77__124_,chained_data_delayed_77__123_,chained_data_delayed_77__122_,
  chained_data_delayed_77__121_,chained_data_delayed_77__120_,
  chained_data_delayed_77__119_,chained_data_delayed_77__118_,chained_data_delayed_77__117_,
  chained_data_delayed_77__116_,chained_data_delayed_77__115_,chained_data_delayed_77__114_,
  chained_data_delayed_77__113_,chained_data_delayed_77__112_,
  chained_data_delayed_77__111_,chained_data_delayed_77__110_,chained_data_delayed_77__109_,
  chained_data_delayed_77__108_,chained_data_delayed_77__107_,chained_data_delayed_77__106_,
  chained_data_delayed_77__105_,chained_data_delayed_77__104_,
  chained_data_delayed_77__103_,chained_data_delayed_77__102_,chained_data_delayed_77__101_,
  chained_data_delayed_77__100_,chained_data_delayed_77__99_,chained_data_delayed_77__98_,
  chained_data_delayed_77__97_,chained_data_delayed_77__96_,chained_data_delayed_77__95_,
  chained_data_delayed_77__94_,chained_data_delayed_77__93_,
  chained_data_delayed_77__92_,chained_data_delayed_77__91_,chained_data_delayed_77__90_,
  chained_data_delayed_77__89_,chained_data_delayed_77__88_,chained_data_delayed_77__87_,
  chained_data_delayed_77__86_,chained_data_delayed_77__85_,chained_data_delayed_77__84_,
  chained_data_delayed_77__83_,chained_data_delayed_77__82_,
  chained_data_delayed_77__81_,chained_data_delayed_77__80_,chained_data_delayed_77__79_,
  chained_data_delayed_77__78_,chained_data_delayed_77__77_,chained_data_delayed_77__76_,
  chained_data_delayed_77__75_,chained_data_delayed_77__74_,chained_data_delayed_77__73_,
  chained_data_delayed_77__72_,chained_data_delayed_77__71_,
  chained_data_delayed_77__70_,chained_data_delayed_77__69_,chained_data_delayed_77__68_,
  chained_data_delayed_77__67_,chained_data_delayed_77__66_,chained_data_delayed_77__65_,
  chained_data_delayed_77__64_,chained_data_delayed_77__63_,chained_data_delayed_77__62_,
  chained_data_delayed_77__61_,chained_data_delayed_77__60_,
  chained_data_delayed_77__59_,chained_data_delayed_77__58_,chained_data_delayed_77__57_,
  chained_data_delayed_77__56_,chained_data_delayed_77__55_,chained_data_delayed_77__54_,
  chained_data_delayed_77__53_,chained_data_delayed_77__52_,chained_data_delayed_77__51_,
  chained_data_delayed_77__50_,chained_data_delayed_77__49_,chained_data_delayed_77__48_,
  chained_data_delayed_77__47_,chained_data_delayed_77__46_,
  chained_data_delayed_77__45_,chained_data_delayed_77__44_,chained_data_delayed_77__43_,
  chained_data_delayed_77__42_,chained_data_delayed_77__41_,chained_data_delayed_77__40_,
  chained_data_delayed_77__39_,chained_data_delayed_77__38_,chained_data_delayed_77__37_,
  chained_data_delayed_77__36_,chained_data_delayed_77__35_,
  chained_data_delayed_77__34_,chained_data_delayed_77__33_,chained_data_delayed_77__32_,
  chained_data_delayed_77__31_,chained_data_delayed_77__30_,chained_data_delayed_77__29_,
  chained_data_delayed_77__28_,chained_data_delayed_77__27_,chained_data_delayed_77__26_,
  chained_data_delayed_77__25_,chained_data_delayed_77__24_,
  chained_data_delayed_77__23_,chained_data_delayed_77__22_,chained_data_delayed_77__21_,
  chained_data_delayed_77__20_,chained_data_delayed_77__19_,chained_data_delayed_77__18_,
  chained_data_delayed_77__17_,chained_data_delayed_77__16_,chained_data_delayed_77__15_,
  chained_data_delayed_77__14_,chained_data_delayed_77__13_,
  chained_data_delayed_77__12_,chained_data_delayed_77__11_,chained_data_delayed_77__10_,
  chained_data_delayed_77__9_,chained_data_delayed_77__8_,chained_data_delayed_77__7_,
  chained_data_delayed_77__6_,chained_data_delayed_77__5_,chained_data_delayed_77__4_,
  chained_data_delayed_77__3_,chained_data_delayed_77__2_,chained_data_delayed_77__1_,
  chained_data_delayed_77__0_,chained_data_delayed_84__127_,
  chained_data_delayed_84__126_,chained_data_delayed_84__125_,chained_data_delayed_84__124_,
  chained_data_delayed_84__123_,chained_data_delayed_84__122_,chained_data_delayed_84__121_,
  chained_data_delayed_84__120_,chained_data_delayed_84__119_,
  chained_data_delayed_84__118_,chained_data_delayed_84__117_,chained_data_delayed_84__116_,
  chained_data_delayed_84__115_,chained_data_delayed_84__114_,chained_data_delayed_84__113_,
  chained_data_delayed_84__112_,chained_data_delayed_84__111_,
  chained_data_delayed_84__110_,chained_data_delayed_84__109_,chained_data_delayed_84__108_,
  chained_data_delayed_84__107_,chained_data_delayed_84__106_,chained_data_delayed_84__105_,
  chained_data_delayed_84__104_,chained_data_delayed_84__103_,
  chained_data_delayed_84__102_,chained_data_delayed_84__101_,chained_data_delayed_84__100_,
  chained_data_delayed_84__99_,chained_data_delayed_84__98_,chained_data_delayed_84__97_,
  chained_data_delayed_84__96_,chained_data_delayed_84__95_,chained_data_delayed_84__94_,
  chained_data_delayed_84__93_,chained_data_delayed_84__92_,
  chained_data_delayed_84__91_,chained_data_delayed_84__90_,chained_data_delayed_84__89_,
  chained_data_delayed_84__88_,chained_data_delayed_84__87_,chained_data_delayed_84__86_,
  chained_data_delayed_84__85_,chained_data_delayed_84__84_,chained_data_delayed_84__83_,
  chained_data_delayed_84__82_,chained_data_delayed_84__81_,
  chained_data_delayed_84__80_,chained_data_delayed_84__79_,chained_data_delayed_84__78_,
  chained_data_delayed_84__77_,chained_data_delayed_84__76_,chained_data_delayed_84__75_,
  chained_data_delayed_84__74_,chained_data_delayed_84__73_,chained_data_delayed_84__72_,
  chained_data_delayed_84__71_,chained_data_delayed_84__70_,
  chained_data_delayed_84__69_,chained_data_delayed_84__68_,chained_data_delayed_84__67_,
  chained_data_delayed_84__66_,chained_data_delayed_84__65_,chained_data_delayed_84__64_,
  chained_data_delayed_84__63_,chained_data_delayed_84__62_,chained_data_delayed_84__61_,
  chained_data_delayed_84__60_,chained_data_delayed_84__59_,chained_data_delayed_84__58_,
  chained_data_delayed_84__57_,chained_data_delayed_84__56_,
  chained_data_delayed_84__55_,chained_data_delayed_84__54_,chained_data_delayed_84__53_,
  chained_data_delayed_84__52_,chained_data_delayed_84__51_,chained_data_delayed_84__50_,
  chained_data_delayed_84__49_,chained_data_delayed_84__48_,chained_data_delayed_84__47_,
  chained_data_delayed_84__46_,chained_data_delayed_84__45_,
  chained_data_delayed_84__44_,chained_data_delayed_84__43_,chained_data_delayed_84__42_,
  chained_data_delayed_84__41_,chained_data_delayed_84__40_,chained_data_delayed_84__39_,
  chained_data_delayed_84__38_,chained_data_delayed_84__37_,chained_data_delayed_84__36_,
  chained_data_delayed_84__35_,chained_data_delayed_84__34_,
  chained_data_delayed_84__33_,chained_data_delayed_84__32_,chained_data_delayed_84__31_,
  chained_data_delayed_84__30_,chained_data_delayed_84__29_,chained_data_delayed_84__28_,
  chained_data_delayed_84__27_,chained_data_delayed_84__26_,chained_data_delayed_84__25_,
  chained_data_delayed_84__24_,chained_data_delayed_84__23_,
  chained_data_delayed_84__22_,chained_data_delayed_84__21_,chained_data_delayed_84__20_,
  chained_data_delayed_84__19_,chained_data_delayed_84__18_,chained_data_delayed_84__17_,
  chained_data_delayed_84__16_,chained_data_delayed_84__15_,chained_data_delayed_84__14_,
  chained_data_delayed_84__13_,chained_data_delayed_84__12_,
  chained_data_delayed_84__11_,chained_data_delayed_84__10_,chained_data_delayed_84__9_,
  chained_data_delayed_84__8_,chained_data_delayed_84__7_,chained_data_delayed_84__6_,
  chained_data_delayed_84__5_,chained_data_delayed_84__4_,chained_data_delayed_84__3_,
  chained_data_delayed_84__2_,chained_data_delayed_84__1_,chained_data_delayed_84__0_,
  chained_data_delayed_83__127_,chained_data_delayed_83__126_,
  chained_data_delayed_83__125_,chained_data_delayed_83__124_,chained_data_delayed_83__123_,
  chained_data_delayed_83__122_,chained_data_delayed_83__121_,chained_data_delayed_83__120_,
  chained_data_delayed_83__119_,chained_data_delayed_83__118_,
  chained_data_delayed_83__117_,chained_data_delayed_83__116_,chained_data_delayed_83__115_,
  chained_data_delayed_83__114_,chained_data_delayed_83__113_,chained_data_delayed_83__112_,
  chained_data_delayed_83__111_,chained_data_delayed_83__110_,
  chained_data_delayed_83__109_,chained_data_delayed_83__108_,chained_data_delayed_83__107_,
  chained_data_delayed_83__106_,chained_data_delayed_83__105_,chained_data_delayed_83__104_,
  chained_data_delayed_83__103_,chained_data_delayed_83__102_,
  chained_data_delayed_83__101_,chained_data_delayed_83__100_,chained_data_delayed_83__99_,
  chained_data_delayed_83__98_,chained_data_delayed_83__97_,chained_data_delayed_83__96_,
  chained_data_delayed_83__95_,chained_data_delayed_83__94_,chained_data_delayed_83__93_,
  chained_data_delayed_83__92_,chained_data_delayed_83__91_,
  chained_data_delayed_83__90_,chained_data_delayed_83__89_,chained_data_delayed_83__88_,
  chained_data_delayed_83__87_,chained_data_delayed_83__86_,chained_data_delayed_83__85_,
  chained_data_delayed_83__84_,chained_data_delayed_83__83_,chained_data_delayed_83__82_,
  chained_data_delayed_83__81_,chained_data_delayed_83__80_,
  chained_data_delayed_83__79_,chained_data_delayed_83__78_,chained_data_delayed_83__77_,
  chained_data_delayed_83__76_,chained_data_delayed_83__75_,chained_data_delayed_83__74_,
  chained_data_delayed_83__73_,chained_data_delayed_83__72_,chained_data_delayed_83__71_,
  chained_data_delayed_83__70_,chained_data_delayed_83__69_,chained_data_delayed_83__68_,
  chained_data_delayed_83__67_,chained_data_delayed_83__66_,
  chained_data_delayed_83__65_,chained_data_delayed_83__64_,chained_data_delayed_83__63_,
  chained_data_delayed_83__62_,chained_data_delayed_83__61_,chained_data_delayed_83__60_,
  chained_data_delayed_83__59_,chained_data_delayed_83__58_,chained_data_delayed_83__57_,
  chained_data_delayed_83__56_,chained_data_delayed_83__55_,
  chained_data_delayed_83__54_,chained_data_delayed_83__53_,chained_data_delayed_83__52_,
  chained_data_delayed_83__51_,chained_data_delayed_83__50_,chained_data_delayed_83__49_,
  chained_data_delayed_83__48_,chained_data_delayed_83__47_,chained_data_delayed_83__46_,
  chained_data_delayed_83__45_,chained_data_delayed_83__44_,
  chained_data_delayed_83__43_,chained_data_delayed_83__42_,chained_data_delayed_83__41_,
  chained_data_delayed_83__40_,chained_data_delayed_83__39_,chained_data_delayed_83__38_,
  chained_data_delayed_83__37_,chained_data_delayed_83__36_,chained_data_delayed_83__35_,
  chained_data_delayed_83__34_,chained_data_delayed_83__33_,
  chained_data_delayed_83__32_,chained_data_delayed_83__31_,chained_data_delayed_83__30_,
  chained_data_delayed_83__29_,chained_data_delayed_83__28_,chained_data_delayed_83__27_,
  chained_data_delayed_83__26_,chained_data_delayed_83__25_,chained_data_delayed_83__24_,
  chained_data_delayed_83__23_,chained_data_delayed_83__22_,
  chained_data_delayed_83__21_,chained_data_delayed_83__20_,chained_data_delayed_83__19_,
  chained_data_delayed_83__18_,chained_data_delayed_83__17_,chained_data_delayed_83__16_,
  chained_data_delayed_83__15_,chained_data_delayed_83__14_,chained_data_delayed_83__13_,
  chained_data_delayed_83__12_,chained_data_delayed_83__11_,
  chained_data_delayed_83__10_,chained_data_delayed_83__9_,chained_data_delayed_83__8_,
  chained_data_delayed_83__7_,chained_data_delayed_83__6_,chained_data_delayed_83__5_,
  chained_data_delayed_83__4_,chained_data_delayed_83__3_,chained_data_delayed_83__2_,
  chained_data_delayed_83__1_,chained_data_delayed_83__0_,chained_data_delayed_82__127_,
  chained_data_delayed_82__126_,chained_data_delayed_82__125_,
  chained_data_delayed_82__124_,chained_data_delayed_82__123_,chained_data_delayed_82__122_,
  chained_data_delayed_82__121_,chained_data_delayed_82__120_,chained_data_delayed_82__119_,
  chained_data_delayed_82__118_,chained_data_delayed_82__117_,
  chained_data_delayed_82__116_,chained_data_delayed_82__115_,chained_data_delayed_82__114_,
  chained_data_delayed_82__113_,chained_data_delayed_82__112_,chained_data_delayed_82__111_,
  chained_data_delayed_82__110_,chained_data_delayed_82__109_,
  chained_data_delayed_82__108_,chained_data_delayed_82__107_,chained_data_delayed_82__106_,
  chained_data_delayed_82__105_,chained_data_delayed_82__104_,chained_data_delayed_82__103_,
  chained_data_delayed_82__102_,chained_data_delayed_82__101_,
  chained_data_delayed_82__100_,chained_data_delayed_82__99_,chained_data_delayed_82__98_,
  chained_data_delayed_82__97_,chained_data_delayed_82__96_,chained_data_delayed_82__95_,
  chained_data_delayed_82__94_,chained_data_delayed_82__93_,chained_data_delayed_82__92_,
  chained_data_delayed_82__91_,chained_data_delayed_82__90_,
  chained_data_delayed_82__89_,chained_data_delayed_82__88_,chained_data_delayed_82__87_,
  chained_data_delayed_82__86_,chained_data_delayed_82__85_,chained_data_delayed_82__84_,
  chained_data_delayed_82__83_,chained_data_delayed_82__82_,chained_data_delayed_82__81_,
  chained_data_delayed_82__80_,chained_data_delayed_82__79_,chained_data_delayed_82__78_,
  chained_data_delayed_82__77_,chained_data_delayed_82__76_,
  chained_data_delayed_82__75_,chained_data_delayed_82__74_,chained_data_delayed_82__73_,
  chained_data_delayed_82__72_,chained_data_delayed_82__71_,chained_data_delayed_82__70_,
  chained_data_delayed_82__69_,chained_data_delayed_82__68_,chained_data_delayed_82__67_,
  chained_data_delayed_82__66_,chained_data_delayed_82__65_,
  chained_data_delayed_82__64_,chained_data_delayed_82__63_,chained_data_delayed_82__62_,
  chained_data_delayed_82__61_,chained_data_delayed_82__60_,chained_data_delayed_82__59_,
  chained_data_delayed_82__58_,chained_data_delayed_82__57_,chained_data_delayed_82__56_,
  chained_data_delayed_82__55_,chained_data_delayed_82__54_,
  chained_data_delayed_82__53_,chained_data_delayed_82__52_,chained_data_delayed_82__51_,
  chained_data_delayed_82__50_,chained_data_delayed_82__49_,chained_data_delayed_82__48_,
  chained_data_delayed_82__47_,chained_data_delayed_82__46_,chained_data_delayed_82__45_,
  chained_data_delayed_82__44_,chained_data_delayed_82__43_,
  chained_data_delayed_82__42_,chained_data_delayed_82__41_,chained_data_delayed_82__40_,
  chained_data_delayed_82__39_,chained_data_delayed_82__38_,chained_data_delayed_82__37_,
  chained_data_delayed_82__36_,chained_data_delayed_82__35_,chained_data_delayed_82__34_,
  chained_data_delayed_82__33_,chained_data_delayed_82__32_,
  chained_data_delayed_82__31_,chained_data_delayed_82__30_,chained_data_delayed_82__29_,
  chained_data_delayed_82__28_,chained_data_delayed_82__27_,chained_data_delayed_82__26_,
  chained_data_delayed_82__25_,chained_data_delayed_82__24_,chained_data_delayed_82__23_,
  chained_data_delayed_82__22_,chained_data_delayed_82__21_,
  chained_data_delayed_82__20_,chained_data_delayed_82__19_,chained_data_delayed_82__18_,
  chained_data_delayed_82__17_,chained_data_delayed_82__16_,chained_data_delayed_82__15_,
  chained_data_delayed_82__14_,chained_data_delayed_82__13_,chained_data_delayed_82__12_,
  chained_data_delayed_82__11_,chained_data_delayed_82__10_,chained_data_delayed_82__9_,
  chained_data_delayed_82__8_,chained_data_delayed_82__7_,
  chained_data_delayed_82__6_,chained_data_delayed_82__5_,chained_data_delayed_82__4_,
  chained_data_delayed_82__3_,chained_data_delayed_82__2_,chained_data_delayed_82__1_,
  chained_data_delayed_82__0_,chained_data_delayed_81__127_,chained_data_delayed_81__126_,
  chained_data_delayed_81__125_,chained_data_delayed_81__124_,
  chained_data_delayed_81__123_,chained_data_delayed_81__122_,chained_data_delayed_81__121_,
  chained_data_delayed_81__120_,chained_data_delayed_81__119_,chained_data_delayed_81__118_,
  chained_data_delayed_81__117_,chained_data_delayed_81__116_,
  chained_data_delayed_81__115_,chained_data_delayed_81__114_,chained_data_delayed_81__113_,
  chained_data_delayed_81__112_,chained_data_delayed_81__111_,chained_data_delayed_81__110_,
  chained_data_delayed_81__109_,chained_data_delayed_81__108_,
  chained_data_delayed_81__107_,chained_data_delayed_81__106_,chained_data_delayed_81__105_,
  chained_data_delayed_81__104_,chained_data_delayed_81__103_,chained_data_delayed_81__102_,
  chained_data_delayed_81__101_,chained_data_delayed_81__100_,
  chained_data_delayed_81__99_,chained_data_delayed_81__98_,chained_data_delayed_81__97_,
  chained_data_delayed_81__96_,chained_data_delayed_81__95_,chained_data_delayed_81__94_,
  chained_data_delayed_81__93_,chained_data_delayed_81__92_,chained_data_delayed_81__91_,
  chained_data_delayed_81__90_,chained_data_delayed_81__89_,chained_data_delayed_81__88_,
  chained_data_delayed_81__87_,chained_data_delayed_81__86_,
  chained_data_delayed_81__85_,chained_data_delayed_81__84_,chained_data_delayed_81__83_,
  chained_data_delayed_81__82_,chained_data_delayed_81__81_,chained_data_delayed_81__80_,
  chained_data_delayed_81__79_,chained_data_delayed_81__78_,chained_data_delayed_81__77_,
  chained_data_delayed_81__76_,chained_data_delayed_81__75_,
  chained_data_delayed_81__74_,chained_data_delayed_81__73_,chained_data_delayed_81__72_,
  chained_data_delayed_81__71_,chained_data_delayed_81__70_,chained_data_delayed_81__69_,
  chained_data_delayed_81__68_,chained_data_delayed_81__67_,chained_data_delayed_81__66_,
  chained_data_delayed_81__65_,chained_data_delayed_81__64_,
  chained_data_delayed_81__63_,chained_data_delayed_81__62_,chained_data_delayed_81__61_,
  chained_data_delayed_81__60_,chained_data_delayed_81__59_,chained_data_delayed_81__58_,
  chained_data_delayed_81__57_,chained_data_delayed_81__56_,chained_data_delayed_81__55_,
  chained_data_delayed_81__54_,chained_data_delayed_81__53_,
  chained_data_delayed_81__52_,chained_data_delayed_81__51_,chained_data_delayed_81__50_,
  chained_data_delayed_81__49_,chained_data_delayed_81__48_,chained_data_delayed_81__47_,
  chained_data_delayed_81__46_,chained_data_delayed_81__45_,chained_data_delayed_81__44_,
  chained_data_delayed_81__43_,chained_data_delayed_81__42_,
  chained_data_delayed_81__41_,chained_data_delayed_81__40_,chained_data_delayed_81__39_,
  chained_data_delayed_81__38_,chained_data_delayed_81__37_,chained_data_delayed_81__36_,
  chained_data_delayed_81__35_,chained_data_delayed_81__34_,chained_data_delayed_81__33_,
  chained_data_delayed_81__32_,chained_data_delayed_81__31_,
  chained_data_delayed_81__30_,chained_data_delayed_81__29_,chained_data_delayed_81__28_,
  chained_data_delayed_81__27_,chained_data_delayed_81__26_,chained_data_delayed_81__25_,
  chained_data_delayed_81__24_,chained_data_delayed_81__23_,chained_data_delayed_81__22_,
  chained_data_delayed_81__21_,chained_data_delayed_81__20_,
  chained_data_delayed_81__19_,chained_data_delayed_81__18_,chained_data_delayed_81__17_,
  chained_data_delayed_81__16_,chained_data_delayed_81__15_,chained_data_delayed_81__14_,
  chained_data_delayed_81__13_,chained_data_delayed_81__12_,chained_data_delayed_81__11_,
  chained_data_delayed_81__10_,chained_data_delayed_81__9_,chained_data_delayed_81__8_,
  chained_data_delayed_81__7_,chained_data_delayed_81__6_,
  chained_data_delayed_81__5_,chained_data_delayed_81__4_,chained_data_delayed_81__3_,
  chained_data_delayed_81__2_,chained_data_delayed_81__1_,chained_data_delayed_81__0_,
  chained_data_delayed_88__127_,chained_data_delayed_88__126_,chained_data_delayed_88__125_,
  chained_data_delayed_88__124_,chained_data_delayed_88__123_,
  chained_data_delayed_88__122_,chained_data_delayed_88__121_,chained_data_delayed_88__120_,
  chained_data_delayed_88__119_,chained_data_delayed_88__118_,chained_data_delayed_88__117_,
  chained_data_delayed_88__116_,chained_data_delayed_88__115_,
  chained_data_delayed_88__114_,chained_data_delayed_88__113_,chained_data_delayed_88__112_,
  chained_data_delayed_88__111_,chained_data_delayed_88__110_,chained_data_delayed_88__109_,
  chained_data_delayed_88__108_,chained_data_delayed_88__107_,
  chained_data_delayed_88__106_,chained_data_delayed_88__105_,chained_data_delayed_88__104_,
  chained_data_delayed_88__103_,chained_data_delayed_88__102_,chained_data_delayed_88__101_,
  chained_data_delayed_88__100_,chained_data_delayed_88__99_,chained_data_delayed_88__98_,
  chained_data_delayed_88__97_,chained_data_delayed_88__96_,
  chained_data_delayed_88__95_,chained_data_delayed_88__94_,chained_data_delayed_88__93_,
  chained_data_delayed_88__92_,chained_data_delayed_88__91_,chained_data_delayed_88__90_,
  chained_data_delayed_88__89_,chained_data_delayed_88__88_,chained_data_delayed_88__87_,
  chained_data_delayed_88__86_,chained_data_delayed_88__85_,
  chained_data_delayed_88__84_,chained_data_delayed_88__83_,chained_data_delayed_88__82_,
  chained_data_delayed_88__81_,chained_data_delayed_88__80_,chained_data_delayed_88__79_,
  chained_data_delayed_88__78_,chained_data_delayed_88__77_,chained_data_delayed_88__76_,
  chained_data_delayed_88__75_,chained_data_delayed_88__74_,
  chained_data_delayed_88__73_,chained_data_delayed_88__72_,chained_data_delayed_88__71_,
  chained_data_delayed_88__70_,chained_data_delayed_88__69_,chained_data_delayed_88__68_,
  chained_data_delayed_88__67_,chained_data_delayed_88__66_,chained_data_delayed_88__65_,
  chained_data_delayed_88__64_,chained_data_delayed_88__63_,
  chained_data_delayed_88__62_,chained_data_delayed_88__61_,chained_data_delayed_88__60_,
  chained_data_delayed_88__59_,chained_data_delayed_88__58_,chained_data_delayed_88__57_,
  chained_data_delayed_88__56_,chained_data_delayed_88__55_,chained_data_delayed_88__54_,
  chained_data_delayed_88__53_,chained_data_delayed_88__52_,
  chained_data_delayed_88__51_,chained_data_delayed_88__50_,chained_data_delayed_88__49_,
  chained_data_delayed_88__48_,chained_data_delayed_88__47_,chained_data_delayed_88__46_,
  chained_data_delayed_88__45_,chained_data_delayed_88__44_,chained_data_delayed_88__43_,
  chained_data_delayed_88__42_,chained_data_delayed_88__41_,
  chained_data_delayed_88__40_,chained_data_delayed_88__39_,chained_data_delayed_88__38_,
  chained_data_delayed_88__37_,chained_data_delayed_88__36_,chained_data_delayed_88__35_,
  chained_data_delayed_88__34_,chained_data_delayed_88__33_,chained_data_delayed_88__32_,
  chained_data_delayed_88__31_,chained_data_delayed_88__30_,
  chained_data_delayed_88__29_,chained_data_delayed_88__28_,chained_data_delayed_88__27_,
  chained_data_delayed_88__26_,chained_data_delayed_88__25_,chained_data_delayed_88__24_,
  chained_data_delayed_88__23_,chained_data_delayed_88__22_,chained_data_delayed_88__21_,
  chained_data_delayed_88__20_,chained_data_delayed_88__19_,chained_data_delayed_88__18_,
  chained_data_delayed_88__17_,chained_data_delayed_88__16_,
  chained_data_delayed_88__15_,chained_data_delayed_88__14_,chained_data_delayed_88__13_,
  chained_data_delayed_88__12_,chained_data_delayed_88__11_,chained_data_delayed_88__10_,
  chained_data_delayed_88__9_,chained_data_delayed_88__8_,chained_data_delayed_88__7_,
  chained_data_delayed_88__6_,chained_data_delayed_88__5_,chained_data_delayed_88__4_,
  chained_data_delayed_88__3_,chained_data_delayed_88__2_,
  chained_data_delayed_88__1_,chained_data_delayed_88__0_,chained_data_delayed_87__127_,
  chained_data_delayed_87__126_,chained_data_delayed_87__125_,chained_data_delayed_87__124_,
  chained_data_delayed_87__123_,chained_data_delayed_87__122_,
  chained_data_delayed_87__121_,chained_data_delayed_87__120_,chained_data_delayed_87__119_,
  chained_data_delayed_87__118_,chained_data_delayed_87__117_,chained_data_delayed_87__116_,
  chained_data_delayed_87__115_,chained_data_delayed_87__114_,
  chained_data_delayed_87__113_,chained_data_delayed_87__112_,chained_data_delayed_87__111_,
  chained_data_delayed_87__110_,chained_data_delayed_87__109_,chained_data_delayed_87__108_,
  chained_data_delayed_87__107_,chained_data_delayed_87__106_,
  chained_data_delayed_87__105_,chained_data_delayed_87__104_,chained_data_delayed_87__103_,
  chained_data_delayed_87__102_,chained_data_delayed_87__101_,chained_data_delayed_87__100_,
  chained_data_delayed_87__99_,chained_data_delayed_87__98_,chained_data_delayed_87__97_,
  chained_data_delayed_87__96_,chained_data_delayed_87__95_,
  chained_data_delayed_87__94_,chained_data_delayed_87__93_,chained_data_delayed_87__92_,
  chained_data_delayed_87__91_,chained_data_delayed_87__90_,chained_data_delayed_87__89_,
  chained_data_delayed_87__88_,chained_data_delayed_87__87_,chained_data_delayed_87__86_,
  chained_data_delayed_87__85_,chained_data_delayed_87__84_,
  chained_data_delayed_87__83_,chained_data_delayed_87__82_,chained_data_delayed_87__81_,
  chained_data_delayed_87__80_,chained_data_delayed_87__79_,chained_data_delayed_87__78_,
  chained_data_delayed_87__77_,chained_data_delayed_87__76_,chained_data_delayed_87__75_,
  chained_data_delayed_87__74_,chained_data_delayed_87__73_,
  chained_data_delayed_87__72_,chained_data_delayed_87__71_,chained_data_delayed_87__70_,
  chained_data_delayed_87__69_,chained_data_delayed_87__68_,chained_data_delayed_87__67_,
  chained_data_delayed_87__66_,chained_data_delayed_87__65_,chained_data_delayed_87__64_,
  chained_data_delayed_87__63_,chained_data_delayed_87__62_,
  chained_data_delayed_87__61_,chained_data_delayed_87__60_,chained_data_delayed_87__59_,
  chained_data_delayed_87__58_,chained_data_delayed_87__57_,chained_data_delayed_87__56_,
  chained_data_delayed_87__55_,chained_data_delayed_87__54_,chained_data_delayed_87__53_,
  chained_data_delayed_87__52_,chained_data_delayed_87__51_,
  chained_data_delayed_87__50_,chained_data_delayed_87__49_,chained_data_delayed_87__48_,
  chained_data_delayed_87__47_,chained_data_delayed_87__46_,chained_data_delayed_87__45_,
  chained_data_delayed_87__44_,chained_data_delayed_87__43_,chained_data_delayed_87__42_,
  chained_data_delayed_87__41_,chained_data_delayed_87__40_,
  chained_data_delayed_87__39_,chained_data_delayed_87__38_,chained_data_delayed_87__37_,
  chained_data_delayed_87__36_,chained_data_delayed_87__35_,chained_data_delayed_87__34_,
  chained_data_delayed_87__33_,chained_data_delayed_87__32_,chained_data_delayed_87__31_,
  chained_data_delayed_87__30_,chained_data_delayed_87__29_,chained_data_delayed_87__28_,
  chained_data_delayed_87__27_,chained_data_delayed_87__26_,
  chained_data_delayed_87__25_,chained_data_delayed_87__24_,chained_data_delayed_87__23_,
  chained_data_delayed_87__22_,chained_data_delayed_87__21_,chained_data_delayed_87__20_,
  chained_data_delayed_87__19_,chained_data_delayed_87__18_,chained_data_delayed_87__17_,
  chained_data_delayed_87__16_,chained_data_delayed_87__15_,
  chained_data_delayed_87__14_,chained_data_delayed_87__13_,chained_data_delayed_87__12_,
  chained_data_delayed_87__11_,chained_data_delayed_87__10_,chained_data_delayed_87__9_,
  chained_data_delayed_87__8_,chained_data_delayed_87__7_,chained_data_delayed_87__6_,
  chained_data_delayed_87__5_,chained_data_delayed_87__4_,chained_data_delayed_87__3_,
  chained_data_delayed_87__2_,chained_data_delayed_87__1_,
  chained_data_delayed_87__0_,chained_data_delayed_86__127_,chained_data_delayed_86__126_,
  chained_data_delayed_86__125_,chained_data_delayed_86__124_,chained_data_delayed_86__123_,
  chained_data_delayed_86__122_,chained_data_delayed_86__121_,
  chained_data_delayed_86__120_,chained_data_delayed_86__119_,chained_data_delayed_86__118_,
  chained_data_delayed_86__117_,chained_data_delayed_86__116_,chained_data_delayed_86__115_,
  chained_data_delayed_86__114_,chained_data_delayed_86__113_,
  chained_data_delayed_86__112_,chained_data_delayed_86__111_,chained_data_delayed_86__110_,
  chained_data_delayed_86__109_,chained_data_delayed_86__108_,chained_data_delayed_86__107_,
  chained_data_delayed_86__106_,chained_data_delayed_86__105_,
  chained_data_delayed_86__104_,chained_data_delayed_86__103_,chained_data_delayed_86__102_,
  chained_data_delayed_86__101_,chained_data_delayed_86__100_,chained_data_delayed_86__99_,
  chained_data_delayed_86__98_,chained_data_delayed_86__97_,chained_data_delayed_86__96_,
  chained_data_delayed_86__95_,chained_data_delayed_86__94_,
  chained_data_delayed_86__93_,chained_data_delayed_86__92_,chained_data_delayed_86__91_,
  chained_data_delayed_86__90_,chained_data_delayed_86__89_,chained_data_delayed_86__88_,
  chained_data_delayed_86__87_,chained_data_delayed_86__86_,chained_data_delayed_86__85_,
  chained_data_delayed_86__84_,chained_data_delayed_86__83_,
  chained_data_delayed_86__82_,chained_data_delayed_86__81_,chained_data_delayed_86__80_,
  chained_data_delayed_86__79_,chained_data_delayed_86__78_,chained_data_delayed_86__77_,
  chained_data_delayed_86__76_,chained_data_delayed_86__75_,chained_data_delayed_86__74_,
  chained_data_delayed_86__73_,chained_data_delayed_86__72_,
  chained_data_delayed_86__71_,chained_data_delayed_86__70_,chained_data_delayed_86__69_,
  chained_data_delayed_86__68_,chained_data_delayed_86__67_,chained_data_delayed_86__66_,
  chained_data_delayed_86__65_,chained_data_delayed_86__64_,chained_data_delayed_86__63_,
  chained_data_delayed_86__62_,chained_data_delayed_86__61_,
  chained_data_delayed_86__60_,chained_data_delayed_86__59_,chained_data_delayed_86__58_,
  chained_data_delayed_86__57_,chained_data_delayed_86__56_,chained_data_delayed_86__55_,
  chained_data_delayed_86__54_,chained_data_delayed_86__53_,chained_data_delayed_86__52_,
  chained_data_delayed_86__51_,chained_data_delayed_86__50_,
  chained_data_delayed_86__49_,chained_data_delayed_86__48_,chained_data_delayed_86__47_,
  chained_data_delayed_86__46_,chained_data_delayed_86__45_,chained_data_delayed_86__44_,
  chained_data_delayed_86__43_,chained_data_delayed_86__42_,chained_data_delayed_86__41_,
  chained_data_delayed_86__40_,chained_data_delayed_86__39_,chained_data_delayed_86__38_,
  chained_data_delayed_86__37_,chained_data_delayed_86__36_,
  chained_data_delayed_86__35_,chained_data_delayed_86__34_,chained_data_delayed_86__33_,
  chained_data_delayed_86__32_,chained_data_delayed_86__31_,chained_data_delayed_86__30_,
  chained_data_delayed_86__29_,chained_data_delayed_86__28_,chained_data_delayed_86__27_,
  chained_data_delayed_86__26_,chained_data_delayed_86__25_,
  chained_data_delayed_86__24_,chained_data_delayed_86__23_,chained_data_delayed_86__22_,
  chained_data_delayed_86__21_,chained_data_delayed_86__20_,chained_data_delayed_86__19_,
  chained_data_delayed_86__18_,chained_data_delayed_86__17_,chained_data_delayed_86__16_,
  chained_data_delayed_86__15_,chained_data_delayed_86__14_,
  chained_data_delayed_86__13_,chained_data_delayed_86__12_,chained_data_delayed_86__11_,
  chained_data_delayed_86__10_,chained_data_delayed_86__9_,chained_data_delayed_86__8_,
  chained_data_delayed_86__7_,chained_data_delayed_86__6_,chained_data_delayed_86__5_,
  chained_data_delayed_86__4_,chained_data_delayed_86__3_,chained_data_delayed_86__2_,
  chained_data_delayed_86__1_,chained_data_delayed_86__0_,
  chained_data_delayed_85__127_,chained_data_delayed_85__126_,chained_data_delayed_85__125_,
  chained_data_delayed_85__124_,chained_data_delayed_85__123_,chained_data_delayed_85__122_,
  chained_data_delayed_85__121_,chained_data_delayed_85__120_,
  chained_data_delayed_85__119_,chained_data_delayed_85__118_,chained_data_delayed_85__117_,
  chained_data_delayed_85__116_,chained_data_delayed_85__115_,chained_data_delayed_85__114_,
  chained_data_delayed_85__113_,chained_data_delayed_85__112_,
  chained_data_delayed_85__111_,chained_data_delayed_85__110_,chained_data_delayed_85__109_,
  chained_data_delayed_85__108_,chained_data_delayed_85__107_,chained_data_delayed_85__106_,
  chained_data_delayed_85__105_,chained_data_delayed_85__104_,
  chained_data_delayed_85__103_,chained_data_delayed_85__102_,chained_data_delayed_85__101_,
  chained_data_delayed_85__100_,chained_data_delayed_85__99_,chained_data_delayed_85__98_,
  chained_data_delayed_85__97_,chained_data_delayed_85__96_,chained_data_delayed_85__95_,
  chained_data_delayed_85__94_,chained_data_delayed_85__93_,
  chained_data_delayed_85__92_,chained_data_delayed_85__91_,chained_data_delayed_85__90_,
  chained_data_delayed_85__89_,chained_data_delayed_85__88_,chained_data_delayed_85__87_,
  chained_data_delayed_85__86_,chained_data_delayed_85__85_,chained_data_delayed_85__84_,
  chained_data_delayed_85__83_,chained_data_delayed_85__82_,
  chained_data_delayed_85__81_,chained_data_delayed_85__80_,chained_data_delayed_85__79_,
  chained_data_delayed_85__78_,chained_data_delayed_85__77_,chained_data_delayed_85__76_,
  chained_data_delayed_85__75_,chained_data_delayed_85__74_,chained_data_delayed_85__73_,
  chained_data_delayed_85__72_,chained_data_delayed_85__71_,
  chained_data_delayed_85__70_,chained_data_delayed_85__69_,chained_data_delayed_85__68_,
  chained_data_delayed_85__67_,chained_data_delayed_85__66_,chained_data_delayed_85__65_,
  chained_data_delayed_85__64_,chained_data_delayed_85__63_,chained_data_delayed_85__62_,
  chained_data_delayed_85__61_,chained_data_delayed_85__60_,
  chained_data_delayed_85__59_,chained_data_delayed_85__58_,chained_data_delayed_85__57_,
  chained_data_delayed_85__56_,chained_data_delayed_85__55_,chained_data_delayed_85__54_,
  chained_data_delayed_85__53_,chained_data_delayed_85__52_,chained_data_delayed_85__51_,
  chained_data_delayed_85__50_,chained_data_delayed_85__49_,chained_data_delayed_85__48_,
  chained_data_delayed_85__47_,chained_data_delayed_85__46_,
  chained_data_delayed_85__45_,chained_data_delayed_85__44_,chained_data_delayed_85__43_,
  chained_data_delayed_85__42_,chained_data_delayed_85__41_,chained_data_delayed_85__40_,
  chained_data_delayed_85__39_,chained_data_delayed_85__38_,chained_data_delayed_85__37_,
  chained_data_delayed_85__36_,chained_data_delayed_85__35_,
  chained_data_delayed_85__34_,chained_data_delayed_85__33_,chained_data_delayed_85__32_,
  chained_data_delayed_85__31_,chained_data_delayed_85__30_,chained_data_delayed_85__29_,
  chained_data_delayed_85__28_,chained_data_delayed_85__27_,chained_data_delayed_85__26_,
  chained_data_delayed_85__25_,chained_data_delayed_85__24_,
  chained_data_delayed_85__23_,chained_data_delayed_85__22_,chained_data_delayed_85__21_,
  chained_data_delayed_85__20_,chained_data_delayed_85__19_,chained_data_delayed_85__18_,
  chained_data_delayed_85__17_,chained_data_delayed_85__16_,chained_data_delayed_85__15_,
  chained_data_delayed_85__14_,chained_data_delayed_85__13_,
  chained_data_delayed_85__12_,chained_data_delayed_85__11_,chained_data_delayed_85__10_,
  chained_data_delayed_85__9_,chained_data_delayed_85__8_,chained_data_delayed_85__7_,
  chained_data_delayed_85__6_,chained_data_delayed_85__5_,chained_data_delayed_85__4_,
  chained_data_delayed_85__3_,chained_data_delayed_85__2_,chained_data_delayed_85__1_,
  chained_data_delayed_85__0_,chained_data_delayed_92__127_,
  chained_data_delayed_92__126_,chained_data_delayed_92__125_,chained_data_delayed_92__124_,
  chained_data_delayed_92__123_,chained_data_delayed_92__122_,chained_data_delayed_92__121_,
  chained_data_delayed_92__120_,chained_data_delayed_92__119_,
  chained_data_delayed_92__118_,chained_data_delayed_92__117_,chained_data_delayed_92__116_,
  chained_data_delayed_92__115_,chained_data_delayed_92__114_,chained_data_delayed_92__113_,
  chained_data_delayed_92__112_,chained_data_delayed_92__111_,
  chained_data_delayed_92__110_,chained_data_delayed_92__109_,chained_data_delayed_92__108_,
  chained_data_delayed_92__107_,chained_data_delayed_92__106_,chained_data_delayed_92__105_,
  chained_data_delayed_92__104_,chained_data_delayed_92__103_,
  chained_data_delayed_92__102_,chained_data_delayed_92__101_,chained_data_delayed_92__100_,
  chained_data_delayed_92__99_,chained_data_delayed_92__98_,chained_data_delayed_92__97_,
  chained_data_delayed_92__96_,chained_data_delayed_92__95_,chained_data_delayed_92__94_,
  chained_data_delayed_92__93_,chained_data_delayed_92__92_,
  chained_data_delayed_92__91_,chained_data_delayed_92__90_,chained_data_delayed_92__89_,
  chained_data_delayed_92__88_,chained_data_delayed_92__87_,chained_data_delayed_92__86_,
  chained_data_delayed_92__85_,chained_data_delayed_92__84_,chained_data_delayed_92__83_,
  chained_data_delayed_92__82_,chained_data_delayed_92__81_,
  chained_data_delayed_92__80_,chained_data_delayed_92__79_,chained_data_delayed_92__78_,
  chained_data_delayed_92__77_,chained_data_delayed_92__76_,chained_data_delayed_92__75_,
  chained_data_delayed_92__74_,chained_data_delayed_92__73_,chained_data_delayed_92__72_,
  chained_data_delayed_92__71_,chained_data_delayed_92__70_,
  chained_data_delayed_92__69_,chained_data_delayed_92__68_,chained_data_delayed_92__67_,
  chained_data_delayed_92__66_,chained_data_delayed_92__65_,chained_data_delayed_92__64_,
  chained_data_delayed_92__63_,chained_data_delayed_92__62_,chained_data_delayed_92__61_,
  chained_data_delayed_92__60_,chained_data_delayed_92__59_,chained_data_delayed_92__58_,
  chained_data_delayed_92__57_,chained_data_delayed_92__56_,
  chained_data_delayed_92__55_,chained_data_delayed_92__54_,chained_data_delayed_92__53_,
  chained_data_delayed_92__52_,chained_data_delayed_92__51_,chained_data_delayed_92__50_,
  chained_data_delayed_92__49_,chained_data_delayed_92__48_,chained_data_delayed_92__47_,
  chained_data_delayed_92__46_,chained_data_delayed_92__45_,
  chained_data_delayed_92__44_,chained_data_delayed_92__43_,chained_data_delayed_92__42_,
  chained_data_delayed_92__41_,chained_data_delayed_92__40_,chained_data_delayed_92__39_,
  chained_data_delayed_92__38_,chained_data_delayed_92__37_,chained_data_delayed_92__36_,
  chained_data_delayed_92__35_,chained_data_delayed_92__34_,
  chained_data_delayed_92__33_,chained_data_delayed_92__32_,chained_data_delayed_92__31_,
  chained_data_delayed_92__30_,chained_data_delayed_92__29_,chained_data_delayed_92__28_,
  chained_data_delayed_92__27_,chained_data_delayed_92__26_,chained_data_delayed_92__25_,
  chained_data_delayed_92__24_,chained_data_delayed_92__23_,
  chained_data_delayed_92__22_,chained_data_delayed_92__21_,chained_data_delayed_92__20_,
  chained_data_delayed_92__19_,chained_data_delayed_92__18_,chained_data_delayed_92__17_,
  chained_data_delayed_92__16_,chained_data_delayed_92__15_,chained_data_delayed_92__14_,
  chained_data_delayed_92__13_,chained_data_delayed_92__12_,
  chained_data_delayed_92__11_,chained_data_delayed_92__10_,chained_data_delayed_92__9_,
  chained_data_delayed_92__8_,chained_data_delayed_92__7_,chained_data_delayed_92__6_,
  chained_data_delayed_92__5_,chained_data_delayed_92__4_,chained_data_delayed_92__3_,
  chained_data_delayed_92__2_,chained_data_delayed_92__1_,chained_data_delayed_92__0_,
  chained_data_delayed_91__127_,chained_data_delayed_91__126_,
  chained_data_delayed_91__125_,chained_data_delayed_91__124_,chained_data_delayed_91__123_,
  chained_data_delayed_91__122_,chained_data_delayed_91__121_,chained_data_delayed_91__120_,
  chained_data_delayed_91__119_,chained_data_delayed_91__118_,
  chained_data_delayed_91__117_,chained_data_delayed_91__116_,chained_data_delayed_91__115_,
  chained_data_delayed_91__114_,chained_data_delayed_91__113_,chained_data_delayed_91__112_,
  chained_data_delayed_91__111_,chained_data_delayed_91__110_,
  chained_data_delayed_91__109_,chained_data_delayed_91__108_,chained_data_delayed_91__107_,
  chained_data_delayed_91__106_,chained_data_delayed_91__105_,chained_data_delayed_91__104_,
  chained_data_delayed_91__103_,chained_data_delayed_91__102_,
  chained_data_delayed_91__101_,chained_data_delayed_91__100_,chained_data_delayed_91__99_,
  chained_data_delayed_91__98_,chained_data_delayed_91__97_,chained_data_delayed_91__96_,
  chained_data_delayed_91__95_,chained_data_delayed_91__94_,chained_data_delayed_91__93_,
  chained_data_delayed_91__92_,chained_data_delayed_91__91_,
  chained_data_delayed_91__90_,chained_data_delayed_91__89_,chained_data_delayed_91__88_,
  chained_data_delayed_91__87_,chained_data_delayed_91__86_,chained_data_delayed_91__85_,
  chained_data_delayed_91__84_,chained_data_delayed_91__83_,chained_data_delayed_91__82_,
  chained_data_delayed_91__81_,chained_data_delayed_91__80_,
  chained_data_delayed_91__79_,chained_data_delayed_91__78_,chained_data_delayed_91__77_,
  chained_data_delayed_91__76_,chained_data_delayed_91__75_,chained_data_delayed_91__74_,
  chained_data_delayed_91__73_,chained_data_delayed_91__72_,chained_data_delayed_91__71_,
  chained_data_delayed_91__70_,chained_data_delayed_91__69_,chained_data_delayed_91__68_,
  chained_data_delayed_91__67_,chained_data_delayed_91__66_,
  chained_data_delayed_91__65_,chained_data_delayed_91__64_,chained_data_delayed_91__63_,
  chained_data_delayed_91__62_,chained_data_delayed_91__61_,chained_data_delayed_91__60_,
  chained_data_delayed_91__59_,chained_data_delayed_91__58_,chained_data_delayed_91__57_,
  chained_data_delayed_91__56_,chained_data_delayed_91__55_,
  chained_data_delayed_91__54_,chained_data_delayed_91__53_,chained_data_delayed_91__52_,
  chained_data_delayed_91__51_,chained_data_delayed_91__50_,chained_data_delayed_91__49_,
  chained_data_delayed_91__48_,chained_data_delayed_91__47_,chained_data_delayed_91__46_,
  chained_data_delayed_91__45_,chained_data_delayed_91__44_,
  chained_data_delayed_91__43_,chained_data_delayed_91__42_,chained_data_delayed_91__41_,
  chained_data_delayed_91__40_,chained_data_delayed_91__39_,chained_data_delayed_91__38_,
  chained_data_delayed_91__37_,chained_data_delayed_91__36_,chained_data_delayed_91__35_,
  chained_data_delayed_91__34_,chained_data_delayed_91__33_,
  chained_data_delayed_91__32_,chained_data_delayed_91__31_,chained_data_delayed_91__30_,
  chained_data_delayed_91__29_,chained_data_delayed_91__28_,chained_data_delayed_91__27_,
  chained_data_delayed_91__26_,chained_data_delayed_91__25_,chained_data_delayed_91__24_,
  chained_data_delayed_91__23_,chained_data_delayed_91__22_,
  chained_data_delayed_91__21_,chained_data_delayed_91__20_,chained_data_delayed_91__19_,
  chained_data_delayed_91__18_,chained_data_delayed_91__17_,chained_data_delayed_91__16_,
  chained_data_delayed_91__15_,chained_data_delayed_91__14_,chained_data_delayed_91__13_,
  chained_data_delayed_91__12_,chained_data_delayed_91__11_,
  chained_data_delayed_91__10_,chained_data_delayed_91__9_,chained_data_delayed_91__8_,
  chained_data_delayed_91__7_,chained_data_delayed_91__6_,chained_data_delayed_91__5_,
  chained_data_delayed_91__4_,chained_data_delayed_91__3_,chained_data_delayed_91__2_,
  chained_data_delayed_91__1_,chained_data_delayed_91__0_,chained_data_delayed_90__127_,
  chained_data_delayed_90__126_,chained_data_delayed_90__125_,
  chained_data_delayed_90__124_,chained_data_delayed_90__123_,chained_data_delayed_90__122_,
  chained_data_delayed_90__121_,chained_data_delayed_90__120_,chained_data_delayed_90__119_,
  chained_data_delayed_90__118_,chained_data_delayed_90__117_,
  chained_data_delayed_90__116_,chained_data_delayed_90__115_,chained_data_delayed_90__114_,
  chained_data_delayed_90__113_,chained_data_delayed_90__112_,chained_data_delayed_90__111_,
  chained_data_delayed_90__110_,chained_data_delayed_90__109_,
  chained_data_delayed_90__108_,chained_data_delayed_90__107_,chained_data_delayed_90__106_,
  chained_data_delayed_90__105_,chained_data_delayed_90__104_,chained_data_delayed_90__103_,
  chained_data_delayed_90__102_,chained_data_delayed_90__101_,
  chained_data_delayed_90__100_,chained_data_delayed_90__99_,chained_data_delayed_90__98_,
  chained_data_delayed_90__97_,chained_data_delayed_90__96_,chained_data_delayed_90__95_,
  chained_data_delayed_90__94_,chained_data_delayed_90__93_,chained_data_delayed_90__92_,
  chained_data_delayed_90__91_,chained_data_delayed_90__90_,
  chained_data_delayed_90__89_,chained_data_delayed_90__88_,chained_data_delayed_90__87_,
  chained_data_delayed_90__86_,chained_data_delayed_90__85_,chained_data_delayed_90__84_,
  chained_data_delayed_90__83_,chained_data_delayed_90__82_,chained_data_delayed_90__81_,
  chained_data_delayed_90__80_,chained_data_delayed_90__79_,chained_data_delayed_90__78_,
  chained_data_delayed_90__77_,chained_data_delayed_90__76_,
  chained_data_delayed_90__75_,chained_data_delayed_90__74_,chained_data_delayed_90__73_,
  chained_data_delayed_90__72_,chained_data_delayed_90__71_,chained_data_delayed_90__70_,
  chained_data_delayed_90__69_,chained_data_delayed_90__68_,chained_data_delayed_90__67_,
  chained_data_delayed_90__66_,chained_data_delayed_90__65_,
  chained_data_delayed_90__64_,chained_data_delayed_90__63_,chained_data_delayed_90__62_,
  chained_data_delayed_90__61_,chained_data_delayed_90__60_,chained_data_delayed_90__59_,
  chained_data_delayed_90__58_,chained_data_delayed_90__57_,chained_data_delayed_90__56_,
  chained_data_delayed_90__55_,chained_data_delayed_90__54_,
  chained_data_delayed_90__53_,chained_data_delayed_90__52_,chained_data_delayed_90__51_,
  chained_data_delayed_90__50_,chained_data_delayed_90__49_,chained_data_delayed_90__48_,
  chained_data_delayed_90__47_,chained_data_delayed_90__46_,chained_data_delayed_90__45_,
  chained_data_delayed_90__44_,chained_data_delayed_90__43_,
  chained_data_delayed_90__42_,chained_data_delayed_90__41_,chained_data_delayed_90__40_,
  chained_data_delayed_90__39_,chained_data_delayed_90__38_,chained_data_delayed_90__37_,
  chained_data_delayed_90__36_,chained_data_delayed_90__35_,chained_data_delayed_90__34_,
  chained_data_delayed_90__33_,chained_data_delayed_90__32_,
  chained_data_delayed_90__31_,chained_data_delayed_90__30_,chained_data_delayed_90__29_,
  chained_data_delayed_90__28_,chained_data_delayed_90__27_,chained_data_delayed_90__26_,
  chained_data_delayed_90__25_,chained_data_delayed_90__24_,chained_data_delayed_90__23_,
  chained_data_delayed_90__22_,chained_data_delayed_90__21_,
  chained_data_delayed_90__20_,chained_data_delayed_90__19_,chained_data_delayed_90__18_,
  chained_data_delayed_90__17_,chained_data_delayed_90__16_,chained_data_delayed_90__15_,
  chained_data_delayed_90__14_,chained_data_delayed_90__13_,chained_data_delayed_90__12_,
  chained_data_delayed_90__11_,chained_data_delayed_90__10_,chained_data_delayed_90__9_,
  chained_data_delayed_90__8_,chained_data_delayed_90__7_,
  chained_data_delayed_90__6_,chained_data_delayed_90__5_,chained_data_delayed_90__4_,
  chained_data_delayed_90__3_,chained_data_delayed_90__2_,chained_data_delayed_90__1_,
  chained_data_delayed_90__0_,chained_data_delayed_89__127_,chained_data_delayed_89__126_,
  chained_data_delayed_89__125_,chained_data_delayed_89__124_,
  chained_data_delayed_89__123_,chained_data_delayed_89__122_,chained_data_delayed_89__121_,
  chained_data_delayed_89__120_,chained_data_delayed_89__119_,chained_data_delayed_89__118_,
  chained_data_delayed_89__117_,chained_data_delayed_89__116_,
  chained_data_delayed_89__115_,chained_data_delayed_89__114_,chained_data_delayed_89__113_,
  chained_data_delayed_89__112_,chained_data_delayed_89__111_,chained_data_delayed_89__110_,
  chained_data_delayed_89__109_,chained_data_delayed_89__108_,
  chained_data_delayed_89__107_,chained_data_delayed_89__106_,chained_data_delayed_89__105_,
  chained_data_delayed_89__104_,chained_data_delayed_89__103_,chained_data_delayed_89__102_,
  chained_data_delayed_89__101_,chained_data_delayed_89__100_,
  chained_data_delayed_89__99_,chained_data_delayed_89__98_,chained_data_delayed_89__97_,
  chained_data_delayed_89__96_,chained_data_delayed_89__95_,chained_data_delayed_89__94_,
  chained_data_delayed_89__93_,chained_data_delayed_89__92_,chained_data_delayed_89__91_,
  chained_data_delayed_89__90_,chained_data_delayed_89__89_,chained_data_delayed_89__88_,
  chained_data_delayed_89__87_,chained_data_delayed_89__86_,
  chained_data_delayed_89__85_,chained_data_delayed_89__84_,chained_data_delayed_89__83_,
  chained_data_delayed_89__82_,chained_data_delayed_89__81_,chained_data_delayed_89__80_,
  chained_data_delayed_89__79_,chained_data_delayed_89__78_,chained_data_delayed_89__77_,
  chained_data_delayed_89__76_,chained_data_delayed_89__75_,
  chained_data_delayed_89__74_,chained_data_delayed_89__73_,chained_data_delayed_89__72_,
  chained_data_delayed_89__71_,chained_data_delayed_89__70_,chained_data_delayed_89__69_,
  chained_data_delayed_89__68_,chained_data_delayed_89__67_,chained_data_delayed_89__66_,
  chained_data_delayed_89__65_,chained_data_delayed_89__64_,
  chained_data_delayed_89__63_,chained_data_delayed_89__62_,chained_data_delayed_89__61_,
  chained_data_delayed_89__60_,chained_data_delayed_89__59_,chained_data_delayed_89__58_,
  chained_data_delayed_89__57_,chained_data_delayed_89__56_,chained_data_delayed_89__55_,
  chained_data_delayed_89__54_,chained_data_delayed_89__53_,
  chained_data_delayed_89__52_,chained_data_delayed_89__51_,chained_data_delayed_89__50_,
  chained_data_delayed_89__49_,chained_data_delayed_89__48_,chained_data_delayed_89__47_,
  chained_data_delayed_89__46_,chained_data_delayed_89__45_,chained_data_delayed_89__44_,
  chained_data_delayed_89__43_,chained_data_delayed_89__42_,
  chained_data_delayed_89__41_,chained_data_delayed_89__40_,chained_data_delayed_89__39_,
  chained_data_delayed_89__38_,chained_data_delayed_89__37_,chained_data_delayed_89__36_,
  chained_data_delayed_89__35_,chained_data_delayed_89__34_,chained_data_delayed_89__33_,
  chained_data_delayed_89__32_,chained_data_delayed_89__31_,
  chained_data_delayed_89__30_,chained_data_delayed_89__29_,chained_data_delayed_89__28_,
  chained_data_delayed_89__27_,chained_data_delayed_89__26_,chained_data_delayed_89__25_,
  chained_data_delayed_89__24_,chained_data_delayed_89__23_,chained_data_delayed_89__22_,
  chained_data_delayed_89__21_,chained_data_delayed_89__20_,
  chained_data_delayed_89__19_,chained_data_delayed_89__18_,chained_data_delayed_89__17_,
  chained_data_delayed_89__16_,chained_data_delayed_89__15_,chained_data_delayed_89__14_,
  chained_data_delayed_89__13_,chained_data_delayed_89__12_,chained_data_delayed_89__11_,
  chained_data_delayed_89__10_,chained_data_delayed_89__9_,chained_data_delayed_89__8_,
  chained_data_delayed_89__7_,chained_data_delayed_89__6_,
  chained_data_delayed_89__5_,chained_data_delayed_89__4_,chained_data_delayed_89__3_,
  chained_data_delayed_89__2_,chained_data_delayed_89__1_,chained_data_delayed_89__0_,
  chained_data_delayed_96__127_,chained_data_delayed_96__126_,chained_data_delayed_96__125_,
  chained_data_delayed_96__124_,chained_data_delayed_96__123_,
  chained_data_delayed_96__122_,chained_data_delayed_96__121_,chained_data_delayed_96__120_,
  chained_data_delayed_96__119_,chained_data_delayed_96__118_,chained_data_delayed_96__117_,
  chained_data_delayed_96__116_,chained_data_delayed_96__115_,
  chained_data_delayed_96__114_,chained_data_delayed_96__113_,chained_data_delayed_96__112_,
  chained_data_delayed_96__111_,chained_data_delayed_96__110_,chained_data_delayed_96__109_,
  chained_data_delayed_96__108_,chained_data_delayed_96__107_,
  chained_data_delayed_96__106_,chained_data_delayed_96__105_,chained_data_delayed_96__104_,
  chained_data_delayed_96__103_,chained_data_delayed_96__102_,chained_data_delayed_96__101_,
  chained_data_delayed_96__100_,chained_data_delayed_96__99_,chained_data_delayed_96__98_,
  chained_data_delayed_96__97_,chained_data_delayed_96__96_,
  chained_data_delayed_96__95_,chained_data_delayed_96__94_,chained_data_delayed_96__93_,
  chained_data_delayed_96__92_,chained_data_delayed_96__91_,chained_data_delayed_96__90_,
  chained_data_delayed_96__89_,chained_data_delayed_96__88_,chained_data_delayed_96__87_,
  chained_data_delayed_96__86_,chained_data_delayed_96__85_,
  chained_data_delayed_96__84_,chained_data_delayed_96__83_,chained_data_delayed_96__82_,
  chained_data_delayed_96__81_,chained_data_delayed_96__80_,chained_data_delayed_96__79_,
  chained_data_delayed_96__78_,chained_data_delayed_96__77_,chained_data_delayed_96__76_,
  chained_data_delayed_96__75_,chained_data_delayed_96__74_,
  chained_data_delayed_96__73_,chained_data_delayed_96__72_,chained_data_delayed_96__71_,
  chained_data_delayed_96__70_,chained_data_delayed_96__69_,chained_data_delayed_96__68_,
  chained_data_delayed_96__67_,chained_data_delayed_96__66_,chained_data_delayed_96__65_,
  chained_data_delayed_96__64_,chained_data_delayed_96__63_,
  chained_data_delayed_96__62_,chained_data_delayed_96__61_,chained_data_delayed_96__60_,
  chained_data_delayed_96__59_,chained_data_delayed_96__58_,chained_data_delayed_96__57_,
  chained_data_delayed_96__56_,chained_data_delayed_96__55_,chained_data_delayed_96__54_,
  chained_data_delayed_96__53_,chained_data_delayed_96__52_,
  chained_data_delayed_96__51_,chained_data_delayed_96__50_,chained_data_delayed_96__49_,
  chained_data_delayed_96__48_,chained_data_delayed_96__47_,chained_data_delayed_96__46_,
  chained_data_delayed_96__45_,chained_data_delayed_96__44_,chained_data_delayed_96__43_,
  chained_data_delayed_96__42_,chained_data_delayed_96__41_,
  chained_data_delayed_96__40_,chained_data_delayed_96__39_,chained_data_delayed_96__38_,
  chained_data_delayed_96__37_,chained_data_delayed_96__36_,chained_data_delayed_96__35_,
  chained_data_delayed_96__34_,chained_data_delayed_96__33_,chained_data_delayed_96__32_,
  chained_data_delayed_96__31_,chained_data_delayed_96__30_,
  chained_data_delayed_96__29_,chained_data_delayed_96__28_,chained_data_delayed_96__27_,
  chained_data_delayed_96__26_,chained_data_delayed_96__25_,chained_data_delayed_96__24_,
  chained_data_delayed_96__23_,chained_data_delayed_96__22_,chained_data_delayed_96__21_,
  chained_data_delayed_96__20_,chained_data_delayed_96__19_,chained_data_delayed_96__18_,
  chained_data_delayed_96__17_,chained_data_delayed_96__16_,
  chained_data_delayed_96__15_,chained_data_delayed_96__14_,chained_data_delayed_96__13_,
  chained_data_delayed_96__12_,chained_data_delayed_96__11_,chained_data_delayed_96__10_,
  chained_data_delayed_96__9_,chained_data_delayed_96__8_,chained_data_delayed_96__7_,
  chained_data_delayed_96__6_,chained_data_delayed_96__5_,chained_data_delayed_96__4_,
  chained_data_delayed_96__3_,chained_data_delayed_96__2_,
  chained_data_delayed_96__1_,chained_data_delayed_96__0_,chained_data_delayed_95__127_,
  chained_data_delayed_95__126_,chained_data_delayed_95__125_,chained_data_delayed_95__124_,
  chained_data_delayed_95__123_,chained_data_delayed_95__122_,
  chained_data_delayed_95__121_,chained_data_delayed_95__120_,chained_data_delayed_95__119_,
  chained_data_delayed_95__118_,chained_data_delayed_95__117_,chained_data_delayed_95__116_,
  chained_data_delayed_95__115_,chained_data_delayed_95__114_,
  chained_data_delayed_95__113_,chained_data_delayed_95__112_,chained_data_delayed_95__111_,
  chained_data_delayed_95__110_,chained_data_delayed_95__109_,chained_data_delayed_95__108_,
  chained_data_delayed_95__107_,chained_data_delayed_95__106_,
  chained_data_delayed_95__105_,chained_data_delayed_95__104_,chained_data_delayed_95__103_,
  chained_data_delayed_95__102_,chained_data_delayed_95__101_,chained_data_delayed_95__100_,
  chained_data_delayed_95__99_,chained_data_delayed_95__98_,chained_data_delayed_95__97_,
  chained_data_delayed_95__96_,chained_data_delayed_95__95_,
  chained_data_delayed_95__94_,chained_data_delayed_95__93_,chained_data_delayed_95__92_,
  chained_data_delayed_95__91_,chained_data_delayed_95__90_,chained_data_delayed_95__89_,
  chained_data_delayed_95__88_,chained_data_delayed_95__87_,chained_data_delayed_95__86_,
  chained_data_delayed_95__85_,chained_data_delayed_95__84_,
  chained_data_delayed_95__83_,chained_data_delayed_95__82_,chained_data_delayed_95__81_,
  chained_data_delayed_95__80_,chained_data_delayed_95__79_,chained_data_delayed_95__78_,
  chained_data_delayed_95__77_,chained_data_delayed_95__76_,chained_data_delayed_95__75_,
  chained_data_delayed_95__74_,chained_data_delayed_95__73_,
  chained_data_delayed_95__72_,chained_data_delayed_95__71_,chained_data_delayed_95__70_,
  chained_data_delayed_95__69_,chained_data_delayed_95__68_,chained_data_delayed_95__67_,
  chained_data_delayed_95__66_,chained_data_delayed_95__65_,chained_data_delayed_95__64_,
  chained_data_delayed_95__63_,chained_data_delayed_95__62_,
  chained_data_delayed_95__61_,chained_data_delayed_95__60_,chained_data_delayed_95__59_,
  chained_data_delayed_95__58_,chained_data_delayed_95__57_,chained_data_delayed_95__56_,
  chained_data_delayed_95__55_,chained_data_delayed_95__54_,chained_data_delayed_95__53_,
  chained_data_delayed_95__52_,chained_data_delayed_95__51_,
  chained_data_delayed_95__50_,chained_data_delayed_95__49_,chained_data_delayed_95__48_,
  chained_data_delayed_95__47_,chained_data_delayed_95__46_,chained_data_delayed_95__45_,
  chained_data_delayed_95__44_,chained_data_delayed_95__43_,chained_data_delayed_95__42_,
  chained_data_delayed_95__41_,chained_data_delayed_95__40_,
  chained_data_delayed_95__39_,chained_data_delayed_95__38_,chained_data_delayed_95__37_,
  chained_data_delayed_95__36_,chained_data_delayed_95__35_,chained_data_delayed_95__34_,
  chained_data_delayed_95__33_,chained_data_delayed_95__32_,chained_data_delayed_95__31_,
  chained_data_delayed_95__30_,chained_data_delayed_95__29_,chained_data_delayed_95__28_,
  chained_data_delayed_95__27_,chained_data_delayed_95__26_,
  chained_data_delayed_95__25_,chained_data_delayed_95__24_,chained_data_delayed_95__23_,
  chained_data_delayed_95__22_,chained_data_delayed_95__21_,chained_data_delayed_95__20_,
  chained_data_delayed_95__19_,chained_data_delayed_95__18_,chained_data_delayed_95__17_,
  chained_data_delayed_95__16_,chained_data_delayed_95__15_,
  chained_data_delayed_95__14_,chained_data_delayed_95__13_,chained_data_delayed_95__12_,
  chained_data_delayed_95__11_,chained_data_delayed_95__10_,chained_data_delayed_95__9_,
  chained_data_delayed_95__8_,chained_data_delayed_95__7_,chained_data_delayed_95__6_,
  chained_data_delayed_95__5_,chained_data_delayed_95__4_,chained_data_delayed_95__3_,
  chained_data_delayed_95__2_,chained_data_delayed_95__1_,
  chained_data_delayed_95__0_,chained_data_delayed_94__127_,chained_data_delayed_94__126_,
  chained_data_delayed_94__125_,chained_data_delayed_94__124_,chained_data_delayed_94__123_,
  chained_data_delayed_94__122_,chained_data_delayed_94__121_,
  chained_data_delayed_94__120_,chained_data_delayed_94__119_,chained_data_delayed_94__118_,
  chained_data_delayed_94__117_,chained_data_delayed_94__116_,chained_data_delayed_94__115_,
  chained_data_delayed_94__114_,chained_data_delayed_94__113_,
  chained_data_delayed_94__112_,chained_data_delayed_94__111_,chained_data_delayed_94__110_,
  chained_data_delayed_94__109_,chained_data_delayed_94__108_,chained_data_delayed_94__107_,
  chained_data_delayed_94__106_,chained_data_delayed_94__105_,
  chained_data_delayed_94__104_,chained_data_delayed_94__103_,chained_data_delayed_94__102_,
  chained_data_delayed_94__101_,chained_data_delayed_94__100_,chained_data_delayed_94__99_,
  chained_data_delayed_94__98_,chained_data_delayed_94__97_,chained_data_delayed_94__96_,
  chained_data_delayed_94__95_,chained_data_delayed_94__94_,
  chained_data_delayed_94__93_,chained_data_delayed_94__92_,chained_data_delayed_94__91_,
  chained_data_delayed_94__90_,chained_data_delayed_94__89_,chained_data_delayed_94__88_,
  chained_data_delayed_94__87_,chained_data_delayed_94__86_,chained_data_delayed_94__85_,
  chained_data_delayed_94__84_,chained_data_delayed_94__83_,
  chained_data_delayed_94__82_,chained_data_delayed_94__81_,chained_data_delayed_94__80_,
  chained_data_delayed_94__79_,chained_data_delayed_94__78_,chained_data_delayed_94__77_,
  chained_data_delayed_94__76_,chained_data_delayed_94__75_,chained_data_delayed_94__74_,
  chained_data_delayed_94__73_,chained_data_delayed_94__72_,
  chained_data_delayed_94__71_,chained_data_delayed_94__70_,chained_data_delayed_94__69_,
  chained_data_delayed_94__68_,chained_data_delayed_94__67_,chained_data_delayed_94__66_,
  chained_data_delayed_94__65_,chained_data_delayed_94__64_,chained_data_delayed_94__63_,
  chained_data_delayed_94__62_,chained_data_delayed_94__61_,
  chained_data_delayed_94__60_,chained_data_delayed_94__59_,chained_data_delayed_94__58_,
  chained_data_delayed_94__57_,chained_data_delayed_94__56_,chained_data_delayed_94__55_,
  chained_data_delayed_94__54_,chained_data_delayed_94__53_,chained_data_delayed_94__52_,
  chained_data_delayed_94__51_,chained_data_delayed_94__50_,
  chained_data_delayed_94__49_,chained_data_delayed_94__48_,chained_data_delayed_94__47_,
  chained_data_delayed_94__46_,chained_data_delayed_94__45_,chained_data_delayed_94__44_,
  chained_data_delayed_94__43_,chained_data_delayed_94__42_,chained_data_delayed_94__41_,
  chained_data_delayed_94__40_,chained_data_delayed_94__39_,chained_data_delayed_94__38_,
  chained_data_delayed_94__37_,chained_data_delayed_94__36_,
  chained_data_delayed_94__35_,chained_data_delayed_94__34_,chained_data_delayed_94__33_,
  chained_data_delayed_94__32_,chained_data_delayed_94__31_,chained_data_delayed_94__30_,
  chained_data_delayed_94__29_,chained_data_delayed_94__28_,chained_data_delayed_94__27_,
  chained_data_delayed_94__26_,chained_data_delayed_94__25_,
  chained_data_delayed_94__24_,chained_data_delayed_94__23_,chained_data_delayed_94__22_,
  chained_data_delayed_94__21_,chained_data_delayed_94__20_,chained_data_delayed_94__19_,
  chained_data_delayed_94__18_,chained_data_delayed_94__17_,chained_data_delayed_94__16_,
  chained_data_delayed_94__15_,chained_data_delayed_94__14_,
  chained_data_delayed_94__13_,chained_data_delayed_94__12_,chained_data_delayed_94__11_,
  chained_data_delayed_94__10_,chained_data_delayed_94__9_,chained_data_delayed_94__8_,
  chained_data_delayed_94__7_,chained_data_delayed_94__6_,chained_data_delayed_94__5_,
  chained_data_delayed_94__4_,chained_data_delayed_94__3_,chained_data_delayed_94__2_,
  chained_data_delayed_94__1_,chained_data_delayed_94__0_,
  chained_data_delayed_93__127_,chained_data_delayed_93__126_,chained_data_delayed_93__125_,
  chained_data_delayed_93__124_,chained_data_delayed_93__123_,chained_data_delayed_93__122_,
  chained_data_delayed_93__121_,chained_data_delayed_93__120_,
  chained_data_delayed_93__119_,chained_data_delayed_93__118_,chained_data_delayed_93__117_,
  chained_data_delayed_93__116_,chained_data_delayed_93__115_,chained_data_delayed_93__114_,
  chained_data_delayed_93__113_,chained_data_delayed_93__112_,
  chained_data_delayed_93__111_,chained_data_delayed_93__110_,chained_data_delayed_93__109_,
  chained_data_delayed_93__108_,chained_data_delayed_93__107_,chained_data_delayed_93__106_,
  chained_data_delayed_93__105_,chained_data_delayed_93__104_,
  chained_data_delayed_93__103_,chained_data_delayed_93__102_,chained_data_delayed_93__101_,
  chained_data_delayed_93__100_,chained_data_delayed_93__99_,chained_data_delayed_93__98_,
  chained_data_delayed_93__97_,chained_data_delayed_93__96_,chained_data_delayed_93__95_,
  chained_data_delayed_93__94_,chained_data_delayed_93__93_,
  chained_data_delayed_93__92_,chained_data_delayed_93__91_,chained_data_delayed_93__90_,
  chained_data_delayed_93__89_,chained_data_delayed_93__88_,chained_data_delayed_93__87_,
  chained_data_delayed_93__86_,chained_data_delayed_93__85_,chained_data_delayed_93__84_,
  chained_data_delayed_93__83_,chained_data_delayed_93__82_,
  chained_data_delayed_93__81_,chained_data_delayed_93__80_,chained_data_delayed_93__79_,
  chained_data_delayed_93__78_,chained_data_delayed_93__77_,chained_data_delayed_93__76_,
  chained_data_delayed_93__75_,chained_data_delayed_93__74_,chained_data_delayed_93__73_,
  chained_data_delayed_93__72_,chained_data_delayed_93__71_,
  chained_data_delayed_93__70_,chained_data_delayed_93__69_,chained_data_delayed_93__68_,
  chained_data_delayed_93__67_,chained_data_delayed_93__66_,chained_data_delayed_93__65_,
  chained_data_delayed_93__64_,chained_data_delayed_93__63_,chained_data_delayed_93__62_,
  chained_data_delayed_93__61_,chained_data_delayed_93__60_,
  chained_data_delayed_93__59_,chained_data_delayed_93__58_,chained_data_delayed_93__57_,
  chained_data_delayed_93__56_,chained_data_delayed_93__55_,chained_data_delayed_93__54_,
  chained_data_delayed_93__53_,chained_data_delayed_93__52_,chained_data_delayed_93__51_,
  chained_data_delayed_93__50_,chained_data_delayed_93__49_,chained_data_delayed_93__48_,
  chained_data_delayed_93__47_,chained_data_delayed_93__46_,
  chained_data_delayed_93__45_,chained_data_delayed_93__44_,chained_data_delayed_93__43_,
  chained_data_delayed_93__42_,chained_data_delayed_93__41_,chained_data_delayed_93__40_,
  chained_data_delayed_93__39_,chained_data_delayed_93__38_,chained_data_delayed_93__37_,
  chained_data_delayed_93__36_,chained_data_delayed_93__35_,
  chained_data_delayed_93__34_,chained_data_delayed_93__33_,chained_data_delayed_93__32_,
  chained_data_delayed_93__31_,chained_data_delayed_93__30_,chained_data_delayed_93__29_,
  chained_data_delayed_93__28_,chained_data_delayed_93__27_,chained_data_delayed_93__26_,
  chained_data_delayed_93__25_,chained_data_delayed_93__24_,
  chained_data_delayed_93__23_,chained_data_delayed_93__22_,chained_data_delayed_93__21_,
  chained_data_delayed_93__20_,chained_data_delayed_93__19_,chained_data_delayed_93__18_,
  chained_data_delayed_93__17_,chained_data_delayed_93__16_,chained_data_delayed_93__15_,
  chained_data_delayed_93__14_,chained_data_delayed_93__13_,
  chained_data_delayed_93__12_,chained_data_delayed_93__11_,chained_data_delayed_93__10_,
  chained_data_delayed_93__9_,chained_data_delayed_93__8_,chained_data_delayed_93__7_,
  chained_data_delayed_93__6_,chained_data_delayed_93__5_,chained_data_delayed_93__4_,
  chained_data_delayed_93__3_,chained_data_delayed_93__2_,chained_data_delayed_93__1_,
  chained_data_delayed_93__0_,chained_data_delayed_100__127_,
  chained_data_delayed_100__126_,chained_data_delayed_100__125_,chained_data_delayed_100__124_,
  chained_data_delayed_100__123_,chained_data_delayed_100__122_,chained_data_delayed_100__121_,
  chained_data_delayed_100__120_,chained_data_delayed_100__119_,
  chained_data_delayed_100__118_,chained_data_delayed_100__117_,chained_data_delayed_100__116_,
  chained_data_delayed_100__115_,chained_data_delayed_100__114_,
  chained_data_delayed_100__113_,chained_data_delayed_100__112_,chained_data_delayed_100__111_,
  chained_data_delayed_100__110_,chained_data_delayed_100__109_,
  chained_data_delayed_100__108_,chained_data_delayed_100__107_,chained_data_delayed_100__106_,
  chained_data_delayed_100__105_,chained_data_delayed_100__104_,chained_data_delayed_100__103_,
  chained_data_delayed_100__102_,chained_data_delayed_100__101_,
  chained_data_delayed_100__100_,chained_data_delayed_100__99_,chained_data_delayed_100__98_,
  chained_data_delayed_100__97_,chained_data_delayed_100__96_,chained_data_delayed_100__95_,
  chained_data_delayed_100__94_,chained_data_delayed_100__93_,
  chained_data_delayed_100__92_,chained_data_delayed_100__91_,chained_data_delayed_100__90_,
  chained_data_delayed_100__89_,chained_data_delayed_100__88_,chained_data_delayed_100__87_,
  chained_data_delayed_100__86_,chained_data_delayed_100__85_,
  chained_data_delayed_100__84_,chained_data_delayed_100__83_,chained_data_delayed_100__82_,
  chained_data_delayed_100__81_,chained_data_delayed_100__80_,chained_data_delayed_100__79_,
  chained_data_delayed_100__78_,chained_data_delayed_100__77_,
  chained_data_delayed_100__76_,chained_data_delayed_100__75_,chained_data_delayed_100__74_,
  chained_data_delayed_100__73_,chained_data_delayed_100__72_,chained_data_delayed_100__71_,
  chained_data_delayed_100__70_,chained_data_delayed_100__69_,
  chained_data_delayed_100__68_,chained_data_delayed_100__67_,chained_data_delayed_100__66_,
  chained_data_delayed_100__65_,chained_data_delayed_100__64_,chained_data_delayed_100__63_,
  chained_data_delayed_100__62_,chained_data_delayed_100__61_,
  chained_data_delayed_100__60_,chained_data_delayed_100__59_,chained_data_delayed_100__58_,
  chained_data_delayed_100__57_,chained_data_delayed_100__56_,chained_data_delayed_100__55_,
  chained_data_delayed_100__54_,chained_data_delayed_100__53_,
  chained_data_delayed_100__52_,chained_data_delayed_100__51_,chained_data_delayed_100__50_,
  chained_data_delayed_100__49_,chained_data_delayed_100__48_,chained_data_delayed_100__47_,
  chained_data_delayed_100__46_,chained_data_delayed_100__45_,
  chained_data_delayed_100__44_,chained_data_delayed_100__43_,chained_data_delayed_100__42_,
  chained_data_delayed_100__41_,chained_data_delayed_100__40_,chained_data_delayed_100__39_,
  chained_data_delayed_100__38_,chained_data_delayed_100__37_,
  chained_data_delayed_100__36_,chained_data_delayed_100__35_,chained_data_delayed_100__34_,
  chained_data_delayed_100__33_,chained_data_delayed_100__32_,chained_data_delayed_100__31_,
  chained_data_delayed_100__30_,chained_data_delayed_100__29_,
  chained_data_delayed_100__28_,chained_data_delayed_100__27_,chained_data_delayed_100__26_,
  chained_data_delayed_100__25_,chained_data_delayed_100__24_,chained_data_delayed_100__23_,
  chained_data_delayed_100__22_,chained_data_delayed_100__21_,
  chained_data_delayed_100__20_,chained_data_delayed_100__19_,chained_data_delayed_100__18_,
  chained_data_delayed_100__17_,chained_data_delayed_100__16_,chained_data_delayed_100__15_,
  chained_data_delayed_100__14_,chained_data_delayed_100__13_,
  chained_data_delayed_100__12_,chained_data_delayed_100__11_,chained_data_delayed_100__10_,
  chained_data_delayed_100__9_,chained_data_delayed_100__8_,chained_data_delayed_100__7_,
  chained_data_delayed_100__6_,chained_data_delayed_100__5_,
  chained_data_delayed_100__4_,chained_data_delayed_100__3_,chained_data_delayed_100__2_,
  chained_data_delayed_100__1_,chained_data_delayed_100__0_,chained_data_delayed_99__127_,
  chained_data_delayed_99__126_,chained_data_delayed_99__125_,chained_data_delayed_99__124_,
  chained_data_delayed_99__123_,chained_data_delayed_99__122_,
  chained_data_delayed_99__121_,chained_data_delayed_99__120_,chained_data_delayed_99__119_,
  chained_data_delayed_99__118_,chained_data_delayed_99__117_,chained_data_delayed_99__116_,
  chained_data_delayed_99__115_,chained_data_delayed_99__114_,
  chained_data_delayed_99__113_,chained_data_delayed_99__112_,chained_data_delayed_99__111_,
  chained_data_delayed_99__110_,chained_data_delayed_99__109_,chained_data_delayed_99__108_,
  chained_data_delayed_99__107_,chained_data_delayed_99__106_,
  chained_data_delayed_99__105_,chained_data_delayed_99__104_,chained_data_delayed_99__103_,
  chained_data_delayed_99__102_,chained_data_delayed_99__101_,chained_data_delayed_99__100_,
  chained_data_delayed_99__99_,chained_data_delayed_99__98_,
  chained_data_delayed_99__97_,chained_data_delayed_99__96_,chained_data_delayed_99__95_,
  chained_data_delayed_99__94_,chained_data_delayed_99__93_,chained_data_delayed_99__92_,
  chained_data_delayed_99__91_,chained_data_delayed_99__90_,chained_data_delayed_99__89_,
  chained_data_delayed_99__88_,chained_data_delayed_99__87_,
  chained_data_delayed_99__86_,chained_data_delayed_99__85_,chained_data_delayed_99__84_,
  chained_data_delayed_99__83_,chained_data_delayed_99__82_,chained_data_delayed_99__81_,
  chained_data_delayed_99__80_,chained_data_delayed_99__79_,chained_data_delayed_99__78_,
  chained_data_delayed_99__77_,chained_data_delayed_99__76_,
  chained_data_delayed_99__75_,chained_data_delayed_99__74_,chained_data_delayed_99__73_,
  chained_data_delayed_99__72_,chained_data_delayed_99__71_,chained_data_delayed_99__70_,
  chained_data_delayed_99__69_,chained_data_delayed_99__68_,chained_data_delayed_99__67_,
  chained_data_delayed_99__66_,chained_data_delayed_99__65_,
  chained_data_delayed_99__64_,chained_data_delayed_99__63_,chained_data_delayed_99__62_,
  chained_data_delayed_99__61_,chained_data_delayed_99__60_,chained_data_delayed_99__59_,
  chained_data_delayed_99__58_,chained_data_delayed_99__57_,chained_data_delayed_99__56_,
  chained_data_delayed_99__55_,chained_data_delayed_99__54_,
  chained_data_delayed_99__53_,chained_data_delayed_99__52_,chained_data_delayed_99__51_,
  chained_data_delayed_99__50_,chained_data_delayed_99__49_,chained_data_delayed_99__48_,
  chained_data_delayed_99__47_,chained_data_delayed_99__46_,chained_data_delayed_99__45_,
  chained_data_delayed_99__44_,chained_data_delayed_99__43_,
  chained_data_delayed_99__42_,chained_data_delayed_99__41_,chained_data_delayed_99__40_,
  chained_data_delayed_99__39_,chained_data_delayed_99__38_,chained_data_delayed_99__37_,
  chained_data_delayed_99__36_,chained_data_delayed_99__35_,chained_data_delayed_99__34_,
  chained_data_delayed_99__33_,chained_data_delayed_99__32_,
  chained_data_delayed_99__31_,chained_data_delayed_99__30_,chained_data_delayed_99__29_,
  chained_data_delayed_99__28_,chained_data_delayed_99__27_,chained_data_delayed_99__26_,
  chained_data_delayed_99__25_,chained_data_delayed_99__24_,chained_data_delayed_99__23_,
  chained_data_delayed_99__22_,chained_data_delayed_99__21_,chained_data_delayed_99__20_,
  chained_data_delayed_99__19_,chained_data_delayed_99__18_,
  chained_data_delayed_99__17_,chained_data_delayed_99__16_,chained_data_delayed_99__15_,
  chained_data_delayed_99__14_,chained_data_delayed_99__13_,chained_data_delayed_99__12_,
  chained_data_delayed_99__11_,chained_data_delayed_99__10_,chained_data_delayed_99__9_,
  chained_data_delayed_99__8_,chained_data_delayed_99__7_,
  chained_data_delayed_99__6_,chained_data_delayed_99__5_,chained_data_delayed_99__4_,
  chained_data_delayed_99__3_,chained_data_delayed_99__2_,chained_data_delayed_99__1_,
  chained_data_delayed_99__0_,chained_data_delayed_98__127_,chained_data_delayed_98__126_,
  chained_data_delayed_98__125_,chained_data_delayed_98__124_,chained_data_delayed_98__123_,
  chained_data_delayed_98__122_,chained_data_delayed_98__121_,
  chained_data_delayed_98__120_,chained_data_delayed_98__119_,chained_data_delayed_98__118_,
  chained_data_delayed_98__117_,chained_data_delayed_98__116_,chained_data_delayed_98__115_,
  chained_data_delayed_98__114_,chained_data_delayed_98__113_,
  chained_data_delayed_98__112_,chained_data_delayed_98__111_,chained_data_delayed_98__110_,
  chained_data_delayed_98__109_,chained_data_delayed_98__108_,chained_data_delayed_98__107_,
  chained_data_delayed_98__106_,chained_data_delayed_98__105_,
  chained_data_delayed_98__104_,chained_data_delayed_98__103_,chained_data_delayed_98__102_,
  chained_data_delayed_98__101_,chained_data_delayed_98__100_,chained_data_delayed_98__99_,
  chained_data_delayed_98__98_,chained_data_delayed_98__97_,
  chained_data_delayed_98__96_,chained_data_delayed_98__95_,chained_data_delayed_98__94_,
  chained_data_delayed_98__93_,chained_data_delayed_98__92_,chained_data_delayed_98__91_,
  chained_data_delayed_98__90_,chained_data_delayed_98__89_,chained_data_delayed_98__88_,
  chained_data_delayed_98__87_,chained_data_delayed_98__86_,
  chained_data_delayed_98__85_,chained_data_delayed_98__84_,chained_data_delayed_98__83_,
  chained_data_delayed_98__82_,chained_data_delayed_98__81_,chained_data_delayed_98__80_,
  chained_data_delayed_98__79_,chained_data_delayed_98__78_,chained_data_delayed_98__77_,
  chained_data_delayed_98__76_,chained_data_delayed_98__75_,
  chained_data_delayed_98__74_,chained_data_delayed_98__73_,chained_data_delayed_98__72_,
  chained_data_delayed_98__71_,chained_data_delayed_98__70_,chained_data_delayed_98__69_,
  chained_data_delayed_98__68_,chained_data_delayed_98__67_,chained_data_delayed_98__66_,
  chained_data_delayed_98__65_,chained_data_delayed_98__64_,
  chained_data_delayed_98__63_,chained_data_delayed_98__62_,chained_data_delayed_98__61_,
  chained_data_delayed_98__60_,chained_data_delayed_98__59_,chained_data_delayed_98__58_,
  chained_data_delayed_98__57_,chained_data_delayed_98__56_,chained_data_delayed_98__55_,
  chained_data_delayed_98__54_,chained_data_delayed_98__53_,
  chained_data_delayed_98__52_,chained_data_delayed_98__51_,chained_data_delayed_98__50_,
  chained_data_delayed_98__49_,chained_data_delayed_98__48_,chained_data_delayed_98__47_,
  chained_data_delayed_98__46_,chained_data_delayed_98__45_,chained_data_delayed_98__44_,
  chained_data_delayed_98__43_,chained_data_delayed_98__42_,
  chained_data_delayed_98__41_,chained_data_delayed_98__40_,chained_data_delayed_98__39_,
  chained_data_delayed_98__38_,chained_data_delayed_98__37_,chained_data_delayed_98__36_,
  chained_data_delayed_98__35_,chained_data_delayed_98__34_,chained_data_delayed_98__33_,
  chained_data_delayed_98__32_,chained_data_delayed_98__31_,chained_data_delayed_98__30_,
  chained_data_delayed_98__29_,chained_data_delayed_98__28_,
  chained_data_delayed_98__27_,chained_data_delayed_98__26_,chained_data_delayed_98__25_,
  chained_data_delayed_98__24_,chained_data_delayed_98__23_,chained_data_delayed_98__22_,
  chained_data_delayed_98__21_,chained_data_delayed_98__20_,chained_data_delayed_98__19_,
  chained_data_delayed_98__18_,chained_data_delayed_98__17_,
  chained_data_delayed_98__16_,chained_data_delayed_98__15_,chained_data_delayed_98__14_,
  chained_data_delayed_98__13_,chained_data_delayed_98__12_,chained_data_delayed_98__11_,
  chained_data_delayed_98__10_,chained_data_delayed_98__9_,chained_data_delayed_98__8_,
  chained_data_delayed_98__7_,chained_data_delayed_98__6_,chained_data_delayed_98__5_,
  chained_data_delayed_98__4_,chained_data_delayed_98__3_,
  chained_data_delayed_98__2_,chained_data_delayed_98__1_,chained_data_delayed_98__0_,
  chained_data_delayed_97__127_,chained_data_delayed_97__126_,chained_data_delayed_97__125_,
  chained_data_delayed_97__124_,chained_data_delayed_97__123_,chained_data_delayed_97__122_,
  chained_data_delayed_97__121_,chained_data_delayed_97__120_,
  chained_data_delayed_97__119_,chained_data_delayed_97__118_,chained_data_delayed_97__117_,
  chained_data_delayed_97__116_,chained_data_delayed_97__115_,chained_data_delayed_97__114_,
  chained_data_delayed_97__113_,chained_data_delayed_97__112_,
  chained_data_delayed_97__111_,chained_data_delayed_97__110_,chained_data_delayed_97__109_,
  chained_data_delayed_97__108_,chained_data_delayed_97__107_,chained_data_delayed_97__106_,
  chained_data_delayed_97__105_,chained_data_delayed_97__104_,
  chained_data_delayed_97__103_,chained_data_delayed_97__102_,chained_data_delayed_97__101_,
  chained_data_delayed_97__100_,chained_data_delayed_97__99_,chained_data_delayed_97__98_,
  chained_data_delayed_97__97_,chained_data_delayed_97__96_,
  chained_data_delayed_97__95_,chained_data_delayed_97__94_,chained_data_delayed_97__93_,
  chained_data_delayed_97__92_,chained_data_delayed_97__91_,chained_data_delayed_97__90_,
  chained_data_delayed_97__89_,chained_data_delayed_97__88_,chained_data_delayed_97__87_,
  chained_data_delayed_97__86_,chained_data_delayed_97__85_,
  chained_data_delayed_97__84_,chained_data_delayed_97__83_,chained_data_delayed_97__82_,
  chained_data_delayed_97__81_,chained_data_delayed_97__80_,chained_data_delayed_97__79_,
  chained_data_delayed_97__78_,chained_data_delayed_97__77_,chained_data_delayed_97__76_,
  chained_data_delayed_97__75_,chained_data_delayed_97__74_,
  chained_data_delayed_97__73_,chained_data_delayed_97__72_,chained_data_delayed_97__71_,
  chained_data_delayed_97__70_,chained_data_delayed_97__69_,chained_data_delayed_97__68_,
  chained_data_delayed_97__67_,chained_data_delayed_97__66_,chained_data_delayed_97__65_,
  chained_data_delayed_97__64_,chained_data_delayed_97__63_,
  chained_data_delayed_97__62_,chained_data_delayed_97__61_,chained_data_delayed_97__60_,
  chained_data_delayed_97__59_,chained_data_delayed_97__58_,chained_data_delayed_97__57_,
  chained_data_delayed_97__56_,chained_data_delayed_97__55_,chained_data_delayed_97__54_,
  chained_data_delayed_97__53_,chained_data_delayed_97__52_,
  chained_data_delayed_97__51_,chained_data_delayed_97__50_,chained_data_delayed_97__49_,
  chained_data_delayed_97__48_,chained_data_delayed_97__47_,chained_data_delayed_97__46_,
  chained_data_delayed_97__45_,chained_data_delayed_97__44_,chained_data_delayed_97__43_,
  chained_data_delayed_97__42_,chained_data_delayed_97__41_,chained_data_delayed_97__40_,
  chained_data_delayed_97__39_,chained_data_delayed_97__38_,
  chained_data_delayed_97__37_,chained_data_delayed_97__36_,chained_data_delayed_97__35_,
  chained_data_delayed_97__34_,chained_data_delayed_97__33_,chained_data_delayed_97__32_,
  chained_data_delayed_97__31_,chained_data_delayed_97__30_,chained_data_delayed_97__29_,
  chained_data_delayed_97__28_,chained_data_delayed_97__27_,
  chained_data_delayed_97__26_,chained_data_delayed_97__25_,chained_data_delayed_97__24_,
  chained_data_delayed_97__23_,chained_data_delayed_97__22_,chained_data_delayed_97__21_,
  chained_data_delayed_97__20_,chained_data_delayed_97__19_,chained_data_delayed_97__18_,
  chained_data_delayed_97__17_,chained_data_delayed_97__16_,
  chained_data_delayed_97__15_,chained_data_delayed_97__14_,chained_data_delayed_97__13_,
  chained_data_delayed_97__12_,chained_data_delayed_97__11_,chained_data_delayed_97__10_,
  chained_data_delayed_97__9_,chained_data_delayed_97__8_,chained_data_delayed_97__7_,
  chained_data_delayed_97__6_,chained_data_delayed_97__5_,chained_data_delayed_97__4_,
  chained_data_delayed_97__3_,chained_data_delayed_97__2_,
  chained_data_delayed_97__1_,chained_data_delayed_97__0_,chained_data_delayed_104__127_,
  chained_data_delayed_104__126_,chained_data_delayed_104__125_,chained_data_delayed_104__124_,
  chained_data_delayed_104__123_,chained_data_delayed_104__122_,
  chained_data_delayed_104__121_,chained_data_delayed_104__120_,chained_data_delayed_104__119_,
  chained_data_delayed_104__118_,chained_data_delayed_104__117_,
  chained_data_delayed_104__116_,chained_data_delayed_104__115_,chained_data_delayed_104__114_,
  chained_data_delayed_104__113_,chained_data_delayed_104__112_,chained_data_delayed_104__111_,
  chained_data_delayed_104__110_,chained_data_delayed_104__109_,
  chained_data_delayed_104__108_,chained_data_delayed_104__107_,chained_data_delayed_104__106_,
  chained_data_delayed_104__105_,chained_data_delayed_104__104_,
  chained_data_delayed_104__103_,chained_data_delayed_104__102_,chained_data_delayed_104__101_,
  chained_data_delayed_104__100_,chained_data_delayed_104__99_,chained_data_delayed_104__98_,
  chained_data_delayed_104__97_,chained_data_delayed_104__96_,
  chained_data_delayed_104__95_,chained_data_delayed_104__94_,chained_data_delayed_104__93_,
  chained_data_delayed_104__92_,chained_data_delayed_104__91_,chained_data_delayed_104__90_,
  chained_data_delayed_104__89_,chained_data_delayed_104__88_,
  chained_data_delayed_104__87_,chained_data_delayed_104__86_,chained_data_delayed_104__85_,
  chained_data_delayed_104__84_,chained_data_delayed_104__83_,chained_data_delayed_104__82_,
  chained_data_delayed_104__81_,chained_data_delayed_104__80_,
  chained_data_delayed_104__79_,chained_data_delayed_104__78_,chained_data_delayed_104__77_,
  chained_data_delayed_104__76_,chained_data_delayed_104__75_,chained_data_delayed_104__74_,
  chained_data_delayed_104__73_,chained_data_delayed_104__72_,
  chained_data_delayed_104__71_,chained_data_delayed_104__70_,chained_data_delayed_104__69_,
  chained_data_delayed_104__68_,chained_data_delayed_104__67_,chained_data_delayed_104__66_,
  chained_data_delayed_104__65_,chained_data_delayed_104__64_,
  chained_data_delayed_104__63_,chained_data_delayed_104__62_,chained_data_delayed_104__61_,
  chained_data_delayed_104__60_,chained_data_delayed_104__59_,chained_data_delayed_104__58_,
  chained_data_delayed_104__57_,chained_data_delayed_104__56_,
  chained_data_delayed_104__55_,chained_data_delayed_104__54_,chained_data_delayed_104__53_,
  chained_data_delayed_104__52_,chained_data_delayed_104__51_,chained_data_delayed_104__50_,
  chained_data_delayed_104__49_,chained_data_delayed_104__48_,
  chained_data_delayed_104__47_,chained_data_delayed_104__46_,chained_data_delayed_104__45_,
  chained_data_delayed_104__44_,chained_data_delayed_104__43_,chained_data_delayed_104__42_,
  chained_data_delayed_104__41_,chained_data_delayed_104__40_,
  chained_data_delayed_104__39_,chained_data_delayed_104__38_,chained_data_delayed_104__37_,
  chained_data_delayed_104__36_,chained_data_delayed_104__35_,chained_data_delayed_104__34_,
  chained_data_delayed_104__33_,chained_data_delayed_104__32_,
  chained_data_delayed_104__31_,chained_data_delayed_104__30_,chained_data_delayed_104__29_,
  chained_data_delayed_104__28_,chained_data_delayed_104__27_,chained_data_delayed_104__26_,
  chained_data_delayed_104__25_,chained_data_delayed_104__24_,
  chained_data_delayed_104__23_,chained_data_delayed_104__22_,chained_data_delayed_104__21_,
  chained_data_delayed_104__20_,chained_data_delayed_104__19_,chained_data_delayed_104__18_,
  chained_data_delayed_104__17_,chained_data_delayed_104__16_,
  chained_data_delayed_104__15_,chained_data_delayed_104__14_,chained_data_delayed_104__13_,
  chained_data_delayed_104__12_,chained_data_delayed_104__11_,chained_data_delayed_104__10_,
  chained_data_delayed_104__9_,chained_data_delayed_104__8_,
  chained_data_delayed_104__7_,chained_data_delayed_104__6_,chained_data_delayed_104__5_,
  chained_data_delayed_104__4_,chained_data_delayed_104__3_,chained_data_delayed_104__2_,
  chained_data_delayed_104__1_,chained_data_delayed_104__0_,chained_data_delayed_103__127_,
  chained_data_delayed_103__126_,chained_data_delayed_103__125_,
  chained_data_delayed_103__124_,chained_data_delayed_103__123_,chained_data_delayed_103__122_,
  chained_data_delayed_103__121_,chained_data_delayed_103__120_,
  chained_data_delayed_103__119_,chained_data_delayed_103__118_,chained_data_delayed_103__117_,
  chained_data_delayed_103__116_,chained_data_delayed_103__115_,
  chained_data_delayed_103__114_,chained_data_delayed_103__113_,chained_data_delayed_103__112_,
  chained_data_delayed_103__111_,chained_data_delayed_103__110_,chained_data_delayed_103__109_,
  chained_data_delayed_103__108_,chained_data_delayed_103__107_,
  chained_data_delayed_103__106_,chained_data_delayed_103__105_,chained_data_delayed_103__104_,
  chained_data_delayed_103__103_,chained_data_delayed_103__102_,
  chained_data_delayed_103__101_,chained_data_delayed_103__100_,chained_data_delayed_103__99_,
  chained_data_delayed_103__98_,chained_data_delayed_103__97_,chained_data_delayed_103__96_,
  chained_data_delayed_103__95_,chained_data_delayed_103__94_,
  chained_data_delayed_103__93_,chained_data_delayed_103__92_,chained_data_delayed_103__91_,
  chained_data_delayed_103__90_,chained_data_delayed_103__89_,chained_data_delayed_103__88_,
  chained_data_delayed_103__87_,chained_data_delayed_103__86_,
  chained_data_delayed_103__85_,chained_data_delayed_103__84_,chained_data_delayed_103__83_,
  chained_data_delayed_103__82_,chained_data_delayed_103__81_,chained_data_delayed_103__80_,
  chained_data_delayed_103__79_,chained_data_delayed_103__78_,
  chained_data_delayed_103__77_,chained_data_delayed_103__76_,chained_data_delayed_103__75_,
  chained_data_delayed_103__74_,chained_data_delayed_103__73_,chained_data_delayed_103__72_,
  chained_data_delayed_103__71_,chained_data_delayed_103__70_,
  chained_data_delayed_103__69_,chained_data_delayed_103__68_,chained_data_delayed_103__67_,
  chained_data_delayed_103__66_,chained_data_delayed_103__65_,chained_data_delayed_103__64_,
  chained_data_delayed_103__63_,chained_data_delayed_103__62_,
  chained_data_delayed_103__61_,chained_data_delayed_103__60_,chained_data_delayed_103__59_,
  chained_data_delayed_103__58_,chained_data_delayed_103__57_,chained_data_delayed_103__56_,
  chained_data_delayed_103__55_,chained_data_delayed_103__54_,
  chained_data_delayed_103__53_,chained_data_delayed_103__52_,chained_data_delayed_103__51_,
  chained_data_delayed_103__50_,chained_data_delayed_103__49_,chained_data_delayed_103__48_,
  chained_data_delayed_103__47_,chained_data_delayed_103__46_,
  chained_data_delayed_103__45_,chained_data_delayed_103__44_,chained_data_delayed_103__43_,
  chained_data_delayed_103__42_,chained_data_delayed_103__41_,chained_data_delayed_103__40_,
  chained_data_delayed_103__39_,chained_data_delayed_103__38_,
  chained_data_delayed_103__37_,chained_data_delayed_103__36_,chained_data_delayed_103__35_,
  chained_data_delayed_103__34_,chained_data_delayed_103__33_,chained_data_delayed_103__32_,
  chained_data_delayed_103__31_,chained_data_delayed_103__30_,
  chained_data_delayed_103__29_,chained_data_delayed_103__28_,chained_data_delayed_103__27_,
  chained_data_delayed_103__26_,chained_data_delayed_103__25_,chained_data_delayed_103__24_,
  chained_data_delayed_103__23_,chained_data_delayed_103__22_,
  chained_data_delayed_103__21_,chained_data_delayed_103__20_,chained_data_delayed_103__19_,
  chained_data_delayed_103__18_,chained_data_delayed_103__17_,chained_data_delayed_103__16_,
  chained_data_delayed_103__15_,chained_data_delayed_103__14_,
  chained_data_delayed_103__13_,chained_data_delayed_103__12_,chained_data_delayed_103__11_,
  chained_data_delayed_103__10_,chained_data_delayed_103__9_,chained_data_delayed_103__8_,
  chained_data_delayed_103__7_,chained_data_delayed_103__6_,
  chained_data_delayed_103__5_,chained_data_delayed_103__4_,chained_data_delayed_103__3_,
  chained_data_delayed_103__2_,chained_data_delayed_103__1_,chained_data_delayed_103__0_,
  chained_data_delayed_102__127_,chained_data_delayed_102__126_,chained_data_delayed_102__125_,
  chained_data_delayed_102__124_,chained_data_delayed_102__123_,
  chained_data_delayed_102__122_,chained_data_delayed_102__121_,chained_data_delayed_102__120_,
  chained_data_delayed_102__119_,chained_data_delayed_102__118_,
  chained_data_delayed_102__117_,chained_data_delayed_102__116_,chained_data_delayed_102__115_,
  chained_data_delayed_102__114_,chained_data_delayed_102__113_,
  chained_data_delayed_102__112_,chained_data_delayed_102__111_,chained_data_delayed_102__110_,
  chained_data_delayed_102__109_,chained_data_delayed_102__108_,chained_data_delayed_102__107_,
  chained_data_delayed_102__106_,chained_data_delayed_102__105_,
  chained_data_delayed_102__104_,chained_data_delayed_102__103_,chained_data_delayed_102__102_,
  chained_data_delayed_102__101_,chained_data_delayed_102__100_,
  chained_data_delayed_102__99_,chained_data_delayed_102__98_,chained_data_delayed_102__97_,
  chained_data_delayed_102__96_,chained_data_delayed_102__95_,chained_data_delayed_102__94_,
  chained_data_delayed_102__93_,chained_data_delayed_102__92_,
  chained_data_delayed_102__91_,chained_data_delayed_102__90_,chained_data_delayed_102__89_,
  chained_data_delayed_102__88_,chained_data_delayed_102__87_,chained_data_delayed_102__86_,
  chained_data_delayed_102__85_,chained_data_delayed_102__84_,
  chained_data_delayed_102__83_,chained_data_delayed_102__82_,chained_data_delayed_102__81_,
  chained_data_delayed_102__80_,chained_data_delayed_102__79_,chained_data_delayed_102__78_,
  chained_data_delayed_102__77_,chained_data_delayed_102__76_,
  chained_data_delayed_102__75_,chained_data_delayed_102__74_,chained_data_delayed_102__73_,
  chained_data_delayed_102__72_,chained_data_delayed_102__71_,chained_data_delayed_102__70_,
  chained_data_delayed_102__69_,chained_data_delayed_102__68_,
  chained_data_delayed_102__67_,chained_data_delayed_102__66_,chained_data_delayed_102__65_,
  chained_data_delayed_102__64_,chained_data_delayed_102__63_,chained_data_delayed_102__62_,
  chained_data_delayed_102__61_,chained_data_delayed_102__60_,
  chained_data_delayed_102__59_,chained_data_delayed_102__58_,chained_data_delayed_102__57_,
  chained_data_delayed_102__56_,chained_data_delayed_102__55_,chained_data_delayed_102__54_,
  chained_data_delayed_102__53_,chained_data_delayed_102__52_,
  chained_data_delayed_102__51_,chained_data_delayed_102__50_,chained_data_delayed_102__49_,
  chained_data_delayed_102__48_,chained_data_delayed_102__47_,chained_data_delayed_102__46_,
  chained_data_delayed_102__45_,chained_data_delayed_102__44_,
  chained_data_delayed_102__43_,chained_data_delayed_102__42_,chained_data_delayed_102__41_,
  chained_data_delayed_102__40_,chained_data_delayed_102__39_,chained_data_delayed_102__38_,
  chained_data_delayed_102__37_,chained_data_delayed_102__36_,
  chained_data_delayed_102__35_,chained_data_delayed_102__34_,chained_data_delayed_102__33_,
  chained_data_delayed_102__32_,chained_data_delayed_102__31_,chained_data_delayed_102__30_,
  chained_data_delayed_102__29_,chained_data_delayed_102__28_,
  chained_data_delayed_102__27_,chained_data_delayed_102__26_,chained_data_delayed_102__25_,
  chained_data_delayed_102__24_,chained_data_delayed_102__23_,chained_data_delayed_102__22_,
  chained_data_delayed_102__21_,chained_data_delayed_102__20_,
  chained_data_delayed_102__19_,chained_data_delayed_102__18_,chained_data_delayed_102__17_,
  chained_data_delayed_102__16_,chained_data_delayed_102__15_,chained_data_delayed_102__14_,
  chained_data_delayed_102__13_,chained_data_delayed_102__12_,
  chained_data_delayed_102__11_,chained_data_delayed_102__10_,chained_data_delayed_102__9_,
  chained_data_delayed_102__8_,chained_data_delayed_102__7_,chained_data_delayed_102__6_,
  chained_data_delayed_102__5_,chained_data_delayed_102__4_,chained_data_delayed_102__3_,
  chained_data_delayed_102__2_,chained_data_delayed_102__1_,
  chained_data_delayed_102__0_,chained_data_delayed_101__127_,chained_data_delayed_101__126_,
  chained_data_delayed_101__125_,chained_data_delayed_101__124_,chained_data_delayed_101__123_,
  chained_data_delayed_101__122_,chained_data_delayed_101__121_,
  chained_data_delayed_101__120_,chained_data_delayed_101__119_,chained_data_delayed_101__118_,
  chained_data_delayed_101__117_,chained_data_delayed_101__116_,
  chained_data_delayed_101__115_,chained_data_delayed_101__114_,chained_data_delayed_101__113_,
  chained_data_delayed_101__112_,chained_data_delayed_101__111_,
  chained_data_delayed_101__110_,chained_data_delayed_101__109_,chained_data_delayed_101__108_,
  chained_data_delayed_101__107_,chained_data_delayed_101__106_,chained_data_delayed_101__105_,
  chained_data_delayed_101__104_,chained_data_delayed_101__103_,
  chained_data_delayed_101__102_,chained_data_delayed_101__101_,chained_data_delayed_101__100_,
  chained_data_delayed_101__99_,chained_data_delayed_101__98_,
  chained_data_delayed_101__97_,chained_data_delayed_101__96_,chained_data_delayed_101__95_,
  chained_data_delayed_101__94_,chained_data_delayed_101__93_,chained_data_delayed_101__92_,
  chained_data_delayed_101__91_,chained_data_delayed_101__90_,
  chained_data_delayed_101__89_,chained_data_delayed_101__88_,chained_data_delayed_101__87_,
  chained_data_delayed_101__86_,chained_data_delayed_101__85_,chained_data_delayed_101__84_,
  chained_data_delayed_101__83_,chained_data_delayed_101__82_,
  chained_data_delayed_101__81_,chained_data_delayed_101__80_,chained_data_delayed_101__79_,
  chained_data_delayed_101__78_,chained_data_delayed_101__77_,chained_data_delayed_101__76_,
  chained_data_delayed_101__75_,chained_data_delayed_101__74_,
  chained_data_delayed_101__73_,chained_data_delayed_101__72_,chained_data_delayed_101__71_,
  chained_data_delayed_101__70_,chained_data_delayed_101__69_,chained_data_delayed_101__68_,
  chained_data_delayed_101__67_,chained_data_delayed_101__66_,
  chained_data_delayed_101__65_,chained_data_delayed_101__64_,chained_data_delayed_101__63_,
  chained_data_delayed_101__62_,chained_data_delayed_101__61_,chained_data_delayed_101__60_,
  chained_data_delayed_101__59_,chained_data_delayed_101__58_,
  chained_data_delayed_101__57_,chained_data_delayed_101__56_,chained_data_delayed_101__55_,
  chained_data_delayed_101__54_,chained_data_delayed_101__53_,chained_data_delayed_101__52_,
  chained_data_delayed_101__51_,chained_data_delayed_101__50_,
  chained_data_delayed_101__49_,chained_data_delayed_101__48_,chained_data_delayed_101__47_,
  chained_data_delayed_101__46_,chained_data_delayed_101__45_,chained_data_delayed_101__44_,
  chained_data_delayed_101__43_,chained_data_delayed_101__42_,
  chained_data_delayed_101__41_,chained_data_delayed_101__40_,chained_data_delayed_101__39_,
  chained_data_delayed_101__38_,chained_data_delayed_101__37_,chained_data_delayed_101__36_,
  chained_data_delayed_101__35_,chained_data_delayed_101__34_,
  chained_data_delayed_101__33_,chained_data_delayed_101__32_,chained_data_delayed_101__31_,
  chained_data_delayed_101__30_,chained_data_delayed_101__29_,chained_data_delayed_101__28_,
  chained_data_delayed_101__27_,chained_data_delayed_101__26_,
  chained_data_delayed_101__25_,chained_data_delayed_101__24_,chained_data_delayed_101__23_,
  chained_data_delayed_101__22_,chained_data_delayed_101__21_,chained_data_delayed_101__20_,
  chained_data_delayed_101__19_,chained_data_delayed_101__18_,
  chained_data_delayed_101__17_,chained_data_delayed_101__16_,chained_data_delayed_101__15_,
  chained_data_delayed_101__14_,chained_data_delayed_101__13_,chained_data_delayed_101__12_,
  chained_data_delayed_101__11_,chained_data_delayed_101__10_,
  chained_data_delayed_101__9_,chained_data_delayed_101__8_,chained_data_delayed_101__7_,
  chained_data_delayed_101__6_,chained_data_delayed_101__5_,chained_data_delayed_101__4_,
  chained_data_delayed_101__3_,chained_data_delayed_101__2_,chained_data_delayed_101__1_,
  chained_data_delayed_101__0_,chained_data_delayed_108__127_,
  chained_data_delayed_108__126_,chained_data_delayed_108__125_,chained_data_delayed_108__124_,
  chained_data_delayed_108__123_,chained_data_delayed_108__122_,chained_data_delayed_108__121_,
  chained_data_delayed_108__120_,chained_data_delayed_108__119_,
  chained_data_delayed_108__118_,chained_data_delayed_108__117_,chained_data_delayed_108__116_,
  chained_data_delayed_108__115_,chained_data_delayed_108__114_,
  chained_data_delayed_108__113_,chained_data_delayed_108__112_,chained_data_delayed_108__111_,
  chained_data_delayed_108__110_,chained_data_delayed_108__109_,
  chained_data_delayed_108__108_,chained_data_delayed_108__107_,chained_data_delayed_108__106_,
  chained_data_delayed_108__105_,chained_data_delayed_108__104_,chained_data_delayed_108__103_,
  chained_data_delayed_108__102_,chained_data_delayed_108__101_,
  chained_data_delayed_108__100_,chained_data_delayed_108__99_,chained_data_delayed_108__98_,
  chained_data_delayed_108__97_,chained_data_delayed_108__96_,chained_data_delayed_108__95_,
  chained_data_delayed_108__94_,chained_data_delayed_108__93_,
  chained_data_delayed_108__92_,chained_data_delayed_108__91_,chained_data_delayed_108__90_,
  chained_data_delayed_108__89_,chained_data_delayed_108__88_,chained_data_delayed_108__87_,
  chained_data_delayed_108__86_,chained_data_delayed_108__85_,
  chained_data_delayed_108__84_,chained_data_delayed_108__83_,chained_data_delayed_108__82_,
  chained_data_delayed_108__81_,chained_data_delayed_108__80_,chained_data_delayed_108__79_,
  chained_data_delayed_108__78_,chained_data_delayed_108__77_,
  chained_data_delayed_108__76_,chained_data_delayed_108__75_,chained_data_delayed_108__74_,
  chained_data_delayed_108__73_,chained_data_delayed_108__72_,chained_data_delayed_108__71_,
  chained_data_delayed_108__70_,chained_data_delayed_108__69_,
  chained_data_delayed_108__68_,chained_data_delayed_108__67_,chained_data_delayed_108__66_,
  chained_data_delayed_108__65_,chained_data_delayed_108__64_,chained_data_delayed_108__63_,
  chained_data_delayed_108__62_,chained_data_delayed_108__61_,
  chained_data_delayed_108__60_,chained_data_delayed_108__59_,chained_data_delayed_108__58_,
  chained_data_delayed_108__57_,chained_data_delayed_108__56_,chained_data_delayed_108__55_,
  chained_data_delayed_108__54_,chained_data_delayed_108__53_,
  chained_data_delayed_108__52_,chained_data_delayed_108__51_,chained_data_delayed_108__50_,
  chained_data_delayed_108__49_,chained_data_delayed_108__48_,chained_data_delayed_108__47_,
  chained_data_delayed_108__46_,chained_data_delayed_108__45_,
  chained_data_delayed_108__44_,chained_data_delayed_108__43_,chained_data_delayed_108__42_,
  chained_data_delayed_108__41_,chained_data_delayed_108__40_,chained_data_delayed_108__39_,
  chained_data_delayed_108__38_,chained_data_delayed_108__37_,
  chained_data_delayed_108__36_,chained_data_delayed_108__35_,chained_data_delayed_108__34_,
  chained_data_delayed_108__33_,chained_data_delayed_108__32_,chained_data_delayed_108__31_,
  chained_data_delayed_108__30_,chained_data_delayed_108__29_,
  chained_data_delayed_108__28_,chained_data_delayed_108__27_,chained_data_delayed_108__26_,
  chained_data_delayed_108__25_,chained_data_delayed_108__24_,chained_data_delayed_108__23_,
  chained_data_delayed_108__22_,chained_data_delayed_108__21_,
  chained_data_delayed_108__20_,chained_data_delayed_108__19_,chained_data_delayed_108__18_,
  chained_data_delayed_108__17_,chained_data_delayed_108__16_,chained_data_delayed_108__15_,
  chained_data_delayed_108__14_,chained_data_delayed_108__13_,
  chained_data_delayed_108__12_,chained_data_delayed_108__11_,chained_data_delayed_108__10_,
  chained_data_delayed_108__9_,chained_data_delayed_108__8_,chained_data_delayed_108__7_,
  chained_data_delayed_108__6_,chained_data_delayed_108__5_,
  chained_data_delayed_108__4_,chained_data_delayed_108__3_,chained_data_delayed_108__2_,
  chained_data_delayed_108__1_,chained_data_delayed_108__0_,chained_data_delayed_107__127_,
  chained_data_delayed_107__126_,chained_data_delayed_107__125_,
  chained_data_delayed_107__124_,chained_data_delayed_107__123_,chained_data_delayed_107__122_,
  chained_data_delayed_107__121_,chained_data_delayed_107__120_,chained_data_delayed_107__119_,
  chained_data_delayed_107__118_,chained_data_delayed_107__117_,
  chained_data_delayed_107__116_,chained_data_delayed_107__115_,chained_data_delayed_107__114_,
  chained_data_delayed_107__113_,chained_data_delayed_107__112_,
  chained_data_delayed_107__111_,chained_data_delayed_107__110_,chained_data_delayed_107__109_,
  chained_data_delayed_107__108_,chained_data_delayed_107__107_,
  chained_data_delayed_107__106_,chained_data_delayed_107__105_,chained_data_delayed_107__104_,
  chained_data_delayed_107__103_,chained_data_delayed_107__102_,chained_data_delayed_107__101_,
  chained_data_delayed_107__100_,chained_data_delayed_107__99_,
  chained_data_delayed_107__98_,chained_data_delayed_107__97_,chained_data_delayed_107__96_,
  chained_data_delayed_107__95_,chained_data_delayed_107__94_,chained_data_delayed_107__93_,
  chained_data_delayed_107__92_,chained_data_delayed_107__91_,
  chained_data_delayed_107__90_,chained_data_delayed_107__89_,chained_data_delayed_107__88_,
  chained_data_delayed_107__87_,chained_data_delayed_107__86_,chained_data_delayed_107__85_,
  chained_data_delayed_107__84_,chained_data_delayed_107__83_,
  chained_data_delayed_107__82_,chained_data_delayed_107__81_,chained_data_delayed_107__80_,
  chained_data_delayed_107__79_,chained_data_delayed_107__78_,chained_data_delayed_107__77_,
  chained_data_delayed_107__76_,chained_data_delayed_107__75_,
  chained_data_delayed_107__74_,chained_data_delayed_107__73_,chained_data_delayed_107__72_,
  chained_data_delayed_107__71_,chained_data_delayed_107__70_,chained_data_delayed_107__69_,
  chained_data_delayed_107__68_,chained_data_delayed_107__67_,
  chained_data_delayed_107__66_,chained_data_delayed_107__65_,chained_data_delayed_107__64_,
  chained_data_delayed_107__63_,chained_data_delayed_107__62_,chained_data_delayed_107__61_,
  chained_data_delayed_107__60_,chained_data_delayed_107__59_,
  chained_data_delayed_107__58_,chained_data_delayed_107__57_,chained_data_delayed_107__56_,
  chained_data_delayed_107__55_,chained_data_delayed_107__54_,chained_data_delayed_107__53_,
  chained_data_delayed_107__52_,chained_data_delayed_107__51_,
  chained_data_delayed_107__50_,chained_data_delayed_107__49_,chained_data_delayed_107__48_,
  chained_data_delayed_107__47_,chained_data_delayed_107__46_,chained_data_delayed_107__45_,
  chained_data_delayed_107__44_,chained_data_delayed_107__43_,
  chained_data_delayed_107__42_,chained_data_delayed_107__41_,chained_data_delayed_107__40_,
  chained_data_delayed_107__39_,chained_data_delayed_107__38_,chained_data_delayed_107__37_,
  chained_data_delayed_107__36_,chained_data_delayed_107__35_,
  chained_data_delayed_107__34_,chained_data_delayed_107__33_,chained_data_delayed_107__32_,
  chained_data_delayed_107__31_,chained_data_delayed_107__30_,chained_data_delayed_107__29_,
  chained_data_delayed_107__28_,chained_data_delayed_107__27_,
  chained_data_delayed_107__26_,chained_data_delayed_107__25_,chained_data_delayed_107__24_,
  chained_data_delayed_107__23_,chained_data_delayed_107__22_,chained_data_delayed_107__21_,
  chained_data_delayed_107__20_,chained_data_delayed_107__19_,
  chained_data_delayed_107__18_,chained_data_delayed_107__17_,chained_data_delayed_107__16_,
  chained_data_delayed_107__15_,chained_data_delayed_107__14_,chained_data_delayed_107__13_,
  chained_data_delayed_107__12_,chained_data_delayed_107__11_,
  chained_data_delayed_107__10_,chained_data_delayed_107__9_,chained_data_delayed_107__8_,
  chained_data_delayed_107__7_,chained_data_delayed_107__6_,chained_data_delayed_107__5_,
  chained_data_delayed_107__4_,chained_data_delayed_107__3_,chained_data_delayed_107__2_,
  chained_data_delayed_107__1_,chained_data_delayed_107__0_,
  chained_data_delayed_106__127_,chained_data_delayed_106__126_,chained_data_delayed_106__125_,
  chained_data_delayed_106__124_,chained_data_delayed_106__123_,
  chained_data_delayed_106__122_,chained_data_delayed_106__121_,chained_data_delayed_106__120_,
  chained_data_delayed_106__119_,chained_data_delayed_106__118_,chained_data_delayed_106__117_,
  chained_data_delayed_106__116_,chained_data_delayed_106__115_,
  chained_data_delayed_106__114_,chained_data_delayed_106__113_,chained_data_delayed_106__112_,
  chained_data_delayed_106__111_,chained_data_delayed_106__110_,
  chained_data_delayed_106__109_,chained_data_delayed_106__108_,chained_data_delayed_106__107_,
  chained_data_delayed_106__106_,chained_data_delayed_106__105_,
  chained_data_delayed_106__104_,chained_data_delayed_106__103_,chained_data_delayed_106__102_,
  chained_data_delayed_106__101_,chained_data_delayed_106__100_,chained_data_delayed_106__99_,
  chained_data_delayed_106__98_,chained_data_delayed_106__97_,
  chained_data_delayed_106__96_,chained_data_delayed_106__95_,chained_data_delayed_106__94_,
  chained_data_delayed_106__93_,chained_data_delayed_106__92_,chained_data_delayed_106__91_,
  chained_data_delayed_106__90_,chained_data_delayed_106__89_,
  chained_data_delayed_106__88_,chained_data_delayed_106__87_,chained_data_delayed_106__86_,
  chained_data_delayed_106__85_,chained_data_delayed_106__84_,chained_data_delayed_106__83_,
  chained_data_delayed_106__82_,chained_data_delayed_106__81_,
  chained_data_delayed_106__80_,chained_data_delayed_106__79_,chained_data_delayed_106__78_,
  chained_data_delayed_106__77_,chained_data_delayed_106__76_,chained_data_delayed_106__75_,
  chained_data_delayed_106__74_,chained_data_delayed_106__73_,
  chained_data_delayed_106__72_,chained_data_delayed_106__71_,chained_data_delayed_106__70_,
  chained_data_delayed_106__69_,chained_data_delayed_106__68_,chained_data_delayed_106__67_,
  chained_data_delayed_106__66_,chained_data_delayed_106__65_,
  chained_data_delayed_106__64_,chained_data_delayed_106__63_,chained_data_delayed_106__62_,
  chained_data_delayed_106__61_,chained_data_delayed_106__60_,chained_data_delayed_106__59_,
  chained_data_delayed_106__58_,chained_data_delayed_106__57_,
  chained_data_delayed_106__56_,chained_data_delayed_106__55_,chained_data_delayed_106__54_,
  chained_data_delayed_106__53_,chained_data_delayed_106__52_,chained_data_delayed_106__51_,
  chained_data_delayed_106__50_,chained_data_delayed_106__49_,
  chained_data_delayed_106__48_,chained_data_delayed_106__47_,chained_data_delayed_106__46_,
  chained_data_delayed_106__45_,chained_data_delayed_106__44_,chained_data_delayed_106__43_,
  chained_data_delayed_106__42_,chained_data_delayed_106__41_,
  chained_data_delayed_106__40_,chained_data_delayed_106__39_,chained_data_delayed_106__38_,
  chained_data_delayed_106__37_,chained_data_delayed_106__36_,chained_data_delayed_106__35_,
  chained_data_delayed_106__34_,chained_data_delayed_106__33_,
  chained_data_delayed_106__32_,chained_data_delayed_106__31_,chained_data_delayed_106__30_,
  chained_data_delayed_106__29_,chained_data_delayed_106__28_,chained_data_delayed_106__27_,
  chained_data_delayed_106__26_,chained_data_delayed_106__25_,
  chained_data_delayed_106__24_,chained_data_delayed_106__23_,chained_data_delayed_106__22_,
  chained_data_delayed_106__21_,chained_data_delayed_106__20_,chained_data_delayed_106__19_,
  chained_data_delayed_106__18_,chained_data_delayed_106__17_,
  chained_data_delayed_106__16_,chained_data_delayed_106__15_,chained_data_delayed_106__14_,
  chained_data_delayed_106__13_,chained_data_delayed_106__12_,chained_data_delayed_106__11_,
  chained_data_delayed_106__10_,chained_data_delayed_106__9_,
  chained_data_delayed_106__8_,chained_data_delayed_106__7_,chained_data_delayed_106__6_,
  chained_data_delayed_106__5_,chained_data_delayed_106__4_,chained_data_delayed_106__3_,
  chained_data_delayed_106__2_,chained_data_delayed_106__1_,chained_data_delayed_106__0_,
  chained_data_delayed_105__127_,chained_data_delayed_105__126_,
  chained_data_delayed_105__125_,chained_data_delayed_105__124_,chained_data_delayed_105__123_,
  chained_data_delayed_105__122_,chained_data_delayed_105__121_,
  chained_data_delayed_105__120_,chained_data_delayed_105__119_,chained_data_delayed_105__118_,
  chained_data_delayed_105__117_,chained_data_delayed_105__116_,chained_data_delayed_105__115_,
  chained_data_delayed_105__114_,chained_data_delayed_105__113_,
  chained_data_delayed_105__112_,chained_data_delayed_105__111_,chained_data_delayed_105__110_,
  chained_data_delayed_105__109_,chained_data_delayed_105__108_,
  chained_data_delayed_105__107_,chained_data_delayed_105__106_,chained_data_delayed_105__105_,
  chained_data_delayed_105__104_,chained_data_delayed_105__103_,
  chained_data_delayed_105__102_,chained_data_delayed_105__101_,chained_data_delayed_105__100_,
  chained_data_delayed_105__99_,chained_data_delayed_105__98_,chained_data_delayed_105__97_,
  chained_data_delayed_105__96_,chained_data_delayed_105__95_,
  chained_data_delayed_105__94_,chained_data_delayed_105__93_,chained_data_delayed_105__92_,
  chained_data_delayed_105__91_,chained_data_delayed_105__90_,chained_data_delayed_105__89_,
  chained_data_delayed_105__88_,chained_data_delayed_105__87_,
  chained_data_delayed_105__86_,chained_data_delayed_105__85_,chained_data_delayed_105__84_,
  chained_data_delayed_105__83_,chained_data_delayed_105__82_,chained_data_delayed_105__81_,
  chained_data_delayed_105__80_,chained_data_delayed_105__79_,
  chained_data_delayed_105__78_,chained_data_delayed_105__77_,chained_data_delayed_105__76_,
  chained_data_delayed_105__75_,chained_data_delayed_105__74_,chained_data_delayed_105__73_,
  chained_data_delayed_105__72_,chained_data_delayed_105__71_,
  chained_data_delayed_105__70_,chained_data_delayed_105__69_,chained_data_delayed_105__68_,
  chained_data_delayed_105__67_,chained_data_delayed_105__66_,chained_data_delayed_105__65_,
  chained_data_delayed_105__64_,chained_data_delayed_105__63_,
  chained_data_delayed_105__62_,chained_data_delayed_105__61_,chained_data_delayed_105__60_,
  chained_data_delayed_105__59_,chained_data_delayed_105__58_,chained_data_delayed_105__57_,
  chained_data_delayed_105__56_,chained_data_delayed_105__55_,
  chained_data_delayed_105__54_,chained_data_delayed_105__53_,chained_data_delayed_105__52_,
  chained_data_delayed_105__51_,chained_data_delayed_105__50_,chained_data_delayed_105__49_,
  chained_data_delayed_105__48_,chained_data_delayed_105__47_,
  chained_data_delayed_105__46_,chained_data_delayed_105__45_,chained_data_delayed_105__44_,
  chained_data_delayed_105__43_,chained_data_delayed_105__42_,chained_data_delayed_105__41_,
  chained_data_delayed_105__40_,chained_data_delayed_105__39_,
  chained_data_delayed_105__38_,chained_data_delayed_105__37_,chained_data_delayed_105__36_,
  chained_data_delayed_105__35_,chained_data_delayed_105__34_,chained_data_delayed_105__33_,
  chained_data_delayed_105__32_,chained_data_delayed_105__31_,
  chained_data_delayed_105__30_,chained_data_delayed_105__29_,chained_data_delayed_105__28_,
  chained_data_delayed_105__27_,chained_data_delayed_105__26_,chained_data_delayed_105__25_,
  chained_data_delayed_105__24_,chained_data_delayed_105__23_,
  chained_data_delayed_105__22_,chained_data_delayed_105__21_,chained_data_delayed_105__20_,
  chained_data_delayed_105__19_,chained_data_delayed_105__18_,chained_data_delayed_105__17_,
  chained_data_delayed_105__16_,chained_data_delayed_105__15_,
  chained_data_delayed_105__14_,chained_data_delayed_105__13_,chained_data_delayed_105__12_,
  chained_data_delayed_105__11_,chained_data_delayed_105__10_,chained_data_delayed_105__9_,
  chained_data_delayed_105__8_,chained_data_delayed_105__7_,chained_data_delayed_105__6_,
  chained_data_delayed_105__5_,chained_data_delayed_105__4_,
  chained_data_delayed_105__3_,chained_data_delayed_105__2_,chained_data_delayed_105__1_,
  chained_data_delayed_105__0_,chained_data_delayed_112__127_,chained_data_delayed_112__126_,
  chained_data_delayed_112__125_,chained_data_delayed_112__124_,
  chained_data_delayed_112__123_,chained_data_delayed_112__122_,chained_data_delayed_112__121_,
  chained_data_delayed_112__120_,chained_data_delayed_112__119_,
  chained_data_delayed_112__118_,chained_data_delayed_112__117_,chained_data_delayed_112__116_,
  chained_data_delayed_112__115_,chained_data_delayed_112__114_,chained_data_delayed_112__113_,
  chained_data_delayed_112__112_,chained_data_delayed_112__111_,
  chained_data_delayed_112__110_,chained_data_delayed_112__109_,chained_data_delayed_112__108_,
  chained_data_delayed_112__107_,chained_data_delayed_112__106_,
  chained_data_delayed_112__105_,chained_data_delayed_112__104_,chained_data_delayed_112__103_,
  chained_data_delayed_112__102_,chained_data_delayed_112__101_,
  chained_data_delayed_112__100_,chained_data_delayed_112__99_,chained_data_delayed_112__98_,
  chained_data_delayed_112__97_,chained_data_delayed_112__96_,chained_data_delayed_112__95_,
  chained_data_delayed_112__94_,chained_data_delayed_112__93_,
  chained_data_delayed_112__92_,chained_data_delayed_112__91_,chained_data_delayed_112__90_,
  chained_data_delayed_112__89_,chained_data_delayed_112__88_,chained_data_delayed_112__87_,
  chained_data_delayed_112__86_,chained_data_delayed_112__85_,
  chained_data_delayed_112__84_,chained_data_delayed_112__83_,chained_data_delayed_112__82_,
  chained_data_delayed_112__81_,chained_data_delayed_112__80_,chained_data_delayed_112__79_,
  chained_data_delayed_112__78_,chained_data_delayed_112__77_,
  chained_data_delayed_112__76_,chained_data_delayed_112__75_,chained_data_delayed_112__74_,
  chained_data_delayed_112__73_,chained_data_delayed_112__72_,chained_data_delayed_112__71_,
  chained_data_delayed_112__70_,chained_data_delayed_112__69_,
  chained_data_delayed_112__68_,chained_data_delayed_112__67_,chained_data_delayed_112__66_,
  chained_data_delayed_112__65_,chained_data_delayed_112__64_,chained_data_delayed_112__63_,
  chained_data_delayed_112__62_,chained_data_delayed_112__61_,
  chained_data_delayed_112__60_,chained_data_delayed_112__59_,chained_data_delayed_112__58_,
  chained_data_delayed_112__57_,chained_data_delayed_112__56_,chained_data_delayed_112__55_,
  chained_data_delayed_112__54_,chained_data_delayed_112__53_,
  chained_data_delayed_112__52_,chained_data_delayed_112__51_,chained_data_delayed_112__50_,
  chained_data_delayed_112__49_,chained_data_delayed_112__48_,chained_data_delayed_112__47_,
  chained_data_delayed_112__46_,chained_data_delayed_112__45_,
  chained_data_delayed_112__44_,chained_data_delayed_112__43_,chained_data_delayed_112__42_,
  chained_data_delayed_112__41_,chained_data_delayed_112__40_,chained_data_delayed_112__39_,
  chained_data_delayed_112__38_,chained_data_delayed_112__37_,
  chained_data_delayed_112__36_,chained_data_delayed_112__35_,chained_data_delayed_112__34_,
  chained_data_delayed_112__33_,chained_data_delayed_112__32_,chained_data_delayed_112__31_,
  chained_data_delayed_112__30_,chained_data_delayed_112__29_,
  chained_data_delayed_112__28_,chained_data_delayed_112__27_,chained_data_delayed_112__26_,
  chained_data_delayed_112__25_,chained_data_delayed_112__24_,chained_data_delayed_112__23_,
  chained_data_delayed_112__22_,chained_data_delayed_112__21_,
  chained_data_delayed_112__20_,chained_data_delayed_112__19_,chained_data_delayed_112__18_,
  chained_data_delayed_112__17_,chained_data_delayed_112__16_,chained_data_delayed_112__15_,
  chained_data_delayed_112__14_,chained_data_delayed_112__13_,
  chained_data_delayed_112__12_,chained_data_delayed_112__11_,chained_data_delayed_112__10_,
  chained_data_delayed_112__9_,chained_data_delayed_112__8_,chained_data_delayed_112__7_,
  chained_data_delayed_112__6_,chained_data_delayed_112__5_,chained_data_delayed_112__4_,
  chained_data_delayed_112__3_,chained_data_delayed_112__2_,
  chained_data_delayed_112__1_,chained_data_delayed_112__0_,chained_data_delayed_111__127_,
  chained_data_delayed_111__126_,chained_data_delayed_111__125_,chained_data_delayed_111__124_,
  chained_data_delayed_111__123_,chained_data_delayed_111__122_,
  chained_data_delayed_111__121_,chained_data_delayed_111__120_,chained_data_delayed_111__119_,
  chained_data_delayed_111__118_,chained_data_delayed_111__117_,
  chained_data_delayed_111__116_,chained_data_delayed_111__115_,chained_data_delayed_111__114_,
  chained_data_delayed_111__113_,chained_data_delayed_111__112_,chained_data_delayed_111__111_,
  chained_data_delayed_111__110_,chained_data_delayed_111__109_,
  chained_data_delayed_111__108_,chained_data_delayed_111__107_,chained_data_delayed_111__106_,
  chained_data_delayed_111__105_,chained_data_delayed_111__104_,
  chained_data_delayed_111__103_,chained_data_delayed_111__102_,chained_data_delayed_111__101_,
  chained_data_delayed_111__100_,chained_data_delayed_111__99_,chained_data_delayed_111__98_,
  chained_data_delayed_111__97_,chained_data_delayed_111__96_,
  chained_data_delayed_111__95_,chained_data_delayed_111__94_,chained_data_delayed_111__93_,
  chained_data_delayed_111__92_,chained_data_delayed_111__91_,chained_data_delayed_111__90_,
  chained_data_delayed_111__89_,chained_data_delayed_111__88_,
  chained_data_delayed_111__87_,chained_data_delayed_111__86_,chained_data_delayed_111__85_,
  chained_data_delayed_111__84_,chained_data_delayed_111__83_,chained_data_delayed_111__82_,
  chained_data_delayed_111__81_,chained_data_delayed_111__80_,
  chained_data_delayed_111__79_,chained_data_delayed_111__78_,chained_data_delayed_111__77_,
  chained_data_delayed_111__76_,chained_data_delayed_111__75_,chained_data_delayed_111__74_,
  chained_data_delayed_111__73_,chained_data_delayed_111__72_,
  chained_data_delayed_111__71_,chained_data_delayed_111__70_,chained_data_delayed_111__69_,
  chained_data_delayed_111__68_,chained_data_delayed_111__67_,chained_data_delayed_111__66_,
  chained_data_delayed_111__65_,chained_data_delayed_111__64_,
  chained_data_delayed_111__63_,chained_data_delayed_111__62_,chained_data_delayed_111__61_,
  chained_data_delayed_111__60_,chained_data_delayed_111__59_,chained_data_delayed_111__58_,
  chained_data_delayed_111__57_,chained_data_delayed_111__56_,
  chained_data_delayed_111__55_,chained_data_delayed_111__54_,chained_data_delayed_111__53_,
  chained_data_delayed_111__52_,chained_data_delayed_111__51_,chained_data_delayed_111__50_,
  chained_data_delayed_111__49_,chained_data_delayed_111__48_,
  chained_data_delayed_111__47_,chained_data_delayed_111__46_,chained_data_delayed_111__45_,
  chained_data_delayed_111__44_,chained_data_delayed_111__43_,chained_data_delayed_111__42_,
  chained_data_delayed_111__41_,chained_data_delayed_111__40_,
  chained_data_delayed_111__39_,chained_data_delayed_111__38_,chained_data_delayed_111__37_,
  chained_data_delayed_111__36_,chained_data_delayed_111__35_,chained_data_delayed_111__34_,
  chained_data_delayed_111__33_,chained_data_delayed_111__32_,
  chained_data_delayed_111__31_,chained_data_delayed_111__30_,chained_data_delayed_111__29_,
  chained_data_delayed_111__28_,chained_data_delayed_111__27_,chained_data_delayed_111__26_,
  chained_data_delayed_111__25_,chained_data_delayed_111__24_,
  chained_data_delayed_111__23_,chained_data_delayed_111__22_,chained_data_delayed_111__21_,
  chained_data_delayed_111__20_,chained_data_delayed_111__19_,chained_data_delayed_111__18_,
  chained_data_delayed_111__17_,chained_data_delayed_111__16_,
  chained_data_delayed_111__15_,chained_data_delayed_111__14_,chained_data_delayed_111__13_,
  chained_data_delayed_111__12_,chained_data_delayed_111__11_,chained_data_delayed_111__10_,
  chained_data_delayed_111__9_,chained_data_delayed_111__8_,
  chained_data_delayed_111__7_,chained_data_delayed_111__6_,chained_data_delayed_111__5_,
  chained_data_delayed_111__4_,chained_data_delayed_111__3_,chained_data_delayed_111__2_,
  chained_data_delayed_111__1_,chained_data_delayed_111__0_,
  chained_data_delayed_110__127_,chained_data_delayed_110__126_,chained_data_delayed_110__125_,
  chained_data_delayed_110__124_,chained_data_delayed_110__123_,chained_data_delayed_110__122_,
  chained_data_delayed_110__121_,chained_data_delayed_110__120_,
  chained_data_delayed_110__119_,chained_data_delayed_110__118_,chained_data_delayed_110__117_,
  chained_data_delayed_110__116_,chained_data_delayed_110__115_,
  chained_data_delayed_110__114_,chained_data_delayed_110__113_,chained_data_delayed_110__112_,
  chained_data_delayed_110__111_,chained_data_delayed_110__110_,chained_data_delayed_110__109_,
  chained_data_delayed_110__108_,chained_data_delayed_110__107_,
  chained_data_delayed_110__106_,chained_data_delayed_110__105_,chained_data_delayed_110__104_,
  chained_data_delayed_110__103_,chained_data_delayed_110__102_,
  chained_data_delayed_110__101_,chained_data_delayed_110__100_,chained_data_delayed_110__99_,
  chained_data_delayed_110__98_,chained_data_delayed_110__97_,chained_data_delayed_110__96_,
  chained_data_delayed_110__95_,chained_data_delayed_110__94_,
  chained_data_delayed_110__93_,chained_data_delayed_110__92_,chained_data_delayed_110__91_,
  chained_data_delayed_110__90_,chained_data_delayed_110__89_,chained_data_delayed_110__88_,
  chained_data_delayed_110__87_,chained_data_delayed_110__86_,
  chained_data_delayed_110__85_,chained_data_delayed_110__84_,chained_data_delayed_110__83_,
  chained_data_delayed_110__82_,chained_data_delayed_110__81_,chained_data_delayed_110__80_,
  chained_data_delayed_110__79_,chained_data_delayed_110__78_,
  chained_data_delayed_110__77_,chained_data_delayed_110__76_,chained_data_delayed_110__75_,
  chained_data_delayed_110__74_,chained_data_delayed_110__73_,chained_data_delayed_110__72_,
  chained_data_delayed_110__71_,chained_data_delayed_110__70_,
  chained_data_delayed_110__69_,chained_data_delayed_110__68_,chained_data_delayed_110__67_,
  chained_data_delayed_110__66_,chained_data_delayed_110__65_,chained_data_delayed_110__64_,
  chained_data_delayed_110__63_,chained_data_delayed_110__62_,
  chained_data_delayed_110__61_,chained_data_delayed_110__60_,chained_data_delayed_110__59_,
  chained_data_delayed_110__58_,chained_data_delayed_110__57_,chained_data_delayed_110__56_,
  chained_data_delayed_110__55_,chained_data_delayed_110__54_,
  chained_data_delayed_110__53_,chained_data_delayed_110__52_,chained_data_delayed_110__51_,
  chained_data_delayed_110__50_,chained_data_delayed_110__49_,chained_data_delayed_110__48_,
  chained_data_delayed_110__47_,chained_data_delayed_110__46_,
  chained_data_delayed_110__45_,chained_data_delayed_110__44_,chained_data_delayed_110__43_,
  chained_data_delayed_110__42_,chained_data_delayed_110__41_,chained_data_delayed_110__40_,
  chained_data_delayed_110__39_,chained_data_delayed_110__38_,
  chained_data_delayed_110__37_,chained_data_delayed_110__36_,chained_data_delayed_110__35_,
  chained_data_delayed_110__34_,chained_data_delayed_110__33_,chained_data_delayed_110__32_,
  chained_data_delayed_110__31_,chained_data_delayed_110__30_,
  chained_data_delayed_110__29_,chained_data_delayed_110__28_,chained_data_delayed_110__27_,
  chained_data_delayed_110__26_,chained_data_delayed_110__25_,chained_data_delayed_110__24_,
  chained_data_delayed_110__23_,chained_data_delayed_110__22_,
  chained_data_delayed_110__21_,chained_data_delayed_110__20_,chained_data_delayed_110__19_,
  chained_data_delayed_110__18_,chained_data_delayed_110__17_,chained_data_delayed_110__16_,
  chained_data_delayed_110__15_,chained_data_delayed_110__14_,
  chained_data_delayed_110__13_,chained_data_delayed_110__12_,chained_data_delayed_110__11_,
  chained_data_delayed_110__10_,chained_data_delayed_110__9_,chained_data_delayed_110__8_,
  chained_data_delayed_110__7_,chained_data_delayed_110__6_,
  chained_data_delayed_110__5_,chained_data_delayed_110__4_,chained_data_delayed_110__3_,
  chained_data_delayed_110__2_,chained_data_delayed_110__1_,chained_data_delayed_110__0_,
  chained_data_delayed_109__127_,chained_data_delayed_109__126_,
  chained_data_delayed_109__125_,chained_data_delayed_109__124_,chained_data_delayed_109__123_,
  chained_data_delayed_109__122_,chained_data_delayed_109__121_,chained_data_delayed_109__120_,
  chained_data_delayed_109__119_,chained_data_delayed_109__118_,
  chained_data_delayed_109__117_,chained_data_delayed_109__116_,chained_data_delayed_109__115_,
  chained_data_delayed_109__114_,chained_data_delayed_109__113_,
  chained_data_delayed_109__112_,chained_data_delayed_109__111_,chained_data_delayed_109__110_,
  chained_data_delayed_109__109_,chained_data_delayed_109__108_,chained_data_delayed_109__107_,
  chained_data_delayed_109__106_,chained_data_delayed_109__105_,
  chained_data_delayed_109__104_,chained_data_delayed_109__103_,chained_data_delayed_109__102_,
  chained_data_delayed_109__101_,chained_data_delayed_109__100_,
  chained_data_delayed_109__99_,chained_data_delayed_109__98_,chained_data_delayed_109__97_,
  chained_data_delayed_109__96_,chained_data_delayed_109__95_,chained_data_delayed_109__94_,
  chained_data_delayed_109__93_,chained_data_delayed_109__92_,
  chained_data_delayed_109__91_,chained_data_delayed_109__90_,chained_data_delayed_109__89_,
  chained_data_delayed_109__88_,chained_data_delayed_109__87_,chained_data_delayed_109__86_,
  chained_data_delayed_109__85_,chained_data_delayed_109__84_,
  chained_data_delayed_109__83_,chained_data_delayed_109__82_,chained_data_delayed_109__81_,
  chained_data_delayed_109__80_,chained_data_delayed_109__79_,chained_data_delayed_109__78_,
  chained_data_delayed_109__77_,chained_data_delayed_109__76_,
  chained_data_delayed_109__75_,chained_data_delayed_109__74_,chained_data_delayed_109__73_,
  chained_data_delayed_109__72_,chained_data_delayed_109__71_,chained_data_delayed_109__70_,
  chained_data_delayed_109__69_,chained_data_delayed_109__68_,
  chained_data_delayed_109__67_,chained_data_delayed_109__66_,chained_data_delayed_109__65_,
  chained_data_delayed_109__64_,chained_data_delayed_109__63_,chained_data_delayed_109__62_,
  chained_data_delayed_109__61_,chained_data_delayed_109__60_,
  chained_data_delayed_109__59_,chained_data_delayed_109__58_,chained_data_delayed_109__57_,
  chained_data_delayed_109__56_,chained_data_delayed_109__55_,chained_data_delayed_109__54_,
  chained_data_delayed_109__53_,chained_data_delayed_109__52_,
  chained_data_delayed_109__51_,chained_data_delayed_109__50_,chained_data_delayed_109__49_,
  chained_data_delayed_109__48_,chained_data_delayed_109__47_,chained_data_delayed_109__46_,
  chained_data_delayed_109__45_,chained_data_delayed_109__44_,
  chained_data_delayed_109__43_,chained_data_delayed_109__42_,chained_data_delayed_109__41_,
  chained_data_delayed_109__40_,chained_data_delayed_109__39_,chained_data_delayed_109__38_,
  chained_data_delayed_109__37_,chained_data_delayed_109__36_,
  chained_data_delayed_109__35_,chained_data_delayed_109__34_,chained_data_delayed_109__33_,
  chained_data_delayed_109__32_,chained_data_delayed_109__31_,chained_data_delayed_109__30_,
  chained_data_delayed_109__29_,chained_data_delayed_109__28_,
  chained_data_delayed_109__27_,chained_data_delayed_109__26_,chained_data_delayed_109__25_,
  chained_data_delayed_109__24_,chained_data_delayed_109__23_,chained_data_delayed_109__22_,
  chained_data_delayed_109__21_,chained_data_delayed_109__20_,
  chained_data_delayed_109__19_,chained_data_delayed_109__18_,chained_data_delayed_109__17_,
  chained_data_delayed_109__16_,chained_data_delayed_109__15_,chained_data_delayed_109__14_,
  chained_data_delayed_109__13_,chained_data_delayed_109__12_,
  chained_data_delayed_109__11_,chained_data_delayed_109__10_,chained_data_delayed_109__9_,
  chained_data_delayed_109__8_,chained_data_delayed_109__7_,chained_data_delayed_109__6_,
  chained_data_delayed_109__5_,chained_data_delayed_109__4_,chained_data_delayed_109__3_,
  chained_data_delayed_109__2_,chained_data_delayed_109__1_,
  chained_data_delayed_109__0_,chained_data_delayed_116__127_,chained_data_delayed_116__126_,
  chained_data_delayed_116__125_,chained_data_delayed_116__124_,
  chained_data_delayed_116__123_,chained_data_delayed_116__122_,chained_data_delayed_116__121_,
  chained_data_delayed_116__120_,chained_data_delayed_116__119_,chained_data_delayed_116__118_,
  chained_data_delayed_116__117_,chained_data_delayed_116__116_,
  chained_data_delayed_116__115_,chained_data_delayed_116__114_,chained_data_delayed_116__113_,
  chained_data_delayed_116__112_,chained_data_delayed_116__111_,
  chained_data_delayed_116__110_,chained_data_delayed_116__109_,chained_data_delayed_116__108_,
  chained_data_delayed_116__107_,chained_data_delayed_116__106_,chained_data_delayed_116__105_,
  chained_data_delayed_116__104_,chained_data_delayed_116__103_,
  chained_data_delayed_116__102_,chained_data_delayed_116__101_,chained_data_delayed_116__100_,
  chained_data_delayed_116__99_,chained_data_delayed_116__98_,
  chained_data_delayed_116__97_,chained_data_delayed_116__96_,chained_data_delayed_116__95_,
  chained_data_delayed_116__94_,chained_data_delayed_116__93_,chained_data_delayed_116__92_,
  chained_data_delayed_116__91_,chained_data_delayed_116__90_,
  chained_data_delayed_116__89_,chained_data_delayed_116__88_,chained_data_delayed_116__87_,
  chained_data_delayed_116__86_,chained_data_delayed_116__85_,chained_data_delayed_116__84_,
  chained_data_delayed_116__83_,chained_data_delayed_116__82_,
  chained_data_delayed_116__81_,chained_data_delayed_116__80_,chained_data_delayed_116__79_,
  chained_data_delayed_116__78_,chained_data_delayed_116__77_,chained_data_delayed_116__76_,
  chained_data_delayed_116__75_,chained_data_delayed_116__74_,
  chained_data_delayed_116__73_,chained_data_delayed_116__72_,chained_data_delayed_116__71_,
  chained_data_delayed_116__70_,chained_data_delayed_116__69_,chained_data_delayed_116__68_,
  chained_data_delayed_116__67_,chained_data_delayed_116__66_,
  chained_data_delayed_116__65_,chained_data_delayed_116__64_,chained_data_delayed_116__63_,
  chained_data_delayed_116__62_,chained_data_delayed_116__61_,chained_data_delayed_116__60_,
  chained_data_delayed_116__59_,chained_data_delayed_116__58_,
  chained_data_delayed_116__57_,chained_data_delayed_116__56_,chained_data_delayed_116__55_,
  chained_data_delayed_116__54_,chained_data_delayed_116__53_,chained_data_delayed_116__52_,
  chained_data_delayed_116__51_,chained_data_delayed_116__50_,
  chained_data_delayed_116__49_,chained_data_delayed_116__48_,chained_data_delayed_116__47_,
  chained_data_delayed_116__46_,chained_data_delayed_116__45_,chained_data_delayed_116__44_,
  chained_data_delayed_116__43_,chained_data_delayed_116__42_,
  chained_data_delayed_116__41_,chained_data_delayed_116__40_,chained_data_delayed_116__39_,
  chained_data_delayed_116__38_,chained_data_delayed_116__37_,chained_data_delayed_116__36_,
  chained_data_delayed_116__35_,chained_data_delayed_116__34_,
  chained_data_delayed_116__33_,chained_data_delayed_116__32_,chained_data_delayed_116__31_,
  chained_data_delayed_116__30_,chained_data_delayed_116__29_,chained_data_delayed_116__28_,
  chained_data_delayed_116__27_,chained_data_delayed_116__26_,
  chained_data_delayed_116__25_,chained_data_delayed_116__24_,chained_data_delayed_116__23_,
  chained_data_delayed_116__22_,chained_data_delayed_116__21_,chained_data_delayed_116__20_,
  chained_data_delayed_116__19_,chained_data_delayed_116__18_,
  chained_data_delayed_116__17_,chained_data_delayed_116__16_,chained_data_delayed_116__15_,
  chained_data_delayed_116__14_,chained_data_delayed_116__13_,chained_data_delayed_116__12_,
  chained_data_delayed_116__11_,chained_data_delayed_116__10_,
  chained_data_delayed_116__9_,chained_data_delayed_116__8_,chained_data_delayed_116__7_,
  chained_data_delayed_116__6_,chained_data_delayed_116__5_,chained_data_delayed_116__4_,
  chained_data_delayed_116__3_,chained_data_delayed_116__2_,chained_data_delayed_116__1_,
  chained_data_delayed_116__0_,chained_data_delayed_115__127_,
  chained_data_delayed_115__126_,chained_data_delayed_115__125_,chained_data_delayed_115__124_,
  chained_data_delayed_115__123_,chained_data_delayed_115__122_,
  chained_data_delayed_115__121_,chained_data_delayed_115__120_,chained_data_delayed_115__119_,
  chained_data_delayed_115__118_,chained_data_delayed_115__117_,chained_data_delayed_115__116_,
  chained_data_delayed_115__115_,chained_data_delayed_115__114_,
  chained_data_delayed_115__113_,chained_data_delayed_115__112_,chained_data_delayed_115__111_,
  chained_data_delayed_115__110_,chained_data_delayed_115__109_,
  chained_data_delayed_115__108_,chained_data_delayed_115__107_,chained_data_delayed_115__106_,
  chained_data_delayed_115__105_,chained_data_delayed_115__104_,chained_data_delayed_115__103_,
  chained_data_delayed_115__102_,chained_data_delayed_115__101_,
  chained_data_delayed_115__100_,chained_data_delayed_115__99_,chained_data_delayed_115__98_,
  chained_data_delayed_115__97_,chained_data_delayed_115__96_,
  chained_data_delayed_115__95_,chained_data_delayed_115__94_,chained_data_delayed_115__93_,
  chained_data_delayed_115__92_,chained_data_delayed_115__91_,chained_data_delayed_115__90_,
  chained_data_delayed_115__89_,chained_data_delayed_115__88_,
  chained_data_delayed_115__87_,chained_data_delayed_115__86_,chained_data_delayed_115__85_,
  chained_data_delayed_115__84_,chained_data_delayed_115__83_,chained_data_delayed_115__82_,
  chained_data_delayed_115__81_,chained_data_delayed_115__80_,
  chained_data_delayed_115__79_,chained_data_delayed_115__78_,chained_data_delayed_115__77_,
  chained_data_delayed_115__76_,chained_data_delayed_115__75_,chained_data_delayed_115__74_,
  chained_data_delayed_115__73_,chained_data_delayed_115__72_,
  chained_data_delayed_115__71_,chained_data_delayed_115__70_,chained_data_delayed_115__69_,
  chained_data_delayed_115__68_,chained_data_delayed_115__67_,chained_data_delayed_115__66_,
  chained_data_delayed_115__65_,chained_data_delayed_115__64_,
  chained_data_delayed_115__63_,chained_data_delayed_115__62_,chained_data_delayed_115__61_,
  chained_data_delayed_115__60_,chained_data_delayed_115__59_,chained_data_delayed_115__58_,
  chained_data_delayed_115__57_,chained_data_delayed_115__56_,
  chained_data_delayed_115__55_,chained_data_delayed_115__54_,chained_data_delayed_115__53_,
  chained_data_delayed_115__52_,chained_data_delayed_115__51_,chained_data_delayed_115__50_,
  chained_data_delayed_115__49_,chained_data_delayed_115__48_,
  chained_data_delayed_115__47_,chained_data_delayed_115__46_,chained_data_delayed_115__45_,
  chained_data_delayed_115__44_,chained_data_delayed_115__43_,chained_data_delayed_115__42_,
  chained_data_delayed_115__41_,chained_data_delayed_115__40_,
  chained_data_delayed_115__39_,chained_data_delayed_115__38_,chained_data_delayed_115__37_,
  chained_data_delayed_115__36_,chained_data_delayed_115__35_,chained_data_delayed_115__34_,
  chained_data_delayed_115__33_,chained_data_delayed_115__32_,
  chained_data_delayed_115__31_,chained_data_delayed_115__30_,chained_data_delayed_115__29_,
  chained_data_delayed_115__28_,chained_data_delayed_115__27_,chained_data_delayed_115__26_,
  chained_data_delayed_115__25_,chained_data_delayed_115__24_,
  chained_data_delayed_115__23_,chained_data_delayed_115__22_,chained_data_delayed_115__21_,
  chained_data_delayed_115__20_,chained_data_delayed_115__19_,chained_data_delayed_115__18_,
  chained_data_delayed_115__17_,chained_data_delayed_115__16_,
  chained_data_delayed_115__15_,chained_data_delayed_115__14_,chained_data_delayed_115__13_,
  chained_data_delayed_115__12_,chained_data_delayed_115__11_,chained_data_delayed_115__10_,
  chained_data_delayed_115__9_,chained_data_delayed_115__8_,chained_data_delayed_115__7_,
  chained_data_delayed_115__6_,chained_data_delayed_115__5_,
  chained_data_delayed_115__4_,chained_data_delayed_115__3_,chained_data_delayed_115__2_,
  chained_data_delayed_115__1_,chained_data_delayed_115__0_,chained_data_delayed_114__127_,
  chained_data_delayed_114__126_,chained_data_delayed_114__125_,
  chained_data_delayed_114__124_,chained_data_delayed_114__123_,chained_data_delayed_114__122_,
  chained_data_delayed_114__121_,chained_data_delayed_114__120_,
  chained_data_delayed_114__119_,chained_data_delayed_114__118_,chained_data_delayed_114__117_,
  chained_data_delayed_114__116_,chained_data_delayed_114__115_,chained_data_delayed_114__114_,
  chained_data_delayed_114__113_,chained_data_delayed_114__112_,
  chained_data_delayed_114__111_,chained_data_delayed_114__110_,chained_data_delayed_114__109_,
  chained_data_delayed_114__108_,chained_data_delayed_114__107_,
  chained_data_delayed_114__106_,chained_data_delayed_114__105_,chained_data_delayed_114__104_,
  chained_data_delayed_114__103_,chained_data_delayed_114__102_,chained_data_delayed_114__101_,
  chained_data_delayed_114__100_,chained_data_delayed_114__99_,
  chained_data_delayed_114__98_,chained_data_delayed_114__97_,chained_data_delayed_114__96_,
  chained_data_delayed_114__95_,chained_data_delayed_114__94_,chained_data_delayed_114__93_,
  chained_data_delayed_114__92_,chained_data_delayed_114__91_,
  chained_data_delayed_114__90_,chained_data_delayed_114__89_,chained_data_delayed_114__88_,
  chained_data_delayed_114__87_,chained_data_delayed_114__86_,chained_data_delayed_114__85_,
  chained_data_delayed_114__84_,chained_data_delayed_114__83_,
  chained_data_delayed_114__82_,chained_data_delayed_114__81_,chained_data_delayed_114__80_,
  chained_data_delayed_114__79_,chained_data_delayed_114__78_,chained_data_delayed_114__77_,
  chained_data_delayed_114__76_,chained_data_delayed_114__75_,
  chained_data_delayed_114__74_,chained_data_delayed_114__73_,chained_data_delayed_114__72_,
  chained_data_delayed_114__71_,chained_data_delayed_114__70_,chained_data_delayed_114__69_,
  chained_data_delayed_114__68_,chained_data_delayed_114__67_,
  chained_data_delayed_114__66_,chained_data_delayed_114__65_,chained_data_delayed_114__64_,
  chained_data_delayed_114__63_,chained_data_delayed_114__62_,chained_data_delayed_114__61_,
  chained_data_delayed_114__60_,chained_data_delayed_114__59_,
  chained_data_delayed_114__58_,chained_data_delayed_114__57_,chained_data_delayed_114__56_,
  chained_data_delayed_114__55_,chained_data_delayed_114__54_,chained_data_delayed_114__53_,
  chained_data_delayed_114__52_,chained_data_delayed_114__51_,
  chained_data_delayed_114__50_,chained_data_delayed_114__49_,chained_data_delayed_114__48_,
  chained_data_delayed_114__47_,chained_data_delayed_114__46_,chained_data_delayed_114__45_,
  chained_data_delayed_114__44_,chained_data_delayed_114__43_,
  chained_data_delayed_114__42_,chained_data_delayed_114__41_,chained_data_delayed_114__40_,
  chained_data_delayed_114__39_,chained_data_delayed_114__38_,chained_data_delayed_114__37_,
  chained_data_delayed_114__36_,chained_data_delayed_114__35_,
  chained_data_delayed_114__34_,chained_data_delayed_114__33_,chained_data_delayed_114__32_,
  chained_data_delayed_114__31_,chained_data_delayed_114__30_,chained_data_delayed_114__29_,
  chained_data_delayed_114__28_,chained_data_delayed_114__27_,
  chained_data_delayed_114__26_,chained_data_delayed_114__25_,chained_data_delayed_114__24_,
  chained_data_delayed_114__23_,chained_data_delayed_114__22_,chained_data_delayed_114__21_,
  chained_data_delayed_114__20_,chained_data_delayed_114__19_,
  chained_data_delayed_114__18_,chained_data_delayed_114__17_,chained_data_delayed_114__16_,
  chained_data_delayed_114__15_,chained_data_delayed_114__14_,chained_data_delayed_114__13_,
  chained_data_delayed_114__12_,chained_data_delayed_114__11_,
  chained_data_delayed_114__10_,chained_data_delayed_114__9_,chained_data_delayed_114__8_,
  chained_data_delayed_114__7_,chained_data_delayed_114__6_,chained_data_delayed_114__5_,
  chained_data_delayed_114__4_,chained_data_delayed_114__3_,
  chained_data_delayed_114__2_,chained_data_delayed_114__1_,chained_data_delayed_114__0_,
  chained_data_delayed_113__127_,chained_data_delayed_113__126_,chained_data_delayed_113__125_,
  chained_data_delayed_113__124_,chained_data_delayed_113__123_,
  chained_data_delayed_113__122_,chained_data_delayed_113__121_,chained_data_delayed_113__120_,
  chained_data_delayed_113__119_,chained_data_delayed_113__118_,
  chained_data_delayed_113__117_,chained_data_delayed_113__116_,chained_data_delayed_113__115_,
  chained_data_delayed_113__114_,chained_data_delayed_113__113_,chained_data_delayed_113__112_,
  chained_data_delayed_113__111_,chained_data_delayed_113__110_,
  chained_data_delayed_113__109_,chained_data_delayed_113__108_,chained_data_delayed_113__107_,
  chained_data_delayed_113__106_,chained_data_delayed_113__105_,
  chained_data_delayed_113__104_,chained_data_delayed_113__103_,chained_data_delayed_113__102_,
  chained_data_delayed_113__101_,chained_data_delayed_113__100_,chained_data_delayed_113__99_,
  chained_data_delayed_113__98_,chained_data_delayed_113__97_,
  chained_data_delayed_113__96_,chained_data_delayed_113__95_,chained_data_delayed_113__94_,
  chained_data_delayed_113__93_,chained_data_delayed_113__92_,chained_data_delayed_113__91_,
  chained_data_delayed_113__90_,chained_data_delayed_113__89_,
  chained_data_delayed_113__88_,chained_data_delayed_113__87_,chained_data_delayed_113__86_,
  chained_data_delayed_113__85_,chained_data_delayed_113__84_,chained_data_delayed_113__83_,
  chained_data_delayed_113__82_,chained_data_delayed_113__81_,
  chained_data_delayed_113__80_,chained_data_delayed_113__79_,chained_data_delayed_113__78_,
  chained_data_delayed_113__77_,chained_data_delayed_113__76_,chained_data_delayed_113__75_,
  chained_data_delayed_113__74_,chained_data_delayed_113__73_,
  chained_data_delayed_113__72_,chained_data_delayed_113__71_,chained_data_delayed_113__70_,
  chained_data_delayed_113__69_,chained_data_delayed_113__68_,chained_data_delayed_113__67_,
  chained_data_delayed_113__66_,chained_data_delayed_113__65_,
  chained_data_delayed_113__64_,chained_data_delayed_113__63_,chained_data_delayed_113__62_,
  chained_data_delayed_113__61_,chained_data_delayed_113__60_,chained_data_delayed_113__59_,
  chained_data_delayed_113__58_,chained_data_delayed_113__57_,
  chained_data_delayed_113__56_,chained_data_delayed_113__55_,chained_data_delayed_113__54_,
  chained_data_delayed_113__53_,chained_data_delayed_113__52_,chained_data_delayed_113__51_,
  chained_data_delayed_113__50_,chained_data_delayed_113__49_,
  chained_data_delayed_113__48_,chained_data_delayed_113__47_,chained_data_delayed_113__46_,
  chained_data_delayed_113__45_,chained_data_delayed_113__44_,chained_data_delayed_113__43_,
  chained_data_delayed_113__42_,chained_data_delayed_113__41_,
  chained_data_delayed_113__40_,chained_data_delayed_113__39_,chained_data_delayed_113__38_,
  chained_data_delayed_113__37_,chained_data_delayed_113__36_,chained_data_delayed_113__35_,
  chained_data_delayed_113__34_,chained_data_delayed_113__33_,
  chained_data_delayed_113__32_,chained_data_delayed_113__31_,chained_data_delayed_113__30_,
  chained_data_delayed_113__29_,chained_data_delayed_113__28_,chained_data_delayed_113__27_,
  chained_data_delayed_113__26_,chained_data_delayed_113__25_,
  chained_data_delayed_113__24_,chained_data_delayed_113__23_,chained_data_delayed_113__22_,
  chained_data_delayed_113__21_,chained_data_delayed_113__20_,chained_data_delayed_113__19_,
  chained_data_delayed_113__18_,chained_data_delayed_113__17_,
  chained_data_delayed_113__16_,chained_data_delayed_113__15_,chained_data_delayed_113__14_,
  chained_data_delayed_113__13_,chained_data_delayed_113__12_,chained_data_delayed_113__11_,
  chained_data_delayed_113__10_,chained_data_delayed_113__9_,
  chained_data_delayed_113__8_,chained_data_delayed_113__7_,chained_data_delayed_113__6_,
  chained_data_delayed_113__5_,chained_data_delayed_113__4_,chained_data_delayed_113__3_,
  chained_data_delayed_113__2_,chained_data_delayed_113__1_,chained_data_delayed_113__0_,
  chained_data_delayed_120__127_,chained_data_delayed_120__126_,
  chained_data_delayed_120__125_,chained_data_delayed_120__124_,chained_data_delayed_120__123_,
  chained_data_delayed_120__122_,chained_data_delayed_120__121_,
  chained_data_delayed_120__120_,chained_data_delayed_120__119_,chained_data_delayed_120__118_,
  chained_data_delayed_120__117_,chained_data_delayed_120__116_,
  chained_data_delayed_120__115_,chained_data_delayed_120__114_,chained_data_delayed_120__113_,
  chained_data_delayed_120__112_,chained_data_delayed_120__111_,chained_data_delayed_120__110_,
  chained_data_delayed_120__109_,chained_data_delayed_120__108_,
  chained_data_delayed_120__107_,chained_data_delayed_120__106_,chained_data_delayed_120__105_,
  chained_data_delayed_120__104_,chained_data_delayed_120__103_,
  chained_data_delayed_120__102_,chained_data_delayed_120__101_,chained_data_delayed_120__100_,
  chained_data_delayed_120__99_,chained_data_delayed_120__98_,chained_data_delayed_120__97_,
  chained_data_delayed_120__96_,chained_data_delayed_120__95_,
  chained_data_delayed_120__94_,chained_data_delayed_120__93_,chained_data_delayed_120__92_,
  chained_data_delayed_120__91_,chained_data_delayed_120__90_,chained_data_delayed_120__89_,
  chained_data_delayed_120__88_,chained_data_delayed_120__87_,
  chained_data_delayed_120__86_,chained_data_delayed_120__85_,chained_data_delayed_120__84_,
  chained_data_delayed_120__83_,chained_data_delayed_120__82_,chained_data_delayed_120__81_,
  chained_data_delayed_120__80_,chained_data_delayed_120__79_,
  chained_data_delayed_120__78_,chained_data_delayed_120__77_,chained_data_delayed_120__76_,
  chained_data_delayed_120__75_,chained_data_delayed_120__74_,chained_data_delayed_120__73_,
  chained_data_delayed_120__72_,chained_data_delayed_120__71_,
  chained_data_delayed_120__70_,chained_data_delayed_120__69_,chained_data_delayed_120__68_,
  chained_data_delayed_120__67_,chained_data_delayed_120__66_,chained_data_delayed_120__65_,
  chained_data_delayed_120__64_,chained_data_delayed_120__63_,
  chained_data_delayed_120__62_,chained_data_delayed_120__61_,chained_data_delayed_120__60_,
  chained_data_delayed_120__59_,chained_data_delayed_120__58_,chained_data_delayed_120__57_,
  chained_data_delayed_120__56_,chained_data_delayed_120__55_,
  chained_data_delayed_120__54_,chained_data_delayed_120__53_,chained_data_delayed_120__52_,
  chained_data_delayed_120__51_,chained_data_delayed_120__50_,chained_data_delayed_120__49_,
  chained_data_delayed_120__48_,chained_data_delayed_120__47_,
  chained_data_delayed_120__46_,chained_data_delayed_120__45_,chained_data_delayed_120__44_,
  chained_data_delayed_120__43_,chained_data_delayed_120__42_,chained_data_delayed_120__41_,
  chained_data_delayed_120__40_,chained_data_delayed_120__39_,
  chained_data_delayed_120__38_,chained_data_delayed_120__37_,chained_data_delayed_120__36_,
  chained_data_delayed_120__35_,chained_data_delayed_120__34_,chained_data_delayed_120__33_,
  chained_data_delayed_120__32_,chained_data_delayed_120__31_,
  chained_data_delayed_120__30_,chained_data_delayed_120__29_,chained_data_delayed_120__28_,
  chained_data_delayed_120__27_,chained_data_delayed_120__26_,chained_data_delayed_120__25_,
  chained_data_delayed_120__24_,chained_data_delayed_120__23_,
  chained_data_delayed_120__22_,chained_data_delayed_120__21_,chained_data_delayed_120__20_,
  chained_data_delayed_120__19_,chained_data_delayed_120__18_,chained_data_delayed_120__17_,
  chained_data_delayed_120__16_,chained_data_delayed_120__15_,
  chained_data_delayed_120__14_,chained_data_delayed_120__13_,chained_data_delayed_120__12_,
  chained_data_delayed_120__11_,chained_data_delayed_120__10_,chained_data_delayed_120__9_,
  chained_data_delayed_120__8_,chained_data_delayed_120__7_,
  chained_data_delayed_120__6_,chained_data_delayed_120__5_,chained_data_delayed_120__4_,
  chained_data_delayed_120__3_,chained_data_delayed_120__2_,chained_data_delayed_120__1_,
  chained_data_delayed_120__0_,chained_data_delayed_119__127_,chained_data_delayed_119__126_,
  chained_data_delayed_119__125_,chained_data_delayed_119__124_,
  chained_data_delayed_119__123_,chained_data_delayed_119__122_,chained_data_delayed_119__121_,
  chained_data_delayed_119__120_,chained_data_delayed_119__119_,
  chained_data_delayed_119__118_,chained_data_delayed_119__117_,chained_data_delayed_119__116_,
  chained_data_delayed_119__115_,chained_data_delayed_119__114_,
  chained_data_delayed_119__113_,chained_data_delayed_119__112_,chained_data_delayed_119__111_,
  chained_data_delayed_119__110_,chained_data_delayed_119__109_,chained_data_delayed_119__108_,
  chained_data_delayed_119__107_,chained_data_delayed_119__106_,
  chained_data_delayed_119__105_,chained_data_delayed_119__104_,chained_data_delayed_119__103_,
  chained_data_delayed_119__102_,chained_data_delayed_119__101_,
  chained_data_delayed_119__100_,chained_data_delayed_119__99_,chained_data_delayed_119__98_,
  chained_data_delayed_119__97_,chained_data_delayed_119__96_,chained_data_delayed_119__95_,
  chained_data_delayed_119__94_,chained_data_delayed_119__93_,
  chained_data_delayed_119__92_,chained_data_delayed_119__91_,chained_data_delayed_119__90_,
  chained_data_delayed_119__89_,chained_data_delayed_119__88_,chained_data_delayed_119__87_,
  chained_data_delayed_119__86_,chained_data_delayed_119__85_,
  chained_data_delayed_119__84_,chained_data_delayed_119__83_,chained_data_delayed_119__82_,
  chained_data_delayed_119__81_,chained_data_delayed_119__80_,chained_data_delayed_119__79_,
  chained_data_delayed_119__78_,chained_data_delayed_119__77_,
  chained_data_delayed_119__76_,chained_data_delayed_119__75_,chained_data_delayed_119__74_,
  chained_data_delayed_119__73_,chained_data_delayed_119__72_,chained_data_delayed_119__71_,
  chained_data_delayed_119__70_,chained_data_delayed_119__69_,
  chained_data_delayed_119__68_,chained_data_delayed_119__67_,chained_data_delayed_119__66_,
  chained_data_delayed_119__65_,chained_data_delayed_119__64_,chained_data_delayed_119__63_,
  chained_data_delayed_119__62_,chained_data_delayed_119__61_,
  chained_data_delayed_119__60_,chained_data_delayed_119__59_,chained_data_delayed_119__58_,
  chained_data_delayed_119__57_,chained_data_delayed_119__56_,chained_data_delayed_119__55_,
  chained_data_delayed_119__54_,chained_data_delayed_119__53_,
  chained_data_delayed_119__52_,chained_data_delayed_119__51_,chained_data_delayed_119__50_,
  chained_data_delayed_119__49_,chained_data_delayed_119__48_,chained_data_delayed_119__47_,
  chained_data_delayed_119__46_,chained_data_delayed_119__45_,
  chained_data_delayed_119__44_,chained_data_delayed_119__43_,chained_data_delayed_119__42_,
  chained_data_delayed_119__41_,chained_data_delayed_119__40_,chained_data_delayed_119__39_,
  chained_data_delayed_119__38_,chained_data_delayed_119__37_,
  chained_data_delayed_119__36_,chained_data_delayed_119__35_,chained_data_delayed_119__34_,
  chained_data_delayed_119__33_,chained_data_delayed_119__32_,chained_data_delayed_119__31_,
  chained_data_delayed_119__30_,chained_data_delayed_119__29_,
  chained_data_delayed_119__28_,chained_data_delayed_119__27_,chained_data_delayed_119__26_,
  chained_data_delayed_119__25_,chained_data_delayed_119__24_,chained_data_delayed_119__23_,
  chained_data_delayed_119__22_,chained_data_delayed_119__21_,
  chained_data_delayed_119__20_,chained_data_delayed_119__19_,chained_data_delayed_119__18_,
  chained_data_delayed_119__17_,chained_data_delayed_119__16_,chained_data_delayed_119__15_,
  chained_data_delayed_119__14_,chained_data_delayed_119__13_,
  chained_data_delayed_119__12_,chained_data_delayed_119__11_,chained_data_delayed_119__10_,
  chained_data_delayed_119__9_,chained_data_delayed_119__8_,chained_data_delayed_119__7_,
  chained_data_delayed_119__6_,chained_data_delayed_119__5_,chained_data_delayed_119__4_,
  chained_data_delayed_119__3_,chained_data_delayed_119__2_,
  chained_data_delayed_119__1_,chained_data_delayed_119__0_,chained_data_delayed_118__127_,
  chained_data_delayed_118__126_,chained_data_delayed_118__125_,chained_data_delayed_118__124_,
  chained_data_delayed_118__123_,chained_data_delayed_118__122_,
  chained_data_delayed_118__121_,chained_data_delayed_118__120_,chained_data_delayed_118__119_,
  chained_data_delayed_118__118_,chained_data_delayed_118__117_,
  chained_data_delayed_118__116_,chained_data_delayed_118__115_,chained_data_delayed_118__114_,
  chained_data_delayed_118__113_,chained_data_delayed_118__112_,
  chained_data_delayed_118__111_,chained_data_delayed_118__110_,chained_data_delayed_118__109_,
  chained_data_delayed_118__108_,chained_data_delayed_118__107_,chained_data_delayed_118__106_,
  chained_data_delayed_118__105_,chained_data_delayed_118__104_,
  chained_data_delayed_118__103_,chained_data_delayed_118__102_,chained_data_delayed_118__101_,
  chained_data_delayed_118__100_,chained_data_delayed_118__99_,
  chained_data_delayed_118__98_,chained_data_delayed_118__97_,chained_data_delayed_118__96_,
  chained_data_delayed_118__95_,chained_data_delayed_118__94_,chained_data_delayed_118__93_,
  chained_data_delayed_118__92_,chained_data_delayed_118__91_,
  chained_data_delayed_118__90_,chained_data_delayed_118__89_,chained_data_delayed_118__88_,
  chained_data_delayed_118__87_,chained_data_delayed_118__86_,chained_data_delayed_118__85_,
  chained_data_delayed_118__84_,chained_data_delayed_118__83_,
  chained_data_delayed_118__82_,chained_data_delayed_118__81_,chained_data_delayed_118__80_,
  chained_data_delayed_118__79_,chained_data_delayed_118__78_,chained_data_delayed_118__77_,
  chained_data_delayed_118__76_,chained_data_delayed_118__75_,
  chained_data_delayed_118__74_,chained_data_delayed_118__73_,chained_data_delayed_118__72_,
  chained_data_delayed_118__71_,chained_data_delayed_118__70_,chained_data_delayed_118__69_,
  chained_data_delayed_118__68_,chained_data_delayed_118__67_,
  chained_data_delayed_118__66_,chained_data_delayed_118__65_,chained_data_delayed_118__64_,
  chained_data_delayed_118__63_,chained_data_delayed_118__62_,chained_data_delayed_118__61_,
  chained_data_delayed_118__60_,chained_data_delayed_118__59_,
  chained_data_delayed_118__58_,chained_data_delayed_118__57_,chained_data_delayed_118__56_,
  chained_data_delayed_118__55_,chained_data_delayed_118__54_,chained_data_delayed_118__53_,
  chained_data_delayed_118__52_,chained_data_delayed_118__51_,
  chained_data_delayed_118__50_,chained_data_delayed_118__49_,chained_data_delayed_118__48_,
  chained_data_delayed_118__47_,chained_data_delayed_118__46_,chained_data_delayed_118__45_,
  chained_data_delayed_118__44_,chained_data_delayed_118__43_,
  chained_data_delayed_118__42_,chained_data_delayed_118__41_,chained_data_delayed_118__40_,
  chained_data_delayed_118__39_,chained_data_delayed_118__38_,chained_data_delayed_118__37_,
  chained_data_delayed_118__36_,chained_data_delayed_118__35_,
  chained_data_delayed_118__34_,chained_data_delayed_118__33_,chained_data_delayed_118__32_,
  chained_data_delayed_118__31_,chained_data_delayed_118__30_,chained_data_delayed_118__29_,
  chained_data_delayed_118__28_,chained_data_delayed_118__27_,
  chained_data_delayed_118__26_,chained_data_delayed_118__25_,chained_data_delayed_118__24_,
  chained_data_delayed_118__23_,chained_data_delayed_118__22_,chained_data_delayed_118__21_,
  chained_data_delayed_118__20_,chained_data_delayed_118__19_,
  chained_data_delayed_118__18_,chained_data_delayed_118__17_,chained_data_delayed_118__16_,
  chained_data_delayed_118__15_,chained_data_delayed_118__14_,chained_data_delayed_118__13_,
  chained_data_delayed_118__12_,chained_data_delayed_118__11_,
  chained_data_delayed_118__10_,chained_data_delayed_118__9_,chained_data_delayed_118__8_,
  chained_data_delayed_118__7_,chained_data_delayed_118__6_,chained_data_delayed_118__5_,
  chained_data_delayed_118__4_,chained_data_delayed_118__3_,chained_data_delayed_118__2_,
  chained_data_delayed_118__1_,chained_data_delayed_118__0_,
  chained_data_delayed_117__127_,chained_data_delayed_117__126_,chained_data_delayed_117__125_,
  chained_data_delayed_117__124_,chained_data_delayed_117__123_,chained_data_delayed_117__122_,
  chained_data_delayed_117__121_,chained_data_delayed_117__120_,
  chained_data_delayed_117__119_,chained_data_delayed_117__118_,chained_data_delayed_117__117_,
  chained_data_delayed_117__116_,chained_data_delayed_117__115_,
  chained_data_delayed_117__114_,chained_data_delayed_117__113_,chained_data_delayed_117__112_,
  chained_data_delayed_117__111_,chained_data_delayed_117__110_,
  chained_data_delayed_117__109_,chained_data_delayed_117__108_,chained_data_delayed_117__107_,
  chained_data_delayed_117__106_,chained_data_delayed_117__105_,chained_data_delayed_117__104_,
  chained_data_delayed_117__103_,chained_data_delayed_117__102_,
  chained_data_delayed_117__101_,chained_data_delayed_117__100_,chained_data_delayed_117__99_,
  chained_data_delayed_117__98_,chained_data_delayed_117__97_,chained_data_delayed_117__96_,
  chained_data_delayed_117__95_,chained_data_delayed_117__94_,
  chained_data_delayed_117__93_,chained_data_delayed_117__92_,chained_data_delayed_117__91_,
  chained_data_delayed_117__90_,chained_data_delayed_117__89_,chained_data_delayed_117__88_,
  chained_data_delayed_117__87_,chained_data_delayed_117__86_,
  chained_data_delayed_117__85_,chained_data_delayed_117__84_,chained_data_delayed_117__83_,
  chained_data_delayed_117__82_,chained_data_delayed_117__81_,chained_data_delayed_117__80_,
  chained_data_delayed_117__79_,chained_data_delayed_117__78_,
  chained_data_delayed_117__77_,chained_data_delayed_117__76_,chained_data_delayed_117__75_,
  chained_data_delayed_117__74_,chained_data_delayed_117__73_,chained_data_delayed_117__72_,
  chained_data_delayed_117__71_,chained_data_delayed_117__70_,
  chained_data_delayed_117__69_,chained_data_delayed_117__68_,chained_data_delayed_117__67_,
  chained_data_delayed_117__66_,chained_data_delayed_117__65_,chained_data_delayed_117__64_,
  chained_data_delayed_117__63_,chained_data_delayed_117__62_,
  chained_data_delayed_117__61_,chained_data_delayed_117__60_,chained_data_delayed_117__59_,
  chained_data_delayed_117__58_,chained_data_delayed_117__57_,chained_data_delayed_117__56_,
  chained_data_delayed_117__55_,chained_data_delayed_117__54_,
  chained_data_delayed_117__53_,chained_data_delayed_117__52_,chained_data_delayed_117__51_,
  chained_data_delayed_117__50_,chained_data_delayed_117__49_,chained_data_delayed_117__48_,
  chained_data_delayed_117__47_,chained_data_delayed_117__46_,
  chained_data_delayed_117__45_,chained_data_delayed_117__44_,chained_data_delayed_117__43_,
  chained_data_delayed_117__42_,chained_data_delayed_117__41_,chained_data_delayed_117__40_,
  chained_data_delayed_117__39_,chained_data_delayed_117__38_,
  chained_data_delayed_117__37_,chained_data_delayed_117__36_,chained_data_delayed_117__35_,
  chained_data_delayed_117__34_,chained_data_delayed_117__33_,chained_data_delayed_117__32_,
  chained_data_delayed_117__31_,chained_data_delayed_117__30_,
  chained_data_delayed_117__29_,chained_data_delayed_117__28_,chained_data_delayed_117__27_,
  chained_data_delayed_117__26_,chained_data_delayed_117__25_,chained_data_delayed_117__24_,
  chained_data_delayed_117__23_,chained_data_delayed_117__22_,
  chained_data_delayed_117__21_,chained_data_delayed_117__20_,chained_data_delayed_117__19_,
  chained_data_delayed_117__18_,chained_data_delayed_117__17_,chained_data_delayed_117__16_,
  chained_data_delayed_117__15_,chained_data_delayed_117__14_,
  chained_data_delayed_117__13_,chained_data_delayed_117__12_,chained_data_delayed_117__11_,
  chained_data_delayed_117__10_,chained_data_delayed_117__9_,chained_data_delayed_117__8_,
  chained_data_delayed_117__7_,chained_data_delayed_117__6_,
  chained_data_delayed_117__5_,chained_data_delayed_117__4_,chained_data_delayed_117__3_,
  chained_data_delayed_117__2_,chained_data_delayed_117__1_,chained_data_delayed_117__0_,
  chained_data_delayed_124__127_,chained_data_delayed_124__126_,
  chained_data_delayed_124__125_,chained_data_delayed_124__124_,chained_data_delayed_124__123_,
  chained_data_delayed_124__122_,chained_data_delayed_124__121_,chained_data_delayed_124__120_,
  chained_data_delayed_124__119_,chained_data_delayed_124__118_,
  chained_data_delayed_124__117_,chained_data_delayed_124__116_,chained_data_delayed_124__115_,
  chained_data_delayed_124__114_,chained_data_delayed_124__113_,
  chained_data_delayed_124__112_,chained_data_delayed_124__111_,chained_data_delayed_124__110_,
  chained_data_delayed_124__109_,chained_data_delayed_124__108_,
  chained_data_delayed_124__107_,chained_data_delayed_124__106_,chained_data_delayed_124__105_,
  chained_data_delayed_124__104_,chained_data_delayed_124__103_,chained_data_delayed_124__102_,
  chained_data_delayed_124__101_,chained_data_delayed_124__100_,
  chained_data_delayed_124__99_,chained_data_delayed_124__98_,chained_data_delayed_124__97_,
  chained_data_delayed_124__96_,chained_data_delayed_124__95_,chained_data_delayed_124__94_,
  chained_data_delayed_124__93_,chained_data_delayed_124__92_,
  chained_data_delayed_124__91_,chained_data_delayed_124__90_,chained_data_delayed_124__89_,
  chained_data_delayed_124__88_,chained_data_delayed_124__87_,chained_data_delayed_124__86_,
  chained_data_delayed_124__85_,chained_data_delayed_124__84_,
  chained_data_delayed_124__83_,chained_data_delayed_124__82_,chained_data_delayed_124__81_,
  chained_data_delayed_124__80_,chained_data_delayed_124__79_,chained_data_delayed_124__78_,
  chained_data_delayed_124__77_,chained_data_delayed_124__76_,
  chained_data_delayed_124__75_,chained_data_delayed_124__74_,chained_data_delayed_124__73_,
  chained_data_delayed_124__72_,chained_data_delayed_124__71_,chained_data_delayed_124__70_,
  chained_data_delayed_124__69_,chained_data_delayed_124__68_,
  chained_data_delayed_124__67_,chained_data_delayed_124__66_,chained_data_delayed_124__65_,
  chained_data_delayed_124__64_,chained_data_delayed_124__63_,chained_data_delayed_124__62_,
  chained_data_delayed_124__61_,chained_data_delayed_124__60_,
  chained_data_delayed_124__59_,chained_data_delayed_124__58_,chained_data_delayed_124__57_,
  chained_data_delayed_124__56_,chained_data_delayed_124__55_,chained_data_delayed_124__54_,
  chained_data_delayed_124__53_,chained_data_delayed_124__52_,
  chained_data_delayed_124__51_,chained_data_delayed_124__50_,chained_data_delayed_124__49_,
  chained_data_delayed_124__48_,chained_data_delayed_124__47_,chained_data_delayed_124__46_,
  chained_data_delayed_124__45_,chained_data_delayed_124__44_,
  chained_data_delayed_124__43_,chained_data_delayed_124__42_,chained_data_delayed_124__41_,
  chained_data_delayed_124__40_,chained_data_delayed_124__39_,chained_data_delayed_124__38_,
  chained_data_delayed_124__37_,chained_data_delayed_124__36_,
  chained_data_delayed_124__35_,chained_data_delayed_124__34_,chained_data_delayed_124__33_,
  chained_data_delayed_124__32_,chained_data_delayed_124__31_,chained_data_delayed_124__30_,
  chained_data_delayed_124__29_,chained_data_delayed_124__28_,
  chained_data_delayed_124__27_,chained_data_delayed_124__26_,chained_data_delayed_124__25_,
  chained_data_delayed_124__24_,chained_data_delayed_124__23_,chained_data_delayed_124__22_,
  chained_data_delayed_124__21_,chained_data_delayed_124__20_,
  chained_data_delayed_124__19_,chained_data_delayed_124__18_,chained_data_delayed_124__17_,
  chained_data_delayed_124__16_,chained_data_delayed_124__15_,chained_data_delayed_124__14_,
  chained_data_delayed_124__13_,chained_data_delayed_124__12_,
  chained_data_delayed_124__11_,chained_data_delayed_124__10_,chained_data_delayed_124__9_,
  chained_data_delayed_124__8_,chained_data_delayed_124__7_,chained_data_delayed_124__6_,
  chained_data_delayed_124__5_,chained_data_delayed_124__4_,
  chained_data_delayed_124__3_,chained_data_delayed_124__2_,chained_data_delayed_124__1_,
  chained_data_delayed_124__0_,chained_data_delayed_123__127_,chained_data_delayed_123__126_,
  chained_data_delayed_123__125_,chained_data_delayed_123__124_,
  chained_data_delayed_123__123_,chained_data_delayed_123__122_,chained_data_delayed_123__121_,
  chained_data_delayed_123__120_,chained_data_delayed_123__119_,chained_data_delayed_123__118_,
  chained_data_delayed_123__117_,chained_data_delayed_123__116_,
  chained_data_delayed_123__115_,chained_data_delayed_123__114_,chained_data_delayed_123__113_,
  chained_data_delayed_123__112_,chained_data_delayed_123__111_,
  chained_data_delayed_123__110_,chained_data_delayed_123__109_,chained_data_delayed_123__108_,
  chained_data_delayed_123__107_,chained_data_delayed_123__106_,
  chained_data_delayed_123__105_,chained_data_delayed_123__104_,chained_data_delayed_123__103_,
  chained_data_delayed_123__102_,chained_data_delayed_123__101_,chained_data_delayed_123__100_,
  chained_data_delayed_123__99_,chained_data_delayed_123__98_,
  chained_data_delayed_123__97_,chained_data_delayed_123__96_,chained_data_delayed_123__95_,
  chained_data_delayed_123__94_,chained_data_delayed_123__93_,chained_data_delayed_123__92_,
  chained_data_delayed_123__91_,chained_data_delayed_123__90_,
  chained_data_delayed_123__89_,chained_data_delayed_123__88_,chained_data_delayed_123__87_,
  chained_data_delayed_123__86_,chained_data_delayed_123__85_,chained_data_delayed_123__84_,
  chained_data_delayed_123__83_,chained_data_delayed_123__82_,
  chained_data_delayed_123__81_,chained_data_delayed_123__80_,chained_data_delayed_123__79_,
  chained_data_delayed_123__78_,chained_data_delayed_123__77_,chained_data_delayed_123__76_,
  chained_data_delayed_123__75_,chained_data_delayed_123__74_,
  chained_data_delayed_123__73_,chained_data_delayed_123__72_,chained_data_delayed_123__71_,
  chained_data_delayed_123__70_,chained_data_delayed_123__69_,chained_data_delayed_123__68_,
  chained_data_delayed_123__67_,chained_data_delayed_123__66_,
  chained_data_delayed_123__65_,chained_data_delayed_123__64_,chained_data_delayed_123__63_,
  chained_data_delayed_123__62_,chained_data_delayed_123__61_,chained_data_delayed_123__60_,
  chained_data_delayed_123__59_,chained_data_delayed_123__58_,
  chained_data_delayed_123__57_,chained_data_delayed_123__56_,chained_data_delayed_123__55_,
  chained_data_delayed_123__54_,chained_data_delayed_123__53_,chained_data_delayed_123__52_,
  chained_data_delayed_123__51_,chained_data_delayed_123__50_,
  chained_data_delayed_123__49_,chained_data_delayed_123__48_,chained_data_delayed_123__47_,
  chained_data_delayed_123__46_,chained_data_delayed_123__45_,chained_data_delayed_123__44_,
  chained_data_delayed_123__43_,chained_data_delayed_123__42_,
  chained_data_delayed_123__41_,chained_data_delayed_123__40_,chained_data_delayed_123__39_,
  chained_data_delayed_123__38_,chained_data_delayed_123__37_,chained_data_delayed_123__36_,
  chained_data_delayed_123__35_,chained_data_delayed_123__34_,
  chained_data_delayed_123__33_,chained_data_delayed_123__32_,chained_data_delayed_123__31_,
  chained_data_delayed_123__30_,chained_data_delayed_123__29_,chained_data_delayed_123__28_,
  chained_data_delayed_123__27_,chained_data_delayed_123__26_,
  chained_data_delayed_123__25_,chained_data_delayed_123__24_,chained_data_delayed_123__23_,
  chained_data_delayed_123__22_,chained_data_delayed_123__21_,chained_data_delayed_123__20_,
  chained_data_delayed_123__19_,chained_data_delayed_123__18_,
  chained_data_delayed_123__17_,chained_data_delayed_123__16_,chained_data_delayed_123__15_,
  chained_data_delayed_123__14_,chained_data_delayed_123__13_,chained_data_delayed_123__12_,
  chained_data_delayed_123__11_,chained_data_delayed_123__10_,
  chained_data_delayed_123__9_,chained_data_delayed_123__8_,chained_data_delayed_123__7_,
  chained_data_delayed_123__6_,chained_data_delayed_123__5_,chained_data_delayed_123__4_,
  chained_data_delayed_123__3_,chained_data_delayed_123__2_,chained_data_delayed_123__1_,
  chained_data_delayed_123__0_,chained_data_delayed_122__127_,
  chained_data_delayed_122__126_,chained_data_delayed_122__125_,chained_data_delayed_122__124_,
  chained_data_delayed_122__123_,chained_data_delayed_122__122_,
  chained_data_delayed_122__121_,chained_data_delayed_122__120_,chained_data_delayed_122__119_,
  chained_data_delayed_122__118_,chained_data_delayed_122__117_,chained_data_delayed_122__116_,
  chained_data_delayed_122__115_,chained_data_delayed_122__114_,
  chained_data_delayed_122__113_,chained_data_delayed_122__112_,chained_data_delayed_122__111_,
  chained_data_delayed_122__110_,chained_data_delayed_122__109_,
  chained_data_delayed_122__108_,chained_data_delayed_122__107_,chained_data_delayed_122__106_,
  chained_data_delayed_122__105_,chained_data_delayed_122__104_,
  chained_data_delayed_122__103_,chained_data_delayed_122__102_,chained_data_delayed_122__101_,
  chained_data_delayed_122__100_,chained_data_delayed_122__99_,chained_data_delayed_122__98_,
  chained_data_delayed_122__97_,chained_data_delayed_122__96_,
  chained_data_delayed_122__95_,chained_data_delayed_122__94_,chained_data_delayed_122__93_,
  chained_data_delayed_122__92_,chained_data_delayed_122__91_,chained_data_delayed_122__90_,
  chained_data_delayed_122__89_,chained_data_delayed_122__88_,
  chained_data_delayed_122__87_,chained_data_delayed_122__86_,chained_data_delayed_122__85_,
  chained_data_delayed_122__84_,chained_data_delayed_122__83_,chained_data_delayed_122__82_,
  chained_data_delayed_122__81_,chained_data_delayed_122__80_,
  chained_data_delayed_122__79_,chained_data_delayed_122__78_,chained_data_delayed_122__77_,
  chained_data_delayed_122__76_,chained_data_delayed_122__75_,chained_data_delayed_122__74_,
  chained_data_delayed_122__73_,chained_data_delayed_122__72_,
  chained_data_delayed_122__71_,chained_data_delayed_122__70_,chained_data_delayed_122__69_,
  chained_data_delayed_122__68_,chained_data_delayed_122__67_,chained_data_delayed_122__66_,
  chained_data_delayed_122__65_,chained_data_delayed_122__64_,
  chained_data_delayed_122__63_,chained_data_delayed_122__62_,chained_data_delayed_122__61_,
  chained_data_delayed_122__60_,chained_data_delayed_122__59_,chained_data_delayed_122__58_,
  chained_data_delayed_122__57_,chained_data_delayed_122__56_,
  chained_data_delayed_122__55_,chained_data_delayed_122__54_,chained_data_delayed_122__53_,
  chained_data_delayed_122__52_,chained_data_delayed_122__51_,chained_data_delayed_122__50_,
  chained_data_delayed_122__49_,chained_data_delayed_122__48_,
  chained_data_delayed_122__47_,chained_data_delayed_122__46_,chained_data_delayed_122__45_,
  chained_data_delayed_122__44_,chained_data_delayed_122__43_,chained_data_delayed_122__42_,
  chained_data_delayed_122__41_,chained_data_delayed_122__40_,
  chained_data_delayed_122__39_,chained_data_delayed_122__38_,chained_data_delayed_122__37_,
  chained_data_delayed_122__36_,chained_data_delayed_122__35_,chained_data_delayed_122__34_,
  chained_data_delayed_122__33_,chained_data_delayed_122__32_,
  chained_data_delayed_122__31_,chained_data_delayed_122__30_,chained_data_delayed_122__29_,
  chained_data_delayed_122__28_,chained_data_delayed_122__27_,chained_data_delayed_122__26_,
  chained_data_delayed_122__25_,chained_data_delayed_122__24_,
  chained_data_delayed_122__23_,chained_data_delayed_122__22_,chained_data_delayed_122__21_,
  chained_data_delayed_122__20_,chained_data_delayed_122__19_,chained_data_delayed_122__18_,
  chained_data_delayed_122__17_,chained_data_delayed_122__16_,
  chained_data_delayed_122__15_,chained_data_delayed_122__14_,chained_data_delayed_122__13_,
  chained_data_delayed_122__12_,chained_data_delayed_122__11_,chained_data_delayed_122__10_,
  chained_data_delayed_122__9_,chained_data_delayed_122__8_,
  chained_data_delayed_122__7_,chained_data_delayed_122__6_,chained_data_delayed_122__5_,
  chained_data_delayed_122__4_,chained_data_delayed_122__3_,chained_data_delayed_122__2_,
  chained_data_delayed_122__1_,chained_data_delayed_122__0_,chained_data_delayed_121__127_,
  chained_data_delayed_121__126_,chained_data_delayed_121__125_,
  chained_data_delayed_121__124_,chained_data_delayed_121__123_,chained_data_delayed_121__122_,
  chained_data_delayed_121__121_,chained_data_delayed_121__120_,
  chained_data_delayed_121__119_,chained_data_delayed_121__118_,chained_data_delayed_121__117_,
  chained_data_delayed_121__116_,chained_data_delayed_121__115_,chained_data_delayed_121__114_,
  chained_data_delayed_121__113_,chained_data_delayed_121__112_,
  chained_data_delayed_121__111_,chained_data_delayed_121__110_,chained_data_delayed_121__109_,
  chained_data_delayed_121__108_,chained_data_delayed_121__107_,
  chained_data_delayed_121__106_,chained_data_delayed_121__105_,chained_data_delayed_121__104_,
  chained_data_delayed_121__103_,chained_data_delayed_121__102_,
  chained_data_delayed_121__101_,chained_data_delayed_121__100_,chained_data_delayed_121__99_,
  chained_data_delayed_121__98_,chained_data_delayed_121__97_,chained_data_delayed_121__96_,
  chained_data_delayed_121__95_,chained_data_delayed_121__94_,
  chained_data_delayed_121__93_,chained_data_delayed_121__92_,chained_data_delayed_121__91_,
  chained_data_delayed_121__90_,chained_data_delayed_121__89_,chained_data_delayed_121__88_,
  chained_data_delayed_121__87_,chained_data_delayed_121__86_,
  chained_data_delayed_121__85_,chained_data_delayed_121__84_,chained_data_delayed_121__83_,
  chained_data_delayed_121__82_,chained_data_delayed_121__81_,chained_data_delayed_121__80_,
  chained_data_delayed_121__79_,chained_data_delayed_121__78_,
  chained_data_delayed_121__77_,chained_data_delayed_121__76_,chained_data_delayed_121__75_,
  chained_data_delayed_121__74_,chained_data_delayed_121__73_,chained_data_delayed_121__72_,
  chained_data_delayed_121__71_,chained_data_delayed_121__70_,
  chained_data_delayed_121__69_,chained_data_delayed_121__68_,chained_data_delayed_121__67_,
  chained_data_delayed_121__66_,chained_data_delayed_121__65_,chained_data_delayed_121__64_,
  chained_data_delayed_121__63_,chained_data_delayed_121__62_,
  chained_data_delayed_121__61_,chained_data_delayed_121__60_,chained_data_delayed_121__59_,
  chained_data_delayed_121__58_,chained_data_delayed_121__57_,chained_data_delayed_121__56_,
  chained_data_delayed_121__55_,chained_data_delayed_121__54_,
  chained_data_delayed_121__53_,chained_data_delayed_121__52_,chained_data_delayed_121__51_,
  chained_data_delayed_121__50_,chained_data_delayed_121__49_,chained_data_delayed_121__48_,
  chained_data_delayed_121__47_,chained_data_delayed_121__46_,
  chained_data_delayed_121__45_,chained_data_delayed_121__44_,chained_data_delayed_121__43_,
  chained_data_delayed_121__42_,chained_data_delayed_121__41_,chained_data_delayed_121__40_,
  chained_data_delayed_121__39_,chained_data_delayed_121__38_,
  chained_data_delayed_121__37_,chained_data_delayed_121__36_,chained_data_delayed_121__35_,
  chained_data_delayed_121__34_,chained_data_delayed_121__33_,chained_data_delayed_121__32_,
  chained_data_delayed_121__31_,chained_data_delayed_121__30_,
  chained_data_delayed_121__29_,chained_data_delayed_121__28_,chained_data_delayed_121__27_,
  chained_data_delayed_121__26_,chained_data_delayed_121__25_,chained_data_delayed_121__24_,
  chained_data_delayed_121__23_,chained_data_delayed_121__22_,
  chained_data_delayed_121__21_,chained_data_delayed_121__20_,chained_data_delayed_121__19_,
  chained_data_delayed_121__18_,chained_data_delayed_121__17_,chained_data_delayed_121__16_,
  chained_data_delayed_121__15_,chained_data_delayed_121__14_,
  chained_data_delayed_121__13_,chained_data_delayed_121__12_,chained_data_delayed_121__11_,
  chained_data_delayed_121__10_,chained_data_delayed_121__9_,chained_data_delayed_121__8_,
  chained_data_delayed_121__7_,chained_data_delayed_121__6_,chained_data_delayed_121__5_,
  chained_data_delayed_121__4_,chained_data_delayed_121__3_,
  chained_data_delayed_121__2_,chained_data_delayed_121__1_,chained_data_delayed_121__0_;

  bsg_dff_width_p128
  chained_genblk1_1__ch_reg
  (
    .clk_i(clk_i),
    .data_i(data_i),
    .data_o({ chained_data_delayed_1__127_, chained_data_delayed_1__126_, chained_data_delayed_1__125_, chained_data_delayed_1__124_, chained_data_delayed_1__123_, chained_data_delayed_1__122_, chained_data_delayed_1__121_, chained_data_delayed_1__120_, chained_data_delayed_1__119_, chained_data_delayed_1__118_, chained_data_delayed_1__117_, chained_data_delayed_1__116_, chained_data_delayed_1__115_, chained_data_delayed_1__114_, chained_data_delayed_1__113_, chained_data_delayed_1__112_, chained_data_delayed_1__111_, chained_data_delayed_1__110_, chained_data_delayed_1__109_, chained_data_delayed_1__108_, chained_data_delayed_1__107_, chained_data_delayed_1__106_, chained_data_delayed_1__105_, chained_data_delayed_1__104_, chained_data_delayed_1__103_, chained_data_delayed_1__102_, chained_data_delayed_1__101_, chained_data_delayed_1__100_, chained_data_delayed_1__99_, chained_data_delayed_1__98_, chained_data_delayed_1__97_, chained_data_delayed_1__96_, chained_data_delayed_1__95_, chained_data_delayed_1__94_, chained_data_delayed_1__93_, chained_data_delayed_1__92_, chained_data_delayed_1__91_, chained_data_delayed_1__90_, chained_data_delayed_1__89_, chained_data_delayed_1__88_, chained_data_delayed_1__87_, chained_data_delayed_1__86_, chained_data_delayed_1__85_, chained_data_delayed_1__84_, chained_data_delayed_1__83_, chained_data_delayed_1__82_, chained_data_delayed_1__81_, chained_data_delayed_1__80_, chained_data_delayed_1__79_, chained_data_delayed_1__78_, chained_data_delayed_1__77_, chained_data_delayed_1__76_, chained_data_delayed_1__75_, chained_data_delayed_1__74_, chained_data_delayed_1__73_, chained_data_delayed_1__72_, chained_data_delayed_1__71_, chained_data_delayed_1__70_, chained_data_delayed_1__69_, chained_data_delayed_1__68_, chained_data_delayed_1__67_, chained_data_delayed_1__66_, chained_data_delayed_1__65_, chained_data_delayed_1__64_, chained_data_delayed_1__63_, chained_data_delayed_1__62_, chained_data_delayed_1__61_, chained_data_delayed_1__60_, chained_data_delayed_1__59_, chained_data_delayed_1__58_, chained_data_delayed_1__57_, chained_data_delayed_1__56_, chained_data_delayed_1__55_, chained_data_delayed_1__54_, chained_data_delayed_1__53_, chained_data_delayed_1__52_, chained_data_delayed_1__51_, chained_data_delayed_1__50_, chained_data_delayed_1__49_, chained_data_delayed_1__48_, chained_data_delayed_1__47_, chained_data_delayed_1__46_, chained_data_delayed_1__45_, chained_data_delayed_1__44_, chained_data_delayed_1__43_, chained_data_delayed_1__42_, chained_data_delayed_1__41_, chained_data_delayed_1__40_, chained_data_delayed_1__39_, chained_data_delayed_1__38_, chained_data_delayed_1__37_, chained_data_delayed_1__36_, chained_data_delayed_1__35_, chained_data_delayed_1__34_, chained_data_delayed_1__33_, chained_data_delayed_1__32_, chained_data_delayed_1__31_, chained_data_delayed_1__30_, chained_data_delayed_1__29_, chained_data_delayed_1__28_, chained_data_delayed_1__27_, chained_data_delayed_1__26_, chained_data_delayed_1__25_, chained_data_delayed_1__24_, chained_data_delayed_1__23_, chained_data_delayed_1__22_, chained_data_delayed_1__21_, chained_data_delayed_1__20_, chained_data_delayed_1__19_, chained_data_delayed_1__18_, chained_data_delayed_1__17_, chained_data_delayed_1__16_, chained_data_delayed_1__15_, chained_data_delayed_1__14_, chained_data_delayed_1__13_, chained_data_delayed_1__12_, chained_data_delayed_1__11_, chained_data_delayed_1__10_, chained_data_delayed_1__9_, chained_data_delayed_1__8_, chained_data_delayed_1__7_, chained_data_delayed_1__6_, chained_data_delayed_1__5_, chained_data_delayed_1__4_, chained_data_delayed_1__3_, chained_data_delayed_1__2_, chained_data_delayed_1__1_, chained_data_delayed_1__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_2__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_1__127_, chained_data_delayed_1__126_, chained_data_delayed_1__125_, chained_data_delayed_1__124_, chained_data_delayed_1__123_, chained_data_delayed_1__122_, chained_data_delayed_1__121_, chained_data_delayed_1__120_, chained_data_delayed_1__119_, chained_data_delayed_1__118_, chained_data_delayed_1__117_, chained_data_delayed_1__116_, chained_data_delayed_1__115_, chained_data_delayed_1__114_, chained_data_delayed_1__113_, chained_data_delayed_1__112_, chained_data_delayed_1__111_, chained_data_delayed_1__110_, chained_data_delayed_1__109_, chained_data_delayed_1__108_, chained_data_delayed_1__107_, chained_data_delayed_1__106_, chained_data_delayed_1__105_, chained_data_delayed_1__104_, chained_data_delayed_1__103_, chained_data_delayed_1__102_, chained_data_delayed_1__101_, chained_data_delayed_1__100_, chained_data_delayed_1__99_, chained_data_delayed_1__98_, chained_data_delayed_1__97_, chained_data_delayed_1__96_, chained_data_delayed_1__95_, chained_data_delayed_1__94_, chained_data_delayed_1__93_, chained_data_delayed_1__92_, chained_data_delayed_1__91_, chained_data_delayed_1__90_, chained_data_delayed_1__89_, chained_data_delayed_1__88_, chained_data_delayed_1__87_, chained_data_delayed_1__86_, chained_data_delayed_1__85_, chained_data_delayed_1__84_, chained_data_delayed_1__83_, chained_data_delayed_1__82_, chained_data_delayed_1__81_, chained_data_delayed_1__80_, chained_data_delayed_1__79_, chained_data_delayed_1__78_, chained_data_delayed_1__77_, chained_data_delayed_1__76_, chained_data_delayed_1__75_, chained_data_delayed_1__74_, chained_data_delayed_1__73_, chained_data_delayed_1__72_, chained_data_delayed_1__71_, chained_data_delayed_1__70_, chained_data_delayed_1__69_, chained_data_delayed_1__68_, chained_data_delayed_1__67_, chained_data_delayed_1__66_, chained_data_delayed_1__65_, chained_data_delayed_1__64_, chained_data_delayed_1__63_, chained_data_delayed_1__62_, chained_data_delayed_1__61_, chained_data_delayed_1__60_, chained_data_delayed_1__59_, chained_data_delayed_1__58_, chained_data_delayed_1__57_, chained_data_delayed_1__56_, chained_data_delayed_1__55_, chained_data_delayed_1__54_, chained_data_delayed_1__53_, chained_data_delayed_1__52_, chained_data_delayed_1__51_, chained_data_delayed_1__50_, chained_data_delayed_1__49_, chained_data_delayed_1__48_, chained_data_delayed_1__47_, chained_data_delayed_1__46_, chained_data_delayed_1__45_, chained_data_delayed_1__44_, chained_data_delayed_1__43_, chained_data_delayed_1__42_, chained_data_delayed_1__41_, chained_data_delayed_1__40_, chained_data_delayed_1__39_, chained_data_delayed_1__38_, chained_data_delayed_1__37_, chained_data_delayed_1__36_, chained_data_delayed_1__35_, chained_data_delayed_1__34_, chained_data_delayed_1__33_, chained_data_delayed_1__32_, chained_data_delayed_1__31_, chained_data_delayed_1__30_, chained_data_delayed_1__29_, chained_data_delayed_1__28_, chained_data_delayed_1__27_, chained_data_delayed_1__26_, chained_data_delayed_1__25_, chained_data_delayed_1__24_, chained_data_delayed_1__23_, chained_data_delayed_1__22_, chained_data_delayed_1__21_, chained_data_delayed_1__20_, chained_data_delayed_1__19_, chained_data_delayed_1__18_, chained_data_delayed_1__17_, chained_data_delayed_1__16_, chained_data_delayed_1__15_, chained_data_delayed_1__14_, chained_data_delayed_1__13_, chained_data_delayed_1__12_, chained_data_delayed_1__11_, chained_data_delayed_1__10_, chained_data_delayed_1__9_, chained_data_delayed_1__8_, chained_data_delayed_1__7_, chained_data_delayed_1__6_, chained_data_delayed_1__5_, chained_data_delayed_1__4_, chained_data_delayed_1__3_, chained_data_delayed_1__2_, chained_data_delayed_1__1_, chained_data_delayed_1__0_ }),
    .data_o({ chained_data_delayed_2__127_, chained_data_delayed_2__126_, chained_data_delayed_2__125_, chained_data_delayed_2__124_, chained_data_delayed_2__123_, chained_data_delayed_2__122_, chained_data_delayed_2__121_, chained_data_delayed_2__120_, chained_data_delayed_2__119_, chained_data_delayed_2__118_, chained_data_delayed_2__117_, chained_data_delayed_2__116_, chained_data_delayed_2__115_, chained_data_delayed_2__114_, chained_data_delayed_2__113_, chained_data_delayed_2__112_, chained_data_delayed_2__111_, chained_data_delayed_2__110_, chained_data_delayed_2__109_, chained_data_delayed_2__108_, chained_data_delayed_2__107_, chained_data_delayed_2__106_, chained_data_delayed_2__105_, chained_data_delayed_2__104_, chained_data_delayed_2__103_, chained_data_delayed_2__102_, chained_data_delayed_2__101_, chained_data_delayed_2__100_, chained_data_delayed_2__99_, chained_data_delayed_2__98_, chained_data_delayed_2__97_, chained_data_delayed_2__96_, chained_data_delayed_2__95_, chained_data_delayed_2__94_, chained_data_delayed_2__93_, chained_data_delayed_2__92_, chained_data_delayed_2__91_, chained_data_delayed_2__90_, chained_data_delayed_2__89_, chained_data_delayed_2__88_, chained_data_delayed_2__87_, chained_data_delayed_2__86_, chained_data_delayed_2__85_, chained_data_delayed_2__84_, chained_data_delayed_2__83_, chained_data_delayed_2__82_, chained_data_delayed_2__81_, chained_data_delayed_2__80_, chained_data_delayed_2__79_, chained_data_delayed_2__78_, chained_data_delayed_2__77_, chained_data_delayed_2__76_, chained_data_delayed_2__75_, chained_data_delayed_2__74_, chained_data_delayed_2__73_, chained_data_delayed_2__72_, chained_data_delayed_2__71_, chained_data_delayed_2__70_, chained_data_delayed_2__69_, chained_data_delayed_2__68_, chained_data_delayed_2__67_, chained_data_delayed_2__66_, chained_data_delayed_2__65_, chained_data_delayed_2__64_, chained_data_delayed_2__63_, chained_data_delayed_2__62_, chained_data_delayed_2__61_, chained_data_delayed_2__60_, chained_data_delayed_2__59_, chained_data_delayed_2__58_, chained_data_delayed_2__57_, chained_data_delayed_2__56_, chained_data_delayed_2__55_, chained_data_delayed_2__54_, chained_data_delayed_2__53_, chained_data_delayed_2__52_, chained_data_delayed_2__51_, chained_data_delayed_2__50_, chained_data_delayed_2__49_, chained_data_delayed_2__48_, chained_data_delayed_2__47_, chained_data_delayed_2__46_, chained_data_delayed_2__45_, chained_data_delayed_2__44_, chained_data_delayed_2__43_, chained_data_delayed_2__42_, chained_data_delayed_2__41_, chained_data_delayed_2__40_, chained_data_delayed_2__39_, chained_data_delayed_2__38_, chained_data_delayed_2__37_, chained_data_delayed_2__36_, chained_data_delayed_2__35_, chained_data_delayed_2__34_, chained_data_delayed_2__33_, chained_data_delayed_2__32_, chained_data_delayed_2__31_, chained_data_delayed_2__30_, chained_data_delayed_2__29_, chained_data_delayed_2__28_, chained_data_delayed_2__27_, chained_data_delayed_2__26_, chained_data_delayed_2__25_, chained_data_delayed_2__24_, chained_data_delayed_2__23_, chained_data_delayed_2__22_, chained_data_delayed_2__21_, chained_data_delayed_2__20_, chained_data_delayed_2__19_, chained_data_delayed_2__18_, chained_data_delayed_2__17_, chained_data_delayed_2__16_, chained_data_delayed_2__15_, chained_data_delayed_2__14_, chained_data_delayed_2__13_, chained_data_delayed_2__12_, chained_data_delayed_2__11_, chained_data_delayed_2__10_, chained_data_delayed_2__9_, chained_data_delayed_2__8_, chained_data_delayed_2__7_, chained_data_delayed_2__6_, chained_data_delayed_2__5_, chained_data_delayed_2__4_, chained_data_delayed_2__3_, chained_data_delayed_2__2_, chained_data_delayed_2__1_, chained_data_delayed_2__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_3__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_2__127_, chained_data_delayed_2__126_, chained_data_delayed_2__125_, chained_data_delayed_2__124_, chained_data_delayed_2__123_, chained_data_delayed_2__122_, chained_data_delayed_2__121_, chained_data_delayed_2__120_, chained_data_delayed_2__119_, chained_data_delayed_2__118_, chained_data_delayed_2__117_, chained_data_delayed_2__116_, chained_data_delayed_2__115_, chained_data_delayed_2__114_, chained_data_delayed_2__113_, chained_data_delayed_2__112_, chained_data_delayed_2__111_, chained_data_delayed_2__110_, chained_data_delayed_2__109_, chained_data_delayed_2__108_, chained_data_delayed_2__107_, chained_data_delayed_2__106_, chained_data_delayed_2__105_, chained_data_delayed_2__104_, chained_data_delayed_2__103_, chained_data_delayed_2__102_, chained_data_delayed_2__101_, chained_data_delayed_2__100_, chained_data_delayed_2__99_, chained_data_delayed_2__98_, chained_data_delayed_2__97_, chained_data_delayed_2__96_, chained_data_delayed_2__95_, chained_data_delayed_2__94_, chained_data_delayed_2__93_, chained_data_delayed_2__92_, chained_data_delayed_2__91_, chained_data_delayed_2__90_, chained_data_delayed_2__89_, chained_data_delayed_2__88_, chained_data_delayed_2__87_, chained_data_delayed_2__86_, chained_data_delayed_2__85_, chained_data_delayed_2__84_, chained_data_delayed_2__83_, chained_data_delayed_2__82_, chained_data_delayed_2__81_, chained_data_delayed_2__80_, chained_data_delayed_2__79_, chained_data_delayed_2__78_, chained_data_delayed_2__77_, chained_data_delayed_2__76_, chained_data_delayed_2__75_, chained_data_delayed_2__74_, chained_data_delayed_2__73_, chained_data_delayed_2__72_, chained_data_delayed_2__71_, chained_data_delayed_2__70_, chained_data_delayed_2__69_, chained_data_delayed_2__68_, chained_data_delayed_2__67_, chained_data_delayed_2__66_, chained_data_delayed_2__65_, chained_data_delayed_2__64_, chained_data_delayed_2__63_, chained_data_delayed_2__62_, chained_data_delayed_2__61_, chained_data_delayed_2__60_, chained_data_delayed_2__59_, chained_data_delayed_2__58_, chained_data_delayed_2__57_, chained_data_delayed_2__56_, chained_data_delayed_2__55_, chained_data_delayed_2__54_, chained_data_delayed_2__53_, chained_data_delayed_2__52_, chained_data_delayed_2__51_, chained_data_delayed_2__50_, chained_data_delayed_2__49_, chained_data_delayed_2__48_, chained_data_delayed_2__47_, chained_data_delayed_2__46_, chained_data_delayed_2__45_, chained_data_delayed_2__44_, chained_data_delayed_2__43_, chained_data_delayed_2__42_, chained_data_delayed_2__41_, chained_data_delayed_2__40_, chained_data_delayed_2__39_, chained_data_delayed_2__38_, chained_data_delayed_2__37_, chained_data_delayed_2__36_, chained_data_delayed_2__35_, chained_data_delayed_2__34_, chained_data_delayed_2__33_, chained_data_delayed_2__32_, chained_data_delayed_2__31_, chained_data_delayed_2__30_, chained_data_delayed_2__29_, chained_data_delayed_2__28_, chained_data_delayed_2__27_, chained_data_delayed_2__26_, chained_data_delayed_2__25_, chained_data_delayed_2__24_, chained_data_delayed_2__23_, chained_data_delayed_2__22_, chained_data_delayed_2__21_, chained_data_delayed_2__20_, chained_data_delayed_2__19_, chained_data_delayed_2__18_, chained_data_delayed_2__17_, chained_data_delayed_2__16_, chained_data_delayed_2__15_, chained_data_delayed_2__14_, chained_data_delayed_2__13_, chained_data_delayed_2__12_, chained_data_delayed_2__11_, chained_data_delayed_2__10_, chained_data_delayed_2__9_, chained_data_delayed_2__8_, chained_data_delayed_2__7_, chained_data_delayed_2__6_, chained_data_delayed_2__5_, chained_data_delayed_2__4_, chained_data_delayed_2__3_, chained_data_delayed_2__2_, chained_data_delayed_2__1_, chained_data_delayed_2__0_ }),
    .data_o({ chained_data_delayed_3__127_, chained_data_delayed_3__126_, chained_data_delayed_3__125_, chained_data_delayed_3__124_, chained_data_delayed_3__123_, chained_data_delayed_3__122_, chained_data_delayed_3__121_, chained_data_delayed_3__120_, chained_data_delayed_3__119_, chained_data_delayed_3__118_, chained_data_delayed_3__117_, chained_data_delayed_3__116_, chained_data_delayed_3__115_, chained_data_delayed_3__114_, chained_data_delayed_3__113_, chained_data_delayed_3__112_, chained_data_delayed_3__111_, chained_data_delayed_3__110_, chained_data_delayed_3__109_, chained_data_delayed_3__108_, chained_data_delayed_3__107_, chained_data_delayed_3__106_, chained_data_delayed_3__105_, chained_data_delayed_3__104_, chained_data_delayed_3__103_, chained_data_delayed_3__102_, chained_data_delayed_3__101_, chained_data_delayed_3__100_, chained_data_delayed_3__99_, chained_data_delayed_3__98_, chained_data_delayed_3__97_, chained_data_delayed_3__96_, chained_data_delayed_3__95_, chained_data_delayed_3__94_, chained_data_delayed_3__93_, chained_data_delayed_3__92_, chained_data_delayed_3__91_, chained_data_delayed_3__90_, chained_data_delayed_3__89_, chained_data_delayed_3__88_, chained_data_delayed_3__87_, chained_data_delayed_3__86_, chained_data_delayed_3__85_, chained_data_delayed_3__84_, chained_data_delayed_3__83_, chained_data_delayed_3__82_, chained_data_delayed_3__81_, chained_data_delayed_3__80_, chained_data_delayed_3__79_, chained_data_delayed_3__78_, chained_data_delayed_3__77_, chained_data_delayed_3__76_, chained_data_delayed_3__75_, chained_data_delayed_3__74_, chained_data_delayed_3__73_, chained_data_delayed_3__72_, chained_data_delayed_3__71_, chained_data_delayed_3__70_, chained_data_delayed_3__69_, chained_data_delayed_3__68_, chained_data_delayed_3__67_, chained_data_delayed_3__66_, chained_data_delayed_3__65_, chained_data_delayed_3__64_, chained_data_delayed_3__63_, chained_data_delayed_3__62_, chained_data_delayed_3__61_, chained_data_delayed_3__60_, chained_data_delayed_3__59_, chained_data_delayed_3__58_, chained_data_delayed_3__57_, chained_data_delayed_3__56_, chained_data_delayed_3__55_, chained_data_delayed_3__54_, chained_data_delayed_3__53_, chained_data_delayed_3__52_, chained_data_delayed_3__51_, chained_data_delayed_3__50_, chained_data_delayed_3__49_, chained_data_delayed_3__48_, chained_data_delayed_3__47_, chained_data_delayed_3__46_, chained_data_delayed_3__45_, chained_data_delayed_3__44_, chained_data_delayed_3__43_, chained_data_delayed_3__42_, chained_data_delayed_3__41_, chained_data_delayed_3__40_, chained_data_delayed_3__39_, chained_data_delayed_3__38_, chained_data_delayed_3__37_, chained_data_delayed_3__36_, chained_data_delayed_3__35_, chained_data_delayed_3__34_, chained_data_delayed_3__33_, chained_data_delayed_3__32_, chained_data_delayed_3__31_, chained_data_delayed_3__30_, chained_data_delayed_3__29_, chained_data_delayed_3__28_, chained_data_delayed_3__27_, chained_data_delayed_3__26_, chained_data_delayed_3__25_, chained_data_delayed_3__24_, chained_data_delayed_3__23_, chained_data_delayed_3__22_, chained_data_delayed_3__21_, chained_data_delayed_3__20_, chained_data_delayed_3__19_, chained_data_delayed_3__18_, chained_data_delayed_3__17_, chained_data_delayed_3__16_, chained_data_delayed_3__15_, chained_data_delayed_3__14_, chained_data_delayed_3__13_, chained_data_delayed_3__12_, chained_data_delayed_3__11_, chained_data_delayed_3__10_, chained_data_delayed_3__9_, chained_data_delayed_3__8_, chained_data_delayed_3__7_, chained_data_delayed_3__6_, chained_data_delayed_3__5_, chained_data_delayed_3__4_, chained_data_delayed_3__3_, chained_data_delayed_3__2_, chained_data_delayed_3__1_, chained_data_delayed_3__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_4__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_3__127_, chained_data_delayed_3__126_, chained_data_delayed_3__125_, chained_data_delayed_3__124_, chained_data_delayed_3__123_, chained_data_delayed_3__122_, chained_data_delayed_3__121_, chained_data_delayed_3__120_, chained_data_delayed_3__119_, chained_data_delayed_3__118_, chained_data_delayed_3__117_, chained_data_delayed_3__116_, chained_data_delayed_3__115_, chained_data_delayed_3__114_, chained_data_delayed_3__113_, chained_data_delayed_3__112_, chained_data_delayed_3__111_, chained_data_delayed_3__110_, chained_data_delayed_3__109_, chained_data_delayed_3__108_, chained_data_delayed_3__107_, chained_data_delayed_3__106_, chained_data_delayed_3__105_, chained_data_delayed_3__104_, chained_data_delayed_3__103_, chained_data_delayed_3__102_, chained_data_delayed_3__101_, chained_data_delayed_3__100_, chained_data_delayed_3__99_, chained_data_delayed_3__98_, chained_data_delayed_3__97_, chained_data_delayed_3__96_, chained_data_delayed_3__95_, chained_data_delayed_3__94_, chained_data_delayed_3__93_, chained_data_delayed_3__92_, chained_data_delayed_3__91_, chained_data_delayed_3__90_, chained_data_delayed_3__89_, chained_data_delayed_3__88_, chained_data_delayed_3__87_, chained_data_delayed_3__86_, chained_data_delayed_3__85_, chained_data_delayed_3__84_, chained_data_delayed_3__83_, chained_data_delayed_3__82_, chained_data_delayed_3__81_, chained_data_delayed_3__80_, chained_data_delayed_3__79_, chained_data_delayed_3__78_, chained_data_delayed_3__77_, chained_data_delayed_3__76_, chained_data_delayed_3__75_, chained_data_delayed_3__74_, chained_data_delayed_3__73_, chained_data_delayed_3__72_, chained_data_delayed_3__71_, chained_data_delayed_3__70_, chained_data_delayed_3__69_, chained_data_delayed_3__68_, chained_data_delayed_3__67_, chained_data_delayed_3__66_, chained_data_delayed_3__65_, chained_data_delayed_3__64_, chained_data_delayed_3__63_, chained_data_delayed_3__62_, chained_data_delayed_3__61_, chained_data_delayed_3__60_, chained_data_delayed_3__59_, chained_data_delayed_3__58_, chained_data_delayed_3__57_, chained_data_delayed_3__56_, chained_data_delayed_3__55_, chained_data_delayed_3__54_, chained_data_delayed_3__53_, chained_data_delayed_3__52_, chained_data_delayed_3__51_, chained_data_delayed_3__50_, chained_data_delayed_3__49_, chained_data_delayed_3__48_, chained_data_delayed_3__47_, chained_data_delayed_3__46_, chained_data_delayed_3__45_, chained_data_delayed_3__44_, chained_data_delayed_3__43_, chained_data_delayed_3__42_, chained_data_delayed_3__41_, chained_data_delayed_3__40_, chained_data_delayed_3__39_, chained_data_delayed_3__38_, chained_data_delayed_3__37_, chained_data_delayed_3__36_, chained_data_delayed_3__35_, chained_data_delayed_3__34_, chained_data_delayed_3__33_, chained_data_delayed_3__32_, chained_data_delayed_3__31_, chained_data_delayed_3__30_, chained_data_delayed_3__29_, chained_data_delayed_3__28_, chained_data_delayed_3__27_, chained_data_delayed_3__26_, chained_data_delayed_3__25_, chained_data_delayed_3__24_, chained_data_delayed_3__23_, chained_data_delayed_3__22_, chained_data_delayed_3__21_, chained_data_delayed_3__20_, chained_data_delayed_3__19_, chained_data_delayed_3__18_, chained_data_delayed_3__17_, chained_data_delayed_3__16_, chained_data_delayed_3__15_, chained_data_delayed_3__14_, chained_data_delayed_3__13_, chained_data_delayed_3__12_, chained_data_delayed_3__11_, chained_data_delayed_3__10_, chained_data_delayed_3__9_, chained_data_delayed_3__8_, chained_data_delayed_3__7_, chained_data_delayed_3__6_, chained_data_delayed_3__5_, chained_data_delayed_3__4_, chained_data_delayed_3__3_, chained_data_delayed_3__2_, chained_data_delayed_3__1_, chained_data_delayed_3__0_ }),
    .data_o({ chained_data_delayed_4__127_, chained_data_delayed_4__126_, chained_data_delayed_4__125_, chained_data_delayed_4__124_, chained_data_delayed_4__123_, chained_data_delayed_4__122_, chained_data_delayed_4__121_, chained_data_delayed_4__120_, chained_data_delayed_4__119_, chained_data_delayed_4__118_, chained_data_delayed_4__117_, chained_data_delayed_4__116_, chained_data_delayed_4__115_, chained_data_delayed_4__114_, chained_data_delayed_4__113_, chained_data_delayed_4__112_, chained_data_delayed_4__111_, chained_data_delayed_4__110_, chained_data_delayed_4__109_, chained_data_delayed_4__108_, chained_data_delayed_4__107_, chained_data_delayed_4__106_, chained_data_delayed_4__105_, chained_data_delayed_4__104_, chained_data_delayed_4__103_, chained_data_delayed_4__102_, chained_data_delayed_4__101_, chained_data_delayed_4__100_, chained_data_delayed_4__99_, chained_data_delayed_4__98_, chained_data_delayed_4__97_, chained_data_delayed_4__96_, chained_data_delayed_4__95_, chained_data_delayed_4__94_, chained_data_delayed_4__93_, chained_data_delayed_4__92_, chained_data_delayed_4__91_, chained_data_delayed_4__90_, chained_data_delayed_4__89_, chained_data_delayed_4__88_, chained_data_delayed_4__87_, chained_data_delayed_4__86_, chained_data_delayed_4__85_, chained_data_delayed_4__84_, chained_data_delayed_4__83_, chained_data_delayed_4__82_, chained_data_delayed_4__81_, chained_data_delayed_4__80_, chained_data_delayed_4__79_, chained_data_delayed_4__78_, chained_data_delayed_4__77_, chained_data_delayed_4__76_, chained_data_delayed_4__75_, chained_data_delayed_4__74_, chained_data_delayed_4__73_, chained_data_delayed_4__72_, chained_data_delayed_4__71_, chained_data_delayed_4__70_, chained_data_delayed_4__69_, chained_data_delayed_4__68_, chained_data_delayed_4__67_, chained_data_delayed_4__66_, chained_data_delayed_4__65_, chained_data_delayed_4__64_, chained_data_delayed_4__63_, chained_data_delayed_4__62_, chained_data_delayed_4__61_, chained_data_delayed_4__60_, chained_data_delayed_4__59_, chained_data_delayed_4__58_, chained_data_delayed_4__57_, chained_data_delayed_4__56_, chained_data_delayed_4__55_, chained_data_delayed_4__54_, chained_data_delayed_4__53_, chained_data_delayed_4__52_, chained_data_delayed_4__51_, chained_data_delayed_4__50_, chained_data_delayed_4__49_, chained_data_delayed_4__48_, chained_data_delayed_4__47_, chained_data_delayed_4__46_, chained_data_delayed_4__45_, chained_data_delayed_4__44_, chained_data_delayed_4__43_, chained_data_delayed_4__42_, chained_data_delayed_4__41_, chained_data_delayed_4__40_, chained_data_delayed_4__39_, chained_data_delayed_4__38_, chained_data_delayed_4__37_, chained_data_delayed_4__36_, chained_data_delayed_4__35_, chained_data_delayed_4__34_, chained_data_delayed_4__33_, chained_data_delayed_4__32_, chained_data_delayed_4__31_, chained_data_delayed_4__30_, chained_data_delayed_4__29_, chained_data_delayed_4__28_, chained_data_delayed_4__27_, chained_data_delayed_4__26_, chained_data_delayed_4__25_, chained_data_delayed_4__24_, chained_data_delayed_4__23_, chained_data_delayed_4__22_, chained_data_delayed_4__21_, chained_data_delayed_4__20_, chained_data_delayed_4__19_, chained_data_delayed_4__18_, chained_data_delayed_4__17_, chained_data_delayed_4__16_, chained_data_delayed_4__15_, chained_data_delayed_4__14_, chained_data_delayed_4__13_, chained_data_delayed_4__12_, chained_data_delayed_4__11_, chained_data_delayed_4__10_, chained_data_delayed_4__9_, chained_data_delayed_4__8_, chained_data_delayed_4__7_, chained_data_delayed_4__6_, chained_data_delayed_4__5_, chained_data_delayed_4__4_, chained_data_delayed_4__3_, chained_data_delayed_4__2_, chained_data_delayed_4__1_, chained_data_delayed_4__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_5__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_4__127_, chained_data_delayed_4__126_, chained_data_delayed_4__125_, chained_data_delayed_4__124_, chained_data_delayed_4__123_, chained_data_delayed_4__122_, chained_data_delayed_4__121_, chained_data_delayed_4__120_, chained_data_delayed_4__119_, chained_data_delayed_4__118_, chained_data_delayed_4__117_, chained_data_delayed_4__116_, chained_data_delayed_4__115_, chained_data_delayed_4__114_, chained_data_delayed_4__113_, chained_data_delayed_4__112_, chained_data_delayed_4__111_, chained_data_delayed_4__110_, chained_data_delayed_4__109_, chained_data_delayed_4__108_, chained_data_delayed_4__107_, chained_data_delayed_4__106_, chained_data_delayed_4__105_, chained_data_delayed_4__104_, chained_data_delayed_4__103_, chained_data_delayed_4__102_, chained_data_delayed_4__101_, chained_data_delayed_4__100_, chained_data_delayed_4__99_, chained_data_delayed_4__98_, chained_data_delayed_4__97_, chained_data_delayed_4__96_, chained_data_delayed_4__95_, chained_data_delayed_4__94_, chained_data_delayed_4__93_, chained_data_delayed_4__92_, chained_data_delayed_4__91_, chained_data_delayed_4__90_, chained_data_delayed_4__89_, chained_data_delayed_4__88_, chained_data_delayed_4__87_, chained_data_delayed_4__86_, chained_data_delayed_4__85_, chained_data_delayed_4__84_, chained_data_delayed_4__83_, chained_data_delayed_4__82_, chained_data_delayed_4__81_, chained_data_delayed_4__80_, chained_data_delayed_4__79_, chained_data_delayed_4__78_, chained_data_delayed_4__77_, chained_data_delayed_4__76_, chained_data_delayed_4__75_, chained_data_delayed_4__74_, chained_data_delayed_4__73_, chained_data_delayed_4__72_, chained_data_delayed_4__71_, chained_data_delayed_4__70_, chained_data_delayed_4__69_, chained_data_delayed_4__68_, chained_data_delayed_4__67_, chained_data_delayed_4__66_, chained_data_delayed_4__65_, chained_data_delayed_4__64_, chained_data_delayed_4__63_, chained_data_delayed_4__62_, chained_data_delayed_4__61_, chained_data_delayed_4__60_, chained_data_delayed_4__59_, chained_data_delayed_4__58_, chained_data_delayed_4__57_, chained_data_delayed_4__56_, chained_data_delayed_4__55_, chained_data_delayed_4__54_, chained_data_delayed_4__53_, chained_data_delayed_4__52_, chained_data_delayed_4__51_, chained_data_delayed_4__50_, chained_data_delayed_4__49_, chained_data_delayed_4__48_, chained_data_delayed_4__47_, chained_data_delayed_4__46_, chained_data_delayed_4__45_, chained_data_delayed_4__44_, chained_data_delayed_4__43_, chained_data_delayed_4__42_, chained_data_delayed_4__41_, chained_data_delayed_4__40_, chained_data_delayed_4__39_, chained_data_delayed_4__38_, chained_data_delayed_4__37_, chained_data_delayed_4__36_, chained_data_delayed_4__35_, chained_data_delayed_4__34_, chained_data_delayed_4__33_, chained_data_delayed_4__32_, chained_data_delayed_4__31_, chained_data_delayed_4__30_, chained_data_delayed_4__29_, chained_data_delayed_4__28_, chained_data_delayed_4__27_, chained_data_delayed_4__26_, chained_data_delayed_4__25_, chained_data_delayed_4__24_, chained_data_delayed_4__23_, chained_data_delayed_4__22_, chained_data_delayed_4__21_, chained_data_delayed_4__20_, chained_data_delayed_4__19_, chained_data_delayed_4__18_, chained_data_delayed_4__17_, chained_data_delayed_4__16_, chained_data_delayed_4__15_, chained_data_delayed_4__14_, chained_data_delayed_4__13_, chained_data_delayed_4__12_, chained_data_delayed_4__11_, chained_data_delayed_4__10_, chained_data_delayed_4__9_, chained_data_delayed_4__8_, chained_data_delayed_4__7_, chained_data_delayed_4__6_, chained_data_delayed_4__5_, chained_data_delayed_4__4_, chained_data_delayed_4__3_, chained_data_delayed_4__2_, chained_data_delayed_4__1_, chained_data_delayed_4__0_ }),
    .data_o({ chained_data_delayed_5__127_, chained_data_delayed_5__126_, chained_data_delayed_5__125_, chained_data_delayed_5__124_, chained_data_delayed_5__123_, chained_data_delayed_5__122_, chained_data_delayed_5__121_, chained_data_delayed_5__120_, chained_data_delayed_5__119_, chained_data_delayed_5__118_, chained_data_delayed_5__117_, chained_data_delayed_5__116_, chained_data_delayed_5__115_, chained_data_delayed_5__114_, chained_data_delayed_5__113_, chained_data_delayed_5__112_, chained_data_delayed_5__111_, chained_data_delayed_5__110_, chained_data_delayed_5__109_, chained_data_delayed_5__108_, chained_data_delayed_5__107_, chained_data_delayed_5__106_, chained_data_delayed_5__105_, chained_data_delayed_5__104_, chained_data_delayed_5__103_, chained_data_delayed_5__102_, chained_data_delayed_5__101_, chained_data_delayed_5__100_, chained_data_delayed_5__99_, chained_data_delayed_5__98_, chained_data_delayed_5__97_, chained_data_delayed_5__96_, chained_data_delayed_5__95_, chained_data_delayed_5__94_, chained_data_delayed_5__93_, chained_data_delayed_5__92_, chained_data_delayed_5__91_, chained_data_delayed_5__90_, chained_data_delayed_5__89_, chained_data_delayed_5__88_, chained_data_delayed_5__87_, chained_data_delayed_5__86_, chained_data_delayed_5__85_, chained_data_delayed_5__84_, chained_data_delayed_5__83_, chained_data_delayed_5__82_, chained_data_delayed_5__81_, chained_data_delayed_5__80_, chained_data_delayed_5__79_, chained_data_delayed_5__78_, chained_data_delayed_5__77_, chained_data_delayed_5__76_, chained_data_delayed_5__75_, chained_data_delayed_5__74_, chained_data_delayed_5__73_, chained_data_delayed_5__72_, chained_data_delayed_5__71_, chained_data_delayed_5__70_, chained_data_delayed_5__69_, chained_data_delayed_5__68_, chained_data_delayed_5__67_, chained_data_delayed_5__66_, chained_data_delayed_5__65_, chained_data_delayed_5__64_, chained_data_delayed_5__63_, chained_data_delayed_5__62_, chained_data_delayed_5__61_, chained_data_delayed_5__60_, chained_data_delayed_5__59_, chained_data_delayed_5__58_, chained_data_delayed_5__57_, chained_data_delayed_5__56_, chained_data_delayed_5__55_, chained_data_delayed_5__54_, chained_data_delayed_5__53_, chained_data_delayed_5__52_, chained_data_delayed_5__51_, chained_data_delayed_5__50_, chained_data_delayed_5__49_, chained_data_delayed_5__48_, chained_data_delayed_5__47_, chained_data_delayed_5__46_, chained_data_delayed_5__45_, chained_data_delayed_5__44_, chained_data_delayed_5__43_, chained_data_delayed_5__42_, chained_data_delayed_5__41_, chained_data_delayed_5__40_, chained_data_delayed_5__39_, chained_data_delayed_5__38_, chained_data_delayed_5__37_, chained_data_delayed_5__36_, chained_data_delayed_5__35_, chained_data_delayed_5__34_, chained_data_delayed_5__33_, chained_data_delayed_5__32_, chained_data_delayed_5__31_, chained_data_delayed_5__30_, chained_data_delayed_5__29_, chained_data_delayed_5__28_, chained_data_delayed_5__27_, chained_data_delayed_5__26_, chained_data_delayed_5__25_, chained_data_delayed_5__24_, chained_data_delayed_5__23_, chained_data_delayed_5__22_, chained_data_delayed_5__21_, chained_data_delayed_5__20_, chained_data_delayed_5__19_, chained_data_delayed_5__18_, chained_data_delayed_5__17_, chained_data_delayed_5__16_, chained_data_delayed_5__15_, chained_data_delayed_5__14_, chained_data_delayed_5__13_, chained_data_delayed_5__12_, chained_data_delayed_5__11_, chained_data_delayed_5__10_, chained_data_delayed_5__9_, chained_data_delayed_5__8_, chained_data_delayed_5__7_, chained_data_delayed_5__6_, chained_data_delayed_5__5_, chained_data_delayed_5__4_, chained_data_delayed_5__3_, chained_data_delayed_5__2_, chained_data_delayed_5__1_, chained_data_delayed_5__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_6__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_5__127_, chained_data_delayed_5__126_, chained_data_delayed_5__125_, chained_data_delayed_5__124_, chained_data_delayed_5__123_, chained_data_delayed_5__122_, chained_data_delayed_5__121_, chained_data_delayed_5__120_, chained_data_delayed_5__119_, chained_data_delayed_5__118_, chained_data_delayed_5__117_, chained_data_delayed_5__116_, chained_data_delayed_5__115_, chained_data_delayed_5__114_, chained_data_delayed_5__113_, chained_data_delayed_5__112_, chained_data_delayed_5__111_, chained_data_delayed_5__110_, chained_data_delayed_5__109_, chained_data_delayed_5__108_, chained_data_delayed_5__107_, chained_data_delayed_5__106_, chained_data_delayed_5__105_, chained_data_delayed_5__104_, chained_data_delayed_5__103_, chained_data_delayed_5__102_, chained_data_delayed_5__101_, chained_data_delayed_5__100_, chained_data_delayed_5__99_, chained_data_delayed_5__98_, chained_data_delayed_5__97_, chained_data_delayed_5__96_, chained_data_delayed_5__95_, chained_data_delayed_5__94_, chained_data_delayed_5__93_, chained_data_delayed_5__92_, chained_data_delayed_5__91_, chained_data_delayed_5__90_, chained_data_delayed_5__89_, chained_data_delayed_5__88_, chained_data_delayed_5__87_, chained_data_delayed_5__86_, chained_data_delayed_5__85_, chained_data_delayed_5__84_, chained_data_delayed_5__83_, chained_data_delayed_5__82_, chained_data_delayed_5__81_, chained_data_delayed_5__80_, chained_data_delayed_5__79_, chained_data_delayed_5__78_, chained_data_delayed_5__77_, chained_data_delayed_5__76_, chained_data_delayed_5__75_, chained_data_delayed_5__74_, chained_data_delayed_5__73_, chained_data_delayed_5__72_, chained_data_delayed_5__71_, chained_data_delayed_5__70_, chained_data_delayed_5__69_, chained_data_delayed_5__68_, chained_data_delayed_5__67_, chained_data_delayed_5__66_, chained_data_delayed_5__65_, chained_data_delayed_5__64_, chained_data_delayed_5__63_, chained_data_delayed_5__62_, chained_data_delayed_5__61_, chained_data_delayed_5__60_, chained_data_delayed_5__59_, chained_data_delayed_5__58_, chained_data_delayed_5__57_, chained_data_delayed_5__56_, chained_data_delayed_5__55_, chained_data_delayed_5__54_, chained_data_delayed_5__53_, chained_data_delayed_5__52_, chained_data_delayed_5__51_, chained_data_delayed_5__50_, chained_data_delayed_5__49_, chained_data_delayed_5__48_, chained_data_delayed_5__47_, chained_data_delayed_5__46_, chained_data_delayed_5__45_, chained_data_delayed_5__44_, chained_data_delayed_5__43_, chained_data_delayed_5__42_, chained_data_delayed_5__41_, chained_data_delayed_5__40_, chained_data_delayed_5__39_, chained_data_delayed_5__38_, chained_data_delayed_5__37_, chained_data_delayed_5__36_, chained_data_delayed_5__35_, chained_data_delayed_5__34_, chained_data_delayed_5__33_, chained_data_delayed_5__32_, chained_data_delayed_5__31_, chained_data_delayed_5__30_, chained_data_delayed_5__29_, chained_data_delayed_5__28_, chained_data_delayed_5__27_, chained_data_delayed_5__26_, chained_data_delayed_5__25_, chained_data_delayed_5__24_, chained_data_delayed_5__23_, chained_data_delayed_5__22_, chained_data_delayed_5__21_, chained_data_delayed_5__20_, chained_data_delayed_5__19_, chained_data_delayed_5__18_, chained_data_delayed_5__17_, chained_data_delayed_5__16_, chained_data_delayed_5__15_, chained_data_delayed_5__14_, chained_data_delayed_5__13_, chained_data_delayed_5__12_, chained_data_delayed_5__11_, chained_data_delayed_5__10_, chained_data_delayed_5__9_, chained_data_delayed_5__8_, chained_data_delayed_5__7_, chained_data_delayed_5__6_, chained_data_delayed_5__5_, chained_data_delayed_5__4_, chained_data_delayed_5__3_, chained_data_delayed_5__2_, chained_data_delayed_5__1_, chained_data_delayed_5__0_ }),
    .data_o({ chained_data_delayed_6__127_, chained_data_delayed_6__126_, chained_data_delayed_6__125_, chained_data_delayed_6__124_, chained_data_delayed_6__123_, chained_data_delayed_6__122_, chained_data_delayed_6__121_, chained_data_delayed_6__120_, chained_data_delayed_6__119_, chained_data_delayed_6__118_, chained_data_delayed_6__117_, chained_data_delayed_6__116_, chained_data_delayed_6__115_, chained_data_delayed_6__114_, chained_data_delayed_6__113_, chained_data_delayed_6__112_, chained_data_delayed_6__111_, chained_data_delayed_6__110_, chained_data_delayed_6__109_, chained_data_delayed_6__108_, chained_data_delayed_6__107_, chained_data_delayed_6__106_, chained_data_delayed_6__105_, chained_data_delayed_6__104_, chained_data_delayed_6__103_, chained_data_delayed_6__102_, chained_data_delayed_6__101_, chained_data_delayed_6__100_, chained_data_delayed_6__99_, chained_data_delayed_6__98_, chained_data_delayed_6__97_, chained_data_delayed_6__96_, chained_data_delayed_6__95_, chained_data_delayed_6__94_, chained_data_delayed_6__93_, chained_data_delayed_6__92_, chained_data_delayed_6__91_, chained_data_delayed_6__90_, chained_data_delayed_6__89_, chained_data_delayed_6__88_, chained_data_delayed_6__87_, chained_data_delayed_6__86_, chained_data_delayed_6__85_, chained_data_delayed_6__84_, chained_data_delayed_6__83_, chained_data_delayed_6__82_, chained_data_delayed_6__81_, chained_data_delayed_6__80_, chained_data_delayed_6__79_, chained_data_delayed_6__78_, chained_data_delayed_6__77_, chained_data_delayed_6__76_, chained_data_delayed_6__75_, chained_data_delayed_6__74_, chained_data_delayed_6__73_, chained_data_delayed_6__72_, chained_data_delayed_6__71_, chained_data_delayed_6__70_, chained_data_delayed_6__69_, chained_data_delayed_6__68_, chained_data_delayed_6__67_, chained_data_delayed_6__66_, chained_data_delayed_6__65_, chained_data_delayed_6__64_, chained_data_delayed_6__63_, chained_data_delayed_6__62_, chained_data_delayed_6__61_, chained_data_delayed_6__60_, chained_data_delayed_6__59_, chained_data_delayed_6__58_, chained_data_delayed_6__57_, chained_data_delayed_6__56_, chained_data_delayed_6__55_, chained_data_delayed_6__54_, chained_data_delayed_6__53_, chained_data_delayed_6__52_, chained_data_delayed_6__51_, chained_data_delayed_6__50_, chained_data_delayed_6__49_, chained_data_delayed_6__48_, chained_data_delayed_6__47_, chained_data_delayed_6__46_, chained_data_delayed_6__45_, chained_data_delayed_6__44_, chained_data_delayed_6__43_, chained_data_delayed_6__42_, chained_data_delayed_6__41_, chained_data_delayed_6__40_, chained_data_delayed_6__39_, chained_data_delayed_6__38_, chained_data_delayed_6__37_, chained_data_delayed_6__36_, chained_data_delayed_6__35_, chained_data_delayed_6__34_, chained_data_delayed_6__33_, chained_data_delayed_6__32_, chained_data_delayed_6__31_, chained_data_delayed_6__30_, chained_data_delayed_6__29_, chained_data_delayed_6__28_, chained_data_delayed_6__27_, chained_data_delayed_6__26_, chained_data_delayed_6__25_, chained_data_delayed_6__24_, chained_data_delayed_6__23_, chained_data_delayed_6__22_, chained_data_delayed_6__21_, chained_data_delayed_6__20_, chained_data_delayed_6__19_, chained_data_delayed_6__18_, chained_data_delayed_6__17_, chained_data_delayed_6__16_, chained_data_delayed_6__15_, chained_data_delayed_6__14_, chained_data_delayed_6__13_, chained_data_delayed_6__12_, chained_data_delayed_6__11_, chained_data_delayed_6__10_, chained_data_delayed_6__9_, chained_data_delayed_6__8_, chained_data_delayed_6__7_, chained_data_delayed_6__6_, chained_data_delayed_6__5_, chained_data_delayed_6__4_, chained_data_delayed_6__3_, chained_data_delayed_6__2_, chained_data_delayed_6__1_, chained_data_delayed_6__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_7__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_6__127_, chained_data_delayed_6__126_, chained_data_delayed_6__125_, chained_data_delayed_6__124_, chained_data_delayed_6__123_, chained_data_delayed_6__122_, chained_data_delayed_6__121_, chained_data_delayed_6__120_, chained_data_delayed_6__119_, chained_data_delayed_6__118_, chained_data_delayed_6__117_, chained_data_delayed_6__116_, chained_data_delayed_6__115_, chained_data_delayed_6__114_, chained_data_delayed_6__113_, chained_data_delayed_6__112_, chained_data_delayed_6__111_, chained_data_delayed_6__110_, chained_data_delayed_6__109_, chained_data_delayed_6__108_, chained_data_delayed_6__107_, chained_data_delayed_6__106_, chained_data_delayed_6__105_, chained_data_delayed_6__104_, chained_data_delayed_6__103_, chained_data_delayed_6__102_, chained_data_delayed_6__101_, chained_data_delayed_6__100_, chained_data_delayed_6__99_, chained_data_delayed_6__98_, chained_data_delayed_6__97_, chained_data_delayed_6__96_, chained_data_delayed_6__95_, chained_data_delayed_6__94_, chained_data_delayed_6__93_, chained_data_delayed_6__92_, chained_data_delayed_6__91_, chained_data_delayed_6__90_, chained_data_delayed_6__89_, chained_data_delayed_6__88_, chained_data_delayed_6__87_, chained_data_delayed_6__86_, chained_data_delayed_6__85_, chained_data_delayed_6__84_, chained_data_delayed_6__83_, chained_data_delayed_6__82_, chained_data_delayed_6__81_, chained_data_delayed_6__80_, chained_data_delayed_6__79_, chained_data_delayed_6__78_, chained_data_delayed_6__77_, chained_data_delayed_6__76_, chained_data_delayed_6__75_, chained_data_delayed_6__74_, chained_data_delayed_6__73_, chained_data_delayed_6__72_, chained_data_delayed_6__71_, chained_data_delayed_6__70_, chained_data_delayed_6__69_, chained_data_delayed_6__68_, chained_data_delayed_6__67_, chained_data_delayed_6__66_, chained_data_delayed_6__65_, chained_data_delayed_6__64_, chained_data_delayed_6__63_, chained_data_delayed_6__62_, chained_data_delayed_6__61_, chained_data_delayed_6__60_, chained_data_delayed_6__59_, chained_data_delayed_6__58_, chained_data_delayed_6__57_, chained_data_delayed_6__56_, chained_data_delayed_6__55_, chained_data_delayed_6__54_, chained_data_delayed_6__53_, chained_data_delayed_6__52_, chained_data_delayed_6__51_, chained_data_delayed_6__50_, chained_data_delayed_6__49_, chained_data_delayed_6__48_, chained_data_delayed_6__47_, chained_data_delayed_6__46_, chained_data_delayed_6__45_, chained_data_delayed_6__44_, chained_data_delayed_6__43_, chained_data_delayed_6__42_, chained_data_delayed_6__41_, chained_data_delayed_6__40_, chained_data_delayed_6__39_, chained_data_delayed_6__38_, chained_data_delayed_6__37_, chained_data_delayed_6__36_, chained_data_delayed_6__35_, chained_data_delayed_6__34_, chained_data_delayed_6__33_, chained_data_delayed_6__32_, chained_data_delayed_6__31_, chained_data_delayed_6__30_, chained_data_delayed_6__29_, chained_data_delayed_6__28_, chained_data_delayed_6__27_, chained_data_delayed_6__26_, chained_data_delayed_6__25_, chained_data_delayed_6__24_, chained_data_delayed_6__23_, chained_data_delayed_6__22_, chained_data_delayed_6__21_, chained_data_delayed_6__20_, chained_data_delayed_6__19_, chained_data_delayed_6__18_, chained_data_delayed_6__17_, chained_data_delayed_6__16_, chained_data_delayed_6__15_, chained_data_delayed_6__14_, chained_data_delayed_6__13_, chained_data_delayed_6__12_, chained_data_delayed_6__11_, chained_data_delayed_6__10_, chained_data_delayed_6__9_, chained_data_delayed_6__8_, chained_data_delayed_6__7_, chained_data_delayed_6__6_, chained_data_delayed_6__5_, chained_data_delayed_6__4_, chained_data_delayed_6__3_, chained_data_delayed_6__2_, chained_data_delayed_6__1_, chained_data_delayed_6__0_ }),
    .data_o({ chained_data_delayed_7__127_, chained_data_delayed_7__126_, chained_data_delayed_7__125_, chained_data_delayed_7__124_, chained_data_delayed_7__123_, chained_data_delayed_7__122_, chained_data_delayed_7__121_, chained_data_delayed_7__120_, chained_data_delayed_7__119_, chained_data_delayed_7__118_, chained_data_delayed_7__117_, chained_data_delayed_7__116_, chained_data_delayed_7__115_, chained_data_delayed_7__114_, chained_data_delayed_7__113_, chained_data_delayed_7__112_, chained_data_delayed_7__111_, chained_data_delayed_7__110_, chained_data_delayed_7__109_, chained_data_delayed_7__108_, chained_data_delayed_7__107_, chained_data_delayed_7__106_, chained_data_delayed_7__105_, chained_data_delayed_7__104_, chained_data_delayed_7__103_, chained_data_delayed_7__102_, chained_data_delayed_7__101_, chained_data_delayed_7__100_, chained_data_delayed_7__99_, chained_data_delayed_7__98_, chained_data_delayed_7__97_, chained_data_delayed_7__96_, chained_data_delayed_7__95_, chained_data_delayed_7__94_, chained_data_delayed_7__93_, chained_data_delayed_7__92_, chained_data_delayed_7__91_, chained_data_delayed_7__90_, chained_data_delayed_7__89_, chained_data_delayed_7__88_, chained_data_delayed_7__87_, chained_data_delayed_7__86_, chained_data_delayed_7__85_, chained_data_delayed_7__84_, chained_data_delayed_7__83_, chained_data_delayed_7__82_, chained_data_delayed_7__81_, chained_data_delayed_7__80_, chained_data_delayed_7__79_, chained_data_delayed_7__78_, chained_data_delayed_7__77_, chained_data_delayed_7__76_, chained_data_delayed_7__75_, chained_data_delayed_7__74_, chained_data_delayed_7__73_, chained_data_delayed_7__72_, chained_data_delayed_7__71_, chained_data_delayed_7__70_, chained_data_delayed_7__69_, chained_data_delayed_7__68_, chained_data_delayed_7__67_, chained_data_delayed_7__66_, chained_data_delayed_7__65_, chained_data_delayed_7__64_, chained_data_delayed_7__63_, chained_data_delayed_7__62_, chained_data_delayed_7__61_, chained_data_delayed_7__60_, chained_data_delayed_7__59_, chained_data_delayed_7__58_, chained_data_delayed_7__57_, chained_data_delayed_7__56_, chained_data_delayed_7__55_, chained_data_delayed_7__54_, chained_data_delayed_7__53_, chained_data_delayed_7__52_, chained_data_delayed_7__51_, chained_data_delayed_7__50_, chained_data_delayed_7__49_, chained_data_delayed_7__48_, chained_data_delayed_7__47_, chained_data_delayed_7__46_, chained_data_delayed_7__45_, chained_data_delayed_7__44_, chained_data_delayed_7__43_, chained_data_delayed_7__42_, chained_data_delayed_7__41_, chained_data_delayed_7__40_, chained_data_delayed_7__39_, chained_data_delayed_7__38_, chained_data_delayed_7__37_, chained_data_delayed_7__36_, chained_data_delayed_7__35_, chained_data_delayed_7__34_, chained_data_delayed_7__33_, chained_data_delayed_7__32_, chained_data_delayed_7__31_, chained_data_delayed_7__30_, chained_data_delayed_7__29_, chained_data_delayed_7__28_, chained_data_delayed_7__27_, chained_data_delayed_7__26_, chained_data_delayed_7__25_, chained_data_delayed_7__24_, chained_data_delayed_7__23_, chained_data_delayed_7__22_, chained_data_delayed_7__21_, chained_data_delayed_7__20_, chained_data_delayed_7__19_, chained_data_delayed_7__18_, chained_data_delayed_7__17_, chained_data_delayed_7__16_, chained_data_delayed_7__15_, chained_data_delayed_7__14_, chained_data_delayed_7__13_, chained_data_delayed_7__12_, chained_data_delayed_7__11_, chained_data_delayed_7__10_, chained_data_delayed_7__9_, chained_data_delayed_7__8_, chained_data_delayed_7__7_, chained_data_delayed_7__6_, chained_data_delayed_7__5_, chained_data_delayed_7__4_, chained_data_delayed_7__3_, chained_data_delayed_7__2_, chained_data_delayed_7__1_, chained_data_delayed_7__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_8__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_7__127_, chained_data_delayed_7__126_, chained_data_delayed_7__125_, chained_data_delayed_7__124_, chained_data_delayed_7__123_, chained_data_delayed_7__122_, chained_data_delayed_7__121_, chained_data_delayed_7__120_, chained_data_delayed_7__119_, chained_data_delayed_7__118_, chained_data_delayed_7__117_, chained_data_delayed_7__116_, chained_data_delayed_7__115_, chained_data_delayed_7__114_, chained_data_delayed_7__113_, chained_data_delayed_7__112_, chained_data_delayed_7__111_, chained_data_delayed_7__110_, chained_data_delayed_7__109_, chained_data_delayed_7__108_, chained_data_delayed_7__107_, chained_data_delayed_7__106_, chained_data_delayed_7__105_, chained_data_delayed_7__104_, chained_data_delayed_7__103_, chained_data_delayed_7__102_, chained_data_delayed_7__101_, chained_data_delayed_7__100_, chained_data_delayed_7__99_, chained_data_delayed_7__98_, chained_data_delayed_7__97_, chained_data_delayed_7__96_, chained_data_delayed_7__95_, chained_data_delayed_7__94_, chained_data_delayed_7__93_, chained_data_delayed_7__92_, chained_data_delayed_7__91_, chained_data_delayed_7__90_, chained_data_delayed_7__89_, chained_data_delayed_7__88_, chained_data_delayed_7__87_, chained_data_delayed_7__86_, chained_data_delayed_7__85_, chained_data_delayed_7__84_, chained_data_delayed_7__83_, chained_data_delayed_7__82_, chained_data_delayed_7__81_, chained_data_delayed_7__80_, chained_data_delayed_7__79_, chained_data_delayed_7__78_, chained_data_delayed_7__77_, chained_data_delayed_7__76_, chained_data_delayed_7__75_, chained_data_delayed_7__74_, chained_data_delayed_7__73_, chained_data_delayed_7__72_, chained_data_delayed_7__71_, chained_data_delayed_7__70_, chained_data_delayed_7__69_, chained_data_delayed_7__68_, chained_data_delayed_7__67_, chained_data_delayed_7__66_, chained_data_delayed_7__65_, chained_data_delayed_7__64_, chained_data_delayed_7__63_, chained_data_delayed_7__62_, chained_data_delayed_7__61_, chained_data_delayed_7__60_, chained_data_delayed_7__59_, chained_data_delayed_7__58_, chained_data_delayed_7__57_, chained_data_delayed_7__56_, chained_data_delayed_7__55_, chained_data_delayed_7__54_, chained_data_delayed_7__53_, chained_data_delayed_7__52_, chained_data_delayed_7__51_, chained_data_delayed_7__50_, chained_data_delayed_7__49_, chained_data_delayed_7__48_, chained_data_delayed_7__47_, chained_data_delayed_7__46_, chained_data_delayed_7__45_, chained_data_delayed_7__44_, chained_data_delayed_7__43_, chained_data_delayed_7__42_, chained_data_delayed_7__41_, chained_data_delayed_7__40_, chained_data_delayed_7__39_, chained_data_delayed_7__38_, chained_data_delayed_7__37_, chained_data_delayed_7__36_, chained_data_delayed_7__35_, chained_data_delayed_7__34_, chained_data_delayed_7__33_, chained_data_delayed_7__32_, chained_data_delayed_7__31_, chained_data_delayed_7__30_, chained_data_delayed_7__29_, chained_data_delayed_7__28_, chained_data_delayed_7__27_, chained_data_delayed_7__26_, chained_data_delayed_7__25_, chained_data_delayed_7__24_, chained_data_delayed_7__23_, chained_data_delayed_7__22_, chained_data_delayed_7__21_, chained_data_delayed_7__20_, chained_data_delayed_7__19_, chained_data_delayed_7__18_, chained_data_delayed_7__17_, chained_data_delayed_7__16_, chained_data_delayed_7__15_, chained_data_delayed_7__14_, chained_data_delayed_7__13_, chained_data_delayed_7__12_, chained_data_delayed_7__11_, chained_data_delayed_7__10_, chained_data_delayed_7__9_, chained_data_delayed_7__8_, chained_data_delayed_7__7_, chained_data_delayed_7__6_, chained_data_delayed_7__5_, chained_data_delayed_7__4_, chained_data_delayed_7__3_, chained_data_delayed_7__2_, chained_data_delayed_7__1_, chained_data_delayed_7__0_ }),
    .data_o({ chained_data_delayed_8__127_, chained_data_delayed_8__126_, chained_data_delayed_8__125_, chained_data_delayed_8__124_, chained_data_delayed_8__123_, chained_data_delayed_8__122_, chained_data_delayed_8__121_, chained_data_delayed_8__120_, chained_data_delayed_8__119_, chained_data_delayed_8__118_, chained_data_delayed_8__117_, chained_data_delayed_8__116_, chained_data_delayed_8__115_, chained_data_delayed_8__114_, chained_data_delayed_8__113_, chained_data_delayed_8__112_, chained_data_delayed_8__111_, chained_data_delayed_8__110_, chained_data_delayed_8__109_, chained_data_delayed_8__108_, chained_data_delayed_8__107_, chained_data_delayed_8__106_, chained_data_delayed_8__105_, chained_data_delayed_8__104_, chained_data_delayed_8__103_, chained_data_delayed_8__102_, chained_data_delayed_8__101_, chained_data_delayed_8__100_, chained_data_delayed_8__99_, chained_data_delayed_8__98_, chained_data_delayed_8__97_, chained_data_delayed_8__96_, chained_data_delayed_8__95_, chained_data_delayed_8__94_, chained_data_delayed_8__93_, chained_data_delayed_8__92_, chained_data_delayed_8__91_, chained_data_delayed_8__90_, chained_data_delayed_8__89_, chained_data_delayed_8__88_, chained_data_delayed_8__87_, chained_data_delayed_8__86_, chained_data_delayed_8__85_, chained_data_delayed_8__84_, chained_data_delayed_8__83_, chained_data_delayed_8__82_, chained_data_delayed_8__81_, chained_data_delayed_8__80_, chained_data_delayed_8__79_, chained_data_delayed_8__78_, chained_data_delayed_8__77_, chained_data_delayed_8__76_, chained_data_delayed_8__75_, chained_data_delayed_8__74_, chained_data_delayed_8__73_, chained_data_delayed_8__72_, chained_data_delayed_8__71_, chained_data_delayed_8__70_, chained_data_delayed_8__69_, chained_data_delayed_8__68_, chained_data_delayed_8__67_, chained_data_delayed_8__66_, chained_data_delayed_8__65_, chained_data_delayed_8__64_, chained_data_delayed_8__63_, chained_data_delayed_8__62_, chained_data_delayed_8__61_, chained_data_delayed_8__60_, chained_data_delayed_8__59_, chained_data_delayed_8__58_, chained_data_delayed_8__57_, chained_data_delayed_8__56_, chained_data_delayed_8__55_, chained_data_delayed_8__54_, chained_data_delayed_8__53_, chained_data_delayed_8__52_, chained_data_delayed_8__51_, chained_data_delayed_8__50_, chained_data_delayed_8__49_, chained_data_delayed_8__48_, chained_data_delayed_8__47_, chained_data_delayed_8__46_, chained_data_delayed_8__45_, chained_data_delayed_8__44_, chained_data_delayed_8__43_, chained_data_delayed_8__42_, chained_data_delayed_8__41_, chained_data_delayed_8__40_, chained_data_delayed_8__39_, chained_data_delayed_8__38_, chained_data_delayed_8__37_, chained_data_delayed_8__36_, chained_data_delayed_8__35_, chained_data_delayed_8__34_, chained_data_delayed_8__33_, chained_data_delayed_8__32_, chained_data_delayed_8__31_, chained_data_delayed_8__30_, chained_data_delayed_8__29_, chained_data_delayed_8__28_, chained_data_delayed_8__27_, chained_data_delayed_8__26_, chained_data_delayed_8__25_, chained_data_delayed_8__24_, chained_data_delayed_8__23_, chained_data_delayed_8__22_, chained_data_delayed_8__21_, chained_data_delayed_8__20_, chained_data_delayed_8__19_, chained_data_delayed_8__18_, chained_data_delayed_8__17_, chained_data_delayed_8__16_, chained_data_delayed_8__15_, chained_data_delayed_8__14_, chained_data_delayed_8__13_, chained_data_delayed_8__12_, chained_data_delayed_8__11_, chained_data_delayed_8__10_, chained_data_delayed_8__9_, chained_data_delayed_8__8_, chained_data_delayed_8__7_, chained_data_delayed_8__6_, chained_data_delayed_8__5_, chained_data_delayed_8__4_, chained_data_delayed_8__3_, chained_data_delayed_8__2_, chained_data_delayed_8__1_, chained_data_delayed_8__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_9__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_8__127_, chained_data_delayed_8__126_, chained_data_delayed_8__125_, chained_data_delayed_8__124_, chained_data_delayed_8__123_, chained_data_delayed_8__122_, chained_data_delayed_8__121_, chained_data_delayed_8__120_, chained_data_delayed_8__119_, chained_data_delayed_8__118_, chained_data_delayed_8__117_, chained_data_delayed_8__116_, chained_data_delayed_8__115_, chained_data_delayed_8__114_, chained_data_delayed_8__113_, chained_data_delayed_8__112_, chained_data_delayed_8__111_, chained_data_delayed_8__110_, chained_data_delayed_8__109_, chained_data_delayed_8__108_, chained_data_delayed_8__107_, chained_data_delayed_8__106_, chained_data_delayed_8__105_, chained_data_delayed_8__104_, chained_data_delayed_8__103_, chained_data_delayed_8__102_, chained_data_delayed_8__101_, chained_data_delayed_8__100_, chained_data_delayed_8__99_, chained_data_delayed_8__98_, chained_data_delayed_8__97_, chained_data_delayed_8__96_, chained_data_delayed_8__95_, chained_data_delayed_8__94_, chained_data_delayed_8__93_, chained_data_delayed_8__92_, chained_data_delayed_8__91_, chained_data_delayed_8__90_, chained_data_delayed_8__89_, chained_data_delayed_8__88_, chained_data_delayed_8__87_, chained_data_delayed_8__86_, chained_data_delayed_8__85_, chained_data_delayed_8__84_, chained_data_delayed_8__83_, chained_data_delayed_8__82_, chained_data_delayed_8__81_, chained_data_delayed_8__80_, chained_data_delayed_8__79_, chained_data_delayed_8__78_, chained_data_delayed_8__77_, chained_data_delayed_8__76_, chained_data_delayed_8__75_, chained_data_delayed_8__74_, chained_data_delayed_8__73_, chained_data_delayed_8__72_, chained_data_delayed_8__71_, chained_data_delayed_8__70_, chained_data_delayed_8__69_, chained_data_delayed_8__68_, chained_data_delayed_8__67_, chained_data_delayed_8__66_, chained_data_delayed_8__65_, chained_data_delayed_8__64_, chained_data_delayed_8__63_, chained_data_delayed_8__62_, chained_data_delayed_8__61_, chained_data_delayed_8__60_, chained_data_delayed_8__59_, chained_data_delayed_8__58_, chained_data_delayed_8__57_, chained_data_delayed_8__56_, chained_data_delayed_8__55_, chained_data_delayed_8__54_, chained_data_delayed_8__53_, chained_data_delayed_8__52_, chained_data_delayed_8__51_, chained_data_delayed_8__50_, chained_data_delayed_8__49_, chained_data_delayed_8__48_, chained_data_delayed_8__47_, chained_data_delayed_8__46_, chained_data_delayed_8__45_, chained_data_delayed_8__44_, chained_data_delayed_8__43_, chained_data_delayed_8__42_, chained_data_delayed_8__41_, chained_data_delayed_8__40_, chained_data_delayed_8__39_, chained_data_delayed_8__38_, chained_data_delayed_8__37_, chained_data_delayed_8__36_, chained_data_delayed_8__35_, chained_data_delayed_8__34_, chained_data_delayed_8__33_, chained_data_delayed_8__32_, chained_data_delayed_8__31_, chained_data_delayed_8__30_, chained_data_delayed_8__29_, chained_data_delayed_8__28_, chained_data_delayed_8__27_, chained_data_delayed_8__26_, chained_data_delayed_8__25_, chained_data_delayed_8__24_, chained_data_delayed_8__23_, chained_data_delayed_8__22_, chained_data_delayed_8__21_, chained_data_delayed_8__20_, chained_data_delayed_8__19_, chained_data_delayed_8__18_, chained_data_delayed_8__17_, chained_data_delayed_8__16_, chained_data_delayed_8__15_, chained_data_delayed_8__14_, chained_data_delayed_8__13_, chained_data_delayed_8__12_, chained_data_delayed_8__11_, chained_data_delayed_8__10_, chained_data_delayed_8__9_, chained_data_delayed_8__8_, chained_data_delayed_8__7_, chained_data_delayed_8__6_, chained_data_delayed_8__5_, chained_data_delayed_8__4_, chained_data_delayed_8__3_, chained_data_delayed_8__2_, chained_data_delayed_8__1_, chained_data_delayed_8__0_ }),
    .data_o({ chained_data_delayed_9__127_, chained_data_delayed_9__126_, chained_data_delayed_9__125_, chained_data_delayed_9__124_, chained_data_delayed_9__123_, chained_data_delayed_9__122_, chained_data_delayed_9__121_, chained_data_delayed_9__120_, chained_data_delayed_9__119_, chained_data_delayed_9__118_, chained_data_delayed_9__117_, chained_data_delayed_9__116_, chained_data_delayed_9__115_, chained_data_delayed_9__114_, chained_data_delayed_9__113_, chained_data_delayed_9__112_, chained_data_delayed_9__111_, chained_data_delayed_9__110_, chained_data_delayed_9__109_, chained_data_delayed_9__108_, chained_data_delayed_9__107_, chained_data_delayed_9__106_, chained_data_delayed_9__105_, chained_data_delayed_9__104_, chained_data_delayed_9__103_, chained_data_delayed_9__102_, chained_data_delayed_9__101_, chained_data_delayed_9__100_, chained_data_delayed_9__99_, chained_data_delayed_9__98_, chained_data_delayed_9__97_, chained_data_delayed_9__96_, chained_data_delayed_9__95_, chained_data_delayed_9__94_, chained_data_delayed_9__93_, chained_data_delayed_9__92_, chained_data_delayed_9__91_, chained_data_delayed_9__90_, chained_data_delayed_9__89_, chained_data_delayed_9__88_, chained_data_delayed_9__87_, chained_data_delayed_9__86_, chained_data_delayed_9__85_, chained_data_delayed_9__84_, chained_data_delayed_9__83_, chained_data_delayed_9__82_, chained_data_delayed_9__81_, chained_data_delayed_9__80_, chained_data_delayed_9__79_, chained_data_delayed_9__78_, chained_data_delayed_9__77_, chained_data_delayed_9__76_, chained_data_delayed_9__75_, chained_data_delayed_9__74_, chained_data_delayed_9__73_, chained_data_delayed_9__72_, chained_data_delayed_9__71_, chained_data_delayed_9__70_, chained_data_delayed_9__69_, chained_data_delayed_9__68_, chained_data_delayed_9__67_, chained_data_delayed_9__66_, chained_data_delayed_9__65_, chained_data_delayed_9__64_, chained_data_delayed_9__63_, chained_data_delayed_9__62_, chained_data_delayed_9__61_, chained_data_delayed_9__60_, chained_data_delayed_9__59_, chained_data_delayed_9__58_, chained_data_delayed_9__57_, chained_data_delayed_9__56_, chained_data_delayed_9__55_, chained_data_delayed_9__54_, chained_data_delayed_9__53_, chained_data_delayed_9__52_, chained_data_delayed_9__51_, chained_data_delayed_9__50_, chained_data_delayed_9__49_, chained_data_delayed_9__48_, chained_data_delayed_9__47_, chained_data_delayed_9__46_, chained_data_delayed_9__45_, chained_data_delayed_9__44_, chained_data_delayed_9__43_, chained_data_delayed_9__42_, chained_data_delayed_9__41_, chained_data_delayed_9__40_, chained_data_delayed_9__39_, chained_data_delayed_9__38_, chained_data_delayed_9__37_, chained_data_delayed_9__36_, chained_data_delayed_9__35_, chained_data_delayed_9__34_, chained_data_delayed_9__33_, chained_data_delayed_9__32_, chained_data_delayed_9__31_, chained_data_delayed_9__30_, chained_data_delayed_9__29_, chained_data_delayed_9__28_, chained_data_delayed_9__27_, chained_data_delayed_9__26_, chained_data_delayed_9__25_, chained_data_delayed_9__24_, chained_data_delayed_9__23_, chained_data_delayed_9__22_, chained_data_delayed_9__21_, chained_data_delayed_9__20_, chained_data_delayed_9__19_, chained_data_delayed_9__18_, chained_data_delayed_9__17_, chained_data_delayed_9__16_, chained_data_delayed_9__15_, chained_data_delayed_9__14_, chained_data_delayed_9__13_, chained_data_delayed_9__12_, chained_data_delayed_9__11_, chained_data_delayed_9__10_, chained_data_delayed_9__9_, chained_data_delayed_9__8_, chained_data_delayed_9__7_, chained_data_delayed_9__6_, chained_data_delayed_9__5_, chained_data_delayed_9__4_, chained_data_delayed_9__3_, chained_data_delayed_9__2_, chained_data_delayed_9__1_, chained_data_delayed_9__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_10__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_9__127_, chained_data_delayed_9__126_, chained_data_delayed_9__125_, chained_data_delayed_9__124_, chained_data_delayed_9__123_, chained_data_delayed_9__122_, chained_data_delayed_9__121_, chained_data_delayed_9__120_, chained_data_delayed_9__119_, chained_data_delayed_9__118_, chained_data_delayed_9__117_, chained_data_delayed_9__116_, chained_data_delayed_9__115_, chained_data_delayed_9__114_, chained_data_delayed_9__113_, chained_data_delayed_9__112_, chained_data_delayed_9__111_, chained_data_delayed_9__110_, chained_data_delayed_9__109_, chained_data_delayed_9__108_, chained_data_delayed_9__107_, chained_data_delayed_9__106_, chained_data_delayed_9__105_, chained_data_delayed_9__104_, chained_data_delayed_9__103_, chained_data_delayed_9__102_, chained_data_delayed_9__101_, chained_data_delayed_9__100_, chained_data_delayed_9__99_, chained_data_delayed_9__98_, chained_data_delayed_9__97_, chained_data_delayed_9__96_, chained_data_delayed_9__95_, chained_data_delayed_9__94_, chained_data_delayed_9__93_, chained_data_delayed_9__92_, chained_data_delayed_9__91_, chained_data_delayed_9__90_, chained_data_delayed_9__89_, chained_data_delayed_9__88_, chained_data_delayed_9__87_, chained_data_delayed_9__86_, chained_data_delayed_9__85_, chained_data_delayed_9__84_, chained_data_delayed_9__83_, chained_data_delayed_9__82_, chained_data_delayed_9__81_, chained_data_delayed_9__80_, chained_data_delayed_9__79_, chained_data_delayed_9__78_, chained_data_delayed_9__77_, chained_data_delayed_9__76_, chained_data_delayed_9__75_, chained_data_delayed_9__74_, chained_data_delayed_9__73_, chained_data_delayed_9__72_, chained_data_delayed_9__71_, chained_data_delayed_9__70_, chained_data_delayed_9__69_, chained_data_delayed_9__68_, chained_data_delayed_9__67_, chained_data_delayed_9__66_, chained_data_delayed_9__65_, chained_data_delayed_9__64_, chained_data_delayed_9__63_, chained_data_delayed_9__62_, chained_data_delayed_9__61_, chained_data_delayed_9__60_, chained_data_delayed_9__59_, chained_data_delayed_9__58_, chained_data_delayed_9__57_, chained_data_delayed_9__56_, chained_data_delayed_9__55_, chained_data_delayed_9__54_, chained_data_delayed_9__53_, chained_data_delayed_9__52_, chained_data_delayed_9__51_, chained_data_delayed_9__50_, chained_data_delayed_9__49_, chained_data_delayed_9__48_, chained_data_delayed_9__47_, chained_data_delayed_9__46_, chained_data_delayed_9__45_, chained_data_delayed_9__44_, chained_data_delayed_9__43_, chained_data_delayed_9__42_, chained_data_delayed_9__41_, chained_data_delayed_9__40_, chained_data_delayed_9__39_, chained_data_delayed_9__38_, chained_data_delayed_9__37_, chained_data_delayed_9__36_, chained_data_delayed_9__35_, chained_data_delayed_9__34_, chained_data_delayed_9__33_, chained_data_delayed_9__32_, chained_data_delayed_9__31_, chained_data_delayed_9__30_, chained_data_delayed_9__29_, chained_data_delayed_9__28_, chained_data_delayed_9__27_, chained_data_delayed_9__26_, chained_data_delayed_9__25_, chained_data_delayed_9__24_, chained_data_delayed_9__23_, chained_data_delayed_9__22_, chained_data_delayed_9__21_, chained_data_delayed_9__20_, chained_data_delayed_9__19_, chained_data_delayed_9__18_, chained_data_delayed_9__17_, chained_data_delayed_9__16_, chained_data_delayed_9__15_, chained_data_delayed_9__14_, chained_data_delayed_9__13_, chained_data_delayed_9__12_, chained_data_delayed_9__11_, chained_data_delayed_9__10_, chained_data_delayed_9__9_, chained_data_delayed_9__8_, chained_data_delayed_9__7_, chained_data_delayed_9__6_, chained_data_delayed_9__5_, chained_data_delayed_9__4_, chained_data_delayed_9__3_, chained_data_delayed_9__2_, chained_data_delayed_9__1_, chained_data_delayed_9__0_ }),
    .data_o({ chained_data_delayed_10__127_, chained_data_delayed_10__126_, chained_data_delayed_10__125_, chained_data_delayed_10__124_, chained_data_delayed_10__123_, chained_data_delayed_10__122_, chained_data_delayed_10__121_, chained_data_delayed_10__120_, chained_data_delayed_10__119_, chained_data_delayed_10__118_, chained_data_delayed_10__117_, chained_data_delayed_10__116_, chained_data_delayed_10__115_, chained_data_delayed_10__114_, chained_data_delayed_10__113_, chained_data_delayed_10__112_, chained_data_delayed_10__111_, chained_data_delayed_10__110_, chained_data_delayed_10__109_, chained_data_delayed_10__108_, chained_data_delayed_10__107_, chained_data_delayed_10__106_, chained_data_delayed_10__105_, chained_data_delayed_10__104_, chained_data_delayed_10__103_, chained_data_delayed_10__102_, chained_data_delayed_10__101_, chained_data_delayed_10__100_, chained_data_delayed_10__99_, chained_data_delayed_10__98_, chained_data_delayed_10__97_, chained_data_delayed_10__96_, chained_data_delayed_10__95_, chained_data_delayed_10__94_, chained_data_delayed_10__93_, chained_data_delayed_10__92_, chained_data_delayed_10__91_, chained_data_delayed_10__90_, chained_data_delayed_10__89_, chained_data_delayed_10__88_, chained_data_delayed_10__87_, chained_data_delayed_10__86_, chained_data_delayed_10__85_, chained_data_delayed_10__84_, chained_data_delayed_10__83_, chained_data_delayed_10__82_, chained_data_delayed_10__81_, chained_data_delayed_10__80_, chained_data_delayed_10__79_, chained_data_delayed_10__78_, chained_data_delayed_10__77_, chained_data_delayed_10__76_, chained_data_delayed_10__75_, chained_data_delayed_10__74_, chained_data_delayed_10__73_, chained_data_delayed_10__72_, chained_data_delayed_10__71_, chained_data_delayed_10__70_, chained_data_delayed_10__69_, chained_data_delayed_10__68_, chained_data_delayed_10__67_, chained_data_delayed_10__66_, chained_data_delayed_10__65_, chained_data_delayed_10__64_, chained_data_delayed_10__63_, chained_data_delayed_10__62_, chained_data_delayed_10__61_, chained_data_delayed_10__60_, chained_data_delayed_10__59_, chained_data_delayed_10__58_, chained_data_delayed_10__57_, chained_data_delayed_10__56_, chained_data_delayed_10__55_, chained_data_delayed_10__54_, chained_data_delayed_10__53_, chained_data_delayed_10__52_, chained_data_delayed_10__51_, chained_data_delayed_10__50_, chained_data_delayed_10__49_, chained_data_delayed_10__48_, chained_data_delayed_10__47_, chained_data_delayed_10__46_, chained_data_delayed_10__45_, chained_data_delayed_10__44_, chained_data_delayed_10__43_, chained_data_delayed_10__42_, chained_data_delayed_10__41_, chained_data_delayed_10__40_, chained_data_delayed_10__39_, chained_data_delayed_10__38_, chained_data_delayed_10__37_, chained_data_delayed_10__36_, chained_data_delayed_10__35_, chained_data_delayed_10__34_, chained_data_delayed_10__33_, chained_data_delayed_10__32_, chained_data_delayed_10__31_, chained_data_delayed_10__30_, chained_data_delayed_10__29_, chained_data_delayed_10__28_, chained_data_delayed_10__27_, chained_data_delayed_10__26_, chained_data_delayed_10__25_, chained_data_delayed_10__24_, chained_data_delayed_10__23_, chained_data_delayed_10__22_, chained_data_delayed_10__21_, chained_data_delayed_10__20_, chained_data_delayed_10__19_, chained_data_delayed_10__18_, chained_data_delayed_10__17_, chained_data_delayed_10__16_, chained_data_delayed_10__15_, chained_data_delayed_10__14_, chained_data_delayed_10__13_, chained_data_delayed_10__12_, chained_data_delayed_10__11_, chained_data_delayed_10__10_, chained_data_delayed_10__9_, chained_data_delayed_10__8_, chained_data_delayed_10__7_, chained_data_delayed_10__6_, chained_data_delayed_10__5_, chained_data_delayed_10__4_, chained_data_delayed_10__3_, chained_data_delayed_10__2_, chained_data_delayed_10__1_, chained_data_delayed_10__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_11__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_10__127_, chained_data_delayed_10__126_, chained_data_delayed_10__125_, chained_data_delayed_10__124_, chained_data_delayed_10__123_, chained_data_delayed_10__122_, chained_data_delayed_10__121_, chained_data_delayed_10__120_, chained_data_delayed_10__119_, chained_data_delayed_10__118_, chained_data_delayed_10__117_, chained_data_delayed_10__116_, chained_data_delayed_10__115_, chained_data_delayed_10__114_, chained_data_delayed_10__113_, chained_data_delayed_10__112_, chained_data_delayed_10__111_, chained_data_delayed_10__110_, chained_data_delayed_10__109_, chained_data_delayed_10__108_, chained_data_delayed_10__107_, chained_data_delayed_10__106_, chained_data_delayed_10__105_, chained_data_delayed_10__104_, chained_data_delayed_10__103_, chained_data_delayed_10__102_, chained_data_delayed_10__101_, chained_data_delayed_10__100_, chained_data_delayed_10__99_, chained_data_delayed_10__98_, chained_data_delayed_10__97_, chained_data_delayed_10__96_, chained_data_delayed_10__95_, chained_data_delayed_10__94_, chained_data_delayed_10__93_, chained_data_delayed_10__92_, chained_data_delayed_10__91_, chained_data_delayed_10__90_, chained_data_delayed_10__89_, chained_data_delayed_10__88_, chained_data_delayed_10__87_, chained_data_delayed_10__86_, chained_data_delayed_10__85_, chained_data_delayed_10__84_, chained_data_delayed_10__83_, chained_data_delayed_10__82_, chained_data_delayed_10__81_, chained_data_delayed_10__80_, chained_data_delayed_10__79_, chained_data_delayed_10__78_, chained_data_delayed_10__77_, chained_data_delayed_10__76_, chained_data_delayed_10__75_, chained_data_delayed_10__74_, chained_data_delayed_10__73_, chained_data_delayed_10__72_, chained_data_delayed_10__71_, chained_data_delayed_10__70_, chained_data_delayed_10__69_, chained_data_delayed_10__68_, chained_data_delayed_10__67_, chained_data_delayed_10__66_, chained_data_delayed_10__65_, chained_data_delayed_10__64_, chained_data_delayed_10__63_, chained_data_delayed_10__62_, chained_data_delayed_10__61_, chained_data_delayed_10__60_, chained_data_delayed_10__59_, chained_data_delayed_10__58_, chained_data_delayed_10__57_, chained_data_delayed_10__56_, chained_data_delayed_10__55_, chained_data_delayed_10__54_, chained_data_delayed_10__53_, chained_data_delayed_10__52_, chained_data_delayed_10__51_, chained_data_delayed_10__50_, chained_data_delayed_10__49_, chained_data_delayed_10__48_, chained_data_delayed_10__47_, chained_data_delayed_10__46_, chained_data_delayed_10__45_, chained_data_delayed_10__44_, chained_data_delayed_10__43_, chained_data_delayed_10__42_, chained_data_delayed_10__41_, chained_data_delayed_10__40_, chained_data_delayed_10__39_, chained_data_delayed_10__38_, chained_data_delayed_10__37_, chained_data_delayed_10__36_, chained_data_delayed_10__35_, chained_data_delayed_10__34_, chained_data_delayed_10__33_, chained_data_delayed_10__32_, chained_data_delayed_10__31_, chained_data_delayed_10__30_, chained_data_delayed_10__29_, chained_data_delayed_10__28_, chained_data_delayed_10__27_, chained_data_delayed_10__26_, chained_data_delayed_10__25_, chained_data_delayed_10__24_, chained_data_delayed_10__23_, chained_data_delayed_10__22_, chained_data_delayed_10__21_, chained_data_delayed_10__20_, chained_data_delayed_10__19_, chained_data_delayed_10__18_, chained_data_delayed_10__17_, chained_data_delayed_10__16_, chained_data_delayed_10__15_, chained_data_delayed_10__14_, chained_data_delayed_10__13_, chained_data_delayed_10__12_, chained_data_delayed_10__11_, chained_data_delayed_10__10_, chained_data_delayed_10__9_, chained_data_delayed_10__8_, chained_data_delayed_10__7_, chained_data_delayed_10__6_, chained_data_delayed_10__5_, chained_data_delayed_10__4_, chained_data_delayed_10__3_, chained_data_delayed_10__2_, chained_data_delayed_10__1_, chained_data_delayed_10__0_ }),
    .data_o({ chained_data_delayed_11__127_, chained_data_delayed_11__126_, chained_data_delayed_11__125_, chained_data_delayed_11__124_, chained_data_delayed_11__123_, chained_data_delayed_11__122_, chained_data_delayed_11__121_, chained_data_delayed_11__120_, chained_data_delayed_11__119_, chained_data_delayed_11__118_, chained_data_delayed_11__117_, chained_data_delayed_11__116_, chained_data_delayed_11__115_, chained_data_delayed_11__114_, chained_data_delayed_11__113_, chained_data_delayed_11__112_, chained_data_delayed_11__111_, chained_data_delayed_11__110_, chained_data_delayed_11__109_, chained_data_delayed_11__108_, chained_data_delayed_11__107_, chained_data_delayed_11__106_, chained_data_delayed_11__105_, chained_data_delayed_11__104_, chained_data_delayed_11__103_, chained_data_delayed_11__102_, chained_data_delayed_11__101_, chained_data_delayed_11__100_, chained_data_delayed_11__99_, chained_data_delayed_11__98_, chained_data_delayed_11__97_, chained_data_delayed_11__96_, chained_data_delayed_11__95_, chained_data_delayed_11__94_, chained_data_delayed_11__93_, chained_data_delayed_11__92_, chained_data_delayed_11__91_, chained_data_delayed_11__90_, chained_data_delayed_11__89_, chained_data_delayed_11__88_, chained_data_delayed_11__87_, chained_data_delayed_11__86_, chained_data_delayed_11__85_, chained_data_delayed_11__84_, chained_data_delayed_11__83_, chained_data_delayed_11__82_, chained_data_delayed_11__81_, chained_data_delayed_11__80_, chained_data_delayed_11__79_, chained_data_delayed_11__78_, chained_data_delayed_11__77_, chained_data_delayed_11__76_, chained_data_delayed_11__75_, chained_data_delayed_11__74_, chained_data_delayed_11__73_, chained_data_delayed_11__72_, chained_data_delayed_11__71_, chained_data_delayed_11__70_, chained_data_delayed_11__69_, chained_data_delayed_11__68_, chained_data_delayed_11__67_, chained_data_delayed_11__66_, chained_data_delayed_11__65_, chained_data_delayed_11__64_, chained_data_delayed_11__63_, chained_data_delayed_11__62_, chained_data_delayed_11__61_, chained_data_delayed_11__60_, chained_data_delayed_11__59_, chained_data_delayed_11__58_, chained_data_delayed_11__57_, chained_data_delayed_11__56_, chained_data_delayed_11__55_, chained_data_delayed_11__54_, chained_data_delayed_11__53_, chained_data_delayed_11__52_, chained_data_delayed_11__51_, chained_data_delayed_11__50_, chained_data_delayed_11__49_, chained_data_delayed_11__48_, chained_data_delayed_11__47_, chained_data_delayed_11__46_, chained_data_delayed_11__45_, chained_data_delayed_11__44_, chained_data_delayed_11__43_, chained_data_delayed_11__42_, chained_data_delayed_11__41_, chained_data_delayed_11__40_, chained_data_delayed_11__39_, chained_data_delayed_11__38_, chained_data_delayed_11__37_, chained_data_delayed_11__36_, chained_data_delayed_11__35_, chained_data_delayed_11__34_, chained_data_delayed_11__33_, chained_data_delayed_11__32_, chained_data_delayed_11__31_, chained_data_delayed_11__30_, chained_data_delayed_11__29_, chained_data_delayed_11__28_, chained_data_delayed_11__27_, chained_data_delayed_11__26_, chained_data_delayed_11__25_, chained_data_delayed_11__24_, chained_data_delayed_11__23_, chained_data_delayed_11__22_, chained_data_delayed_11__21_, chained_data_delayed_11__20_, chained_data_delayed_11__19_, chained_data_delayed_11__18_, chained_data_delayed_11__17_, chained_data_delayed_11__16_, chained_data_delayed_11__15_, chained_data_delayed_11__14_, chained_data_delayed_11__13_, chained_data_delayed_11__12_, chained_data_delayed_11__11_, chained_data_delayed_11__10_, chained_data_delayed_11__9_, chained_data_delayed_11__8_, chained_data_delayed_11__7_, chained_data_delayed_11__6_, chained_data_delayed_11__5_, chained_data_delayed_11__4_, chained_data_delayed_11__3_, chained_data_delayed_11__2_, chained_data_delayed_11__1_, chained_data_delayed_11__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_12__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_11__127_, chained_data_delayed_11__126_, chained_data_delayed_11__125_, chained_data_delayed_11__124_, chained_data_delayed_11__123_, chained_data_delayed_11__122_, chained_data_delayed_11__121_, chained_data_delayed_11__120_, chained_data_delayed_11__119_, chained_data_delayed_11__118_, chained_data_delayed_11__117_, chained_data_delayed_11__116_, chained_data_delayed_11__115_, chained_data_delayed_11__114_, chained_data_delayed_11__113_, chained_data_delayed_11__112_, chained_data_delayed_11__111_, chained_data_delayed_11__110_, chained_data_delayed_11__109_, chained_data_delayed_11__108_, chained_data_delayed_11__107_, chained_data_delayed_11__106_, chained_data_delayed_11__105_, chained_data_delayed_11__104_, chained_data_delayed_11__103_, chained_data_delayed_11__102_, chained_data_delayed_11__101_, chained_data_delayed_11__100_, chained_data_delayed_11__99_, chained_data_delayed_11__98_, chained_data_delayed_11__97_, chained_data_delayed_11__96_, chained_data_delayed_11__95_, chained_data_delayed_11__94_, chained_data_delayed_11__93_, chained_data_delayed_11__92_, chained_data_delayed_11__91_, chained_data_delayed_11__90_, chained_data_delayed_11__89_, chained_data_delayed_11__88_, chained_data_delayed_11__87_, chained_data_delayed_11__86_, chained_data_delayed_11__85_, chained_data_delayed_11__84_, chained_data_delayed_11__83_, chained_data_delayed_11__82_, chained_data_delayed_11__81_, chained_data_delayed_11__80_, chained_data_delayed_11__79_, chained_data_delayed_11__78_, chained_data_delayed_11__77_, chained_data_delayed_11__76_, chained_data_delayed_11__75_, chained_data_delayed_11__74_, chained_data_delayed_11__73_, chained_data_delayed_11__72_, chained_data_delayed_11__71_, chained_data_delayed_11__70_, chained_data_delayed_11__69_, chained_data_delayed_11__68_, chained_data_delayed_11__67_, chained_data_delayed_11__66_, chained_data_delayed_11__65_, chained_data_delayed_11__64_, chained_data_delayed_11__63_, chained_data_delayed_11__62_, chained_data_delayed_11__61_, chained_data_delayed_11__60_, chained_data_delayed_11__59_, chained_data_delayed_11__58_, chained_data_delayed_11__57_, chained_data_delayed_11__56_, chained_data_delayed_11__55_, chained_data_delayed_11__54_, chained_data_delayed_11__53_, chained_data_delayed_11__52_, chained_data_delayed_11__51_, chained_data_delayed_11__50_, chained_data_delayed_11__49_, chained_data_delayed_11__48_, chained_data_delayed_11__47_, chained_data_delayed_11__46_, chained_data_delayed_11__45_, chained_data_delayed_11__44_, chained_data_delayed_11__43_, chained_data_delayed_11__42_, chained_data_delayed_11__41_, chained_data_delayed_11__40_, chained_data_delayed_11__39_, chained_data_delayed_11__38_, chained_data_delayed_11__37_, chained_data_delayed_11__36_, chained_data_delayed_11__35_, chained_data_delayed_11__34_, chained_data_delayed_11__33_, chained_data_delayed_11__32_, chained_data_delayed_11__31_, chained_data_delayed_11__30_, chained_data_delayed_11__29_, chained_data_delayed_11__28_, chained_data_delayed_11__27_, chained_data_delayed_11__26_, chained_data_delayed_11__25_, chained_data_delayed_11__24_, chained_data_delayed_11__23_, chained_data_delayed_11__22_, chained_data_delayed_11__21_, chained_data_delayed_11__20_, chained_data_delayed_11__19_, chained_data_delayed_11__18_, chained_data_delayed_11__17_, chained_data_delayed_11__16_, chained_data_delayed_11__15_, chained_data_delayed_11__14_, chained_data_delayed_11__13_, chained_data_delayed_11__12_, chained_data_delayed_11__11_, chained_data_delayed_11__10_, chained_data_delayed_11__9_, chained_data_delayed_11__8_, chained_data_delayed_11__7_, chained_data_delayed_11__6_, chained_data_delayed_11__5_, chained_data_delayed_11__4_, chained_data_delayed_11__3_, chained_data_delayed_11__2_, chained_data_delayed_11__1_, chained_data_delayed_11__0_ }),
    .data_o({ chained_data_delayed_12__127_, chained_data_delayed_12__126_, chained_data_delayed_12__125_, chained_data_delayed_12__124_, chained_data_delayed_12__123_, chained_data_delayed_12__122_, chained_data_delayed_12__121_, chained_data_delayed_12__120_, chained_data_delayed_12__119_, chained_data_delayed_12__118_, chained_data_delayed_12__117_, chained_data_delayed_12__116_, chained_data_delayed_12__115_, chained_data_delayed_12__114_, chained_data_delayed_12__113_, chained_data_delayed_12__112_, chained_data_delayed_12__111_, chained_data_delayed_12__110_, chained_data_delayed_12__109_, chained_data_delayed_12__108_, chained_data_delayed_12__107_, chained_data_delayed_12__106_, chained_data_delayed_12__105_, chained_data_delayed_12__104_, chained_data_delayed_12__103_, chained_data_delayed_12__102_, chained_data_delayed_12__101_, chained_data_delayed_12__100_, chained_data_delayed_12__99_, chained_data_delayed_12__98_, chained_data_delayed_12__97_, chained_data_delayed_12__96_, chained_data_delayed_12__95_, chained_data_delayed_12__94_, chained_data_delayed_12__93_, chained_data_delayed_12__92_, chained_data_delayed_12__91_, chained_data_delayed_12__90_, chained_data_delayed_12__89_, chained_data_delayed_12__88_, chained_data_delayed_12__87_, chained_data_delayed_12__86_, chained_data_delayed_12__85_, chained_data_delayed_12__84_, chained_data_delayed_12__83_, chained_data_delayed_12__82_, chained_data_delayed_12__81_, chained_data_delayed_12__80_, chained_data_delayed_12__79_, chained_data_delayed_12__78_, chained_data_delayed_12__77_, chained_data_delayed_12__76_, chained_data_delayed_12__75_, chained_data_delayed_12__74_, chained_data_delayed_12__73_, chained_data_delayed_12__72_, chained_data_delayed_12__71_, chained_data_delayed_12__70_, chained_data_delayed_12__69_, chained_data_delayed_12__68_, chained_data_delayed_12__67_, chained_data_delayed_12__66_, chained_data_delayed_12__65_, chained_data_delayed_12__64_, chained_data_delayed_12__63_, chained_data_delayed_12__62_, chained_data_delayed_12__61_, chained_data_delayed_12__60_, chained_data_delayed_12__59_, chained_data_delayed_12__58_, chained_data_delayed_12__57_, chained_data_delayed_12__56_, chained_data_delayed_12__55_, chained_data_delayed_12__54_, chained_data_delayed_12__53_, chained_data_delayed_12__52_, chained_data_delayed_12__51_, chained_data_delayed_12__50_, chained_data_delayed_12__49_, chained_data_delayed_12__48_, chained_data_delayed_12__47_, chained_data_delayed_12__46_, chained_data_delayed_12__45_, chained_data_delayed_12__44_, chained_data_delayed_12__43_, chained_data_delayed_12__42_, chained_data_delayed_12__41_, chained_data_delayed_12__40_, chained_data_delayed_12__39_, chained_data_delayed_12__38_, chained_data_delayed_12__37_, chained_data_delayed_12__36_, chained_data_delayed_12__35_, chained_data_delayed_12__34_, chained_data_delayed_12__33_, chained_data_delayed_12__32_, chained_data_delayed_12__31_, chained_data_delayed_12__30_, chained_data_delayed_12__29_, chained_data_delayed_12__28_, chained_data_delayed_12__27_, chained_data_delayed_12__26_, chained_data_delayed_12__25_, chained_data_delayed_12__24_, chained_data_delayed_12__23_, chained_data_delayed_12__22_, chained_data_delayed_12__21_, chained_data_delayed_12__20_, chained_data_delayed_12__19_, chained_data_delayed_12__18_, chained_data_delayed_12__17_, chained_data_delayed_12__16_, chained_data_delayed_12__15_, chained_data_delayed_12__14_, chained_data_delayed_12__13_, chained_data_delayed_12__12_, chained_data_delayed_12__11_, chained_data_delayed_12__10_, chained_data_delayed_12__9_, chained_data_delayed_12__8_, chained_data_delayed_12__7_, chained_data_delayed_12__6_, chained_data_delayed_12__5_, chained_data_delayed_12__4_, chained_data_delayed_12__3_, chained_data_delayed_12__2_, chained_data_delayed_12__1_, chained_data_delayed_12__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_13__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_12__127_, chained_data_delayed_12__126_, chained_data_delayed_12__125_, chained_data_delayed_12__124_, chained_data_delayed_12__123_, chained_data_delayed_12__122_, chained_data_delayed_12__121_, chained_data_delayed_12__120_, chained_data_delayed_12__119_, chained_data_delayed_12__118_, chained_data_delayed_12__117_, chained_data_delayed_12__116_, chained_data_delayed_12__115_, chained_data_delayed_12__114_, chained_data_delayed_12__113_, chained_data_delayed_12__112_, chained_data_delayed_12__111_, chained_data_delayed_12__110_, chained_data_delayed_12__109_, chained_data_delayed_12__108_, chained_data_delayed_12__107_, chained_data_delayed_12__106_, chained_data_delayed_12__105_, chained_data_delayed_12__104_, chained_data_delayed_12__103_, chained_data_delayed_12__102_, chained_data_delayed_12__101_, chained_data_delayed_12__100_, chained_data_delayed_12__99_, chained_data_delayed_12__98_, chained_data_delayed_12__97_, chained_data_delayed_12__96_, chained_data_delayed_12__95_, chained_data_delayed_12__94_, chained_data_delayed_12__93_, chained_data_delayed_12__92_, chained_data_delayed_12__91_, chained_data_delayed_12__90_, chained_data_delayed_12__89_, chained_data_delayed_12__88_, chained_data_delayed_12__87_, chained_data_delayed_12__86_, chained_data_delayed_12__85_, chained_data_delayed_12__84_, chained_data_delayed_12__83_, chained_data_delayed_12__82_, chained_data_delayed_12__81_, chained_data_delayed_12__80_, chained_data_delayed_12__79_, chained_data_delayed_12__78_, chained_data_delayed_12__77_, chained_data_delayed_12__76_, chained_data_delayed_12__75_, chained_data_delayed_12__74_, chained_data_delayed_12__73_, chained_data_delayed_12__72_, chained_data_delayed_12__71_, chained_data_delayed_12__70_, chained_data_delayed_12__69_, chained_data_delayed_12__68_, chained_data_delayed_12__67_, chained_data_delayed_12__66_, chained_data_delayed_12__65_, chained_data_delayed_12__64_, chained_data_delayed_12__63_, chained_data_delayed_12__62_, chained_data_delayed_12__61_, chained_data_delayed_12__60_, chained_data_delayed_12__59_, chained_data_delayed_12__58_, chained_data_delayed_12__57_, chained_data_delayed_12__56_, chained_data_delayed_12__55_, chained_data_delayed_12__54_, chained_data_delayed_12__53_, chained_data_delayed_12__52_, chained_data_delayed_12__51_, chained_data_delayed_12__50_, chained_data_delayed_12__49_, chained_data_delayed_12__48_, chained_data_delayed_12__47_, chained_data_delayed_12__46_, chained_data_delayed_12__45_, chained_data_delayed_12__44_, chained_data_delayed_12__43_, chained_data_delayed_12__42_, chained_data_delayed_12__41_, chained_data_delayed_12__40_, chained_data_delayed_12__39_, chained_data_delayed_12__38_, chained_data_delayed_12__37_, chained_data_delayed_12__36_, chained_data_delayed_12__35_, chained_data_delayed_12__34_, chained_data_delayed_12__33_, chained_data_delayed_12__32_, chained_data_delayed_12__31_, chained_data_delayed_12__30_, chained_data_delayed_12__29_, chained_data_delayed_12__28_, chained_data_delayed_12__27_, chained_data_delayed_12__26_, chained_data_delayed_12__25_, chained_data_delayed_12__24_, chained_data_delayed_12__23_, chained_data_delayed_12__22_, chained_data_delayed_12__21_, chained_data_delayed_12__20_, chained_data_delayed_12__19_, chained_data_delayed_12__18_, chained_data_delayed_12__17_, chained_data_delayed_12__16_, chained_data_delayed_12__15_, chained_data_delayed_12__14_, chained_data_delayed_12__13_, chained_data_delayed_12__12_, chained_data_delayed_12__11_, chained_data_delayed_12__10_, chained_data_delayed_12__9_, chained_data_delayed_12__8_, chained_data_delayed_12__7_, chained_data_delayed_12__6_, chained_data_delayed_12__5_, chained_data_delayed_12__4_, chained_data_delayed_12__3_, chained_data_delayed_12__2_, chained_data_delayed_12__1_, chained_data_delayed_12__0_ }),
    .data_o({ chained_data_delayed_13__127_, chained_data_delayed_13__126_, chained_data_delayed_13__125_, chained_data_delayed_13__124_, chained_data_delayed_13__123_, chained_data_delayed_13__122_, chained_data_delayed_13__121_, chained_data_delayed_13__120_, chained_data_delayed_13__119_, chained_data_delayed_13__118_, chained_data_delayed_13__117_, chained_data_delayed_13__116_, chained_data_delayed_13__115_, chained_data_delayed_13__114_, chained_data_delayed_13__113_, chained_data_delayed_13__112_, chained_data_delayed_13__111_, chained_data_delayed_13__110_, chained_data_delayed_13__109_, chained_data_delayed_13__108_, chained_data_delayed_13__107_, chained_data_delayed_13__106_, chained_data_delayed_13__105_, chained_data_delayed_13__104_, chained_data_delayed_13__103_, chained_data_delayed_13__102_, chained_data_delayed_13__101_, chained_data_delayed_13__100_, chained_data_delayed_13__99_, chained_data_delayed_13__98_, chained_data_delayed_13__97_, chained_data_delayed_13__96_, chained_data_delayed_13__95_, chained_data_delayed_13__94_, chained_data_delayed_13__93_, chained_data_delayed_13__92_, chained_data_delayed_13__91_, chained_data_delayed_13__90_, chained_data_delayed_13__89_, chained_data_delayed_13__88_, chained_data_delayed_13__87_, chained_data_delayed_13__86_, chained_data_delayed_13__85_, chained_data_delayed_13__84_, chained_data_delayed_13__83_, chained_data_delayed_13__82_, chained_data_delayed_13__81_, chained_data_delayed_13__80_, chained_data_delayed_13__79_, chained_data_delayed_13__78_, chained_data_delayed_13__77_, chained_data_delayed_13__76_, chained_data_delayed_13__75_, chained_data_delayed_13__74_, chained_data_delayed_13__73_, chained_data_delayed_13__72_, chained_data_delayed_13__71_, chained_data_delayed_13__70_, chained_data_delayed_13__69_, chained_data_delayed_13__68_, chained_data_delayed_13__67_, chained_data_delayed_13__66_, chained_data_delayed_13__65_, chained_data_delayed_13__64_, chained_data_delayed_13__63_, chained_data_delayed_13__62_, chained_data_delayed_13__61_, chained_data_delayed_13__60_, chained_data_delayed_13__59_, chained_data_delayed_13__58_, chained_data_delayed_13__57_, chained_data_delayed_13__56_, chained_data_delayed_13__55_, chained_data_delayed_13__54_, chained_data_delayed_13__53_, chained_data_delayed_13__52_, chained_data_delayed_13__51_, chained_data_delayed_13__50_, chained_data_delayed_13__49_, chained_data_delayed_13__48_, chained_data_delayed_13__47_, chained_data_delayed_13__46_, chained_data_delayed_13__45_, chained_data_delayed_13__44_, chained_data_delayed_13__43_, chained_data_delayed_13__42_, chained_data_delayed_13__41_, chained_data_delayed_13__40_, chained_data_delayed_13__39_, chained_data_delayed_13__38_, chained_data_delayed_13__37_, chained_data_delayed_13__36_, chained_data_delayed_13__35_, chained_data_delayed_13__34_, chained_data_delayed_13__33_, chained_data_delayed_13__32_, chained_data_delayed_13__31_, chained_data_delayed_13__30_, chained_data_delayed_13__29_, chained_data_delayed_13__28_, chained_data_delayed_13__27_, chained_data_delayed_13__26_, chained_data_delayed_13__25_, chained_data_delayed_13__24_, chained_data_delayed_13__23_, chained_data_delayed_13__22_, chained_data_delayed_13__21_, chained_data_delayed_13__20_, chained_data_delayed_13__19_, chained_data_delayed_13__18_, chained_data_delayed_13__17_, chained_data_delayed_13__16_, chained_data_delayed_13__15_, chained_data_delayed_13__14_, chained_data_delayed_13__13_, chained_data_delayed_13__12_, chained_data_delayed_13__11_, chained_data_delayed_13__10_, chained_data_delayed_13__9_, chained_data_delayed_13__8_, chained_data_delayed_13__7_, chained_data_delayed_13__6_, chained_data_delayed_13__5_, chained_data_delayed_13__4_, chained_data_delayed_13__3_, chained_data_delayed_13__2_, chained_data_delayed_13__1_, chained_data_delayed_13__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_14__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_13__127_, chained_data_delayed_13__126_, chained_data_delayed_13__125_, chained_data_delayed_13__124_, chained_data_delayed_13__123_, chained_data_delayed_13__122_, chained_data_delayed_13__121_, chained_data_delayed_13__120_, chained_data_delayed_13__119_, chained_data_delayed_13__118_, chained_data_delayed_13__117_, chained_data_delayed_13__116_, chained_data_delayed_13__115_, chained_data_delayed_13__114_, chained_data_delayed_13__113_, chained_data_delayed_13__112_, chained_data_delayed_13__111_, chained_data_delayed_13__110_, chained_data_delayed_13__109_, chained_data_delayed_13__108_, chained_data_delayed_13__107_, chained_data_delayed_13__106_, chained_data_delayed_13__105_, chained_data_delayed_13__104_, chained_data_delayed_13__103_, chained_data_delayed_13__102_, chained_data_delayed_13__101_, chained_data_delayed_13__100_, chained_data_delayed_13__99_, chained_data_delayed_13__98_, chained_data_delayed_13__97_, chained_data_delayed_13__96_, chained_data_delayed_13__95_, chained_data_delayed_13__94_, chained_data_delayed_13__93_, chained_data_delayed_13__92_, chained_data_delayed_13__91_, chained_data_delayed_13__90_, chained_data_delayed_13__89_, chained_data_delayed_13__88_, chained_data_delayed_13__87_, chained_data_delayed_13__86_, chained_data_delayed_13__85_, chained_data_delayed_13__84_, chained_data_delayed_13__83_, chained_data_delayed_13__82_, chained_data_delayed_13__81_, chained_data_delayed_13__80_, chained_data_delayed_13__79_, chained_data_delayed_13__78_, chained_data_delayed_13__77_, chained_data_delayed_13__76_, chained_data_delayed_13__75_, chained_data_delayed_13__74_, chained_data_delayed_13__73_, chained_data_delayed_13__72_, chained_data_delayed_13__71_, chained_data_delayed_13__70_, chained_data_delayed_13__69_, chained_data_delayed_13__68_, chained_data_delayed_13__67_, chained_data_delayed_13__66_, chained_data_delayed_13__65_, chained_data_delayed_13__64_, chained_data_delayed_13__63_, chained_data_delayed_13__62_, chained_data_delayed_13__61_, chained_data_delayed_13__60_, chained_data_delayed_13__59_, chained_data_delayed_13__58_, chained_data_delayed_13__57_, chained_data_delayed_13__56_, chained_data_delayed_13__55_, chained_data_delayed_13__54_, chained_data_delayed_13__53_, chained_data_delayed_13__52_, chained_data_delayed_13__51_, chained_data_delayed_13__50_, chained_data_delayed_13__49_, chained_data_delayed_13__48_, chained_data_delayed_13__47_, chained_data_delayed_13__46_, chained_data_delayed_13__45_, chained_data_delayed_13__44_, chained_data_delayed_13__43_, chained_data_delayed_13__42_, chained_data_delayed_13__41_, chained_data_delayed_13__40_, chained_data_delayed_13__39_, chained_data_delayed_13__38_, chained_data_delayed_13__37_, chained_data_delayed_13__36_, chained_data_delayed_13__35_, chained_data_delayed_13__34_, chained_data_delayed_13__33_, chained_data_delayed_13__32_, chained_data_delayed_13__31_, chained_data_delayed_13__30_, chained_data_delayed_13__29_, chained_data_delayed_13__28_, chained_data_delayed_13__27_, chained_data_delayed_13__26_, chained_data_delayed_13__25_, chained_data_delayed_13__24_, chained_data_delayed_13__23_, chained_data_delayed_13__22_, chained_data_delayed_13__21_, chained_data_delayed_13__20_, chained_data_delayed_13__19_, chained_data_delayed_13__18_, chained_data_delayed_13__17_, chained_data_delayed_13__16_, chained_data_delayed_13__15_, chained_data_delayed_13__14_, chained_data_delayed_13__13_, chained_data_delayed_13__12_, chained_data_delayed_13__11_, chained_data_delayed_13__10_, chained_data_delayed_13__9_, chained_data_delayed_13__8_, chained_data_delayed_13__7_, chained_data_delayed_13__6_, chained_data_delayed_13__5_, chained_data_delayed_13__4_, chained_data_delayed_13__3_, chained_data_delayed_13__2_, chained_data_delayed_13__1_, chained_data_delayed_13__0_ }),
    .data_o({ chained_data_delayed_14__127_, chained_data_delayed_14__126_, chained_data_delayed_14__125_, chained_data_delayed_14__124_, chained_data_delayed_14__123_, chained_data_delayed_14__122_, chained_data_delayed_14__121_, chained_data_delayed_14__120_, chained_data_delayed_14__119_, chained_data_delayed_14__118_, chained_data_delayed_14__117_, chained_data_delayed_14__116_, chained_data_delayed_14__115_, chained_data_delayed_14__114_, chained_data_delayed_14__113_, chained_data_delayed_14__112_, chained_data_delayed_14__111_, chained_data_delayed_14__110_, chained_data_delayed_14__109_, chained_data_delayed_14__108_, chained_data_delayed_14__107_, chained_data_delayed_14__106_, chained_data_delayed_14__105_, chained_data_delayed_14__104_, chained_data_delayed_14__103_, chained_data_delayed_14__102_, chained_data_delayed_14__101_, chained_data_delayed_14__100_, chained_data_delayed_14__99_, chained_data_delayed_14__98_, chained_data_delayed_14__97_, chained_data_delayed_14__96_, chained_data_delayed_14__95_, chained_data_delayed_14__94_, chained_data_delayed_14__93_, chained_data_delayed_14__92_, chained_data_delayed_14__91_, chained_data_delayed_14__90_, chained_data_delayed_14__89_, chained_data_delayed_14__88_, chained_data_delayed_14__87_, chained_data_delayed_14__86_, chained_data_delayed_14__85_, chained_data_delayed_14__84_, chained_data_delayed_14__83_, chained_data_delayed_14__82_, chained_data_delayed_14__81_, chained_data_delayed_14__80_, chained_data_delayed_14__79_, chained_data_delayed_14__78_, chained_data_delayed_14__77_, chained_data_delayed_14__76_, chained_data_delayed_14__75_, chained_data_delayed_14__74_, chained_data_delayed_14__73_, chained_data_delayed_14__72_, chained_data_delayed_14__71_, chained_data_delayed_14__70_, chained_data_delayed_14__69_, chained_data_delayed_14__68_, chained_data_delayed_14__67_, chained_data_delayed_14__66_, chained_data_delayed_14__65_, chained_data_delayed_14__64_, chained_data_delayed_14__63_, chained_data_delayed_14__62_, chained_data_delayed_14__61_, chained_data_delayed_14__60_, chained_data_delayed_14__59_, chained_data_delayed_14__58_, chained_data_delayed_14__57_, chained_data_delayed_14__56_, chained_data_delayed_14__55_, chained_data_delayed_14__54_, chained_data_delayed_14__53_, chained_data_delayed_14__52_, chained_data_delayed_14__51_, chained_data_delayed_14__50_, chained_data_delayed_14__49_, chained_data_delayed_14__48_, chained_data_delayed_14__47_, chained_data_delayed_14__46_, chained_data_delayed_14__45_, chained_data_delayed_14__44_, chained_data_delayed_14__43_, chained_data_delayed_14__42_, chained_data_delayed_14__41_, chained_data_delayed_14__40_, chained_data_delayed_14__39_, chained_data_delayed_14__38_, chained_data_delayed_14__37_, chained_data_delayed_14__36_, chained_data_delayed_14__35_, chained_data_delayed_14__34_, chained_data_delayed_14__33_, chained_data_delayed_14__32_, chained_data_delayed_14__31_, chained_data_delayed_14__30_, chained_data_delayed_14__29_, chained_data_delayed_14__28_, chained_data_delayed_14__27_, chained_data_delayed_14__26_, chained_data_delayed_14__25_, chained_data_delayed_14__24_, chained_data_delayed_14__23_, chained_data_delayed_14__22_, chained_data_delayed_14__21_, chained_data_delayed_14__20_, chained_data_delayed_14__19_, chained_data_delayed_14__18_, chained_data_delayed_14__17_, chained_data_delayed_14__16_, chained_data_delayed_14__15_, chained_data_delayed_14__14_, chained_data_delayed_14__13_, chained_data_delayed_14__12_, chained_data_delayed_14__11_, chained_data_delayed_14__10_, chained_data_delayed_14__9_, chained_data_delayed_14__8_, chained_data_delayed_14__7_, chained_data_delayed_14__6_, chained_data_delayed_14__5_, chained_data_delayed_14__4_, chained_data_delayed_14__3_, chained_data_delayed_14__2_, chained_data_delayed_14__1_, chained_data_delayed_14__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_15__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_14__127_, chained_data_delayed_14__126_, chained_data_delayed_14__125_, chained_data_delayed_14__124_, chained_data_delayed_14__123_, chained_data_delayed_14__122_, chained_data_delayed_14__121_, chained_data_delayed_14__120_, chained_data_delayed_14__119_, chained_data_delayed_14__118_, chained_data_delayed_14__117_, chained_data_delayed_14__116_, chained_data_delayed_14__115_, chained_data_delayed_14__114_, chained_data_delayed_14__113_, chained_data_delayed_14__112_, chained_data_delayed_14__111_, chained_data_delayed_14__110_, chained_data_delayed_14__109_, chained_data_delayed_14__108_, chained_data_delayed_14__107_, chained_data_delayed_14__106_, chained_data_delayed_14__105_, chained_data_delayed_14__104_, chained_data_delayed_14__103_, chained_data_delayed_14__102_, chained_data_delayed_14__101_, chained_data_delayed_14__100_, chained_data_delayed_14__99_, chained_data_delayed_14__98_, chained_data_delayed_14__97_, chained_data_delayed_14__96_, chained_data_delayed_14__95_, chained_data_delayed_14__94_, chained_data_delayed_14__93_, chained_data_delayed_14__92_, chained_data_delayed_14__91_, chained_data_delayed_14__90_, chained_data_delayed_14__89_, chained_data_delayed_14__88_, chained_data_delayed_14__87_, chained_data_delayed_14__86_, chained_data_delayed_14__85_, chained_data_delayed_14__84_, chained_data_delayed_14__83_, chained_data_delayed_14__82_, chained_data_delayed_14__81_, chained_data_delayed_14__80_, chained_data_delayed_14__79_, chained_data_delayed_14__78_, chained_data_delayed_14__77_, chained_data_delayed_14__76_, chained_data_delayed_14__75_, chained_data_delayed_14__74_, chained_data_delayed_14__73_, chained_data_delayed_14__72_, chained_data_delayed_14__71_, chained_data_delayed_14__70_, chained_data_delayed_14__69_, chained_data_delayed_14__68_, chained_data_delayed_14__67_, chained_data_delayed_14__66_, chained_data_delayed_14__65_, chained_data_delayed_14__64_, chained_data_delayed_14__63_, chained_data_delayed_14__62_, chained_data_delayed_14__61_, chained_data_delayed_14__60_, chained_data_delayed_14__59_, chained_data_delayed_14__58_, chained_data_delayed_14__57_, chained_data_delayed_14__56_, chained_data_delayed_14__55_, chained_data_delayed_14__54_, chained_data_delayed_14__53_, chained_data_delayed_14__52_, chained_data_delayed_14__51_, chained_data_delayed_14__50_, chained_data_delayed_14__49_, chained_data_delayed_14__48_, chained_data_delayed_14__47_, chained_data_delayed_14__46_, chained_data_delayed_14__45_, chained_data_delayed_14__44_, chained_data_delayed_14__43_, chained_data_delayed_14__42_, chained_data_delayed_14__41_, chained_data_delayed_14__40_, chained_data_delayed_14__39_, chained_data_delayed_14__38_, chained_data_delayed_14__37_, chained_data_delayed_14__36_, chained_data_delayed_14__35_, chained_data_delayed_14__34_, chained_data_delayed_14__33_, chained_data_delayed_14__32_, chained_data_delayed_14__31_, chained_data_delayed_14__30_, chained_data_delayed_14__29_, chained_data_delayed_14__28_, chained_data_delayed_14__27_, chained_data_delayed_14__26_, chained_data_delayed_14__25_, chained_data_delayed_14__24_, chained_data_delayed_14__23_, chained_data_delayed_14__22_, chained_data_delayed_14__21_, chained_data_delayed_14__20_, chained_data_delayed_14__19_, chained_data_delayed_14__18_, chained_data_delayed_14__17_, chained_data_delayed_14__16_, chained_data_delayed_14__15_, chained_data_delayed_14__14_, chained_data_delayed_14__13_, chained_data_delayed_14__12_, chained_data_delayed_14__11_, chained_data_delayed_14__10_, chained_data_delayed_14__9_, chained_data_delayed_14__8_, chained_data_delayed_14__7_, chained_data_delayed_14__6_, chained_data_delayed_14__5_, chained_data_delayed_14__4_, chained_data_delayed_14__3_, chained_data_delayed_14__2_, chained_data_delayed_14__1_, chained_data_delayed_14__0_ }),
    .data_o({ chained_data_delayed_15__127_, chained_data_delayed_15__126_, chained_data_delayed_15__125_, chained_data_delayed_15__124_, chained_data_delayed_15__123_, chained_data_delayed_15__122_, chained_data_delayed_15__121_, chained_data_delayed_15__120_, chained_data_delayed_15__119_, chained_data_delayed_15__118_, chained_data_delayed_15__117_, chained_data_delayed_15__116_, chained_data_delayed_15__115_, chained_data_delayed_15__114_, chained_data_delayed_15__113_, chained_data_delayed_15__112_, chained_data_delayed_15__111_, chained_data_delayed_15__110_, chained_data_delayed_15__109_, chained_data_delayed_15__108_, chained_data_delayed_15__107_, chained_data_delayed_15__106_, chained_data_delayed_15__105_, chained_data_delayed_15__104_, chained_data_delayed_15__103_, chained_data_delayed_15__102_, chained_data_delayed_15__101_, chained_data_delayed_15__100_, chained_data_delayed_15__99_, chained_data_delayed_15__98_, chained_data_delayed_15__97_, chained_data_delayed_15__96_, chained_data_delayed_15__95_, chained_data_delayed_15__94_, chained_data_delayed_15__93_, chained_data_delayed_15__92_, chained_data_delayed_15__91_, chained_data_delayed_15__90_, chained_data_delayed_15__89_, chained_data_delayed_15__88_, chained_data_delayed_15__87_, chained_data_delayed_15__86_, chained_data_delayed_15__85_, chained_data_delayed_15__84_, chained_data_delayed_15__83_, chained_data_delayed_15__82_, chained_data_delayed_15__81_, chained_data_delayed_15__80_, chained_data_delayed_15__79_, chained_data_delayed_15__78_, chained_data_delayed_15__77_, chained_data_delayed_15__76_, chained_data_delayed_15__75_, chained_data_delayed_15__74_, chained_data_delayed_15__73_, chained_data_delayed_15__72_, chained_data_delayed_15__71_, chained_data_delayed_15__70_, chained_data_delayed_15__69_, chained_data_delayed_15__68_, chained_data_delayed_15__67_, chained_data_delayed_15__66_, chained_data_delayed_15__65_, chained_data_delayed_15__64_, chained_data_delayed_15__63_, chained_data_delayed_15__62_, chained_data_delayed_15__61_, chained_data_delayed_15__60_, chained_data_delayed_15__59_, chained_data_delayed_15__58_, chained_data_delayed_15__57_, chained_data_delayed_15__56_, chained_data_delayed_15__55_, chained_data_delayed_15__54_, chained_data_delayed_15__53_, chained_data_delayed_15__52_, chained_data_delayed_15__51_, chained_data_delayed_15__50_, chained_data_delayed_15__49_, chained_data_delayed_15__48_, chained_data_delayed_15__47_, chained_data_delayed_15__46_, chained_data_delayed_15__45_, chained_data_delayed_15__44_, chained_data_delayed_15__43_, chained_data_delayed_15__42_, chained_data_delayed_15__41_, chained_data_delayed_15__40_, chained_data_delayed_15__39_, chained_data_delayed_15__38_, chained_data_delayed_15__37_, chained_data_delayed_15__36_, chained_data_delayed_15__35_, chained_data_delayed_15__34_, chained_data_delayed_15__33_, chained_data_delayed_15__32_, chained_data_delayed_15__31_, chained_data_delayed_15__30_, chained_data_delayed_15__29_, chained_data_delayed_15__28_, chained_data_delayed_15__27_, chained_data_delayed_15__26_, chained_data_delayed_15__25_, chained_data_delayed_15__24_, chained_data_delayed_15__23_, chained_data_delayed_15__22_, chained_data_delayed_15__21_, chained_data_delayed_15__20_, chained_data_delayed_15__19_, chained_data_delayed_15__18_, chained_data_delayed_15__17_, chained_data_delayed_15__16_, chained_data_delayed_15__15_, chained_data_delayed_15__14_, chained_data_delayed_15__13_, chained_data_delayed_15__12_, chained_data_delayed_15__11_, chained_data_delayed_15__10_, chained_data_delayed_15__9_, chained_data_delayed_15__8_, chained_data_delayed_15__7_, chained_data_delayed_15__6_, chained_data_delayed_15__5_, chained_data_delayed_15__4_, chained_data_delayed_15__3_, chained_data_delayed_15__2_, chained_data_delayed_15__1_, chained_data_delayed_15__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_16__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_15__127_, chained_data_delayed_15__126_, chained_data_delayed_15__125_, chained_data_delayed_15__124_, chained_data_delayed_15__123_, chained_data_delayed_15__122_, chained_data_delayed_15__121_, chained_data_delayed_15__120_, chained_data_delayed_15__119_, chained_data_delayed_15__118_, chained_data_delayed_15__117_, chained_data_delayed_15__116_, chained_data_delayed_15__115_, chained_data_delayed_15__114_, chained_data_delayed_15__113_, chained_data_delayed_15__112_, chained_data_delayed_15__111_, chained_data_delayed_15__110_, chained_data_delayed_15__109_, chained_data_delayed_15__108_, chained_data_delayed_15__107_, chained_data_delayed_15__106_, chained_data_delayed_15__105_, chained_data_delayed_15__104_, chained_data_delayed_15__103_, chained_data_delayed_15__102_, chained_data_delayed_15__101_, chained_data_delayed_15__100_, chained_data_delayed_15__99_, chained_data_delayed_15__98_, chained_data_delayed_15__97_, chained_data_delayed_15__96_, chained_data_delayed_15__95_, chained_data_delayed_15__94_, chained_data_delayed_15__93_, chained_data_delayed_15__92_, chained_data_delayed_15__91_, chained_data_delayed_15__90_, chained_data_delayed_15__89_, chained_data_delayed_15__88_, chained_data_delayed_15__87_, chained_data_delayed_15__86_, chained_data_delayed_15__85_, chained_data_delayed_15__84_, chained_data_delayed_15__83_, chained_data_delayed_15__82_, chained_data_delayed_15__81_, chained_data_delayed_15__80_, chained_data_delayed_15__79_, chained_data_delayed_15__78_, chained_data_delayed_15__77_, chained_data_delayed_15__76_, chained_data_delayed_15__75_, chained_data_delayed_15__74_, chained_data_delayed_15__73_, chained_data_delayed_15__72_, chained_data_delayed_15__71_, chained_data_delayed_15__70_, chained_data_delayed_15__69_, chained_data_delayed_15__68_, chained_data_delayed_15__67_, chained_data_delayed_15__66_, chained_data_delayed_15__65_, chained_data_delayed_15__64_, chained_data_delayed_15__63_, chained_data_delayed_15__62_, chained_data_delayed_15__61_, chained_data_delayed_15__60_, chained_data_delayed_15__59_, chained_data_delayed_15__58_, chained_data_delayed_15__57_, chained_data_delayed_15__56_, chained_data_delayed_15__55_, chained_data_delayed_15__54_, chained_data_delayed_15__53_, chained_data_delayed_15__52_, chained_data_delayed_15__51_, chained_data_delayed_15__50_, chained_data_delayed_15__49_, chained_data_delayed_15__48_, chained_data_delayed_15__47_, chained_data_delayed_15__46_, chained_data_delayed_15__45_, chained_data_delayed_15__44_, chained_data_delayed_15__43_, chained_data_delayed_15__42_, chained_data_delayed_15__41_, chained_data_delayed_15__40_, chained_data_delayed_15__39_, chained_data_delayed_15__38_, chained_data_delayed_15__37_, chained_data_delayed_15__36_, chained_data_delayed_15__35_, chained_data_delayed_15__34_, chained_data_delayed_15__33_, chained_data_delayed_15__32_, chained_data_delayed_15__31_, chained_data_delayed_15__30_, chained_data_delayed_15__29_, chained_data_delayed_15__28_, chained_data_delayed_15__27_, chained_data_delayed_15__26_, chained_data_delayed_15__25_, chained_data_delayed_15__24_, chained_data_delayed_15__23_, chained_data_delayed_15__22_, chained_data_delayed_15__21_, chained_data_delayed_15__20_, chained_data_delayed_15__19_, chained_data_delayed_15__18_, chained_data_delayed_15__17_, chained_data_delayed_15__16_, chained_data_delayed_15__15_, chained_data_delayed_15__14_, chained_data_delayed_15__13_, chained_data_delayed_15__12_, chained_data_delayed_15__11_, chained_data_delayed_15__10_, chained_data_delayed_15__9_, chained_data_delayed_15__8_, chained_data_delayed_15__7_, chained_data_delayed_15__6_, chained_data_delayed_15__5_, chained_data_delayed_15__4_, chained_data_delayed_15__3_, chained_data_delayed_15__2_, chained_data_delayed_15__1_, chained_data_delayed_15__0_ }),
    .data_o({ chained_data_delayed_16__127_, chained_data_delayed_16__126_, chained_data_delayed_16__125_, chained_data_delayed_16__124_, chained_data_delayed_16__123_, chained_data_delayed_16__122_, chained_data_delayed_16__121_, chained_data_delayed_16__120_, chained_data_delayed_16__119_, chained_data_delayed_16__118_, chained_data_delayed_16__117_, chained_data_delayed_16__116_, chained_data_delayed_16__115_, chained_data_delayed_16__114_, chained_data_delayed_16__113_, chained_data_delayed_16__112_, chained_data_delayed_16__111_, chained_data_delayed_16__110_, chained_data_delayed_16__109_, chained_data_delayed_16__108_, chained_data_delayed_16__107_, chained_data_delayed_16__106_, chained_data_delayed_16__105_, chained_data_delayed_16__104_, chained_data_delayed_16__103_, chained_data_delayed_16__102_, chained_data_delayed_16__101_, chained_data_delayed_16__100_, chained_data_delayed_16__99_, chained_data_delayed_16__98_, chained_data_delayed_16__97_, chained_data_delayed_16__96_, chained_data_delayed_16__95_, chained_data_delayed_16__94_, chained_data_delayed_16__93_, chained_data_delayed_16__92_, chained_data_delayed_16__91_, chained_data_delayed_16__90_, chained_data_delayed_16__89_, chained_data_delayed_16__88_, chained_data_delayed_16__87_, chained_data_delayed_16__86_, chained_data_delayed_16__85_, chained_data_delayed_16__84_, chained_data_delayed_16__83_, chained_data_delayed_16__82_, chained_data_delayed_16__81_, chained_data_delayed_16__80_, chained_data_delayed_16__79_, chained_data_delayed_16__78_, chained_data_delayed_16__77_, chained_data_delayed_16__76_, chained_data_delayed_16__75_, chained_data_delayed_16__74_, chained_data_delayed_16__73_, chained_data_delayed_16__72_, chained_data_delayed_16__71_, chained_data_delayed_16__70_, chained_data_delayed_16__69_, chained_data_delayed_16__68_, chained_data_delayed_16__67_, chained_data_delayed_16__66_, chained_data_delayed_16__65_, chained_data_delayed_16__64_, chained_data_delayed_16__63_, chained_data_delayed_16__62_, chained_data_delayed_16__61_, chained_data_delayed_16__60_, chained_data_delayed_16__59_, chained_data_delayed_16__58_, chained_data_delayed_16__57_, chained_data_delayed_16__56_, chained_data_delayed_16__55_, chained_data_delayed_16__54_, chained_data_delayed_16__53_, chained_data_delayed_16__52_, chained_data_delayed_16__51_, chained_data_delayed_16__50_, chained_data_delayed_16__49_, chained_data_delayed_16__48_, chained_data_delayed_16__47_, chained_data_delayed_16__46_, chained_data_delayed_16__45_, chained_data_delayed_16__44_, chained_data_delayed_16__43_, chained_data_delayed_16__42_, chained_data_delayed_16__41_, chained_data_delayed_16__40_, chained_data_delayed_16__39_, chained_data_delayed_16__38_, chained_data_delayed_16__37_, chained_data_delayed_16__36_, chained_data_delayed_16__35_, chained_data_delayed_16__34_, chained_data_delayed_16__33_, chained_data_delayed_16__32_, chained_data_delayed_16__31_, chained_data_delayed_16__30_, chained_data_delayed_16__29_, chained_data_delayed_16__28_, chained_data_delayed_16__27_, chained_data_delayed_16__26_, chained_data_delayed_16__25_, chained_data_delayed_16__24_, chained_data_delayed_16__23_, chained_data_delayed_16__22_, chained_data_delayed_16__21_, chained_data_delayed_16__20_, chained_data_delayed_16__19_, chained_data_delayed_16__18_, chained_data_delayed_16__17_, chained_data_delayed_16__16_, chained_data_delayed_16__15_, chained_data_delayed_16__14_, chained_data_delayed_16__13_, chained_data_delayed_16__12_, chained_data_delayed_16__11_, chained_data_delayed_16__10_, chained_data_delayed_16__9_, chained_data_delayed_16__8_, chained_data_delayed_16__7_, chained_data_delayed_16__6_, chained_data_delayed_16__5_, chained_data_delayed_16__4_, chained_data_delayed_16__3_, chained_data_delayed_16__2_, chained_data_delayed_16__1_, chained_data_delayed_16__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_17__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_16__127_, chained_data_delayed_16__126_, chained_data_delayed_16__125_, chained_data_delayed_16__124_, chained_data_delayed_16__123_, chained_data_delayed_16__122_, chained_data_delayed_16__121_, chained_data_delayed_16__120_, chained_data_delayed_16__119_, chained_data_delayed_16__118_, chained_data_delayed_16__117_, chained_data_delayed_16__116_, chained_data_delayed_16__115_, chained_data_delayed_16__114_, chained_data_delayed_16__113_, chained_data_delayed_16__112_, chained_data_delayed_16__111_, chained_data_delayed_16__110_, chained_data_delayed_16__109_, chained_data_delayed_16__108_, chained_data_delayed_16__107_, chained_data_delayed_16__106_, chained_data_delayed_16__105_, chained_data_delayed_16__104_, chained_data_delayed_16__103_, chained_data_delayed_16__102_, chained_data_delayed_16__101_, chained_data_delayed_16__100_, chained_data_delayed_16__99_, chained_data_delayed_16__98_, chained_data_delayed_16__97_, chained_data_delayed_16__96_, chained_data_delayed_16__95_, chained_data_delayed_16__94_, chained_data_delayed_16__93_, chained_data_delayed_16__92_, chained_data_delayed_16__91_, chained_data_delayed_16__90_, chained_data_delayed_16__89_, chained_data_delayed_16__88_, chained_data_delayed_16__87_, chained_data_delayed_16__86_, chained_data_delayed_16__85_, chained_data_delayed_16__84_, chained_data_delayed_16__83_, chained_data_delayed_16__82_, chained_data_delayed_16__81_, chained_data_delayed_16__80_, chained_data_delayed_16__79_, chained_data_delayed_16__78_, chained_data_delayed_16__77_, chained_data_delayed_16__76_, chained_data_delayed_16__75_, chained_data_delayed_16__74_, chained_data_delayed_16__73_, chained_data_delayed_16__72_, chained_data_delayed_16__71_, chained_data_delayed_16__70_, chained_data_delayed_16__69_, chained_data_delayed_16__68_, chained_data_delayed_16__67_, chained_data_delayed_16__66_, chained_data_delayed_16__65_, chained_data_delayed_16__64_, chained_data_delayed_16__63_, chained_data_delayed_16__62_, chained_data_delayed_16__61_, chained_data_delayed_16__60_, chained_data_delayed_16__59_, chained_data_delayed_16__58_, chained_data_delayed_16__57_, chained_data_delayed_16__56_, chained_data_delayed_16__55_, chained_data_delayed_16__54_, chained_data_delayed_16__53_, chained_data_delayed_16__52_, chained_data_delayed_16__51_, chained_data_delayed_16__50_, chained_data_delayed_16__49_, chained_data_delayed_16__48_, chained_data_delayed_16__47_, chained_data_delayed_16__46_, chained_data_delayed_16__45_, chained_data_delayed_16__44_, chained_data_delayed_16__43_, chained_data_delayed_16__42_, chained_data_delayed_16__41_, chained_data_delayed_16__40_, chained_data_delayed_16__39_, chained_data_delayed_16__38_, chained_data_delayed_16__37_, chained_data_delayed_16__36_, chained_data_delayed_16__35_, chained_data_delayed_16__34_, chained_data_delayed_16__33_, chained_data_delayed_16__32_, chained_data_delayed_16__31_, chained_data_delayed_16__30_, chained_data_delayed_16__29_, chained_data_delayed_16__28_, chained_data_delayed_16__27_, chained_data_delayed_16__26_, chained_data_delayed_16__25_, chained_data_delayed_16__24_, chained_data_delayed_16__23_, chained_data_delayed_16__22_, chained_data_delayed_16__21_, chained_data_delayed_16__20_, chained_data_delayed_16__19_, chained_data_delayed_16__18_, chained_data_delayed_16__17_, chained_data_delayed_16__16_, chained_data_delayed_16__15_, chained_data_delayed_16__14_, chained_data_delayed_16__13_, chained_data_delayed_16__12_, chained_data_delayed_16__11_, chained_data_delayed_16__10_, chained_data_delayed_16__9_, chained_data_delayed_16__8_, chained_data_delayed_16__7_, chained_data_delayed_16__6_, chained_data_delayed_16__5_, chained_data_delayed_16__4_, chained_data_delayed_16__3_, chained_data_delayed_16__2_, chained_data_delayed_16__1_, chained_data_delayed_16__0_ }),
    .data_o({ chained_data_delayed_17__127_, chained_data_delayed_17__126_, chained_data_delayed_17__125_, chained_data_delayed_17__124_, chained_data_delayed_17__123_, chained_data_delayed_17__122_, chained_data_delayed_17__121_, chained_data_delayed_17__120_, chained_data_delayed_17__119_, chained_data_delayed_17__118_, chained_data_delayed_17__117_, chained_data_delayed_17__116_, chained_data_delayed_17__115_, chained_data_delayed_17__114_, chained_data_delayed_17__113_, chained_data_delayed_17__112_, chained_data_delayed_17__111_, chained_data_delayed_17__110_, chained_data_delayed_17__109_, chained_data_delayed_17__108_, chained_data_delayed_17__107_, chained_data_delayed_17__106_, chained_data_delayed_17__105_, chained_data_delayed_17__104_, chained_data_delayed_17__103_, chained_data_delayed_17__102_, chained_data_delayed_17__101_, chained_data_delayed_17__100_, chained_data_delayed_17__99_, chained_data_delayed_17__98_, chained_data_delayed_17__97_, chained_data_delayed_17__96_, chained_data_delayed_17__95_, chained_data_delayed_17__94_, chained_data_delayed_17__93_, chained_data_delayed_17__92_, chained_data_delayed_17__91_, chained_data_delayed_17__90_, chained_data_delayed_17__89_, chained_data_delayed_17__88_, chained_data_delayed_17__87_, chained_data_delayed_17__86_, chained_data_delayed_17__85_, chained_data_delayed_17__84_, chained_data_delayed_17__83_, chained_data_delayed_17__82_, chained_data_delayed_17__81_, chained_data_delayed_17__80_, chained_data_delayed_17__79_, chained_data_delayed_17__78_, chained_data_delayed_17__77_, chained_data_delayed_17__76_, chained_data_delayed_17__75_, chained_data_delayed_17__74_, chained_data_delayed_17__73_, chained_data_delayed_17__72_, chained_data_delayed_17__71_, chained_data_delayed_17__70_, chained_data_delayed_17__69_, chained_data_delayed_17__68_, chained_data_delayed_17__67_, chained_data_delayed_17__66_, chained_data_delayed_17__65_, chained_data_delayed_17__64_, chained_data_delayed_17__63_, chained_data_delayed_17__62_, chained_data_delayed_17__61_, chained_data_delayed_17__60_, chained_data_delayed_17__59_, chained_data_delayed_17__58_, chained_data_delayed_17__57_, chained_data_delayed_17__56_, chained_data_delayed_17__55_, chained_data_delayed_17__54_, chained_data_delayed_17__53_, chained_data_delayed_17__52_, chained_data_delayed_17__51_, chained_data_delayed_17__50_, chained_data_delayed_17__49_, chained_data_delayed_17__48_, chained_data_delayed_17__47_, chained_data_delayed_17__46_, chained_data_delayed_17__45_, chained_data_delayed_17__44_, chained_data_delayed_17__43_, chained_data_delayed_17__42_, chained_data_delayed_17__41_, chained_data_delayed_17__40_, chained_data_delayed_17__39_, chained_data_delayed_17__38_, chained_data_delayed_17__37_, chained_data_delayed_17__36_, chained_data_delayed_17__35_, chained_data_delayed_17__34_, chained_data_delayed_17__33_, chained_data_delayed_17__32_, chained_data_delayed_17__31_, chained_data_delayed_17__30_, chained_data_delayed_17__29_, chained_data_delayed_17__28_, chained_data_delayed_17__27_, chained_data_delayed_17__26_, chained_data_delayed_17__25_, chained_data_delayed_17__24_, chained_data_delayed_17__23_, chained_data_delayed_17__22_, chained_data_delayed_17__21_, chained_data_delayed_17__20_, chained_data_delayed_17__19_, chained_data_delayed_17__18_, chained_data_delayed_17__17_, chained_data_delayed_17__16_, chained_data_delayed_17__15_, chained_data_delayed_17__14_, chained_data_delayed_17__13_, chained_data_delayed_17__12_, chained_data_delayed_17__11_, chained_data_delayed_17__10_, chained_data_delayed_17__9_, chained_data_delayed_17__8_, chained_data_delayed_17__7_, chained_data_delayed_17__6_, chained_data_delayed_17__5_, chained_data_delayed_17__4_, chained_data_delayed_17__3_, chained_data_delayed_17__2_, chained_data_delayed_17__1_, chained_data_delayed_17__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_18__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_17__127_, chained_data_delayed_17__126_, chained_data_delayed_17__125_, chained_data_delayed_17__124_, chained_data_delayed_17__123_, chained_data_delayed_17__122_, chained_data_delayed_17__121_, chained_data_delayed_17__120_, chained_data_delayed_17__119_, chained_data_delayed_17__118_, chained_data_delayed_17__117_, chained_data_delayed_17__116_, chained_data_delayed_17__115_, chained_data_delayed_17__114_, chained_data_delayed_17__113_, chained_data_delayed_17__112_, chained_data_delayed_17__111_, chained_data_delayed_17__110_, chained_data_delayed_17__109_, chained_data_delayed_17__108_, chained_data_delayed_17__107_, chained_data_delayed_17__106_, chained_data_delayed_17__105_, chained_data_delayed_17__104_, chained_data_delayed_17__103_, chained_data_delayed_17__102_, chained_data_delayed_17__101_, chained_data_delayed_17__100_, chained_data_delayed_17__99_, chained_data_delayed_17__98_, chained_data_delayed_17__97_, chained_data_delayed_17__96_, chained_data_delayed_17__95_, chained_data_delayed_17__94_, chained_data_delayed_17__93_, chained_data_delayed_17__92_, chained_data_delayed_17__91_, chained_data_delayed_17__90_, chained_data_delayed_17__89_, chained_data_delayed_17__88_, chained_data_delayed_17__87_, chained_data_delayed_17__86_, chained_data_delayed_17__85_, chained_data_delayed_17__84_, chained_data_delayed_17__83_, chained_data_delayed_17__82_, chained_data_delayed_17__81_, chained_data_delayed_17__80_, chained_data_delayed_17__79_, chained_data_delayed_17__78_, chained_data_delayed_17__77_, chained_data_delayed_17__76_, chained_data_delayed_17__75_, chained_data_delayed_17__74_, chained_data_delayed_17__73_, chained_data_delayed_17__72_, chained_data_delayed_17__71_, chained_data_delayed_17__70_, chained_data_delayed_17__69_, chained_data_delayed_17__68_, chained_data_delayed_17__67_, chained_data_delayed_17__66_, chained_data_delayed_17__65_, chained_data_delayed_17__64_, chained_data_delayed_17__63_, chained_data_delayed_17__62_, chained_data_delayed_17__61_, chained_data_delayed_17__60_, chained_data_delayed_17__59_, chained_data_delayed_17__58_, chained_data_delayed_17__57_, chained_data_delayed_17__56_, chained_data_delayed_17__55_, chained_data_delayed_17__54_, chained_data_delayed_17__53_, chained_data_delayed_17__52_, chained_data_delayed_17__51_, chained_data_delayed_17__50_, chained_data_delayed_17__49_, chained_data_delayed_17__48_, chained_data_delayed_17__47_, chained_data_delayed_17__46_, chained_data_delayed_17__45_, chained_data_delayed_17__44_, chained_data_delayed_17__43_, chained_data_delayed_17__42_, chained_data_delayed_17__41_, chained_data_delayed_17__40_, chained_data_delayed_17__39_, chained_data_delayed_17__38_, chained_data_delayed_17__37_, chained_data_delayed_17__36_, chained_data_delayed_17__35_, chained_data_delayed_17__34_, chained_data_delayed_17__33_, chained_data_delayed_17__32_, chained_data_delayed_17__31_, chained_data_delayed_17__30_, chained_data_delayed_17__29_, chained_data_delayed_17__28_, chained_data_delayed_17__27_, chained_data_delayed_17__26_, chained_data_delayed_17__25_, chained_data_delayed_17__24_, chained_data_delayed_17__23_, chained_data_delayed_17__22_, chained_data_delayed_17__21_, chained_data_delayed_17__20_, chained_data_delayed_17__19_, chained_data_delayed_17__18_, chained_data_delayed_17__17_, chained_data_delayed_17__16_, chained_data_delayed_17__15_, chained_data_delayed_17__14_, chained_data_delayed_17__13_, chained_data_delayed_17__12_, chained_data_delayed_17__11_, chained_data_delayed_17__10_, chained_data_delayed_17__9_, chained_data_delayed_17__8_, chained_data_delayed_17__7_, chained_data_delayed_17__6_, chained_data_delayed_17__5_, chained_data_delayed_17__4_, chained_data_delayed_17__3_, chained_data_delayed_17__2_, chained_data_delayed_17__1_, chained_data_delayed_17__0_ }),
    .data_o({ chained_data_delayed_18__127_, chained_data_delayed_18__126_, chained_data_delayed_18__125_, chained_data_delayed_18__124_, chained_data_delayed_18__123_, chained_data_delayed_18__122_, chained_data_delayed_18__121_, chained_data_delayed_18__120_, chained_data_delayed_18__119_, chained_data_delayed_18__118_, chained_data_delayed_18__117_, chained_data_delayed_18__116_, chained_data_delayed_18__115_, chained_data_delayed_18__114_, chained_data_delayed_18__113_, chained_data_delayed_18__112_, chained_data_delayed_18__111_, chained_data_delayed_18__110_, chained_data_delayed_18__109_, chained_data_delayed_18__108_, chained_data_delayed_18__107_, chained_data_delayed_18__106_, chained_data_delayed_18__105_, chained_data_delayed_18__104_, chained_data_delayed_18__103_, chained_data_delayed_18__102_, chained_data_delayed_18__101_, chained_data_delayed_18__100_, chained_data_delayed_18__99_, chained_data_delayed_18__98_, chained_data_delayed_18__97_, chained_data_delayed_18__96_, chained_data_delayed_18__95_, chained_data_delayed_18__94_, chained_data_delayed_18__93_, chained_data_delayed_18__92_, chained_data_delayed_18__91_, chained_data_delayed_18__90_, chained_data_delayed_18__89_, chained_data_delayed_18__88_, chained_data_delayed_18__87_, chained_data_delayed_18__86_, chained_data_delayed_18__85_, chained_data_delayed_18__84_, chained_data_delayed_18__83_, chained_data_delayed_18__82_, chained_data_delayed_18__81_, chained_data_delayed_18__80_, chained_data_delayed_18__79_, chained_data_delayed_18__78_, chained_data_delayed_18__77_, chained_data_delayed_18__76_, chained_data_delayed_18__75_, chained_data_delayed_18__74_, chained_data_delayed_18__73_, chained_data_delayed_18__72_, chained_data_delayed_18__71_, chained_data_delayed_18__70_, chained_data_delayed_18__69_, chained_data_delayed_18__68_, chained_data_delayed_18__67_, chained_data_delayed_18__66_, chained_data_delayed_18__65_, chained_data_delayed_18__64_, chained_data_delayed_18__63_, chained_data_delayed_18__62_, chained_data_delayed_18__61_, chained_data_delayed_18__60_, chained_data_delayed_18__59_, chained_data_delayed_18__58_, chained_data_delayed_18__57_, chained_data_delayed_18__56_, chained_data_delayed_18__55_, chained_data_delayed_18__54_, chained_data_delayed_18__53_, chained_data_delayed_18__52_, chained_data_delayed_18__51_, chained_data_delayed_18__50_, chained_data_delayed_18__49_, chained_data_delayed_18__48_, chained_data_delayed_18__47_, chained_data_delayed_18__46_, chained_data_delayed_18__45_, chained_data_delayed_18__44_, chained_data_delayed_18__43_, chained_data_delayed_18__42_, chained_data_delayed_18__41_, chained_data_delayed_18__40_, chained_data_delayed_18__39_, chained_data_delayed_18__38_, chained_data_delayed_18__37_, chained_data_delayed_18__36_, chained_data_delayed_18__35_, chained_data_delayed_18__34_, chained_data_delayed_18__33_, chained_data_delayed_18__32_, chained_data_delayed_18__31_, chained_data_delayed_18__30_, chained_data_delayed_18__29_, chained_data_delayed_18__28_, chained_data_delayed_18__27_, chained_data_delayed_18__26_, chained_data_delayed_18__25_, chained_data_delayed_18__24_, chained_data_delayed_18__23_, chained_data_delayed_18__22_, chained_data_delayed_18__21_, chained_data_delayed_18__20_, chained_data_delayed_18__19_, chained_data_delayed_18__18_, chained_data_delayed_18__17_, chained_data_delayed_18__16_, chained_data_delayed_18__15_, chained_data_delayed_18__14_, chained_data_delayed_18__13_, chained_data_delayed_18__12_, chained_data_delayed_18__11_, chained_data_delayed_18__10_, chained_data_delayed_18__9_, chained_data_delayed_18__8_, chained_data_delayed_18__7_, chained_data_delayed_18__6_, chained_data_delayed_18__5_, chained_data_delayed_18__4_, chained_data_delayed_18__3_, chained_data_delayed_18__2_, chained_data_delayed_18__1_, chained_data_delayed_18__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_19__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_18__127_, chained_data_delayed_18__126_, chained_data_delayed_18__125_, chained_data_delayed_18__124_, chained_data_delayed_18__123_, chained_data_delayed_18__122_, chained_data_delayed_18__121_, chained_data_delayed_18__120_, chained_data_delayed_18__119_, chained_data_delayed_18__118_, chained_data_delayed_18__117_, chained_data_delayed_18__116_, chained_data_delayed_18__115_, chained_data_delayed_18__114_, chained_data_delayed_18__113_, chained_data_delayed_18__112_, chained_data_delayed_18__111_, chained_data_delayed_18__110_, chained_data_delayed_18__109_, chained_data_delayed_18__108_, chained_data_delayed_18__107_, chained_data_delayed_18__106_, chained_data_delayed_18__105_, chained_data_delayed_18__104_, chained_data_delayed_18__103_, chained_data_delayed_18__102_, chained_data_delayed_18__101_, chained_data_delayed_18__100_, chained_data_delayed_18__99_, chained_data_delayed_18__98_, chained_data_delayed_18__97_, chained_data_delayed_18__96_, chained_data_delayed_18__95_, chained_data_delayed_18__94_, chained_data_delayed_18__93_, chained_data_delayed_18__92_, chained_data_delayed_18__91_, chained_data_delayed_18__90_, chained_data_delayed_18__89_, chained_data_delayed_18__88_, chained_data_delayed_18__87_, chained_data_delayed_18__86_, chained_data_delayed_18__85_, chained_data_delayed_18__84_, chained_data_delayed_18__83_, chained_data_delayed_18__82_, chained_data_delayed_18__81_, chained_data_delayed_18__80_, chained_data_delayed_18__79_, chained_data_delayed_18__78_, chained_data_delayed_18__77_, chained_data_delayed_18__76_, chained_data_delayed_18__75_, chained_data_delayed_18__74_, chained_data_delayed_18__73_, chained_data_delayed_18__72_, chained_data_delayed_18__71_, chained_data_delayed_18__70_, chained_data_delayed_18__69_, chained_data_delayed_18__68_, chained_data_delayed_18__67_, chained_data_delayed_18__66_, chained_data_delayed_18__65_, chained_data_delayed_18__64_, chained_data_delayed_18__63_, chained_data_delayed_18__62_, chained_data_delayed_18__61_, chained_data_delayed_18__60_, chained_data_delayed_18__59_, chained_data_delayed_18__58_, chained_data_delayed_18__57_, chained_data_delayed_18__56_, chained_data_delayed_18__55_, chained_data_delayed_18__54_, chained_data_delayed_18__53_, chained_data_delayed_18__52_, chained_data_delayed_18__51_, chained_data_delayed_18__50_, chained_data_delayed_18__49_, chained_data_delayed_18__48_, chained_data_delayed_18__47_, chained_data_delayed_18__46_, chained_data_delayed_18__45_, chained_data_delayed_18__44_, chained_data_delayed_18__43_, chained_data_delayed_18__42_, chained_data_delayed_18__41_, chained_data_delayed_18__40_, chained_data_delayed_18__39_, chained_data_delayed_18__38_, chained_data_delayed_18__37_, chained_data_delayed_18__36_, chained_data_delayed_18__35_, chained_data_delayed_18__34_, chained_data_delayed_18__33_, chained_data_delayed_18__32_, chained_data_delayed_18__31_, chained_data_delayed_18__30_, chained_data_delayed_18__29_, chained_data_delayed_18__28_, chained_data_delayed_18__27_, chained_data_delayed_18__26_, chained_data_delayed_18__25_, chained_data_delayed_18__24_, chained_data_delayed_18__23_, chained_data_delayed_18__22_, chained_data_delayed_18__21_, chained_data_delayed_18__20_, chained_data_delayed_18__19_, chained_data_delayed_18__18_, chained_data_delayed_18__17_, chained_data_delayed_18__16_, chained_data_delayed_18__15_, chained_data_delayed_18__14_, chained_data_delayed_18__13_, chained_data_delayed_18__12_, chained_data_delayed_18__11_, chained_data_delayed_18__10_, chained_data_delayed_18__9_, chained_data_delayed_18__8_, chained_data_delayed_18__7_, chained_data_delayed_18__6_, chained_data_delayed_18__5_, chained_data_delayed_18__4_, chained_data_delayed_18__3_, chained_data_delayed_18__2_, chained_data_delayed_18__1_, chained_data_delayed_18__0_ }),
    .data_o({ chained_data_delayed_19__127_, chained_data_delayed_19__126_, chained_data_delayed_19__125_, chained_data_delayed_19__124_, chained_data_delayed_19__123_, chained_data_delayed_19__122_, chained_data_delayed_19__121_, chained_data_delayed_19__120_, chained_data_delayed_19__119_, chained_data_delayed_19__118_, chained_data_delayed_19__117_, chained_data_delayed_19__116_, chained_data_delayed_19__115_, chained_data_delayed_19__114_, chained_data_delayed_19__113_, chained_data_delayed_19__112_, chained_data_delayed_19__111_, chained_data_delayed_19__110_, chained_data_delayed_19__109_, chained_data_delayed_19__108_, chained_data_delayed_19__107_, chained_data_delayed_19__106_, chained_data_delayed_19__105_, chained_data_delayed_19__104_, chained_data_delayed_19__103_, chained_data_delayed_19__102_, chained_data_delayed_19__101_, chained_data_delayed_19__100_, chained_data_delayed_19__99_, chained_data_delayed_19__98_, chained_data_delayed_19__97_, chained_data_delayed_19__96_, chained_data_delayed_19__95_, chained_data_delayed_19__94_, chained_data_delayed_19__93_, chained_data_delayed_19__92_, chained_data_delayed_19__91_, chained_data_delayed_19__90_, chained_data_delayed_19__89_, chained_data_delayed_19__88_, chained_data_delayed_19__87_, chained_data_delayed_19__86_, chained_data_delayed_19__85_, chained_data_delayed_19__84_, chained_data_delayed_19__83_, chained_data_delayed_19__82_, chained_data_delayed_19__81_, chained_data_delayed_19__80_, chained_data_delayed_19__79_, chained_data_delayed_19__78_, chained_data_delayed_19__77_, chained_data_delayed_19__76_, chained_data_delayed_19__75_, chained_data_delayed_19__74_, chained_data_delayed_19__73_, chained_data_delayed_19__72_, chained_data_delayed_19__71_, chained_data_delayed_19__70_, chained_data_delayed_19__69_, chained_data_delayed_19__68_, chained_data_delayed_19__67_, chained_data_delayed_19__66_, chained_data_delayed_19__65_, chained_data_delayed_19__64_, chained_data_delayed_19__63_, chained_data_delayed_19__62_, chained_data_delayed_19__61_, chained_data_delayed_19__60_, chained_data_delayed_19__59_, chained_data_delayed_19__58_, chained_data_delayed_19__57_, chained_data_delayed_19__56_, chained_data_delayed_19__55_, chained_data_delayed_19__54_, chained_data_delayed_19__53_, chained_data_delayed_19__52_, chained_data_delayed_19__51_, chained_data_delayed_19__50_, chained_data_delayed_19__49_, chained_data_delayed_19__48_, chained_data_delayed_19__47_, chained_data_delayed_19__46_, chained_data_delayed_19__45_, chained_data_delayed_19__44_, chained_data_delayed_19__43_, chained_data_delayed_19__42_, chained_data_delayed_19__41_, chained_data_delayed_19__40_, chained_data_delayed_19__39_, chained_data_delayed_19__38_, chained_data_delayed_19__37_, chained_data_delayed_19__36_, chained_data_delayed_19__35_, chained_data_delayed_19__34_, chained_data_delayed_19__33_, chained_data_delayed_19__32_, chained_data_delayed_19__31_, chained_data_delayed_19__30_, chained_data_delayed_19__29_, chained_data_delayed_19__28_, chained_data_delayed_19__27_, chained_data_delayed_19__26_, chained_data_delayed_19__25_, chained_data_delayed_19__24_, chained_data_delayed_19__23_, chained_data_delayed_19__22_, chained_data_delayed_19__21_, chained_data_delayed_19__20_, chained_data_delayed_19__19_, chained_data_delayed_19__18_, chained_data_delayed_19__17_, chained_data_delayed_19__16_, chained_data_delayed_19__15_, chained_data_delayed_19__14_, chained_data_delayed_19__13_, chained_data_delayed_19__12_, chained_data_delayed_19__11_, chained_data_delayed_19__10_, chained_data_delayed_19__9_, chained_data_delayed_19__8_, chained_data_delayed_19__7_, chained_data_delayed_19__6_, chained_data_delayed_19__5_, chained_data_delayed_19__4_, chained_data_delayed_19__3_, chained_data_delayed_19__2_, chained_data_delayed_19__1_, chained_data_delayed_19__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_20__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_19__127_, chained_data_delayed_19__126_, chained_data_delayed_19__125_, chained_data_delayed_19__124_, chained_data_delayed_19__123_, chained_data_delayed_19__122_, chained_data_delayed_19__121_, chained_data_delayed_19__120_, chained_data_delayed_19__119_, chained_data_delayed_19__118_, chained_data_delayed_19__117_, chained_data_delayed_19__116_, chained_data_delayed_19__115_, chained_data_delayed_19__114_, chained_data_delayed_19__113_, chained_data_delayed_19__112_, chained_data_delayed_19__111_, chained_data_delayed_19__110_, chained_data_delayed_19__109_, chained_data_delayed_19__108_, chained_data_delayed_19__107_, chained_data_delayed_19__106_, chained_data_delayed_19__105_, chained_data_delayed_19__104_, chained_data_delayed_19__103_, chained_data_delayed_19__102_, chained_data_delayed_19__101_, chained_data_delayed_19__100_, chained_data_delayed_19__99_, chained_data_delayed_19__98_, chained_data_delayed_19__97_, chained_data_delayed_19__96_, chained_data_delayed_19__95_, chained_data_delayed_19__94_, chained_data_delayed_19__93_, chained_data_delayed_19__92_, chained_data_delayed_19__91_, chained_data_delayed_19__90_, chained_data_delayed_19__89_, chained_data_delayed_19__88_, chained_data_delayed_19__87_, chained_data_delayed_19__86_, chained_data_delayed_19__85_, chained_data_delayed_19__84_, chained_data_delayed_19__83_, chained_data_delayed_19__82_, chained_data_delayed_19__81_, chained_data_delayed_19__80_, chained_data_delayed_19__79_, chained_data_delayed_19__78_, chained_data_delayed_19__77_, chained_data_delayed_19__76_, chained_data_delayed_19__75_, chained_data_delayed_19__74_, chained_data_delayed_19__73_, chained_data_delayed_19__72_, chained_data_delayed_19__71_, chained_data_delayed_19__70_, chained_data_delayed_19__69_, chained_data_delayed_19__68_, chained_data_delayed_19__67_, chained_data_delayed_19__66_, chained_data_delayed_19__65_, chained_data_delayed_19__64_, chained_data_delayed_19__63_, chained_data_delayed_19__62_, chained_data_delayed_19__61_, chained_data_delayed_19__60_, chained_data_delayed_19__59_, chained_data_delayed_19__58_, chained_data_delayed_19__57_, chained_data_delayed_19__56_, chained_data_delayed_19__55_, chained_data_delayed_19__54_, chained_data_delayed_19__53_, chained_data_delayed_19__52_, chained_data_delayed_19__51_, chained_data_delayed_19__50_, chained_data_delayed_19__49_, chained_data_delayed_19__48_, chained_data_delayed_19__47_, chained_data_delayed_19__46_, chained_data_delayed_19__45_, chained_data_delayed_19__44_, chained_data_delayed_19__43_, chained_data_delayed_19__42_, chained_data_delayed_19__41_, chained_data_delayed_19__40_, chained_data_delayed_19__39_, chained_data_delayed_19__38_, chained_data_delayed_19__37_, chained_data_delayed_19__36_, chained_data_delayed_19__35_, chained_data_delayed_19__34_, chained_data_delayed_19__33_, chained_data_delayed_19__32_, chained_data_delayed_19__31_, chained_data_delayed_19__30_, chained_data_delayed_19__29_, chained_data_delayed_19__28_, chained_data_delayed_19__27_, chained_data_delayed_19__26_, chained_data_delayed_19__25_, chained_data_delayed_19__24_, chained_data_delayed_19__23_, chained_data_delayed_19__22_, chained_data_delayed_19__21_, chained_data_delayed_19__20_, chained_data_delayed_19__19_, chained_data_delayed_19__18_, chained_data_delayed_19__17_, chained_data_delayed_19__16_, chained_data_delayed_19__15_, chained_data_delayed_19__14_, chained_data_delayed_19__13_, chained_data_delayed_19__12_, chained_data_delayed_19__11_, chained_data_delayed_19__10_, chained_data_delayed_19__9_, chained_data_delayed_19__8_, chained_data_delayed_19__7_, chained_data_delayed_19__6_, chained_data_delayed_19__5_, chained_data_delayed_19__4_, chained_data_delayed_19__3_, chained_data_delayed_19__2_, chained_data_delayed_19__1_, chained_data_delayed_19__0_ }),
    .data_o({ chained_data_delayed_20__127_, chained_data_delayed_20__126_, chained_data_delayed_20__125_, chained_data_delayed_20__124_, chained_data_delayed_20__123_, chained_data_delayed_20__122_, chained_data_delayed_20__121_, chained_data_delayed_20__120_, chained_data_delayed_20__119_, chained_data_delayed_20__118_, chained_data_delayed_20__117_, chained_data_delayed_20__116_, chained_data_delayed_20__115_, chained_data_delayed_20__114_, chained_data_delayed_20__113_, chained_data_delayed_20__112_, chained_data_delayed_20__111_, chained_data_delayed_20__110_, chained_data_delayed_20__109_, chained_data_delayed_20__108_, chained_data_delayed_20__107_, chained_data_delayed_20__106_, chained_data_delayed_20__105_, chained_data_delayed_20__104_, chained_data_delayed_20__103_, chained_data_delayed_20__102_, chained_data_delayed_20__101_, chained_data_delayed_20__100_, chained_data_delayed_20__99_, chained_data_delayed_20__98_, chained_data_delayed_20__97_, chained_data_delayed_20__96_, chained_data_delayed_20__95_, chained_data_delayed_20__94_, chained_data_delayed_20__93_, chained_data_delayed_20__92_, chained_data_delayed_20__91_, chained_data_delayed_20__90_, chained_data_delayed_20__89_, chained_data_delayed_20__88_, chained_data_delayed_20__87_, chained_data_delayed_20__86_, chained_data_delayed_20__85_, chained_data_delayed_20__84_, chained_data_delayed_20__83_, chained_data_delayed_20__82_, chained_data_delayed_20__81_, chained_data_delayed_20__80_, chained_data_delayed_20__79_, chained_data_delayed_20__78_, chained_data_delayed_20__77_, chained_data_delayed_20__76_, chained_data_delayed_20__75_, chained_data_delayed_20__74_, chained_data_delayed_20__73_, chained_data_delayed_20__72_, chained_data_delayed_20__71_, chained_data_delayed_20__70_, chained_data_delayed_20__69_, chained_data_delayed_20__68_, chained_data_delayed_20__67_, chained_data_delayed_20__66_, chained_data_delayed_20__65_, chained_data_delayed_20__64_, chained_data_delayed_20__63_, chained_data_delayed_20__62_, chained_data_delayed_20__61_, chained_data_delayed_20__60_, chained_data_delayed_20__59_, chained_data_delayed_20__58_, chained_data_delayed_20__57_, chained_data_delayed_20__56_, chained_data_delayed_20__55_, chained_data_delayed_20__54_, chained_data_delayed_20__53_, chained_data_delayed_20__52_, chained_data_delayed_20__51_, chained_data_delayed_20__50_, chained_data_delayed_20__49_, chained_data_delayed_20__48_, chained_data_delayed_20__47_, chained_data_delayed_20__46_, chained_data_delayed_20__45_, chained_data_delayed_20__44_, chained_data_delayed_20__43_, chained_data_delayed_20__42_, chained_data_delayed_20__41_, chained_data_delayed_20__40_, chained_data_delayed_20__39_, chained_data_delayed_20__38_, chained_data_delayed_20__37_, chained_data_delayed_20__36_, chained_data_delayed_20__35_, chained_data_delayed_20__34_, chained_data_delayed_20__33_, chained_data_delayed_20__32_, chained_data_delayed_20__31_, chained_data_delayed_20__30_, chained_data_delayed_20__29_, chained_data_delayed_20__28_, chained_data_delayed_20__27_, chained_data_delayed_20__26_, chained_data_delayed_20__25_, chained_data_delayed_20__24_, chained_data_delayed_20__23_, chained_data_delayed_20__22_, chained_data_delayed_20__21_, chained_data_delayed_20__20_, chained_data_delayed_20__19_, chained_data_delayed_20__18_, chained_data_delayed_20__17_, chained_data_delayed_20__16_, chained_data_delayed_20__15_, chained_data_delayed_20__14_, chained_data_delayed_20__13_, chained_data_delayed_20__12_, chained_data_delayed_20__11_, chained_data_delayed_20__10_, chained_data_delayed_20__9_, chained_data_delayed_20__8_, chained_data_delayed_20__7_, chained_data_delayed_20__6_, chained_data_delayed_20__5_, chained_data_delayed_20__4_, chained_data_delayed_20__3_, chained_data_delayed_20__2_, chained_data_delayed_20__1_, chained_data_delayed_20__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_21__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_20__127_, chained_data_delayed_20__126_, chained_data_delayed_20__125_, chained_data_delayed_20__124_, chained_data_delayed_20__123_, chained_data_delayed_20__122_, chained_data_delayed_20__121_, chained_data_delayed_20__120_, chained_data_delayed_20__119_, chained_data_delayed_20__118_, chained_data_delayed_20__117_, chained_data_delayed_20__116_, chained_data_delayed_20__115_, chained_data_delayed_20__114_, chained_data_delayed_20__113_, chained_data_delayed_20__112_, chained_data_delayed_20__111_, chained_data_delayed_20__110_, chained_data_delayed_20__109_, chained_data_delayed_20__108_, chained_data_delayed_20__107_, chained_data_delayed_20__106_, chained_data_delayed_20__105_, chained_data_delayed_20__104_, chained_data_delayed_20__103_, chained_data_delayed_20__102_, chained_data_delayed_20__101_, chained_data_delayed_20__100_, chained_data_delayed_20__99_, chained_data_delayed_20__98_, chained_data_delayed_20__97_, chained_data_delayed_20__96_, chained_data_delayed_20__95_, chained_data_delayed_20__94_, chained_data_delayed_20__93_, chained_data_delayed_20__92_, chained_data_delayed_20__91_, chained_data_delayed_20__90_, chained_data_delayed_20__89_, chained_data_delayed_20__88_, chained_data_delayed_20__87_, chained_data_delayed_20__86_, chained_data_delayed_20__85_, chained_data_delayed_20__84_, chained_data_delayed_20__83_, chained_data_delayed_20__82_, chained_data_delayed_20__81_, chained_data_delayed_20__80_, chained_data_delayed_20__79_, chained_data_delayed_20__78_, chained_data_delayed_20__77_, chained_data_delayed_20__76_, chained_data_delayed_20__75_, chained_data_delayed_20__74_, chained_data_delayed_20__73_, chained_data_delayed_20__72_, chained_data_delayed_20__71_, chained_data_delayed_20__70_, chained_data_delayed_20__69_, chained_data_delayed_20__68_, chained_data_delayed_20__67_, chained_data_delayed_20__66_, chained_data_delayed_20__65_, chained_data_delayed_20__64_, chained_data_delayed_20__63_, chained_data_delayed_20__62_, chained_data_delayed_20__61_, chained_data_delayed_20__60_, chained_data_delayed_20__59_, chained_data_delayed_20__58_, chained_data_delayed_20__57_, chained_data_delayed_20__56_, chained_data_delayed_20__55_, chained_data_delayed_20__54_, chained_data_delayed_20__53_, chained_data_delayed_20__52_, chained_data_delayed_20__51_, chained_data_delayed_20__50_, chained_data_delayed_20__49_, chained_data_delayed_20__48_, chained_data_delayed_20__47_, chained_data_delayed_20__46_, chained_data_delayed_20__45_, chained_data_delayed_20__44_, chained_data_delayed_20__43_, chained_data_delayed_20__42_, chained_data_delayed_20__41_, chained_data_delayed_20__40_, chained_data_delayed_20__39_, chained_data_delayed_20__38_, chained_data_delayed_20__37_, chained_data_delayed_20__36_, chained_data_delayed_20__35_, chained_data_delayed_20__34_, chained_data_delayed_20__33_, chained_data_delayed_20__32_, chained_data_delayed_20__31_, chained_data_delayed_20__30_, chained_data_delayed_20__29_, chained_data_delayed_20__28_, chained_data_delayed_20__27_, chained_data_delayed_20__26_, chained_data_delayed_20__25_, chained_data_delayed_20__24_, chained_data_delayed_20__23_, chained_data_delayed_20__22_, chained_data_delayed_20__21_, chained_data_delayed_20__20_, chained_data_delayed_20__19_, chained_data_delayed_20__18_, chained_data_delayed_20__17_, chained_data_delayed_20__16_, chained_data_delayed_20__15_, chained_data_delayed_20__14_, chained_data_delayed_20__13_, chained_data_delayed_20__12_, chained_data_delayed_20__11_, chained_data_delayed_20__10_, chained_data_delayed_20__9_, chained_data_delayed_20__8_, chained_data_delayed_20__7_, chained_data_delayed_20__6_, chained_data_delayed_20__5_, chained_data_delayed_20__4_, chained_data_delayed_20__3_, chained_data_delayed_20__2_, chained_data_delayed_20__1_, chained_data_delayed_20__0_ }),
    .data_o({ chained_data_delayed_21__127_, chained_data_delayed_21__126_, chained_data_delayed_21__125_, chained_data_delayed_21__124_, chained_data_delayed_21__123_, chained_data_delayed_21__122_, chained_data_delayed_21__121_, chained_data_delayed_21__120_, chained_data_delayed_21__119_, chained_data_delayed_21__118_, chained_data_delayed_21__117_, chained_data_delayed_21__116_, chained_data_delayed_21__115_, chained_data_delayed_21__114_, chained_data_delayed_21__113_, chained_data_delayed_21__112_, chained_data_delayed_21__111_, chained_data_delayed_21__110_, chained_data_delayed_21__109_, chained_data_delayed_21__108_, chained_data_delayed_21__107_, chained_data_delayed_21__106_, chained_data_delayed_21__105_, chained_data_delayed_21__104_, chained_data_delayed_21__103_, chained_data_delayed_21__102_, chained_data_delayed_21__101_, chained_data_delayed_21__100_, chained_data_delayed_21__99_, chained_data_delayed_21__98_, chained_data_delayed_21__97_, chained_data_delayed_21__96_, chained_data_delayed_21__95_, chained_data_delayed_21__94_, chained_data_delayed_21__93_, chained_data_delayed_21__92_, chained_data_delayed_21__91_, chained_data_delayed_21__90_, chained_data_delayed_21__89_, chained_data_delayed_21__88_, chained_data_delayed_21__87_, chained_data_delayed_21__86_, chained_data_delayed_21__85_, chained_data_delayed_21__84_, chained_data_delayed_21__83_, chained_data_delayed_21__82_, chained_data_delayed_21__81_, chained_data_delayed_21__80_, chained_data_delayed_21__79_, chained_data_delayed_21__78_, chained_data_delayed_21__77_, chained_data_delayed_21__76_, chained_data_delayed_21__75_, chained_data_delayed_21__74_, chained_data_delayed_21__73_, chained_data_delayed_21__72_, chained_data_delayed_21__71_, chained_data_delayed_21__70_, chained_data_delayed_21__69_, chained_data_delayed_21__68_, chained_data_delayed_21__67_, chained_data_delayed_21__66_, chained_data_delayed_21__65_, chained_data_delayed_21__64_, chained_data_delayed_21__63_, chained_data_delayed_21__62_, chained_data_delayed_21__61_, chained_data_delayed_21__60_, chained_data_delayed_21__59_, chained_data_delayed_21__58_, chained_data_delayed_21__57_, chained_data_delayed_21__56_, chained_data_delayed_21__55_, chained_data_delayed_21__54_, chained_data_delayed_21__53_, chained_data_delayed_21__52_, chained_data_delayed_21__51_, chained_data_delayed_21__50_, chained_data_delayed_21__49_, chained_data_delayed_21__48_, chained_data_delayed_21__47_, chained_data_delayed_21__46_, chained_data_delayed_21__45_, chained_data_delayed_21__44_, chained_data_delayed_21__43_, chained_data_delayed_21__42_, chained_data_delayed_21__41_, chained_data_delayed_21__40_, chained_data_delayed_21__39_, chained_data_delayed_21__38_, chained_data_delayed_21__37_, chained_data_delayed_21__36_, chained_data_delayed_21__35_, chained_data_delayed_21__34_, chained_data_delayed_21__33_, chained_data_delayed_21__32_, chained_data_delayed_21__31_, chained_data_delayed_21__30_, chained_data_delayed_21__29_, chained_data_delayed_21__28_, chained_data_delayed_21__27_, chained_data_delayed_21__26_, chained_data_delayed_21__25_, chained_data_delayed_21__24_, chained_data_delayed_21__23_, chained_data_delayed_21__22_, chained_data_delayed_21__21_, chained_data_delayed_21__20_, chained_data_delayed_21__19_, chained_data_delayed_21__18_, chained_data_delayed_21__17_, chained_data_delayed_21__16_, chained_data_delayed_21__15_, chained_data_delayed_21__14_, chained_data_delayed_21__13_, chained_data_delayed_21__12_, chained_data_delayed_21__11_, chained_data_delayed_21__10_, chained_data_delayed_21__9_, chained_data_delayed_21__8_, chained_data_delayed_21__7_, chained_data_delayed_21__6_, chained_data_delayed_21__5_, chained_data_delayed_21__4_, chained_data_delayed_21__3_, chained_data_delayed_21__2_, chained_data_delayed_21__1_, chained_data_delayed_21__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_22__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_21__127_, chained_data_delayed_21__126_, chained_data_delayed_21__125_, chained_data_delayed_21__124_, chained_data_delayed_21__123_, chained_data_delayed_21__122_, chained_data_delayed_21__121_, chained_data_delayed_21__120_, chained_data_delayed_21__119_, chained_data_delayed_21__118_, chained_data_delayed_21__117_, chained_data_delayed_21__116_, chained_data_delayed_21__115_, chained_data_delayed_21__114_, chained_data_delayed_21__113_, chained_data_delayed_21__112_, chained_data_delayed_21__111_, chained_data_delayed_21__110_, chained_data_delayed_21__109_, chained_data_delayed_21__108_, chained_data_delayed_21__107_, chained_data_delayed_21__106_, chained_data_delayed_21__105_, chained_data_delayed_21__104_, chained_data_delayed_21__103_, chained_data_delayed_21__102_, chained_data_delayed_21__101_, chained_data_delayed_21__100_, chained_data_delayed_21__99_, chained_data_delayed_21__98_, chained_data_delayed_21__97_, chained_data_delayed_21__96_, chained_data_delayed_21__95_, chained_data_delayed_21__94_, chained_data_delayed_21__93_, chained_data_delayed_21__92_, chained_data_delayed_21__91_, chained_data_delayed_21__90_, chained_data_delayed_21__89_, chained_data_delayed_21__88_, chained_data_delayed_21__87_, chained_data_delayed_21__86_, chained_data_delayed_21__85_, chained_data_delayed_21__84_, chained_data_delayed_21__83_, chained_data_delayed_21__82_, chained_data_delayed_21__81_, chained_data_delayed_21__80_, chained_data_delayed_21__79_, chained_data_delayed_21__78_, chained_data_delayed_21__77_, chained_data_delayed_21__76_, chained_data_delayed_21__75_, chained_data_delayed_21__74_, chained_data_delayed_21__73_, chained_data_delayed_21__72_, chained_data_delayed_21__71_, chained_data_delayed_21__70_, chained_data_delayed_21__69_, chained_data_delayed_21__68_, chained_data_delayed_21__67_, chained_data_delayed_21__66_, chained_data_delayed_21__65_, chained_data_delayed_21__64_, chained_data_delayed_21__63_, chained_data_delayed_21__62_, chained_data_delayed_21__61_, chained_data_delayed_21__60_, chained_data_delayed_21__59_, chained_data_delayed_21__58_, chained_data_delayed_21__57_, chained_data_delayed_21__56_, chained_data_delayed_21__55_, chained_data_delayed_21__54_, chained_data_delayed_21__53_, chained_data_delayed_21__52_, chained_data_delayed_21__51_, chained_data_delayed_21__50_, chained_data_delayed_21__49_, chained_data_delayed_21__48_, chained_data_delayed_21__47_, chained_data_delayed_21__46_, chained_data_delayed_21__45_, chained_data_delayed_21__44_, chained_data_delayed_21__43_, chained_data_delayed_21__42_, chained_data_delayed_21__41_, chained_data_delayed_21__40_, chained_data_delayed_21__39_, chained_data_delayed_21__38_, chained_data_delayed_21__37_, chained_data_delayed_21__36_, chained_data_delayed_21__35_, chained_data_delayed_21__34_, chained_data_delayed_21__33_, chained_data_delayed_21__32_, chained_data_delayed_21__31_, chained_data_delayed_21__30_, chained_data_delayed_21__29_, chained_data_delayed_21__28_, chained_data_delayed_21__27_, chained_data_delayed_21__26_, chained_data_delayed_21__25_, chained_data_delayed_21__24_, chained_data_delayed_21__23_, chained_data_delayed_21__22_, chained_data_delayed_21__21_, chained_data_delayed_21__20_, chained_data_delayed_21__19_, chained_data_delayed_21__18_, chained_data_delayed_21__17_, chained_data_delayed_21__16_, chained_data_delayed_21__15_, chained_data_delayed_21__14_, chained_data_delayed_21__13_, chained_data_delayed_21__12_, chained_data_delayed_21__11_, chained_data_delayed_21__10_, chained_data_delayed_21__9_, chained_data_delayed_21__8_, chained_data_delayed_21__7_, chained_data_delayed_21__6_, chained_data_delayed_21__5_, chained_data_delayed_21__4_, chained_data_delayed_21__3_, chained_data_delayed_21__2_, chained_data_delayed_21__1_, chained_data_delayed_21__0_ }),
    .data_o({ chained_data_delayed_22__127_, chained_data_delayed_22__126_, chained_data_delayed_22__125_, chained_data_delayed_22__124_, chained_data_delayed_22__123_, chained_data_delayed_22__122_, chained_data_delayed_22__121_, chained_data_delayed_22__120_, chained_data_delayed_22__119_, chained_data_delayed_22__118_, chained_data_delayed_22__117_, chained_data_delayed_22__116_, chained_data_delayed_22__115_, chained_data_delayed_22__114_, chained_data_delayed_22__113_, chained_data_delayed_22__112_, chained_data_delayed_22__111_, chained_data_delayed_22__110_, chained_data_delayed_22__109_, chained_data_delayed_22__108_, chained_data_delayed_22__107_, chained_data_delayed_22__106_, chained_data_delayed_22__105_, chained_data_delayed_22__104_, chained_data_delayed_22__103_, chained_data_delayed_22__102_, chained_data_delayed_22__101_, chained_data_delayed_22__100_, chained_data_delayed_22__99_, chained_data_delayed_22__98_, chained_data_delayed_22__97_, chained_data_delayed_22__96_, chained_data_delayed_22__95_, chained_data_delayed_22__94_, chained_data_delayed_22__93_, chained_data_delayed_22__92_, chained_data_delayed_22__91_, chained_data_delayed_22__90_, chained_data_delayed_22__89_, chained_data_delayed_22__88_, chained_data_delayed_22__87_, chained_data_delayed_22__86_, chained_data_delayed_22__85_, chained_data_delayed_22__84_, chained_data_delayed_22__83_, chained_data_delayed_22__82_, chained_data_delayed_22__81_, chained_data_delayed_22__80_, chained_data_delayed_22__79_, chained_data_delayed_22__78_, chained_data_delayed_22__77_, chained_data_delayed_22__76_, chained_data_delayed_22__75_, chained_data_delayed_22__74_, chained_data_delayed_22__73_, chained_data_delayed_22__72_, chained_data_delayed_22__71_, chained_data_delayed_22__70_, chained_data_delayed_22__69_, chained_data_delayed_22__68_, chained_data_delayed_22__67_, chained_data_delayed_22__66_, chained_data_delayed_22__65_, chained_data_delayed_22__64_, chained_data_delayed_22__63_, chained_data_delayed_22__62_, chained_data_delayed_22__61_, chained_data_delayed_22__60_, chained_data_delayed_22__59_, chained_data_delayed_22__58_, chained_data_delayed_22__57_, chained_data_delayed_22__56_, chained_data_delayed_22__55_, chained_data_delayed_22__54_, chained_data_delayed_22__53_, chained_data_delayed_22__52_, chained_data_delayed_22__51_, chained_data_delayed_22__50_, chained_data_delayed_22__49_, chained_data_delayed_22__48_, chained_data_delayed_22__47_, chained_data_delayed_22__46_, chained_data_delayed_22__45_, chained_data_delayed_22__44_, chained_data_delayed_22__43_, chained_data_delayed_22__42_, chained_data_delayed_22__41_, chained_data_delayed_22__40_, chained_data_delayed_22__39_, chained_data_delayed_22__38_, chained_data_delayed_22__37_, chained_data_delayed_22__36_, chained_data_delayed_22__35_, chained_data_delayed_22__34_, chained_data_delayed_22__33_, chained_data_delayed_22__32_, chained_data_delayed_22__31_, chained_data_delayed_22__30_, chained_data_delayed_22__29_, chained_data_delayed_22__28_, chained_data_delayed_22__27_, chained_data_delayed_22__26_, chained_data_delayed_22__25_, chained_data_delayed_22__24_, chained_data_delayed_22__23_, chained_data_delayed_22__22_, chained_data_delayed_22__21_, chained_data_delayed_22__20_, chained_data_delayed_22__19_, chained_data_delayed_22__18_, chained_data_delayed_22__17_, chained_data_delayed_22__16_, chained_data_delayed_22__15_, chained_data_delayed_22__14_, chained_data_delayed_22__13_, chained_data_delayed_22__12_, chained_data_delayed_22__11_, chained_data_delayed_22__10_, chained_data_delayed_22__9_, chained_data_delayed_22__8_, chained_data_delayed_22__7_, chained_data_delayed_22__6_, chained_data_delayed_22__5_, chained_data_delayed_22__4_, chained_data_delayed_22__3_, chained_data_delayed_22__2_, chained_data_delayed_22__1_, chained_data_delayed_22__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_23__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_22__127_, chained_data_delayed_22__126_, chained_data_delayed_22__125_, chained_data_delayed_22__124_, chained_data_delayed_22__123_, chained_data_delayed_22__122_, chained_data_delayed_22__121_, chained_data_delayed_22__120_, chained_data_delayed_22__119_, chained_data_delayed_22__118_, chained_data_delayed_22__117_, chained_data_delayed_22__116_, chained_data_delayed_22__115_, chained_data_delayed_22__114_, chained_data_delayed_22__113_, chained_data_delayed_22__112_, chained_data_delayed_22__111_, chained_data_delayed_22__110_, chained_data_delayed_22__109_, chained_data_delayed_22__108_, chained_data_delayed_22__107_, chained_data_delayed_22__106_, chained_data_delayed_22__105_, chained_data_delayed_22__104_, chained_data_delayed_22__103_, chained_data_delayed_22__102_, chained_data_delayed_22__101_, chained_data_delayed_22__100_, chained_data_delayed_22__99_, chained_data_delayed_22__98_, chained_data_delayed_22__97_, chained_data_delayed_22__96_, chained_data_delayed_22__95_, chained_data_delayed_22__94_, chained_data_delayed_22__93_, chained_data_delayed_22__92_, chained_data_delayed_22__91_, chained_data_delayed_22__90_, chained_data_delayed_22__89_, chained_data_delayed_22__88_, chained_data_delayed_22__87_, chained_data_delayed_22__86_, chained_data_delayed_22__85_, chained_data_delayed_22__84_, chained_data_delayed_22__83_, chained_data_delayed_22__82_, chained_data_delayed_22__81_, chained_data_delayed_22__80_, chained_data_delayed_22__79_, chained_data_delayed_22__78_, chained_data_delayed_22__77_, chained_data_delayed_22__76_, chained_data_delayed_22__75_, chained_data_delayed_22__74_, chained_data_delayed_22__73_, chained_data_delayed_22__72_, chained_data_delayed_22__71_, chained_data_delayed_22__70_, chained_data_delayed_22__69_, chained_data_delayed_22__68_, chained_data_delayed_22__67_, chained_data_delayed_22__66_, chained_data_delayed_22__65_, chained_data_delayed_22__64_, chained_data_delayed_22__63_, chained_data_delayed_22__62_, chained_data_delayed_22__61_, chained_data_delayed_22__60_, chained_data_delayed_22__59_, chained_data_delayed_22__58_, chained_data_delayed_22__57_, chained_data_delayed_22__56_, chained_data_delayed_22__55_, chained_data_delayed_22__54_, chained_data_delayed_22__53_, chained_data_delayed_22__52_, chained_data_delayed_22__51_, chained_data_delayed_22__50_, chained_data_delayed_22__49_, chained_data_delayed_22__48_, chained_data_delayed_22__47_, chained_data_delayed_22__46_, chained_data_delayed_22__45_, chained_data_delayed_22__44_, chained_data_delayed_22__43_, chained_data_delayed_22__42_, chained_data_delayed_22__41_, chained_data_delayed_22__40_, chained_data_delayed_22__39_, chained_data_delayed_22__38_, chained_data_delayed_22__37_, chained_data_delayed_22__36_, chained_data_delayed_22__35_, chained_data_delayed_22__34_, chained_data_delayed_22__33_, chained_data_delayed_22__32_, chained_data_delayed_22__31_, chained_data_delayed_22__30_, chained_data_delayed_22__29_, chained_data_delayed_22__28_, chained_data_delayed_22__27_, chained_data_delayed_22__26_, chained_data_delayed_22__25_, chained_data_delayed_22__24_, chained_data_delayed_22__23_, chained_data_delayed_22__22_, chained_data_delayed_22__21_, chained_data_delayed_22__20_, chained_data_delayed_22__19_, chained_data_delayed_22__18_, chained_data_delayed_22__17_, chained_data_delayed_22__16_, chained_data_delayed_22__15_, chained_data_delayed_22__14_, chained_data_delayed_22__13_, chained_data_delayed_22__12_, chained_data_delayed_22__11_, chained_data_delayed_22__10_, chained_data_delayed_22__9_, chained_data_delayed_22__8_, chained_data_delayed_22__7_, chained_data_delayed_22__6_, chained_data_delayed_22__5_, chained_data_delayed_22__4_, chained_data_delayed_22__3_, chained_data_delayed_22__2_, chained_data_delayed_22__1_, chained_data_delayed_22__0_ }),
    .data_o({ chained_data_delayed_23__127_, chained_data_delayed_23__126_, chained_data_delayed_23__125_, chained_data_delayed_23__124_, chained_data_delayed_23__123_, chained_data_delayed_23__122_, chained_data_delayed_23__121_, chained_data_delayed_23__120_, chained_data_delayed_23__119_, chained_data_delayed_23__118_, chained_data_delayed_23__117_, chained_data_delayed_23__116_, chained_data_delayed_23__115_, chained_data_delayed_23__114_, chained_data_delayed_23__113_, chained_data_delayed_23__112_, chained_data_delayed_23__111_, chained_data_delayed_23__110_, chained_data_delayed_23__109_, chained_data_delayed_23__108_, chained_data_delayed_23__107_, chained_data_delayed_23__106_, chained_data_delayed_23__105_, chained_data_delayed_23__104_, chained_data_delayed_23__103_, chained_data_delayed_23__102_, chained_data_delayed_23__101_, chained_data_delayed_23__100_, chained_data_delayed_23__99_, chained_data_delayed_23__98_, chained_data_delayed_23__97_, chained_data_delayed_23__96_, chained_data_delayed_23__95_, chained_data_delayed_23__94_, chained_data_delayed_23__93_, chained_data_delayed_23__92_, chained_data_delayed_23__91_, chained_data_delayed_23__90_, chained_data_delayed_23__89_, chained_data_delayed_23__88_, chained_data_delayed_23__87_, chained_data_delayed_23__86_, chained_data_delayed_23__85_, chained_data_delayed_23__84_, chained_data_delayed_23__83_, chained_data_delayed_23__82_, chained_data_delayed_23__81_, chained_data_delayed_23__80_, chained_data_delayed_23__79_, chained_data_delayed_23__78_, chained_data_delayed_23__77_, chained_data_delayed_23__76_, chained_data_delayed_23__75_, chained_data_delayed_23__74_, chained_data_delayed_23__73_, chained_data_delayed_23__72_, chained_data_delayed_23__71_, chained_data_delayed_23__70_, chained_data_delayed_23__69_, chained_data_delayed_23__68_, chained_data_delayed_23__67_, chained_data_delayed_23__66_, chained_data_delayed_23__65_, chained_data_delayed_23__64_, chained_data_delayed_23__63_, chained_data_delayed_23__62_, chained_data_delayed_23__61_, chained_data_delayed_23__60_, chained_data_delayed_23__59_, chained_data_delayed_23__58_, chained_data_delayed_23__57_, chained_data_delayed_23__56_, chained_data_delayed_23__55_, chained_data_delayed_23__54_, chained_data_delayed_23__53_, chained_data_delayed_23__52_, chained_data_delayed_23__51_, chained_data_delayed_23__50_, chained_data_delayed_23__49_, chained_data_delayed_23__48_, chained_data_delayed_23__47_, chained_data_delayed_23__46_, chained_data_delayed_23__45_, chained_data_delayed_23__44_, chained_data_delayed_23__43_, chained_data_delayed_23__42_, chained_data_delayed_23__41_, chained_data_delayed_23__40_, chained_data_delayed_23__39_, chained_data_delayed_23__38_, chained_data_delayed_23__37_, chained_data_delayed_23__36_, chained_data_delayed_23__35_, chained_data_delayed_23__34_, chained_data_delayed_23__33_, chained_data_delayed_23__32_, chained_data_delayed_23__31_, chained_data_delayed_23__30_, chained_data_delayed_23__29_, chained_data_delayed_23__28_, chained_data_delayed_23__27_, chained_data_delayed_23__26_, chained_data_delayed_23__25_, chained_data_delayed_23__24_, chained_data_delayed_23__23_, chained_data_delayed_23__22_, chained_data_delayed_23__21_, chained_data_delayed_23__20_, chained_data_delayed_23__19_, chained_data_delayed_23__18_, chained_data_delayed_23__17_, chained_data_delayed_23__16_, chained_data_delayed_23__15_, chained_data_delayed_23__14_, chained_data_delayed_23__13_, chained_data_delayed_23__12_, chained_data_delayed_23__11_, chained_data_delayed_23__10_, chained_data_delayed_23__9_, chained_data_delayed_23__8_, chained_data_delayed_23__7_, chained_data_delayed_23__6_, chained_data_delayed_23__5_, chained_data_delayed_23__4_, chained_data_delayed_23__3_, chained_data_delayed_23__2_, chained_data_delayed_23__1_, chained_data_delayed_23__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_24__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_23__127_, chained_data_delayed_23__126_, chained_data_delayed_23__125_, chained_data_delayed_23__124_, chained_data_delayed_23__123_, chained_data_delayed_23__122_, chained_data_delayed_23__121_, chained_data_delayed_23__120_, chained_data_delayed_23__119_, chained_data_delayed_23__118_, chained_data_delayed_23__117_, chained_data_delayed_23__116_, chained_data_delayed_23__115_, chained_data_delayed_23__114_, chained_data_delayed_23__113_, chained_data_delayed_23__112_, chained_data_delayed_23__111_, chained_data_delayed_23__110_, chained_data_delayed_23__109_, chained_data_delayed_23__108_, chained_data_delayed_23__107_, chained_data_delayed_23__106_, chained_data_delayed_23__105_, chained_data_delayed_23__104_, chained_data_delayed_23__103_, chained_data_delayed_23__102_, chained_data_delayed_23__101_, chained_data_delayed_23__100_, chained_data_delayed_23__99_, chained_data_delayed_23__98_, chained_data_delayed_23__97_, chained_data_delayed_23__96_, chained_data_delayed_23__95_, chained_data_delayed_23__94_, chained_data_delayed_23__93_, chained_data_delayed_23__92_, chained_data_delayed_23__91_, chained_data_delayed_23__90_, chained_data_delayed_23__89_, chained_data_delayed_23__88_, chained_data_delayed_23__87_, chained_data_delayed_23__86_, chained_data_delayed_23__85_, chained_data_delayed_23__84_, chained_data_delayed_23__83_, chained_data_delayed_23__82_, chained_data_delayed_23__81_, chained_data_delayed_23__80_, chained_data_delayed_23__79_, chained_data_delayed_23__78_, chained_data_delayed_23__77_, chained_data_delayed_23__76_, chained_data_delayed_23__75_, chained_data_delayed_23__74_, chained_data_delayed_23__73_, chained_data_delayed_23__72_, chained_data_delayed_23__71_, chained_data_delayed_23__70_, chained_data_delayed_23__69_, chained_data_delayed_23__68_, chained_data_delayed_23__67_, chained_data_delayed_23__66_, chained_data_delayed_23__65_, chained_data_delayed_23__64_, chained_data_delayed_23__63_, chained_data_delayed_23__62_, chained_data_delayed_23__61_, chained_data_delayed_23__60_, chained_data_delayed_23__59_, chained_data_delayed_23__58_, chained_data_delayed_23__57_, chained_data_delayed_23__56_, chained_data_delayed_23__55_, chained_data_delayed_23__54_, chained_data_delayed_23__53_, chained_data_delayed_23__52_, chained_data_delayed_23__51_, chained_data_delayed_23__50_, chained_data_delayed_23__49_, chained_data_delayed_23__48_, chained_data_delayed_23__47_, chained_data_delayed_23__46_, chained_data_delayed_23__45_, chained_data_delayed_23__44_, chained_data_delayed_23__43_, chained_data_delayed_23__42_, chained_data_delayed_23__41_, chained_data_delayed_23__40_, chained_data_delayed_23__39_, chained_data_delayed_23__38_, chained_data_delayed_23__37_, chained_data_delayed_23__36_, chained_data_delayed_23__35_, chained_data_delayed_23__34_, chained_data_delayed_23__33_, chained_data_delayed_23__32_, chained_data_delayed_23__31_, chained_data_delayed_23__30_, chained_data_delayed_23__29_, chained_data_delayed_23__28_, chained_data_delayed_23__27_, chained_data_delayed_23__26_, chained_data_delayed_23__25_, chained_data_delayed_23__24_, chained_data_delayed_23__23_, chained_data_delayed_23__22_, chained_data_delayed_23__21_, chained_data_delayed_23__20_, chained_data_delayed_23__19_, chained_data_delayed_23__18_, chained_data_delayed_23__17_, chained_data_delayed_23__16_, chained_data_delayed_23__15_, chained_data_delayed_23__14_, chained_data_delayed_23__13_, chained_data_delayed_23__12_, chained_data_delayed_23__11_, chained_data_delayed_23__10_, chained_data_delayed_23__9_, chained_data_delayed_23__8_, chained_data_delayed_23__7_, chained_data_delayed_23__6_, chained_data_delayed_23__5_, chained_data_delayed_23__4_, chained_data_delayed_23__3_, chained_data_delayed_23__2_, chained_data_delayed_23__1_, chained_data_delayed_23__0_ }),
    .data_o({ chained_data_delayed_24__127_, chained_data_delayed_24__126_, chained_data_delayed_24__125_, chained_data_delayed_24__124_, chained_data_delayed_24__123_, chained_data_delayed_24__122_, chained_data_delayed_24__121_, chained_data_delayed_24__120_, chained_data_delayed_24__119_, chained_data_delayed_24__118_, chained_data_delayed_24__117_, chained_data_delayed_24__116_, chained_data_delayed_24__115_, chained_data_delayed_24__114_, chained_data_delayed_24__113_, chained_data_delayed_24__112_, chained_data_delayed_24__111_, chained_data_delayed_24__110_, chained_data_delayed_24__109_, chained_data_delayed_24__108_, chained_data_delayed_24__107_, chained_data_delayed_24__106_, chained_data_delayed_24__105_, chained_data_delayed_24__104_, chained_data_delayed_24__103_, chained_data_delayed_24__102_, chained_data_delayed_24__101_, chained_data_delayed_24__100_, chained_data_delayed_24__99_, chained_data_delayed_24__98_, chained_data_delayed_24__97_, chained_data_delayed_24__96_, chained_data_delayed_24__95_, chained_data_delayed_24__94_, chained_data_delayed_24__93_, chained_data_delayed_24__92_, chained_data_delayed_24__91_, chained_data_delayed_24__90_, chained_data_delayed_24__89_, chained_data_delayed_24__88_, chained_data_delayed_24__87_, chained_data_delayed_24__86_, chained_data_delayed_24__85_, chained_data_delayed_24__84_, chained_data_delayed_24__83_, chained_data_delayed_24__82_, chained_data_delayed_24__81_, chained_data_delayed_24__80_, chained_data_delayed_24__79_, chained_data_delayed_24__78_, chained_data_delayed_24__77_, chained_data_delayed_24__76_, chained_data_delayed_24__75_, chained_data_delayed_24__74_, chained_data_delayed_24__73_, chained_data_delayed_24__72_, chained_data_delayed_24__71_, chained_data_delayed_24__70_, chained_data_delayed_24__69_, chained_data_delayed_24__68_, chained_data_delayed_24__67_, chained_data_delayed_24__66_, chained_data_delayed_24__65_, chained_data_delayed_24__64_, chained_data_delayed_24__63_, chained_data_delayed_24__62_, chained_data_delayed_24__61_, chained_data_delayed_24__60_, chained_data_delayed_24__59_, chained_data_delayed_24__58_, chained_data_delayed_24__57_, chained_data_delayed_24__56_, chained_data_delayed_24__55_, chained_data_delayed_24__54_, chained_data_delayed_24__53_, chained_data_delayed_24__52_, chained_data_delayed_24__51_, chained_data_delayed_24__50_, chained_data_delayed_24__49_, chained_data_delayed_24__48_, chained_data_delayed_24__47_, chained_data_delayed_24__46_, chained_data_delayed_24__45_, chained_data_delayed_24__44_, chained_data_delayed_24__43_, chained_data_delayed_24__42_, chained_data_delayed_24__41_, chained_data_delayed_24__40_, chained_data_delayed_24__39_, chained_data_delayed_24__38_, chained_data_delayed_24__37_, chained_data_delayed_24__36_, chained_data_delayed_24__35_, chained_data_delayed_24__34_, chained_data_delayed_24__33_, chained_data_delayed_24__32_, chained_data_delayed_24__31_, chained_data_delayed_24__30_, chained_data_delayed_24__29_, chained_data_delayed_24__28_, chained_data_delayed_24__27_, chained_data_delayed_24__26_, chained_data_delayed_24__25_, chained_data_delayed_24__24_, chained_data_delayed_24__23_, chained_data_delayed_24__22_, chained_data_delayed_24__21_, chained_data_delayed_24__20_, chained_data_delayed_24__19_, chained_data_delayed_24__18_, chained_data_delayed_24__17_, chained_data_delayed_24__16_, chained_data_delayed_24__15_, chained_data_delayed_24__14_, chained_data_delayed_24__13_, chained_data_delayed_24__12_, chained_data_delayed_24__11_, chained_data_delayed_24__10_, chained_data_delayed_24__9_, chained_data_delayed_24__8_, chained_data_delayed_24__7_, chained_data_delayed_24__6_, chained_data_delayed_24__5_, chained_data_delayed_24__4_, chained_data_delayed_24__3_, chained_data_delayed_24__2_, chained_data_delayed_24__1_, chained_data_delayed_24__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_25__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_24__127_, chained_data_delayed_24__126_, chained_data_delayed_24__125_, chained_data_delayed_24__124_, chained_data_delayed_24__123_, chained_data_delayed_24__122_, chained_data_delayed_24__121_, chained_data_delayed_24__120_, chained_data_delayed_24__119_, chained_data_delayed_24__118_, chained_data_delayed_24__117_, chained_data_delayed_24__116_, chained_data_delayed_24__115_, chained_data_delayed_24__114_, chained_data_delayed_24__113_, chained_data_delayed_24__112_, chained_data_delayed_24__111_, chained_data_delayed_24__110_, chained_data_delayed_24__109_, chained_data_delayed_24__108_, chained_data_delayed_24__107_, chained_data_delayed_24__106_, chained_data_delayed_24__105_, chained_data_delayed_24__104_, chained_data_delayed_24__103_, chained_data_delayed_24__102_, chained_data_delayed_24__101_, chained_data_delayed_24__100_, chained_data_delayed_24__99_, chained_data_delayed_24__98_, chained_data_delayed_24__97_, chained_data_delayed_24__96_, chained_data_delayed_24__95_, chained_data_delayed_24__94_, chained_data_delayed_24__93_, chained_data_delayed_24__92_, chained_data_delayed_24__91_, chained_data_delayed_24__90_, chained_data_delayed_24__89_, chained_data_delayed_24__88_, chained_data_delayed_24__87_, chained_data_delayed_24__86_, chained_data_delayed_24__85_, chained_data_delayed_24__84_, chained_data_delayed_24__83_, chained_data_delayed_24__82_, chained_data_delayed_24__81_, chained_data_delayed_24__80_, chained_data_delayed_24__79_, chained_data_delayed_24__78_, chained_data_delayed_24__77_, chained_data_delayed_24__76_, chained_data_delayed_24__75_, chained_data_delayed_24__74_, chained_data_delayed_24__73_, chained_data_delayed_24__72_, chained_data_delayed_24__71_, chained_data_delayed_24__70_, chained_data_delayed_24__69_, chained_data_delayed_24__68_, chained_data_delayed_24__67_, chained_data_delayed_24__66_, chained_data_delayed_24__65_, chained_data_delayed_24__64_, chained_data_delayed_24__63_, chained_data_delayed_24__62_, chained_data_delayed_24__61_, chained_data_delayed_24__60_, chained_data_delayed_24__59_, chained_data_delayed_24__58_, chained_data_delayed_24__57_, chained_data_delayed_24__56_, chained_data_delayed_24__55_, chained_data_delayed_24__54_, chained_data_delayed_24__53_, chained_data_delayed_24__52_, chained_data_delayed_24__51_, chained_data_delayed_24__50_, chained_data_delayed_24__49_, chained_data_delayed_24__48_, chained_data_delayed_24__47_, chained_data_delayed_24__46_, chained_data_delayed_24__45_, chained_data_delayed_24__44_, chained_data_delayed_24__43_, chained_data_delayed_24__42_, chained_data_delayed_24__41_, chained_data_delayed_24__40_, chained_data_delayed_24__39_, chained_data_delayed_24__38_, chained_data_delayed_24__37_, chained_data_delayed_24__36_, chained_data_delayed_24__35_, chained_data_delayed_24__34_, chained_data_delayed_24__33_, chained_data_delayed_24__32_, chained_data_delayed_24__31_, chained_data_delayed_24__30_, chained_data_delayed_24__29_, chained_data_delayed_24__28_, chained_data_delayed_24__27_, chained_data_delayed_24__26_, chained_data_delayed_24__25_, chained_data_delayed_24__24_, chained_data_delayed_24__23_, chained_data_delayed_24__22_, chained_data_delayed_24__21_, chained_data_delayed_24__20_, chained_data_delayed_24__19_, chained_data_delayed_24__18_, chained_data_delayed_24__17_, chained_data_delayed_24__16_, chained_data_delayed_24__15_, chained_data_delayed_24__14_, chained_data_delayed_24__13_, chained_data_delayed_24__12_, chained_data_delayed_24__11_, chained_data_delayed_24__10_, chained_data_delayed_24__9_, chained_data_delayed_24__8_, chained_data_delayed_24__7_, chained_data_delayed_24__6_, chained_data_delayed_24__5_, chained_data_delayed_24__4_, chained_data_delayed_24__3_, chained_data_delayed_24__2_, chained_data_delayed_24__1_, chained_data_delayed_24__0_ }),
    .data_o({ chained_data_delayed_25__127_, chained_data_delayed_25__126_, chained_data_delayed_25__125_, chained_data_delayed_25__124_, chained_data_delayed_25__123_, chained_data_delayed_25__122_, chained_data_delayed_25__121_, chained_data_delayed_25__120_, chained_data_delayed_25__119_, chained_data_delayed_25__118_, chained_data_delayed_25__117_, chained_data_delayed_25__116_, chained_data_delayed_25__115_, chained_data_delayed_25__114_, chained_data_delayed_25__113_, chained_data_delayed_25__112_, chained_data_delayed_25__111_, chained_data_delayed_25__110_, chained_data_delayed_25__109_, chained_data_delayed_25__108_, chained_data_delayed_25__107_, chained_data_delayed_25__106_, chained_data_delayed_25__105_, chained_data_delayed_25__104_, chained_data_delayed_25__103_, chained_data_delayed_25__102_, chained_data_delayed_25__101_, chained_data_delayed_25__100_, chained_data_delayed_25__99_, chained_data_delayed_25__98_, chained_data_delayed_25__97_, chained_data_delayed_25__96_, chained_data_delayed_25__95_, chained_data_delayed_25__94_, chained_data_delayed_25__93_, chained_data_delayed_25__92_, chained_data_delayed_25__91_, chained_data_delayed_25__90_, chained_data_delayed_25__89_, chained_data_delayed_25__88_, chained_data_delayed_25__87_, chained_data_delayed_25__86_, chained_data_delayed_25__85_, chained_data_delayed_25__84_, chained_data_delayed_25__83_, chained_data_delayed_25__82_, chained_data_delayed_25__81_, chained_data_delayed_25__80_, chained_data_delayed_25__79_, chained_data_delayed_25__78_, chained_data_delayed_25__77_, chained_data_delayed_25__76_, chained_data_delayed_25__75_, chained_data_delayed_25__74_, chained_data_delayed_25__73_, chained_data_delayed_25__72_, chained_data_delayed_25__71_, chained_data_delayed_25__70_, chained_data_delayed_25__69_, chained_data_delayed_25__68_, chained_data_delayed_25__67_, chained_data_delayed_25__66_, chained_data_delayed_25__65_, chained_data_delayed_25__64_, chained_data_delayed_25__63_, chained_data_delayed_25__62_, chained_data_delayed_25__61_, chained_data_delayed_25__60_, chained_data_delayed_25__59_, chained_data_delayed_25__58_, chained_data_delayed_25__57_, chained_data_delayed_25__56_, chained_data_delayed_25__55_, chained_data_delayed_25__54_, chained_data_delayed_25__53_, chained_data_delayed_25__52_, chained_data_delayed_25__51_, chained_data_delayed_25__50_, chained_data_delayed_25__49_, chained_data_delayed_25__48_, chained_data_delayed_25__47_, chained_data_delayed_25__46_, chained_data_delayed_25__45_, chained_data_delayed_25__44_, chained_data_delayed_25__43_, chained_data_delayed_25__42_, chained_data_delayed_25__41_, chained_data_delayed_25__40_, chained_data_delayed_25__39_, chained_data_delayed_25__38_, chained_data_delayed_25__37_, chained_data_delayed_25__36_, chained_data_delayed_25__35_, chained_data_delayed_25__34_, chained_data_delayed_25__33_, chained_data_delayed_25__32_, chained_data_delayed_25__31_, chained_data_delayed_25__30_, chained_data_delayed_25__29_, chained_data_delayed_25__28_, chained_data_delayed_25__27_, chained_data_delayed_25__26_, chained_data_delayed_25__25_, chained_data_delayed_25__24_, chained_data_delayed_25__23_, chained_data_delayed_25__22_, chained_data_delayed_25__21_, chained_data_delayed_25__20_, chained_data_delayed_25__19_, chained_data_delayed_25__18_, chained_data_delayed_25__17_, chained_data_delayed_25__16_, chained_data_delayed_25__15_, chained_data_delayed_25__14_, chained_data_delayed_25__13_, chained_data_delayed_25__12_, chained_data_delayed_25__11_, chained_data_delayed_25__10_, chained_data_delayed_25__9_, chained_data_delayed_25__8_, chained_data_delayed_25__7_, chained_data_delayed_25__6_, chained_data_delayed_25__5_, chained_data_delayed_25__4_, chained_data_delayed_25__3_, chained_data_delayed_25__2_, chained_data_delayed_25__1_, chained_data_delayed_25__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_26__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_25__127_, chained_data_delayed_25__126_, chained_data_delayed_25__125_, chained_data_delayed_25__124_, chained_data_delayed_25__123_, chained_data_delayed_25__122_, chained_data_delayed_25__121_, chained_data_delayed_25__120_, chained_data_delayed_25__119_, chained_data_delayed_25__118_, chained_data_delayed_25__117_, chained_data_delayed_25__116_, chained_data_delayed_25__115_, chained_data_delayed_25__114_, chained_data_delayed_25__113_, chained_data_delayed_25__112_, chained_data_delayed_25__111_, chained_data_delayed_25__110_, chained_data_delayed_25__109_, chained_data_delayed_25__108_, chained_data_delayed_25__107_, chained_data_delayed_25__106_, chained_data_delayed_25__105_, chained_data_delayed_25__104_, chained_data_delayed_25__103_, chained_data_delayed_25__102_, chained_data_delayed_25__101_, chained_data_delayed_25__100_, chained_data_delayed_25__99_, chained_data_delayed_25__98_, chained_data_delayed_25__97_, chained_data_delayed_25__96_, chained_data_delayed_25__95_, chained_data_delayed_25__94_, chained_data_delayed_25__93_, chained_data_delayed_25__92_, chained_data_delayed_25__91_, chained_data_delayed_25__90_, chained_data_delayed_25__89_, chained_data_delayed_25__88_, chained_data_delayed_25__87_, chained_data_delayed_25__86_, chained_data_delayed_25__85_, chained_data_delayed_25__84_, chained_data_delayed_25__83_, chained_data_delayed_25__82_, chained_data_delayed_25__81_, chained_data_delayed_25__80_, chained_data_delayed_25__79_, chained_data_delayed_25__78_, chained_data_delayed_25__77_, chained_data_delayed_25__76_, chained_data_delayed_25__75_, chained_data_delayed_25__74_, chained_data_delayed_25__73_, chained_data_delayed_25__72_, chained_data_delayed_25__71_, chained_data_delayed_25__70_, chained_data_delayed_25__69_, chained_data_delayed_25__68_, chained_data_delayed_25__67_, chained_data_delayed_25__66_, chained_data_delayed_25__65_, chained_data_delayed_25__64_, chained_data_delayed_25__63_, chained_data_delayed_25__62_, chained_data_delayed_25__61_, chained_data_delayed_25__60_, chained_data_delayed_25__59_, chained_data_delayed_25__58_, chained_data_delayed_25__57_, chained_data_delayed_25__56_, chained_data_delayed_25__55_, chained_data_delayed_25__54_, chained_data_delayed_25__53_, chained_data_delayed_25__52_, chained_data_delayed_25__51_, chained_data_delayed_25__50_, chained_data_delayed_25__49_, chained_data_delayed_25__48_, chained_data_delayed_25__47_, chained_data_delayed_25__46_, chained_data_delayed_25__45_, chained_data_delayed_25__44_, chained_data_delayed_25__43_, chained_data_delayed_25__42_, chained_data_delayed_25__41_, chained_data_delayed_25__40_, chained_data_delayed_25__39_, chained_data_delayed_25__38_, chained_data_delayed_25__37_, chained_data_delayed_25__36_, chained_data_delayed_25__35_, chained_data_delayed_25__34_, chained_data_delayed_25__33_, chained_data_delayed_25__32_, chained_data_delayed_25__31_, chained_data_delayed_25__30_, chained_data_delayed_25__29_, chained_data_delayed_25__28_, chained_data_delayed_25__27_, chained_data_delayed_25__26_, chained_data_delayed_25__25_, chained_data_delayed_25__24_, chained_data_delayed_25__23_, chained_data_delayed_25__22_, chained_data_delayed_25__21_, chained_data_delayed_25__20_, chained_data_delayed_25__19_, chained_data_delayed_25__18_, chained_data_delayed_25__17_, chained_data_delayed_25__16_, chained_data_delayed_25__15_, chained_data_delayed_25__14_, chained_data_delayed_25__13_, chained_data_delayed_25__12_, chained_data_delayed_25__11_, chained_data_delayed_25__10_, chained_data_delayed_25__9_, chained_data_delayed_25__8_, chained_data_delayed_25__7_, chained_data_delayed_25__6_, chained_data_delayed_25__5_, chained_data_delayed_25__4_, chained_data_delayed_25__3_, chained_data_delayed_25__2_, chained_data_delayed_25__1_, chained_data_delayed_25__0_ }),
    .data_o({ chained_data_delayed_26__127_, chained_data_delayed_26__126_, chained_data_delayed_26__125_, chained_data_delayed_26__124_, chained_data_delayed_26__123_, chained_data_delayed_26__122_, chained_data_delayed_26__121_, chained_data_delayed_26__120_, chained_data_delayed_26__119_, chained_data_delayed_26__118_, chained_data_delayed_26__117_, chained_data_delayed_26__116_, chained_data_delayed_26__115_, chained_data_delayed_26__114_, chained_data_delayed_26__113_, chained_data_delayed_26__112_, chained_data_delayed_26__111_, chained_data_delayed_26__110_, chained_data_delayed_26__109_, chained_data_delayed_26__108_, chained_data_delayed_26__107_, chained_data_delayed_26__106_, chained_data_delayed_26__105_, chained_data_delayed_26__104_, chained_data_delayed_26__103_, chained_data_delayed_26__102_, chained_data_delayed_26__101_, chained_data_delayed_26__100_, chained_data_delayed_26__99_, chained_data_delayed_26__98_, chained_data_delayed_26__97_, chained_data_delayed_26__96_, chained_data_delayed_26__95_, chained_data_delayed_26__94_, chained_data_delayed_26__93_, chained_data_delayed_26__92_, chained_data_delayed_26__91_, chained_data_delayed_26__90_, chained_data_delayed_26__89_, chained_data_delayed_26__88_, chained_data_delayed_26__87_, chained_data_delayed_26__86_, chained_data_delayed_26__85_, chained_data_delayed_26__84_, chained_data_delayed_26__83_, chained_data_delayed_26__82_, chained_data_delayed_26__81_, chained_data_delayed_26__80_, chained_data_delayed_26__79_, chained_data_delayed_26__78_, chained_data_delayed_26__77_, chained_data_delayed_26__76_, chained_data_delayed_26__75_, chained_data_delayed_26__74_, chained_data_delayed_26__73_, chained_data_delayed_26__72_, chained_data_delayed_26__71_, chained_data_delayed_26__70_, chained_data_delayed_26__69_, chained_data_delayed_26__68_, chained_data_delayed_26__67_, chained_data_delayed_26__66_, chained_data_delayed_26__65_, chained_data_delayed_26__64_, chained_data_delayed_26__63_, chained_data_delayed_26__62_, chained_data_delayed_26__61_, chained_data_delayed_26__60_, chained_data_delayed_26__59_, chained_data_delayed_26__58_, chained_data_delayed_26__57_, chained_data_delayed_26__56_, chained_data_delayed_26__55_, chained_data_delayed_26__54_, chained_data_delayed_26__53_, chained_data_delayed_26__52_, chained_data_delayed_26__51_, chained_data_delayed_26__50_, chained_data_delayed_26__49_, chained_data_delayed_26__48_, chained_data_delayed_26__47_, chained_data_delayed_26__46_, chained_data_delayed_26__45_, chained_data_delayed_26__44_, chained_data_delayed_26__43_, chained_data_delayed_26__42_, chained_data_delayed_26__41_, chained_data_delayed_26__40_, chained_data_delayed_26__39_, chained_data_delayed_26__38_, chained_data_delayed_26__37_, chained_data_delayed_26__36_, chained_data_delayed_26__35_, chained_data_delayed_26__34_, chained_data_delayed_26__33_, chained_data_delayed_26__32_, chained_data_delayed_26__31_, chained_data_delayed_26__30_, chained_data_delayed_26__29_, chained_data_delayed_26__28_, chained_data_delayed_26__27_, chained_data_delayed_26__26_, chained_data_delayed_26__25_, chained_data_delayed_26__24_, chained_data_delayed_26__23_, chained_data_delayed_26__22_, chained_data_delayed_26__21_, chained_data_delayed_26__20_, chained_data_delayed_26__19_, chained_data_delayed_26__18_, chained_data_delayed_26__17_, chained_data_delayed_26__16_, chained_data_delayed_26__15_, chained_data_delayed_26__14_, chained_data_delayed_26__13_, chained_data_delayed_26__12_, chained_data_delayed_26__11_, chained_data_delayed_26__10_, chained_data_delayed_26__9_, chained_data_delayed_26__8_, chained_data_delayed_26__7_, chained_data_delayed_26__6_, chained_data_delayed_26__5_, chained_data_delayed_26__4_, chained_data_delayed_26__3_, chained_data_delayed_26__2_, chained_data_delayed_26__1_, chained_data_delayed_26__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_27__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_26__127_, chained_data_delayed_26__126_, chained_data_delayed_26__125_, chained_data_delayed_26__124_, chained_data_delayed_26__123_, chained_data_delayed_26__122_, chained_data_delayed_26__121_, chained_data_delayed_26__120_, chained_data_delayed_26__119_, chained_data_delayed_26__118_, chained_data_delayed_26__117_, chained_data_delayed_26__116_, chained_data_delayed_26__115_, chained_data_delayed_26__114_, chained_data_delayed_26__113_, chained_data_delayed_26__112_, chained_data_delayed_26__111_, chained_data_delayed_26__110_, chained_data_delayed_26__109_, chained_data_delayed_26__108_, chained_data_delayed_26__107_, chained_data_delayed_26__106_, chained_data_delayed_26__105_, chained_data_delayed_26__104_, chained_data_delayed_26__103_, chained_data_delayed_26__102_, chained_data_delayed_26__101_, chained_data_delayed_26__100_, chained_data_delayed_26__99_, chained_data_delayed_26__98_, chained_data_delayed_26__97_, chained_data_delayed_26__96_, chained_data_delayed_26__95_, chained_data_delayed_26__94_, chained_data_delayed_26__93_, chained_data_delayed_26__92_, chained_data_delayed_26__91_, chained_data_delayed_26__90_, chained_data_delayed_26__89_, chained_data_delayed_26__88_, chained_data_delayed_26__87_, chained_data_delayed_26__86_, chained_data_delayed_26__85_, chained_data_delayed_26__84_, chained_data_delayed_26__83_, chained_data_delayed_26__82_, chained_data_delayed_26__81_, chained_data_delayed_26__80_, chained_data_delayed_26__79_, chained_data_delayed_26__78_, chained_data_delayed_26__77_, chained_data_delayed_26__76_, chained_data_delayed_26__75_, chained_data_delayed_26__74_, chained_data_delayed_26__73_, chained_data_delayed_26__72_, chained_data_delayed_26__71_, chained_data_delayed_26__70_, chained_data_delayed_26__69_, chained_data_delayed_26__68_, chained_data_delayed_26__67_, chained_data_delayed_26__66_, chained_data_delayed_26__65_, chained_data_delayed_26__64_, chained_data_delayed_26__63_, chained_data_delayed_26__62_, chained_data_delayed_26__61_, chained_data_delayed_26__60_, chained_data_delayed_26__59_, chained_data_delayed_26__58_, chained_data_delayed_26__57_, chained_data_delayed_26__56_, chained_data_delayed_26__55_, chained_data_delayed_26__54_, chained_data_delayed_26__53_, chained_data_delayed_26__52_, chained_data_delayed_26__51_, chained_data_delayed_26__50_, chained_data_delayed_26__49_, chained_data_delayed_26__48_, chained_data_delayed_26__47_, chained_data_delayed_26__46_, chained_data_delayed_26__45_, chained_data_delayed_26__44_, chained_data_delayed_26__43_, chained_data_delayed_26__42_, chained_data_delayed_26__41_, chained_data_delayed_26__40_, chained_data_delayed_26__39_, chained_data_delayed_26__38_, chained_data_delayed_26__37_, chained_data_delayed_26__36_, chained_data_delayed_26__35_, chained_data_delayed_26__34_, chained_data_delayed_26__33_, chained_data_delayed_26__32_, chained_data_delayed_26__31_, chained_data_delayed_26__30_, chained_data_delayed_26__29_, chained_data_delayed_26__28_, chained_data_delayed_26__27_, chained_data_delayed_26__26_, chained_data_delayed_26__25_, chained_data_delayed_26__24_, chained_data_delayed_26__23_, chained_data_delayed_26__22_, chained_data_delayed_26__21_, chained_data_delayed_26__20_, chained_data_delayed_26__19_, chained_data_delayed_26__18_, chained_data_delayed_26__17_, chained_data_delayed_26__16_, chained_data_delayed_26__15_, chained_data_delayed_26__14_, chained_data_delayed_26__13_, chained_data_delayed_26__12_, chained_data_delayed_26__11_, chained_data_delayed_26__10_, chained_data_delayed_26__9_, chained_data_delayed_26__8_, chained_data_delayed_26__7_, chained_data_delayed_26__6_, chained_data_delayed_26__5_, chained_data_delayed_26__4_, chained_data_delayed_26__3_, chained_data_delayed_26__2_, chained_data_delayed_26__1_, chained_data_delayed_26__0_ }),
    .data_o({ chained_data_delayed_27__127_, chained_data_delayed_27__126_, chained_data_delayed_27__125_, chained_data_delayed_27__124_, chained_data_delayed_27__123_, chained_data_delayed_27__122_, chained_data_delayed_27__121_, chained_data_delayed_27__120_, chained_data_delayed_27__119_, chained_data_delayed_27__118_, chained_data_delayed_27__117_, chained_data_delayed_27__116_, chained_data_delayed_27__115_, chained_data_delayed_27__114_, chained_data_delayed_27__113_, chained_data_delayed_27__112_, chained_data_delayed_27__111_, chained_data_delayed_27__110_, chained_data_delayed_27__109_, chained_data_delayed_27__108_, chained_data_delayed_27__107_, chained_data_delayed_27__106_, chained_data_delayed_27__105_, chained_data_delayed_27__104_, chained_data_delayed_27__103_, chained_data_delayed_27__102_, chained_data_delayed_27__101_, chained_data_delayed_27__100_, chained_data_delayed_27__99_, chained_data_delayed_27__98_, chained_data_delayed_27__97_, chained_data_delayed_27__96_, chained_data_delayed_27__95_, chained_data_delayed_27__94_, chained_data_delayed_27__93_, chained_data_delayed_27__92_, chained_data_delayed_27__91_, chained_data_delayed_27__90_, chained_data_delayed_27__89_, chained_data_delayed_27__88_, chained_data_delayed_27__87_, chained_data_delayed_27__86_, chained_data_delayed_27__85_, chained_data_delayed_27__84_, chained_data_delayed_27__83_, chained_data_delayed_27__82_, chained_data_delayed_27__81_, chained_data_delayed_27__80_, chained_data_delayed_27__79_, chained_data_delayed_27__78_, chained_data_delayed_27__77_, chained_data_delayed_27__76_, chained_data_delayed_27__75_, chained_data_delayed_27__74_, chained_data_delayed_27__73_, chained_data_delayed_27__72_, chained_data_delayed_27__71_, chained_data_delayed_27__70_, chained_data_delayed_27__69_, chained_data_delayed_27__68_, chained_data_delayed_27__67_, chained_data_delayed_27__66_, chained_data_delayed_27__65_, chained_data_delayed_27__64_, chained_data_delayed_27__63_, chained_data_delayed_27__62_, chained_data_delayed_27__61_, chained_data_delayed_27__60_, chained_data_delayed_27__59_, chained_data_delayed_27__58_, chained_data_delayed_27__57_, chained_data_delayed_27__56_, chained_data_delayed_27__55_, chained_data_delayed_27__54_, chained_data_delayed_27__53_, chained_data_delayed_27__52_, chained_data_delayed_27__51_, chained_data_delayed_27__50_, chained_data_delayed_27__49_, chained_data_delayed_27__48_, chained_data_delayed_27__47_, chained_data_delayed_27__46_, chained_data_delayed_27__45_, chained_data_delayed_27__44_, chained_data_delayed_27__43_, chained_data_delayed_27__42_, chained_data_delayed_27__41_, chained_data_delayed_27__40_, chained_data_delayed_27__39_, chained_data_delayed_27__38_, chained_data_delayed_27__37_, chained_data_delayed_27__36_, chained_data_delayed_27__35_, chained_data_delayed_27__34_, chained_data_delayed_27__33_, chained_data_delayed_27__32_, chained_data_delayed_27__31_, chained_data_delayed_27__30_, chained_data_delayed_27__29_, chained_data_delayed_27__28_, chained_data_delayed_27__27_, chained_data_delayed_27__26_, chained_data_delayed_27__25_, chained_data_delayed_27__24_, chained_data_delayed_27__23_, chained_data_delayed_27__22_, chained_data_delayed_27__21_, chained_data_delayed_27__20_, chained_data_delayed_27__19_, chained_data_delayed_27__18_, chained_data_delayed_27__17_, chained_data_delayed_27__16_, chained_data_delayed_27__15_, chained_data_delayed_27__14_, chained_data_delayed_27__13_, chained_data_delayed_27__12_, chained_data_delayed_27__11_, chained_data_delayed_27__10_, chained_data_delayed_27__9_, chained_data_delayed_27__8_, chained_data_delayed_27__7_, chained_data_delayed_27__6_, chained_data_delayed_27__5_, chained_data_delayed_27__4_, chained_data_delayed_27__3_, chained_data_delayed_27__2_, chained_data_delayed_27__1_, chained_data_delayed_27__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_28__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_27__127_, chained_data_delayed_27__126_, chained_data_delayed_27__125_, chained_data_delayed_27__124_, chained_data_delayed_27__123_, chained_data_delayed_27__122_, chained_data_delayed_27__121_, chained_data_delayed_27__120_, chained_data_delayed_27__119_, chained_data_delayed_27__118_, chained_data_delayed_27__117_, chained_data_delayed_27__116_, chained_data_delayed_27__115_, chained_data_delayed_27__114_, chained_data_delayed_27__113_, chained_data_delayed_27__112_, chained_data_delayed_27__111_, chained_data_delayed_27__110_, chained_data_delayed_27__109_, chained_data_delayed_27__108_, chained_data_delayed_27__107_, chained_data_delayed_27__106_, chained_data_delayed_27__105_, chained_data_delayed_27__104_, chained_data_delayed_27__103_, chained_data_delayed_27__102_, chained_data_delayed_27__101_, chained_data_delayed_27__100_, chained_data_delayed_27__99_, chained_data_delayed_27__98_, chained_data_delayed_27__97_, chained_data_delayed_27__96_, chained_data_delayed_27__95_, chained_data_delayed_27__94_, chained_data_delayed_27__93_, chained_data_delayed_27__92_, chained_data_delayed_27__91_, chained_data_delayed_27__90_, chained_data_delayed_27__89_, chained_data_delayed_27__88_, chained_data_delayed_27__87_, chained_data_delayed_27__86_, chained_data_delayed_27__85_, chained_data_delayed_27__84_, chained_data_delayed_27__83_, chained_data_delayed_27__82_, chained_data_delayed_27__81_, chained_data_delayed_27__80_, chained_data_delayed_27__79_, chained_data_delayed_27__78_, chained_data_delayed_27__77_, chained_data_delayed_27__76_, chained_data_delayed_27__75_, chained_data_delayed_27__74_, chained_data_delayed_27__73_, chained_data_delayed_27__72_, chained_data_delayed_27__71_, chained_data_delayed_27__70_, chained_data_delayed_27__69_, chained_data_delayed_27__68_, chained_data_delayed_27__67_, chained_data_delayed_27__66_, chained_data_delayed_27__65_, chained_data_delayed_27__64_, chained_data_delayed_27__63_, chained_data_delayed_27__62_, chained_data_delayed_27__61_, chained_data_delayed_27__60_, chained_data_delayed_27__59_, chained_data_delayed_27__58_, chained_data_delayed_27__57_, chained_data_delayed_27__56_, chained_data_delayed_27__55_, chained_data_delayed_27__54_, chained_data_delayed_27__53_, chained_data_delayed_27__52_, chained_data_delayed_27__51_, chained_data_delayed_27__50_, chained_data_delayed_27__49_, chained_data_delayed_27__48_, chained_data_delayed_27__47_, chained_data_delayed_27__46_, chained_data_delayed_27__45_, chained_data_delayed_27__44_, chained_data_delayed_27__43_, chained_data_delayed_27__42_, chained_data_delayed_27__41_, chained_data_delayed_27__40_, chained_data_delayed_27__39_, chained_data_delayed_27__38_, chained_data_delayed_27__37_, chained_data_delayed_27__36_, chained_data_delayed_27__35_, chained_data_delayed_27__34_, chained_data_delayed_27__33_, chained_data_delayed_27__32_, chained_data_delayed_27__31_, chained_data_delayed_27__30_, chained_data_delayed_27__29_, chained_data_delayed_27__28_, chained_data_delayed_27__27_, chained_data_delayed_27__26_, chained_data_delayed_27__25_, chained_data_delayed_27__24_, chained_data_delayed_27__23_, chained_data_delayed_27__22_, chained_data_delayed_27__21_, chained_data_delayed_27__20_, chained_data_delayed_27__19_, chained_data_delayed_27__18_, chained_data_delayed_27__17_, chained_data_delayed_27__16_, chained_data_delayed_27__15_, chained_data_delayed_27__14_, chained_data_delayed_27__13_, chained_data_delayed_27__12_, chained_data_delayed_27__11_, chained_data_delayed_27__10_, chained_data_delayed_27__9_, chained_data_delayed_27__8_, chained_data_delayed_27__7_, chained_data_delayed_27__6_, chained_data_delayed_27__5_, chained_data_delayed_27__4_, chained_data_delayed_27__3_, chained_data_delayed_27__2_, chained_data_delayed_27__1_, chained_data_delayed_27__0_ }),
    .data_o({ chained_data_delayed_28__127_, chained_data_delayed_28__126_, chained_data_delayed_28__125_, chained_data_delayed_28__124_, chained_data_delayed_28__123_, chained_data_delayed_28__122_, chained_data_delayed_28__121_, chained_data_delayed_28__120_, chained_data_delayed_28__119_, chained_data_delayed_28__118_, chained_data_delayed_28__117_, chained_data_delayed_28__116_, chained_data_delayed_28__115_, chained_data_delayed_28__114_, chained_data_delayed_28__113_, chained_data_delayed_28__112_, chained_data_delayed_28__111_, chained_data_delayed_28__110_, chained_data_delayed_28__109_, chained_data_delayed_28__108_, chained_data_delayed_28__107_, chained_data_delayed_28__106_, chained_data_delayed_28__105_, chained_data_delayed_28__104_, chained_data_delayed_28__103_, chained_data_delayed_28__102_, chained_data_delayed_28__101_, chained_data_delayed_28__100_, chained_data_delayed_28__99_, chained_data_delayed_28__98_, chained_data_delayed_28__97_, chained_data_delayed_28__96_, chained_data_delayed_28__95_, chained_data_delayed_28__94_, chained_data_delayed_28__93_, chained_data_delayed_28__92_, chained_data_delayed_28__91_, chained_data_delayed_28__90_, chained_data_delayed_28__89_, chained_data_delayed_28__88_, chained_data_delayed_28__87_, chained_data_delayed_28__86_, chained_data_delayed_28__85_, chained_data_delayed_28__84_, chained_data_delayed_28__83_, chained_data_delayed_28__82_, chained_data_delayed_28__81_, chained_data_delayed_28__80_, chained_data_delayed_28__79_, chained_data_delayed_28__78_, chained_data_delayed_28__77_, chained_data_delayed_28__76_, chained_data_delayed_28__75_, chained_data_delayed_28__74_, chained_data_delayed_28__73_, chained_data_delayed_28__72_, chained_data_delayed_28__71_, chained_data_delayed_28__70_, chained_data_delayed_28__69_, chained_data_delayed_28__68_, chained_data_delayed_28__67_, chained_data_delayed_28__66_, chained_data_delayed_28__65_, chained_data_delayed_28__64_, chained_data_delayed_28__63_, chained_data_delayed_28__62_, chained_data_delayed_28__61_, chained_data_delayed_28__60_, chained_data_delayed_28__59_, chained_data_delayed_28__58_, chained_data_delayed_28__57_, chained_data_delayed_28__56_, chained_data_delayed_28__55_, chained_data_delayed_28__54_, chained_data_delayed_28__53_, chained_data_delayed_28__52_, chained_data_delayed_28__51_, chained_data_delayed_28__50_, chained_data_delayed_28__49_, chained_data_delayed_28__48_, chained_data_delayed_28__47_, chained_data_delayed_28__46_, chained_data_delayed_28__45_, chained_data_delayed_28__44_, chained_data_delayed_28__43_, chained_data_delayed_28__42_, chained_data_delayed_28__41_, chained_data_delayed_28__40_, chained_data_delayed_28__39_, chained_data_delayed_28__38_, chained_data_delayed_28__37_, chained_data_delayed_28__36_, chained_data_delayed_28__35_, chained_data_delayed_28__34_, chained_data_delayed_28__33_, chained_data_delayed_28__32_, chained_data_delayed_28__31_, chained_data_delayed_28__30_, chained_data_delayed_28__29_, chained_data_delayed_28__28_, chained_data_delayed_28__27_, chained_data_delayed_28__26_, chained_data_delayed_28__25_, chained_data_delayed_28__24_, chained_data_delayed_28__23_, chained_data_delayed_28__22_, chained_data_delayed_28__21_, chained_data_delayed_28__20_, chained_data_delayed_28__19_, chained_data_delayed_28__18_, chained_data_delayed_28__17_, chained_data_delayed_28__16_, chained_data_delayed_28__15_, chained_data_delayed_28__14_, chained_data_delayed_28__13_, chained_data_delayed_28__12_, chained_data_delayed_28__11_, chained_data_delayed_28__10_, chained_data_delayed_28__9_, chained_data_delayed_28__8_, chained_data_delayed_28__7_, chained_data_delayed_28__6_, chained_data_delayed_28__5_, chained_data_delayed_28__4_, chained_data_delayed_28__3_, chained_data_delayed_28__2_, chained_data_delayed_28__1_, chained_data_delayed_28__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_29__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_28__127_, chained_data_delayed_28__126_, chained_data_delayed_28__125_, chained_data_delayed_28__124_, chained_data_delayed_28__123_, chained_data_delayed_28__122_, chained_data_delayed_28__121_, chained_data_delayed_28__120_, chained_data_delayed_28__119_, chained_data_delayed_28__118_, chained_data_delayed_28__117_, chained_data_delayed_28__116_, chained_data_delayed_28__115_, chained_data_delayed_28__114_, chained_data_delayed_28__113_, chained_data_delayed_28__112_, chained_data_delayed_28__111_, chained_data_delayed_28__110_, chained_data_delayed_28__109_, chained_data_delayed_28__108_, chained_data_delayed_28__107_, chained_data_delayed_28__106_, chained_data_delayed_28__105_, chained_data_delayed_28__104_, chained_data_delayed_28__103_, chained_data_delayed_28__102_, chained_data_delayed_28__101_, chained_data_delayed_28__100_, chained_data_delayed_28__99_, chained_data_delayed_28__98_, chained_data_delayed_28__97_, chained_data_delayed_28__96_, chained_data_delayed_28__95_, chained_data_delayed_28__94_, chained_data_delayed_28__93_, chained_data_delayed_28__92_, chained_data_delayed_28__91_, chained_data_delayed_28__90_, chained_data_delayed_28__89_, chained_data_delayed_28__88_, chained_data_delayed_28__87_, chained_data_delayed_28__86_, chained_data_delayed_28__85_, chained_data_delayed_28__84_, chained_data_delayed_28__83_, chained_data_delayed_28__82_, chained_data_delayed_28__81_, chained_data_delayed_28__80_, chained_data_delayed_28__79_, chained_data_delayed_28__78_, chained_data_delayed_28__77_, chained_data_delayed_28__76_, chained_data_delayed_28__75_, chained_data_delayed_28__74_, chained_data_delayed_28__73_, chained_data_delayed_28__72_, chained_data_delayed_28__71_, chained_data_delayed_28__70_, chained_data_delayed_28__69_, chained_data_delayed_28__68_, chained_data_delayed_28__67_, chained_data_delayed_28__66_, chained_data_delayed_28__65_, chained_data_delayed_28__64_, chained_data_delayed_28__63_, chained_data_delayed_28__62_, chained_data_delayed_28__61_, chained_data_delayed_28__60_, chained_data_delayed_28__59_, chained_data_delayed_28__58_, chained_data_delayed_28__57_, chained_data_delayed_28__56_, chained_data_delayed_28__55_, chained_data_delayed_28__54_, chained_data_delayed_28__53_, chained_data_delayed_28__52_, chained_data_delayed_28__51_, chained_data_delayed_28__50_, chained_data_delayed_28__49_, chained_data_delayed_28__48_, chained_data_delayed_28__47_, chained_data_delayed_28__46_, chained_data_delayed_28__45_, chained_data_delayed_28__44_, chained_data_delayed_28__43_, chained_data_delayed_28__42_, chained_data_delayed_28__41_, chained_data_delayed_28__40_, chained_data_delayed_28__39_, chained_data_delayed_28__38_, chained_data_delayed_28__37_, chained_data_delayed_28__36_, chained_data_delayed_28__35_, chained_data_delayed_28__34_, chained_data_delayed_28__33_, chained_data_delayed_28__32_, chained_data_delayed_28__31_, chained_data_delayed_28__30_, chained_data_delayed_28__29_, chained_data_delayed_28__28_, chained_data_delayed_28__27_, chained_data_delayed_28__26_, chained_data_delayed_28__25_, chained_data_delayed_28__24_, chained_data_delayed_28__23_, chained_data_delayed_28__22_, chained_data_delayed_28__21_, chained_data_delayed_28__20_, chained_data_delayed_28__19_, chained_data_delayed_28__18_, chained_data_delayed_28__17_, chained_data_delayed_28__16_, chained_data_delayed_28__15_, chained_data_delayed_28__14_, chained_data_delayed_28__13_, chained_data_delayed_28__12_, chained_data_delayed_28__11_, chained_data_delayed_28__10_, chained_data_delayed_28__9_, chained_data_delayed_28__8_, chained_data_delayed_28__7_, chained_data_delayed_28__6_, chained_data_delayed_28__5_, chained_data_delayed_28__4_, chained_data_delayed_28__3_, chained_data_delayed_28__2_, chained_data_delayed_28__1_, chained_data_delayed_28__0_ }),
    .data_o({ chained_data_delayed_29__127_, chained_data_delayed_29__126_, chained_data_delayed_29__125_, chained_data_delayed_29__124_, chained_data_delayed_29__123_, chained_data_delayed_29__122_, chained_data_delayed_29__121_, chained_data_delayed_29__120_, chained_data_delayed_29__119_, chained_data_delayed_29__118_, chained_data_delayed_29__117_, chained_data_delayed_29__116_, chained_data_delayed_29__115_, chained_data_delayed_29__114_, chained_data_delayed_29__113_, chained_data_delayed_29__112_, chained_data_delayed_29__111_, chained_data_delayed_29__110_, chained_data_delayed_29__109_, chained_data_delayed_29__108_, chained_data_delayed_29__107_, chained_data_delayed_29__106_, chained_data_delayed_29__105_, chained_data_delayed_29__104_, chained_data_delayed_29__103_, chained_data_delayed_29__102_, chained_data_delayed_29__101_, chained_data_delayed_29__100_, chained_data_delayed_29__99_, chained_data_delayed_29__98_, chained_data_delayed_29__97_, chained_data_delayed_29__96_, chained_data_delayed_29__95_, chained_data_delayed_29__94_, chained_data_delayed_29__93_, chained_data_delayed_29__92_, chained_data_delayed_29__91_, chained_data_delayed_29__90_, chained_data_delayed_29__89_, chained_data_delayed_29__88_, chained_data_delayed_29__87_, chained_data_delayed_29__86_, chained_data_delayed_29__85_, chained_data_delayed_29__84_, chained_data_delayed_29__83_, chained_data_delayed_29__82_, chained_data_delayed_29__81_, chained_data_delayed_29__80_, chained_data_delayed_29__79_, chained_data_delayed_29__78_, chained_data_delayed_29__77_, chained_data_delayed_29__76_, chained_data_delayed_29__75_, chained_data_delayed_29__74_, chained_data_delayed_29__73_, chained_data_delayed_29__72_, chained_data_delayed_29__71_, chained_data_delayed_29__70_, chained_data_delayed_29__69_, chained_data_delayed_29__68_, chained_data_delayed_29__67_, chained_data_delayed_29__66_, chained_data_delayed_29__65_, chained_data_delayed_29__64_, chained_data_delayed_29__63_, chained_data_delayed_29__62_, chained_data_delayed_29__61_, chained_data_delayed_29__60_, chained_data_delayed_29__59_, chained_data_delayed_29__58_, chained_data_delayed_29__57_, chained_data_delayed_29__56_, chained_data_delayed_29__55_, chained_data_delayed_29__54_, chained_data_delayed_29__53_, chained_data_delayed_29__52_, chained_data_delayed_29__51_, chained_data_delayed_29__50_, chained_data_delayed_29__49_, chained_data_delayed_29__48_, chained_data_delayed_29__47_, chained_data_delayed_29__46_, chained_data_delayed_29__45_, chained_data_delayed_29__44_, chained_data_delayed_29__43_, chained_data_delayed_29__42_, chained_data_delayed_29__41_, chained_data_delayed_29__40_, chained_data_delayed_29__39_, chained_data_delayed_29__38_, chained_data_delayed_29__37_, chained_data_delayed_29__36_, chained_data_delayed_29__35_, chained_data_delayed_29__34_, chained_data_delayed_29__33_, chained_data_delayed_29__32_, chained_data_delayed_29__31_, chained_data_delayed_29__30_, chained_data_delayed_29__29_, chained_data_delayed_29__28_, chained_data_delayed_29__27_, chained_data_delayed_29__26_, chained_data_delayed_29__25_, chained_data_delayed_29__24_, chained_data_delayed_29__23_, chained_data_delayed_29__22_, chained_data_delayed_29__21_, chained_data_delayed_29__20_, chained_data_delayed_29__19_, chained_data_delayed_29__18_, chained_data_delayed_29__17_, chained_data_delayed_29__16_, chained_data_delayed_29__15_, chained_data_delayed_29__14_, chained_data_delayed_29__13_, chained_data_delayed_29__12_, chained_data_delayed_29__11_, chained_data_delayed_29__10_, chained_data_delayed_29__9_, chained_data_delayed_29__8_, chained_data_delayed_29__7_, chained_data_delayed_29__6_, chained_data_delayed_29__5_, chained_data_delayed_29__4_, chained_data_delayed_29__3_, chained_data_delayed_29__2_, chained_data_delayed_29__1_, chained_data_delayed_29__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_30__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_29__127_, chained_data_delayed_29__126_, chained_data_delayed_29__125_, chained_data_delayed_29__124_, chained_data_delayed_29__123_, chained_data_delayed_29__122_, chained_data_delayed_29__121_, chained_data_delayed_29__120_, chained_data_delayed_29__119_, chained_data_delayed_29__118_, chained_data_delayed_29__117_, chained_data_delayed_29__116_, chained_data_delayed_29__115_, chained_data_delayed_29__114_, chained_data_delayed_29__113_, chained_data_delayed_29__112_, chained_data_delayed_29__111_, chained_data_delayed_29__110_, chained_data_delayed_29__109_, chained_data_delayed_29__108_, chained_data_delayed_29__107_, chained_data_delayed_29__106_, chained_data_delayed_29__105_, chained_data_delayed_29__104_, chained_data_delayed_29__103_, chained_data_delayed_29__102_, chained_data_delayed_29__101_, chained_data_delayed_29__100_, chained_data_delayed_29__99_, chained_data_delayed_29__98_, chained_data_delayed_29__97_, chained_data_delayed_29__96_, chained_data_delayed_29__95_, chained_data_delayed_29__94_, chained_data_delayed_29__93_, chained_data_delayed_29__92_, chained_data_delayed_29__91_, chained_data_delayed_29__90_, chained_data_delayed_29__89_, chained_data_delayed_29__88_, chained_data_delayed_29__87_, chained_data_delayed_29__86_, chained_data_delayed_29__85_, chained_data_delayed_29__84_, chained_data_delayed_29__83_, chained_data_delayed_29__82_, chained_data_delayed_29__81_, chained_data_delayed_29__80_, chained_data_delayed_29__79_, chained_data_delayed_29__78_, chained_data_delayed_29__77_, chained_data_delayed_29__76_, chained_data_delayed_29__75_, chained_data_delayed_29__74_, chained_data_delayed_29__73_, chained_data_delayed_29__72_, chained_data_delayed_29__71_, chained_data_delayed_29__70_, chained_data_delayed_29__69_, chained_data_delayed_29__68_, chained_data_delayed_29__67_, chained_data_delayed_29__66_, chained_data_delayed_29__65_, chained_data_delayed_29__64_, chained_data_delayed_29__63_, chained_data_delayed_29__62_, chained_data_delayed_29__61_, chained_data_delayed_29__60_, chained_data_delayed_29__59_, chained_data_delayed_29__58_, chained_data_delayed_29__57_, chained_data_delayed_29__56_, chained_data_delayed_29__55_, chained_data_delayed_29__54_, chained_data_delayed_29__53_, chained_data_delayed_29__52_, chained_data_delayed_29__51_, chained_data_delayed_29__50_, chained_data_delayed_29__49_, chained_data_delayed_29__48_, chained_data_delayed_29__47_, chained_data_delayed_29__46_, chained_data_delayed_29__45_, chained_data_delayed_29__44_, chained_data_delayed_29__43_, chained_data_delayed_29__42_, chained_data_delayed_29__41_, chained_data_delayed_29__40_, chained_data_delayed_29__39_, chained_data_delayed_29__38_, chained_data_delayed_29__37_, chained_data_delayed_29__36_, chained_data_delayed_29__35_, chained_data_delayed_29__34_, chained_data_delayed_29__33_, chained_data_delayed_29__32_, chained_data_delayed_29__31_, chained_data_delayed_29__30_, chained_data_delayed_29__29_, chained_data_delayed_29__28_, chained_data_delayed_29__27_, chained_data_delayed_29__26_, chained_data_delayed_29__25_, chained_data_delayed_29__24_, chained_data_delayed_29__23_, chained_data_delayed_29__22_, chained_data_delayed_29__21_, chained_data_delayed_29__20_, chained_data_delayed_29__19_, chained_data_delayed_29__18_, chained_data_delayed_29__17_, chained_data_delayed_29__16_, chained_data_delayed_29__15_, chained_data_delayed_29__14_, chained_data_delayed_29__13_, chained_data_delayed_29__12_, chained_data_delayed_29__11_, chained_data_delayed_29__10_, chained_data_delayed_29__9_, chained_data_delayed_29__8_, chained_data_delayed_29__7_, chained_data_delayed_29__6_, chained_data_delayed_29__5_, chained_data_delayed_29__4_, chained_data_delayed_29__3_, chained_data_delayed_29__2_, chained_data_delayed_29__1_, chained_data_delayed_29__0_ }),
    .data_o({ chained_data_delayed_30__127_, chained_data_delayed_30__126_, chained_data_delayed_30__125_, chained_data_delayed_30__124_, chained_data_delayed_30__123_, chained_data_delayed_30__122_, chained_data_delayed_30__121_, chained_data_delayed_30__120_, chained_data_delayed_30__119_, chained_data_delayed_30__118_, chained_data_delayed_30__117_, chained_data_delayed_30__116_, chained_data_delayed_30__115_, chained_data_delayed_30__114_, chained_data_delayed_30__113_, chained_data_delayed_30__112_, chained_data_delayed_30__111_, chained_data_delayed_30__110_, chained_data_delayed_30__109_, chained_data_delayed_30__108_, chained_data_delayed_30__107_, chained_data_delayed_30__106_, chained_data_delayed_30__105_, chained_data_delayed_30__104_, chained_data_delayed_30__103_, chained_data_delayed_30__102_, chained_data_delayed_30__101_, chained_data_delayed_30__100_, chained_data_delayed_30__99_, chained_data_delayed_30__98_, chained_data_delayed_30__97_, chained_data_delayed_30__96_, chained_data_delayed_30__95_, chained_data_delayed_30__94_, chained_data_delayed_30__93_, chained_data_delayed_30__92_, chained_data_delayed_30__91_, chained_data_delayed_30__90_, chained_data_delayed_30__89_, chained_data_delayed_30__88_, chained_data_delayed_30__87_, chained_data_delayed_30__86_, chained_data_delayed_30__85_, chained_data_delayed_30__84_, chained_data_delayed_30__83_, chained_data_delayed_30__82_, chained_data_delayed_30__81_, chained_data_delayed_30__80_, chained_data_delayed_30__79_, chained_data_delayed_30__78_, chained_data_delayed_30__77_, chained_data_delayed_30__76_, chained_data_delayed_30__75_, chained_data_delayed_30__74_, chained_data_delayed_30__73_, chained_data_delayed_30__72_, chained_data_delayed_30__71_, chained_data_delayed_30__70_, chained_data_delayed_30__69_, chained_data_delayed_30__68_, chained_data_delayed_30__67_, chained_data_delayed_30__66_, chained_data_delayed_30__65_, chained_data_delayed_30__64_, chained_data_delayed_30__63_, chained_data_delayed_30__62_, chained_data_delayed_30__61_, chained_data_delayed_30__60_, chained_data_delayed_30__59_, chained_data_delayed_30__58_, chained_data_delayed_30__57_, chained_data_delayed_30__56_, chained_data_delayed_30__55_, chained_data_delayed_30__54_, chained_data_delayed_30__53_, chained_data_delayed_30__52_, chained_data_delayed_30__51_, chained_data_delayed_30__50_, chained_data_delayed_30__49_, chained_data_delayed_30__48_, chained_data_delayed_30__47_, chained_data_delayed_30__46_, chained_data_delayed_30__45_, chained_data_delayed_30__44_, chained_data_delayed_30__43_, chained_data_delayed_30__42_, chained_data_delayed_30__41_, chained_data_delayed_30__40_, chained_data_delayed_30__39_, chained_data_delayed_30__38_, chained_data_delayed_30__37_, chained_data_delayed_30__36_, chained_data_delayed_30__35_, chained_data_delayed_30__34_, chained_data_delayed_30__33_, chained_data_delayed_30__32_, chained_data_delayed_30__31_, chained_data_delayed_30__30_, chained_data_delayed_30__29_, chained_data_delayed_30__28_, chained_data_delayed_30__27_, chained_data_delayed_30__26_, chained_data_delayed_30__25_, chained_data_delayed_30__24_, chained_data_delayed_30__23_, chained_data_delayed_30__22_, chained_data_delayed_30__21_, chained_data_delayed_30__20_, chained_data_delayed_30__19_, chained_data_delayed_30__18_, chained_data_delayed_30__17_, chained_data_delayed_30__16_, chained_data_delayed_30__15_, chained_data_delayed_30__14_, chained_data_delayed_30__13_, chained_data_delayed_30__12_, chained_data_delayed_30__11_, chained_data_delayed_30__10_, chained_data_delayed_30__9_, chained_data_delayed_30__8_, chained_data_delayed_30__7_, chained_data_delayed_30__6_, chained_data_delayed_30__5_, chained_data_delayed_30__4_, chained_data_delayed_30__3_, chained_data_delayed_30__2_, chained_data_delayed_30__1_, chained_data_delayed_30__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_31__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_30__127_, chained_data_delayed_30__126_, chained_data_delayed_30__125_, chained_data_delayed_30__124_, chained_data_delayed_30__123_, chained_data_delayed_30__122_, chained_data_delayed_30__121_, chained_data_delayed_30__120_, chained_data_delayed_30__119_, chained_data_delayed_30__118_, chained_data_delayed_30__117_, chained_data_delayed_30__116_, chained_data_delayed_30__115_, chained_data_delayed_30__114_, chained_data_delayed_30__113_, chained_data_delayed_30__112_, chained_data_delayed_30__111_, chained_data_delayed_30__110_, chained_data_delayed_30__109_, chained_data_delayed_30__108_, chained_data_delayed_30__107_, chained_data_delayed_30__106_, chained_data_delayed_30__105_, chained_data_delayed_30__104_, chained_data_delayed_30__103_, chained_data_delayed_30__102_, chained_data_delayed_30__101_, chained_data_delayed_30__100_, chained_data_delayed_30__99_, chained_data_delayed_30__98_, chained_data_delayed_30__97_, chained_data_delayed_30__96_, chained_data_delayed_30__95_, chained_data_delayed_30__94_, chained_data_delayed_30__93_, chained_data_delayed_30__92_, chained_data_delayed_30__91_, chained_data_delayed_30__90_, chained_data_delayed_30__89_, chained_data_delayed_30__88_, chained_data_delayed_30__87_, chained_data_delayed_30__86_, chained_data_delayed_30__85_, chained_data_delayed_30__84_, chained_data_delayed_30__83_, chained_data_delayed_30__82_, chained_data_delayed_30__81_, chained_data_delayed_30__80_, chained_data_delayed_30__79_, chained_data_delayed_30__78_, chained_data_delayed_30__77_, chained_data_delayed_30__76_, chained_data_delayed_30__75_, chained_data_delayed_30__74_, chained_data_delayed_30__73_, chained_data_delayed_30__72_, chained_data_delayed_30__71_, chained_data_delayed_30__70_, chained_data_delayed_30__69_, chained_data_delayed_30__68_, chained_data_delayed_30__67_, chained_data_delayed_30__66_, chained_data_delayed_30__65_, chained_data_delayed_30__64_, chained_data_delayed_30__63_, chained_data_delayed_30__62_, chained_data_delayed_30__61_, chained_data_delayed_30__60_, chained_data_delayed_30__59_, chained_data_delayed_30__58_, chained_data_delayed_30__57_, chained_data_delayed_30__56_, chained_data_delayed_30__55_, chained_data_delayed_30__54_, chained_data_delayed_30__53_, chained_data_delayed_30__52_, chained_data_delayed_30__51_, chained_data_delayed_30__50_, chained_data_delayed_30__49_, chained_data_delayed_30__48_, chained_data_delayed_30__47_, chained_data_delayed_30__46_, chained_data_delayed_30__45_, chained_data_delayed_30__44_, chained_data_delayed_30__43_, chained_data_delayed_30__42_, chained_data_delayed_30__41_, chained_data_delayed_30__40_, chained_data_delayed_30__39_, chained_data_delayed_30__38_, chained_data_delayed_30__37_, chained_data_delayed_30__36_, chained_data_delayed_30__35_, chained_data_delayed_30__34_, chained_data_delayed_30__33_, chained_data_delayed_30__32_, chained_data_delayed_30__31_, chained_data_delayed_30__30_, chained_data_delayed_30__29_, chained_data_delayed_30__28_, chained_data_delayed_30__27_, chained_data_delayed_30__26_, chained_data_delayed_30__25_, chained_data_delayed_30__24_, chained_data_delayed_30__23_, chained_data_delayed_30__22_, chained_data_delayed_30__21_, chained_data_delayed_30__20_, chained_data_delayed_30__19_, chained_data_delayed_30__18_, chained_data_delayed_30__17_, chained_data_delayed_30__16_, chained_data_delayed_30__15_, chained_data_delayed_30__14_, chained_data_delayed_30__13_, chained_data_delayed_30__12_, chained_data_delayed_30__11_, chained_data_delayed_30__10_, chained_data_delayed_30__9_, chained_data_delayed_30__8_, chained_data_delayed_30__7_, chained_data_delayed_30__6_, chained_data_delayed_30__5_, chained_data_delayed_30__4_, chained_data_delayed_30__3_, chained_data_delayed_30__2_, chained_data_delayed_30__1_, chained_data_delayed_30__0_ }),
    .data_o({ chained_data_delayed_31__127_, chained_data_delayed_31__126_, chained_data_delayed_31__125_, chained_data_delayed_31__124_, chained_data_delayed_31__123_, chained_data_delayed_31__122_, chained_data_delayed_31__121_, chained_data_delayed_31__120_, chained_data_delayed_31__119_, chained_data_delayed_31__118_, chained_data_delayed_31__117_, chained_data_delayed_31__116_, chained_data_delayed_31__115_, chained_data_delayed_31__114_, chained_data_delayed_31__113_, chained_data_delayed_31__112_, chained_data_delayed_31__111_, chained_data_delayed_31__110_, chained_data_delayed_31__109_, chained_data_delayed_31__108_, chained_data_delayed_31__107_, chained_data_delayed_31__106_, chained_data_delayed_31__105_, chained_data_delayed_31__104_, chained_data_delayed_31__103_, chained_data_delayed_31__102_, chained_data_delayed_31__101_, chained_data_delayed_31__100_, chained_data_delayed_31__99_, chained_data_delayed_31__98_, chained_data_delayed_31__97_, chained_data_delayed_31__96_, chained_data_delayed_31__95_, chained_data_delayed_31__94_, chained_data_delayed_31__93_, chained_data_delayed_31__92_, chained_data_delayed_31__91_, chained_data_delayed_31__90_, chained_data_delayed_31__89_, chained_data_delayed_31__88_, chained_data_delayed_31__87_, chained_data_delayed_31__86_, chained_data_delayed_31__85_, chained_data_delayed_31__84_, chained_data_delayed_31__83_, chained_data_delayed_31__82_, chained_data_delayed_31__81_, chained_data_delayed_31__80_, chained_data_delayed_31__79_, chained_data_delayed_31__78_, chained_data_delayed_31__77_, chained_data_delayed_31__76_, chained_data_delayed_31__75_, chained_data_delayed_31__74_, chained_data_delayed_31__73_, chained_data_delayed_31__72_, chained_data_delayed_31__71_, chained_data_delayed_31__70_, chained_data_delayed_31__69_, chained_data_delayed_31__68_, chained_data_delayed_31__67_, chained_data_delayed_31__66_, chained_data_delayed_31__65_, chained_data_delayed_31__64_, chained_data_delayed_31__63_, chained_data_delayed_31__62_, chained_data_delayed_31__61_, chained_data_delayed_31__60_, chained_data_delayed_31__59_, chained_data_delayed_31__58_, chained_data_delayed_31__57_, chained_data_delayed_31__56_, chained_data_delayed_31__55_, chained_data_delayed_31__54_, chained_data_delayed_31__53_, chained_data_delayed_31__52_, chained_data_delayed_31__51_, chained_data_delayed_31__50_, chained_data_delayed_31__49_, chained_data_delayed_31__48_, chained_data_delayed_31__47_, chained_data_delayed_31__46_, chained_data_delayed_31__45_, chained_data_delayed_31__44_, chained_data_delayed_31__43_, chained_data_delayed_31__42_, chained_data_delayed_31__41_, chained_data_delayed_31__40_, chained_data_delayed_31__39_, chained_data_delayed_31__38_, chained_data_delayed_31__37_, chained_data_delayed_31__36_, chained_data_delayed_31__35_, chained_data_delayed_31__34_, chained_data_delayed_31__33_, chained_data_delayed_31__32_, chained_data_delayed_31__31_, chained_data_delayed_31__30_, chained_data_delayed_31__29_, chained_data_delayed_31__28_, chained_data_delayed_31__27_, chained_data_delayed_31__26_, chained_data_delayed_31__25_, chained_data_delayed_31__24_, chained_data_delayed_31__23_, chained_data_delayed_31__22_, chained_data_delayed_31__21_, chained_data_delayed_31__20_, chained_data_delayed_31__19_, chained_data_delayed_31__18_, chained_data_delayed_31__17_, chained_data_delayed_31__16_, chained_data_delayed_31__15_, chained_data_delayed_31__14_, chained_data_delayed_31__13_, chained_data_delayed_31__12_, chained_data_delayed_31__11_, chained_data_delayed_31__10_, chained_data_delayed_31__9_, chained_data_delayed_31__8_, chained_data_delayed_31__7_, chained_data_delayed_31__6_, chained_data_delayed_31__5_, chained_data_delayed_31__4_, chained_data_delayed_31__3_, chained_data_delayed_31__2_, chained_data_delayed_31__1_, chained_data_delayed_31__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_32__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_31__127_, chained_data_delayed_31__126_, chained_data_delayed_31__125_, chained_data_delayed_31__124_, chained_data_delayed_31__123_, chained_data_delayed_31__122_, chained_data_delayed_31__121_, chained_data_delayed_31__120_, chained_data_delayed_31__119_, chained_data_delayed_31__118_, chained_data_delayed_31__117_, chained_data_delayed_31__116_, chained_data_delayed_31__115_, chained_data_delayed_31__114_, chained_data_delayed_31__113_, chained_data_delayed_31__112_, chained_data_delayed_31__111_, chained_data_delayed_31__110_, chained_data_delayed_31__109_, chained_data_delayed_31__108_, chained_data_delayed_31__107_, chained_data_delayed_31__106_, chained_data_delayed_31__105_, chained_data_delayed_31__104_, chained_data_delayed_31__103_, chained_data_delayed_31__102_, chained_data_delayed_31__101_, chained_data_delayed_31__100_, chained_data_delayed_31__99_, chained_data_delayed_31__98_, chained_data_delayed_31__97_, chained_data_delayed_31__96_, chained_data_delayed_31__95_, chained_data_delayed_31__94_, chained_data_delayed_31__93_, chained_data_delayed_31__92_, chained_data_delayed_31__91_, chained_data_delayed_31__90_, chained_data_delayed_31__89_, chained_data_delayed_31__88_, chained_data_delayed_31__87_, chained_data_delayed_31__86_, chained_data_delayed_31__85_, chained_data_delayed_31__84_, chained_data_delayed_31__83_, chained_data_delayed_31__82_, chained_data_delayed_31__81_, chained_data_delayed_31__80_, chained_data_delayed_31__79_, chained_data_delayed_31__78_, chained_data_delayed_31__77_, chained_data_delayed_31__76_, chained_data_delayed_31__75_, chained_data_delayed_31__74_, chained_data_delayed_31__73_, chained_data_delayed_31__72_, chained_data_delayed_31__71_, chained_data_delayed_31__70_, chained_data_delayed_31__69_, chained_data_delayed_31__68_, chained_data_delayed_31__67_, chained_data_delayed_31__66_, chained_data_delayed_31__65_, chained_data_delayed_31__64_, chained_data_delayed_31__63_, chained_data_delayed_31__62_, chained_data_delayed_31__61_, chained_data_delayed_31__60_, chained_data_delayed_31__59_, chained_data_delayed_31__58_, chained_data_delayed_31__57_, chained_data_delayed_31__56_, chained_data_delayed_31__55_, chained_data_delayed_31__54_, chained_data_delayed_31__53_, chained_data_delayed_31__52_, chained_data_delayed_31__51_, chained_data_delayed_31__50_, chained_data_delayed_31__49_, chained_data_delayed_31__48_, chained_data_delayed_31__47_, chained_data_delayed_31__46_, chained_data_delayed_31__45_, chained_data_delayed_31__44_, chained_data_delayed_31__43_, chained_data_delayed_31__42_, chained_data_delayed_31__41_, chained_data_delayed_31__40_, chained_data_delayed_31__39_, chained_data_delayed_31__38_, chained_data_delayed_31__37_, chained_data_delayed_31__36_, chained_data_delayed_31__35_, chained_data_delayed_31__34_, chained_data_delayed_31__33_, chained_data_delayed_31__32_, chained_data_delayed_31__31_, chained_data_delayed_31__30_, chained_data_delayed_31__29_, chained_data_delayed_31__28_, chained_data_delayed_31__27_, chained_data_delayed_31__26_, chained_data_delayed_31__25_, chained_data_delayed_31__24_, chained_data_delayed_31__23_, chained_data_delayed_31__22_, chained_data_delayed_31__21_, chained_data_delayed_31__20_, chained_data_delayed_31__19_, chained_data_delayed_31__18_, chained_data_delayed_31__17_, chained_data_delayed_31__16_, chained_data_delayed_31__15_, chained_data_delayed_31__14_, chained_data_delayed_31__13_, chained_data_delayed_31__12_, chained_data_delayed_31__11_, chained_data_delayed_31__10_, chained_data_delayed_31__9_, chained_data_delayed_31__8_, chained_data_delayed_31__7_, chained_data_delayed_31__6_, chained_data_delayed_31__5_, chained_data_delayed_31__4_, chained_data_delayed_31__3_, chained_data_delayed_31__2_, chained_data_delayed_31__1_, chained_data_delayed_31__0_ }),
    .data_o({ chained_data_delayed_32__127_, chained_data_delayed_32__126_, chained_data_delayed_32__125_, chained_data_delayed_32__124_, chained_data_delayed_32__123_, chained_data_delayed_32__122_, chained_data_delayed_32__121_, chained_data_delayed_32__120_, chained_data_delayed_32__119_, chained_data_delayed_32__118_, chained_data_delayed_32__117_, chained_data_delayed_32__116_, chained_data_delayed_32__115_, chained_data_delayed_32__114_, chained_data_delayed_32__113_, chained_data_delayed_32__112_, chained_data_delayed_32__111_, chained_data_delayed_32__110_, chained_data_delayed_32__109_, chained_data_delayed_32__108_, chained_data_delayed_32__107_, chained_data_delayed_32__106_, chained_data_delayed_32__105_, chained_data_delayed_32__104_, chained_data_delayed_32__103_, chained_data_delayed_32__102_, chained_data_delayed_32__101_, chained_data_delayed_32__100_, chained_data_delayed_32__99_, chained_data_delayed_32__98_, chained_data_delayed_32__97_, chained_data_delayed_32__96_, chained_data_delayed_32__95_, chained_data_delayed_32__94_, chained_data_delayed_32__93_, chained_data_delayed_32__92_, chained_data_delayed_32__91_, chained_data_delayed_32__90_, chained_data_delayed_32__89_, chained_data_delayed_32__88_, chained_data_delayed_32__87_, chained_data_delayed_32__86_, chained_data_delayed_32__85_, chained_data_delayed_32__84_, chained_data_delayed_32__83_, chained_data_delayed_32__82_, chained_data_delayed_32__81_, chained_data_delayed_32__80_, chained_data_delayed_32__79_, chained_data_delayed_32__78_, chained_data_delayed_32__77_, chained_data_delayed_32__76_, chained_data_delayed_32__75_, chained_data_delayed_32__74_, chained_data_delayed_32__73_, chained_data_delayed_32__72_, chained_data_delayed_32__71_, chained_data_delayed_32__70_, chained_data_delayed_32__69_, chained_data_delayed_32__68_, chained_data_delayed_32__67_, chained_data_delayed_32__66_, chained_data_delayed_32__65_, chained_data_delayed_32__64_, chained_data_delayed_32__63_, chained_data_delayed_32__62_, chained_data_delayed_32__61_, chained_data_delayed_32__60_, chained_data_delayed_32__59_, chained_data_delayed_32__58_, chained_data_delayed_32__57_, chained_data_delayed_32__56_, chained_data_delayed_32__55_, chained_data_delayed_32__54_, chained_data_delayed_32__53_, chained_data_delayed_32__52_, chained_data_delayed_32__51_, chained_data_delayed_32__50_, chained_data_delayed_32__49_, chained_data_delayed_32__48_, chained_data_delayed_32__47_, chained_data_delayed_32__46_, chained_data_delayed_32__45_, chained_data_delayed_32__44_, chained_data_delayed_32__43_, chained_data_delayed_32__42_, chained_data_delayed_32__41_, chained_data_delayed_32__40_, chained_data_delayed_32__39_, chained_data_delayed_32__38_, chained_data_delayed_32__37_, chained_data_delayed_32__36_, chained_data_delayed_32__35_, chained_data_delayed_32__34_, chained_data_delayed_32__33_, chained_data_delayed_32__32_, chained_data_delayed_32__31_, chained_data_delayed_32__30_, chained_data_delayed_32__29_, chained_data_delayed_32__28_, chained_data_delayed_32__27_, chained_data_delayed_32__26_, chained_data_delayed_32__25_, chained_data_delayed_32__24_, chained_data_delayed_32__23_, chained_data_delayed_32__22_, chained_data_delayed_32__21_, chained_data_delayed_32__20_, chained_data_delayed_32__19_, chained_data_delayed_32__18_, chained_data_delayed_32__17_, chained_data_delayed_32__16_, chained_data_delayed_32__15_, chained_data_delayed_32__14_, chained_data_delayed_32__13_, chained_data_delayed_32__12_, chained_data_delayed_32__11_, chained_data_delayed_32__10_, chained_data_delayed_32__9_, chained_data_delayed_32__8_, chained_data_delayed_32__7_, chained_data_delayed_32__6_, chained_data_delayed_32__5_, chained_data_delayed_32__4_, chained_data_delayed_32__3_, chained_data_delayed_32__2_, chained_data_delayed_32__1_, chained_data_delayed_32__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_33__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_32__127_, chained_data_delayed_32__126_, chained_data_delayed_32__125_, chained_data_delayed_32__124_, chained_data_delayed_32__123_, chained_data_delayed_32__122_, chained_data_delayed_32__121_, chained_data_delayed_32__120_, chained_data_delayed_32__119_, chained_data_delayed_32__118_, chained_data_delayed_32__117_, chained_data_delayed_32__116_, chained_data_delayed_32__115_, chained_data_delayed_32__114_, chained_data_delayed_32__113_, chained_data_delayed_32__112_, chained_data_delayed_32__111_, chained_data_delayed_32__110_, chained_data_delayed_32__109_, chained_data_delayed_32__108_, chained_data_delayed_32__107_, chained_data_delayed_32__106_, chained_data_delayed_32__105_, chained_data_delayed_32__104_, chained_data_delayed_32__103_, chained_data_delayed_32__102_, chained_data_delayed_32__101_, chained_data_delayed_32__100_, chained_data_delayed_32__99_, chained_data_delayed_32__98_, chained_data_delayed_32__97_, chained_data_delayed_32__96_, chained_data_delayed_32__95_, chained_data_delayed_32__94_, chained_data_delayed_32__93_, chained_data_delayed_32__92_, chained_data_delayed_32__91_, chained_data_delayed_32__90_, chained_data_delayed_32__89_, chained_data_delayed_32__88_, chained_data_delayed_32__87_, chained_data_delayed_32__86_, chained_data_delayed_32__85_, chained_data_delayed_32__84_, chained_data_delayed_32__83_, chained_data_delayed_32__82_, chained_data_delayed_32__81_, chained_data_delayed_32__80_, chained_data_delayed_32__79_, chained_data_delayed_32__78_, chained_data_delayed_32__77_, chained_data_delayed_32__76_, chained_data_delayed_32__75_, chained_data_delayed_32__74_, chained_data_delayed_32__73_, chained_data_delayed_32__72_, chained_data_delayed_32__71_, chained_data_delayed_32__70_, chained_data_delayed_32__69_, chained_data_delayed_32__68_, chained_data_delayed_32__67_, chained_data_delayed_32__66_, chained_data_delayed_32__65_, chained_data_delayed_32__64_, chained_data_delayed_32__63_, chained_data_delayed_32__62_, chained_data_delayed_32__61_, chained_data_delayed_32__60_, chained_data_delayed_32__59_, chained_data_delayed_32__58_, chained_data_delayed_32__57_, chained_data_delayed_32__56_, chained_data_delayed_32__55_, chained_data_delayed_32__54_, chained_data_delayed_32__53_, chained_data_delayed_32__52_, chained_data_delayed_32__51_, chained_data_delayed_32__50_, chained_data_delayed_32__49_, chained_data_delayed_32__48_, chained_data_delayed_32__47_, chained_data_delayed_32__46_, chained_data_delayed_32__45_, chained_data_delayed_32__44_, chained_data_delayed_32__43_, chained_data_delayed_32__42_, chained_data_delayed_32__41_, chained_data_delayed_32__40_, chained_data_delayed_32__39_, chained_data_delayed_32__38_, chained_data_delayed_32__37_, chained_data_delayed_32__36_, chained_data_delayed_32__35_, chained_data_delayed_32__34_, chained_data_delayed_32__33_, chained_data_delayed_32__32_, chained_data_delayed_32__31_, chained_data_delayed_32__30_, chained_data_delayed_32__29_, chained_data_delayed_32__28_, chained_data_delayed_32__27_, chained_data_delayed_32__26_, chained_data_delayed_32__25_, chained_data_delayed_32__24_, chained_data_delayed_32__23_, chained_data_delayed_32__22_, chained_data_delayed_32__21_, chained_data_delayed_32__20_, chained_data_delayed_32__19_, chained_data_delayed_32__18_, chained_data_delayed_32__17_, chained_data_delayed_32__16_, chained_data_delayed_32__15_, chained_data_delayed_32__14_, chained_data_delayed_32__13_, chained_data_delayed_32__12_, chained_data_delayed_32__11_, chained_data_delayed_32__10_, chained_data_delayed_32__9_, chained_data_delayed_32__8_, chained_data_delayed_32__7_, chained_data_delayed_32__6_, chained_data_delayed_32__5_, chained_data_delayed_32__4_, chained_data_delayed_32__3_, chained_data_delayed_32__2_, chained_data_delayed_32__1_, chained_data_delayed_32__0_ }),
    .data_o({ chained_data_delayed_33__127_, chained_data_delayed_33__126_, chained_data_delayed_33__125_, chained_data_delayed_33__124_, chained_data_delayed_33__123_, chained_data_delayed_33__122_, chained_data_delayed_33__121_, chained_data_delayed_33__120_, chained_data_delayed_33__119_, chained_data_delayed_33__118_, chained_data_delayed_33__117_, chained_data_delayed_33__116_, chained_data_delayed_33__115_, chained_data_delayed_33__114_, chained_data_delayed_33__113_, chained_data_delayed_33__112_, chained_data_delayed_33__111_, chained_data_delayed_33__110_, chained_data_delayed_33__109_, chained_data_delayed_33__108_, chained_data_delayed_33__107_, chained_data_delayed_33__106_, chained_data_delayed_33__105_, chained_data_delayed_33__104_, chained_data_delayed_33__103_, chained_data_delayed_33__102_, chained_data_delayed_33__101_, chained_data_delayed_33__100_, chained_data_delayed_33__99_, chained_data_delayed_33__98_, chained_data_delayed_33__97_, chained_data_delayed_33__96_, chained_data_delayed_33__95_, chained_data_delayed_33__94_, chained_data_delayed_33__93_, chained_data_delayed_33__92_, chained_data_delayed_33__91_, chained_data_delayed_33__90_, chained_data_delayed_33__89_, chained_data_delayed_33__88_, chained_data_delayed_33__87_, chained_data_delayed_33__86_, chained_data_delayed_33__85_, chained_data_delayed_33__84_, chained_data_delayed_33__83_, chained_data_delayed_33__82_, chained_data_delayed_33__81_, chained_data_delayed_33__80_, chained_data_delayed_33__79_, chained_data_delayed_33__78_, chained_data_delayed_33__77_, chained_data_delayed_33__76_, chained_data_delayed_33__75_, chained_data_delayed_33__74_, chained_data_delayed_33__73_, chained_data_delayed_33__72_, chained_data_delayed_33__71_, chained_data_delayed_33__70_, chained_data_delayed_33__69_, chained_data_delayed_33__68_, chained_data_delayed_33__67_, chained_data_delayed_33__66_, chained_data_delayed_33__65_, chained_data_delayed_33__64_, chained_data_delayed_33__63_, chained_data_delayed_33__62_, chained_data_delayed_33__61_, chained_data_delayed_33__60_, chained_data_delayed_33__59_, chained_data_delayed_33__58_, chained_data_delayed_33__57_, chained_data_delayed_33__56_, chained_data_delayed_33__55_, chained_data_delayed_33__54_, chained_data_delayed_33__53_, chained_data_delayed_33__52_, chained_data_delayed_33__51_, chained_data_delayed_33__50_, chained_data_delayed_33__49_, chained_data_delayed_33__48_, chained_data_delayed_33__47_, chained_data_delayed_33__46_, chained_data_delayed_33__45_, chained_data_delayed_33__44_, chained_data_delayed_33__43_, chained_data_delayed_33__42_, chained_data_delayed_33__41_, chained_data_delayed_33__40_, chained_data_delayed_33__39_, chained_data_delayed_33__38_, chained_data_delayed_33__37_, chained_data_delayed_33__36_, chained_data_delayed_33__35_, chained_data_delayed_33__34_, chained_data_delayed_33__33_, chained_data_delayed_33__32_, chained_data_delayed_33__31_, chained_data_delayed_33__30_, chained_data_delayed_33__29_, chained_data_delayed_33__28_, chained_data_delayed_33__27_, chained_data_delayed_33__26_, chained_data_delayed_33__25_, chained_data_delayed_33__24_, chained_data_delayed_33__23_, chained_data_delayed_33__22_, chained_data_delayed_33__21_, chained_data_delayed_33__20_, chained_data_delayed_33__19_, chained_data_delayed_33__18_, chained_data_delayed_33__17_, chained_data_delayed_33__16_, chained_data_delayed_33__15_, chained_data_delayed_33__14_, chained_data_delayed_33__13_, chained_data_delayed_33__12_, chained_data_delayed_33__11_, chained_data_delayed_33__10_, chained_data_delayed_33__9_, chained_data_delayed_33__8_, chained_data_delayed_33__7_, chained_data_delayed_33__6_, chained_data_delayed_33__5_, chained_data_delayed_33__4_, chained_data_delayed_33__3_, chained_data_delayed_33__2_, chained_data_delayed_33__1_, chained_data_delayed_33__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_34__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_33__127_, chained_data_delayed_33__126_, chained_data_delayed_33__125_, chained_data_delayed_33__124_, chained_data_delayed_33__123_, chained_data_delayed_33__122_, chained_data_delayed_33__121_, chained_data_delayed_33__120_, chained_data_delayed_33__119_, chained_data_delayed_33__118_, chained_data_delayed_33__117_, chained_data_delayed_33__116_, chained_data_delayed_33__115_, chained_data_delayed_33__114_, chained_data_delayed_33__113_, chained_data_delayed_33__112_, chained_data_delayed_33__111_, chained_data_delayed_33__110_, chained_data_delayed_33__109_, chained_data_delayed_33__108_, chained_data_delayed_33__107_, chained_data_delayed_33__106_, chained_data_delayed_33__105_, chained_data_delayed_33__104_, chained_data_delayed_33__103_, chained_data_delayed_33__102_, chained_data_delayed_33__101_, chained_data_delayed_33__100_, chained_data_delayed_33__99_, chained_data_delayed_33__98_, chained_data_delayed_33__97_, chained_data_delayed_33__96_, chained_data_delayed_33__95_, chained_data_delayed_33__94_, chained_data_delayed_33__93_, chained_data_delayed_33__92_, chained_data_delayed_33__91_, chained_data_delayed_33__90_, chained_data_delayed_33__89_, chained_data_delayed_33__88_, chained_data_delayed_33__87_, chained_data_delayed_33__86_, chained_data_delayed_33__85_, chained_data_delayed_33__84_, chained_data_delayed_33__83_, chained_data_delayed_33__82_, chained_data_delayed_33__81_, chained_data_delayed_33__80_, chained_data_delayed_33__79_, chained_data_delayed_33__78_, chained_data_delayed_33__77_, chained_data_delayed_33__76_, chained_data_delayed_33__75_, chained_data_delayed_33__74_, chained_data_delayed_33__73_, chained_data_delayed_33__72_, chained_data_delayed_33__71_, chained_data_delayed_33__70_, chained_data_delayed_33__69_, chained_data_delayed_33__68_, chained_data_delayed_33__67_, chained_data_delayed_33__66_, chained_data_delayed_33__65_, chained_data_delayed_33__64_, chained_data_delayed_33__63_, chained_data_delayed_33__62_, chained_data_delayed_33__61_, chained_data_delayed_33__60_, chained_data_delayed_33__59_, chained_data_delayed_33__58_, chained_data_delayed_33__57_, chained_data_delayed_33__56_, chained_data_delayed_33__55_, chained_data_delayed_33__54_, chained_data_delayed_33__53_, chained_data_delayed_33__52_, chained_data_delayed_33__51_, chained_data_delayed_33__50_, chained_data_delayed_33__49_, chained_data_delayed_33__48_, chained_data_delayed_33__47_, chained_data_delayed_33__46_, chained_data_delayed_33__45_, chained_data_delayed_33__44_, chained_data_delayed_33__43_, chained_data_delayed_33__42_, chained_data_delayed_33__41_, chained_data_delayed_33__40_, chained_data_delayed_33__39_, chained_data_delayed_33__38_, chained_data_delayed_33__37_, chained_data_delayed_33__36_, chained_data_delayed_33__35_, chained_data_delayed_33__34_, chained_data_delayed_33__33_, chained_data_delayed_33__32_, chained_data_delayed_33__31_, chained_data_delayed_33__30_, chained_data_delayed_33__29_, chained_data_delayed_33__28_, chained_data_delayed_33__27_, chained_data_delayed_33__26_, chained_data_delayed_33__25_, chained_data_delayed_33__24_, chained_data_delayed_33__23_, chained_data_delayed_33__22_, chained_data_delayed_33__21_, chained_data_delayed_33__20_, chained_data_delayed_33__19_, chained_data_delayed_33__18_, chained_data_delayed_33__17_, chained_data_delayed_33__16_, chained_data_delayed_33__15_, chained_data_delayed_33__14_, chained_data_delayed_33__13_, chained_data_delayed_33__12_, chained_data_delayed_33__11_, chained_data_delayed_33__10_, chained_data_delayed_33__9_, chained_data_delayed_33__8_, chained_data_delayed_33__7_, chained_data_delayed_33__6_, chained_data_delayed_33__5_, chained_data_delayed_33__4_, chained_data_delayed_33__3_, chained_data_delayed_33__2_, chained_data_delayed_33__1_, chained_data_delayed_33__0_ }),
    .data_o({ chained_data_delayed_34__127_, chained_data_delayed_34__126_, chained_data_delayed_34__125_, chained_data_delayed_34__124_, chained_data_delayed_34__123_, chained_data_delayed_34__122_, chained_data_delayed_34__121_, chained_data_delayed_34__120_, chained_data_delayed_34__119_, chained_data_delayed_34__118_, chained_data_delayed_34__117_, chained_data_delayed_34__116_, chained_data_delayed_34__115_, chained_data_delayed_34__114_, chained_data_delayed_34__113_, chained_data_delayed_34__112_, chained_data_delayed_34__111_, chained_data_delayed_34__110_, chained_data_delayed_34__109_, chained_data_delayed_34__108_, chained_data_delayed_34__107_, chained_data_delayed_34__106_, chained_data_delayed_34__105_, chained_data_delayed_34__104_, chained_data_delayed_34__103_, chained_data_delayed_34__102_, chained_data_delayed_34__101_, chained_data_delayed_34__100_, chained_data_delayed_34__99_, chained_data_delayed_34__98_, chained_data_delayed_34__97_, chained_data_delayed_34__96_, chained_data_delayed_34__95_, chained_data_delayed_34__94_, chained_data_delayed_34__93_, chained_data_delayed_34__92_, chained_data_delayed_34__91_, chained_data_delayed_34__90_, chained_data_delayed_34__89_, chained_data_delayed_34__88_, chained_data_delayed_34__87_, chained_data_delayed_34__86_, chained_data_delayed_34__85_, chained_data_delayed_34__84_, chained_data_delayed_34__83_, chained_data_delayed_34__82_, chained_data_delayed_34__81_, chained_data_delayed_34__80_, chained_data_delayed_34__79_, chained_data_delayed_34__78_, chained_data_delayed_34__77_, chained_data_delayed_34__76_, chained_data_delayed_34__75_, chained_data_delayed_34__74_, chained_data_delayed_34__73_, chained_data_delayed_34__72_, chained_data_delayed_34__71_, chained_data_delayed_34__70_, chained_data_delayed_34__69_, chained_data_delayed_34__68_, chained_data_delayed_34__67_, chained_data_delayed_34__66_, chained_data_delayed_34__65_, chained_data_delayed_34__64_, chained_data_delayed_34__63_, chained_data_delayed_34__62_, chained_data_delayed_34__61_, chained_data_delayed_34__60_, chained_data_delayed_34__59_, chained_data_delayed_34__58_, chained_data_delayed_34__57_, chained_data_delayed_34__56_, chained_data_delayed_34__55_, chained_data_delayed_34__54_, chained_data_delayed_34__53_, chained_data_delayed_34__52_, chained_data_delayed_34__51_, chained_data_delayed_34__50_, chained_data_delayed_34__49_, chained_data_delayed_34__48_, chained_data_delayed_34__47_, chained_data_delayed_34__46_, chained_data_delayed_34__45_, chained_data_delayed_34__44_, chained_data_delayed_34__43_, chained_data_delayed_34__42_, chained_data_delayed_34__41_, chained_data_delayed_34__40_, chained_data_delayed_34__39_, chained_data_delayed_34__38_, chained_data_delayed_34__37_, chained_data_delayed_34__36_, chained_data_delayed_34__35_, chained_data_delayed_34__34_, chained_data_delayed_34__33_, chained_data_delayed_34__32_, chained_data_delayed_34__31_, chained_data_delayed_34__30_, chained_data_delayed_34__29_, chained_data_delayed_34__28_, chained_data_delayed_34__27_, chained_data_delayed_34__26_, chained_data_delayed_34__25_, chained_data_delayed_34__24_, chained_data_delayed_34__23_, chained_data_delayed_34__22_, chained_data_delayed_34__21_, chained_data_delayed_34__20_, chained_data_delayed_34__19_, chained_data_delayed_34__18_, chained_data_delayed_34__17_, chained_data_delayed_34__16_, chained_data_delayed_34__15_, chained_data_delayed_34__14_, chained_data_delayed_34__13_, chained_data_delayed_34__12_, chained_data_delayed_34__11_, chained_data_delayed_34__10_, chained_data_delayed_34__9_, chained_data_delayed_34__8_, chained_data_delayed_34__7_, chained_data_delayed_34__6_, chained_data_delayed_34__5_, chained_data_delayed_34__4_, chained_data_delayed_34__3_, chained_data_delayed_34__2_, chained_data_delayed_34__1_, chained_data_delayed_34__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_35__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_34__127_, chained_data_delayed_34__126_, chained_data_delayed_34__125_, chained_data_delayed_34__124_, chained_data_delayed_34__123_, chained_data_delayed_34__122_, chained_data_delayed_34__121_, chained_data_delayed_34__120_, chained_data_delayed_34__119_, chained_data_delayed_34__118_, chained_data_delayed_34__117_, chained_data_delayed_34__116_, chained_data_delayed_34__115_, chained_data_delayed_34__114_, chained_data_delayed_34__113_, chained_data_delayed_34__112_, chained_data_delayed_34__111_, chained_data_delayed_34__110_, chained_data_delayed_34__109_, chained_data_delayed_34__108_, chained_data_delayed_34__107_, chained_data_delayed_34__106_, chained_data_delayed_34__105_, chained_data_delayed_34__104_, chained_data_delayed_34__103_, chained_data_delayed_34__102_, chained_data_delayed_34__101_, chained_data_delayed_34__100_, chained_data_delayed_34__99_, chained_data_delayed_34__98_, chained_data_delayed_34__97_, chained_data_delayed_34__96_, chained_data_delayed_34__95_, chained_data_delayed_34__94_, chained_data_delayed_34__93_, chained_data_delayed_34__92_, chained_data_delayed_34__91_, chained_data_delayed_34__90_, chained_data_delayed_34__89_, chained_data_delayed_34__88_, chained_data_delayed_34__87_, chained_data_delayed_34__86_, chained_data_delayed_34__85_, chained_data_delayed_34__84_, chained_data_delayed_34__83_, chained_data_delayed_34__82_, chained_data_delayed_34__81_, chained_data_delayed_34__80_, chained_data_delayed_34__79_, chained_data_delayed_34__78_, chained_data_delayed_34__77_, chained_data_delayed_34__76_, chained_data_delayed_34__75_, chained_data_delayed_34__74_, chained_data_delayed_34__73_, chained_data_delayed_34__72_, chained_data_delayed_34__71_, chained_data_delayed_34__70_, chained_data_delayed_34__69_, chained_data_delayed_34__68_, chained_data_delayed_34__67_, chained_data_delayed_34__66_, chained_data_delayed_34__65_, chained_data_delayed_34__64_, chained_data_delayed_34__63_, chained_data_delayed_34__62_, chained_data_delayed_34__61_, chained_data_delayed_34__60_, chained_data_delayed_34__59_, chained_data_delayed_34__58_, chained_data_delayed_34__57_, chained_data_delayed_34__56_, chained_data_delayed_34__55_, chained_data_delayed_34__54_, chained_data_delayed_34__53_, chained_data_delayed_34__52_, chained_data_delayed_34__51_, chained_data_delayed_34__50_, chained_data_delayed_34__49_, chained_data_delayed_34__48_, chained_data_delayed_34__47_, chained_data_delayed_34__46_, chained_data_delayed_34__45_, chained_data_delayed_34__44_, chained_data_delayed_34__43_, chained_data_delayed_34__42_, chained_data_delayed_34__41_, chained_data_delayed_34__40_, chained_data_delayed_34__39_, chained_data_delayed_34__38_, chained_data_delayed_34__37_, chained_data_delayed_34__36_, chained_data_delayed_34__35_, chained_data_delayed_34__34_, chained_data_delayed_34__33_, chained_data_delayed_34__32_, chained_data_delayed_34__31_, chained_data_delayed_34__30_, chained_data_delayed_34__29_, chained_data_delayed_34__28_, chained_data_delayed_34__27_, chained_data_delayed_34__26_, chained_data_delayed_34__25_, chained_data_delayed_34__24_, chained_data_delayed_34__23_, chained_data_delayed_34__22_, chained_data_delayed_34__21_, chained_data_delayed_34__20_, chained_data_delayed_34__19_, chained_data_delayed_34__18_, chained_data_delayed_34__17_, chained_data_delayed_34__16_, chained_data_delayed_34__15_, chained_data_delayed_34__14_, chained_data_delayed_34__13_, chained_data_delayed_34__12_, chained_data_delayed_34__11_, chained_data_delayed_34__10_, chained_data_delayed_34__9_, chained_data_delayed_34__8_, chained_data_delayed_34__7_, chained_data_delayed_34__6_, chained_data_delayed_34__5_, chained_data_delayed_34__4_, chained_data_delayed_34__3_, chained_data_delayed_34__2_, chained_data_delayed_34__1_, chained_data_delayed_34__0_ }),
    .data_o({ chained_data_delayed_35__127_, chained_data_delayed_35__126_, chained_data_delayed_35__125_, chained_data_delayed_35__124_, chained_data_delayed_35__123_, chained_data_delayed_35__122_, chained_data_delayed_35__121_, chained_data_delayed_35__120_, chained_data_delayed_35__119_, chained_data_delayed_35__118_, chained_data_delayed_35__117_, chained_data_delayed_35__116_, chained_data_delayed_35__115_, chained_data_delayed_35__114_, chained_data_delayed_35__113_, chained_data_delayed_35__112_, chained_data_delayed_35__111_, chained_data_delayed_35__110_, chained_data_delayed_35__109_, chained_data_delayed_35__108_, chained_data_delayed_35__107_, chained_data_delayed_35__106_, chained_data_delayed_35__105_, chained_data_delayed_35__104_, chained_data_delayed_35__103_, chained_data_delayed_35__102_, chained_data_delayed_35__101_, chained_data_delayed_35__100_, chained_data_delayed_35__99_, chained_data_delayed_35__98_, chained_data_delayed_35__97_, chained_data_delayed_35__96_, chained_data_delayed_35__95_, chained_data_delayed_35__94_, chained_data_delayed_35__93_, chained_data_delayed_35__92_, chained_data_delayed_35__91_, chained_data_delayed_35__90_, chained_data_delayed_35__89_, chained_data_delayed_35__88_, chained_data_delayed_35__87_, chained_data_delayed_35__86_, chained_data_delayed_35__85_, chained_data_delayed_35__84_, chained_data_delayed_35__83_, chained_data_delayed_35__82_, chained_data_delayed_35__81_, chained_data_delayed_35__80_, chained_data_delayed_35__79_, chained_data_delayed_35__78_, chained_data_delayed_35__77_, chained_data_delayed_35__76_, chained_data_delayed_35__75_, chained_data_delayed_35__74_, chained_data_delayed_35__73_, chained_data_delayed_35__72_, chained_data_delayed_35__71_, chained_data_delayed_35__70_, chained_data_delayed_35__69_, chained_data_delayed_35__68_, chained_data_delayed_35__67_, chained_data_delayed_35__66_, chained_data_delayed_35__65_, chained_data_delayed_35__64_, chained_data_delayed_35__63_, chained_data_delayed_35__62_, chained_data_delayed_35__61_, chained_data_delayed_35__60_, chained_data_delayed_35__59_, chained_data_delayed_35__58_, chained_data_delayed_35__57_, chained_data_delayed_35__56_, chained_data_delayed_35__55_, chained_data_delayed_35__54_, chained_data_delayed_35__53_, chained_data_delayed_35__52_, chained_data_delayed_35__51_, chained_data_delayed_35__50_, chained_data_delayed_35__49_, chained_data_delayed_35__48_, chained_data_delayed_35__47_, chained_data_delayed_35__46_, chained_data_delayed_35__45_, chained_data_delayed_35__44_, chained_data_delayed_35__43_, chained_data_delayed_35__42_, chained_data_delayed_35__41_, chained_data_delayed_35__40_, chained_data_delayed_35__39_, chained_data_delayed_35__38_, chained_data_delayed_35__37_, chained_data_delayed_35__36_, chained_data_delayed_35__35_, chained_data_delayed_35__34_, chained_data_delayed_35__33_, chained_data_delayed_35__32_, chained_data_delayed_35__31_, chained_data_delayed_35__30_, chained_data_delayed_35__29_, chained_data_delayed_35__28_, chained_data_delayed_35__27_, chained_data_delayed_35__26_, chained_data_delayed_35__25_, chained_data_delayed_35__24_, chained_data_delayed_35__23_, chained_data_delayed_35__22_, chained_data_delayed_35__21_, chained_data_delayed_35__20_, chained_data_delayed_35__19_, chained_data_delayed_35__18_, chained_data_delayed_35__17_, chained_data_delayed_35__16_, chained_data_delayed_35__15_, chained_data_delayed_35__14_, chained_data_delayed_35__13_, chained_data_delayed_35__12_, chained_data_delayed_35__11_, chained_data_delayed_35__10_, chained_data_delayed_35__9_, chained_data_delayed_35__8_, chained_data_delayed_35__7_, chained_data_delayed_35__6_, chained_data_delayed_35__5_, chained_data_delayed_35__4_, chained_data_delayed_35__3_, chained_data_delayed_35__2_, chained_data_delayed_35__1_, chained_data_delayed_35__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_36__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_35__127_, chained_data_delayed_35__126_, chained_data_delayed_35__125_, chained_data_delayed_35__124_, chained_data_delayed_35__123_, chained_data_delayed_35__122_, chained_data_delayed_35__121_, chained_data_delayed_35__120_, chained_data_delayed_35__119_, chained_data_delayed_35__118_, chained_data_delayed_35__117_, chained_data_delayed_35__116_, chained_data_delayed_35__115_, chained_data_delayed_35__114_, chained_data_delayed_35__113_, chained_data_delayed_35__112_, chained_data_delayed_35__111_, chained_data_delayed_35__110_, chained_data_delayed_35__109_, chained_data_delayed_35__108_, chained_data_delayed_35__107_, chained_data_delayed_35__106_, chained_data_delayed_35__105_, chained_data_delayed_35__104_, chained_data_delayed_35__103_, chained_data_delayed_35__102_, chained_data_delayed_35__101_, chained_data_delayed_35__100_, chained_data_delayed_35__99_, chained_data_delayed_35__98_, chained_data_delayed_35__97_, chained_data_delayed_35__96_, chained_data_delayed_35__95_, chained_data_delayed_35__94_, chained_data_delayed_35__93_, chained_data_delayed_35__92_, chained_data_delayed_35__91_, chained_data_delayed_35__90_, chained_data_delayed_35__89_, chained_data_delayed_35__88_, chained_data_delayed_35__87_, chained_data_delayed_35__86_, chained_data_delayed_35__85_, chained_data_delayed_35__84_, chained_data_delayed_35__83_, chained_data_delayed_35__82_, chained_data_delayed_35__81_, chained_data_delayed_35__80_, chained_data_delayed_35__79_, chained_data_delayed_35__78_, chained_data_delayed_35__77_, chained_data_delayed_35__76_, chained_data_delayed_35__75_, chained_data_delayed_35__74_, chained_data_delayed_35__73_, chained_data_delayed_35__72_, chained_data_delayed_35__71_, chained_data_delayed_35__70_, chained_data_delayed_35__69_, chained_data_delayed_35__68_, chained_data_delayed_35__67_, chained_data_delayed_35__66_, chained_data_delayed_35__65_, chained_data_delayed_35__64_, chained_data_delayed_35__63_, chained_data_delayed_35__62_, chained_data_delayed_35__61_, chained_data_delayed_35__60_, chained_data_delayed_35__59_, chained_data_delayed_35__58_, chained_data_delayed_35__57_, chained_data_delayed_35__56_, chained_data_delayed_35__55_, chained_data_delayed_35__54_, chained_data_delayed_35__53_, chained_data_delayed_35__52_, chained_data_delayed_35__51_, chained_data_delayed_35__50_, chained_data_delayed_35__49_, chained_data_delayed_35__48_, chained_data_delayed_35__47_, chained_data_delayed_35__46_, chained_data_delayed_35__45_, chained_data_delayed_35__44_, chained_data_delayed_35__43_, chained_data_delayed_35__42_, chained_data_delayed_35__41_, chained_data_delayed_35__40_, chained_data_delayed_35__39_, chained_data_delayed_35__38_, chained_data_delayed_35__37_, chained_data_delayed_35__36_, chained_data_delayed_35__35_, chained_data_delayed_35__34_, chained_data_delayed_35__33_, chained_data_delayed_35__32_, chained_data_delayed_35__31_, chained_data_delayed_35__30_, chained_data_delayed_35__29_, chained_data_delayed_35__28_, chained_data_delayed_35__27_, chained_data_delayed_35__26_, chained_data_delayed_35__25_, chained_data_delayed_35__24_, chained_data_delayed_35__23_, chained_data_delayed_35__22_, chained_data_delayed_35__21_, chained_data_delayed_35__20_, chained_data_delayed_35__19_, chained_data_delayed_35__18_, chained_data_delayed_35__17_, chained_data_delayed_35__16_, chained_data_delayed_35__15_, chained_data_delayed_35__14_, chained_data_delayed_35__13_, chained_data_delayed_35__12_, chained_data_delayed_35__11_, chained_data_delayed_35__10_, chained_data_delayed_35__9_, chained_data_delayed_35__8_, chained_data_delayed_35__7_, chained_data_delayed_35__6_, chained_data_delayed_35__5_, chained_data_delayed_35__4_, chained_data_delayed_35__3_, chained_data_delayed_35__2_, chained_data_delayed_35__1_, chained_data_delayed_35__0_ }),
    .data_o({ chained_data_delayed_36__127_, chained_data_delayed_36__126_, chained_data_delayed_36__125_, chained_data_delayed_36__124_, chained_data_delayed_36__123_, chained_data_delayed_36__122_, chained_data_delayed_36__121_, chained_data_delayed_36__120_, chained_data_delayed_36__119_, chained_data_delayed_36__118_, chained_data_delayed_36__117_, chained_data_delayed_36__116_, chained_data_delayed_36__115_, chained_data_delayed_36__114_, chained_data_delayed_36__113_, chained_data_delayed_36__112_, chained_data_delayed_36__111_, chained_data_delayed_36__110_, chained_data_delayed_36__109_, chained_data_delayed_36__108_, chained_data_delayed_36__107_, chained_data_delayed_36__106_, chained_data_delayed_36__105_, chained_data_delayed_36__104_, chained_data_delayed_36__103_, chained_data_delayed_36__102_, chained_data_delayed_36__101_, chained_data_delayed_36__100_, chained_data_delayed_36__99_, chained_data_delayed_36__98_, chained_data_delayed_36__97_, chained_data_delayed_36__96_, chained_data_delayed_36__95_, chained_data_delayed_36__94_, chained_data_delayed_36__93_, chained_data_delayed_36__92_, chained_data_delayed_36__91_, chained_data_delayed_36__90_, chained_data_delayed_36__89_, chained_data_delayed_36__88_, chained_data_delayed_36__87_, chained_data_delayed_36__86_, chained_data_delayed_36__85_, chained_data_delayed_36__84_, chained_data_delayed_36__83_, chained_data_delayed_36__82_, chained_data_delayed_36__81_, chained_data_delayed_36__80_, chained_data_delayed_36__79_, chained_data_delayed_36__78_, chained_data_delayed_36__77_, chained_data_delayed_36__76_, chained_data_delayed_36__75_, chained_data_delayed_36__74_, chained_data_delayed_36__73_, chained_data_delayed_36__72_, chained_data_delayed_36__71_, chained_data_delayed_36__70_, chained_data_delayed_36__69_, chained_data_delayed_36__68_, chained_data_delayed_36__67_, chained_data_delayed_36__66_, chained_data_delayed_36__65_, chained_data_delayed_36__64_, chained_data_delayed_36__63_, chained_data_delayed_36__62_, chained_data_delayed_36__61_, chained_data_delayed_36__60_, chained_data_delayed_36__59_, chained_data_delayed_36__58_, chained_data_delayed_36__57_, chained_data_delayed_36__56_, chained_data_delayed_36__55_, chained_data_delayed_36__54_, chained_data_delayed_36__53_, chained_data_delayed_36__52_, chained_data_delayed_36__51_, chained_data_delayed_36__50_, chained_data_delayed_36__49_, chained_data_delayed_36__48_, chained_data_delayed_36__47_, chained_data_delayed_36__46_, chained_data_delayed_36__45_, chained_data_delayed_36__44_, chained_data_delayed_36__43_, chained_data_delayed_36__42_, chained_data_delayed_36__41_, chained_data_delayed_36__40_, chained_data_delayed_36__39_, chained_data_delayed_36__38_, chained_data_delayed_36__37_, chained_data_delayed_36__36_, chained_data_delayed_36__35_, chained_data_delayed_36__34_, chained_data_delayed_36__33_, chained_data_delayed_36__32_, chained_data_delayed_36__31_, chained_data_delayed_36__30_, chained_data_delayed_36__29_, chained_data_delayed_36__28_, chained_data_delayed_36__27_, chained_data_delayed_36__26_, chained_data_delayed_36__25_, chained_data_delayed_36__24_, chained_data_delayed_36__23_, chained_data_delayed_36__22_, chained_data_delayed_36__21_, chained_data_delayed_36__20_, chained_data_delayed_36__19_, chained_data_delayed_36__18_, chained_data_delayed_36__17_, chained_data_delayed_36__16_, chained_data_delayed_36__15_, chained_data_delayed_36__14_, chained_data_delayed_36__13_, chained_data_delayed_36__12_, chained_data_delayed_36__11_, chained_data_delayed_36__10_, chained_data_delayed_36__9_, chained_data_delayed_36__8_, chained_data_delayed_36__7_, chained_data_delayed_36__6_, chained_data_delayed_36__5_, chained_data_delayed_36__4_, chained_data_delayed_36__3_, chained_data_delayed_36__2_, chained_data_delayed_36__1_, chained_data_delayed_36__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_37__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_36__127_, chained_data_delayed_36__126_, chained_data_delayed_36__125_, chained_data_delayed_36__124_, chained_data_delayed_36__123_, chained_data_delayed_36__122_, chained_data_delayed_36__121_, chained_data_delayed_36__120_, chained_data_delayed_36__119_, chained_data_delayed_36__118_, chained_data_delayed_36__117_, chained_data_delayed_36__116_, chained_data_delayed_36__115_, chained_data_delayed_36__114_, chained_data_delayed_36__113_, chained_data_delayed_36__112_, chained_data_delayed_36__111_, chained_data_delayed_36__110_, chained_data_delayed_36__109_, chained_data_delayed_36__108_, chained_data_delayed_36__107_, chained_data_delayed_36__106_, chained_data_delayed_36__105_, chained_data_delayed_36__104_, chained_data_delayed_36__103_, chained_data_delayed_36__102_, chained_data_delayed_36__101_, chained_data_delayed_36__100_, chained_data_delayed_36__99_, chained_data_delayed_36__98_, chained_data_delayed_36__97_, chained_data_delayed_36__96_, chained_data_delayed_36__95_, chained_data_delayed_36__94_, chained_data_delayed_36__93_, chained_data_delayed_36__92_, chained_data_delayed_36__91_, chained_data_delayed_36__90_, chained_data_delayed_36__89_, chained_data_delayed_36__88_, chained_data_delayed_36__87_, chained_data_delayed_36__86_, chained_data_delayed_36__85_, chained_data_delayed_36__84_, chained_data_delayed_36__83_, chained_data_delayed_36__82_, chained_data_delayed_36__81_, chained_data_delayed_36__80_, chained_data_delayed_36__79_, chained_data_delayed_36__78_, chained_data_delayed_36__77_, chained_data_delayed_36__76_, chained_data_delayed_36__75_, chained_data_delayed_36__74_, chained_data_delayed_36__73_, chained_data_delayed_36__72_, chained_data_delayed_36__71_, chained_data_delayed_36__70_, chained_data_delayed_36__69_, chained_data_delayed_36__68_, chained_data_delayed_36__67_, chained_data_delayed_36__66_, chained_data_delayed_36__65_, chained_data_delayed_36__64_, chained_data_delayed_36__63_, chained_data_delayed_36__62_, chained_data_delayed_36__61_, chained_data_delayed_36__60_, chained_data_delayed_36__59_, chained_data_delayed_36__58_, chained_data_delayed_36__57_, chained_data_delayed_36__56_, chained_data_delayed_36__55_, chained_data_delayed_36__54_, chained_data_delayed_36__53_, chained_data_delayed_36__52_, chained_data_delayed_36__51_, chained_data_delayed_36__50_, chained_data_delayed_36__49_, chained_data_delayed_36__48_, chained_data_delayed_36__47_, chained_data_delayed_36__46_, chained_data_delayed_36__45_, chained_data_delayed_36__44_, chained_data_delayed_36__43_, chained_data_delayed_36__42_, chained_data_delayed_36__41_, chained_data_delayed_36__40_, chained_data_delayed_36__39_, chained_data_delayed_36__38_, chained_data_delayed_36__37_, chained_data_delayed_36__36_, chained_data_delayed_36__35_, chained_data_delayed_36__34_, chained_data_delayed_36__33_, chained_data_delayed_36__32_, chained_data_delayed_36__31_, chained_data_delayed_36__30_, chained_data_delayed_36__29_, chained_data_delayed_36__28_, chained_data_delayed_36__27_, chained_data_delayed_36__26_, chained_data_delayed_36__25_, chained_data_delayed_36__24_, chained_data_delayed_36__23_, chained_data_delayed_36__22_, chained_data_delayed_36__21_, chained_data_delayed_36__20_, chained_data_delayed_36__19_, chained_data_delayed_36__18_, chained_data_delayed_36__17_, chained_data_delayed_36__16_, chained_data_delayed_36__15_, chained_data_delayed_36__14_, chained_data_delayed_36__13_, chained_data_delayed_36__12_, chained_data_delayed_36__11_, chained_data_delayed_36__10_, chained_data_delayed_36__9_, chained_data_delayed_36__8_, chained_data_delayed_36__7_, chained_data_delayed_36__6_, chained_data_delayed_36__5_, chained_data_delayed_36__4_, chained_data_delayed_36__3_, chained_data_delayed_36__2_, chained_data_delayed_36__1_, chained_data_delayed_36__0_ }),
    .data_o({ chained_data_delayed_37__127_, chained_data_delayed_37__126_, chained_data_delayed_37__125_, chained_data_delayed_37__124_, chained_data_delayed_37__123_, chained_data_delayed_37__122_, chained_data_delayed_37__121_, chained_data_delayed_37__120_, chained_data_delayed_37__119_, chained_data_delayed_37__118_, chained_data_delayed_37__117_, chained_data_delayed_37__116_, chained_data_delayed_37__115_, chained_data_delayed_37__114_, chained_data_delayed_37__113_, chained_data_delayed_37__112_, chained_data_delayed_37__111_, chained_data_delayed_37__110_, chained_data_delayed_37__109_, chained_data_delayed_37__108_, chained_data_delayed_37__107_, chained_data_delayed_37__106_, chained_data_delayed_37__105_, chained_data_delayed_37__104_, chained_data_delayed_37__103_, chained_data_delayed_37__102_, chained_data_delayed_37__101_, chained_data_delayed_37__100_, chained_data_delayed_37__99_, chained_data_delayed_37__98_, chained_data_delayed_37__97_, chained_data_delayed_37__96_, chained_data_delayed_37__95_, chained_data_delayed_37__94_, chained_data_delayed_37__93_, chained_data_delayed_37__92_, chained_data_delayed_37__91_, chained_data_delayed_37__90_, chained_data_delayed_37__89_, chained_data_delayed_37__88_, chained_data_delayed_37__87_, chained_data_delayed_37__86_, chained_data_delayed_37__85_, chained_data_delayed_37__84_, chained_data_delayed_37__83_, chained_data_delayed_37__82_, chained_data_delayed_37__81_, chained_data_delayed_37__80_, chained_data_delayed_37__79_, chained_data_delayed_37__78_, chained_data_delayed_37__77_, chained_data_delayed_37__76_, chained_data_delayed_37__75_, chained_data_delayed_37__74_, chained_data_delayed_37__73_, chained_data_delayed_37__72_, chained_data_delayed_37__71_, chained_data_delayed_37__70_, chained_data_delayed_37__69_, chained_data_delayed_37__68_, chained_data_delayed_37__67_, chained_data_delayed_37__66_, chained_data_delayed_37__65_, chained_data_delayed_37__64_, chained_data_delayed_37__63_, chained_data_delayed_37__62_, chained_data_delayed_37__61_, chained_data_delayed_37__60_, chained_data_delayed_37__59_, chained_data_delayed_37__58_, chained_data_delayed_37__57_, chained_data_delayed_37__56_, chained_data_delayed_37__55_, chained_data_delayed_37__54_, chained_data_delayed_37__53_, chained_data_delayed_37__52_, chained_data_delayed_37__51_, chained_data_delayed_37__50_, chained_data_delayed_37__49_, chained_data_delayed_37__48_, chained_data_delayed_37__47_, chained_data_delayed_37__46_, chained_data_delayed_37__45_, chained_data_delayed_37__44_, chained_data_delayed_37__43_, chained_data_delayed_37__42_, chained_data_delayed_37__41_, chained_data_delayed_37__40_, chained_data_delayed_37__39_, chained_data_delayed_37__38_, chained_data_delayed_37__37_, chained_data_delayed_37__36_, chained_data_delayed_37__35_, chained_data_delayed_37__34_, chained_data_delayed_37__33_, chained_data_delayed_37__32_, chained_data_delayed_37__31_, chained_data_delayed_37__30_, chained_data_delayed_37__29_, chained_data_delayed_37__28_, chained_data_delayed_37__27_, chained_data_delayed_37__26_, chained_data_delayed_37__25_, chained_data_delayed_37__24_, chained_data_delayed_37__23_, chained_data_delayed_37__22_, chained_data_delayed_37__21_, chained_data_delayed_37__20_, chained_data_delayed_37__19_, chained_data_delayed_37__18_, chained_data_delayed_37__17_, chained_data_delayed_37__16_, chained_data_delayed_37__15_, chained_data_delayed_37__14_, chained_data_delayed_37__13_, chained_data_delayed_37__12_, chained_data_delayed_37__11_, chained_data_delayed_37__10_, chained_data_delayed_37__9_, chained_data_delayed_37__8_, chained_data_delayed_37__7_, chained_data_delayed_37__6_, chained_data_delayed_37__5_, chained_data_delayed_37__4_, chained_data_delayed_37__3_, chained_data_delayed_37__2_, chained_data_delayed_37__1_, chained_data_delayed_37__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_38__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_37__127_, chained_data_delayed_37__126_, chained_data_delayed_37__125_, chained_data_delayed_37__124_, chained_data_delayed_37__123_, chained_data_delayed_37__122_, chained_data_delayed_37__121_, chained_data_delayed_37__120_, chained_data_delayed_37__119_, chained_data_delayed_37__118_, chained_data_delayed_37__117_, chained_data_delayed_37__116_, chained_data_delayed_37__115_, chained_data_delayed_37__114_, chained_data_delayed_37__113_, chained_data_delayed_37__112_, chained_data_delayed_37__111_, chained_data_delayed_37__110_, chained_data_delayed_37__109_, chained_data_delayed_37__108_, chained_data_delayed_37__107_, chained_data_delayed_37__106_, chained_data_delayed_37__105_, chained_data_delayed_37__104_, chained_data_delayed_37__103_, chained_data_delayed_37__102_, chained_data_delayed_37__101_, chained_data_delayed_37__100_, chained_data_delayed_37__99_, chained_data_delayed_37__98_, chained_data_delayed_37__97_, chained_data_delayed_37__96_, chained_data_delayed_37__95_, chained_data_delayed_37__94_, chained_data_delayed_37__93_, chained_data_delayed_37__92_, chained_data_delayed_37__91_, chained_data_delayed_37__90_, chained_data_delayed_37__89_, chained_data_delayed_37__88_, chained_data_delayed_37__87_, chained_data_delayed_37__86_, chained_data_delayed_37__85_, chained_data_delayed_37__84_, chained_data_delayed_37__83_, chained_data_delayed_37__82_, chained_data_delayed_37__81_, chained_data_delayed_37__80_, chained_data_delayed_37__79_, chained_data_delayed_37__78_, chained_data_delayed_37__77_, chained_data_delayed_37__76_, chained_data_delayed_37__75_, chained_data_delayed_37__74_, chained_data_delayed_37__73_, chained_data_delayed_37__72_, chained_data_delayed_37__71_, chained_data_delayed_37__70_, chained_data_delayed_37__69_, chained_data_delayed_37__68_, chained_data_delayed_37__67_, chained_data_delayed_37__66_, chained_data_delayed_37__65_, chained_data_delayed_37__64_, chained_data_delayed_37__63_, chained_data_delayed_37__62_, chained_data_delayed_37__61_, chained_data_delayed_37__60_, chained_data_delayed_37__59_, chained_data_delayed_37__58_, chained_data_delayed_37__57_, chained_data_delayed_37__56_, chained_data_delayed_37__55_, chained_data_delayed_37__54_, chained_data_delayed_37__53_, chained_data_delayed_37__52_, chained_data_delayed_37__51_, chained_data_delayed_37__50_, chained_data_delayed_37__49_, chained_data_delayed_37__48_, chained_data_delayed_37__47_, chained_data_delayed_37__46_, chained_data_delayed_37__45_, chained_data_delayed_37__44_, chained_data_delayed_37__43_, chained_data_delayed_37__42_, chained_data_delayed_37__41_, chained_data_delayed_37__40_, chained_data_delayed_37__39_, chained_data_delayed_37__38_, chained_data_delayed_37__37_, chained_data_delayed_37__36_, chained_data_delayed_37__35_, chained_data_delayed_37__34_, chained_data_delayed_37__33_, chained_data_delayed_37__32_, chained_data_delayed_37__31_, chained_data_delayed_37__30_, chained_data_delayed_37__29_, chained_data_delayed_37__28_, chained_data_delayed_37__27_, chained_data_delayed_37__26_, chained_data_delayed_37__25_, chained_data_delayed_37__24_, chained_data_delayed_37__23_, chained_data_delayed_37__22_, chained_data_delayed_37__21_, chained_data_delayed_37__20_, chained_data_delayed_37__19_, chained_data_delayed_37__18_, chained_data_delayed_37__17_, chained_data_delayed_37__16_, chained_data_delayed_37__15_, chained_data_delayed_37__14_, chained_data_delayed_37__13_, chained_data_delayed_37__12_, chained_data_delayed_37__11_, chained_data_delayed_37__10_, chained_data_delayed_37__9_, chained_data_delayed_37__8_, chained_data_delayed_37__7_, chained_data_delayed_37__6_, chained_data_delayed_37__5_, chained_data_delayed_37__4_, chained_data_delayed_37__3_, chained_data_delayed_37__2_, chained_data_delayed_37__1_, chained_data_delayed_37__0_ }),
    .data_o({ chained_data_delayed_38__127_, chained_data_delayed_38__126_, chained_data_delayed_38__125_, chained_data_delayed_38__124_, chained_data_delayed_38__123_, chained_data_delayed_38__122_, chained_data_delayed_38__121_, chained_data_delayed_38__120_, chained_data_delayed_38__119_, chained_data_delayed_38__118_, chained_data_delayed_38__117_, chained_data_delayed_38__116_, chained_data_delayed_38__115_, chained_data_delayed_38__114_, chained_data_delayed_38__113_, chained_data_delayed_38__112_, chained_data_delayed_38__111_, chained_data_delayed_38__110_, chained_data_delayed_38__109_, chained_data_delayed_38__108_, chained_data_delayed_38__107_, chained_data_delayed_38__106_, chained_data_delayed_38__105_, chained_data_delayed_38__104_, chained_data_delayed_38__103_, chained_data_delayed_38__102_, chained_data_delayed_38__101_, chained_data_delayed_38__100_, chained_data_delayed_38__99_, chained_data_delayed_38__98_, chained_data_delayed_38__97_, chained_data_delayed_38__96_, chained_data_delayed_38__95_, chained_data_delayed_38__94_, chained_data_delayed_38__93_, chained_data_delayed_38__92_, chained_data_delayed_38__91_, chained_data_delayed_38__90_, chained_data_delayed_38__89_, chained_data_delayed_38__88_, chained_data_delayed_38__87_, chained_data_delayed_38__86_, chained_data_delayed_38__85_, chained_data_delayed_38__84_, chained_data_delayed_38__83_, chained_data_delayed_38__82_, chained_data_delayed_38__81_, chained_data_delayed_38__80_, chained_data_delayed_38__79_, chained_data_delayed_38__78_, chained_data_delayed_38__77_, chained_data_delayed_38__76_, chained_data_delayed_38__75_, chained_data_delayed_38__74_, chained_data_delayed_38__73_, chained_data_delayed_38__72_, chained_data_delayed_38__71_, chained_data_delayed_38__70_, chained_data_delayed_38__69_, chained_data_delayed_38__68_, chained_data_delayed_38__67_, chained_data_delayed_38__66_, chained_data_delayed_38__65_, chained_data_delayed_38__64_, chained_data_delayed_38__63_, chained_data_delayed_38__62_, chained_data_delayed_38__61_, chained_data_delayed_38__60_, chained_data_delayed_38__59_, chained_data_delayed_38__58_, chained_data_delayed_38__57_, chained_data_delayed_38__56_, chained_data_delayed_38__55_, chained_data_delayed_38__54_, chained_data_delayed_38__53_, chained_data_delayed_38__52_, chained_data_delayed_38__51_, chained_data_delayed_38__50_, chained_data_delayed_38__49_, chained_data_delayed_38__48_, chained_data_delayed_38__47_, chained_data_delayed_38__46_, chained_data_delayed_38__45_, chained_data_delayed_38__44_, chained_data_delayed_38__43_, chained_data_delayed_38__42_, chained_data_delayed_38__41_, chained_data_delayed_38__40_, chained_data_delayed_38__39_, chained_data_delayed_38__38_, chained_data_delayed_38__37_, chained_data_delayed_38__36_, chained_data_delayed_38__35_, chained_data_delayed_38__34_, chained_data_delayed_38__33_, chained_data_delayed_38__32_, chained_data_delayed_38__31_, chained_data_delayed_38__30_, chained_data_delayed_38__29_, chained_data_delayed_38__28_, chained_data_delayed_38__27_, chained_data_delayed_38__26_, chained_data_delayed_38__25_, chained_data_delayed_38__24_, chained_data_delayed_38__23_, chained_data_delayed_38__22_, chained_data_delayed_38__21_, chained_data_delayed_38__20_, chained_data_delayed_38__19_, chained_data_delayed_38__18_, chained_data_delayed_38__17_, chained_data_delayed_38__16_, chained_data_delayed_38__15_, chained_data_delayed_38__14_, chained_data_delayed_38__13_, chained_data_delayed_38__12_, chained_data_delayed_38__11_, chained_data_delayed_38__10_, chained_data_delayed_38__9_, chained_data_delayed_38__8_, chained_data_delayed_38__7_, chained_data_delayed_38__6_, chained_data_delayed_38__5_, chained_data_delayed_38__4_, chained_data_delayed_38__3_, chained_data_delayed_38__2_, chained_data_delayed_38__1_, chained_data_delayed_38__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_39__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_38__127_, chained_data_delayed_38__126_, chained_data_delayed_38__125_, chained_data_delayed_38__124_, chained_data_delayed_38__123_, chained_data_delayed_38__122_, chained_data_delayed_38__121_, chained_data_delayed_38__120_, chained_data_delayed_38__119_, chained_data_delayed_38__118_, chained_data_delayed_38__117_, chained_data_delayed_38__116_, chained_data_delayed_38__115_, chained_data_delayed_38__114_, chained_data_delayed_38__113_, chained_data_delayed_38__112_, chained_data_delayed_38__111_, chained_data_delayed_38__110_, chained_data_delayed_38__109_, chained_data_delayed_38__108_, chained_data_delayed_38__107_, chained_data_delayed_38__106_, chained_data_delayed_38__105_, chained_data_delayed_38__104_, chained_data_delayed_38__103_, chained_data_delayed_38__102_, chained_data_delayed_38__101_, chained_data_delayed_38__100_, chained_data_delayed_38__99_, chained_data_delayed_38__98_, chained_data_delayed_38__97_, chained_data_delayed_38__96_, chained_data_delayed_38__95_, chained_data_delayed_38__94_, chained_data_delayed_38__93_, chained_data_delayed_38__92_, chained_data_delayed_38__91_, chained_data_delayed_38__90_, chained_data_delayed_38__89_, chained_data_delayed_38__88_, chained_data_delayed_38__87_, chained_data_delayed_38__86_, chained_data_delayed_38__85_, chained_data_delayed_38__84_, chained_data_delayed_38__83_, chained_data_delayed_38__82_, chained_data_delayed_38__81_, chained_data_delayed_38__80_, chained_data_delayed_38__79_, chained_data_delayed_38__78_, chained_data_delayed_38__77_, chained_data_delayed_38__76_, chained_data_delayed_38__75_, chained_data_delayed_38__74_, chained_data_delayed_38__73_, chained_data_delayed_38__72_, chained_data_delayed_38__71_, chained_data_delayed_38__70_, chained_data_delayed_38__69_, chained_data_delayed_38__68_, chained_data_delayed_38__67_, chained_data_delayed_38__66_, chained_data_delayed_38__65_, chained_data_delayed_38__64_, chained_data_delayed_38__63_, chained_data_delayed_38__62_, chained_data_delayed_38__61_, chained_data_delayed_38__60_, chained_data_delayed_38__59_, chained_data_delayed_38__58_, chained_data_delayed_38__57_, chained_data_delayed_38__56_, chained_data_delayed_38__55_, chained_data_delayed_38__54_, chained_data_delayed_38__53_, chained_data_delayed_38__52_, chained_data_delayed_38__51_, chained_data_delayed_38__50_, chained_data_delayed_38__49_, chained_data_delayed_38__48_, chained_data_delayed_38__47_, chained_data_delayed_38__46_, chained_data_delayed_38__45_, chained_data_delayed_38__44_, chained_data_delayed_38__43_, chained_data_delayed_38__42_, chained_data_delayed_38__41_, chained_data_delayed_38__40_, chained_data_delayed_38__39_, chained_data_delayed_38__38_, chained_data_delayed_38__37_, chained_data_delayed_38__36_, chained_data_delayed_38__35_, chained_data_delayed_38__34_, chained_data_delayed_38__33_, chained_data_delayed_38__32_, chained_data_delayed_38__31_, chained_data_delayed_38__30_, chained_data_delayed_38__29_, chained_data_delayed_38__28_, chained_data_delayed_38__27_, chained_data_delayed_38__26_, chained_data_delayed_38__25_, chained_data_delayed_38__24_, chained_data_delayed_38__23_, chained_data_delayed_38__22_, chained_data_delayed_38__21_, chained_data_delayed_38__20_, chained_data_delayed_38__19_, chained_data_delayed_38__18_, chained_data_delayed_38__17_, chained_data_delayed_38__16_, chained_data_delayed_38__15_, chained_data_delayed_38__14_, chained_data_delayed_38__13_, chained_data_delayed_38__12_, chained_data_delayed_38__11_, chained_data_delayed_38__10_, chained_data_delayed_38__9_, chained_data_delayed_38__8_, chained_data_delayed_38__7_, chained_data_delayed_38__6_, chained_data_delayed_38__5_, chained_data_delayed_38__4_, chained_data_delayed_38__3_, chained_data_delayed_38__2_, chained_data_delayed_38__1_, chained_data_delayed_38__0_ }),
    .data_o({ chained_data_delayed_39__127_, chained_data_delayed_39__126_, chained_data_delayed_39__125_, chained_data_delayed_39__124_, chained_data_delayed_39__123_, chained_data_delayed_39__122_, chained_data_delayed_39__121_, chained_data_delayed_39__120_, chained_data_delayed_39__119_, chained_data_delayed_39__118_, chained_data_delayed_39__117_, chained_data_delayed_39__116_, chained_data_delayed_39__115_, chained_data_delayed_39__114_, chained_data_delayed_39__113_, chained_data_delayed_39__112_, chained_data_delayed_39__111_, chained_data_delayed_39__110_, chained_data_delayed_39__109_, chained_data_delayed_39__108_, chained_data_delayed_39__107_, chained_data_delayed_39__106_, chained_data_delayed_39__105_, chained_data_delayed_39__104_, chained_data_delayed_39__103_, chained_data_delayed_39__102_, chained_data_delayed_39__101_, chained_data_delayed_39__100_, chained_data_delayed_39__99_, chained_data_delayed_39__98_, chained_data_delayed_39__97_, chained_data_delayed_39__96_, chained_data_delayed_39__95_, chained_data_delayed_39__94_, chained_data_delayed_39__93_, chained_data_delayed_39__92_, chained_data_delayed_39__91_, chained_data_delayed_39__90_, chained_data_delayed_39__89_, chained_data_delayed_39__88_, chained_data_delayed_39__87_, chained_data_delayed_39__86_, chained_data_delayed_39__85_, chained_data_delayed_39__84_, chained_data_delayed_39__83_, chained_data_delayed_39__82_, chained_data_delayed_39__81_, chained_data_delayed_39__80_, chained_data_delayed_39__79_, chained_data_delayed_39__78_, chained_data_delayed_39__77_, chained_data_delayed_39__76_, chained_data_delayed_39__75_, chained_data_delayed_39__74_, chained_data_delayed_39__73_, chained_data_delayed_39__72_, chained_data_delayed_39__71_, chained_data_delayed_39__70_, chained_data_delayed_39__69_, chained_data_delayed_39__68_, chained_data_delayed_39__67_, chained_data_delayed_39__66_, chained_data_delayed_39__65_, chained_data_delayed_39__64_, chained_data_delayed_39__63_, chained_data_delayed_39__62_, chained_data_delayed_39__61_, chained_data_delayed_39__60_, chained_data_delayed_39__59_, chained_data_delayed_39__58_, chained_data_delayed_39__57_, chained_data_delayed_39__56_, chained_data_delayed_39__55_, chained_data_delayed_39__54_, chained_data_delayed_39__53_, chained_data_delayed_39__52_, chained_data_delayed_39__51_, chained_data_delayed_39__50_, chained_data_delayed_39__49_, chained_data_delayed_39__48_, chained_data_delayed_39__47_, chained_data_delayed_39__46_, chained_data_delayed_39__45_, chained_data_delayed_39__44_, chained_data_delayed_39__43_, chained_data_delayed_39__42_, chained_data_delayed_39__41_, chained_data_delayed_39__40_, chained_data_delayed_39__39_, chained_data_delayed_39__38_, chained_data_delayed_39__37_, chained_data_delayed_39__36_, chained_data_delayed_39__35_, chained_data_delayed_39__34_, chained_data_delayed_39__33_, chained_data_delayed_39__32_, chained_data_delayed_39__31_, chained_data_delayed_39__30_, chained_data_delayed_39__29_, chained_data_delayed_39__28_, chained_data_delayed_39__27_, chained_data_delayed_39__26_, chained_data_delayed_39__25_, chained_data_delayed_39__24_, chained_data_delayed_39__23_, chained_data_delayed_39__22_, chained_data_delayed_39__21_, chained_data_delayed_39__20_, chained_data_delayed_39__19_, chained_data_delayed_39__18_, chained_data_delayed_39__17_, chained_data_delayed_39__16_, chained_data_delayed_39__15_, chained_data_delayed_39__14_, chained_data_delayed_39__13_, chained_data_delayed_39__12_, chained_data_delayed_39__11_, chained_data_delayed_39__10_, chained_data_delayed_39__9_, chained_data_delayed_39__8_, chained_data_delayed_39__7_, chained_data_delayed_39__6_, chained_data_delayed_39__5_, chained_data_delayed_39__4_, chained_data_delayed_39__3_, chained_data_delayed_39__2_, chained_data_delayed_39__1_, chained_data_delayed_39__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_40__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_39__127_, chained_data_delayed_39__126_, chained_data_delayed_39__125_, chained_data_delayed_39__124_, chained_data_delayed_39__123_, chained_data_delayed_39__122_, chained_data_delayed_39__121_, chained_data_delayed_39__120_, chained_data_delayed_39__119_, chained_data_delayed_39__118_, chained_data_delayed_39__117_, chained_data_delayed_39__116_, chained_data_delayed_39__115_, chained_data_delayed_39__114_, chained_data_delayed_39__113_, chained_data_delayed_39__112_, chained_data_delayed_39__111_, chained_data_delayed_39__110_, chained_data_delayed_39__109_, chained_data_delayed_39__108_, chained_data_delayed_39__107_, chained_data_delayed_39__106_, chained_data_delayed_39__105_, chained_data_delayed_39__104_, chained_data_delayed_39__103_, chained_data_delayed_39__102_, chained_data_delayed_39__101_, chained_data_delayed_39__100_, chained_data_delayed_39__99_, chained_data_delayed_39__98_, chained_data_delayed_39__97_, chained_data_delayed_39__96_, chained_data_delayed_39__95_, chained_data_delayed_39__94_, chained_data_delayed_39__93_, chained_data_delayed_39__92_, chained_data_delayed_39__91_, chained_data_delayed_39__90_, chained_data_delayed_39__89_, chained_data_delayed_39__88_, chained_data_delayed_39__87_, chained_data_delayed_39__86_, chained_data_delayed_39__85_, chained_data_delayed_39__84_, chained_data_delayed_39__83_, chained_data_delayed_39__82_, chained_data_delayed_39__81_, chained_data_delayed_39__80_, chained_data_delayed_39__79_, chained_data_delayed_39__78_, chained_data_delayed_39__77_, chained_data_delayed_39__76_, chained_data_delayed_39__75_, chained_data_delayed_39__74_, chained_data_delayed_39__73_, chained_data_delayed_39__72_, chained_data_delayed_39__71_, chained_data_delayed_39__70_, chained_data_delayed_39__69_, chained_data_delayed_39__68_, chained_data_delayed_39__67_, chained_data_delayed_39__66_, chained_data_delayed_39__65_, chained_data_delayed_39__64_, chained_data_delayed_39__63_, chained_data_delayed_39__62_, chained_data_delayed_39__61_, chained_data_delayed_39__60_, chained_data_delayed_39__59_, chained_data_delayed_39__58_, chained_data_delayed_39__57_, chained_data_delayed_39__56_, chained_data_delayed_39__55_, chained_data_delayed_39__54_, chained_data_delayed_39__53_, chained_data_delayed_39__52_, chained_data_delayed_39__51_, chained_data_delayed_39__50_, chained_data_delayed_39__49_, chained_data_delayed_39__48_, chained_data_delayed_39__47_, chained_data_delayed_39__46_, chained_data_delayed_39__45_, chained_data_delayed_39__44_, chained_data_delayed_39__43_, chained_data_delayed_39__42_, chained_data_delayed_39__41_, chained_data_delayed_39__40_, chained_data_delayed_39__39_, chained_data_delayed_39__38_, chained_data_delayed_39__37_, chained_data_delayed_39__36_, chained_data_delayed_39__35_, chained_data_delayed_39__34_, chained_data_delayed_39__33_, chained_data_delayed_39__32_, chained_data_delayed_39__31_, chained_data_delayed_39__30_, chained_data_delayed_39__29_, chained_data_delayed_39__28_, chained_data_delayed_39__27_, chained_data_delayed_39__26_, chained_data_delayed_39__25_, chained_data_delayed_39__24_, chained_data_delayed_39__23_, chained_data_delayed_39__22_, chained_data_delayed_39__21_, chained_data_delayed_39__20_, chained_data_delayed_39__19_, chained_data_delayed_39__18_, chained_data_delayed_39__17_, chained_data_delayed_39__16_, chained_data_delayed_39__15_, chained_data_delayed_39__14_, chained_data_delayed_39__13_, chained_data_delayed_39__12_, chained_data_delayed_39__11_, chained_data_delayed_39__10_, chained_data_delayed_39__9_, chained_data_delayed_39__8_, chained_data_delayed_39__7_, chained_data_delayed_39__6_, chained_data_delayed_39__5_, chained_data_delayed_39__4_, chained_data_delayed_39__3_, chained_data_delayed_39__2_, chained_data_delayed_39__1_, chained_data_delayed_39__0_ }),
    .data_o({ chained_data_delayed_40__127_, chained_data_delayed_40__126_, chained_data_delayed_40__125_, chained_data_delayed_40__124_, chained_data_delayed_40__123_, chained_data_delayed_40__122_, chained_data_delayed_40__121_, chained_data_delayed_40__120_, chained_data_delayed_40__119_, chained_data_delayed_40__118_, chained_data_delayed_40__117_, chained_data_delayed_40__116_, chained_data_delayed_40__115_, chained_data_delayed_40__114_, chained_data_delayed_40__113_, chained_data_delayed_40__112_, chained_data_delayed_40__111_, chained_data_delayed_40__110_, chained_data_delayed_40__109_, chained_data_delayed_40__108_, chained_data_delayed_40__107_, chained_data_delayed_40__106_, chained_data_delayed_40__105_, chained_data_delayed_40__104_, chained_data_delayed_40__103_, chained_data_delayed_40__102_, chained_data_delayed_40__101_, chained_data_delayed_40__100_, chained_data_delayed_40__99_, chained_data_delayed_40__98_, chained_data_delayed_40__97_, chained_data_delayed_40__96_, chained_data_delayed_40__95_, chained_data_delayed_40__94_, chained_data_delayed_40__93_, chained_data_delayed_40__92_, chained_data_delayed_40__91_, chained_data_delayed_40__90_, chained_data_delayed_40__89_, chained_data_delayed_40__88_, chained_data_delayed_40__87_, chained_data_delayed_40__86_, chained_data_delayed_40__85_, chained_data_delayed_40__84_, chained_data_delayed_40__83_, chained_data_delayed_40__82_, chained_data_delayed_40__81_, chained_data_delayed_40__80_, chained_data_delayed_40__79_, chained_data_delayed_40__78_, chained_data_delayed_40__77_, chained_data_delayed_40__76_, chained_data_delayed_40__75_, chained_data_delayed_40__74_, chained_data_delayed_40__73_, chained_data_delayed_40__72_, chained_data_delayed_40__71_, chained_data_delayed_40__70_, chained_data_delayed_40__69_, chained_data_delayed_40__68_, chained_data_delayed_40__67_, chained_data_delayed_40__66_, chained_data_delayed_40__65_, chained_data_delayed_40__64_, chained_data_delayed_40__63_, chained_data_delayed_40__62_, chained_data_delayed_40__61_, chained_data_delayed_40__60_, chained_data_delayed_40__59_, chained_data_delayed_40__58_, chained_data_delayed_40__57_, chained_data_delayed_40__56_, chained_data_delayed_40__55_, chained_data_delayed_40__54_, chained_data_delayed_40__53_, chained_data_delayed_40__52_, chained_data_delayed_40__51_, chained_data_delayed_40__50_, chained_data_delayed_40__49_, chained_data_delayed_40__48_, chained_data_delayed_40__47_, chained_data_delayed_40__46_, chained_data_delayed_40__45_, chained_data_delayed_40__44_, chained_data_delayed_40__43_, chained_data_delayed_40__42_, chained_data_delayed_40__41_, chained_data_delayed_40__40_, chained_data_delayed_40__39_, chained_data_delayed_40__38_, chained_data_delayed_40__37_, chained_data_delayed_40__36_, chained_data_delayed_40__35_, chained_data_delayed_40__34_, chained_data_delayed_40__33_, chained_data_delayed_40__32_, chained_data_delayed_40__31_, chained_data_delayed_40__30_, chained_data_delayed_40__29_, chained_data_delayed_40__28_, chained_data_delayed_40__27_, chained_data_delayed_40__26_, chained_data_delayed_40__25_, chained_data_delayed_40__24_, chained_data_delayed_40__23_, chained_data_delayed_40__22_, chained_data_delayed_40__21_, chained_data_delayed_40__20_, chained_data_delayed_40__19_, chained_data_delayed_40__18_, chained_data_delayed_40__17_, chained_data_delayed_40__16_, chained_data_delayed_40__15_, chained_data_delayed_40__14_, chained_data_delayed_40__13_, chained_data_delayed_40__12_, chained_data_delayed_40__11_, chained_data_delayed_40__10_, chained_data_delayed_40__9_, chained_data_delayed_40__8_, chained_data_delayed_40__7_, chained_data_delayed_40__6_, chained_data_delayed_40__5_, chained_data_delayed_40__4_, chained_data_delayed_40__3_, chained_data_delayed_40__2_, chained_data_delayed_40__1_, chained_data_delayed_40__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_41__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_40__127_, chained_data_delayed_40__126_, chained_data_delayed_40__125_, chained_data_delayed_40__124_, chained_data_delayed_40__123_, chained_data_delayed_40__122_, chained_data_delayed_40__121_, chained_data_delayed_40__120_, chained_data_delayed_40__119_, chained_data_delayed_40__118_, chained_data_delayed_40__117_, chained_data_delayed_40__116_, chained_data_delayed_40__115_, chained_data_delayed_40__114_, chained_data_delayed_40__113_, chained_data_delayed_40__112_, chained_data_delayed_40__111_, chained_data_delayed_40__110_, chained_data_delayed_40__109_, chained_data_delayed_40__108_, chained_data_delayed_40__107_, chained_data_delayed_40__106_, chained_data_delayed_40__105_, chained_data_delayed_40__104_, chained_data_delayed_40__103_, chained_data_delayed_40__102_, chained_data_delayed_40__101_, chained_data_delayed_40__100_, chained_data_delayed_40__99_, chained_data_delayed_40__98_, chained_data_delayed_40__97_, chained_data_delayed_40__96_, chained_data_delayed_40__95_, chained_data_delayed_40__94_, chained_data_delayed_40__93_, chained_data_delayed_40__92_, chained_data_delayed_40__91_, chained_data_delayed_40__90_, chained_data_delayed_40__89_, chained_data_delayed_40__88_, chained_data_delayed_40__87_, chained_data_delayed_40__86_, chained_data_delayed_40__85_, chained_data_delayed_40__84_, chained_data_delayed_40__83_, chained_data_delayed_40__82_, chained_data_delayed_40__81_, chained_data_delayed_40__80_, chained_data_delayed_40__79_, chained_data_delayed_40__78_, chained_data_delayed_40__77_, chained_data_delayed_40__76_, chained_data_delayed_40__75_, chained_data_delayed_40__74_, chained_data_delayed_40__73_, chained_data_delayed_40__72_, chained_data_delayed_40__71_, chained_data_delayed_40__70_, chained_data_delayed_40__69_, chained_data_delayed_40__68_, chained_data_delayed_40__67_, chained_data_delayed_40__66_, chained_data_delayed_40__65_, chained_data_delayed_40__64_, chained_data_delayed_40__63_, chained_data_delayed_40__62_, chained_data_delayed_40__61_, chained_data_delayed_40__60_, chained_data_delayed_40__59_, chained_data_delayed_40__58_, chained_data_delayed_40__57_, chained_data_delayed_40__56_, chained_data_delayed_40__55_, chained_data_delayed_40__54_, chained_data_delayed_40__53_, chained_data_delayed_40__52_, chained_data_delayed_40__51_, chained_data_delayed_40__50_, chained_data_delayed_40__49_, chained_data_delayed_40__48_, chained_data_delayed_40__47_, chained_data_delayed_40__46_, chained_data_delayed_40__45_, chained_data_delayed_40__44_, chained_data_delayed_40__43_, chained_data_delayed_40__42_, chained_data_delayed_40__41_, chained_data_delayed_40__40_, chained_data_delayed_40__39_, chained_data_delayed_40__38_, chained_data_delayed_40__37_, chained_data_delayed_40__36_, chained_data_delayed_40__35_, chained_data_delayed_40__34_, chained_data_delayed_40__33_, chained_data_delayed_40__32_, chained_data_delayed_40__31_, chained_data_delayed_40__30_, chained_data_delayed_40__29_, chained_data_delayed_40__28_, chained_data_delayed_40__27_, chained_data_delayed_40__26_, chained_data_delayed_40__25_, chained_data_delayed_40__24_, chained_data_delayed_40__23_, chained_data_delayed_40__22_, chained_data_delayed_40__21_, chained_data_delayed_40__20_, chained_data_delayed_40__19_, chained_data_delayed_40__18_, chained_data_delayed_40__17_, chained_data_delayed_40__16_, chained_data_delayed_40__15_, chained_data_delayed_40__14_, chained_data_delayed_40__13_, chained_data_delayed_40__12_, chained_data_delayed_40__11_, chained_data_delayed_40__10_, chained_data_delayed_40__9_, chained_data_delayed_40__8_, chained_data_delayed_40__7_, chained_data_delayed_40__6_, chained_data_delayed_40__5_, chained_data_delayed_40__4_, chained_data_delayed_40__3_, chained_data_delayed_40__2_, chained_data_delayed_40__1_, chained_data_delayed_40__0_ }),
    .data_o({ chained_data_delayed_41__127_, chained_data_delayed_41__126_, chained_data_delayed_41__125_, chained_data_delayed_41__124_, chained_data_delayed_41__123_, chained_data_delayed_41__122_, chained_data_delayed_41__121_, chained_data_delayed_41__120_, chained_data_delayed_41__119_, chained_data_delayed_41__118_, chained_data_delayed_41__117_, chained_data_delayed_41__116_, chained_data_delayed_41__115_, chained_data_delayed_41__114_, chained_data_delayed_41__113_, chained_data_delayed_41__112_, chained_data_delayed_41__111_, chained_data_delayed_41__110_, chained_data_delayed_41__109_, chained_data_delayed_41__108_, chained_data_delayed_41__107_, chained_data_delayed_41__106_, chained_data_delayed_41__105_, chained_data_delayed_41__104_, chained_data_delayed_41__103_, chained_data_delayed_41__102_, chained_data_delayed_41__101_, chained_data_delayed_41__100_, chained_data_delayed_41__99_, chained_data_delayed_41__98_, chained_data_delayed_41__97_, chained_data_delayed_41__96_, chained_data_delayed_41__95_, chained_data_delayed_41__94_, chained_data_delayed_41__93_, chained_data_delayed_41__92_, chained_data_delayed_41__91_, chained_data_delayed_41__90_, chained_data_delayed_41__89_, chained_data_delayed_41__88_, chained_data_delayed_41__87_, chained_data_delayed_41__86_, chained_data_delayed_41__85_, chained_data_delayed_41__84_, chained_data_delayed_41__83_, chained_data_delayed_41__82_, chained_data_delayed_41__81_, chained_data_delayed_41__80_, chained_data_delayed_41__79_, chained_data_delayed_41__78_, chained_data_delayed_41__77_, chained_data_delayed_41__76_, chained_data_delayed_41__75_, chained_data_delayed_41__74_, chained_data_delayed_41__73_, chained_data_delayed_41__72_, chained_data_delayed_41__71_, chained_data_delayed_41__70_, chained_data_delayed_41__69_, chained_data_delayed_41__68_, chained_data_delayed_41__67_, chained_data_delayed_41__66_, chained_data_delayed_41__65_, chained_data_delayed_41__64_, chained_data_delayed_41__63_, chained_data_delayed_41__62_, chained_data_delayed_41__61_, chained_data_delayed_41__60_, chained_data_delayed_41__59_, chained_data_delayed_41__58_, chained_data_delayed_41__57_, chained_data_delayed_41__56_, chained_data_delayed_41__55_, chained_data_delayed_41__54_, chained_data_delayed_41__53_, chained_data_delayed_41__52_, chained_data_delayed_41__51_, chained_data_delayed_41__50_, chained_data_delayed_41__49_, chained_data_delayed_41__48_, chained_data_delayed_41__47_, chained_data_delayed_41__46_, chained_data_delayed_41__45_, chained_data_delayed_41__44_, chained_data_delayed_41__43_, chained_data_delayed_41__42_, chained_data_delayed_41__41_, chained_data_delayed_41__40_, chained_data_delayed_41__39_, chained_data_delayed_41__38_, chained_data_delayed_41__37_, chained_data_delayed_41__36_, chained_data_delayed_41__35_, chained_data_delayed_41__34_, chained_data_delayed_41__33_, chained_data_delayed_41__32_, chained_data_delayed_41__31_, chained_data_delayed_41__30_, chained_data_delayed_41__29_, chained_data_delayed_41__28_, chained_data_delayed_41__27_, chained_data_delayed_41__26_, chained_data_delayed_41__25_, chained_data_delayed_41__24_, chained_data_delayed_41__23_, chained_data_delayed_41__22_, chained_data_delayed_41__21_, chained_data_delayed_41__20_, chained_data_delayed_41__19_, chained_data_delayed_41__18_, chained_data_delayed_41__17_, chained_data_delayed_41__16_, chained_data_delayed_41__15_, chained_data_delayed_41__14_, chained_data_delayed_41__13_, chained_data_delayed_41__12_, chained_data_delayed_41__11_, chained_data_delayed_41__10_, chained_data_delayed_41__9_, chained_data_delayed_41__8_, chained_data_delayed_41__7_, chained_data_delayed_41__6_, chained_data_delayed_41__5_, chained_data_delayed_41__4_, chained_data_delayed_41__3_, chained_data_delayed_41__2_, chained_data_delayed_41__1_, chained_data_delayed_41__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_42__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_41__127_, chained_data_delayed_41__126_, chained_data_delayed_41__125_, chained_data_delayed_41__124_, chained_data_delayed_41__123_, chained_data_delayed_41__122_, chained_data_delayed_41__121_, chained_data_delayed_41__120_, chained_data_delayed_41__119_, chained_data_delayed_41__118_, chained_data_delayed_41__117_, chained_data_delayed_41__116_, chained_data_delayed_41__115_, chained_data_delayed_41__114_, chained_data_delayed_41__113_, chained_data_delayed_41__112_, chained_data_delayed_41__111_, chained_data_delayed_41__110_, chained_data_delayed_41__109_, chained_data_delayed_41__108_, chained_data_delayed_41__107_, chained_data_delayed_41__106_, chained_data_delayed_41__105_, chained_data_delayed_41__104_, chained_data_delayed_41__103_, chained_data_delayed_41__102_, chained_data_delayed_41__101_, chained_data_delayed_41__100_, chained_data_delayed_41__99_, chained_data_delayed_41__98_, chained_data_delayed_41__97_, chained_data_delayed_41__96_, chained_data_delayed_41__95_, chained_data_delayed_41__94_, chained_data_delayed_41__93_, chained_data_delayed_41__92_, chained_data_delayed_41__91_, chained_data_delayed_41__90_, chained_data_delayed_41__89_, chained_data_delayed_41__88_, chained_data_delayed_41__87_, chained_data_delayed_41__86_, chained_data_delayed_41__85_, chained_data_delayed_41__84_, chained_data_delayed_41__83_, chained_data_delayed_41__82_, chained_data_delayed_41__81_, chained_data_delayed_41__80_, chained_data_delayed_41__79_, chained_data_delayed_41__78_, chained_data_delayed_41__77_, chained_data_delayed_41__76_, chained_data_delayed_41__75_, chained_data_delayed_41__74_, chained_data_delayed_41__73_, chained_data_delayed_41__72_, chained_data_delayed_41__71_, chained_data_delayed_41__70_, chained_data_delayed_41__69_, chained_data_delayed_41__68_, chained_data_delayed_41__67_, chained_data_delayed_41__66_, chained_data_delayed_41__65_, chained_data_delayed_41__64_, chained_data_delayed_41__63_, chained_data_delayed_41__62_, chained_data_delayed_41__61_, chained_data_delayed_41__60_, chained_data_delayed_41__59_, chained_data_delayed_41__58_, chained_data_delayed_41__57_, chained_data_delayed_41__56_, chained_data_delayed_41__55_, chained_data_delayed_41__54_, chained_data_delayed_41__53_, chained_data_delayed_41__52_, chained_data_delayed_41__51_, chained_data_delayed_41__50_, chained_data_delayed_41__49_, chained_data_delayed_41__48_, chained_data_delayed_41__47_, chained_data_delayed_41__46_, chained_data_delayed_41__45_, chained_data_delayed_41__44_, chained_data_delayed_41__43_, chained_data_delayed_41__42_, chained_data_delayed_41__41_, chained_data_delayed_41__40_, chained_data_delayed_41__39_, chained_data_delayed_41__38_, chained_data_delayed_41__37_, chained_data_delayed_41__36_, chained_data_delayed_41__35_, chained_data_delayed_41__34_, chained_data_delayed_41__33_, chained_data_delayed_41__32_, chained_data_delayed_41__31_, chained_data_delayed_41__30_, chained_data_delayed_41__29_, chained_data_delayed_41__28_, chained_data_delayed_41__27_, chained_data_delayed_41__26_, chained_data_delayed_41__25_, chained_data_delayed_41__24_, chained_data_delayed_41__23_, chained_data_delayed_41__22_, chained_data_delayed_41__21_, chained_data_delayed_41__20_, chained_data_delayed_41__19_, chained_data_delayed_41__18_, chained_data_delayed_41__17_, chained_data_delayed_41__16_, chained_data_delayed_41__15_, chained_data_delayed_41__14_, chained_data_delayed_41__13_, chained_data_delayed_41__12_, chained_data_delayed_41__11_, chained_data_delayed_41__10_, chained_data_delayed_41__9_, chained_data_delayed_41__8_, chained_data_delayed_41__7_, chained_data_delayed_41__6_, chained_data_delayed_41__5_, chained_data_delayed_41__4_, chained_data_delayed_41__3_, chained_data_delayed_41__2_, chained_data_delayed_41__1_, chained_data_delayed_41__0_ }),
    .data_o({ chained_data_delayed_42__127_, chained_data_delayed_42__126_, chained_data_delayed_42__125_, chained_data_delayed_42__124_, chained_data_delayed_42__123_, chained_data_delayed_42__122_, chained_data_delayed_42__121_, chained_data_delayed_42__120_, chained_data_delayed_42__119_, chained_data_delayed_42__118_, chained_data_delayed_42__117_, chained_data_delayed_42__116_, chained_data_delayed_42__115_, chained_data_delayed_42__114_, chained_data_delayed_42__113_, chained_data_delayed_42__112_, chained_data_delayed_42__111_, chained_data_delayed_42__110_, chained_data_delayed_42__109_, chained_data_delayed_42__108_, chained_data_delayed_42__107_, chained_data_delayed_42__106_, chained_data_delayed_42__105_, chained_data_delayed_42__104_, chained_data_delayed_42__103_, chained_data_delayed_42__102_, chained_data_delayed_42__101_, chained_data_delayed_42__100_, chained_data_delayed_42__99_, chained_data_delayed_42__98_, chained_data_delayed_42__97_, chained_data_delayed_42__96_, chained_data_delayed_42__95_, chained_data_delayed_42__94_, chained_data_delayed_42__93_, chained_data_delayed_42__92_, chained_data_delayed_42__91_, chained_data_delayed_42__90_, chained_data_delayed_42__89_, chained_data_delayed_42__88_, chained_data_delayed_42__87_, chained_data_delayed_42__86_, chained_data_delayed_42__85_, chained_data_delayed_42__84_, chained_data_delayed_42__83_, chained_data_delayed_42__82_, chained_data_delayed_42__81_, chained_data_delayed_42__80_, chained_data_delayed_42__79_, chained_data_delayed_42__78_, chained_data_delayed_42__77_, chained_data_delayed_42__76_, chained_data_delayed_42__75_, chained_data_delayed_42__74_, chained_data_delayed_42__73_, chained_data_delayed_42__72_, chained_data_delayed_42__71_, chained_data_delayed_42__70_, chained_data_delayed_42__69_, chained_data_delayed_42__68_, chained_data_delayed_42__67_, chained_data_delayed_42__66_, chained_data_delayed_42__65_, chained_data_delayed_42__64_, chained_data_delayed_42__63_, chained_data_delayed_42__62_, chained_data_delayed_42__61_, chained_data_delayed_42__60_, chained_data_delayed_42__59_, chained_data_delayed_42__58_, chained_data_delayed_42__57_, chained_data_delayed_42__56_, chained_data_delayed_42__55_, chained_data_delayed_42__54_, chained_data_delayed_42__53_, chained_data_delayed_42__52_, chained_data_delayed_42__51_, chained_data_delayed_42__50_, chained_data_delayed_42__49_, chained_data_delayed_42__48_, chained_data_delayed_42__47_, chained_data_delayed_42__46_, chained_data_delayed_42__45_, chained_data_delayed_42__44_, chained_data_delayed_42__43_, chained_data_delayed_42__42_, chained_data_delayed_42__41_, chained_data_delayed_42__40_, chained_data_delayed_42__39_, chained_data_delayed_42__38_, chained_data_delayed_42__37_, chained_data_delayed_42__36_, chained_data_delayed_42__35_, chained_data_delayed_42__34_, chained_data_delayed_42__33_, chained_data_delayed_42__32_, chained_data_delayed_42__31_, chained_data_delayed_42__30_, chained_data_delayed_42__29_, chained_data_delayed_42__28_, chained_data_delayed_42__27_, chained_data_delayed_42__26_, chained_data_delayed_42__25_, chained_data_delayed_42__24_, chained_data_delayed_42__23_, chained_data_delayed_42__22_, chained_data_delayed_42__21_, chained_data_delayed_42__20_, chained_data_delayed_42__19_, chained_data_delayed_42__18_, chained_data_delayed_42__17_, chained_data_delayed_42__16_, chained_data_delayed_42__15_, chained_data_delayed_42__14_, chained_data_delayed_42__13_, chained_data_delayed_42__12_, chained_data_delayed_42__11_, chained_data_delayed_42__10_, chained_data_delayed_42__9_, chained_data_delayed_42__8_, chained_data_delayed_42__7_, chained_data_delayed_42__6_, chained_data_delayed_42__5_, chained_data_delayed_42__4_, chained_data_delayed_42__3_, chained_data_delayed_42__2_, chained_data_delayed_42__1_, chained_data_delayed_42__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_43__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_42__127_, chained_data_delayed_42__126_, chained_data_delayed_42__125_, chained_data_delayed_42__124_, chained_data_delayed_42__123_, chained_data_delayed_42__122_, chained_data_delayed_42__121_, chained_data_delayed_42__120_, chained_data_delayed_42__119_, chained_data_delayed_42__118_, chained_data_delayed_42__117_, chained_data_delayed_42__116_, chained_data_delayed_42__115_, chained_data_delayed_42__114_, chained_data_delayed_42__113_, chained_data_delayed_42__112_, chained_data_delayed_42__111_, chained_data_delayed_42__110_, chained_data_delayed_42__109_, chained_data_delayed_42__108_, chained_data_delayed_42__107_, chained_data_delayed_42__106_, chained_data_delayed_42__105_, chained_data_delayed_42__104_, chained_data_delayed_42__103_, chained_data_delayed_42__102_, chained_data_delayed_42__101_, chained_data_delayed_42__100_, chained_data_delayed_42__99_, chained_data_delayed_42__98_, chained_data_delayed_42__97_, chained_data_delayed_42__96_, chained_data_delayed_42__95_, chained_data_delayed_42__94_, chained_data_delayed_42__93_, chained_data_delayed_42__92_, chained_data_delayed_42__91_, chained_data_delayed_42__90_, chained_data_delayed_42__89_, chained_data_delayed_42__88_, chained_data_delayed_42__87_, chained_data_delayed_42__86_, chained_data_delayed_42__85_, chained_data_delayed_42__84_, chained_data_delayed_42__83_, chained_data_delayed_42__82_, chained_data_delayed_42__81_, chained_data_delayed_42__80_, chained_data_delayed_42__79_, chained_data_delayed_42__78_, chained_data_delayed_42__77_, chained_data_delayed_42__76_, chained_data_delayed_42__75_, chained_data_delayed_42__74_, chained_data_delayed_42__73_, chained_data_delayed_42__72_, chained_data_delayed_42__71_, chained_data_delayed_42__70_, chained_data_delayed_42__69_, chained_data_delayed_42__68_, chained_data_delayed_42__67_, chained_data_delayed_42__66_, chained_data_delayed_42__65_, chained_data_delayed_42__64_, chained_data_delayed_42__63_, chained_data_delayed_42__62_, chained_data_delayed_42__61_, chained_data_delayed_42__60_, chained_data_delayed_42__59_, chained_data_delayed_42__58_, chained_data_delayed_42__57_, chained_data_delayed_42__56_, chained_data_delayed_42__55_, chained_data_delayed_42__54_, chained_data_delayed_42__53_, chained_data_delayed_42__52_, chained_data_delayed_42__51_, chained_data_delayed_42__50_, chained_data_delayed_42__49_, chained_data_delayed_42__48_, chained_data_delayed_42__47_, chained_data_delayed_42__46_, chained_data_delayed_42__45_, chained_data_delayed_42__44_, chained_data_delayed_42__43_, chained_data_delayed_42__42_, chained_data_delayed_42__41_, chained_data_delayed_42__40_, chained_data_delayed_42__39_, chained_data_delayed_42__38_, chained_data_delayed_42__37_, chained_data_delayed_42__36_, chained_data_delayed_42__35_, chained_data_delayed_42__34_, chained_data_delayed_42__33_, chained_data_delayed_42__32_, chained_data_delayed_42__31_, chained_data_delayed_42__30_, chained_data_delayed_42__29_, chained_data_delayed_42__28_, chained_data_delayed_42__27_, chained_data_delayed_42__26_, chained_data_delayed_42__25_, chained_data_delayed_42__24_, chained_data_delayed_42__23_, chained_data_delayed_42__22_, chained_data_delayed_42__21_, chained_data_delayed_42__20_, chained_data_delayed_42__19_, chained_data_delayed_42__18_, chained_data_delayed_42__17_, chained_data_delayed_42__16_, chained_data_delayed_42__15_, chained_data_delayed_42__14_, chained_data_delayed_42__13_, chained_data_delayed_42__12_, chained_data_delayed_42__11_, chained_data_delayed_42__10_, chained_data_delayed_42__9_, chained_data_delayed_42__8_, chained_data_delayed_42__7_, chained_data_delayed_42__6_, chained_data_delayed_42__5_, chained_data_delayed_42__4_, chained_data_delayed_42__3_, chained_data_delayed_42__2_, chained_data_delayed_42__1_, chained_data_delayed_42__0_ }),
    .data_o({ chained_data_delayed_43__127_, chained_data_delayed_43__126_, chained_data_delayed_43__125_, chained_data_delayed_43__124_, chained_data_delayed_43__123_, chained_data_delayed_43__122_, chained_data_delayed_43__121_, chained_data_delayed_43__120_, chained_data_delayed_43__119_, chained_data_delayed_43__118_, chained_data_delayed_43__117_, chained_data_delayed_43__116_, chained_data_delayed_43__115_, chained_data_delayed_43__114_, chained_data_delayed_43__113_, chained_data_delayed_43__112_, chained_data_delayed_43__111_, chained_data_delayed_43__110_, chained_data_delayed_43__109_, chained_data_delayed_43__108_, chained_data_delayed_43__107_, chained_data_delayed_43__106_, chained_data_delayed_43__105_, chained_data_delayed_43__104_, chained_data_delayed_43__103_, chained_data_delayed_43__102_, chained_data_delayed_43__101_, chained_data_delayed_43__100_, chained_data_delayed_43__99_, chained_data_delayed_43__98_, chained_data_delayed_43__97_, chained_data_delayed_43__96_, chained_data_delayed_43__95_, chained_data_delayed_43__94_, chained_data_delayed_43__93_, chained_data_delayed_43__92_, chained_data_delayed_43__91_, chained_data_delayed_43__90_, chained_data_delayed_43__89_, chained_data_delayed_43__88_, chained_data_delayed_43__87_, chained_data_delayed_43__86_, chained_data_delayed_43__85_, chained_data_delayed_43__84_, chained_data_delayed_43__83_, chained_data_delayed_43__82_, chained_data_delayed_43__81_, chained_data_delayed_43__80_, chained_data_delayed_43__79_, chained_data_delayed_43__78_, chained_data_delayed_43__77_, chained_data_delayed_43__76_, chained_data_delayed_43__75_, chained_data_delayed_43__74_, chained_data_delayed_43__73_, chained_data_delayed_43__72_, chained_data_delayed_43__71_, chained_data_delayed_43__70_, chained_data_delayed_43__69_, chained_data_delayed_43__68_, chained_data_delayed_43__67_, chained_data_delayed_43__66_, chained_data_delayed_43__65_, chained_data_delayed_43__64_, chained_data_delayed_43__63_, chained_data_delayed_43__62_, chained_data_delayed_43__61_, chained_data_delayed_43__60_, chained_data_delayed_43__59_, chained_data_delayed_43__58_, chained_data_delayed_43__57_, chained_data_delayed_43__56_, chained_data_delayed_43__55_, chained_data_delayed_43__54_, chained_data_delayed_43__53_, chained_data_delayed_43__52_, chained_data_delayed_43__51_, chained_data_delayed_43__50_, chained_data_delayed_43__49_, chained_data_delayed_43__48_, chained_data_delayed_43__47_, chained_data_delayed_43__46_, chained_data_delayed_43__45_, chained_data_delayed_43__44_, chained_data_delayed_43__43_, chained_data_delayed_43__42_, chained_data_delayed_43__41_, chained_data_delayed_43__40_, chained_data_delayed_43__39_, chained_data_delayed_43__38_, chained_data_delayed_43__37_, chained_data_delayed_43__36_, chained_data_delayed_43__35_, chained_data_delayed_43__34_, chained_data_delayed_43__33_, chained_data_delayed_43__32_, chained_data_delayed_43__31_, chained_data_delayed_43__30_, chained_data_delayed_43__29_, chained_data_delayed_43__28_, chained_data_delayed_43__27_, chained_data_delayed_43__26_, chained_data_delayed_43__25_, chained_data_delayed_43__24_, chained_data_delayed_43__23_, chained_data_delayed_43__22_, chained_data_delayed_43__21_, chained_data_delayed_43__20_, chained_data_delayed_43__19_, chained_data_delayed_43__18_, chained_data_delayed_43__17_, chained_data_delayed_43__16_, chained_data_delayed_43__15_, chained_data_delayed_43__14_, chained_data_delayed_43__13_, chained_data_delayed_43__12_, chained_data_delayed_43__11_, chained_data_delayed_43__10_, chained_data_delayed_43__9_, chained_data_delayed_43__8_, chained_data_delayed_43__7_, chained_data_delayed_43__6_, chained_data_delayed_43__5_, chained_data_delayed_43__4_, chained_data_delayed_43__3_, chained_data_delayed_43__2_, chained_data_delayed_43__1_, chained_data_delayed_43__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_44__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_43__127_, chained_data_delayed_43__126_, chained_data_delayed_43__125_, chained_data_delayed_43__124_, chained_data_delayed_43__123_, chained_data_delayed_43__122_, chained_data_delayed_43__121_, chained_data_delayed_43__120_, chained_data_delayed_43__119_, chained_data_delayed_43__118_, chained_data_delayed_43__117_, chained_data_delayed_43__116_, chained_data_delayed_43__115_, chained_data_delayed_43__114_, chained_data_delayed_43__113_, chained_data_delayed_43__112_, chained_data_delayed_43__111_, chained_data_delayed_43__110_, chained_data_delayed_43__109_, chained_data_delayed_43__108_, chained_data_delayed_43__107_, chained_data_delayed_43__106_, chained_data_delayed_43__105_, chained_data_delayed_43__104_, chained_data_delayed_43__103_, chained_data_delayed_43__102_, chained_data_delayed_43__101_, chained_data_delayed_43__100_, chained_data_delayed_43__99_, chained_data_delayed_43__98_, chained_data_delayed_43__97_, chained_data_delayed_43__96_, chained_data_delayed_43__95_, chained_data_delayed_43__94_, chained_data_delayed_43__93_, chained_data_delayed_43__92_, chained_data_delayed_43__91_, chained_data_delayed_43__90_, chained_data_delayed_43__89_, chained_data_delayed_43__88_, chained_data_delayed_43__87_, chained_data_delayed_43__86_, chained_data_delayed_43__85_, chained_data_delayed_43__84_, chained_data_delayed_43__83_, chained_data_delayed_43__82_, chained_data_delayed_43__81_, chained_data_delayed_43__80_, chained_data_delayed_43__79_, chained_data_delayed_43__78_, chained_data_delayed_43__77_, chained_data_delayed_43__76_, chained_data_delayed_43__75_, chained_data_delayed_43__74_, chained_data_delayed_43__73_, chained_data_delayed_43__72_, chained_data_delayed_43__71_, chained_data_delayed_43__70_, chained_data_delayed_43__69_, chained_data_delayed_43__68_, chained_data_delayed_43__67_, chained_data_delayed_43__66_, chained_data_delayed_43__65_, chained_data_delayed_43__64_, chained_data_delayed_43__63_, chained_data_delayed_43__62_, chained_data_delayed_43__61_, chained_data_delayed_43__60_, chained_data_delayed_43__59_, chained_data_delayed_43__58_, chained_data_delayed_43__57_, chained_data_delayed_43__56_, chained_data_delayed_43__55_, chained_data_delayed_43__54_, chained_data_delayed_43__53_, chained_data_delayed_43__52_, chained_data_delayed_43__51_, chained_data_delayed_43__50_, chained_data_delayed_43__49_, chained_data_delayed_43__48_, chained_data_delayed_43__47_, chained_data_delayed_43__46_, chained_data_delayed_43__45_, chained_data_delayed_43__44_, chained_data_delayed_43__43_, chained_data_delayed_43__42_, chained_data_delayed_43__41_, chained_data_delayed_43__40_, chained_data_delayed_43__39_, chained_data_delayed_43__38_, chained_data_delayed_43__37_, chained_data_delayed_43__36_, chained_data_delayed_43__35_, chained_data_delayed_43__34_, chained_data_delayed_43__33_, chained_data_delayed_43__32_, chained_data_delayed_43__31_, chained_data_delayed_43__30_, chained_data_delayed_43__29_, chained_data_delayed_43__28_, chained_data_delayed_43__27_, chained_data_delayed_43__26_, chained_data_delayed_43__25_, chained_data_delayed_43__24_, chained_data_delayed_43__23_, chained_data_delayed_43__22_, chained_data_delayed_43__21_, chained_data_delayed_43__20_, chained_data_delayed_43__19_, chained_data_delayed_43__18_, chained_data_delayed_43__17_, chained_data_delayed_43__16_, chained_data_delayed_43__15_, chained_data_delayed_43__14_, chained_data_delayed_43__13_, chained_data_delayed_43__12_, chained_data_delayed_43__11_, chained_data_delayed_43__10_, chained_data_delayed_43__9_, chained_data_delayed_43__8_, chained_data_delayed_43__7_, chained_data_delayed_43__6_, chained_data_delayed_43__5_, chained_data_delayed_43__4_, chained_data_delayed_43__3_, chained_data_delayed_43__2_, chained_data_delayed_43__1_, chained_data_delayed_43__0_ }),
    .data_o({ chained_data_delayed_44__127_, chained_data_delayed_44__126_, chained_data_delayed_44__125_, chained_data_delayed_44__124_, chained_data_delayed_44__123_, chained_data_delayed_44__122_, chained_data_delayed_44__121_, chained_data_delayed_44__120_, chained_data_delayed_44__119_, chained_data_delayed_44__118_, chained_data_delayed_44__117_, chained_data_delayed_44__116_, chained_data_delayed_44__115_, chained_data_delayed_44__114_, chained_data_delayed_44__113_, chained_data_delayed_44__112_, chained_data_delayed_44__111_, chained_data_delayed_44__110_, chained_data_delayed_44__109_, chained_data_delayed_44__108_, chained_data_delayed_44__107_, chained_data_delayed_44__106_, chained_data_delayed_44__105_, chained_data_delayed_44__104_, chained_data_delayed_44__103_, chained_data_delayed_44__102_, chained_data_delayed_44__101_, chained_data_delayed_44__100_, chained_data_delayed_44__99_, chained_data_delayed_44__98_, chained_data_delayed_44__97_, chained_data_delayed_44__96_, chained_data_delayed_44__95_, chained_data_delayed_44__94_, chained_data_delayed_44__93_, chained_data_delayed_44__92_, chained_data_delayed_44__91_, chained_data_delayed_44__90_, chained_data_delayed_44__89_, chained_data_delayed_44__88_, chained_data_delayed_44__87_, chained_data_delayed_44__86_, chained_data_delayed_44__85_, chained_data_delayed_44__84_, chained_data_delayed_44__83_, chained_data_delayed_44__82_, chained_data_delayed_44__81_, chained_data_delayed_44__80_, chained_data_delayed_44__79_, chained_data_delayed_44__78_, chained_data_delayed_44__77_, chained_data_delayed_44__76_, chained_data_delayed_44__75_, chained_data_delayed_44__74_, chained_data_delayed_44__73_, chained_data_delayed_44__72_, chained_data_delayed_44__71_, chained_data_delayed_44__70_, chained_data_delayed_44__69_, chained_data_delayed_44__68_, chained_data_delayed_44__67_, chained_data_delayed_44__66_, chained_data_delayed_44__65_, chained_data_delayed_44__64_, chained_data_delayed_44__63_, chained_data_delayed_44__62_, chained_data_delayed_44__61_, chained_data_delayed_44__60_, chained_data_delayed_44__59_, chained_data_delayed_44__58_, chained_data_delayed_44__57_, chained_data_delayed_44__56_, chained_data_delayed_44__55_, chained_data_delayed_44__54_, chained_data_delayed_44__53_, chained_data_delayed_44__52_, chained_data_delayed_44__51_, chained_data_delayed_44__50_, chained_data_delayed_44__49_, chained_data_delayed_44__48_, chained_data_delayed_44__47_, chained_data_delayed_44__46_, chained_data_delayed_44__45_, chained_data_delayed_44__44_, chained_data_delayed_44__43_, chained_data_delayed_44__42_, chained_data_delayed_44__41_, chained_data_delayed_44__40_, chained_data_delayed_44__39_, chained_data_delayed_44__38_, chained_data_delayed_44__37_, chained_data_delayed_44__36_, chained_data_delayed_44__35_, chained_data_delayed_44__34_, chained_data_delayed_44__33_, chained_data_delayed_44__32_, chained_data_delayed_44__31_, chained_data_delayed_44__30_, chained_data_delayed_44__29_, chained_data_delayed_44__28_, chained_data_delayed_44__27_, chained_data_delayed_44__26_, chained_data_delayed_44__25_, chained_data_delayed_44__24_, chained_data_delayed_44__23_, chained_data_delayed_44__22_, chained_data_delayed_44__21_, chained_data_delayed_44__20_, chained_data_delayed_44__19_, chained_data_delayed_44__18_, chained_data_delayed_44__17_, chained_data_delayed_44__16_, chained_data_delayed_44__15_, chained_data_delayed_44__14_, chained_data_delayed_44__13_, chained_data_delayed_44__12_, chained_data_delayed_44__11_, chained_data_delayed_44__10_, chained_data_delayed_44__9_, chained_data_delayed_44__8_, chained_data_delayed_44__7_, chained_data_delayed_44__6_, chained_data_delayed_44__5_, chained_data_delayed_44__4_, chained_data_delayed_44__3_, chained_data_delayed_44__2_, chained_data_delayed_44__1_, chained_data_delayed_44__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_45__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_44__127_, chained_data_delayed_44__126_, chained_data_delayed_44__125_, chained_data_delayed_44__124_, chained_data_delayed_44__123_, chained_data_delayed_44__122_, chained_data_delayed_44__121_, chained_data_delayed_44__120_, chained_data_delayed_44__119_, chained_data_delayed_44__118_, chained_data_delayed_44__117_, chained_data_delayed_44__116_, chained_data_delayed_44__115_, chained_data_delayed_44__114_, chained_data_delayed_44__113_, chained_data_delayed_44__112_, chained_data_delayed_44__111_, chained_data_delayed_44__110_, chained_data_delayed_44__109_, chained_data_delayed_44__108_, chained_data_delayed_44__107_, chained_data_delayed_44__106_, chained_data_delayed_44__105_, chained_data_delayed_44__104_, chained_data_delayed_44__103_, chained_data_delayed_44__102_, chained_data_delayed_44__101_, chained_data_delayed_44__100_, chained_data_delayed_44__99_, chained_data_delayed_44__98_, chained_data_delayed_44__97_, chained_data_delayed_44__96_, chained_data_delayed_44__95_, chained_data_delayed_44__94_, chained_data_delayed_44__93_, chained_data_delayed_44__92_, chained_data_delayed_44__91_, chained_data_delayed_44__90_, chained_data_delayed_44__89_, chained_data_delayed_44__88_, chained_data_delayed_44__87_, chained_data_delayed_44__86_, chained_data_delayed_44__85_, chained_data_delayed_44__84_, chained_data_delayed_44__83_, chained_data_delayed_44__82_, chained_data_delayed_44__81_, chained_data_delayed_44__80_, chained_data_delayed_44__79_, chained_data_delayed_44__78_, chained_data_delayed_44__77_, chained_data_delayed_44__76_, chained_data_delayed_44__75_, chained_data_delayed_44__74_, chained_data_delayed_44__73_, chained_data_delayed_44__72_, chained_data_delayed_44__71_, chained_data_delayed_44__70_, chained_data_delayed_44__69_, chained_data_delayed_44__68_, chained_data_delayed_44__67_, chained_data_delayed_44__66_, chained_data_delayed_44__65_, chained_data_delayed_44__64_, chained_data_delayed_44__63_, chained_data_delayed_44__62_, chained_data_delayed_44__61_, chained_data_delayed_44__60_, chained_data_delayed_44__59_, chained_data_delayed_44__58_, chained_data_delayed_44__57_, chained_data_delayed_44__56_, chained_data_delayed_44__55_, chained_data_delayed_44__54_, chained_data_delayed_44__53_, chained_data_delayed_44__52_, chained_data_delayed_44__51_, chained_data_delayed_44__50_, chained_data_delayed_44__49_, chained_data_delayed_44__48_, chained_data_delayed_44__47_, chained_data_delayed_44__46_, chained_data_delayed_44__45_, chained_data_delayed_44__44_, chained_data_delayed_44__43_, chained_data_delayed_44__42_, chained_data_delayed_44__41_, chained_data_delayed_44__40_, chained_data_delayed_44__39_, chained_data_delayed_44__38_, chained_data_delayed_44__37_, chained_data_delayed_44__36_, chained_data_delayed_44__35_, chained_data_delayed_44__34_, chained_data_delayed_44__33_, chained_data_delayed_44__32_, chained_data_delayed_44__31_, chained_data_delayed_44__30_, chained_data_delayed_44__29_, chained_data_delayed_44__28_, chained_data_delayed_44__27_, chained_data_delayed_44__26_, chained_data_delayed_44__25_, chained_data_delayed_44__24_, chained_data_delayed_44__23_, chained_data_delayed_44__22_, chained_data_delayed_44__21_, chained_data_delayed_44__20_, chained_data_delayed_44__19_, chained_data_delayed_44__18_, chained_data_delayed_44__17_, chained_data_delayed_44__16_, chained_data_delayed_44__15_, chained_data_delayed_44__14_, chained_data_delayed_44__13_, chained_data_delayed_44__12_, chained_data_delayed_44__11_, chained_data_delayed_44__10_, chained_data_delayed_44__9_, chained_data_delayed_44__8_, chained_data_delayed_44__7_, chained_data_delayed_44__6_, chained_data_delayed_44__5_, chained_data_delayed_44__4_, chained_data_delayed_44__3_, chained_data_delayed_44__2_, chained_data_delayed_44__1_, chained_data_delayed_44__0_ }),
    .data_o({ chained_data_delayed_45__127_, chained_data_delayed_45__126_, chained_data_delayed_45__125_, chained_data_delayed_45__124_, chained_data_delayed_45__123_, chained_data_delayed_45__122_, chained_data_delayed_45__121_, chained_data_delayed_45__120_, chained_data_delayed_45__119_, chained_data_delayed_45__118_, chained_data_delayed_45__117_, chained_data_delayed_45__116_, chained_data_delayed_45__115_, chained_data_delayed_45__114_, chained_data_delayed_45__113_, chained_data_delayed_45__112_, chained_data_delayed_45__111_, chained_data_delayed_45__110_, chained_data_delayed_45__109_, chained_data_delayed_45__108_, chained_data_delayed_45__107_, chained_data_delayed_45__106_, chained_data_delayed_45__105_, chained_data_delayed_45__104_, chained_data_delayed_45__103_, chained_data_delayed_45__102_, chained_data_delayed_45__101_, chained_data_delayed_45__100_, chained_data_delayed_45__99_, chained_data_delayed_45__98_, chained_data_delayed_45__97_, chained_data_delayed_45__96_, chained_data_delayed_45__95_, chained_data_delayed_45__94_, chained_data_delayed_45__93_, chained_data_delayed_45__92_, chained_data_delayed_45__91_, chained_data_delayed_45__90_, chained_data_delayed_45__89_, chained_data_delayed_45__88_, chained_data_delayed_45__87_, chained_data_delayed_45__86_, chained_data_delayed_45__85_, chained_data_delayed_45__84_, chained_data_delayed_45__83_, chained_data_delayed_45__82_, chained_data_delayed_45__81_, chained_data_delayed_45__80_, chained_data_delayed_45__79_, chained_data_delayed_45__78_, chained_data_delayed_45__77_, chained_data_delayed_45__76_, chained_data_delayed_45__75_, chained_data_delayed_45__74_, chained_data_delayed_45__73_, chained_data_delayed_45__72_, chained_data_delayed_45__71_, chained_data_delayed_45__70_, chained_data_delayed_45__69_, chained_data_delayed_45__68_, chained_data_delayed_45__67_, chained_data_delayed_45__66_, chained_data_delayed_45__65_, chained_data_delayed_45__64_, chained_data_delayed_45__63_, chained_data_delayed_45__62_, chained_data_delayed_45__61_, chained_data_delayed_45__60_, chained_data_delayed_45__59_, chained_data_delayed_45__58_, chained_data_delayed_45__57_, chained_data_delayed_45__56_, chained_data_delayed_45__55_, chained_data_delayed_45__54_, chained_data_delayed_45__53_, chained_data_delayed_45__52_, chained_data_delayed_45__51_, chained_data_delayed_45__50_, chained_data_delayed_45__49_, chained_data_delayed_45__48_, chained_data_delayed_45__47_, chained_data_delayed_45__46_, chained_data_delayed_45__45_, chained_data_delayed_45__44_, chained_data_delayed_45__43_, chained_data_delayed_45__42_, chained_data_delayed_45__41_, chained_data_delayed_45__40_, chained_data_delayed_45__39_, chained_data_delayed_45__38_, chained_data_delayed_45__37_, chained_data_delayed_45__36_, chained_data_delayed_45__35_, chained_data_delayed_45__34_, chained_data_delayed_45__33_, chained_data_delayed_45__32_, chained_data_delayed_45__31_, chained_data_delayed_45__30_, chained_data_delayed_45__29_, chained_data_delayed_45__28_, chained_data_delayed_45__27_, chained_data_delayed_45__26_, chained_data_delayed_45__25_, chained_data_delayed_45__24_, chained_data_delayed_45__23_, chained_data_delayed_45__22_, chained_data_delayed_45__21_, chained_data_delayed_45__20_, chained_data_delayed_45__19_, chained_data_delayed_45__18_, chained_data_delayed_45__17_, chained_data_delayed_45__16_, chained_data_delayed_45__15_, chained_data_delayed_45__14_, chained_data_delayed_45__13_, chained_data_delayed_45__12_, chained_data_delayed_45__11_, chained_data_delayed_45__10_, chained_data_delayed_45__9_, chained_data_delayed_45__8_, chained_data_delayed_45__7_, chained_data_delayed_45__6_, chained_data_delayed_45__5_, chained_data_delayed_45__4_, chained_data_delayed_45__3_, chained_data_delayed_45__2_, chained_data_delayed_45__1_, chained_data_delayed_45__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_46__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_45__127_, chained_data_delayed_45__126_, chained_data_delayed_45__125_, chained_data_delayed_45__124_, chained_data_delayed_45__123_, chained_data_delayed_45__122_, chained_data_delayed_45__121_, chained_data_delayed_45__120_, chained_data_delayed_45__119_, chained_data_delayed_45__118_, chained_data_delayed_45__117_, chained_data_delayed_45__116_, chained_data_delayed_45__115_, chained_data_delayed_45__114_, chained_data_delayed_45__113_, chained_data_delayed_45__112_, chained_data_delayed_45__111_, chained_data_delayed_45__110_, chained_data_delayed_45__109_, chained_data_delayed_45__108_, chained_data_delayed_45__107_, chained_data_delayed_45__106_, chained_data_delayed_45__105_, chained_data_delayed_45__104_, chained_data_delayed_45__103_, chained_data_delayed_45__102_, chained_data_delayed_45__101_, chained_data_delayed_45__100_, chained_data_delayed_45__99_, chained_data_delayed_45__98_, chained_data_delayed_45__97_, chained_data_delayed_45__96_, chained_data_delayed_45__95_, chained_data_delayed_45__94_, chained_data_delayed_45__93_, chained_data_delayed_45__92_, chained_data_delayed_45__91_, chained_data_delayed_45__90_, chained_data_delayed_45__89_, chained_data_delayed_45__88_, chained_data_delayed_45__87_, chained_data_delayed_45__86_, chained_data_delayed_45__85_, chained_data_delayed_45__84_, chained_data_delayed_45__83_, chained_data_delayed_45__82_, chained_data_delayed_45__81_, chained_data_delayed_45__80_, chained_data_delayed_45__79_, chained_data_delayed_45__78_, chained_data_delayed_45__77_, chained_data_delayed_45__76_, chained_data_delayed_45__75_, chained_data_delayed_45__74_, chained_data_delayed_45__73_, chained_data_delayed_45__72_, chained_data_delayed_45__71_, chained_data_delayed_45__70_, chained_data_delayed_45__69_, chained_data_delayed_45__68_, chained_data_delayed_45__67_, chained_data_delayed_45__66_, chained_data_delayed_45__65_, chained_data_delayed_45__64_, chained_data_delayed_45__63_, chained_data_delayed_45__62_, chained_data_delayed_45__61_, chained_data_delayed_45__60_, chained_data_delayed_45__59_, chained_data_delayed_45__58_, chained_data_delayed_45__57_, chained_data_delayed_45__56_, chained_data_delayed_45__55_, chained_data_delayed_45__54_, chained_data_delayed_45__53_, chained_data_delayed_45__52_, chained_data_delayed_45__51_, chained_data_delayed_45__50_, chained_data_delayed_45__49_, chained_data_delayed_45__48_, chained_data_delayed_45__47_, chained_data_delayed_45__46_, chained_data_delayed_45__45_, chained_data_delayed_45__44_, chained_data_delayed_45__43_, chained_data_delayed_45__42_, chained_data_delayed_45__41_, chained_data_delayed_45__40_, chained_data_delayed_45__39_, chained_data_delayed_45__38_, chained_data_delayed_45__37_, chained_data_delayed_45__36_, chained_data_delayed_45__35_, chained_data_delayed_45__34_, chained_data_delayed_45__33_, chained_data_delayed_45__32_, chained_data_delayed_45__31_, chained_data_delayed_45__30_, chained_data_delayed_45__29_, chained_data_delayed_45__28_, chained_data_delayed_45__27_, chained_data_delayed_45__26_, chained_data_delayed_45__25_, chained_data_delayed_45__24_, chained_data_delayed_45__23_, chained_data_delayed_45__22_, chained_data_delayed_45__21_, chained_data_delayed_45__20_, chained_data_delayed_45__19_, chained_data_delayed_45__18_, chained_data_delayed_45__17_, chained_data_delayed_45__16_, chained_data_delayed_45__15_, chained_data_delayed_45__14_, chained_data_delayed_45__13_, chained_data_delayed_45__12_, chained_data_delayed_45__11_, chained_data_delayed_45__10_, chained_data_delayed_45__9_, chained_data_delayed_45__8_, chained_data_delayed_45__7_, chained_data_delayed_45__6_, chained_data_delayed_45__5_, chained_data_delayed_45__4_, chained_data_delayed_45__3_, chained_data_delayed_45__2_, chained_data_delayed_45__1_, chained_data_delayed_45__0_ }),
    .data_o({ chained_data_delayed_46__127_, chained_data_delayed_46__126_, chained_data_delayed_46__125_, chained_data_delayed_46__124_, chained_data_delayed_46__123_, chained_data_delayed_46__122_, chained_data_delayed_46__121_, chained_data_delayed_46__120_, chained_data_delayed_46__119_, chained_data_delayed_46__118_, chained_data_delayed_46__117_, chained_data_delayed_46__116_, chained_data_delayed_46__115_, chained_data_delayed_46__114_, chained_data_delayed_46__113_, chained_data_delayed_46__112_, chained_data_delayed_46__111_, chained_data_delayed_46__110_, chained_data_delayed_46__109_, chained_data_delayed_46__108_, chained_data_delayed_46__107_, chained_data_delayed_46__106_, chained_data_delayed_46__105_, chained_data_delayed_46__104_, chained_data_delayed_46__103_, chained_data_delayed_46__102_, chained_data_delayed_46__101_, chained_data_delayed_46__100_, chained_data_delayed_46__99_, chained_data_delayed_46__98_, chained_data_delayed_46__97_, chained_data_delayed_46__96_, chained_data_delayed_46__95_, chained_data_delayed_46__94_, chained_data_delayed_46__93_, chained_data_delayed_46__92_, chained_data_delayed_46__91_, chained_data_delayed_46__90_, chained_data_delayed_46__89_, chained_data_delayed_46__88_, chained_data_delayed_46__87_, chained_data_delayed_46__86_, chained_data_delayed_46__85_, chained_data_delayed_46__84_, chained_data_delayed_46__83_, chained_data_delayed_46__82_, chained_data_delayed_46__81_, chained_data_delayed_46__80_, chained_data_delayed_46__79_, chained_data_delayed_46__78_, chained_data_delayed_46__77_, chained_data_delayed_46__76_, chained_data_delayed_46__75_, chained_data_delayed_46__74_, chained_data_delayed_46__73_, chained_data_delayed_46__72_, chained_data_delayed_46__71_, chained_data_delayed_46__70_, chained_data_delayed_46__69_, chained_data_delayed_46__68_, chained_data_delayed_46__67_, chained_data_delayed_46__66_, chained_data_delayed_46__65_, chained_data_delayed_46__64_, chained_data_delayed_46__63_, chained_data_delayed_46__62_, chained_data_delayed_46__61_, chained_data_delayed_46__60_, chained_data_delayed_46__59_, chained_data_delayed_46__58_, chained_data_delayed_46__57_, chained_data_delayed_46__56_, chained_data_delayed_46__55_, chained_data_delayed_46__54_, chained_data_delayed_46__53_, chained_data_delayed_46__52_, chained_data_delayed_46__51_, chained_data_delayed_46__50_, chained_data_delayed_46__49_, chained_data_delayed_46__48_, chained_data_delayed_46__47_, chained_data_delayed_46__46_, chained_data_delayed_46__45_, chained_data_delayed_46__44_, chained_data_delayed_46__43_, chained_data_delayed_46__42_, chained_data_delayed_46__41_, chained_data_delayed_46__40_, chained_data_delayed_46__39_, chained_data_delayed_46__38_, chained_data_delayed_46__37_, chained_data_delayed_46__36_, chained_data_delayed_46__35_, chained_data_delayed_46__34_, chained_data_delayed_46__33_, chained_data_delayed_46__32_, chained_data_delayed_46__31_, chained_data_delayed_46__30_, chained_data_delayed_46__29_, chained_data_delayed_46__28_, chained_data_delayed_46__27_, chained_data_delayed_46__26_, chained_data_delayed_46__25_, chained_data_delayed_46__24_, chained_data_delayed_46__23_, chained_data_delayed_46__22_, chained_data_delayed_46__21_, chained_data_delayed_46__20_, chained_data_delayed_46__19_, chained_data_delayed_46__18_, chained_data_delayed_46__17_, chained_data_delayed_46__16_, chained_data_delayed_46__15_, chained_data_delayed_46__14_, chained_data_delayed_46__13_, chained_data_delayed_46__12_, chained_data_delayed_46__11_, chained_data_delayed_46__10_, chained_data_delayed_46__9_, chained_data_delayed_46__8_, chained_data_delayed_46__7_, chained_data_delayed_46__6_, chained_data_delayed_46__5_, chained_data_delayed_46__4_, chained_data_delayed_46__3_, chained_data_delayed_46__2_, chained_data_delayed_46__1_, chained_data_delayed_46__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_47__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_46__127_, chained_data_delayed_46__126_, chained_data_delayed_46__125_, chained_data_delayed_46__124_, chained_data_delayed_46__123_, chained_data_delayed_46__122_, chained_data_delayed_46__121_, chained_data_delayed_46__120_, chained_data_delayed_46__119_, chained_data_delayed_46__118_, chained_data_delayed_46__117_, chained_data_delayed_46__116_, chained_data_delayed_46__115_, chained_data_delayed_46__114_, chained_data_delayed_46__113_, chained_data_delayed_46__112_, chained_data_delayed_46__111_, chained_data_delayed_46__110_, chained_data_delayed_46__109_, chained_data_delayed_46__108_, chained_data_delayed_46__107_, chained_data_delayed_46__106_, chained_data_delayed_46__105_, chained_data_delayed_46__104_, chained_data_delayed_46__103_, chained_data_delayed_46__102_, chained_data_delayed_46__101_, chained_data_delayed_46__100_, chained_data_delayed_46__99_, chained_data_delayed_46__98_, chained_data_delayed_46__97_, chained_data_delayed_46__96_, chained_data_delayed_46__95_, chained_data_delayed_46__94_, chained_data_delayed_46__93_, chained_data_delayed_46__92_, chained_data_delayed_46__91_, chained_data_delayed_46__90_, chained_data_delayed_46__89_, chained_data_delayed_46__88_, chained_data_delayed_46__87_, chained_data_delayed_46__86_, chained_data_delayed_46__85_, chained_data_delayed_46__84_, chained_data_delayed_46__83_, chained_data_delayed_46__82_, chained_data_delayed_46__81_, chained_data_delayed_46__80_, chained_data_delayed_46__79_, chained_data_delayed_46__78_, chained_data_delayed_46__77_, chained_data_delayed_46__76_, chained_data_delayed_46__75_, chained_data_delayed_46__74_, chained_data_delayed_46__73_, chained_data_delayed_46__72_, chained_data_delayed_46__71_, chained_data_delayed_46__70_, chained_data_delayed_46__69_, chained_data_delayed_46__68_, chained_data_delayed_46__67_, chained_data_delayed_46__66_, chained_data_delayed_46__65_, chained_data_delayed_46__64_, chained_data_delayed_46__63_, chained_data_delayed_46__62_, chained_data_delayed_46__61_, chained_data_delayed_46__60_, chained_data_delayed_46__59_, chained_data_delayed_46__58_, chained_data_delayed_46__57_, chained_data_delayed_46__56_, chained_data_delayed_46__55_, chained_data_delayed_46__54_, chained_data_delayed_46__53_, chained_data_delayed_46__52_, chained_data_delayed_46__51_, chained_data_delayed_46__50_, chained_data_delayed_46__49_, chained_data_delayed_46__48_, chained_data_delayed_46__47_, chained_data_delayed_46__46_, chained_data_delayed_46__45_, chained_data_delayed_46__44_, chained_data_delayed_46__43_, chained_data_delayed_46__42_, chained_data_delayed_46__41_, chained_data_delayed_46__40_, chained_data_delayed_46__39_, chained_data_delayed_46__38_, chained_data_delayed_46__37_, chained_data_delayed_46__36_, chained_data_delayed_46__35_, chained_data_delayed_46__34_, chained_data_delayed_46__33_, chained_data_delayed_46__32_, chained_data_delayed_46__31_, chained_data_delayed_46__30_, chained_data_delayed_46__29_, chained_data_delayed_46__28_, chained_data_delayed_46__27_, chained_data_delayed_46__26_, chained_data_delayed_46__25_, chained_data_delayed_46__24_, chained_data_delayed_46__23_, chained_data_delayed_46__22_, chained_data_delayed_46__21_, chained_data_delayed_46__20_, chained_data_delayed_46__19_, chained_data_delayed_46__18_, chained_data_delayed_46__17_, chained_data_delayed_46__16_, chained_data_delayed_46__15_, chained_data_delayed_46__14_, chained_data_delayed_46__13_, chained_data_delayed_46__12_, chained_data_delayed_46__11_, chained_data_delayed_46__10_, chained_data_delayed_46__9_, chained_data_delayed_46__8_, chained_data_delayed_46__7_, chained_data_delayed_46__6_, chained_data_delayed_46__5_, chained_data_delayed_46__4_, chained_data_delayed_46__3_, chained_data_delayed_46__2_, chained_data_delayed_46__1_, chained_data_delayed_46__0_ }),
    .data_o({ chained_data_delayed_47__127_, chained_data_delayed_47__126_, chained_data_delayed_47__125_, chained_data_delayed_47__124_, chained_data_delayed_47__123_, chained_data_delayed_47__122_, chained_data_delayed_47__121_, chained_data_delayed_47__120_, chained_data_delayed_47__119_, chained_data_delayed_47__118_, chained_data_delayed_47__117_, chained_data_delayed_47__116_, chained_data_delayed_47__115_, chained_data_delayed_47__114_, chained_data_delayed_47__113_, chained_data_delayed_47__112_, chained_data_delayed_47__111_, chained_data_delayed_47__110_, chained_data_delayed_47__109_, chained_data_delayed_47__108_, chained_data_delayed_47__107_, chained_data_delayed_47__106_, chained_data_delayed_47__105_, chained_data_delayed_47__104_, chained_data_delayed_47__103_, chained_data_delayed_47__102_, chained_data_delayed_47__101_, chained_data_delayed_47__100_, chained_data_delayed_47__99_, chained_data_delayed_47__98_, chained_data_delayed_47__97_, chained_data_delayed_47__96_, chained_data_delayed_47__95_, chained_data_delayed_47__94_, chained_data_delayed_47__93_, chained_data_delayed_47__92_, chained_data_delayed_47__91_, chained_data_delayed_47__90_, chained_data_delayed_47__89_, chained_data_delayed_47__88_, chained_data_delayed_47__87_, chained_data_delayed_47__86_, chained_data_delayed_47__85_, chained_data_delayed_47__84_, chained_data_delayed_47__83_, chained_data_delayed_47__82_, chained_data_delayed_47__81_, chained_data_delayed_47__80_, chained_data_delayed_47__79_, chained_data_delayed_47__78_, chained_data_delayed_47__77_, chained_data_delayed_47__76_, chained_data_delayed_47__75_, chained_data_delayed_47__74_, chained_data_delayed_47__73_, chained_data_delayed_47__72_, chained_data_delayed_47__71_, chained_data_delayed_47__70_, chained_data_delayed_47__69_, chained_data_delayed_47__68_, chained_data_delayed_47__67_, chained_data_delayed_47__66_, chained_data_delayed_47__65_, chained_data_delayed_47__64_, chained_data_delayed_47__63_, chained_data_delayed_47__62_, chained_data_delayed_47__61_, chained_data_delayed_47__60_, chained_data_delayed_47__59_, chained_data_delayed_47__58_, chained_data_delayed_47__57_, chained_data_delayed_47__56_, chained_data_delayed_47__55_, chained_data_delayed_47__54_, chained_data_delayed_47__53_, chained_data_delayed_47__52_, chained_data_delayed_47__51_, chained_data_delayed_47__50_, chained_data_delayed_47__49_, chained_data_delayed_47__48_, chained_data_delayed_47__47_, chained_data_delayed_47__46_, chained_data_delayed_47__45_, chained_data_delayed_47__44_, chained_data_delayed_47__43_, chained_data_delayed_47__42_, chained_data_delayed_47__41_, chained_data_delayed_47__40_, chained_data_delayed_47__39_, chained_data_delayed_47__38_, chained_data_delayed_47__37_, chained_data_delayed_47__36_, chained_data_delayed_47__35_, chained_data_delayed_47__34_, chained_data_delayed_47__33_, chained_data_delayed_47__32_, chained_data_delayed_47__31_, chained_data_delayed_47__30_, chained_data_delayed_47__29_, chained_data_delayed_47__28_, chained_data_delayed_47__27_, chained_data_delayed_47__26_, chained_data_delayed_47__25_, chained_data_delayed_47__24_, chained_data_delayed_47__23_, chained_data_delayed_47__22_, chained_data_delayed_47__21_, chained_data_delayed_47__20_, chained_data_delayed_47__19_, chained_data_delayed_47__18_, chained_data_delayed_47__17_, chained_data_delayed_47__16_, chained_data_delayed_47__15_, chained_data_delayed_47__14_, chained_data_delayed_47__13_, chained_data_delayed_47__12_, chained_data_delayed_47__11_, chained_data_delayed_47__10_, chained_data_delayed_47__9_, chained_data_delayed_47__8_, chained_data_delayed_47__7_, chained_data_delayed_47__6_, chained_data_delayed_47__5_, chained_data_delayed_47__4_, chained_data_delayed_47__3_, chained_data_delayed_47__2_, chained_data_delayed_47__1_, chained_data_delayed_47__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_48__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_47__127_, chained_data_delayed_47__126_, chained_data_delayed_47__125_, chained_data_delayed_47__124_, chained_data_delayed_47__123_, chained_data_delayed_47__122_, chained_data_delayed_47__121_, chained_data_delayed_47__120_, chained_data_delayed_47__119_, chained_data_delayed_47__118_, chained_data_delayed_47__117_, chained_data_delayed_47__116_, chained_data_delayed_47__115_, chained_data_delayed_47__114_, chained_data_delayed_47__113_, chained_data_delayed_47__112_, chained_data_delayed_47__111_, chained_data_delayed_47__110_, chained_data_delayed_47__109_, chained_data_delayed_47__108_, chained_data_delayed_47__107_, chained_data_delayed_47__106_, chained_data_delayed_47__105_, chained_data_delayed_47__104_, chained_data_delayed_47__103_, chained_data_delayed_47__102_, chained_data_delayed_47__101_, chained_data_delayed_47__100_, chained_data_delayed_47__99_, chained_data_delayed_47__98_, chained_data_delayed_47__97_, chained_data_delayed_47__96_, chained_data_delayed_47__95_, chained_data_delayed_47__94_, chained_data_delayed_47__93_, chained_data_delayed_47__92_, chained_data_delayed_47__91_, chained_data_delayed_47__90_, chained_data_delayed_47__89_, chained_data_delayed_47__88_, chained_data_delayed_47__87_, chained_data_delayed_47__86_, chained_data_delayed_47__85_, chained_data_delayed_47__84_, chained_data_delayed_47__83_, chained_data_delayed_47__82_, chained_data_delayed_47__81_, chained_data_delayed_47__80_, chained_data_delayed_47__79_, chained_data_delayed_47__78_, chained_data_delayed_47__77_, chained_data_delayed_47__76_, chained_data_delayed_47__75_, chained_data_delayed_47__74_, chained_data_delayed_47__73_, chained_data_delayed_47__72_, chained_data_delayed_47__71_, chained_data_delayed_47__70_, chained_data_delayed_47__69_, chained_data_delayed_47__68_, chained_data_delayed_47__67_, chained_data_delayed_47__66_, chained_data_delayed_47__65_, chained_data_delayed_47__64_, chained_data_delayed_47__63_, chained_data_delayed_47__62_, chained_data_delayed_47__61_, chained_data_delayed_47__60_, chained_data_delayed_47__59_, chained_data_delayed_47__58_, chained_data_delayed_47__57_, chained_data_delayed_47__56_, chained_data_delayed_47__55_, chained_data_delayed_47__54_, chained_data_delayed_47__53_, chained_data_delayed_47__52_, chained_data_delayed_47__51_, chained_data_delayed_47__50_, chained_data_delayed_47__49_, chained_data_delayed_47__48_, chained_data_delayed_47__47_, chained_data_delayed_47__46_, chained_data_delayed_47__45_, chained_data_delayed_47__44_, chained_data_delayed_47__43_, chained_data_delayed_47__42_, chained_data_delayed_47__41_, chained_data_delayed_47__40_, chained_data_delayed_47__39_, chained_data_delayed_47__38_, chained_data_delayed_47__37_, chained_data_delayed_47__36_, chained_data_delayed_47__35_, chained_data_delayed_47__34_, chained_data_delayed_47__33_, chained_data_delayed_47__32_, chained_data_delayed_47__31_, chained_data_delayed_47__30_, chained_data_delayed_47__29_, chained_data_delayed_47__28_, chained_data_delayed_47__27_, chained_data_delayed_47__26_, chained_data_delayed_47__25_, chained_data_delayed_47__24_, chained_data_delayed_47__23_, chained_data_delayed_47__22_, chained_data_delayed_47__21_, chained_data_delayed_47__20_, chained_data_delayed_47__19_, chained_data_delayed_47__18_, chained_data_delayed_47__17_, chained_data_delayed_47__16_, chained_data_delayed_47__15_, chained_data_delayed_47__14_, chained_data_delayed_47__13_, chained_data_delayed_47__12_, chained_data_delayed_47__11_, chained_data_delayed_47__10_, chained_data_delayed_47__9_, chained_data_delayed_47__8_, chained_data_delayed_47__7_, chained_data_delayed_47__6_, chained_data_delayed_47__5_, chained_data_delayed_47__4_, chained_data_delayed_47__3_, chained_data_delayed_47__2_, chained_data_delayed_47__1_, chained_data_delayed_47__0_ }),
    .data_o({ chained_data_delayed_48__127_, chained_data_delayed_48__126_, chained_data_delayed_48__125_, chained_data_delayed_48__124_, chained_data_delayed_48__123_, chained_data_delayed_48__122_, chained_data_delayed_48__121_, chained_data_delayed_48__120_, chained_data_delayed_48__119_, chained_data_delayed_48__118_, chained_data_delayed_48__117_, chained_data_delayed_48__116_, chained_data_delayed_48__115_, chained_data_delayed_48__114_, chained_data_delayed_48__113_, chained_data_delayed_48__112_, chained_data_delayed_48__111_, chained_data_delayed_48__110_, chained_data_delayed_48__109_, chained_data_delayed_48__108_, chained_data_delayed_48__107_, chained_data_delayed_48__106_, chained_data_delayed_48__105_, chained_data_delayed_48__104_, chained_data_delayed_48__103_, chained_data_delayed_48__102_, chained_data_delayed_48__101_, chained_data_delayed_48__100_, chained_data_delayed_48__99_, chained_data_delayed_48__98_, chained_data_delayed_48__97_, chained_data_delayed_48__96_, chained_data_delayed_48__95_, chained_data_delayed_48__94_, chained_data_delayed_48__93_, chained_data_delayed_48__92_, chained_data_delayed_48__91_, chained_data_delayed_48__90_, chained_data_delayed_48__89_, chained_data_delayed_48__88_, chained_data_delayed_48__87_, chained_data_delayed_48__86_, chained_data_delayed_48__85_, chained_data_delayed_48__84_, chained_data_delayed_48__83_, chained_data_delayed_48__82_, chained_data_delayed_48__81_, chained_data_delayed_48__80_, chained_data_delayed_48__79_, chained_data_delayed_48__78_, chained_data_delayed_48__77_, chained_data_delayed_48__76_, chained_data_delayed_48__75_, chained_data_delayed_48__74_, chained_data_delayed_48__73_, chained_data_delayed_48__72_, chained_data_delayed_48__71_, chained_data_delayed_48__70_, chained_data_delayed_48__69_, chained_data_delayed_48__68_, chained_data_delayed_48__67_, chained_data_delayed_48__66_, chained_data_delayed_48__65_, chained_data_delayed_48__64_, chained_data_delayed_48__63_, chained_data_delayed_48__62_, chained_data_delayed_48__61_, chained_data_delayed_48__60_, chained_data_delayed_48__59_, chained_data_delayed_48__58_, chained_data_delayed_48__57_, chained_data_delayed_48__56_, chained_data_delayed_48__55_, chained_data_delayed_48__54_, chained_data_delayed_48__53_, chained_data_delayed_48__52_, chained_data_delayed_48__51_, chained_data_delayed_48__50_, chained_data_delayed_48__49_, chained_data_delayed_48__48_, chained_data_delayed_48__47_, chained_data_delayed_48__46_, chained_data_delayed_48__45_, chained_data_delayed_48__44_, chained_data_delayed_48__43_, chained_data_delayed_48__42_, chained_data_delayed_48__41_, chained_data_delayed_48__40_, chained_data_delayed_48__39_, chained_data_delayed_48__38_, chained_data_delayed_48__37_, chained_data_delayed_48__36_, chained_data_delayed_48__35_, chained_data_delayed_48__34_, chained_data_delayed_48__33_, chained_data_delayed_48__32_, chained_data_delayed_48__31_, chained_data_delayed_48__30_, chained_data_delayed_48__29_, chained_data_delayed_48__28_, chained_data_delayed_48__27_, chained_data_delayed_48__26_, chained_data_delayed_48__25_, chained_data_delayed_48__24_, chained_data_delayed_48__23_, chained_data_delayed_48__22_, chained_data_delayed_48__21_, chained_data_delayed_48__20_, chained_data_delayed_48__19_, chained_data_delayed_48__18_, chained_data_delayed_48__17_, chained_data_delayed_48__16_, chained_data_delayed_48__15_, chained_data_delayed_48__14_, chained_data_delayed_48__13_, chained_data_delayed_48__12_, chained_data_delayed_48__11_, chained_data_delayed_48__10_, chained_data_delayed_48__9_, chained_data_delayed_48__8_, chained_data_delayed_48__7_, chained_data_delayed_48__6_, chained_data_delayed_48__5_, chained_data_delayed_48__4_, chained_data_delayed_48__3_, chained_data_delayed_48__2_, chained_data_delayed_48__1_, chained_data_delayed_48__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_49__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_48__127_, chained_data_delayed_48__126_, chained_data_delayed_48__125_, chained_data_delayed_48__124_, chained_data_delayed_48__123_, chained_data_delayed_48__122_, chained_data_delayed_48__121_, chained_data_delayed_48__120_, chained_data_delayed_48__119_, chained_data_delayed_48__118_, chained_data_delayed_48__117_, chained_data_delayed_48__116_, chained_data_delayed_48__115_, chained_data_delayed_48__114_, chained_data_delayed_48__113_, chained_data_delayed_48__112_, chained_data_delayed_48__111_, chained_data_delayed_48__110_, chained_data_delayed_48__109_, chained_data_delayed_48__108_, chained_data_delayed_48__107_, chained_data_delayed_48__106_, chained_data_delayed_48__105_, chained_data_delayed_48__104_, chained_data_delayed_48__103_, chained_data_delayed_48__102_, chained_data_delayed_48__101_, chained_data_delayed_48__100_, chained_data_delayed_48__99_, chained_data_delayed_48__98_, chained_data_delayed_48__97_, chained_data_delayed_48__96_, chained_data_delayed_48__95_, chained_data_delayed_48__94_, chained_data_delayed_48__93_, chained_data_delayed_48__92_, chained_data_delayed_48__91_, chained_data_delayed_48__90_, chained_data_delayed_48__89_, chained_data_delayed_48__88_, chained_data_delayed_48__87_, chained_data_delayed_48__86_, chained_data_delayed_48__85_, chained_data_delayed_48__84_, chained_data_delayed_48__83_, chained_data_delayed_48__82_, chained_data_delayed_48__81_, chained_data_delayed_48__80_, chained_data_delayed_48__79_, chained_data_delayed_48__78_, chained_data_delayed_48__77_, chained_data_delayed_48__76_, chained_data_delayed_48__75_, chained_data_delayed_48__74_, chained_data_delayed_48__73_, chained_data_delayed_48__72_, chained_data_delayed_48__71_, chained_data_delayed_48__70_, chained_data_delayed_48__69_, chained_data_delayed_48__68_, chained_data_delayed_48__67_, chained_data_delayed_48__66_, chained_data_delayed_48__65_, chained_data_delayed_48__64_, chained_data_delayed_48__63_, chained_data_delayed_48__62_, chained_data_delayed_48__61_, chained_data_delayed_48__60_, chained_data_delayed_48__59_, chained_data_delayed_48__58_, chained_data_delayed_48__57_, chained_data_delayed_48__56_, chained_data_delayed_48__55_, chained_data_delayed_48__54_, chained_data_delayed_48__53_, chained_data_delayed_48__52_, chained_data_delayed_48__51_, chained_data_delayed_48__50_, chained_data_delayed_48__49_, chained_data_delayed_48__48_, chained_data_delayed_48__47_, chained_data_delayed_48__46_, chained_data_delayed_48__45_, chained_data_delayed_48__44_, chained_data_delayed_48__43_, chained_data_delayed_48__42_, chained_data_delayed_48__41_, chained_data_delayed_48__40_, chained_data_delayed_48__39_, chained_data_delayed_48__38_, chained_data_delayed_48__37_, chained_data_delayed_48__36_, chained_data_delayed_48__35_, chained_data_delayed_48__34_, chained_data_delayed_48__33_, chained_data_delayed_48__32_, chained_data_delayed_48__31_, chained_data_delayed_48__30_, chained_data_delayed_48__29_, chained_data_delayed_48__28_, chained_data_delayed_48__27_, chained_data_delayed_48__26_, chained_data_delayed_48__25_, chained_data_delayed_48__24_, chained_data_delayed_48__23_, chained_data_delayed_48__22_, chained_data_delayed_48__21_, chained_data_delayed_48__20_, chained_data_delayed_48__19_, chained_data_delayed_48__18_, chained_data_delayed_48__17_, chained_data_delayed_48__16_, chained_data_delayed_48__15_, chained_data_delayed_48__14_, chained_data_delayed_48__13_, chained_data_delayed_48__12_, chained_data_delayed_48__11_, chained_data_delayed_48__10_, chained_data_delayed_48__9_, chained_data_delayed_48__8_, chained_data_delayed_48__7_, chained_data_delayed_48__6_, chained_data_delayed_48__5_, chained_data_delayed_48__4_, chained_data_delayed_48__3_, chained_data_delayed_48__2_, chained_data_delayed_48__1_, chained_data_delayed_48__0_ }),
    .data_o({ chained_data_delayed_49__127_, chained_data_delayed_49__126_, chained_data_delayed_49__125_, chained_data_delayed_49__124_, chained_data_delayed_49__123_, chained_data_delayed_49__122_, chained_data_delayed_49__121_, chained_data_delayed_49__120_, chained_data_delayed_49__119_, chained_data_delayed_49__118_, chained_data_delayed_49__117_, chained_data_delayed_49__116_, chained_data_delayed_49__115_, chained_data_delayed_49__114_, chained_data_delayed_49__113_, chained_data_delayed_49__112_, chained_data_delayed_49__111_, chained_data_delayed_49__110_, chained_data_delayed_49__109_, chained_data_delayed_49__108_, chained_data_delayed_49__107_, chained_data_delayed_49__106_, chained_data_delayed_49__105_, chained_data_delayed_49__104_, chained_data_delayed_49__103_, chained_data_delayed_49__102_, chained_data_delayed_49__101_, chained_data_delayed_49__100_, chained_data_delayed_49__99_, chained_data_delayed_49__98_, chained_data_delayed_49__97_, chained_data_delayed_49__96_, chained_data_delayed_49__95_, chained_data_delayed_49__94_, chained_data_delayed_49__93_, chained_data_delayed_49__92_, chained_data_delayed_49__91_, chained_data_delayed_49__90_, chained_data_delayed_49__89_, chained_data_delayed_49__88_, chained_data_delayed_49__87_, chained_data_delayed_49__86_, chained_data_delayed_49__85_, chained_data_delayed_49__84_, chained_data_delayed_49__83_, chained_data_delayed_49__82_, chained_data_delayed_49__81_, chained_data_delayed_49__80_, chained_data_delayed_49__79_, chained_data_delayed_49__78_, chained_data_delayed_49__77_, chained_data_delayed_49__76_, chained_data_delayed_49__75_, chained_data_delayed_49__74_, chained_data_delayed_49__73_, chained_data_delayed_49__72_, chained_data_delayed_49__71_, chained_data_delayed_49__70_, chained_data_delayed_49__69_, chained_data_delayed_49__68_, chained_data_delayed_49__67_, chained_data_delayed_49__66_, chained_data_delayed_49__65_, chained_data_delayed_49__64_, chained_data_delayed_49__63_, chained_data_delayed_49__62_, chained_data_delayed_49__61_, chained_data_delayed_49__60_, chained_data_delayed_49__59_, chained_data_delayed_49__58_, chained_data_delayed_49__57_, chained_data_delayed_49__56_, chained_data_delayed_49__55_, chained_data_delayed_49__54_, chained_data_delayed_49__53_, chained_data_delayed_49__52_, chained_data_delayed_49__51_, chained_data_delayed_49__50_, chained_data_delayed_49__49_, chained_data_delayed_49__48_, chained_data_delayed_49__47_, chained_data_delayed_49__46_, chained_data_delayed_49__45_, chained_data_delayed_49__44_, chained_data_delayed_49__43_, chained_data_delayed_49__42_, chained_data_delayed_49__41_, chained_data_delayed_49__40_, chained_data_delayed_49__39_, chained_data_delayed_49__38_, chained_data_delayed_49__37_, chained_data_delayed_49__36_, chained_data_delayed_49__35_, chained_data_delayed_49__34_, chained_data_delayed_49__33_, chained_data_delayed_49__32_, chained_data_delayed_49__31_, chained_data_delayed_49__30_, chained_data_delayed_49__29_, chained_data_delayed_49__28_, chained_data_delayed_49__27_, chained_data_delayed_49__26_, chained_data_delayed_49__25_, chained_data_delayed_49__24_, chained_data_delayed_49__23_, chained_data_delayed_49__22_, chained_data_delayed_49__21_, chained_data_delayed_49__20_, chained_data_delayed_49__19_, chained_data_delayed_49__18_, chained_data_delayed_49__17_, chained_data_delayed_49__16_, chained_data_delayed_49__15_, chained_data_delayed_49__14_, chained_data_delayed_49__13_, chained_data_delayed_49__12_, chained_data_delayed_49__11_, chained_data_delayed_49__10_, chained_data_delayed_49__9_, chained_data_delayed_49__8_, chained_data_delayed_49__7_, chained_data_delayed_49__6_, chained_data_delayed_49__5_, chained_data_delayed_49__4_, chained_data_delayed_49__3_, chained_data_delayed_49__2_, chained_data_delayed_49__1_, chained_data_delayed_49__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_50__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_49__127_, chained_data_delayed_49__126_, chained_data_delayed_49__125_, chained_data_delayed_49__124_, chained_data_delayed_49__123_, chained_data_delayed_49__122_, chained_data_delayed_49__121_, chained_data_delayed_49__120_, chained_data_delayed_49__119_, chained_data_delayed_49__118_, chained_data_delayed_49__117_, chained_data_delayed_49__116_, chained_data_delayed_49__115_, chained_data_delayed_49__114_, chained_data_delayed_49__113_, chained_data_delayed_49__112_, chained_data_delayed_49__111_, chained_data_delayed_49__110_, chained_data_delayed_49__109_, chained_data_delayed_49__108_, chained_data_delayed_49__107_, chained_data_delayed_49__106_, chained_data_delayed_49__105_, chained_data_delayed_49__104_, chained_data_delayed_49__103_, chained_data_delayed_49__102_, chained_data_delayed_49__101_, chained_data_delayed_49__100_, chained_data_delayed_49__99_, chained_data_delayed_49__98_, chained_data_delayed_49__97_, chained_data_delayed_49__96_, chained_data_delayed_49__95_, chained_data_delayed_49__94_, chained_data_delayed_49__93_, chained_data_delayed_49__92_, chained_data_delayed_49__91_, chained_data_delayed_49__90_, chained_data_delayed_49__89_, chained_data_delayed_49__88_, chained_data_delayed_49__87_, chained_data_delayed_49__86_, chained_data_delayed_49__85_, chained_data_delayed_49__84_, chained_data_delayed_49__83_, chained_data_delayed_49__82_, chained_data_delayed_49__81_, chained_data_delayed_49__80_, chained_data_delayed_49__79_, chained_data_delayed_49__78_, chained_data_delayed_49__77_, chained_data_delayed_49__76_, chained_data_delayed_49__75_, chained_data_delayed_49__74_, chained_data_delayed_49__73_, chained_data_delayed_49__72_, chained_data_delayed_49__71_, chained_data_delayed_49__70_, chained_data_delayed_49__69_, chained_data_delayed_49__68_, chained_data_delayed_49__67_, chained_data_delayed_49__66_, chained_data_delayed_49__65_, chained_data_delayed_49__64_, chained_data_delayed_49__63_, chained_data_delayed_49__62_, chained_data_delayed_49__61_, chained_data_delayed_49__60_, chained_data_delayed_49__59_, chained_data_delayed_49__58_, chained_data_delayed_49__57_, chained_data_delayed_49__56_, chained_data_delayed_49__55_, chained_data_delayed_49__54_, chained_data_delayed_49__53_, chained_data_delayed_49__52_, chained_data_delayed_49__51_, chained_data_delayed_49__50_, chained_data_delayed_49__49_, chained_data_delayed_49__48_, chained_data_delayed_49__47_, chained_data_delayed_49__46_, chained_data_delayed_49__45_, chained_data_delayed_49__44_, chained_data_delayed_49__43_, chained_data_delayed_49__42_, chained_data_delayed_49__41_, chained_data_delayed_49__40_, chained_data_delayed_49__39_, chained_data_delayed_49__38_, chained_data_delayed_49__37_, chained_data_delayed_49__36_, chained_data_delayed_49__35_, chained_data_delayed_49__34_, chained_data_delayed_49__33_, chained_data_delayed_49__32_, chained_data_delayed_49__31_, chained_data_delayed_49__30_, chained_data_delayed_49__29_, chained_data_delayed_49__28_, chained_data_delayed_49__27_, chained_data_delayed_49__26_, chained_data_delayed_49__25_, chained_data_delayed_49__24_, chained_data_delayed_49__23_, chained_data_delayed_49__22_, chained_data_delayed_49__21_, chained_data_delayed_49__20_, chained_data_delayed_49__19_, chained_data_delayed_49__18_, chained_data_delayed_49__17_, chained_data_delayed_49__16_, chained_data_delayed_49__15_, chained_data_delayed_49__14_, chained_data_delayed_49__13_, chained_data_delayed_49__12_, chained_data_delayed_49__11_, chained_data_delayed_49__10_, chained_data_delayed_49__9_, chained_data_delayed_49__8_, chained_data_delayed_49__7_, chained_data_delayed_49__6_, chained_data_delayed_49__5_, chained_data_delayed_49__4_, chained_data_delayed_49__3_, chained_data_delayed_49__2_, chained_data_delayed_49__1_, chained_data_delayed_49__0_ }),
    .data_o({ chained_data_delayed_50__127_, chained_data_delayed_50__126_, chained_data_delayed_50__125_, chained_data_delayed_50__124_, chained_data_delayed_50__123_, chained_data_delayed_50__122_, chained_data_delayed_50__121_, chained_data_delayed_50__120_, chained_data_delayed_50__119_, chained_data_delayed_50__118_, chained_data_delayed_50__117_, chained_data_delayed_50__116_, chained_data_delayed_50__115_, chained_data_delayed_50__114_, chained_data_delayed_50__113_, chained_data_delayed_50__112_, chained_data_delayed_50__111_, chained_data_delayed_50__110_, chained_data_delayed_50__109_, chained_data_delayed_50__108_, chained_data_delayed_50__107_, chained_data_delayed_50__106_, chained_data_delayed_50__105_, chained_data_delayed_50__104_, chained_data_delayed_50__103_, chained_data_delayed_50__102_, chained_data_delayed_50__101_, chained_data_delayed_50__100_, chained_data_delayed_50__99_, chained_data_delayed_50__98_, chained_data_delayed_50__97_, chained_data_delayed_50__96_, chained_data_delayed_50__95_, chained_data_delayed_50__94_, chained_data_delayed_50__93_, chained_data_delayed_50__92_, chained_data_delayed_50__91_, chained_data_delayed_50__90_, chained_data_delayed_50__89_, chained_data_delayed_50__88_, chained_data_delayed_50__87_, chained_data_delayed_50__86_, chained_data_delayed_50__85_, chained_data_delayed_50__84_, chained_data_delayed_50__83_, chained_data_delayed_50__82_, chained_data_delayed_50__81_, chained_data_delayed_50__80_, chained_data_delayed_50__79_, chained_data_delayed_50__78_, chained_data_delayed_50__77_, chained_data_delayed_50__76_, chained_data_delayed_50__75_, chained_data_delayed_50__74_, chained_data_delayed_50__73_, chained_data_delayed_50__72_, chained_data_delayed_50__71_, chained_data_delayed_50__70_, chained_data_delayed_50__69_, chained_data_delayed_50__68_, chained_data_delayed_50__67_, chained_data_delayed_50__66_, chained_data_delayed_50__65_, chained_data_delayed_50__64_, chained_data_delayed_50__63_, chained_data_delayed_50__62_, chained_data_delayed_50__61_, chained_data_delayed_50__60_, chained_data_delayed_50__59_, chained_data_delayed_50__58_, chained_data_delayed_50__57_, chained_data_delayed_50__56_, chained_data_delayed_50__55_, chained_data_delayed_50__54_, chained_data_delayed_50__53_, chained_data_delayed_50__52_, chained_data_delayed_50__51_, chained_data_delayed_50__50_, chained_data_delayed_50__49_, chained_data_delayed_50__48_, chained_data_delayed_50__47_, chained_data_delayed_50__46_, chained_data_delayed_50__45_, chained_data_delayed_50__44_, chained_data_delayed_50__43_, chained_data_delayed_50__42_, chained_data_delayed_50__41_, chained_data_delayed_50__40_, chained_data_delayed_50__39_, chained_data_delayed_50__38_, chained_data_delayed_50__37_, chained_data_delayed_50__36_, chained_data_delayed_50__35_, chained_data_delayed_50__34_, chained_data_delayed_50__33_, chained_data_delayed_50__32_, chained_data_delayed_50__31_, chained_data_delayed_50__30_, chained_data_delayed_50__29_, chained_data_delayed_50__28_, chained_data_delayed_50__27_, chained_data_delayed_50__26_, chained_data_delayed_50__25_, chained_data_delayed_50__24_, chained_data_delayed_50__23_, chained_data_delayed_50__22_, chained_data_delayed_50__21_, chained_data_delayed_50__20_, chained_data_delayed_50__19_, chained_data_delayed_50__18_, chained_data_delayed_50__17_, chained_data_delayed_50__16_, chained_data_delayed_50__15_, chained_data_delayed_50__14_, chained_data_delayed_50__13_, chained_data_delayed_50__12_, chained_data_delayed_50__11_, chained_data_delayed_50__10_, chained_data_delayed_50__9_, chained_data_delayed_50__8_, chained_data_delayed_50__7_, chained_data_delayed_50__6_, chained_data_delayed_50__5_, chained_data_delayed_50__4_, chained_data_delayed_50__3_, chained_data_delayed_50__2_, chained_data_delayed_50__1_, chained_data_delayed_50__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_51__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_50__127_, chained_data_delayed_50__126_, chained_data_delayed_50__125_, chained_data_delayed_50__124_, chained_data_delayed_50__123_, chained_data_delayed_50__122_, chained_data_delayed_50__121_, chained_data_delayed_50__120_, chained_data_delayed_50__119_, chained_data_delayed_50__118_, chained_data_delayed_50__117_, chained_data_delayed_50__116_, chained_data_delayed_50__115_, chained_data_delayed_50__114_, chained_data_delayed_50__113_, chained_data_delayed_50__112_, chained_data_delayed_50__111_, chained_data_delayed_50__110_, chained_data_delayed_50__109_, chained_data_delayed_50__108_, chained_data_delayed_50__107_, chained_data_delayed_50__106_, chained_data_delayed_50__105_, chained_data_delayed_50__104_, chained_data_delayed_50__103_, chained_data_delayed_50__102_, chained_data_delayed_50__101_, chained_data_delayed_50__100_, chained_data_delayed_50__99_, chained_data_delayed_50__98_, chained_data_delayed_50__97_, chained_data_delayed_50__96_, chained_data_delayed_50__95_, chained_data_delayed_50__94_, chained_data_delayed_50__93_, chained_data_delayed_50__92_, chained_data_delayed_50__91_, chained_data_delayed_50__90_, chained_data_delayed_50__89_, chained_data_delayed_50__88_, chained_data_delayed_50__87_, chained_data_delayed_50__86_, chained_data_delayed_50__85_, chained_data_delayed_50__84_, chained_data_delayed_50__83_, chained_data_delayed_50__82_, chained_data_delayed_50__81_, chained_data_delayed_50__80_, chained_data_delayed_50__79_, chained_data_delayed_50__78_, chained_data_delayed_50__77_, chained_data_delayed_50__76_, chained_data_delayed_50__75_, chained_data_delayed_50__74_, chained_data_delayed_50__73_, chained_data_delayed_50__72_, chained_data_delayed_50__71_, chained_data_delayed_50__70_, chained_data_delayed_50__69_, chained_data_delayed_50__68_, chained_data_delayed_50__67_, chained_data_delayed_50__66_, chained_data_delayed_50__65_, chained_data_delayed_50__64_, chained_data_delayed_50__63_, chained_data_delayed_50__62_, chained_data_delayed_50__61_, chained_data_delayed_50__60_, chained_data_delayed_50__59_, chained_data_delayed_50__58_, chained_data_delayed_50__57_, chained_data_delayed_50__56_, chained_data_delayed_50__55_, chained_data_delayed_50__54_, chained_data_delayed_50__53_, chained_data_delayed_50__52_, chained_data_delayed_50__51_, chained_data_delayed_50__50_, chained_data_delayed_50__49_, chained_data_delayed_50__48_, chained_data_delayed_50__47_, chained_data_delayed_50__46_, chained_data_delayed_50__45_, chained_data_delayed_50__44_, chained_data_delayed_50__43_, chained_data_delayed_50__42_, chained_data_delayed_50__41_, chained_data_delayed_50__40_, chained_data_delayed_50__39_, chained_data_delayed_50__38_, chained_data_delayed_50__37_, chained_data_delayed_50__36_, chained_data_delayed_50__35_, chained_data_delayed_50__34_, chained_data_delayed_50__33_, chained_data_delayed_50__32_, chained_data_delayed_50__31_, chained_data_delayed_50__30_, chained_data_delayed_50__29_, chained_data_delayed_50__28_, chained_data_delayed_50__27_, chained_data_delayed_50__26_, chained_data_delayed_50__25_, chained_data_delayed_50__24_, chained_data_delayed_50__23_, chained_data_delayed_50__22_, chained_data_delayed_50__21_, chained_data_delayed_50__20_, chained_data_delayed_50__19_, chained_data_delayed_50__18_, chained_data_delayed_50__17_, chained_data_delayed_50__16_, chained_data_delayed_50__15_, chained_data_delayed_50__14_, chained_data_delayed_50__13_, chained_data_delayed_50__12_, chained_data_delayed_50__11_, chained_data_delayed_50__10_, chained_data_delayed_50__9_, chained_data_delayed_50__8_, chained_data_delayed_50__7_, chained_data_delayed_50__6_, chained_data_delayed_50__5_, chained_data_delayed_50__4_, chained_data_delayed_50__3_, chained_data_delayed_50__2_, chained_data_delayed_50__1_, chained_data_delayed_50__0_ }),
    .data_o({ chained_data_delayed_51__127_, chained_data_delayed_51__126_, chained_data_delayed_51__125_, chained_data_delayed_51__124_, chained_data_delayed_51__123_, chained_data_delayed_51__122_, chained_data_delayed_51__121_, chained_data_delayed_51__120_, chained_data_delayed_51__119_, chained_data_delayed_51__118_, chained_data_delayed_51__117_, chained_data_delayed_51__116_, chained_data_delayed_51__115_, chained_data_delayed_51__114_, chained_data_delayed_51__113_, chained_data_delayed_51__112_, chained_data_delayed_51__111_, chained_data_delayed_51__110_, chained_data_delayed_51__109_, chained_data_delayed_51__108_, chained_data_delayed_51__107_, chained_data_delayed_51__106_, chained_data_delayed_51__105_, chained_data_delayed_51__104_, chained_data_delayed_51__103_, chained_data_delayed_51__102_, chained_data_delayed_51__101_, chained_data_delayed_51__100_, chained_data_delayed_51__99_, chained_data_delayed_51__98_, chained_data_delayed_51__97_, chained_data_delayed_51__96_, chained_data_delayed_51__95_, chained_data_delayed_51__94_, chained_data_delayed_51__93_, chained_data_delayed_51__92_, chained_data_delayed_51__91_, chained_data_delayed_51__90_, chained_data_delayed_51__89_, chained_data_delayed_51__88_, chained_data_delayed_51__87_, chained_data_delayed_51__86_, chained_data_delayed_51__85_, chained_data_delayed_51__84_, chained_data_delayed_51__83_, chained_data_delayed_51__82_, chained_data_delayed_51__81_, chained_data_delayed_51__80_, chained_data_delayed_51__79_, chained_data_delayed_51__78_, chained_data_delayed_51__77_, chained_data_delayed_51__76_, chained_data_delayed_51__75_, chained_data_delayed_51__74_, chained_data_delayed_51__73_, chained_data_delayed_51__72_, chained_data_delayed_51__71_, chained_data_delayed_51__70_, chained_data_delayed_51__69_, chained_data_delayed_51__68_, chained_data_delayed_51__67_, chained_data_delayed_51__66_, chained_data_delayed_51__65_, chained_data_delayed_51__64_, chained_data_delayed_51__63_, chained_data_delayed_51__62_, chained_data_delayed_51__61_, chained_data_delayed_51__60_, chained_data_delayed_51__59_, chained_data_delayed_51__58_, chained_data_delayed_51__57_, chained_data_delayed_51__56_, chained_data_delayed_51__55_, chained_data_delayed_51__54_, chained_data_delayed_51__53_, chained_data_delayed_51__52_, chained_data_delayed_51__51_, chained_data_delayed_51__50_, chained_data_delayed_51__49_, chained_data_delayed_51__48_, chained_data_delayed_51__47_, chained_data_delayed_51__46_, chained_data_delayed_51__45_, chained_data_delayed_51__44_, chained_data_delayed_51__43_, chained_data_delayed_51__42_, chained_data_delayed_51__41_, chained_data_delayed_51__40_, chained_data_delayed_51__39_, chained_data_delayed_51__38_, chained_data_delayed_51__37_, chained_data_delayed_51__36_, chained_data_delayed_51__35_, chained_data_delayed_51__34_, chained_data_delayed_51__33_, chained_data_delayed_51__32_, chained_data_delayed_51__31_, chained_data_delayed_51__30_, chained_data_delayed_51__29_, chained_data_delayed_51__28_, chained_data_delayed_51__27_, chained_data_delayed_51__26_, chained_data_delayed_51__25_, chained_data_delayed_51__24_, chained_data_delayed_51__23_, chained_data_delayed_51__22_, chained_data_delayed_51__21_, chained_data_delayed_51__20_, chained_data_delayed_51__19_, chained_data_delayed_51__18_, chained_data_delayed_51__17_, chained_data_delayed_51__16_, chained_data_delayed_51__15_, chained_data_delayed_51__14_, chained_data_delayed_51__13_, chained_data_delayed_51__12_, chained_data_delayed_51__11_, chained_data_delayed_51__10_, chained_data_delayed_51__9_, chained_data_delayed_51__8_, chained_data_delayed_51__7_, chained_data_delayed_51__6_, chained_data_delayed_51__5_, chained_data_delayed_51__4_, chained_data_delayed_51__3_, chained_data_delayed_51__2_, chained_data_delayed_51__1_, chained_data_delayed_51__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_52__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_51__127_, chained_data_delayed_51__126_, chained_data_delayed_51__125_, chained_data_delayed_51__124_, chained_data_delayed_51__123_, chained_data_delayed_51__122_, chained_data_delayed_51__121_, chained_data_delayed_51__120_, chained_data_delayed_51__119_, chained_data_delayed_51__118_, chained_data_delayed_51__117_, chained_data_delayed_51__116_, chained_data_delayed_51__115_, chained_data_delayed_51__114_, chained_data_delayed_51__113_, chained_data_delayed_51__112_, chained_data_delayed_51__111_, chained_data_delayed_51__110_, chained_data_delayed_51__109_, chained_data_delayed_51__108_, chained_data_delayed_51__107_, chained_data_delayed_51__106_, chained_data_delayed_51__105_, chained_data_delayed_51__104_, chained_data_delayed_51__103_, chained_data_delayed_51__102_, chained_data_delayed_51__101_, chained_data_delayed_51__100_, chained_data_delayed_51__99_, chained_data_delayed_51__98_, chained_data_delayed_51__97_, chained_data_delayed_51__96_, chained_data_delayed_51__95_, chained_data_delayed_51__94_, chained_data_delayed_51__93_, chained_data_delayed_51__92_, chained_data_delayed_51__91_, chained_data_delayed_51__90_, chained_data_delayed_51__89_, chained_data_delayed_51__88_, chained_data_delayed_51__87_, chained_data_delayed_51__86_, chained_data_delayed_51__85_, chained_data_delayed_51__84_, chained_data_delayed_51__83_, chained_data_delayed_51__82_, chained_data_delayed_51__81_, chained_data_delayed_51__80_, chained_data_delayed_51__79_, chained_data_delayed_51__78_, chained_data_delayed_51__77_, chained_data_delayed_51__76_, chained_data_delayed_51__75_, chained_data_delayed_51__74_, chained_data_delayed_51__73_, chained_data_delayed_51__72_, chained_data_delayed_51__71_, chained_data_delayed_51__70_, chained_data_delayed_51__69_, chained_data_delayed_51__68_, chained_data_delayed_51__67_, chained_data_delayed_51__66_, chained_data_delayed_51__65_, chained_data_delayed_51__64_, chained_data_delayed_51__63_, chained_data_delayed_51__62_, chained_data_delayed_51__61_, chained_data_delayed_51__60_, chained_data_delayed_51__59_, chained_data_delayed_51__58_, chained_data_delayed_51__57_, chained_data_delayed_51__56_, chained_data_delayed_51__55_, chained_data_delayed_51__54_, chained_data_delayed_51__53_, chained_data_delayed_51__52_, chained_data_delayed_51__51_, chained_data_delayed_51__50_, chained_data_delayed_51__49_, chained_data_delayed_51__48_, chained_data_delayed_51__47_, chained_data_delayed_51__46_, chained_data_delayed_51__45_, chained_data_delayed_51__44_, chained_data_delayed_51__43_, chained_data_delayed_51__42_, chained_data_delayed_51__41_, chained_data_delayed_51__40_, chained_data_delayed_51__39_, chained_data_delayed_51__38_, chained_data_delayed_51__37_, chained_data_delayed_51__36_, chained_data_delayed_51__35_, chained_data_delayed_51__34_, chained_data_delayed_51__33_, chained_data_delayed_51__32_, chained_data_delayed_51__31_, chained_data_delayed_51__30_, chained_data_delayed_51__29_, chained_data_delayed_51__28_, chained_data_delayed_51__27_, chained_data_delayed_51__26_, chained_data_delayed_51__25_, chained_data_delayed_51__24_, chained_data_delayed_51__23_, chained_data_delayed_51__22_, chained_data_delayed_51__21_, chained_data_delayed_51__20_, chained_data_delayed_51__19_, chained_data_delayed_51__18_, chained_data_delayed_51__17_, chained_data_delayed_51__16_, chained_data_delayed_51__15_, chained_data_delayed_51__14_, chained_data_delayed_51__13_, chained_data_delayed_51__12_, chained_data_delayed_51__11_, chained_data_delayed_51__10_, chained_data_delayed_51__9_, chained_data_delayed_51__8_, chained_data_delayed_51__7_, chained_data_delayed_51__6_, chained_data_delayed_51__5_, chained_data_delayed_51__4_, chained_data_delayed_51__3_, chained_data_delayed_51__2_, chained_data_delayed_51__1_, chained_data_delayed_51__0_ }),
    .data_o({ chained_data_delayed_52__127_, chained_data_delayed_52__126_, chained_data_delayed_52__125_, chained_data_delayed_52__124_, chained_data_delayed_52__123_, chained_data_delayed_52__122_, chained_data_delayed_52__121_, chained_data_delayed_52__120_, chained_data_delayed_52__119_, chained_data_delayed_52__118_, chained_data_delayed_52__117_, chained_data_delayed_52__116_, chained_data_delayed_52__115_, chained_data_delayed_52__114_, chained_data_delayed_52__113_, chained_data_delayed_52__112_, chained_data_delayed_52__111_, chained_data_delayed_52__110_, chained_data_delayed_52__109_, chained_data_delayed_52__108_, chained_data_delayed_52__107_, chained_data_delayed_52__106_, chained_data_delayed_52__105_, chained_data_delayed_52__104_, chained_data_delayed_52__103_, chained_data_delayed_52__102_, chained_data_delayed_52__101_, chained_data_delayed_52__100_, chained_data_delayed_52__99_, chained_data_delayed_52__98_, chained_data_delayed_52__97_, chained_data_delayed_52__96_, chained_data_delayed_52__95_, chained_data_delayed_52__94_, chained_data_delayed_52__93_, chained_data_delayed_52__92_, chained_data_delayed_52__91_, chained_data_delayed_52__90_, chained_data_delayed_52__89_, chained_data_delayed_52__88_, chained_data_delayed_52__87_, chained_data_delayed_52__86_, chained_data_delayed_52__85_, chained_data_delayed_52__84_, chained_data_delayed_52__83_, chained_data_delayed_52__82_, chained_data_delayed_52__81_, chained_data_delayed_52__80_, chained_data_delayed_52__79_, chained_data_delayed_52__78_, chained_data_delayed_52__77_, chained_data_delayed_52__76_, chained_data_delayed_52__75_, chained_data_delayed_52__74_, chained_data_delayed_52__73_, chained_data_delayed_52__72_, chained_data_delayed_52__71_, chained_data_delayed_52__70_, chained_data_delayed_52__69_, chained_data_delayed_52__68_, chained_data_delayed_52__67_, chained_data_delayed_52__66_, chained_data_delayed_52__65_, chained_data_delayed_52__64_, chained_data_delayed_52__63_, chained_data_delayed_52__62_, chained_data_delayed_52__61_, chained_data_delayed_52__60_, chained_data_delayed_52__59_, chained_data_delayed_52__58_, chained_data_delayed_52__57_, chained_data_delayed_52__56_, chained_data_delayed_52__55_, chained_data_delayed_52__54_, chained_data_delayed_52__53_, chained_data_delayed_52__52_, chained_data_delayed_52__51_, chained_data_delayed_52__50_, chained_data_delayed_52__49_, chained_data_delayed_52__48_, chained_data_delayed_52__47_, chained_data_delayed_52__46_, chained_data_delayed_52__45_, chained_data_delayed_52__44_, chained_data_delayed_52__43_, chained_data_delayed_52__42_, chained_data_delayed_52__41_, chained_data_delayed_52__40_, chained_data_delayed_52__39_, chained_data_delayed_52__38_, chained_data_delayed_52__37_, chained_data_delayed_52__36_, chained_data_delayed_52__35_, chained_data_delayed_52__34_, chained_data_delayed_52__33_, chained_data_delayed_52__32_, chained_data_delayed_52__31_, chained_data_delayed_52__30_, chained_data_delayed_52__29_, chained_data_delayed_52__28_, chained_data_delayed_52__27_, chained_data_delayed_52__26_, chained_data_delayed_52__25_, chained_data_delayed_52__24_, chained_data_delayed_52__23_, chained_data_delayed_52__22_, chained_data_delayed_52__21_, chained_data_delayed_52__20_, chained_data_delayed_52__19_, chained_data_delayed_52__18_, chained_data_delayed_52__17_, chained_data_delayed_52__16_, chained_data_delayed_52__15_, chained_data_delayed_52__14_, chained_data_delayed_52__13_, chained_data_delayed_52__12_, chained_data_delayed_52__11_, chained_data_delayed_52__10_, chained_data_delayed_52__9_, chained_data_delayed_52__8_, chained_data_delayed_52__7_, chained_data_delayed_52__6_, chained_data_delayed_52__5_, chained_data_delayed_52__4_, chained_data_delayed_52__3_, chained_data_delayed_52__2_, chained_data_delayed_52__1_, chained_data_delayed_52__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_53__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_52__127_, chained_data_delayed_52__126_, chained_data_delayed_52__125_, chained_data_delayed_52__124_, chained_data_delayed_52__123_, chained_data_delayed_52__122_, chained_data_delayed_52__121_, chained_data_delayed_52__120_, chained_data_delayed_52__119_, chained_data_delayed_52__118_, chained_data_delayed_52__117_, chained_data_delayed_52__116_, chained_data_delayed_52__115_, chained_data_delayed_52__114_, chained_data_delayed_52__113_, chained_data_delayed_52__112_, chained_data_delayed_52__111_, chained_data_delayed_52__110_, chained_data_delayed_52__109_, chained_data_delayed_52__108_, chained_data_delayed_52__107_, chained_data_delayed_52__106_, chained_data_delayed_52__105_, chained_data_delayed_52__104_, chained_data_delayed_52__103_, chained_data_delayed_52__102_, chained_data_delayed_52__101_, chained_data_delayed_52__100_, chained_data_delayed_52__99_, chained_data_delayed_52__98_, chained_data_delayed_52__97_, chained_data_delayed_52__96_, chained_data_delayed_52__95_, chained_data_delayed_52__94_, chained_data_delayed_52__93_, chained_data_delayed_52__92_, chained_data_delayed_52__91_, chained_data_delayed_52__90_, chained_data_delayed_52__89_, chained_data_delayed_52__88_, chained_data_delayed_52__87_, chained_data_delayed_52__86_, chained_data_delayed_52__85_, chained_data_delayed_52__84_, chained_data_delayed_52__83_, chained_data_delayed_52__82_, chained_data_delayed_52__81_, chained_data_delayed_52__80_, chained_data_delayed_52__79_, chained_data_delayed_52__78_, chained_data_delayed_52__77_, chained_data_delayed_52__76_, chained_data_delayed_52__75_, chained_data_delayed_52__74_, chained_data_delayed_52__73_, chained_data_delayed_52__72_, chained_data_delayed_52__71_, chained_data_delayed_52__70_, chained_data_delayed_52__69_, chained_data_delayed_52__68_, chained_data_delayed_52__67_, chained_data_delayed_52__66_, chained_data_delayed_52__65_, chained_data_delayed_52__64_, chained_data_delayed_52__63_, chained_data_delayed_52__62_, chained_data_delayed_52__61_, chained_data_delayed_52__60_, chained_data_delayed_52__59_, chained_data_delayed_52__58_, chained_data_delayed_52__57_, chained_data_delayed_52__56_, chained_data_delayed_52__55_, chained_data_delayed_52__54_, chained_data_delayed_52__53_, chained_data_delayed_52__52_, chained_data_delayed_52__51_, chained_data_delayed_52__50_, chained_data_delayed_52__49_, chained_data_delayed_52__48_, chained_data_delayed_52__47_, chained_data_delayed_52__46_, chained_data_delayed_52__45_, chained_data_delayed_52__44_, chained_data_delayed_52__43_, chained_data_delayed_52__42_, chained_data_delayed_52__41_, chained_data_delayed_52__40_, chained_data_delayed_52__39_, chained_data_delayed_52__38_, chained_data_delayed_52__37_, chained_data_delayed_52__36_, chained_data_delayed_52__35_, chained_data_delayed_52__34_, chained_data_delayed_52__33_, chained_data_delayed_52__32_, chained_data_delayed_52__31_, chained_data_delayed_52__30_, chained_data_delayed_52__29_, chained_data_delayed_52__28_, chained_data_delayed_52__27_, chained_data_delayed_52__26_, chained_data_delayed_52__25_, chained_data_delayed_52__24_, chained_data_delayed_52__23_, chained_data_delayed_52__22_, chained_data_delayed_52__21_, chained_data_delayed_52__20_, chained_data_delayed_52__19_, chained_data_delayed_52__18_, chained_data_delayed_52__17_, chained_data_delayed_52__16_, chained_data_delayed_52__15_, chained_data_delayed_52__14_, chained_data_delayed_52__13_, chained_data_delayed_52__12_, chained_data_delayed_52__11_, chained_data_delayed_52__10_, chained_data_delayed_52__9_, chained_data_delayed_52__8_, chained_data_delayed_52__7_, chained_data_delayed_52__6_, chained_data_delayed_52__5_, chained_data_delayed_52__4_, chained_data_delayed_52__3_, chained_data_delayed_52__2_, chained_data_delayed_52__1_, chained_data_delayed_52__0_ }),
    .data_o({ chained_data_delayed_53__127_, chained_data_delayed_53__126_, chained_data_delayed_53__125_, chained_data_delayed_53__124_, chained_data_delayed_53__123_, chained_data_delayed_53__122_, chained_data_delayed_53__121_, chained_data_delayed_53__120_, chained_data_delayed_53__119_, chained_data_delayed_53__118_, chained_data_delayed_53__117_, chained_data_delayed_53__116_, chained_data_delayed_53__115_, chained_data_delayed_53__114_, chained_data_delayed_53__113_, chained_data_delayed_53__112_, chained_data_delayed_53__111_, chained_data_delayed_53__110_, chained_data_delayed_53__109_, chained_data_delayed_53__108_, chained_data_delayed_53__107_, chained_data_delayed_53__106_, chained_data_delayed_53__105_, chained_data_delayed_53__104_, chained_data_delayed_53__103_, chained_data_delayed_53__102_, chained_data_delayed_53__101_, chained_data_delayed_53__100_, chained_data_delayed_53__99_, chained_data_delayed_53__98_, chained_data_delayed_53__97_, chained_data_delayed_53__96_, chained_data_delayed_53__95_, chained_data_delayed_53__94_, chained_data_delayed_53__93_, chained_data_delayed_53__92_, chained_data_delayed_53__91_, chained_data_delayed_53__90_, chained_data_delayed_53__89_, chained_data_delayed_53__88_, chained_data_delayed_53__87_, chained_data_delayed_53__86_, chained_data_delayed_53__85_, chained_data_delayed_53__84_, chained_data_delayed_53__83_, chained_data_delayed_53__82_, chained_data_delayed_53__81_, chained_data_delayed_53__80_, chained_data_delayed_53__79_, chained_data_delayed_53__78_, chained_data_delayed_53__77_, chained_data_delayed_53__76_, chained_data_delayed_53__75_, chained_data_delayed_53__74_, chained_data_delayed_53__73_, chained_data_delayed_53__72_, chained_data_delayed_53__71_, chained_data_delayed_53__70_, chained_data_delayed_53__69_, chained_data_delayed_53__68_, chained_data_delayed_53__67_, chained_data_delayed_53__66_, chained_data_delayed_53__65_, chained_data_delayed_53__64_, chained_data_delayed_53__63_, chained_data_delayed_53__62_, chained_data_delayed_53__61_, chained_data_delayed_53__60_, chained_data_delayed_53__59_, chained_data_delayed_53__58_, chained_data_delayed_53__57_, chained_data_delayed_53__56_, chained_data_delayed_53__55_, chained_data_delayed_53__54_, chained_data_delayed_53__53_, chained_data_delayed_53__52_, chained_data_delayed_53__51_, chained_data_delayed_53__50_, chained_data_delayed_53__49_, chained_data_delayed_53__48_, chained_data_delayed_53__47_, chained_data_delayed_53__46_, chained_data_delayed_53__45_, chained_data_delayed_53__44_, chained_data_delayed_53__43_, chained_data_delayed_53__42_, chained_data_delayed_53__41_, chained_data_delayed_53__40_, chained_data_delayed_53__39_, chained_data_delayed_53__38_, chained_data_delayed_53__37_, chained_data_delayed_53__36_, chained_data_delayed_53__35_, chained_data_delayed_53__34_, chained_data_delayed_53__33_, chained_data_delayed_53__32_, chained_data_delayed_53__31_, chained_data_delayed_53__30_, chained_data_delayed_53__29_, chained_data_delayed_53__28_, chained_data_delayed_53__27_, chained_data_delayed_53__26_, chained_data_delayed_53__25_, chained_data_delayed_53__24_, chained_data_delayed_53__23_, chained_data_delayed_53__22_, chained_data_delayed_53__21_, chained_data_delayed_53__20_, chained_data_delayed_53__19_, chained_data_delayed_53__18_, chained_data_delayed_53__17_, chained_data_delayed_53__16_, chained_data_delayed_53__15_, chained_data_delayed_53__14_, chained_data_delayed_53__13_, chained_data_delayed_53__12_, chained_data_delayed_53__11_, chained_data_delayed_53__10_, chained_data_delayed_53__9_, chained_data_delayed_53__8_, chained_data_delayed_53__7_, chained_data_delayed_53__6_, chained_data_delayed_53__5_, chained_data_delayed_53__4_, chained_data_delayed_53__3_, chained_data_delayed_53__2_, chained_data_delayed_53__1_, chained_data_delayed_53__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_54__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_53__127_, chained_data_delayed_53__126_, chained_data_delayed_53__125_, chained_data_delayed_53__124_, chained_data_delayed_53__123_, chained_data_delayed_53__122_, chained_data_delayed_53__121_, chained_data_delayed_53__120_, chained_data_delayed_53__119_, chained_data_delayed_53__118_, chained_data_delayed_53__117_, chained_data_delayed_53__116_, chained_data_delayed_53__115_, chained_data_delayed_53__114_, chained_data_delayed_53__113_, chained_data_delayed_53__112_, chained_data_delayed_53__111_, chained_data_delayed_53__110_, chained_data_delayed_53__109_, chained_data_delayed_53__108_, chained_data_delayed_53__107_, chained_data_delayed_53__106_, chained_data_delayed_53__105_, chained_data_delayed_53__104_, chained_data_delayed_53__103_, chained_data_delayed_53__102_, chained_data_delayed_53__101_, chained_data_delayed_53__100_, chained_data_delayed_53__99_, chained_data_delayed_53__98_, chained_data_delayed_53__97_, chained_data_delayed_53__96_, chained_data_delayed_53__95_, chained_data_delayed_53__94_, chained_data_delayed_53__93_, chained_data_delayed_53__92_, chained_data_delayed_53__91_, chained_data_delayed_53__90_, chained_data_delayed_53__89_, chained_data_delayed_53__88_, chained_data_delayed_53__87_, chained_data_delayed_53__86_, chained_data_delayed_53__85_, chained_data_delayed_53__84_, chained_data_delayed_53__83_, chained_data_delayed_53__82_, chained_data_delayed_53__81_, chained_data_delayed_53__80_, chained_data_delayed_53__79_, chained_data_delayed_53__78_, chained_data_delayed_53__77_, chained_data_delayed_53__76_, chained_data_delayed_53__75_, chained_data_delayed_53__74_, chained_data_delayed_53__73_, chained_data_delayed_53__72_, chained_data_delayed_53__71_, chained_data_delayed_53__70_, chained_data_delayed_53__69_, chained_data_delayed_53__68_, chained_data_delayed_53__67_, chained_data_delayed_53__66_, chained_data_delayed_53__65_, chained_data_delayed_53__64_, chained_data_delayed_53__63_, chained_data_delayed_53__62_, chained_data_delayed_53__61_, chained_data_delayed_53__60_, chained_data_delayed_53__59_, chained_data_delayed_53__58_, chained_data_delayed_53__57_, chained_data_delayed_53__56_, chained_data_delayed_53__55_, chained_data_delayed_53__54_, chained_data_delayed_53__53_, chained_data_delayed_53__52_, chained_data_delayed_53__51_, chained_data_delayed_53__50_, chained_data_delayed_53__49_, chained_data_delayed_53__48_, chained_data_delayed_53__47_, chained_data_delayed_53__46_, chained_data_delayed_53__45_, chained_data_delayed_53__44_, chained_data_delayed_53__43_, chained_data_delayed_53__42_, chained_data_delayed_53__41_, chained_data_delayed_53__40_, chained_data_delayed_53__39_, chained_data_delayed_53__38_, chained_data_delayed_53__37_, chained_data_delayed_53__36_, chained_data_delayed_53__35_, chained_data_delayed_53__34_, chained_data_delayed_53__33_, chained_data_delayed_53__32_, chained_data_delayed_53__31_, chained_data_delayed_53__30_, chained_data_delayed_53__29_, chained_data_delayed_53__28_, chained_data_delayed_53__27_, chained_data_delayed_53__26_, chained_data_delayed_53__25_, chained_data_delayed_53__24_, chained_data_delayed_53__23_, chained_data_delayed_53__22_, chained_data_delayed_53__21_, chained_data_delayed_53__20_, chained_data_delayed_53__19_, chained_data_delayed_53__18_, chained_data_delayed_53__17_, chained_data_delayed_53__16_, chained_data_delayed_53__15_, chained_data_delayed_53__14_, chained_data_delayed_53__13_, chained_data_delayed_53__12_, chained_data_delayed_53__11_, chained_data_delayed_53__10_, chained_data_delayed_53__9_, chained_data_delayed_53__8_, chained_data_delayed_53__7_, chained_data_delayed_53__6_, chained_data_delayed_53__5_, chained_data_delayed_53__4_, chained_data_delayed_53__3_, chained_data_delayed_53__2_, chained_data_delayed_53__1_, chained_data_delayed_53__0_ }),
    .data_o({ chained_data_delayed_54__127_, chained_data_delayed_54__126_, chained_data_delayed_54__125_, chained_data_delayed_54__124_, chained_data_delayed_54__123_, chained_data_delayed_54__122_, chained_data_delayed_54__121_, chained_data_delayed_54__120_, chained_data_delayed_54__119_, chained_data_delayed_54__118_, chained_data_delayed_54__117_, chained_data_delayed_54__116_, chained_data_delayed_54__115_, chained_data_delayed_54__114_, chained_data_delayed_54__113_, chained_data_delayed_54__112_, chained_data_delayed_54__111_, chained_data_delayed_54__110_, chained_data_delayed_54__109_, chained_data_delayed_54__108_, chained_data_delayed_54__107_, chained_data_delayed_54__106_, chained_data_delayed_54__105_, chained_data_delayed_54__104_, chained_data_delayed_54__103_, chained_data_delayed_54__102_, chained_data_delayed_54__101_, chained_data_delayed_54__100_, chained_data_delayed_54__99_, chained_data_delayed_54__98_, chained_data_delayed_54__97_, chained_data_delayed_54__96_, chained_data_delayed_54__95_, chained_data_delayed_54__94_, chained_data_delayed_54__93_, chained_data_delayed_54__92_, chained_data_delayed_54__91_, chained_data_delayed_54__90_, chained_data_delayed_54__89_, chained_data_delayed_54__88_, chained_data_delayed_54__87_, chained_data_delayed_54__86_, chained_data_delayed_54__85_, chained_data_delayed_54__84_, chained_data_delayed_54__83_, chained_data_delayed_54__82_, chained_data_delayed_54__81_, chained_data_delayed_54__80_, chained_data_delayed_54__79_, chained_data_delayed_54__78_, chained_data_delayed_54__77_, chained_data_delayed_54__76_, chained_data_delayed_54__75_, chained_data_delayed_54__74_, chained_data_delayed_54__73_, chained_data_delayed_54__72_, chained_data_delayed_54__71_, chained_data_delayed_54__70_, chained_data_delayed_54__69_, chained_data_delayed_54__68_, chained_data_delayed_54__67_, chained_data_delayed_54__66_, chained_data_delayed_54__65_, chained_data_delayed_54__64_, chained_data_delayed_54__63_, chained_data_delayed_54__62_, chained_data_delayed_54__61_, chained_data_delayed_54__60_, chained_data_delayed_54__59_, chained_data_delayed_54__58_, chained_data_delayed_54__57_, chained_data_delayed_54__56_, chained_data_delayed_54__55_, chained_data_delayed_54__54_, chained_data_delayed_54__53_, chained_data_delayed_54__52_, chained_data_delayed_54__51_, chained_data_delayed_54__50_, chained_data_delayed_54__49_, chained_data_delayed_54__48_, chained_data_delayed_54__47_, chained_data_delayed_54__46_, chained_data_delayed_54__45_, chained_data_delayed_54__44_, chained_data_delayed_54__43_, chained_data_delayed_54__42_, chained_data_delayed_54__41_, chained_data_delayed_54__40_, chained_data_delayed_54__39_, chained_data_delayed_54__38_, chained_data_delayed_54__37_, chained_data_delayed_54__36_, chained_data_delayed_54__35_, chained_data_delayed_54__34_, chained_data_delayed_54__33_, chained_data_delayed_54__32_, chained_data_delayed_54__31_, chained_data_delayed_54__30_, chained_data_delayed_54__29_, chained_data_delayed_54__28_, chained_data_delayed_54__27_, chained_data_delayed_54__26_, chained_data_delayed_54__25_, chained_data_delayed_54__24_, chained_data_delayed_54__23_, chained_data_delayed_54__22_, chained_data_delayed_54__21_, chained_data_delayed_54__20_, chained_data_delayed_54__19_, chained_data_delayed_54__18_, chained_data_delayed_54__17_, chained_data_delayed_54__16_, chained_data_delayed_54__15_, chained_data_delayed_54__14_, chained_data_delayed_54__13_, chained_data_delayed_54__12_, chained_data_delayed_54__11_, chained_data_delayed_54__10_, chained_data_delayed_54__9_, chained_data_delayed_54__8_, chained_data_delayed_54__7_, chained_data_delayed_54__6_, chained_data_delayed_54__5_, chained_data_delayed_54__4_, chained_data_delayed_54__3_, chained_data_delayed_54__2_, chained_data_delayed_54__1_, chained_data_delayed_54__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_55__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_54__127_, chained_data_delayed_54__126_, chained_data_delayed_54__125_, chained_data_delayed_54__124_, chained_data_delayed_54__123_, chained_data_delayed_54__122_, chained_data_delayed_54__121_, chained_data_delayed_54__120_, chained_data_delayed_54__119_, chained_data_delayed_54__118_, chained_data_delayed_54__117_, chained_data_delayed_54__116_, chained_data_delayed_54__115_, chained_data_delayed_54__114_, chained_data_delayed_54__113_, chained_data_delayed_54__112_, chained_data_delayed_54__111_, chained_data_delayed_54__110_, chained_data_delayed_54__109_, chained_data_delayed_54__108_, chained_data_delayed_54__107_, chained_data_delayed_54__106_, chained_data_delayed_54__105_, chained_data_delayed_54__104_, chained_data_delayed_54__103_, chained_data_delayed_54__102_, chained_data_delayed_54__101_, chained_data_delayed_54__100_, chained_data_delayed_54__99_, chained_data_delayed_54__98_, chained_data_delayed_54__97_, chained_data_delayed_54__96_, chained_data_delayed_54__95_, chained_data_delayed_54__94_, chained_data_delayed_54__93_, chained_data_delayed_54__92_, chained_data_delayed_54__91_, chained_data_delayed_54__90_, chained_data_delayed_54__89_, chained_data_delayed_54__88_, chained_data_delayed_54__87_, chained_data_delayed_54__86_, chained_data_delayed_54__85_, chained_data_delayed_54__84_, chained_data_delayed_54__83_, chained_data_delayed_54__82_, chained_data_delayed_54__81_, chained_data_delayed_54__80_, chained_data_delayed_54__79_, chained_data_delayed_54__78_, chained_data_delayed_54__77_, chained_data_delayed_54__76_, chained_data_delayed_54__75_, chained_data_delayed_54__74_, chained_data_delayed_54__73_, chained_data_delayed_54__72_, chained_data_delayed_54__71_, chained_data_delayed_54__70_, chained_data_delayed_54__69_, chained_data_delayed_54__68_, chained_data_delayed_54__67_, chained_data_delayed_54__66_, chained_data_delayed_54__65_, chained_data_delayed_54__64_, chained_data_delayed_54__63_, chained_data_delayed_54__62_, chained_data_delayed_54__61_, chained_data_delayed_54__60_, chained_data_delayed_54__59_, chained_data_delayed_54__58_, chained_data_delayed_54__57_, chained_data_delayed_54__56_, chained_data_delayed_54__55_, chained_data_delayed_54__54_, chained_data_delayed_54__53_, chained_data_delayed_54__52_, chained_data_delayed_54__51_, chained_data_delayed_54__50_, chained_data_delayed_54__49_, chained_data_delayed_54__48_, chained_data_delayed_54__47_, chained_data_delayed_54__46_, chained_data_delayed_54__45_, chained_data_delayed_54__44_, chained_data_delayed_54__43_, chained_data_delayed_54__42_, chained_data_delayed_54__41_, chained_data_delayed_54__40_, chained_data_delayed_54__39_, chained_data_delayed_54__38_, chained_data_delayed_54__37_, chained_data_delayed_54__36_, chained_data_delayed_54__35_, chained_data_delayed_54__34_, chained_data_delayed_54__33_, chained_data_delayed_54__32_, chained_data_delayed_54__31_, chained_data_delayed_54__30_, chained_data_delayed_54__29_, chained_data_delayed_54__28_, chained_data_delayed_54__27_, chained_data_delayed_54__26_, chained_data_delayed_54__25_, chained_data_delayed_54__24_, chained_data_delayed_54__23_, chained_data_delayed_54__22_, chained_data_delayed_54__21_, chained_data_delayed_54__20_, chained_data_delayed_54__19_, chained_data_delayed_54__18_, chained_data_delayed_54__17_, chained_data_delayed_54__16_, chained_data_delayed_54__15_, chained_data_delayed_54__14_, chained_data_delayed_54__13_, chained_data_delayed_54__12_, chained_data_delayed_54__11_, chained_data_delayed_54__10_, chained_data_delayed_54__9_, chained_data_delayed_54__8_, chained_data_delayed_54__7_, chained_data_delayed_54__6_, chained_data_delayed_54__5_, chained_data_delayed_54__4_, chained_data_delayed_54__3_, chained_data_delayed_54__2_, chained_data_delayed_54__1_, chained_data_delayed_54__0_ }),
    .data_o({ chained_data_delayed_55__127_, chained_data_delayed_55__126_, chained_data_delayed_55__125_, chained_data_delayed_55__124_, chained_data_delayed_55__123_, chained_data_delayed_55__122_, chained_data_delayed_55__121_, chained_data_delayed_55__120_, chained_data_delayed_55__119_, chained_data_delayed_55__118_, chained_data_delayed_55__117_, chained_data_delayed_55__116_, chained_data_delayed_55__115_, chained_data_delayed_55__114_, chained_data_delayed_55__113_, chained_data_delayed_55__112_, chained_data_delayed_55__111_, chained_data_delayed_55__110_, chained_data_delayed_55__109_, chained_data_delayed_55__108_, chained_data_delayed_55__107_, chained_data_delayed_55__106_, chained_data_delayed_55__105_, chained_data_delayed_55__104_, chained_data_delayed_55__103_, chained_data_delayed_55__102_, chained_data_delayed_55__101_, chained_data_delayed_55__100_, chained_data_delayed_55__99_, chained_data_delayed_55__98_, chained_data_delayed_55__97_, chained_data_delayed_55__96_, chained_data_delayed_55__95_, chained_data_delayed_55__94_, chained_data_delayed_55__93_, chained_data_delayed_55__92_, chained_data_delayed_55__91_, chained_data_delayed_55__90_, chained_data_delayed_55__89_, chained_data_delayed_55__88_, chained_data_delayed_55__87_, chained_data_delayed_55__86_, chained_data_delayed_55__85_, chained_data_delayed_55__84_, chained_data_delayed_55__83_, chained_data_delayed_55__82_, chained_data_delayed_55__81_, chained_data_delayed_55__80_, chained_data_delayed_55__79_, chained_data_delayed_55__78_, chained_data_delayed_55__77_, chained_data_delayed_55__76_, chained_data_delayed_55__75_, chained_data_delayed_55__74_, chained_data_delayed_55__73_, chained_data_delayed_55__72_, chained_data_delayed_55__71_, chained_data_delayed_55__70_, chained_data_delayed_55__69_, chained_data_delayed_55__68_, chained_data_delayed_55__67_, chained_data_delayed_55__66_, chained_data_delayed_55__65_, chained_data_delayed_55__64_, chained_data_delayed_55__63_, chained_data_delayed_55__62_, chained_data_delayed_55__61_, chained_data_delayed_55__60_, chained_data_delayed_55__59_, chained_data_delayed_55__58_, chained_data_delayed_55__57_, chained_data_delayed_55__56_, chained_data_delayed_55__55_, chained_data_delayed_55__54_, chained_data_delayed_55__53_, chained_data_delayed_55__52_, chained_data_delayed_55__51_, chained_data_delayed_55__50_, chained_data_delayed_55__49_, chained_data_delayed_55__48_, chained_data_delayed_55__47_, chained_data_delayed_55__46_, chained_data_delayed_55__45_, chained_data_delayed_55__44_, chained_data_delayed_55__43_, chained_data_delayed_55__42_, chained_data_delayed_55__41_, chained_data_delayed_55__40_, chained_data_delayed_55__39_, chained_data_delayed_55__38_, chained_data_delayed_55__37_, chained_data_delayed_55__36_, chained_data_delayed_55__35_, chained_data_delayed_55__34_, chained_data_delayed_55__33_, chained_data_delayed_55__32_, chained_data_delayed_55__31_, chained_data_delayed_55__30_, chained_data_delayed_55__29_, chained_data_delayed_55__28_, chained_data_delayed_55__27_, chained_data_delayed_55__26_, chained_data_delayed_55__25_, chained_data_delayed_55__24_, chained_data_delayed_55__23_, chained_data_delayed_55__22_, chained_data_delayed_55__21_, chained_data_delayed_55__20_, chained_data_delayed_55__19_, chained_data_delayed_55__18_, chained_data_delayed_55__17_, chained_data_delayed_55__16_, chained_data_delayed_55__15_, chained_data_delayed_55__14_, chained_data_delayed_55__13_, chained_data_delayed_55__12_, chained_data_delayed_55__11_, chained_data_delayed_55__10_, chained_data_delayed_55__9_, chained_data_delayed_55__8_, chained_data_delayed_55__7_, chained_data_delayed_55__6_, chained_data_delayed_55__5_, chained_data_delayed_55__4_, chained_data_delayed_55__3_, chained_data_delayed_55__2_, chained_data_delayed_55__1_, chained_data_delayed_55__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_56__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_55__127_, chained_data_delayed_55__126_, chained_data_delayed_55__125_, chained_data_delayed_55__124_, chained_data_delayed_55__123_, chained_data_delayed_55__122_, chained_data_delayed_55__121_, chained_data_delayed_55__120_, chained_data_delayed_55__119_, chained_data_delayed_55__118_, chained_data_delayed_55__117_, chained_data_delayed_55__116_, chained_data_delayed_55__115_, chained_data_delayed_55__114_, chained_data_delayed_55__113_, chained_data_delayed_55__112_, chained_data_delayed_55__111_, chained_data_delayed_55__110_, chained_data_delayed_55__109_, chained_data_delayed_55__108_, chained_data_delayed_55__107_, chained_data_delayed_55__106_, chained_data_delayed_55__105_, chained_data_delayed_55__104_, chained_data_delayed_55__103_, chained_data_delayed_55__102_, chained_data_delayed_55__101_, chained_data_delayed_55__100_, chained_data_delayed_55__99_, chained_data_delayed_55__98_, chained_data_delayed_55__97_, chained_data_delayed_55__96_, chained_data_delayed_55__95_, chained_data_delayed_55__94_, chained_data_delayed_55__93_, chained_data_delayed_55__92_, chained_data_delayed_55__91_, chained_data_delayed_55__90_, chained_data_delayed_55__89_, chained_data_delayed_55__88_, chained_data_delayed_55__87_, chained_data_delayed_55__86_, chained_data_delayed_55__85_, chained_data_delayed_55__84_, chained_data_delayed_55__83_, chained_data_delayed_55__82_, chained_data_delayed_55__81_, chained_data_delayed_55__80_, chained_data_delayed_55__79_, chained_data_delayed_55__78_, chained_data_delayed_55__77_, chained_data_delayed_55__76_, chained_data_delayed_55__75_, chained_data_delayed_55__74_, chained_data_delayed_55__73_, chained_data_delayed_55__72_, chained_data_delayed_55__71_, chained_data_delayed_55__70_, chained_data_delayed_55__69_, chained_data_delayed_55__68_, chained_data_delayed_55__67_, chained_data_delayed_55__66_, chained_data_delayed_55__65_, chained_data_delayed_55__64_, chained_data_delayed_55__63_, chained_data_delayed_55__62_, chained_data_delayed_55__61_, chained_data_delayed_55__60_, chained_data_delayed_55__59_, chained_data_delayed_55__58_, chained_data_delayed_55__57_, chained_data_delayed_55__56_, chained_data_delayed_55__55_, chained_data_delayed_55__54_, chained_data_delayed_55__53_, chained_data_delayed_55__52_, chained_data_delayed_55__51_, chained_data_delayed_55__50_, chained_data_delayed_55__49_, chained_data_delayed_55__48_, chained_data_delayed_55__47_, chained_data_delayed_55__46_, chained_data_delayed_55__45_, chained_data_delayed_55__44_, chained_data_delayed_55__43_, chained_data_delayed_55__42_, chained_data_delayed_55__41_, chained_data_delayed_55__40_, chained_data_delayed_55__39_, chained_data_delayed_55__38_, chained_data_delayed_55__37_, chained_data_delayed_55__36_, chained_data_delayed_55__35_, chained_data_delayed_55__34_, chained_data_delayed_55__33_, chained_data_delayed_55__32_, chained_data_delayed_55__31_, chained_data_delayed_55__30_, chained_data_delayed_55__29_, chained_data_delayed_55__28_, chained_data_delayed_55__27_, chained_data_delayed_55__26_, chained_data_delayed_55__25_, chained_data_delayed_55__24_, chained_data_delayed_55__23_, chained_data_delayed_55__22_, chained_data_delayed_55__21_, chained_data_delayed_55__20_, chained_data_delayed_55__19_, chained_data_delayed_55__18_, chained_data_delayed_55__17_, chained_data_delayed_55__16_, chained_data_delayed_55__15_, chained_data_delayed_55__14_, chained_data_delayed_55__13_, chained_data_delayed_55__12_, chained_data_delayed_55__11_, chained_data_delayed_55__10_, chained_data_delayed_55__9_, chained_data_delayed_55__8_, chained_data_delayed_55__7_, chained_data_delayed_55__6_, chained_data_delayed_55__5_, chained_data_delayed_55__4_, chained_data_delayed_55__3_, chained_data_delayed_55__2_, chained_data_delayed_55__1_, chained_data_delayed_55__0_ }),
    .data_o({ chained_data_delayed_56__127_, chained_data_delayed_56__126_, chained_data_delayed_56__125_, chained_data_delayed_56__124_, chained_data_delayed_56__123_, chained_data_delayed_56__122_, chained_data_delayed_56__121_, chained_data_delayed_56__120_, chained_data_delayed_56__119_, chained_data_delayed_56__118_, chained_data_delayed_56__117_, chained_data_delayed_56__116_, chained_data_delayed_56__115_, chained_data_delayed_56__114_, chained_data_delayed_56__113_, chained_data_delayed_56__112_, chained_data_delayed_56__111_, chained_data_delayed_56__110_, chained_data_delayed_56__109_, chained_data_delayed_56__108_, chained_data_delayed_56__107_, chained_data_delayed_56__106_, chained_data_delayed_56__105_, chained_data_delayed_56__104_, chained_data_delayed_56__103_, chained_data_delayed_56__102_, chained_data_delayed_56__101_, chained_data_delayed_56__100_, chained_data_delayed_56__99_, chained_data_delayed_56__98_, chained_data_delayed_56__97_, chained_data_delayed_56__96_, chained_data_delayed_56__95_, chained_data_delayed_56__94_, chained_data_delayed_56__93_, chained_data_delayed_56__92_, chained_data_delayed_56__91_, chained_data_delayed_56__90_, chained_data_delayed_56__89_, chained_data_delayed_56__88_, chained_data_delayed_56__87_, chained_data_delayed_56__86_, chained_data_delayed_56__85_, chained_data_delayed_56__84_, chained_data_delayed_56__83_, chained_data_delayed_56__82_, chained_data_delayed_56__81_, chained_data_delayed_56__80_, chained_data_delayed_56__79_, chained_data_delayed_56__78_, chained_data_delayed_56__77_, chained_data_delayed_56__76_, chained_data_delayed_56__75_, chained_data_delayed_56__74_, chained_data_delayed_56__73_, chained_data_delayed_56__72_, chained_data_delayed_56__71_, chained_data_delayed_56__70_, chained_data_delayed_56__69_, chained_data_delayed_56__68_, chained_data_delayed_56__67_, chained_data_delayed_56__66_, chained_data_delayed_56__65_, chained_data_delayed_56__64_, chained_data_delayed_56__63_, chained_data_delayed_56__62_, chained_data_delayed_56__61_, chained_data_delayed_56__60_, chained_data_delayed_56__59_, chained_data_delayed_56__58_, chained_data_delayed_56__57_, chained_data_delayed_56__56_, chained_data_delayed_56__55_, chained_data_delayed_56__54_, chained_data_delayed_56__53_, chained_data_delayed_56__52_, chained_data_delayed_56__51_, chained_data_delayed_56__50_, chained_data_delayed_56__49_, chained_data_delayed_56__48_, chained_data_delayed_56__47_, chained_data_delayed_56__46_, chained_data_delayed_56__45_, chained_data_delayed_56__44_, chained_data_delayed_56__43_, chained_data_delayed_56__42_, chained_data_delayed_56__41_, chained_data_delayed_56__40_, chained_data_delayed_56__39_, chained_data_delayed_56__38_, chained_data_delayed_56__37_, chained_data_delayed_56__36_, chained_data_delayed_56__35_, chained_data_delayed_56__34_, chained_data_delayed_56__33_, chained_data_delayed_56__32_, chained_data_delayed_56__31_, chained_data_delayed_56__30_, chained_data_delayed_56__29_, chained_data_delayed_56__28_, chained_data_delayed_56__27_, chained_data_delayed_56__26_, chained_data_delayed_56__25_, chained_data_delayed_56__24_, chained_data_delayed_56__23_, chained_data_delayed_56__22_, chained_data_delayed_56__21_, chained_data_delayed_56__20_, chained_data_delayed_56__19_, chained_data_delayed_56__18_, chained_data_delayed_56__17_, chained_data_delayed_56__16_, chained_data_delayed_56__15_, chained_data_delayed_56__14_, chained_data_delayed_56__13_, chained_data_delayed_56__12_, chained_data_delayed_56__11_, chained_data_delayed_56__10_, chained_data_delayed_56__9_, chained_data_delayed_56__8_, chained_data_delayed_56__7_, chained_data_delayed_56__6_, chained_data_delayed_56__5_, chained_data_delayed_56__4_, chained_data_delayed_56__3_, chained_data_delayed_56__2_, chained_data_delayed_56__1_, chained_data_delayed_56__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_57__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_56__127_, chained_data_delayed_56__126_, chained_data_delayed_56__125_, chained_data_delayed_56__124_, chained_data_delayed_56__123_, chained_data_delayed_56__122_, chained_data_delayed_56__121_, chained_data_delayed_56__120_, chained_data_delayed_56__119_, chained_data_delayed_56__118_, chained_data_delayed_56__117_, chained_data_delayed_56__116_, chained_data_delayed_56__115_, chained_data_delayed_56__114_, chained_data_delayed_56__113_, chained_data_delayed_56__112_, chained_data_delayed_56__111_, chained_data_delayed_56__110_, chained_data_delayed_56__109_, chained_data_delayed_56__108_, chained_data_delayed_56__107_, chained_data_delayed_56__106_, chained_data_delayed_56__105_, chained_data_delayed_56__104_, chained_data_delayed_56__103_, chained_data_delayed_56__102_, chained_data_delayed_56__101_, chained_data_delayed_56__100_, chained_data_delayed_56__99_, chained_data_delayed_56__98_, chained_data_delayed_56__97_, chained_data_delayed_56__96_, chained_data_delayed_56__95_, chained_data_delayed_56__94_, chained_data_delayed_56__93_, chained_data_delayed_56__92_, chained_data_delayed_56__91_, chained_data_delayed_56__90_, chained_data_delayed_56__89_, chained_data_delayed_56__88_, chained_data_delayed_56__87_, chained_data_delayed_56__86_, chained_data_delayed_56__85_, chained_data_delayed_56__84_, chained_data_delayed_56__83_, chained_data_delayed_56__82_, chained_data_delayed_56__81_, chained_data_delayed_56__80_, chained_data_delayed_56__79_, chained_data_delayed_56__78_, chained_data_delayed_56__77_, chained_data_delayed_56__76_, chained_data_delayed_56__75_, chained_data_delayed_56__74_, chained_data_delayed_56__73_, chained_data_delayed_56__72_, chained_data_delayed_56__71_, chained_data_delayed_56__70_, chained_data_delayed_56__69_, chained_data_delayed_56__68_, chained_data_delayed_56__67_, chained_data_delayed_56__66_, chained_data_delayed_56__65_, chained_data_delayed_56__64_, chained_data_delayed_56__63_, chained_data_delayed_56__62_, chained_data_delayed_56__61_, chained_data_delayed_56__60_, chained_data_delayed_56__59_, chained_data_delayed_56__58_, chained_data_delayed_56__57_, chained_data_delayed_56__56_, chained_data_delayed_56__55_, chained_data_delayed_56__54_, chained_data_delayed_56__53_, chained_data_delayed_56__52_, chained_data_delayed_56__51_, chained_data_delayed_56__50_, chained_data_delayed_56__49_, chained_data_delayed_56__48_, chained_data_delayed_56__47_, chained_data_delayed_56__46_, chained_data_delayed_56__45_, chained_data_delayed_56__44_, chained_data_delayed_56__43_, chained_data_delayed_56__42_, chained_data_delayed_56__41_, chained_data_delayed_56__40_, chained_data_delayed_56__39_, chained_data_delayed_56__38_, chained_data_delayed_56__37_, chained_data_delayed_56__36_, chained_data_delayed_56__35_, chained_data_delayed_56__34_, chained_data_delayed_56__33_, chained_data_delayed_56__32_, chained_data_delayed_56__31_, chained_data_delayed_56__30_, chained_data_delayed_56__29_, chained_data_delayed_56__28_, chained_data_delayed_56__27_, chained_data_delayed_56__26_, chained_data_delayed_56__25_, chained_data_delayed_56__24_, chained_data_delayed_56__23_, chained_data_delayed_56__22_, chained_data_delayed_56__21_, chained_data_delayed_56__20_, chained_data_delayed_56__19_, chained_data_delayed_56__18_, chained_data_delayed_56__17_, chained_data_delayed_56__16_, chained_data_delayed_56__15_, chained_data_delayed_56__14_, chained_data_delayed_56__13_, chained_data_delayed_56__12_, chained_data_delayed_56__11_, chained_data_delayed_56__10_, chained_data_delayed_56__9_, chained_data_delayed_56__8_, chained_data_delayed_56__7_, chained_data_delayed_56__6_, chained_data_delayed_56__5_, chained_data_delayed_56__4_, chained_data_delayed_56__3_, chained_data_delayed_56__2_, chained_data_delayed_56__1_, chained_data_delayed_56__0_ }),
    .data_o({ chained_data_delayed_57__127_, chained_data_delayed_57__126_, chained_data_delayed_57__125_, chained_data_delayed_57__124_, chained_data_delayed_57__123_, chained_data_delayed_57__122_, chained_data_delayed_57__121_, chained_data_delayed_57__120_, chained_data_delayed_57__119_, chained_data_delayed_57__118_, chained_data_delayed_57__117_, chained_data_delayed_57__116_, chained_data_delayed_57__115_, chained_data_delayed_57__114_, chained_data_delayed_57__113_, chained_data_delayed_57__112_, chained_data_delayed_57__111_, chained_data_delayed_57__110_, chained_data_delayed_57__109_, chained_data_delayed_57__108_, chained_data_delayed_57__107_, chained_data_delayed_57__106_, chained_data_delayed_57__105_, chained_data_delayed_57__104_, chained_data_delayed_57__103_, chained_data_delayed_57__102_, chained_data_delayed_57__101_, chained_data_delayed_57__100_, chained_data_delayed_57__99_, chained_data_delayed_57__98_, chained_data_delayed_57__97_, chained_data_delayed_57__96_, chained_data_delayed_57__95_, chained_data_delayed_57__94_, chained_data_delayed_57__93_, chained_data_delayed_57__92_, chained_data_delayed_57__91_, chained_data_delayed_57__90_, chained_data_delayed_57__89_, chained_data_delayed_57__88_, chained_data_delayed_57__87_, chained_data_delayed_57__86_, chained_data_delayed_57__85_, chained_data_delayed_57__84_, chained_data_delayed_57__83_, chained_data_delayed_57__82_, chained_data_delayed_57__81_, chained_data_delayed_57__80_, chained_data_delayed_57__79_, chained_data_delayed_57__78_, chained_data_delayed_57__77_, chained_data_delayed_57__76_, chained_data_delayed_57__75_, chained_data_delayed_57__74_, chained_data_delayed_57__73_, chained_data_delayed_57__72_, chained_data_delayed_57__71_, chained_data_delayed_57__70_, chained_data_delayed_57__69_, chained_data_delayed_57__68_, chained_data_delayed_57__67_, chained_data_delayed_57__66_, chained_data_delayed_57__65_, chained_data_delayed_57__64_, chained_data_delayed_57__63_, chained_data_delayed_57__62_, chained_data_delayed_57__61_, chained_data_delayed_57__60_, chained_data_delayed_57__59_, chained_data_delayed_57__58_, chained_data_delayed_57__57_, chained_data_delayed_57__56_, chained_data_delayed_57__55_, chained_data_delayed_57__54_, chained_data_delayed_57__53_, chained_data_delayed_57__52_, chained_data_delayed_57__51_, chained_data_delayed_57__50_, chained_data_delayed_57__49_, chained_data_delayed_57__48_, chained_data_delayed_57__47_, chained_data_delayed_57__46_, chained_data_delayed_57__45_, chained_data_delayed_57__44_, chained_data_delayed_57__43_, chained_data_delayed_57__42_, chained_data_delayed_57__41_, chained_data_delayed_57__40_, chained_data_delayed_57__39_, chained_data_delayed_57__38_, chained_data_delayed_57__37_, chained_data_delayed_57__36_, chained_data_delayed_57__35_, chained_data_delayed_57__34_, chained_data_delayed_57__33_, chained_data_delayed_57__32_, chained_data_delayed_57__31_, chained_data_delayed_57__30_, chained_data_delayed_57__29_, chained_data_delayed_57__28_, chained_data_delayed_57__27_, chained_data_delayed_57__26_, chained_data_delayed_57__25_, chained_data_delayed_57__24_, chained_data_delayed_57__23_, chained_data_delayed_57__22_, chained_data_delayed_57__21_, chained_data_delayed_57__20_, chained_data_delayed_57__19_, chained_data_delayed_57__18_, chained_data_delayed_57__17_, chained_data_delayed_57__16_, chained_data_delayed_57__15_, chained_data_delayed_57__14_, chained_data_delayed_57__13_, chained_data_delayed_57__12_, chained_data_delayed_57__11_, chained_data_delayed_57__10_, chained_data_delayed_57__9_, chained_data_delayed_57__8_, chained_data_delayed_57__7_, chained_data_delayed_57__6_, chained_data_delayed_57__5_, chained_data_delayed_57__4_, chained_data_delayed_57__3_, chained_data_delayed_57__2_, chained_data_delayed_57__1_, chained_data_delayed_57__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_58__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_57__127_, chained_data_delayed_57__126_, chained_data_delayed_57__125_, chained_data_delayed_57__124_, chained_data_delayed_57__123_, chained_data_delayed_57__122_, chained_data_delayed_57__121_, chained_data_delayed_57__120_, chained_data_delayed_57__119_, chained_data_delayed_57__118_, chained_data_delayed_57__117_, chained_data_delayed_57__116_, chained_data_delayed_57__115_, chained_data_delayed_57__114_, chained_data_delayed_57__113_, chained_data_delayed_57__112_, chained_data_delayed_57__111_, chained_data_delayed_57__110_, chained_data_delayed_57__109_, chained_data_delayed_57__108_, chained_data_delayed_57__107_, chained_data_delayed_57__106_, chained_data_delayed_57__105_, chained_data_delayed_57__104_, chained_data_delayed_57__103_, chained_data_delayed_57__102_, chained_data_delayed_57__101_, chained_data_delayed_57__100_, chained_data_delayed_57__99_, chained_data_delayed_57__98_, chained_data_delayed_57__97_, chained_data_delayed_57__96_, chained_data_delayed_57__95_, chained_data_delayed_57__94_, chained_data_delayed_57__93_, chained_data_delayed_57__92_, chained_data_delayed_57__91_, chained_data_delayed_57__90_, chained_data_delayed_57__89_, chained_data_delayed_57__88_, chained_data_delayed_57__87_, chained_data_delayed_57__86_, chained_data_delayed_57__85_, chained_data_delayed_57__84_, chained_data_delayed_57__83_, chained_data_delayed_57__82_, chained_data_delayed_57__81_, chained_data_delayed_57__80_, chained_data_delayed_57__79_, chained_data_delayed_57__78_, chained_data_delayed_57__77_, chained_data_delayed_57__76_, chained_data_delayed_57__75_, chained_data_delayed_57__74_, chained_data_delayed_57__73_, chained_data_delayed_57__72_, chained_data_delayed_57__71_, chained_data_delayed_57__70_, chained_data_delayed_57__69_, chained_data_delayed_57__68_, chained_data_delayed_57__67_, chained_data_delayed_57__66_, chained_data_delayed_57__65_, chained_data_delayed_57__64_, chained_data_delayed_57__63_, chained_data_delayed_57__62_, chained_data_delayed_57__61_, chained_data_delayed_57__60_, chained_data_delayed_57__59_, chained_data_delayed_57__58_, chained_data_delayed_57__57_, chained_data_delayed_57__56_, chained_data_delayed_57__55_, chained_data_delayed_57__54_, chained_data_delayed_57__53_, chained_data_delayed_57__52_, chained_data_delayed_57__51_, chained_data_delayed_57__50_, chained_data_delayed_57__49_, chained_data_delayed_57__48_, chained_data_delayed_57__47_, chained_data_delayed_57__46_, chained_data_delayed_57__45_, chained_data_delayed_57__44_, chained_data_delayed_57__43_, chained_data_delayed_57__42_, chained_data_delayed_57__41_, chained_data_delayed_57__40_, chained_data_delayed_57__39_, chained_data_delayed_57__38_, chained_data_delayed_57__37_, chained_data_delayed_57__36_, chained_data_delayed_57__35_, chained_data_delayed_57__34_, chained_data_delayed_57__33_, chained_data_delayed_57__32_, chained_data_delayed_57__31_, chained_data_delayed_57__30_, chained_data_delayed_57__29_, chained_data_delayed_57__28_, chained_data_delayed_57__27_, chained_data_delayed_57__26_, chained_data_delayed_57__25_, chained_data_delayed_57__24_, chained_data_delayed_57__23_, chained_data_delayed_57__22_, chained_data_delayed_57__21_, chained_data_delayed_57__20_, chained_data_delayed_57__19_, chained_data_delayed_57__18_, chained_data_delayed_57__17_, chained_data_delayed_57__16_, chained_data_delayed_57__15_, chained_data_delayed_57__14_, chained_data_delayed_57__13_, chained_data_delayed_57__12_, chained_data_delayed_57__11_, chained_data_delayed_57__10_, chained_data_delayed_57__9_, chained_data_delayed_57__8_, chained_data_delayed_57__7_, chained_data_delayed_57__6_, chained_data_delayed_57__5_, chained_data_delayed_57__4_, chained_data_delayed_57__3_, chained_data_delayed_57__2_, chained_data_delayed_57__1_, chained_data_delayed_57__0_ }),
    .data_o({ chained_data_delayed_58__127_, chained_data_delayed_58__126_, chained_data_delayed_58__125_, chained_data_delayed_58__124_, chained_data_delayed_58__123_, chained_data_delayed_58__122_, chained_data_delayed_58__121_, chained_data_delayed_58__120_, chained_data_delayed_58__119_, chained_data_delayed_58__118_, chained_data_delayed_58__117_, chained_data_delayed_58__116_, chained_data_delayed_58__115_, chained_data_delayed_58__114_, chained_data_delayed_58__113_, chained_data_delayed_58__112_, chained_data_delayed_58__111_, chained_data_delayed_58__110_, chained_data_delayed_58__109_, chained_data_delayed_58__108_, chained_data_delayed_58__107_, chained_data_delayed_58__106_, chained_data_delayed_58__105_, chained_data_delayed_58__104_, chained_data_delayed_58__103_, chained_data_delayed_58__102_, chained_data_delayed_58__101_, chained_data_delayed_58__100_, chained_data_delayed_58__99_, chained_data_delayed_58__98_, chained_data_delayed_58__97_, chained_data_delayed_58__96_, chained_data_delayed_58__95_, chained_data_delayed_58__94_, chained_data_delayed_58__93_, chained_data_delayed_58__92_, chained_data_delayed_58__91_, chained_data_delayed_58__90_, chained_data_delayed_58__89_, chained_data_delayed_58__88_, chained_data_delayed_58__87_, chained_data_delayed_58__86_, chained_data_delayed_58__85_, chained_data_delayed_58__84_, chained_data_delayed_58__83_, chained_data_delayed_58__82_, chained_data_delayed_58__81_, chained_data_delayed_58__80_, chained_data_delayed_58__79_, chained_data_delayed_58__78_, chained_data_delayed_58__77_, chained_data_delayed_58__76_, chained_data_delayed_58__75_, chained_data_delayed_58__74_, chained_data_delayed_58__73_, chained_data_delayed_58__72_, chained_data_delayed_58__71_, chained_data_delayed_58__70_, chained_data_delayed_58__69_, chained_data_delayed_58__68_, chained_data_delayed_58__67_, chained_data_delayed_58__66_, chained_data_delayed_58__65_, chained_data_delayed_58__64_, chained_data_delayed_58__63_, chained_data_delayed_58__62_, chained_data_delayed_58__61_, chained_data_delayed_58__60_, chained_data_delayed_58__59_, chained_data_delayed_58__58_, chained_data_delayed_58__57_, chained_data_delayed_58__56_, chained_data_delayed_58__55_, chained_data_delayed_58__54_, chained_data_delayed_58__53_, chained_data_delayed_58__52_, chained_data_delayed_58__51_, chained_data_delayed_58__50_, chained_data_delayed_58__49_, chained_data_delayed_58__48_, chained_data_delayed_58__47_, chained_data_delayed_58__46_, chained_data_delayed_58__45_, chained_data_delayed_58__44_, chained_data_delayed_58__43_, chained_data_delayed_58__42_, chained_data_delayed_58__41_, chained_data_delayed_58__40_, chained_data_delayed_58__39_, chained_data_delayed_58__38_, chained_data_delayed_58__37_, chained_data_delayed_58__36_, chained_data_delayed_58__35_, chained_data_delayed_58__34_, chained_data_delayed_58__33_, chained_data_delayed_58__32_, chained_data_delayed_58__31_, chained_data_delayed_58__30_, chained_data_delayed_58__29_, chained_data_delayed_58__28_, chained_data_delayed_58__27_, chained_data_delayed_58__26_, chained_data_delayed_58__25_, chained_data_delayed_58__24_, chained_data_delayed_58__23_, chained_data_delayed_58__22_, chained_data_delayed_58__21_, chained_data_delayed_58__20_, chained_data_delayed_58__19_, chained_data_delayed_58__18_, chained_data_delayed_58__17_, chained_data_delayed_58__16_, chained_data_delayed_58__15_, chained_data_delayed_58__14_, chained_data_delayed_58__13_, chained_data_delayed_58__12_, chained_data_delayed_58__11_, chained_data_delayed_58__10_, chained_data_delayed_58__9_, chained_data_delayed_58__8_, chained_data_delayed_58__7_, chained_data_delayed_58__6_, chained_data_delayed_58__5_, chained_data_delayed_58__4_, chained_data_delayed_58__3_, chained_data_delayed_58__2_, chained_data_delayed_58__1_, chained_data_delayed_58__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_59__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_58__127_, chained_data_delayed_58__126_, chained_data_delayed_58__125_, chained_data_delayed_58__124_, chained_data_delayed_58__123_, chained_data_delayed_58__122_, chained_data_delayed_58__121_, chained_data_delayed_58__120_, chained_data_delayed_58__119_, chained_data_delayed_58__118_, chained_data_delayed_58__117_, chained_data_delayed_58__116_, chained_data_delayed_58__115_, chained_data_delayed_58__114_, chained_data_delayed_58__113_, chained_data_delayed_58__112_, chained_data_delayed_58__111_, chained_data_delayed_58__110_, chained_data_delayed_58__109_, chained_data_delayed_58__108_, chained_data_delayed_58__107_, chained_data_delayed_58__106_, chained_data_delayed_58__105_, chained_data_delayed_58__104_, chained_data_delayed_58__103_, chained_data_delayed_58__102_, chained_data_delayed_58__101_, chained_data_delayed_58__100_, chained_data_delayed_58__99_, chained_data_delayed_58__98_, chained_data_delayed_58__97_, chained_data_delayed_58__96_, chained_data_delayed_58__95_, chained_data_delayed_58__94_, chained_data_delayed_58__93_, chained_data_delayed_58__92_, chained_data_delayed_58__91_, chained_data_delayed_58__90_, chained_data_delayed_58__89_, chained_data_delayed_58__88_, chained_data_delayed_58__87_, chained_data_delayed_58__86_, chained_data_delayed_58__85_, chained_data_delayed_58__84_, chained_data_delayed_58__83_, chained_data_delayed_58__82_, chained_data_delayed_58__81_, chained_data_delayed_58__80_, chained_data_delayed_58__79_, chained_data_delayed_58__78_, chained_data_delayed_58__77_, chained_data_delayed_58__76_, chained_data_delayed_58__75_, chained_data_delayed_58__74_, chained_data_delayed_58__73_, chained_data_delayed_58__72_, chained_data_delayed_58__71_, chained_data_delayed_58__70_, chained_data_delayed_58__69_, chained_data_delayed_58__68_, chained_data_delayed_58__67_, chained_data_delayed_58__66_, chained_data_delayed_58__65_, chained_data_delayed_58__64_, chained_data_delayed_58__63_, chained_data_delayed_58__62_, chained_data_delayed_58__61_, chained_data_delayed_58__60_, chained_data_delayed_58__59_, chained_data_delayed_58__58_, chained_data_delayed_58__57_, chained_data_delayed_58__56_, chained_data_delayed_58__55_, chained_data_delayed_58__54_, chained_data_delayed_58__53_, chained_data_delayed_58__52_, chained_data_delayed_58__51_, chained_data_delayed_58__50_, chained_data_delayed_58__49_, chained_data_delayed_58__48_, chained_data_delayed_58__47_, chained_data_delayed_58__46_, chained_data_delayed_58__45_, chained_data_delayed_58__44_, chained_data_delayed_58__43_, chained_data_delayed_58__42_, chained_data_delayed_58__41_, chained_data_delayed_58__40_, chained_data_delayed_58__39_, chained_data_delayed_58__38_, chained_data_delayed_58__37_, chained_data_delayed_58__36_, chained_data_delayed_58__35_, chained_data_delayed_58__34_, chained_data_delayed_58__33_, chained_data_delayed_58__32_, chained_data_delayed_58__31_, chained_data_delayed_58__30_, chained_data_delayed_58__29_, chained_data_delayed_58__28_, chained_data_delayed_58__27_, chained_data_delayed_58__26_, chained_data_delayed_58__25_, chained_data_delayed_58__24_, chained_data_delayed_58__23_, chained_data_delayed_58__22_, chained_data_delayed_58__21_, chained_data_delayed_58__20_, chained_data_delayed_58__19_, chained_data_delayed_58__18_, chained_data_delayed_58__17_, chained_data_delayed_58__16_, chained_data_delayed_58__15_, chained_data_delayed_58__14_, chained_data_delayed_58__13_, chained_data_delayed_58__12_, chained_data_delayed_58__11_, chained_data_delayed_58__10_, chained_data_delayed_58__9_, chained_data_delayed_58__8_, chained_data_delayed_58__7_, chained_data_delayed_58__6_, chained_data_delayed_58__5_, chained_data_delayed_58__4_, chained_data_delayed_58__3_, chained_data_delayed_58__2_, chained_data_delayed_58__1_, chained_data_delayed_58__0_ }),
    .data_o({ chained_data_delayed_59__127_, chained_data_delayed_59__126_, chained_data_delayed_59__125_, chained_data_delayed_59__124_, chained_data_delayed_59__123_, chained_data_delayed_59__122_, chained_data_delayed_59__121_, chained_data_delayed_59__120_, chained_data_delayed_59__119_, chained_data_delayed_59__118_, chained_data_delayed_59__117_, chained_data_delayed_59__116_, chained_data_delayed_59__115_, chained_data_delayed_59__114_, chained_data_delayed_59__113_, chained_data_delayed_59__112_, chained_data_delayed_59__111_, chained_data_delayed_59__110_, chained_data_delayed_59__109_, chained_data_delayed_59__108_, chained_data_delayed_59__107_, chained_data_delayed_59__106_, chained_data_delayed_59__105_, chained_data_delayed_59__104_, chained_data_delayed_59__103_, chained_data_delayed_59__102_, chained_data_delayed_59__101_, chained_data_delayed_59__100_, chained_data_delayed_59__99_, chained_data_delayed_59__98_, chained_data_delayed_59__97_, chained_data_delayed_59__96_, chained_data_delayed_59__95_, chained_data_delayed_59__94_, chained_data_delayed_59__93_, chained_data_delayed_59__92_, chained_data_delayed_59__91_, chained_data_delayed_59__90_, chained_data_delayed_59__89_, chained_data_delayed_59__88_, chained_data_delayed_59__87_, chained_data_delayed_59__86_, chained_data_delayed_59__85_, chained_data_delayed_59__84_, chained_data_delayed_59__83_, chained_data_delayed_59__82_, chained_data_delayed_59__81_, chained_data_delayed_59__80_, chained_data_delayed_59__79_, chained_data_delayed_59__78_, chained_data_delayed_59__77_, chained_data_delayed_59__76_, chained_data_delayed_59__75_, chained_data_delayed_59__74_, chained_data_delayed_59__73_, chained_data_delayed_59__72_, chained_data_delayed_59__71_, chained_data_delayed_59__70_, chained_data_delayed_59__69_, chained_data_delayed_59__68_, chained_data_delayed_59__67_, chained_data_delayed_59__66_, chained_data_delayed_59__65_, chained_data_delayed_59__64_, chained_data_delayed_59__63_, chained_data_delayed_59__62_, chained_data_delayed_59__61_, chained_data_delayed_59__60_, chained_data_delayed_59__59_, chained_data_delayed_59__58_, chained_data_delayed_59__57_, chained_data_delayed_59__56_, chained_data_delayed_59__55_, chained_data_delayed_59__54_, chained_data_delayed_59__53_, chained_data_delayed_59__52_, chained_data_delayed_59__51_, chained_data_delayed_59__50_, chained_data_delayed_59__49_, chained_data_delayed_59__48_, chained_data_delayed_59__47_, chained_data_delayed_59__46_, chained_data_delayed_59__45_, chained_data_delayed_59__44_, chained_data_delayed_59__43_, chained_data_delayed_59__42_, chained_data_delayed_59__41_, chained_data_delayed_59__40_, chained_data_delayed_59__39_, chained_data_delayed_59__38_, chained_data_delayed_59__37_, chained_data_delayed_59__36_, chained_data_delayed_59__35_, chained_data_delayed_59__34_, chained_data_delayed_59__33_, chained_data_delayed_59__32_, chained_data_delayed_59__31_, chained_data_delayed_59__30_, chained_data_delayed_59__29_, chained_data_delayed_59__28_, chained_data_delayed_59__27_, chained_data_delayed_59__26_, chained_data_delayed_59__25_, chained_data_delayed_59__24_, chained_data_delayed_59__23_, chained_data_delayed_59__22_, chained_data_delayed_59__21_, chained_data_delayed_59__20_, chained_data_delayed_59__19_, chained_data_delayed_59__18_, chained_data_delayed_59__17_, chained_data_delayed_59__16_, chained_data_delayed_59__15_, chained_data_delayed_59__14_, chained_data_delayed_59__13_, chained_data_delayed_59__12_, chained_data_delayed_59__11_, chained_data_delayed_59__10_, chained_data_delayed_59__9_, chained_data_delayed_59__8_, chained_data_delayed_59__7_, chained_data_delayed_59__6_, chained_data_delayed_59__5_, chained_data_delayed_59__4_, chained_data_delayed_59__3_, chained_data_delayed_59__2_, chained_data_delayed_59__1_, chained_data_delayed_59__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_60__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_59__127_, chained_data_delayed_59__126_, chained_data_delayed_59__125_, chained_data_delayed_59__124_, chained_data_delayed_59__123_, chained_data_delayed_59__122_, chained_data_delayed_59__121_, chained_data_delayed_59__120_, chained_data_delayed_59__119_, chained_data_delayed_59__118_, chained_data_delayed_59__117_, chained_data_delayed_59__116_, chained_data_delayed_59__115_, chained_data_delayed_59__114_, chained_data_delayed_59__113_, chained_data_delayed_59__112_, chained_data_delayed_59__111_, chained_data_delayed_59__110_, chained_data_delayed_59__109_, chained_data_delayed_59__108_, chained_data_delayed_59__107_, chained_data_delayed_59__106_, chained_data_delayed_59__105_, chained_data_delayed_59__104_, chained_data_delayed_59__103_, chained_data_delayed_59__102_, chained_data_delayed_59__101_, chained_data_delayed_59__100_, chained_data_delayed_59__99_, chained_data_delayed_59__98_, chained_data_delayed_59__97_, chained_data_delayed_59__96_, chained_data_delayed_59__95_, chained_data_delayed_59__94_, chained_data_delayed_59__93_, chained_data_delayed_59__92_, chained_data_delayed_59__91_, chained_data_delayed_59__90_, chained_data_delayed_59__89_, chained_data_delayed_59__88_, chained_data_delayed_59__87_, chained_data_delayed_59__86_, chained_data_delayed_59__85_, chained_data_delayed_59__84_, chained_data_delayed_59__83_, chained_data_delayed_59__82_, chained_data_delayed_59__81_, chained_data_delayed_59__80_, chained_data_delayed_59__79_, chained_data_delayed_59__78_, chained_data_delayed_59__77_, chained_data_delayed_59__76_, chained_data_delayed_59__75_, chained_data_delayed_59__74_, chained_data_delayed_59__73_, chained_data_delayed_59__72_, chained_data_delayed_59__71_, chained_data_delayed_59__70_, chained_data_delayed_59__69_, chained_data_delayed_59__68_, chained_data_delayed_59__67_, chained_data_delayed_59__66_, chained_data_delayed_59__65_, chained_data_delayed_59__64_, chained_data_delayed_59__63_, chained_data_delayed_59__62_, chained_data_delayed_59__61_, chained_data_delayed_59__60_, chained_data_delayed_59__59_, chained_data_delayed_59__58_, chained_data_delayed_59__57_, chained_data_delayed_59__56_, chained_data_delayed_59__55_, chained_data_delayed_59__54_, chained_data_delayed_59__53_, chained_data_delayed_59__52_, chained_data_delayed_59__51_, chained_data_delayed_59__50_, chained_data_delayed_59__49_, chained_data_delayed_59__48_, chained_data_delayed_59__47_, chained_data_delayed_59__46_, chained_data_delayed_59__45_, chained_data_delayed_59__44_, chained_data_delayed_59__43_, chained_data_delayed_59__42_, chained_data_delayed_59__41_, chained_data_delayed_59__40_, chained_data_delayed_59__39_, chained_data_delayed_59__38_, chained_data_delayed_59__37_, chained_data_delayed_59__36_, chained_data_delayed_59__35_, chained_data_delayed_59__34_, chained_data_delayed_59__33_, chained_data_delayed_59__32_, chained_data_delayed_59__31_, chained_data_delayed_59__30_, chained_data_delayed_59__29_, chained_data_delayed_59__28_, chained_data_delayed_59__27_, chained_data_delayed_59__26_, chained_data_delayed_59__25_, chained_data_delayed_59__24_, chained_data_delayed_59__23_, chained_data_delayed_59__22_, chained_data_delayed_59__21_, chained_data_delayed_59__20_, chained_data_delayed_59__19_, chained_data_delayed_59__18_, chained_data_delayed_59__17_, chained_data_delayed_59__16_, chained_data_delayed_59__15_, chained_data_delayed_59__14_, chained_data_delayed_59__13_, chained_data_delayed_59__12_, chained_data_delayed_59__11_, chained_data_delayed_59__10_, chained_data_delayed_59__9_, chained_data_delayed_59__8_, chained_data_delayed_59__7_, chained_data_delayed_59__6_, chained_data_delayed_59__5_, chained_data_delayed_59__4_, chained_data_delayed_59__3_, chained_data_delayed_59__2_, chained_data_delayed_59__1_, chained_data_delayed_59__0_ }),
    .data_o({ chained_data_delayed_60__127_, chained_data_delayed_60__126_, chained_data_delayed_60__125_, chained_data_delayed_60__124_, chained_data_delayed_60__123_, chained_data_delayed_60__122_, chained_data_delayed_60__121_, chained_data_delayed_60__120_, chained_data_delayed_60__119_, chained_data_delayed_60__118_, chained_data_delayed_60__117_, chained_data_delayed_60__116_, chained_data_delayed_60__115_, chained_data_delayed_60__114_, chained_data_delayed_60__113_, chained_data_delayed_60__112_, chained_data_delayed_60__111_, chained_data_delayed_60__110_, chained_data_delayed_60__109_, chained_data_delayed_60__108_, chained_data_delayed_60__107_, chained_data_delayed_60__106_, chained_data_delayed_60__105_, chained_data_delayed_60__104_, chained_data_delayed_60__103_, chained_data_delayed_60__102_, chained_data_delayed_60__101_, chained_data_delayed_60__100_, chained_data_delayed_60__99_, chained_data_delayed_60__98_, chained_data_delayed_60__97_, chained_data_delayed_60__96_, chained_data_delayed_60__95_, chained_data_delayed_60__94_, chained_data_delayed_60__93_, chained_data_delayed_60__92_, chained_data_delayed_60__91_, chained_data_delayed_60__90_, chained_data_delayed_60__89_, chained_data_delayed_60__88_, chained_data_delayed_60__87_, chained_data_delayed_60__86_, chained_data_delayed_60__85_, chained_data_delayed_60__84_, chained_data_delayed_60__83_, chained_data_delayed_60__82_, chained_data_delayed_60__81_, chained_data_delayed_60__80_, chained_data_delayed_60__79_, chained_data_delayed_60__78_, chained_data_delayed_60__77_, chained_data_delayed_60__76_, chained_data_delayed_60__75_, chained_data_delayed_60__74_, chained_data_delayed_60__73_, chained_data_delayed_60__72_, chained_data_delayed_60__71_, chained_data_delayed_60__70_, chained_data_delayed_60__69_, chained_data_delayed_60__68_, chained_data_delayed_60__67_, chained_data_delayed_60__66_, chained_data_delayed_60__65_, chained_data_delayed_60__64_, chained_data_delayed_60__63_, chained_data_delayed_60__62_, chained_data_delayed_60__61_, chained_data_delayed_60__60_, chained_data_delayed_60__59_, chained_data_delayed_60__58_, chained_data_delayed_60__57_, chained_data_delayed_60__56_, chained_data_delayed_60__55_, chained_data_delayed_60__54_, chained_data_delayed_60__53_, chained_data_delayed_60__52_, chained_data_delayed_60__51_, chained_data_delayed_60__50_, chained_data_delayed_60__49_, chained_data_delayed_60__48_, chained_data_delayed_60__47_, chained_data_delayed_60__46_, chained_data_delayed_60__45_, chained_data_delayed_60__44_, chained_data_delayed_60__43_, chained_data_delayed_60__42_, chained_data_delayed_60__41_, chained_data_delayed_60__40_, chained_data_delayed_60__39_, chained_data_delayed_60__38_, chained_data_delayed_60__37_, chained_data_delayed_60__36_, chained_data_delayed_60__35_, chained_data_delayed_60__34_, chained_data_delayed_60__33_, chained_data_delayed_60__32_, chained_data_delayed_60__31_, chained_data_delayed_60__30_, chained_data_delayed_60__29_, chained_data_delayed_60__28_, chained_data_delayed_60__27_, chained_data_delayed_60__26_, chained_data_delayed_60__25_, chained_data_delayed_60__24_, chained_data_delayed_60__23_, chained_data_delayed_60__22_, chained_data_delayed_60__21_, chained_data_delayed_60__20_, chained_data_delayed_60__19_, chained_data_delayed_60__18_, chained_data_delayed_60__17_, chained_data_delayed_60__16_, chained_data_delayed_60__15_, chained_data_delayed_60__14_, chained_data_delayed_60__13_, chained_data_delayed_60__12_, chained_data_delayed_60__11_, chained_data_delayed_60__10_, chained_data_delayed_60__9_, chained_data_delayed_60__8_, chained_data_delayed_60__7_, chained_data_delayed_60__6_, chained_data_delayed_60__5_, chained_data_delayed_60__4_, chained_data_delayed_60__3_, chained_data_delayed_60__2_, chained_data_delayed_60__1_, chained_data_delayed_60__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_61__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_60__127_, chained_data_delayed_60__126_, chained_data_delayed_60__125_, chained_data_delayed_60__124_, chained_data_delayed_60__123_, chained_data_delayed_60__122_, chained_data_delayed_60__121_, chained_data_delayed_60__120_, chained_data_delayed_60__119_, chained_data_delayed_60__118_, chained_data_delayed_60__117_, chained_data_delayed_60__116_, chained_data_delayed_60__115_, chained_data_delayed_60__114_, chained_data_delayed_60__113_, chained_data_delayed_60__112_, chained_data_delayed_60__111_, chained_data_delayed_60__110_, chained_data_delayed_60__109_, chained_data_delayed_60__108_, chained_data_delayed_60__107_, chained_data_delayed_60__106_, chained_data_delayed_60__105_, chained_data_delayed_60__104_, chained_data_delayed_60__103_, chained_data_delayed_60__102_, chained_data_delayed_60__101_, chained_data_delayed_60__100_, chained_data_delayed_60__99_, chained_data_delayed_60__98_, chained_data_delayed_60__97_, chained_data_delayed_60__96_, chained_data_delayed_60__95_, chained_data_delayed_60__94_, chained_data_delayed_60__93_, chained_data_delayed_60__92_, chained_data_delayed_60__91_, chained_data_delayed_60__90_, chained_data_delayed_60__89_, chained_data_delayed_60__88_, chained_data_delayed_60__87_, chained_data_delayed_60__86_, chained_data_delayed_60__85_, chained_data_delayed_60__84_, chained_data_delayed_60__83_, chained_data_delayed_60__82_, chained_data_delayed_60__81_, chained_data_delayed_60__80_, chained_data_delayed_60__79_, chained_data_delayed_60__78_, chained_data_delayed_60__77_, chained_data_delayed_60__76_, chained_data_delayed_60__75_, chained_data_delayed_60__74_, chained_data_delayed_60__73_, chained_data_delayed_60__72_, chained_data_delayed_60__71_, chained_data_delayed_60__70_, chained_data_delayed_60__69_, chained_data_delayed_60__68_, chained_data_delayed_60__67_, chained_data_delayed_60__66_, chained_data_delayed_60__65_, chained_data_delayed_60__64_, chained_data_delayed_60__63_, chained_data_delayed_60__62_, chained_data_delayed_60__61_, chained_data_delayed_60__60_, chained_data_delayed_60__59_, chained_data_delayed_60__58_, chained_data_delayed_60__57_, chained_data_delayed_60__56_, chained_data_delayed_60__55_, chained_data_delayed_60__54_, chained_data_delayed_60__53_, chained_data_delayed_60__52_, chained_data_delayed_60__51_, chained_data_delayed_60__50_, chained_data_delayed_60__49_, chained_data_delayed_60__48_, chained_data_delayed_60__47_, chained_data_delayed_60__46_, chained_data_delayed_60__45_, chained_data_delayed_60__44_, chained_data_delayed_60__43_, chained_data_delayed_60__42_, chained_data_delayed_60__41_, chained_data_delayed_60__40_, chained_data_delayed_60__39_, chained_data_delayed_60__38_, chained_data_delayed_60__37_, chained_data_delayed_60__36_, chained_data_delayed_60__35_, chained_data_delayed_60__34_, chained_data_delayed_60__33_, chained_data_delayed_60__32_, chained_data_delayed_60__31_, chained_data_delayed_60__30_, chained_data_delayed_60__29_, chained_data_delayed_60__28_, chained_data_delayed_60__27_, chained_data_delayed_60__26_, chained_data_delayed_60__25_, chained_data_delayed_60__24_, chained_data_delayed_60__23_, chained_data_delayed_60__22_, chained_data_delayed_60__21_, chained_data_delayed_60__20_, chained_data_delayed_60__19_, chained_data_delayed_60__18_, chained_data_delayed_60__17_, chained_data_delayed_60__16_, chained_data_delayed_60__15_, chained_data_delayed_60__14_, chained_data_delayed_60__13_, chained_data_delayed_60__12_, chained_data_delayed_60__11_, chained_data_delayed_60__10_, chained_data_delayed_60__9_, chained_data_delayed_60__8_, chained_data_delayed_60__7_, chained_data_delayed_60__6_, chained_data_delayed_60__5_, chained_data_delayed_60__4_, chained_data_delayed_60__3_, chained_data_delayed_60__2_, chained_data_delayed_60__1_, chained_data_delayed_60__0_ }),
    .data_o({ chained_data_delayed_61__127_, chained_data_delayed_61__126_, chained_data_delayed_61__125_, chained_data_delayed_61__124_, chained_data_delayed_61__123_, chained_data_delayed_61__122_, chained_data_delayed_61__121_, chained_data_delayed_61__120_, chained_data_delayed_61__119_, chained_data_delayed_61__118_, chained_data_delayed_61__117_, chained_data_delayed_61__116_, chained_data_delayed_61__115_, chained_data_delayed_61__114_, chained_data_delayed_61__113_, chained_data_delayed_61__112_, chained_data_delayed_61__111_, chained_data_delayed_61__110_, chained_data_delayed_61__109_, chained_data_delayed_61__108_, chained_data_delayed_61__107_, chained_data_delayed_61__106_, chained_data_delayed_61__105_, chained_data_delayed_61__104_, chained_data_delayed_61__103_, chained_data_delayed_61__102_, chained_data_delayed_61__101_, chained_data_delayed_61__100_, chained_data_delayed_61__99_, chained_data_delayed_61__98_, chained_data_delayed_61__97_, chained_data_delayed_61__96_, chained_data_delayed_61__95_, chained_data_delayed_61__94_, chained_data_delayed_61__93_, chained_data_delayed_61__92_, chained_data_delayed_61__91_, chained_data_delayed_61__90_, chained_data_delayed_61__89_, chained_data_delayed_61__88_, chained_data_delayed_61__87_, chained_data_delayed_61__86_, chained_data_delayed_61__85_, chained_data_delayed_61__84_, chained_data_delayed_61__83_, chained_data_delayed_61__82_, chained_data_delayed_61__81_, chained_data_delayed_61__80_, chained_data_delayed_61__79_, chained_data_delayed_61__78_, chained_data_delayed_61__77_, chained_data_delayed_61__76_, chained_data_delayed_61__75_, chained_data_delayed_61__74_, chained_data_delayed_61__73_, chained_data_delayed_61__72_, chained_data_delayed_61__71_, chained_data_delayed_61__70_, chained_data_delayed_61__69_, chained_data_delayed_61__68_, chained_data_delayed_61__67_, chained_data_delayed_61__66_, chained_data_delayed_61__65_, chained_data_delayed_61__64_, chained_data_delayed_61__63_, chained_data_delayed_61__62_, chained_data_delayed_61__61_, chained_data_delayed_61__60_, chained_data_delayed_61__59_, chained_data_delayed_61__58_, chained_data_delayed_61__57_, chained_data_delayed_61__56_, chained_data_delayed_61__55_, chained_data_delayed_61__54_, chained_data_delayed_61__53_, chained_data_delayed_61__52_, chained_data_delayed_61__51_, chained_data_delayed_61__50_, chained_data_delayed_61__49_, chained_data_delayed_61__48_, chained_data_delayed_61__47_, chained_data_delayed_61__46_, chained_data_delayed_61__45_, chained_data_delayed_61__44_, chained_data_delayed_61__43_, chained_data_delayed_61__42_, chained_data_delayed_61__41_, chained_data_delayed_61__40_, chained_data_delayed_61__39_, chained_data_delayed_61__38_, chained_data_delayed_61__37_, chained_data_delayed_61__36_, chained_data_delayed_61__35_, chained_data_delayed_61__34_, chained_data_delayed_61__33_, chained_data_delayed_61__32_, chained_data_delayed_61__31_, chained_data_delayed_61__30_, chained_data_delayed_61__29_, chained_data_delayed_61__28_, chained_data_delayed_61__27_, chained_data_delayed_61__26_, chained_data_delayed_61__25_, chained_data_delayed_61__24_, chained_data_delayed_61__23_, chained_data_delayed_61__22_, chained_data_delayed_61__21_, chained_data_delayed_61__20_, chained_data_delayed_61__19_, chained_data_delayed_61__18_, chained_data_delayed_61__17_, chained_data_delayed_61__16_, chained_data_delayed_61__15_, chained_data_delayed_61__14_, chained_data_delayed_61__13_, chained_data_delayed_61__12_, chained_data_delayed_61__11_, chained_data_delayed_61__10_, chained_data_delayed_61__9_, chained_data_delayed_61__8_, chained_data_delayed_61__7_, chained_data_delayed_61__6_, chained_data_delayed_61__5_, chained_data_delayed_61__4_, chained_data_delayed_61__3_, chained_data_delayed_61__2_, chained_data_delayed_61__1_, chained_data_delayed_61__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_62__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_61__127_, chained_data_delayed_61__126_, chained_data_delayed_61__125_, chained_data_delayed_61__124_, chained_data_delayed_61__123_, chained_data_delayed_61__122_, chained_data_delayed_61__121_, chained_data_delayed_61__120_, chained_data_delayed_61__119_, chained_data_delayed_61__118_, chained_data_delayed_61__117_, chained_data_delayed_61__116_, chained_data_delayed_61__115_, chained_data_delayed_61__114_, chained_data_delayed_61__113_, chained_data_delayed_61__112_, chained_data_delayed_61__111_, chained_data_delayed_61__110_, chained_data_delayed_61__109_, chained_data_delayed_61__108_, chained_data_delayed_61__107_, chained_data_delayed_61__106_, chained_data_delayed_61__105_, chained_data_delayed_61__104_, chained_data_delayed_61__103_, chained_data_delayed_61__102_, chained_data_delayed_61__101_, chained_data_delayed_61__100_, chained_data_delayed_61__99_, chained_data_delayed_61__98_, chained_data_delayed_61__97_, chained_data_delayed_61__96_, chained_data_delayed_61__95_, chained_data_delayed_61__94_, chained_data_delayed_61__93_, chained_data_delayed_61__92_, chained_data_delayed_61__91_, chained_data_delayed_61__90_, chained_data_delayed_61__89_, chained_data_delayed_61__88_, chained_data_delayed_61__87_, chained_data_delayed_61__86_, chained_data_delayed_61__85_, chained_data_delayed_61__84_, chained_data_delayed_61__83_, chained_data_delayed_61__82_, chained_data_delayed_61__81_, chained_data_delayed_61__80_, chained_data_delayed_61__79_, chained_data_delayed_61__78_, chained_data_delayed_61__77_, chained_data_delayed_61__76_, chained_data_delayed_61__75_, chained_data_delayed_61__74_, chained_data_delayed_61__73_, chained_data_delayed_61__72_, chained_data_delayed_61__71_, chained_data_delayed_61__70_, chained_data_delayed_61__69_, chained_data_delayed_61__68_, chained_data_delayed_61__67_, chained_data_delayed_61__66_, chained_data_delayed_61__65_, chained_data_delayed_61__64_, chained_data_delayed_61__63_, chained_data_delayed_61__62_, chained_data_delayed_61__61_, chained_data_delayed_61__60_, chained_data_delayed_61__59_, chained_data_delayed_61__58_, chained_data_delayed_61__57_, chained_data_delayed_61__56_, chained_data_delayed_61__55_, chained_data_delayed_61__54_, chained_data_delayed_61__53_, chained_data_delayed_61__52_, chained_data_delayed_61__51_, chained_data_delayed_61__50_, chained_data_delayed_61__49_, chained_data_delayed_61__48_, chained_data_delayed_61__47_, chained_data_delayed_61__46_, chained_data_delayed_61__45_, chained_data_delayed_61__44_, chained_data_delayed_61__43_, chained_data_delayed_61__42_, chained_data_delayed_61__41_, chained_data_delayed_61__40_, chained_data_delayed_61__39_, chained_data_delayed_61__38_, chained_data_delayed_61__37_, chained_data_delayed_61__36_, chained_data_delayed_61__35_, chained_data_delayed_61__34_, chained_data_delayed_61__33_, chained_data_delayed_61__32_, chained_data_delayed_61__31_, chained_data_delayed_61__30_, chained_data_delayed_61__29_, chained_data_delayed_61__28_, chained_data_delayed_61__27_, chained_data_delayed_61__26_, chained_data_delayed_61__25_, chained_data_delayed_61__24_, chained_data_delayed_61__23_, chained_data_delayed_61__22_, chained_data_delayed_61__21_, chained_data_delayed_61__20_, chained_data_delayed_61__19_, chained_data_delayed_61__18_, chained_data_delayed_61__17_, chained_data_delayed_61__16_, chained_data_delayed_61__15_, chained_data_delayed_61__14_, chained_data_delayed_61__13_, chained_data_delayed_61__12_, chained_data_delayed_61__11_, chained_data_delayed_61__10_, chained_data_delayed_61__9_, chained_data_delayed_61__8_, chained_data_delayed_61__7_, chained_data_delayed_61__6_, chained_data_delayed_61__5_, chained_data_delayed_61__4_, chained_data_delayed_61__3_, chained_data_delayed_61__2_, chained_data_delayed_61__1_, chained_data_delayed_61__0_ }),
    .data_o({ chained_data_delayed_62__127_, chained_data_delayed_62__126_, chained_data_delayed_62__125_, chained_data_delayed_62__124_, chained_data_delayed_62__123_, chained_data_delayed_62__122_, chained_data_delayed_62__121_, chained_data_delayed_62__120_, chained_data_delayed_62__119_, chained_data_delayed_62__118_, chained_data_delayed_62__117_, chained_data_delayed_62__116_, chained_data_delayed_62__115_, chained_data_delayed_62__114_, chained_data_delayed_62__113_, chained_data_delayed_62__112_, chained_data_delayed_62__111_, chained_data_delayed_62__110_, chained_data_delayed_62__109_, chained_data_delayed_62__108_, chained_data_delayed_62__107_, chained_data_delayed_62__106_, chained_data_delayed_62__105_, chained_data_delayed_62__104_, chained_data_delayed_62__103_, chained_data_delayed_62__102_, chained_data_delayed_62__101_, chained_data_delayed_62__100_, chained_data_delayed_62__99_, chained_data_delayed_62__98_, chained_data_delayed_62__97_, chained_data_delayed_62__96_, chained_data_delayed_62__95_, chained_data_delayed_62__94_, chained_data_delayed_62__93_, chained_data_delayed_62__92_, chained_data_delayed_62__91_, chained_data_delayed_62__90_, chained_data_delayed_62__89_, chained_data_delayed_62__88_, chained_data_delayed_62__87_, chained_data_delayed_62__86_, chained_data_delayed_62__85_, chained_data_delayed_62__84_, chained_data_delayed_62__83_, chained_data_delayed_62__82_, chained_data_delayed_62__81_, chained_data_delayed_62__80_, chained_data_delayed_62__79_, chained_data_delayed_62__78_, chained_data_delayed_62__77_, chained_data_delayed_62__76_, chained_data_delayed_62__75_, chained_data_delayed_62__74_, chained_data_delayed_62__73_, chained_data_delayed_62__72_, chained_data_delayed_62__71_, chained_data_delayed_62__70_, chained_data_delayed_62__69_, chained_data_delayed_62__68_, chained_data_delayed_62__67_, chained_data_delayed_62__66_, chained_data_delayed_62__65_, chained_data_delayed_62__64_, chained_data_delayed_62__63_, chained_data_delayed_62__62_, chained_data_delayed_62__61_, chained_data_delayed_62__60_, chained_data_delayed_62__59_, chained_data_delayed_62__58_, chained_data_delayed_62__57_, chained_data_delayed_62__56_, chained_data_delayed_62__55_, chained_data_delayed_62__54_, chained_data_delayed_62__53_, chained_data_delayed_62__52_, chained_data_delayed_62__51_, chained_data_delayed_62__50_, chained_data_delayed_62__49_, chained_data_delayed_62__48_, chained_data_delayed_62__47_, chained_data_delayed_62__46_, chained_data_delayed_62__45_, chained_data_delayed_62__44_, chained_data_delayed_62__43_, chained_data_delayed_62__42_, chained_data_delayed_62__41_, chained_data_delayed_62__40_, chained_data_delayed_62__39_, chained_data_delayed_62__38_, chained_data_delayed_62__37_, chained_data_delayed_62__36_, chained_data_delayed_62__35_, chained_data_delayed_62__34_, chained_data_delayed_62__33_, chained_data_delayed_62__32_, chained_data_delayed_62__31_, chained_data_delayed_62__30_, chained_data_delayed_62__29_, chained_data_delayed_62__28_, chained_data_delayed_62__27_, chained_data_delayed_62__26_, chained_data_delayed_62__25_, chained_data_delayed_62__24_, chained_data_delayed_62__23_, chained_data_delayed_62__22_, chained_data_delayed_62__21_, chained_data_delayed_62__20_, chained_data_delayed_62__19_, chained_data_delayed_62__18_, chained_data_delayed_62__17_, chained_data_delayed_62__16_, chained_data_delayed_62__15_, chained_data_delayed_62__14_, chained_data_delayed_62__13_, chained_data_delayed_62__12_, chained_data_delayed_62__11_, chained_data_delayed_62__10_, chained_data_delayed_62__9_, chained_data_delayed_62__8_, chained_data_delayed_62__7_, chained_data_delayed_62__6_, chained_data_delayed_62__5_, chained_data_delayed_62__4_, chained_data_delayed_62__3_, chained_data_delayed_62__2_, chained_data_delayed_62__1_, chained_data_delayed_62__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_63__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_62__127_, chained_data_delayed_62__126_, chained_data_delayed_62__125_, chained_data_delayed_62__124_, chained_data_delayed_62__123_, chained_data_delayed_62__122_, chained_data_delayed_62__121_, chained_data_delayed_62__120_, chained_data_delayed_62__119_, chained_data_delayed_62__118_, chained_data_delayed_62__117_, chained_data_delayed_62__116_, chained_data_delayed_62__115_, chained_data_delayed_62__114_, chained_data_delayed_62__113_, chained_data_delayed_62__112_, chained_data_delayed_62__111_, chained_data_delayed_62__110_, chained_data_delayed_62__109_, chained_data_delayed_62__108_, chained_data_delayed_62__107_, chained_data_delayed_62__106_, chained_data_delayed_62__105_, chained_data_delayed_62__104_, chained_data_delayed_62__103_, chained_data_delayed_62__102_, chained_data_delayed_62__101_, chained_data_delayed_62__100_, chained_data_delayed_62__99_, chained_data_delayed_62__98_, chained_data_delayed_62__97_, chained_data_delayed_62__96_, chained_data_delayed_62__95_, chained_data_delayed_62__94_, chained_data_delayed_62__93_, chained_data_delayed_62__92_, chained_data_delayed_62__91_, chained_data_delayed_62__90_, chained_data_delayed_62__89_, chained_data_delayed_62__88_, chained_data_delayed_62__87_, chained_data_delayed_62__86_, chained_data_delayed_62__85_, chained_data_delayed_62__84_, chained_data_delayed_62__83_, chained_data_delayed_62__82_, chained_data_delayed_62__81_, chained_data_delayed_62__80_, chained_data_delayed_62__79_, chained_data_delayed_62__78_, chained_data_delayed_62__77_, chained_data_delayed_62__76_, chained_data_delayed_62__75_, chained_data_delayed_62__74_, chained_data_delayed_62__73_, chained_data_delayed_62__72_, chained_data_delayed_62__71_, chained_data_delayed_62__70_, chained_data_delayed_62__69_, chained_data_delayed_62__68_, chained_data_delayed_62__67_, chained_data_delayed_62__66_, chained_data_delayed_62__65_, chained_data_delayed_62__64_, chained_data_delayed_62__63_, chained_data_delayed_62__62_, chained_data_delayed_62__61_, chained_data_delayed_62__60_, chained_data_delayed_62__59_, chained_data_delayed_62__58_, chained_data_delayed_62__57_, chained_data_delayed_62__56_, chained_data_delayed_62__55_, chained_data_delayed_62__54_, chained_data_delayed_62__53_, chained_data_delayed_62__52_, chained_data_delayed_62__51_, chained_data_delayed_62__50_, chained_data_delayed_62__49_, chained_data_delayed_62__48_, chained_data_delayed_62__47_, chained_data_delayed_62__46_, chained_data_delayed_62__45_, chained_data_delayed_62__44_, chained_data_delayed_62__43_, chained_data_delayed_62__42_, chained_data_delayed_62__41_, chained_data_delayed_62__40_, chained_data_delayed_62__39_, chained_data_delayed_62__38_, chained_data_delayed_62__37_, chained_data_delayed_62__36_, chained_data_delayed_62__35_, chained_data_delayed_62__34_, chained_data_delayed_62__33_, chained_data_delayed_62__32_, chained_data_delayed_62__31_, chained_data_delayed_62__30_, chained_data_delayed_62__29_, chained_data_delayed_62__28_, chained_data_delayed_62__27_, chained_data_delayed_62__26_, chained_data_delayed_62__25_, chained_data_delayed_62__24_, chained_data_delayed_62__23_, chained_data_delayed_62__22_, chained_data_delayed_62__21_, chained_data_delayed_62__20_, chained_data_delayed_62__19_, chained_data_delayed_62__18_, chained_data_delayed_62__17_, chained_data_delayed_62__16_, chained_data_delayed_62__15_, chained_data_delayed_62__14_, chained_data_delayed_62__13_, chained_data_delayed_62__12_, chained_data_delayed_62__11_, chained_data_delayed_62__10_, chained_data_delayed_62__9_, chained_data_delayed_62__8_, chained_data_delayed_62__7_, chained_data_delayed_62__6_, chained_data_delayed_62__5_, chained_data_delayed_62__4_, chained_data_delayed_62__3_, chained_data_delayed_62__2_, chained_data_delayed_62__1_, chained_data_delayed_62__0_ }),
    .data_o({ chained_data_delayed_63__127_, chained_data_delayed_63__126_, chained_data_delayed_63__125_, chained_data_delayed_63__124_, chained_data_delayed_63__123_, chained_data_delayed_63__122_, chained_data_delayed_63__121_, chained_data_delayed_63__120_, chained_data_delayed_63__119_, chained_data_delayed_63__118_, chained_data_delayed_63__117_, chained_data_delayed_63__116_, chained_data_delayed_63__115_, chained_data_delayed_63__114_, chained_data_delayed_63__113_, chained_data_delayed_63__112_, chained_data_delayed_63__111_, chained_data_delayed_63__110_, chained_data_delayed_63__109_, chained_data_delayed_63__108_, chained_data_delayed_63__107_, chained_data_delayed_63__106_, chained_data_delayed_63__105_, chained_data_delayed_63__104_, chained_data_delayed_63__103_, chained_data_delayed_63__102_, chained_data_delayed_63__101_, chained_data_delayed_63__100_, chained_data_delayed_63__99_, chained_data_delayed_63__98_, chained_data_delayed_63__97_, chained_data_delayed_63__96_, chained_data_delayed_63__95_, chained_data_delayed_63__94_, chained_data_delayed_63__93_, chained_data_delayed_63__92_, chained_data_delayed_63__91_, chained_data_delayed_63__90_, chained_data_delayed_63__89_, chained_data_delayed_63__88_, chained_data_delayed_63__87_, chained_data_delayed_63__86_, chained_data_delayed_63__85_, chained_data_delayed_63__84_, chained_data_delayed_63__83_, chained_data_delayed_63__82_, chained_data_delayed_63__81_, chained_data_delayed_63__80_, chained_data_delayed_63__79_, chained_data_delayed_63__78_, chained_data_delayed_63__77_, chained_data_delayed_63__76_, chained_data_delayed_63__75_, chained_data_delayed_63__74_, chained_data_delayed_63__73_, chained_data_delayed_63__72_, chained_data_delayed_63__71_, chained_data_delayed_63__70_, chained_data_delayed_63__69_, chained_data_delayed_63__68_, chained_data_delayed_63__67_, chained_data_delayed_63__66_, chained_data_delayed_63__65_, chained_data_delayed_63__64_, chained_data_delayed_63__63_, chained_data_delayed_63__62_, chained_data_delayed_63__61_, chained_data_delayed_63__60_, chained_data_delayed_63__59_, chained_data_delayed_63__58_, chained_data_delayed_63__57_, chained_data_delayed_63__56_, chained_data_delayed_63__55_, chained_data_delayed_63__54_, chained_data_delayed_63__53_, chained_data_delayed_63__52_, chained_data_delayed_63__51_, chained_data_delayed_63__50_, chained_data_delayed_63__49_, chained_data_delayed_63__48_, chained_data_delayed_63__47_, chained_data_delayed_63__46_, chained_data_delayed_63__45_, chained_data_delayed_63__44_, chained_data_delayed_63__43_, chained_data_delayed_63__42_, chained_data_delayed_63__41_, chained_data_delayed_63__40_, chained_data_delayed_63__39_, chained_data_delayed_63__38_, chained_data_delayed_63__37_, chained_data_delayed_63__36_, chained_data_delayed_63__35_, chained_data_delayed_63__34_, chained_data_delayed_63__33_, chained_data_delayed_63__32_, chained_data_delayed_63__31_, chained_data_delayed_63__30_, chained_data_delayed_63__29_, chained_data_delayed_63__28_, chained_data_delayed_63__27_, chained_data_delayed_63__26_, chained_data_delayed_63__25_, chained_data_delayed_63__24_, chained_data_delayed_63__23_, chained_data_delayed_63__22_, chained_data_delayed_63__21_, chained_data_delayed_63__20_, chained_data_delayed_63__19_, chained_data_delayed_63__18_, chained_data_delayed_63__17_, chained_data_delayed_63__16_, chained_data_delayed_63__15_, chained_data_delayed_63__14_, chained_data_delayed_63__13_, chained_data_delayed_63__12_, chained_data_delayed_63__11_, chained_data_delayed_63__10_, chained_data_delayed_63__9_, chained_data_delayed_63__8_, chained_data_delayed_63__7_, chained_data_delayed_63__6_, chained_data_delayed_63__5_, chained_data_delayed_63__4_, chained_data_delayed_63__3_, chained_data_delayed_63__2_, chained_data_delayed_63__1_, chained_data_delayed_63__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_64__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_63__127_, chained_data_delayed_63__126_, chained_data_delayed_63__125_, chained_data_delayed_63__124_, chained_data_delayed_63__123_, chained_data_delayed_63__122_, chained_data_delayed_63__121_, chained_data_delayed_63__120_, chained_data_delayed_63__119_, chained_data_delayed_63__118_, chained_data_delayed_63__117_, chained_data_delayed_63__116_, chained_data_delayed_63__115_, chained_data_delayed_63__114_, chained_data_delayed_63__113_, chained_data_delayed_63__112_, chained_data_delayed_63__111_, chained_data_delayed_63__110_, chained_data_delayed_63__109_, chained_data_delayed_63__108_, chained_data_delayed_63__107_, chained_data_delayed_63__106_, chained_data_delayed_63__105_, chained_data_delayed_63__104_, chained_data_delayed_63__103_, chained_data_delayed_63__102_, chained_data_delayed_63__101_, chained_data_delayed_63__100_, chained_data_delayed_63__99_, chained_data_delayed_63__98_, chained_data_delayed_63__97_, chained_data_delayed_63__96_, chained_data_delayed_63__95_, chained_data_delayed_63__94_, chained_data_delayed_63__93_, chained_data_delayed_63__92_, chained_data_delayed_63__91_, chained_data_delayed_63__90_, chained_data_delayed_63__89_, chained_data_delayed_63__88_, chained_data_delayed_63__87_, chained_data_delayed_63__86_, chained_data_delayed_63__85_, chained_data_delayed_63__84_, chained_data_delayed_63__83_, chained_data_delayed_63__82_, chained_data_delayed_63__81_, chained_data_delayed_63__80_, chained_data_delayed_63__79_, chained_data_delayed_63__78_, chained_data_delayed_63__77_, chained_data_delayed_63__76_, chained_data_delayed_63__75_, chained_data_delayed_63__74_, chained_data_delayed_63__73_, chained_data_delayed_63__72_, chained_data_delayed_63__71_, chained_data_delayed_63__70_, chained_data_delayed_63__69_, chained_data_delayed_63__68_, chained_data_delayed_63__67_, chained_data_delayed_63__66_, chained_data_delayed_63__65_, chained_data_delayed_63__64_, chained_data_delayed_63__63_, chained_data_delayed_63__62_, chained_data_delayed_63__61_, chained_data_delayed_63__60_, chained_data_delayed_63__59_, chained_data_delayed_63__58_, chained_data_delayed_63__57_, chained_data_delayed_63__56_, chained_data_delayed_63__55_, chained_data_delayed_63__54_, chained_data_delayed_63__53_, chained_data_delayed_63__52_, chained_data_delayed_63__51_, chained_data_delayed_63__50_, chained_data_delayed_63__49_, chained_data_delayed_63__48_, chained_data_delayed_63__47_, chained_data_delayed_63__46_, chained_data_delayed_63__45_, chained_data_delayed_63__44_, chained_data_delayed_63__43_, chained_data_delayed_63__42_, chained_data_delayed_63__41_, chained_data_delayed_63__40_, chained_data_delayed_63__39_, chained_data_delayed_63__38_, chained_data_delayed_63__37_, chained_data_delayed_63__36_, chained_data_delayed_63__35_, chained_data_delayed_63__34_, chained_data_delayed_63__33_, chained_data_delayed_63__32_, chained_data_delayed_63__31_, chained_data_delayed_63__30_, chained_data_delayed_63__29_, chained_data_delayed_63__28_, chained_data_delayed_63__27_, chained_data_delayed_63__26_, chained_data_delayed_63__25_, chained_data_delayed_63__24_, chained_data_delayed_63__23_, chained_data_delayed_63__22_, chained_data_delayed_63__21_, chained_data_delayed_63__20_, chained_data_delayed_63__19_, chained_data_delayed_63__18_, chained_data_delayed_63__17_, chained_data_delayed_63__16_, chained_data_delayed_63__15_, chained_data_delayed_63__14_, chained_data_delayed_63__13_, chained_data_delayed_63__12_, chained_data_delayed_63__11_, chained_data_delayed_63__10_, chained_data_delayed_63__9_, chained_data_delayed_63__8_, chained_data_delayed_63__7_, chained_data_delayed_63__6_, chained_data_delayed_63__5_, chained_data_delayed_63__4_, chained_data_delayed_63__3_, chained_data_delayed_63__2_, chained_data_delayed_63__1_, chained_data_delayed_63__0_ }),
    .data_o({ chained_data_delayed_64__127_, chained_data_delayed_64__126_, chained_data_delayed_64__125_, chained_data_delayed_64__124_, chained_data_delayed_64__123_, chained_data_delayed_64__122_, chained_data_delayed_64__121_, chained_data_delayed_64__120_, chained_data_delayed_64__119_, chained_data_delayed_64__118_, chained_data_delayed_64__117_, chained_data_delayed_64__116_, chained_data_delayed_64__115_, chained_data_delayed_64__114_, chained_data_delayed_64__113_, chained_data_delayed_64__112_, chained_data_delayed_64__111_, chained_data_delayed_64__110_, chained_data_delayed_64__109_, chained_data_delayed_64__108_, chained_data_delayed_64__107_, chained_data_delayed_64__106_, chained_data_delayed_64__105_, chained_data_delayed_64__104_, chained_data_delayed_64__103_, chained_data_delayed_64__102_, chained_data_delayed_64__101_, chained_data_delayed_64__100_, chained_data_delayed_64__99_, chained_data_delayed_64__98_, chained_data_delayed_64__97_, chained_data_delayed_64__96_, chained_data_delayed_64__95_, chained_data_delayed_64__94_, chained_data_delayed_64__93_, chained_data_delayed_64__92_, chained_data_delayed_64__91_, chained_data_delayed_64__90_, chained_data_delayed_64__89_, chained_data_delayed_64__88_, chained_data_delayed_64__87_, chained_data_delayed_64__86_, chained_data_delayed_64__85_, chained_data_delayed_64__84_, chained_data_delayed_64__83_, chained_data_delayed_64__82_, chained_data_delayed_64__81_, chained_data_delayed_64__80_, chained_data_delayed_64__79_, chained_data_delayed_64__78_, chained_data_delayed_64__77_, chained_data_delayed_64__76_, chained_data_delayed_64__75_, chained_data_delayed_64__74_, chained_data_delayed_64__73_, chained_data_delayed_64__72_, chained_data_delayed_64__71_, chained_data_delayed_64__70_, chained_data_delayed_64__69_, chained_data_delayed_64__68_, chained_data_delayed_64__67_, chained_data_delayed_64__66_, chained_data_delayed_64__65_, chained_data_delayed_64__64_, chained_data_delayed_64__63_, chained_data_delayed_64__62_, chained_data_delayed_64__61_, chained_data_delayed_64__60_, chained_data_delayed_64__59_, chained_data_delayed_64__58_, chained_data_delayed_64__57_, chained_data_delayed_64__56_, chained_data_delayed_64__55_, chained_data_delayed_64__54_, chained_data_delayed_64__53_, chained_data_delayed_64__52_, chained_data_delayed_64__51_, chained_data_delayed_64__50_, chained_data_delayed_64__49_, chained_data_delayed_64__48_, chained_data_delayed_64__47_, chained_data_delayed_64__46_, chained_data_delayed_64__45_, chained_data_delayed_64__44_, chained_data_delayed_64__43_, chained_data_delayed_64__42_, chained_data_delayed_64__41_, chained_data_delayed_64__40_, chained_data_delayed_64__39_, chained_data_delayed_64__38_, chained_data_delayed_64__37_, chained_data_delayed_64__36_, chained_data_delayed_64__35_, chained_data_delayed_64__34_, chained_data_delayed_64__33_, chained_data_delayed_64__32_, chained_data_delayed_64__31_, chained_data_delayed_64__30_, chained_data_delayed_64__29_, chained_data_delayed_64__28_, chained_data_delayed_64__27_, chained_data_delayed_64__26_, chained_data_delayed_64__25_, chained_data_delayed_64__24_, chained_data_delayed_64__23_, chained_data_delayed_64__22_, chained_data_delayed_64__21_, chained_data_delayed_64__20_, chained_data_delayed_64__19_, chained_data_delayed_64__18_, chained_data_delayed_64__17_, chained_data_delayed_64__16_, chained_data_delayed_64__15_, chained_data_delayed_64__14_, chained_data_delayed_64__13_, chained_data_delayed_64__12_, chained_data_delayed_64__11_, chained_data_delayed_64__10_, chained_data_delayed_64__9_, chained_data_delayed_64__8_, chained_data_delayed_64__7_, chained_data_delayed_64__6_, chained_data_delayed_64__5_, chained_data_delayed_64__4_, chained_data_delayed_64__3_, chained_data_delayed_64__2_, chained_data_delayed_64__1_, chained_data_delayed_64__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_65__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_64__127_, chained_data_delayed_64__126_, chained_data_delayed_64__125_, chained_data_delayed_64__124_, chained_data_delayed_64__123_, chained_data_delayed_64__122_, chained_data_delayed_64__121_, chained_data_delayed_64__120_, chained_data_delayed_64__119_, chained_data_delayed_64__118_, chained_data_delayed_64__117_, chained_data_delayed_64__116_, chained_data_delayed_64__115_, chained_data_delayed_64__114_, chained_data_delayed_64__113_, chained_data_delayed_64__112_, chained_data_delayed_64__111_, chained_data_delayed_64__110_, chained_data_delayed_64__109_, chained_data_delayed_64__108_, chained_data_delayed_64__107_, chained_data_delayed_64__106_, chained_data_delayed_64__105_, chained_data_delayed_64__104_, chained_data_delayed_64__103_, chained_data_delayed_64__102_, chained_data_delayed_64__101_, chained_data_delayed_64__100_, chained_data_delayed_64__99_, chained_data_delayed_64__98_, chained_data_delayed_64__97_, chained_data_delayed_64__96_, chained_data_delayed_64__95_, chained_data_delayed_64__94_, chained_data_delayed_64__93_, chained_data_delayed_64__92_, chained_data_delayed_64__91_, chained_data_delayed_64__90_, chained_data_delayed_64__89_, chained_data_delayed_64__88_, chained_data_delayed_64__87_, chained_data_delayed_64__86_, chained_data_delayed_64__85_, chained_data_delayed_64__84_, chained_data_delayed_64__83_, chained_data_delayed_64__82_, chained_data_delayed_64__81_, chained_data_delayed_64__80_, chained_data_delayed_64__79_, chained_data_delayed_64__78_, chained_data_delayed_64__77_, chained_data_delayed_64__76_, chained_data_delayed_64__75_, chained_data_delayed_64__74_, chained_data_delayed_64__73_, chained_data_delayed_64__72_, chained_data_delayed_64__71_, chained_data_delayed_64__70_, chained_data_delayed_64__69_, chained_data_delayed_64__68_, chained_data_delayed_64__67_, chained_data_delayed_64__66_, chained_data_delayed_64__65_, chained_data_delayed_64__64_, chained_data_delayed_64__63_, chained_data_delayed_64__62_, chained_data_delayed_64__61_, chained_data_delayed_64__60_, chained_data_delayed_64__59_, chained_data_delayed_64__58_, chained_data_delayed_64__57_, chained_data_delayed_64__56_, chained_data_delayed_64__55_, chained_data_delayed_64__54_, chained_data_delayed_64__53_, chained_data_delayed_64__52_, chained_data_delayed_64__51_, chained_data_delayed_64__50_, chained_data_delayed_64__49_, chained_data_delayed_64__48_, chained_data_delayed_64__47_, chained_data_delayed_64__46_, chained_data_delayed_64__45_, chained_data_delayed_64__44_, chained_data_delayed_64__43_, chained_data_delayed_64__42_, chained_data_delayed_64__41_, chained_data_delayed_64__40_, chained_data_delayed_64__39_, chained_data_delayed_64__38_, chained_data_delayed_64__37_, chained_data_delayed_64__36_, chained_data_delayed_64__35_, chained_data_delayed_64__34_, chained_data_delayed_64__33_, chained_data_delayed_64__32_, chained_data_delayed_64__31_, chained_data_delayed_64__30_, chained_data_delayed_64__29_, chained_data_delayed_64__28_, chained_data_delayed_64__27_, chained_data_delayed_64__26_, chained_data_delayed_64__25_, chained_data_delayed_64__24_, chained_data_delayed_64__23_, chained_data_delayed_64__22_, chained_data_delayed_64__21_, chained_data_delayed_64__20_, chained_data_delayed_64__19_, chained_data_delayed_64__18_, chained_data_delayed_64__17_, chained_data_delayed_64__16_, chained_data_delayed_64__15_, chained_data_delayed_64__14_, chained_data_delayed_64__13_, chained_data_delayed_64__12_, chained_data_delayed_64__11_, chained_data_delayed_64__10_, chained_data_delayed_64__9_, chained_data_delayed_64__8_, chained_data_delayed_64__7_, chained_data_delayed_64__6_, chained_data_delayed_64__5_, chained_data_delayed_64__4_, chained_data_delayed_64__3_, chained_data_delayed_64__2_, chained_data_delayed_64__1_, chained_data_delayed_64__0_ }),
    .data_o({ chained_data_delayed_65__127_, chained_data_delayed_65__126_, chained_data_delayed_65__125_, chained_data_delayed_65__124_, chained_data_delayed_65__123_, chained_data_delayed_65__122_, chained_data_delayed_65__121_, chained_data_delayed_65__120_, chained_data_delayed_65__119_, chained_data_delayed_65__118_, chained_data_delayed_65__117_, chained_data_delayed_65__116_, chained_data_delayed_65__115_, chained_data_delayed_65__114_, chained_data_delayed_65__113_, chained_data_delayed_65__112_, chained_data_delayed_65__111_, chained_data_delayed_65__110_, chained_data_delayed_65__109_, chained_data_delayed_65__108_, chained_data_delayed_65__107_, chained_data_delayed_65__106_, chained_data_delayed_65__105_, chained_data_delayed_65__104_, chained_data_delayed_65__103_, chained_data_delayed_65__102_, chained_data_delayed_65__101_, chained_data_delayed_65__100_, chained_data_delayed_65__99_, chained_data_delayed_65__98_, chained_data_delayed_65__97_, chained_data_delayed_65__96_, chained_data_delayed_65__95_, chained_data_delayed_65__94_, chained_data_delayed_65__93_, chained_data_delayed_65__92_, chained_data_delayed_65__91_, chained_data_delayed_65__90_, chained_data_delayed_65__89_, chained_data_delayed_65__88_, chained_data_delayed_65__87_, chained_data_delayed_65__86_, chained_data_delayed_65__85_, chained_data_delayed_65__84_, chained_data_delayed_65__83_, chained_data_delayed_65__82_, chained_data_delayed_65__81_, chained_data_delayed_65__80_, chained_data_delayed_65__79_, chained_data_delayed_65__78_, chained_data_delayed_65__77_, chained_data_delayed_65__76_, chained_data_delayed_65__75_, chained_data_delayed_65__74_, chained_data_delayed_65__73_, chained_data_delayed_65__72_, chained_data_delayed_65__71_, chained_data_delayed_65__70_, chained_data_delayed_65__69_, chained_data_delayed_65__68_, chained_data_delayed_65__67_, chained_data_delayed_65__66_, chained_data_delayed_65__65_, chained_data_delayed_65__64_, chained_data_delayed_65__63_, chained_data_delayed_65__62_, chained_data_delayed_65__61_, chained_data_delayed_65__60_, chained_data_delayed_65__59_, chained_data_delayed_65__58_, chained_data_delayed_65__57_, chained_data_delayed_65__56_, chained_data_delayed_65__55_, chained_data_delayed_65__54_, chained_data_delayed_65__53_, chained_data_delayed_65__52_, chained_data_delayed_65__51_, chained_data_delayed_65__50_, chained_data_delayed_65__49_, chained_data_delayed_65__48_, chained_data_delayed_65__47_, chained_data_delayed_65__46_, chained_data_delayed_65__45_, chained_data_delayed_65__44_, chained_data_delayed_65__43_, chained_data_delayed_65__42_, chained_data_delayed_65__41_, chained_data_delayed_65__40_, chained_data_delayed_65__39_, chained_data_delayed_65__38_, chained_data_delayed_65__37_, chained_data_delayed_65__36_, chained_data_delayed_65__35_, chained_data_delayed_65__34_, chained_data_delayed_65__33_, chained_data_delayed_65__32_, chained_data_delayed_65__31_, chained_data_delayed_65__30_, chained_data_delayed_65__29_, chained_data_delayed_65__28_, chained_data_delayed_65__27_, chained_data_delayed_65__26_, chained_data_delayed_65__25_, chained_data_delayed_65__24_, chained_data_delayed_65__23_, chained_data_delayed_65__22_, chained_data_delayed_65__21_, chained_data_delayed_65__20_, chained_data_delayed_65__19_, chained_data_delayed_65__18_, chained_data_delayed_65__17_, chained_data_delayed_65__16_, chained_data_delayed_65__15_, chained_data_delayed_65__14_, chained_data_delayed_65__13_, chained_data_delayed_65__12_, chained_data_delayed_65__11_, chained_data_delayed_65__10_, chained_data_delayed_65__9_, chained_data_delayed_65__8_, chained_data_delayed_65__7_, chained_data_delayed_65__6_, chained_data_delayed_65__5_, chained_data_delayed_65__4_, chained_data_delayed_65__3_, chained_data_delayed_65__2_, chained_data_delayed_65__1_, chained_data_delayed_65__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_66__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_65__127_, chained_data_delayed_65__126_, chained_data_delayed_65__125_, chained_data_delayed_65__124_, chained_data_delayed_65__123_, chained_data_delayed_65__122_, chained_data_delayed_65__121_, chained_data_delayed_65__120_, chained_data_delayed_65__119_, chained_data_delayed_65__118_, chained_data_delayed_65__117_, chained_data_delayed_65__116_, chained_data_delayed_65__115_, chained_data_delayed_65__114_, chained_data_delayed_65__113_, chained_data_delayed_65__112_, chained_data_delayed_65__111_, chained_data_delayed_65__110_, chained_data_delayed_65__109_, chained_data_delayed_65__108_, chained_data_delayed_65__107_, chained_data_delayed_65__106_, chained_data_delayed_65__105_, chained_data_delayed_65__104_, chained_data_delayed_65__103_, chained_data_delayed_65__102_, chained_data_delayed_65__101_, chained_data_delayed_65__100_, chained_data_delayed_65__99_, chained_data_delayed_65__98_, chained_data_delayed_65__97_, chained_data_delayed_65__96_, chained_data_delayed_65__95_, chained_data_delayed_65__94_, chained_data_delayed_65__93_, chained_data_delayed_65__92_, chained_data_delayed_65__91_, chained_data_delayed_65__90_, chained_data_delayed_65__89_, chained_data_delayed_65__88_, chained_data_delayed_65__87_, chained_data_delayed_65__86_, chained_data_delayed_65__85_, chained_data_delayed_65__84_, chained_data_delayed_65__83_, chained_data_delayed_65__82_, chained_data_delayed_65__81_, chained_data_delayed_65__80_, chained_data_delayed_65__79_, chained_data_delayed_65__78_, chained_data_delayed_65__77_, chained_data_delayed_65__76_, chained_data_delayed_65__75_, chained_data_delayed_65__74_, chained_data_delayed_65__73_, chained_data_delayed_65__72_, chained_data_delayed_65__71_, chained_data_delayed_65__70_, chained_data_delayed_65__69_, chained_data_delayed_65__68_, chained_data_delayed_65__67_, chained_data_delayed_65__66_, chained_data_delayed_65__65_, chained_data_delayed_65__64_, chained_data_delayed_65__63_, chained_data_delayed_65__62_, chained_data_delayed_65__61_, chained_data_delayed_65__60_, chained_data_delayed_65__59_, chained_data_delayed_65__58_, chained_data_delayed_65__57_, chained_data_delayed_65__56_, chained_data_delayed_65__55_, chained_data_delayed_65__54_, chained_data_delayed_65__53_, chained_data_delayed_65__52_, chained_data_delayed_65__51_, chained_data_delayed_65__50_, chained_data_delayed_65__49_, chained_data_delayed_65__48_, chained_data_delayed_65__47_, chained_data_delayed_65__46_, chained_data_delayed_65__45_, chained_data_delayed_65__44_, chained_data_delayed_65__43_, chained_data_delayed_65__42_, chained_data_delayed_65__41_, chained_data_delayed_65__40_, chained_data_delayed_65__39_, chained_data_delayed_65__38_, chained_data_delayed_65__37_, chained_data_delayed_65__36_, chained_data_delayed_65__35_, chained_data_delayed_65__34_, chained_data_delayed_65__33_, chained_data_delayed_65__32_, chained_data_delayed_65__31_, chained_data_delayed_65__30_, chained_data_delayed_65__29_, chained_data_delayed_65__28_, chained_data_delayed_65__27_, chained_data_delayed_65__26_, chained_data_delayed_65__25_, chained_data_delayed_65__24_, chained_data_delayed_65__23_, chained_data_delayed_65__22_, chained_data_delayed_65__21_, chained_data_delayed_65__20_, chained_data_delayed_65__19_, chained_data_delayed_65__18_, chained_data_delayed_65__17_, chained_data_delayed_65__16_, chained_data_delayed_65__15_, chained_data_delayed_65__14_, chained_data_delayed_65__13_, chained_data_delayed_65__12_, chained_data_delayed_65__11_, chained_data_delayed_65__10_, chained_data_delayed_65__9_, chained_data_delayed_65__8_, chained_data_delayed_65__7_, chained_data_delayed_65__6_, chained_data_delayed_65__5_, chained_data_delayed_65__4_, chained_data_delayed_65__3_, chained_data_delayed_65__2_, chained_data_delayed_65__1_, chained_data_delayed_65__0_ }),
    .data_o({ chained_data_delayed_66__127_, chained_data_delayed_66__126_, chained_data_delayed_66__125_, chained_data_delayed_66__124_, chained_data_delayed_66__123_, chained_data_delayed_66__122_, chained_data_delayed_66__121_, chained_data_delayed_66__120_, chained_data_delayed_66__119_, chained_data_delayed_66__118_, chained_data_delayed_66__117_, chained_data_delayed_66__116_, chained_data_delayed_66__115_, chained_data_delayed_66__114_, chained_data_delayed_66__113_, chained_data_delayed_66__112_, chained_data_delayed_66__111_, chained_data_delayed_66__110_, chained_data_delayed_66__109_, chained_data_delayed_66__108_, chained_data_delayed_66__107_, chained_data_delayed_66__106_, chained_data_delayed_66__105_, chained_data_delayed_66__104_, chained_data_delayed_66__103_, chained_data_delayed_66__102_, chained_data_delayed_66__101_, chained_data_delayed_66__100_, chained_data_delayed_66__99_, chained_data_delayed_66__98_, chained_data_delayed_66__97_, chained_data_delayed_66__96_, chained_data_delayed_66__95_, chained_data_delayed_66__94_, chained_data_delayed_66__93_, chained_data_delayed_66__92_, chained_data_delayed_66__91_, chained_data_delayed_66__90_, chained_data_delayed_66__89_, chained_data_delayed_66__88_, chained_data_delayed_66__87_, chained_data_delayed_66__86_, chained_data_delayed_66__85_, chained_data_delayed_66__84_, chained_data_delayed_66__83_, chained_data_delayed_66__82_, chained_data_delayed_66__81_, chained_data_delayed_66__80_, chained_data_delayed_66__79_, chained_data_delayed_66__78_, chained_data_delayed_66__77_, chained_data_delayed_66__76_, chained_data_delayed_66__75_, chained_data_delayed_66__74_, chained_data_delayed_66__73_, chained_data_delayed_66__72_, chained_data_delayed_66__71_, chained_data_delayed_66__70_, chained_data_delayed_66__69_, chained_data_delayed_66__68_, chained_data_delayed_66__67_, chained_data_delayed_66__66_, chained_data_delayed_66__65_, chained_data_delayed_66__64_, chained_data_delayed_66__63_, chained_data_delayed_66__62_, chained_data_delayed_66__61_, chained_data_delayed_66__60_, chained_data_delayed_66__59_, chained_data_delayed_66__58_, chained_data_delayed_66__57_, chained_data_delayed_66__56_, chained_data_delayed_66__55_, chained_data_delayed_66__54_, chained_data_delayed_66__53_, chained_data_delayed_66__52_, chained_data_delayed_66__51_, chained_data_delayed_66__50_, chained_data_delayed_66__49_, chained_data_delayed_66__48_, chained_data_delayed_66__47_, chained_data_delayed_66__46_, chained_data_delayed_66__45_, chained_data_delayed_66__44_, chained_data_delayed_66__43_, chained_data_delayed_66__42_, chained_data_delayed_66__41_, chained_data_delayed_66__40_, chained_data_delayed_66__39_, chained_data_delayed_66__38_, chained_data_delayed_66__37_, chained_data_delayed_66__36_, chained_data_delayed_66__35_, chained_data_delayed_66__34_, chained_data_delayed_66__33_, chained_data_delayed_66__32_, chained_data_delayed_66__31_, chained_data_delayed_66__30_, chained_data_delayed_66__29_, chained_data_delayed_66__28_, chained_data_delayed_66__27_, chained_data_delayed_66__26_, chained_data_delayed_66__25_, chained_data_delayed_66__24_, chained_data_delayed_66__23_, chained_data_delayed_66__22_, chained_data_delayed_66__21_, chained_data_delayed_66__20_, chained_data_delayed_66__19_, chained_data_delayed_66__18_, chained_data_delayed_66__17_, chained_data_delayed_66__16_, chained_data_delayed_66__15_, chained_data_delayed_66__14_, chained_data_delayed_66__13_, chained_data_delayed_66__12_, chained_data_delayed_66__11_, chained_data_delayed_66__10_, chained_data_delayed_66__9_, chained_data_delayed_66__8_, chained_data_delayed_66__7_, chained_data_delayed_66__6_, chained_data_delayed_66__5_, chained_data_delayed_66__4_, chained_data_delayed_66__3_, chained_data_delayed_66__2_, chained_data_delayed_66__1_, chained_data_delayed_66__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_67__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_66__127_, chained_data_delayed_66__126_, chained_data_delayed_66__125_, chained_data_delayed_66__124_, chained_data_delayed_66__123_, chained_data_delayed_66__122_, chained_data_delayed_66__121_, chained_data_delayed_66__120_, chained_data_delayed_66__119_, chained_data_delayed_66__118_, chained_data_delayed_66__117_, chained_data_delayed_66__116_, chained_data_delayed_66__115_, chained_data_delayed_66__114_, chained_data_delayed_66__113_, chained_data_delayed_66__112_, chained_data_delayed_66__111_, chained_data_delayed_66__110_, chained_data_delayed_66__109_, chained_data_delayed_66__108_, chained_data_delayed_66__107_, chained_data_delayed_66__106_, chained_data_delayed_66__105_, chained_data_delayed_66__104_, chained_data_delayed_66__103_, chained_data_delayed_66__102_, chained_data_delayed_66__101_, chained_data_delayed_66__100_, chained_data_delayed_66__99_, chained_data_delayed_66__98_, chained_data_delayed_66__97_, chained_data_delayed_66__96_, chained_data_delayed_66__95_, chained_data_delayed_66__94_, chained_data_delayed_66__93_, chained_data_delayed_66__92_, chained_data_delayed_66__91_, chained_data_delayed_66__90_, chained_data_delayed_66__89_, chained_data_delayed_66__88_, chained_data_delayed_66__87_, chained_data_delayed_66__86_, chained_data_delayed_66__85_, chained_data_delayed_66__84_, chained_data_delayed_66__83_, chained_data_delayed_66__82_, chained_data_delayed_66__81_, chained_data_delayed_66__80_, chained_data_delayed_66__79_, chained_data_delayed_66__78_, chained_data_delayed_66__77_, chained_data_delayed_66__76_, chained_data_delayed_66__75_, chained_data_delayed_66__74_, chained_data_delayed_66__73_, chained_data_delayed_66__72_, chained_data_delayed_66__71_, chained_data_delayed_66__70_, chained_data_delayed_66__69_, chained_data_delayed_66__68_, chained_data_delayed_66__67_, chained_data_delayed_66__66_, chained_data_delayed_66__65_, chained_data_delayed_66__64_, chained_data_delayed_66__63_, chained_data_delayed_66__62_, chained_data_delayed_66__61_, chained_data_delayed_66__60_, chained_data_delayed_66__59_, chained_data_delayed_66__58_, chained_data_delayed_66__57_, chained_data_delayed_66__56_, chained_data_delayed_66__55_, chained_data_delayed_66__54_, chained_data_delayed_66__53_, chained_data_delayed_66__52_, chained_data_delayed_66__51_, chained_data_delayed_66__50_, chained_data_delayed_66__49_, chained_data_delayed_66__48_, chained_data_delayed_66__47_, chained_data_delayed_66__46_, chained_data_delayed_66__45_, chained_data_delayed_66__44_, chained_data_delayed_66__43_, chained_data_delayed_66__42_, chained_data_delayed_66__41_, chained_data_delayed_66__40_, chained_data_delayed_66__39_, chained_data_delayed_66__38_, chained_data_delayed_66__37_, chained_data_delayed_66__36_, chained_data_delayed_66__35_, chained_data_delayed_66__34_, chained_data_delayed_66__33_, chained_data_delayed_66__32_, chained_data_delayed_66__31_, chained_data_delayed_66__30_, chained_data_delayed_66__29_, chained_data_delayed_66__28_, chained_data_delayed_66__27_, chained_data_delayed_66__26_, chained_data_delayed_66__25_, chained_data_delayed_66__24_, chained_data_delayed_66__23_, chained_data_delayed_66__22_, chained_data_delayed_66__21_, chained_data_delayed_66__20_, chained_data_delayed_66__19_, chained_data_delayed_66__18_, chained_data_delayed_66__17_, chained_data_delayed_66__16_, chained_data_delayed_66__15_, chained_data_delayed_66__14_, chained_data_delayed_66__13_, chained_data_delayed_66__12_, chained_data_delayed_66__11_, chained_data_delayed_66__10_, chained_data_delayed_66__9_, chained_data_delayed_66__8_, chained_data_delayed_66__7_, chained_data_delayed_66__6_, chained_data_delayed_66__5_, chained_data_delayed_66__4_, chained_data_delayed_66__3_, chained_data_delayed_66__2_, chained_data_delayed_66__1_, chained_data_delayed_66__0_ }),
    .data_o({ chained_data_delayed_67__127_, chained_data_delayed_67__126_, chained_data_delayed_67__125_, chained_data_delayed_67__124_, chained_data_delayed_67__123_, chained_data_delayed_67__122_, chained_data_delayed_67__121_, chained_data_delayed_67__120_, chained_data_delayed_67__119_, chained_data_delayed_67__118_, chained_data_delayed_67__117_, chained_data_delayed_67__116_, chained_data_delayed_67__115_, chained_data_delayed_67__114_, chained_data_delayed_67__113_, chained_data_delayed_67__112_, chained_data_delayed_67__111_, chained_data_delayed_67__110_, chained_data_delayed_67__109_, chained_data_delayed_67__108_, chained_data_delayed_67__107_, chained_data_delayed_67__106_, chained_data_delayed_67__105_, chained_data_delayed_67__104_, chained_data_delayed_67__103_, chained_data_delayed_67__102_, chained_data_delayed_67__101_, chained_data_delayed_67__100_, chained_data_delayed_67__99_, chained_data_delayed_67__98_, chained_data_delayed_67__97_, chained_data_delayed_67__96_, chained_data_delayed_67__95_, chained_data_delayed_67__94_, chained_data_delayed_67__93_, chained_data_delayed_67__92_, chained_data_delayed_67__91_, chained_data_delayed_67__90_, chained_data_delayed_67__89_, chained_data_delayed_67__88_, chained_data_delayed_67__87_, chained_data_delayed_67__86_, chained_data_delayed_67__85_, chained_data_delayed_67__84_, chained_data_delayed_67__83_, chained_data_delayed_67__82_, chained_data_delayed_67__81_, chained_data_delayed_67__80_, chained_data_delayed_67__79_, chained_data_delayed_67__78_, chained_data_delayed_67__77_, chained_data_delayed_67__76_, chained_data_delayed_67__75_, chained_data_delayed_67__74_, chained_data_delayed_67__73_, chained_data_delayed_67__72_, chained_data_delayed_67__71_, chained_data_delayed_67__70_, chained_data_delayed_67__69_, chained_data_delayed_67__68_, chained_data_delayed_67__67_, chained_data_delayed_67__66_, chained_data_delayed_67__65_, chained_data_delayed_67__64_, chained_data_delayed_67__63_, chained_data_delayed_67__62_, chained_data_delayed_67__61_, chained_data_delayed_67__60_, chained_data_delayed_67__59_, chained_data_delayed_67__58_, chained_data_delayed_67__57_, chained_data_delayed_67__56_, chained_data_delayed_67__55_, chained_data_delayed_67__54_, chained_data_delayed_67__53_, chained_data_delayed_67__52_, chained_data_delayed_67__51_, chained_data_delayed_67__50_, chained_data_delayed_67__49_, chained_data_delayed_67__48_, chained_data_delayed_67__47_, chained_data_delayed_67__46_, chained_data_delayed_67__45_, chained_data_delayed_67__44_, chained_data_delayed_67__43_, chained_data_delayed_67__42_, chained_data_delayed_67__41_, chained_data_delayed_67__40_, chained_data_delayed_67__39_, chained_data_delayed_67__38_, chained_data_delayed_67__37_, chained_data_delayed_67__36_, chained_data_delayed_67__35_, chained_data_delayed_67__34_, chained_data_delayed_67__33_, chained_data_delayed_67__32_, chained_data_delayed_67__31_, chained_data_delayed_67__30_, chained_data_delayed_67__29_, chained_data_delayed_67__28_, chained_data_delayed_67__27_, chained_data_delayed_67__26_, chained_data_delayed_67__25_, chained_data_delayed_67__24_, chained_data_delayed_67__23_, chained_data_delayed_67__22_, chained_data_delayed_67__21_, chained_data_delayed_67__20_, chained_data_delayed_67__19_, chained_data_delayed_67__18_, chained_data_delayed_67__17_, chained_data_delayed_67__16_, chained_data_delayed_67__15_, chained_data_delayed_67__14_, chained_data_delayed_67__13_, chained_data_delayed_67__12_, chained_data_delayed_67__11_, chained_data_delayed_67__10_, chained_data_delayed_67__9_, chained_data_delayed_67__8_, chained_data_delayed_67__7_, chained_data_delayed_67__6_, chained_data_delayed_67__5_, chained_data_delayed_67__4_, chained_data_delayed_67__3_, chained_data_delayed_67__2_, chained_data_delayed_67__1_, chained_data_delayed_67__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_68__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_67__127_, chained_data_delayed_67__126_, chained_data_delayed_67__125_, chained_data_delayed_67__124_, chained_data_delayed_67__123_, chained_data_delayed_67__122_, chained_data_delayed_67__121_, chained_data_delayed_67__120_, chained_data_delayed_67__119_, chained_data_delayed_67__118_, chained_data_delayed_67__117_, chained_data_delayed_67__116_, chained_data_delayed_67__115_, chained_data_delayed_67__114_, chained_data_delayed_67__113_, chained_data_delayed_67__112_, chained_data_delayed_67__111_, chained_data_delayed_67__110_, chained_data_delayed_67__109_, chained_data_delayed_67__108_, chained_data_delayed_67__107_, chained_data_delayed_67__106_, chained_data_delayed_67__105_, chained_data_delayed_67__104_, chained_data_delayed_67__103_, chained_data_delayed_67__102_, chained_data_delayed_67__101_, chained_data_delayed_67__100_, chained_data_delayed_67__99_, chained_data_delayed_67__98_, chained_data_delayed_67__97_, chained_data_delayed_67__96_, chained_data_delayed_67__95_, chained_data_delayed_67__94_, chained_data_delayed_67__93_, chained_data_delayed_67__92_, chained_data_delayed_67__91_, chained_data_delayed_67__90_, chained_data_delayed_67__89_, chained_data_delayed_67__88_, chained_data_delayed_67__87_, chained_data_delayed_67__86_, chained_data_delayed_67__85_, chained_data_delayed_67__84_, chained_data_delayed_67__83_, chained_data_delayed_67__82_, chained_data_delayed_67__81_, chained_data_delayed_67__80_, chained_data_delayed_67__79_, chained_data_delayed_67__78_, chained_data_delayed_67__77_, chained_data_delayed_67__76_, chained_data_delayed_67__75_, chained_data_delayed_67__74_, chained_data_delayed_67__73_, chained_data_delayed_67__72_, chained_data_delayed_67__71_, chained_data_delayed_67__70_, chained_data_delayed_67__69_, chained_data_delayed_67__68_, chained_data_delayed_67__67_, chained_data_delayed_67__66_, chained_data_delayed_67__65_, chained_data_delayed_67__64_, chained_data_delayed_67__63_, chained_data_delayed_67__62_, chained_data_delayed_67__61_, chained_data_delayed_67__60_, chained_data_delayed_67__59_, chained_data_delayed_67__58_, chained_data_delayed_67__57_, chained_data_delayed_67__56_, chained_data_delayed_67__55_, chained_data_delayed_67__54_, chained_data_delayed_67__53_, chained_data_delayed_67__52_, chained_data_delayed_67__51_, chained_data_delayed_67__50_, chained_data_delayed_67__49_, chained_data_delayed_67__48_, chained_data_delayed_67__47_, chained_data_delayed_67__46_, chained_data_delayed_67__45_, chained_data_delayed_67__44_, chained_data_delayed_67__43_, chained_data_delayed_67__42_, chained_data_delayed_67__41_, chained_data_delayed_67__40_, chained_data_delayed_67__39_, chained_data_delayed_67__38_, chained_data_delayed_67__37_, chained_data_delayed_67__36_, chained_data_delayed_67__35_, chained_data_delayed_67__34_, chained_data_delayed_67__33_, chained_data_delayed_67__32_, chained_data_delayed_67__31_, chained_data_delayed_67__30_, chained_data_delayed_67__29_, chained_data_delayed_67__28_, chained_data_delayed_67__27_, chained_data_delayed_67__26_, chained_data_delayed_67__25_, chained_data_delayed_67__24_, chained_data_delayed_67__23_, chained_data_delayed_67__22_, chained_data_delayed_67__21_, chained_data_delayed_67__20_, chained_data_delayed_67__19_, chained_data_delayed_67__18_, chained_data_delayed_67__17_, chained_data_delayed_67__16_, chained_data_delayed_67__15_, chained_data_delayed_67__14_, chained_data_delayed_67__13_, chained_data_delayed_67__12_, chained_data_delayed_67__11_, chained_data_delayed_67__10_, chained_data_delayed_67__9_, chained_data_delayed_67__8_, chained_data_delayed_67__7_, chained_data_delayed_67__6_, chained_data_delayed_67__5_, chained_data_delayed_67__4_, chained_data_delayed_67__3_, chained_data_delayed_67__2_, chained_data_delayed_67__1_, chained_data_delayed_67__0_ }),
    .data_o({ chained_data_delayed_68__127_, chained_data_delayed_68__126_, chained_data_delayed_68__125_, chained_data_delayed_68__124_, chained_data_delayed_68__123_, chained_data_delayed_68__122_, chained_data_delayed_68__121_, chained_data_delayed_68__120_, chained_data_delayed_68__119_, chained_data_delayed_68__118_, chained_data_delayed_68__117_, chained_data_delayed_68__116_, chained_data_delayed_68__115_, chained_data_delayed_68__114_, chained_data_delayed_68__113_, chained_data_delayed_68__112_, chained_data_delayed_68__111_, chained_data_delayed_68__110_, chained_data_delayed_68__109_, chained_data_delayed_68__108_, chained_data_delayed_68__107_, chained_data_delayed_68__106_, chained_data_delayed_68__105_, chained_data_delayed_68__104_, chained_data_delayed_68__103_, chained_data_delayed_68__102_, chained_data_delayed_68__101_, chained_data_delayed_68__100_, chained_data_delayed_68__99_, chained_data_delayed_68__98_, chained_data_delayed_68__97_, chained_data_delayed_68__96_, chained_data_delayed_68__95_, chained_data_delayed_68__94_, chained_data_delayed_68__93_, chained_data_delayed_68__92_, chained_data_delayed_68__91_, chained_data_delayed_68__90_, chained_data_delayed_68__89_, chained_data_delayed_68__88_, chained_data_delayed_68__87_, chained_data_delayed_68__86_, chained_data_delayed_68__85_, chained_data_delayed_68__84_, chained_data_delayed_68__83_, chained_data_delayed_68__82_, chained_data_delayed_68__81_, chained_data_delayed_68__80_, chained_data_delayed_68__79_, chained_data_delayed_68__78_, chained_data_delayed_68__77_, chained_data_delayed_68__76_, chained_data_delayed_68__75_, chained_data_delayed_68__74_, chained_data_delayed_68__73_, chained_data_delayed_68__72_, chained_data_delayed_68__71_, chained_data_delayed_68__70_, chained_data_delayed_68__69_, chained_data_delayed_68__68_, chained_data_delayed_68__67_, chained_data_delayed_68__66_, chained_data_delayed_68__65_, chained_data_delayed_68__64_, chained_data_delayed_68__63_, chained_data_delayed_68__62_, chained_data_delayed_68__61_, chained_data_delayed_68__60_, chained_data_delayed_68__59_, chained_data_delayed_68__58_, chained_data_delayed_68__57_, chained_data_delayed_68__56_, chained_data_delayed_68__55_, chained_data_delayed_68__54_, chained_data_delayed_68__53_, chained_data_delayed_68__52_, chained_data_delayed_68__51_, chained_data_delayed_68__50_, chained_data_delayed_68__49_, chained_data_delayed_68__48_, chained_data_delayed_68__47_, chained_data_delayed_68__46_, chained_data_delayed_68__45_, chained_data_delayed_68__44_, chained_data_delayed_68__43_, chained_data_delayed_68__42_, chained_data_delayed_68__41_, chained_data_delayed_68__40_, chained_data_delayed_68__39_, chained_data_delayed_68__38_, chained_data_delayed_68__37_, chained_data_delayed_68__36_, chained_data_delayed_68__35_, chained_data_delayed_68__34_, chained_data_delayed_68__33_, chained_data_delayed_68__32_, chained_data_delayed_68__31_, chained_data_delayed_68__30_, chained_data_delayed_68__29_, chained_data_delayed_68__28_, chained_data_delayed_68__27_, chained_data_delayed_68__26_, chained_data_delayed_68__25_, chained_data_delayed_68__24_, chained_data_delayed_68__23_, chained_data_delayed_68__22_, chained_data_delayed_68__21_, chained_data_delayed_68__20_, chained_data_delayed_68__19_, chained_data_delayed_68__18_, chained_data_delayed_68__17_, chained_data_delayed_68__16_, chained_data_delayed_68__15_, chained_data_delayed_68__14_, chained_data_delayed_68__13_, chained_data_delayed_68__12_, chained_data_delayed_68__11_, chained_data_delayed_68__10_, chained_data_delayed_68__9_, chained_data_delayed_68__8_, chained_data_delayed_68__7_, chained_data_delayed_68__6_, chained_data_delayed_68__5_, chained_data_delayed_68__4_, chained_data_delayed_68__3_, chained_data_delayed_68__2_, chained_data_delayed_68__1_, chained_data_delayed_68__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_69__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_68__127_, chained_data_delayed_68__126_, chained_data_delayed_68__125_, chained_data_delayed_68__124_, chained_data_delayed_68__123_, chained_data_delayed_68__122_, chained_data_delayed_68__121_, chained_data_delayed_68__120_, chained_data_delayed_68__119_, chained_data_delayed_68__118_, chained_data_delayed_68__117_, chained_data_delayed_68__116_, chained_data_delayed_68__115_, chained_data_delayed_68__114_, chained_data_delayed_68__113_, chained_data_delayed_68__112_, chained_data_delayed_68__111_, chained_data_delayed_68__110_, chained_data_delayed_68__109_, chained_data_delayed_68__108_, chained_data_delayed_68__107_, chained_data_delayed_68__106_, chained_data_delayed_68__105_, chained_data_delayed_68__104_, chained_data_delayed_68__103_, chained_data_delayed_68__102_, chained_data_delayed_68__101_, chained_data_delayed_68__100_, chained_data_delayed_68__99_, chained_data_delayed_68__98_, chained_data_delayed_68__97_, chained_data_delayed_68__96_, chained_data_delayed_68__95_, chained_data_delayed_68__94_, chained_data_delayed_68__93_, chained_data_delayed_68__92_, chained_data_delayed_68__91_, chained_data_delayed_68__90_, chained_data_delayed_68__89_, chained_data_delayed_68__88_, chained_data_delayed_68__87_, chained_data_delayed_68__86_, chained_data_delayed_68__85_, chained_data_delayed_68__84_, chained_data_delayed_68__83_, chained_data_delayed_68__82_, chained_data_delayed_68__81_, chained_data_delayed_68__80_, chained_data_delayed_68__79_, chained_data_delayed_68__78_, chained_data_delayed_68__77_, chained_data_delayed_68__76_, chained_data_delayed_68__75_, chained_data_delayed_68__74_, chained_data_delayed_68__73_, chained_data_delayed_68__72_, chained_data_delayed_68__71_, chained_data_delayed_68__70_, chained_data_delayed_68__69_, chained_data_delayed_68__68_, chained_data_delayed_68__67_, chained_data_delayed_68__66_, chained_data_delayed_68__65_, chained_data_delayed_68__64_, chained_data_delayed_68__63_, chained_data_delayed_68__62_, chained_data_delayed_68__61_, chained_data_delayed_68__60_, chained_data_delayed_68__59_, chained_data_delayed_68__58_, chained_data_delayed_68__57_, chained_data_delayed_68__56_, chained_data_delayed_68__55_, chained_data_delayed_68__54_, chained_data_delayed_68__53_, chained_data_delayed_68__52_, chained_data_delayed_68__51_, chained_data_delayed_68__50_, chained_data_delayed_68__49_, chained_data_delayed_68__48_, chained_data_delayed_68__47_, chained_data_delayed_68__46_, chained_data_delayed_68__45_, chained_data_delayed_68__44_, chained_data_delayed_68__43_, chained_data_delayed_68__42_, chained_data_delayed_68__41_, chained_data_delayed_68__40_, chained_data_delayed_68__39_, chained_data_delayed_68__38_, chained_data_delayed_68__37_, chained_data_delayed_68__36_, chained_data_delayed_68__35_, chained_data_delayed_68__34_, chained_data_delayed_68__33_, chained_data_delayed_68__32_, chained_data_delayed_68__31_, chained_data_delayed_68__30_, chained_data_delayed_68__29_, chained_data_delayed_68__28_, chained_data_delayed_68__27_, chained_data_delayed_68__26_, chained_data_delayed_68__25_, chained_data_delayed_68__24_, chained_data_delayed_68__23_, chained_data_delayed_68__22_, chained_data_delayed_68__21_, chained_data_delayed_68__20_, chained_data_delayed_68__19_, chained_data_delayed_68__18_, chained_data_delayed_68__17_, chained_data_delayed_68__16_, chained_data_delayed_68__15_, chained_data_delayed_68__14_, chained_data_delayed_68__13_, chained_data_delayed_68__12_, chained_data_delayed_68__11_, chained_data_delayed_68__10_, chained_data_delayed_68__9_, chained_data_delayed_68__8_, chained_data_delayed_68__7_, chained_data_delayed_68__6_, chained_data_delayed_68__5_, chained_data_delayed_68__4_, chained_data_delayed_68__3_, chained_data_delayed_68__2_, chained_data_delayed_68__1_, chained_data_delayed_68__0_ }),
    .data_o({ chained_data_delayed_69__127_, chained_data_delayed_69__126_, chained_data_delayed_69__125_, chained_data_delayed_69__124_, chained_data_delayed_69__123_, chained_data_delayed_69__122_, chained_data_delayed_69__121_, chained_data_delayed_69__120_, chained_data_delayed_69__119_, chained_data_delayed_69__118_, chained_data_delayed_69__117_, chained_data_delayed_69__116_, chained_data_delayed_69__115_, chained_data_delayed_69__114_, chained_data_delayed_69__113_, chained_data_delayed_69__112_, chained_data_delayed_69__111_, chained_data_delayed_69__110_, chained_data_delayed_69__109_, chained_data_delayed_69__108_, chained_data_delayed_69__107_, chained_data_delayed_69__106_, chained_data_delayed_69__105_, chained_data_delayed_69__104_, chained_data_delayed_69__103_, chained_data_delayed_69__102_, chained_data_delayed_69__101_, chained_data_delayed_69__100_, chained_data_delayed_69__99_, chained_data_delayed_69__98_, chained_data_delayed_69__97_, chained_data_delayed_69__96_, chained_data_delayed_69__95_, chained_data_delayed_69__94_, chained_data_delayed_69__93_, chained_data_delayed_69__92_, chained_data_delayed_69__91_, chained_data_delayed_69__90_, chained_data_delayed_69__89_, chained_data_delayed_69__88_, chained_data_delayed_69__87_, chained_data_delayed_69__86_, chained_data_delayed_69__85_, chained_data_delayed_69__84_, chained_data_delayed_69__83_, chained_data_delayed_69__82_, chained_data_delayed_69__81_, chained_data_delayed_69__80_, chained_data_delayed_69__79_, chained_data_delayed_69__78_, chained_data_delayed_69__77_, chained_data_delayed_69__76_, chained_data_delayed_69__75_, chained_data_delayed_69__74_, chained_data_delayed_69__73_, chained_data_delayed_69__72_, chained_data_delayed_69__71_, chained_data_delayed_69__70_, chained_data_delayed_69__69_, chained_data_delayed_69__68_, chained_data_delayed_69__67_, chained_data_delayed_69__66_, chained_data_delayed_69__65_, chained_data_delayed_69__64_, chained_data_delayed_69__63_, chained_data_delayed_69__62_, chained_data_delayed_69__61_, chained_data_delayed_69__60_, chained_data_delayed_69__59_, chained_data_delayed_69__58_, chained_data_delayed_69__57_, chained_data_delayed_69__56_, chained_data_delayed_69__55_, chained_data_delayed_69__54_, chained_data_delayed_69__53_, chained_data_delayed_69__52_, chained_data_delayed_69__51_, chained_data_delayed_69__50_, chained_data_delayed_69__49_, chained_data_delayed_69__48_, chained_data_delayed_69__47_, chained_data_delayed_69__46_, chained_data_delayed_69__45_, chained_data_delayed_69__44_, chained_data_delayed_69__43_, chained_data_delayed_69__42_, chained_data_delayed_69__41_, chained_data_delayed_69__40_, chained_data_delayed_69__39_, chained_data_delayed_69__38_, chained_data_delayed_69__37_, chained_data_delayed_69__36_, chained_data_delayed_69__35_, chained_data_delayed_69__34_, chained_data_delayed_69__33_, chained_data_delayed_69__32_, chained_data_delayed_69__31_, chained_data_delayed_69__30_, chained_data_delayed_69__29_, chained_data_delayed_69__28_, chained_data_delayed_69__27_, chained_data_delayed_69__26_, chained_data_delayed_69__25_, chained_data_delayed_69__24_, chained_data_delayed_69__23_, chained_data_delayed_69__22_, chained_data_delayed_69__21_, chained_data_delayed_69__20_, chained_data_delayed_69__19_, chained_data_delayed_69__18_, chained_data_delayed_69__17_, chained_data_delayed_69__16_, chained_data_delayed_69__15_, chained_data_delayed_69__14_, chained_data_delayed_69__13_, chained_data_delayed_69__12_, chained_data_delayed_69__11_, chained_data_delayed_69__10_, chained_data_delayed_69__9_, chained_data_delayed_69__8_, chained_data_delayed_69__7_, chained_data_delayed_69__6_, chained_data_delayed_69__5_, chained_data_delayed_69__4_, chained_data_delayed_69__3_, chained_data_delayed_69__2_, chained_data_delayed_69__1_, chained_data_delayed_69__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_70__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_69__127_, chained_data_delayed_69__126_, chained_data_delayed_69__125_, chained_data_delayed_69__124_, chained_data_delayed_69__123_, chained_data_delayed_69__122_, chained_data_delayed_69__121_, chained_data_delayed_69__120_, chained_data_delayed_69__119_, chained_data_delayed_69__118_, chained_data_delayed_69__117_, chained_data_delayed_69__116_, chained_data_delayed_69__115_, chained_data_delayed_69__114_, chained_data_delayed_69__113_, chained_data_delayed_69__112_, chained_data_delayed_69__111_, chained_data_delayed_69__110_, chained_data_delayed_69__109_, chained_data_delayed_69__108_, chained_data_delayed_69__107_, chained_data_delayed_69__106_, chained_data_delayed_69__105_, chained_data_delayed_69__104_, chained_data_delayed_69__103_, chained_data_delayed_69__102_, chained_data_delayed_69__101_, chained_data_delayed_69__100_, chained_data_delayed_69__99_, chained_data_delayed_69__98_, chained_data_delayed_69__97_, chained_data_delayed_69__96_, chained_data_delayed_69__95_, chained_data_delayed_69__94_, chained_data_delayed_69__93_, chained_data_delayed_69__92_, chained_data_delayed_69__91_, chained_data_delayed_69__90_, chained_data_delayed_69__89_, chained_data_delayed_69__88_, chained_data_delayed_69__87_, chained_data_delayed_69__86_, chained_data_delayed_69__85_, chained_data_delayed_69__84_, chained_data_delayed_69__83_, chained_data_delayed_69__82_, chained_data_delayed_69__81_, chained_data_delayed_69__80_, chained_data_delayed_69__79_, chained_data_delayed_69__78_, chained_data_delayed_69__77_, chained_data_delayed_69__76_, chained_data_delayed_69__75_, chained_data_delayed_69__74_, chained_data_delayed_69__73_, chained_data_delayed_69__72_, chained_data_delayed_69__71_, chained_data_delayed_69__70_, chained_data_delayed_69__69_, chained_data_delayed_69__68_, chained_data_delayed_69__67_, chained_data_delayed_69__66_, chained_data_delayed_69__65_, chained_data_delayed_69__64_, chained_data_delayed_69__63_, chained_data_delayed_69__62_, chained_data_delayed_69__61_, chained_data_delayed_69__60_, chained_data_delayed_69__59_, chained_data_delayed_69__58_, chained_data_delayed_69__57_, chained_data_delayed_69__56_, chained_data_delayed_69__55_, chained_data_delayed_69__54_, chained_data_delayed_69__53_, chained_data_delayed_69__52_, chained_data_delayed_69__51_, chained_data_delayed_69__50_, chained_data_delayed_69__49_, chained_data_delayed_69__48_, chained_data_delayed_69__47_, chained_data_delayed_69__46_, chained_data_delayed_69__45_, chained_data_delayed_69__44_, chained_data_delayed_69__43_, chained_data_delayed_69__42_, chained_data_delayed_69__41_, chained_data_delayed_69__40_, chained_data_delayed_69__39_, chained_data_delayed_69__38_, chained_data_delayed_69__37_, chained_data_delayed_69__36_, chained_data_delayed_69__35_, chained_data_delayed_69__34_, chained_data_delayed_69__33_, chained_data_delayed_69__32_, chained_data_delayed_69__31_, chained_data_delayed_69__30_, chained_data_delayed_69__29_, chained_data_delayed_69__28_, chained_data_delayed_69__27_, chained_data_delayed_69__26_, chained_data_delayed_69__25_, chained_data_delayed_69__24_, chained_data_delayed_69__23_, chained_data_delayed_69__22_, chained_data_delayed_69__21_, chained_data_delayed_69__20_, chained_data_delayed_69__19_, chained_data_delayed_69__18_, chained_data_delayed_69__17_, chained_data_delayed_69__16_, chained_data_delayed_69__15_, chained_data_delayed_69__14_, chained_data_delayed_69__13_, chained_data_delayed_69__12_, chained_data_delayed_69__11_, chained_data_delayed_69__10_, chained_data_delayed_69__9_, chained_data_delayed_69__8_, chained_data_delayed_69__7_, chained_data_delayed_69__6_, chained_data_delayed_69__5_, chained_data_delayed_69__4_, chained_data_delayed_69__3_, chained_data_delayed_69__2_, chained_data_delayed_69__1_, chained_data_delayed_69__0_ }),
    .data_o({ chained_data_delayed_70__127_, chained_data_delayed_70__126_, chained_data_delayed_70__125_, chained_data_delayed_70__124_, chained_data_delayed_70__123_, chained_data_delayed_70__122_, chained_data_delayed_70__121_, chained_data_delayed_70__120_, chained_data_delayed_70__119_, chained_data_delayed_70__118_, chained_data_delayed_70__117_, chained_data_delayed_70__116_, chained_data_delayed_70__115_, chained_data_delayed_70__114_, chained_data_delayed_70__113_, chained_data_delayed_70__112_, chained_data_delayed_70__111_, chained_data_delayed_70__110_, chained_data_delayed_70__109_, chained_data_delayed_70__108_, chained_data_delayed_70__107_, chained_data_delayed_70__106_, chained_data_delayed_70__105_, chained_data_delayed_70__104_, chained_data_delayed_70__103_, chained_data_delayed_70__102_, chained_data_delayed_70__101_, chained_data_delayed_70__100_, chained_data_delayed_70__99_, chained_data_delayed_70__98_, chained_data_delayed_70__97_, chained_data_delayed_70__96_, chained_data_delayed_70__95_, chained_data_delayed_70__94_, chained_data_delayed_70__93_, chained_data_delayed_70__92_, chained_data_delayed_70__91_, chained_data_delayed_70__90_, chained_data_delayed_70__89_, chained_data_delayed_70__88_, chained_data_delayed_70__87_, chained_data_delayed_70__86_, chained_data_delayed_70__85_, chained_data_delayed_70__84_, chained_data_delayed_70__83_, chained_data_delayed_70__82_, chained_data_delayed_70__81_, chained_data_delayed_70__80_, chained_data_delayed_70__79_, chained_data_delayed_70__78_, chained_data_delayed_70__77_, chained_data_delayed_70__76_, chained_data_delayed_70__75_, chained_data_delayed_70__74_, chained_data_delayed_70__73_, chained_data_delayed_70__72_, chained_data_delayed_70__71_, chained_data_delayed_70__70_, chained_data_delayed_70__69_, chained_data_delayed_70__68_, chained_data_delayed_70__67_, chained_data_delayed_70__66_, chained_data_delayed_70__65_, chained_data_delayed_70__64_, chained_data_delayed_70__63_, chained_data_delayed_70__62_, chained_data_delayed_70__61_, chained_data_delayed_70__60_, chained_data_delayed_70__59_, chained_data_delayed_70__58_, chained_data_delayed_70__57_, chained_data_delayed_70__56_, chained_data_delayed_70__55_, chained_data_delayed_70__54_, chained_data_delayed_70__53_, chained_data_delayed_70__52_, chained_data_delayed_70__51_, chained_data_delayed_70__50_, chained_data_delayed_70__49_, chained_data_delayed_70__48_, chained_data_delayed_70__47_, chained_data_delayed_70__46_, chained_data_delayed_70__45_, chained_data_delayed_70__44_, chained_data_delayed_70__43_, chained_data_delayed_70__42_, chained_data_delayed_70__41_, chained_data_delayed_70__40_, chained_data_delayed_70__39_, chained_data_delayed_70__38_, chained_data_delayed_70__37_, chained_data_delayed_70__36_, chained_data_delayed_70__35_, chained_data_delayed_70__34_, chained_data_delayed_70__33_, chained_data_delayed_70__32_, chained_data_delayed_70__31_, chained_data_delayed_70__30_, chained_data_delayed_70__29_, chained_data_delayed_70__28_, chained_data_delayed_70__27_, chained_data_delayed_70__26_, chained_data_delayed_70__25_, chained_data_delayed_70__24_, chained_data_delayed_70__23_, chained_data_delayed_70__22_, chained_data_delayed_70__21_, chained_data_delayed_70__20_, chained_data_delayed_70__19_, chained_data_delayed_70__18_, chained_data_delayed_70__17_, chained_data_delayed_70__16_, chained_data_delayed_70__15_, chained_data_delayed_70__14_, chained_data_delayed_70__13_, chained_data_delayed_70__12_, chained_data_delayed_70__11_, chained_data_delayed_70__10_, chained_data_delayed_70__9_, chained_data_delayed_70__8_, chained_data_delayed_70__7_, chained_data_delayed_70__6_, chained_data_delayed_70__5_, chained_data_delayed_70__4_, chained_data_delayed_70__3_, chained_data_delayed_70__2_, chained_data_delayed_70__1_, chained_data_delayed_70__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_71__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_70__127_, chained_data_delayed_70__126_, chained_data_delayed_70__125_, chained_data_delayed_70__124_, chained_data_delayed_70__123_, chained_data_delayed_70__122_, chained_data_delayed_70__121_, chained_data_delayed_70__120_, chained_data_delayed_70__119_, chained_data_delayed_70__118_, chained_data_delayed_70__117_, chained_data_delayed_70__116_, chained_data_delayed_70__115_, chained_data_delayed_70__114_, chained_data_delayed_70__113_, chained_data_delayed_70__112_, chained_data_delayed_70__111_, chained_data_delayed_70__110_, chained_data_delayed_70__109_, chained_data_delayed_70__108_, chained_data_delayed_70__107_, chained_data_delayed_70__106_, chained_data_delayed_70__105_, chained_data_delayed_70__104_, chained_data_delayed_70__103_, chained_data_delayed_70__102_, chained_data_delayed_70__101_, chained_data_delayed_70__100_, chained_data_delayed_70__99_, chained_data_delayed_70__98_, chained_data_delayed_70__97_, chained_data_delayed_70__96_, chained_data_delayed_70__95_, chained_data_delayed_70__94_, chained_data_delayed_70__93_, chained_data_delayed_70__92_, chained_data_delayed_70__91_, chained_data_delayed_70__90_, chained_data_delayed_70__89_, chained_data_delayed_70__88_, chained_data_delayed_70__87_, chained_data_delayed_70__86_, chained_data_delayed_70__85_, chained_data_delayed_70__84_, chained_data_delayed_70__83_, chained_data_delayed_70__82_, chained_data_delayed_70__81_, chained_data_delayed_70__80_, chained_data_delayed_70__79_, chained_data_delayed_70__78_, chained_data_delayed_70__77_, chained_data_delayed_70__76_, chained_data_delayed_70__75_, chained_data_delayed_70__74_, chained_data_delayed_70__73_, chained_data_delayed_70__72_, chained_data_delayed_70__71_, chained_data_delayed_70__70_, chained_data_delayed_70__69_, chained_data_delayed_70__68_, chained_data_delayed_70__67_, chained_data_delayed_70__66_, chained_data_delayed_70__65_, chained_data_delayed_70__64_, chained_data_delayed_70__63_, chained_data_delayed_70__62_, chained_data_delayed_70__61_, chained_data_delayed_70__60_, chained_data_delayed_70__59_, chained_data_delayed_70__58_, chained_data_delayed_70__57_, chained_data_delayed_70__56_, chained_data_delayed_70__55_, chained_data_delayed_70__54_, chained_data_delayed_70__53_, chained_data_delayed_70__52_, chained_data_delayed_70__51_, chained_data_delayed_70__50_, chained_data_delayed_70__49_, chained_data_delayed_70__48_, chained_data_delayed_70__47_, chained_data_delayed_70__46_, chained_data_delayed_70__45_, chained_data_delayed_70__44_, chained_data_delayed_70__43_, chained_data_delayed_70__42_, chained_data_delayed_70__41_, chained_data_delayed_70__40_, chained_data_delayed_70__39_, chained_data_delayed_70__38_, chained_data_delayed_70__37_, chained_data_delayed_70__36_, chained_data_delayed_70__35_, chained_data_delayed_70__34_, chained_data_delayed_70__33_, chained_data_delayed_70__32_, chained_data_delayed_70__31_, chained_data_delayed_70__30_, chained_data_delayed_70__29_, chained_data_delayed_70__28_, chained_data_delayed_70__27_, chained_data_delayed_70__26_, chained_data_delayed_70__25_, chained_data_delayed_70__24_, chained_data_delayed_70__23_, chained_data_delayed_70__22_, chained_data_delayed_70__21_, chained_data_delayed_70__20_, chained_data_delayed_70__19_, chained_data_delayed_70__18_, chained_data_delayed_70__17_, chained_data_delayed_70__16_, chained_data_delayed_70__15_, chained_data_delayed_70__14_, chained_data_delayed_70__13_, chained_data_delayed_70__12_, chained_data_delayed_70__11_, chained_data_delayed_70__10_, chained_data_delayed_70__9_, chained_data_delayed_70__8_, chained_data_delayed_70__7_, chained_data_delayed_70__6_, chained_data_delayed_70__5_, chained_data_delayed_70__4_, chained_data_delayed_70__3_, chained_data_delayed_70__2_, chained_data_delayed_70__1_, chained_data_delayed_70__0_ }),
    .data_o({ chained_data_delayed_71__127_, chained_data_delayed_71__126_, chained_data_delayed_71__125_, chained_data_delayed_71__124_, chained_data_delayed_71__123_, chained_data_delayed_71__122_, chained_data_delayed_71__121_, chained_data_delayed_71__120_, chained_data_delayed_71__119_, chained_data_delayed_71__118_, chained_data_delayed_71__117_, chained_data_delayed_71__116_, chained_data_delayed_71__115_, chained_data_delayed_71__114_, chained_data_delayed_71__113_, chained_data_delayed_71__112_, chained_data_delayed_71__111_, chained_data_delayed_71__110_, chained_data_delayed_71__109_, chained_data_delayed_71__108_, chained_data_delayed_71__107_, chained_data_delayed_71__106_, chained_data_delayed_71__105_, chained_data_delayed_71__104_, chained_data_delayed_71__103_, chained_data_delayed_71__102_, chained_data_delayed_71__101_, chained_data_delayed_71__100_, chained_data_delayed_71__99_, chained_data_delayed_71__98_, chained_data_delayed_71__97_, chained_data_delayed_71__96_, chained_data_delayed_71__95_, chained_data_delayed_71__94_, chained_data_delayed_71__93_, chained_data_delayed_71__92_, chained_data_delayed_71__91_, chained_data_delayed_71__90_, chained_data_delayed_71__89_, chained_data_delayed_71__88_, chained_data_delayed_71__87_, chained_data_delayed_71__86_, chained_data_delayed_71__85_, chained_data_delayed_71__84_, chained_data_delayed_71__83_, chained_data_delayed_71__82_, chained_data_delayed_71__81_, chained_data_delayed_71__80_, chained_data_delayed_71__79_, chained_data_delayed_71__78_, chained_data_delayed_71__77_, chained_data_delayed_71__76_, chained_data_delayed_71__75_, chained_data_delayed_71__74_, chained_data_delayed_71__73_, chained_data_delayed_71__72_, chained_data_delayed_71__71_, chained_data_delayed_71__70_, chained_data_delayed_71__69_, chained_data_delayed_71__68_, chained_data_delayed_71__67_, chained_data_delayed_71__66_, chained_data_delayed_71__65_, chained_data_delayed_71__64_, chained_data_delayed_71__63_, chained_data_delayed_71__62_, chained_data_delayed_71__61_, chained_data_delayed_71__60_, chained_data_delayed_71__59_, chained_data_delayed_71__58_, chained_data_delayed_71__57_, chained_data_delayed_71__56_, chained_data_delayed_71__55_, chained_data_delayed_71__54_, chained_data_delayed_71__53_, chained_data_delayed_71__52_, chained_data_delayed_71__51_, chained_data_delayed_71__50_, chained_data_delayed_71__49_, chained_data_delayed_71__48_, chained_data_delayed_71__47_, chained_data_delayed_71__46_, chained_data_delayed_71__45_, chained_data_delayed_71__44_, chained_data_delayed_71__43_, chained_data_delayed_71__42_, chained_data_delayed_71__41_, chained_data_delayed_71__40_, chained_data_delayed_71__39_, chained_data_delayed_71__38_, chained_data_delayed_71__37_, chained_data_delayed_71__36_, chained_data_delayed_71__35_, chained_data_delayed_71__34_, chained_data_delayed_71__33_, chained_data_delayed_71__32_, chained_data_delayed_71__31_, chained_data_delayed_71__30_, chained_data_delayed_71__29_, chained_data_delayed_71__28_, chained_data_delayed_71__27_, chained_data_delayed_71__26_, chained_data_delayed_71__25_, chained_data_delayed_71__24_, chained_data_delayed_71__23_, chained_data_delayed_71__22_, chained_data_delayed_71__21_, chained_data_delayed_71__20_, chained_data_delayed_71__19_, chained_data_delayed_71__18_, chained_data_delayed_71__17_, chained_data_delayed_71__16_, chained_data_delayed_71__15_, chained_data_delayed_71__14_, chained_data_delayed_71__13_, chained_data_delayed_71__12_, chained_data_delayed_71__11_, chained_data_delayed_71__10_, chained_data_delayed_71__9_, chained_data_delayed_71__8_, chained_data_delayed_71__7_, chained_data_delayed_71__6_, chained_data_delayed_71__5_, chained_data_delayed_71__4_, chained_data_delayed_71__3_, chained_data_delayed_71__2_, chained_data_delayed_71__1_, chained_data_delayed_71__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_72__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_71__127_, chained_data_delayed_71__126_, chained_data_delayed_71__125_, chained_data_delayed_71__124_, chained_data_delayed_71__123_, chained_data_delayed_71__122_, chained_data_delayed_71__121_, chained_data_delayed_71__120_, chained_data_delayed_71__119_, chained_data_delayed_71__118_, chained_data_delayed_71__117_, chained_data_delayed_71__116_, chained_data_delayed_71__115_, chained_data_delayed_71__114_, chained_data_delayed_71__113_, chained_data_delayed_71__112_, chained_data_delayed_71__111_, chained_data_delayed_71__110_, chained_data_delayed_71__109_, chained_data_delayed_71__108_, chained_data_delayed_71__107_, chained_data_delayed_71__106_, chained_data_delayed_71__105_, chained_data_delayed_71__104_, chained_data_delayed_71__103_, chained_data_delayed_71__102_, chained_data_delayed_71__101_, chained_data_delayed_71__100_, chained_data_delayed_71__99_, chained_data_delayed_71__98_, chained_data_delayed_71__97_, chained_data_delayed_71__96_, chained_data_delayed_71__95_, chained_data_delayed_71__94_, chained_data_delayed_71__93_, chained_data_delayed_71__92_, chained_data_delayed_71__91_, chained_data_delayed_71__90_, chained_data_delayed_71__89_, chained_data_delayed_71__88_, chained_data_delayed_71__87_, chained_data_delayed_71__86_, chained_data_delayed_71__85_, chained_data_delayed_71__84_, chained_data_delayed_71__83_, chained_data_delayed_71__82_, chained_data_delayed_71__81_, chained_data_delayed_71__80_, chained_data_delayed_71__79_, chained_data_delayed_71__78_, chained_data_delayed_71__77_, chained_data_delayed_71__76_, chained_data_delayed_71__75_, chained_data_delayed_71__74_, chained_data_delayed_71__73_, chained_data_delayed_71__72_, chained_data_delayed_71__71_, chained_data_delayed_71__70_, chained_data_delayed_71__69_, chained_data_delayed_71__68_, chained_data_delayed_71__67_, chained_data_delayed_71__66_, chained_data_delayed_71__65_, chained_data_delayed_71__64_, chained_data_delayed_71__63_, chained_data_delayed_71__62_, chained_data_delayed_71__61_, chained_data_delayed_71__60_, chained_data_delayed_71__59_, chained_data_delayed_71__58_, chained_data_delayed_71__57_, chained_data_delayed_71__56_, chained_data_delayed_71__55_, chained_data_delayed_71__54_, chained_data_delayed_71__53_, chained_data_delayed_71__52_, chained_data_delayed_71__51_, chained_data_delayed_71__50_, chained_data_delayed_71__49_, chained_data_delayed_71__48_, chained_data_delayed_71__47_, chained_data_delayed_71__46_, chained_data_delayed_71__45_, chained_data_delayed_71__44_, chained_data_delayed_71__43_, chained_data_delayed_71__42_, chained_data_delayed_71__41_, chained_data_delayed_71__40_, chained_data_delayed_71__39_, chained_data_delayed_71__38_, chained_data_delayed_71__37_, chained_data_delayed_71__36_, chained_data_delayed_71__35_, chained_data_delayed_71__34_, chained_data_delayed_71__33_, chained_data_delayed_71__32_, chained_data_delayed_71__31_, chained_data_delayed_71__30_, chained_data_delayed_71__29_, chained_data_delayed_71__28_, chained_data_delayed_71__27_, chained_data_delayed_71__26_, chained_data_delayed_71__25_, chained_data_delayed_71__24_, chained_data_delayed_71__23_, chained_data_delayed_71__22_, chained_data_delayed_71__21_, chained_data_delayed_71__20_, chained_data_delayed_71__19_, chained_data_delayed_71__18_, chained_data_delayed_71__17_, chained_data_delayed_71__16_, chained_data_delayed_71__15_, chained_data_delayed_71__14_, chained_data_delayed_71__13_, chained_data_delayed_71__12_, chained_data_delayed_71__11_, chained_data_delayed_71__10_, chained_data_delayed_71__9_, chained_data_delayed_71__8_, chained_data_delayed_71__7_, chained_data_delayed_71__6_, chained_data_delayed_71__5_, chained_data_delayed_71__4_, chained_data_delayed_71__3_, chained_data_delayed_71__2_, chained_data_delayed_71__1_, chained_data_delayed_71__0_ }),
    .data_o({ chained_data_delayed_72__127_, chained_data_delayed_72__126_, chained_data_delayed_72__125_, chained_data_delayed_72__124_, chained_data_delayed_72__123_, chained_data_delayed_72__122_, chained_data_delayed_72__121_, chained_data_delayed_72__120_, chained_data_delayed_72__119_, chained_data_delayed_72__118_, chained_data_delayed_72__117_, chained_data_delayed_72__116_, chained_data_delayed_72__115_, chained_data_delayed_72__114_, chained_data_delayed_72__113_, chained_data_delayed_72__112_, chained_data_delayed_72__111_, chained_data_delayed_72__110_, chained_data_delayed_72__109_, chained_data_delayed_72__108_, chained_data_delayed_72__107_, chained_data_delayed_72__106_, chained_data_delayed_72__105_, chained_data_delayed_72__104_, chained_data_delayed_72__103_, chained_data_delayed_72__102_, chained_data_delayed_72__101_, chained_data_delayed_72__100_, chained_data_delayed_72__99_, chained_data_delayed_72__98_, chained_data_delayed_72__97_, chained_data_delayed_72__96_, chained_data_delayed_72__95_, chained_data_delayed_72__94_, chained_data_delayed_72__93_, chained_data_delayed_72__92_, chained_data_delayed_72__91_, chained_data_delayed_72__90_, chained_data_delayed_72__89_, chained_data_delayed_72__88_, chained_data_delayed_72__87_, chained_data_delayed_72__86_, chained_data_delayed_72__85_, chained_data_delayed_72__84_, chained_data_delayed_72__83_, chained_data_delayed_72__82_, chained_data_delayed_72__81_, chained_data_delayed_72__80_, chained_data_delayed_72__79_, chained_data_delayed_72__78_, chained_data_delayed_72__77_, chained_data_delayed_72__76_, chained_data_delayed_72__75_, chained_data_delayed_72__74_, chained_data_delayed_72__73_, chained_data_delayed_72__72_, chained_data_delayed_72__71_, chained_data_delayed_72__70_, chained_data_delayed_72__69_, chained_data_delayed_72__68_, chained_data_delayed_72__67_, chained_data_delayed_72__66_, chained_data_delayed_72__65_, chained_data_delayed_72__64_, chained_data_delayed_72__63_, chained_data_delayed_72__62_, chained_data_delayed_72__61_, chained_data_delayed_72__60_, chained_data_delayed_72__59_, chained_data_delayed_72__58_, chained_data_delayed_72__57_, chained_data_delayed_72__56_, chained_data_delayed_72__55_, chained_data_delayed_72__54_, chained_data_delayed_72__53_, chained_data_delayed_72__52_, chained_data_delayed_72__51_, chained_data_delayed_72__50_, chained_data_delayed_72__49_, chained_data_delayed_72__48_, chained_data_delayed_72__47_, chained_data_delayed_72__46_, chained_data_delayed_72__45_, chained_data_delayed_72__44_, chained_data_delayed_72__43_, chained_data_delayed_72__42_, chained_data_delayed_72__41_, chained_data_delayed_72__40_, chained_data_delayed_72__39_, chained_data_delayed_72__38_, chained_data_delayed_72__37_, chained_data_delayed_72__36_, chained_data_delayed_72__35_, chained_data_delayed_72__34_, chained_data_delayed_72__33_, chained_data_delayed_72__32_, chained_data_delayed_72__31_, chained_data_delayed_72__30_, chained_data_delayed_72__29_, chained_data_delayed_72__28_, chained_data_delayed_72__27_, chained_data_delayed_72__26_, chained_data_delayed_72__25_, chained_data_delayed_72__24_, chained_data_delayed_72__23_, chained_data_delayed_72__22_, chained_data_delayed_72__21_, chained_data_delayed_72__20_, chained_data_delayed_72__19_, chained_data_delayed_72__18_, chained_data_delayed_72__17_, chained_data_delayed_72__16_, chained_data_delayed_72__15_, chained_data_delayed_72__14_, chained_data_delayed_72__13_, chained_data_delayed_72__12_, chained_data_delayed_72__11_, chained_data_delayed_72__10_, chained_data_delayed_72__9_, chained_data_delayed_72__8_, chained_data_delayed_72__7_, chained_data_delayed_72__6_, chained_data_delayed_72__5_, chained_data_delayed_72__4_, chained_data_delayed_72__3_, chained_data_delayed_72__2_, chained_data_delayed_72__1_, chained_data_delayed_72__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_73__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_72__127_, chained_data_delayed_72__126_, chained_data_delayed_72__125_, chained_data_delayed_72__124_, chained_data_delayed_72__123_, chained_data_delayed_72__122_, chained_data_delayed_72__121_, chained_data_delayed_72__120_, chained_data_delayed_72__119_, chained_data_delayed_72__118_, chained_data_delayed_72__117_, chained_data_delayed_72__116_, chained_data_delayed_72__115_, chained_data_delayed_72__114_, chained_data_delayed_72__113_, chained_data_delayed_72__112_, chained_data_delayed_72__111_, chained_data_delayed_72__110_, chained_data_delayed_72__109_, chained_data_delayed_72__108_, chained_data_delayed_72__107_, chained_data_delayed_72__106_, chained_data_delayed_72__105_, chained_data_delayed_72__104_, chained_data_delayed_72__103_, chained_data_delayed_72__102_, chained_data_delayed_72__101_, chained_data_delayed_72__100_, chained_data_delayed_72__99_, chained_data_delayed_72__98_, chained_data_delayed_72__97_, chained_data_delayed_72__96_, chained_data_delayed_72__95_, chained_data_delayed_72__94_, chained_data_delayed_72__93_, chained_data_delayed_72__92_, chained_data_delayed_72__91_, chained_data_delayed_72__90_, chained_data_delayed_72__89_, chained_data_delayed_72__88_, chained_data_delayed_72__87_, chained_data_delayed_72__86_, chained_data_delayed_72__85_, chained_data_delayed_72__84_, chained_data_delayed_72__83_, chained_data_delayed_72__82_, chained_data_delayed_72__81_, chained_data_delayed_72__80_, chained_data_delayed_72__79_, chained_data_delayed_72__78_, chained_data_delayed_72__77_, chained_data_delayed_72__76_, chained_data_delayed_72__75_, chained_data_delayed_72__74_, chained_data_delayed_72__73_, chained_data_delayed_72__72_, chained_data_delayed_72__71_, chained_data_delayed_72__70_, chained_data_delayed_72__69_, chained_data_delayed_72__68_, chained_data_delayed_72__67_, chained_data_delayed_72__66_, chained_data_delayed_72__65_, chained_data_delayed_72__64_, chained_data_delayed_72__63_, chained_data_delayed_72__62_, chained_data_delayed_72__61_, chained_data_delayed_72__60_, chained_data_delayed_72__59_, chained_data_delayed_72__58_, chained_data_delayed_72__57_, chained_data_delayed_72__56_, chained_data_delayed_72__55_, chained_data_delayed_72__54_, chained_data_delayed_72__53_, chained_data_delayed_72__52_, chained_data_delayed_72__51_, chained_data_delayed_72__50_, chained_data_delayed_72__49_, chained_data_delayed_72__48_, chained_data_delayed_72__47_, chained_data_delayed_72__46_, chained_data_delayed_72__45_, chained_data_delayed_72__44_, chained_data_delayed_72__43_, chained_data_delayed_72__42_, chained_data_delayed_72__41_, chained_data_delayed_72__40_, chained_data_delayed_72__39_, chained_data_delayed_72__38_, chained_data_delayed_72__37_, chained_data_delayed_72__36_, chained_data_delayed_72__35_, chained_data_delayed_72__34_, chained_data_delayed_72__33_, chained_data_delayed_72__32_, chained_data_delayed_72__31_, chained_data_delayed_72__30_, chained_data_delayed_72__29_, chained_data_delayed_72__28_, chained_data_delayed_72__27_, chained_data_delayed_72__26_, chained_data_delayed_72__25_, chained_data_delayed_72__24_, chained_data_delayed_72__23_, chained_data_delayed_72__22_, chained_data_delayed_72__21_, chained_data_delayed_72__20_, chained_data_delayed_72__19_, chained_data_delayed_72__18_, chained_data_delayed_72__17_, chained_data_delayed_72__16_, chained_data_delayed_72__15_, chained_data_delayed_72__14_, chained_data_delayed_72__13_, chained_data_delayed_72__12_, chained_data_delayed_72__11_, chained_data_delayed_72__10_, chained_data_delayed_72__9_, chained_data_delayed_72__8_, chained_data_delayed_72__7_, chained_data_delayed_72__6_, chained_data_delayed_72__5_, chained_data_delayed_72__4_, chained_data_delayed_72__3_, chained_data_delayed_72__2_, chained_data_delayed_72__1_, chained_data_delayed_72__0_ }),
    .data_o({ chained_data_delayed_73__127_, chained_data_delayed_73__126_, chained_data_delayed_73__125_, chained_data_delayed_73__124_, chained_data_delayed_73__123_, chained_data_delayed_73__122_, chained_data_delayed_73__121_, chained_data_delayed_73__120_, chained_data_delayed_73__119_, chained_data_delayed_73__118_, chained_data_delayed_73__117_, chained_data_delayed_73__116_, chained_data_delayed_73__115_, chained_data_delayed_73__114_, chained_data_delayed_73__113_, chained_data_delayed_73__112_, chained_data_delayed_73__111_, chained_data_delayed_73__110_, chained_data_delayed_73__109_, chained_data_delayed_73__108_, chained_data_delayed_73__107_, chained_data_delayed_73__106_, chained_data_delayed_73__105_, chained_data_delayed_73__104_, chained_data_delayed_73__103_, chained_data_delayed_73__102_, chained_data_delayed_73__101_, chained_data_delayed_73__100_, chained_data_delayed_73__99_, chained_data_delayed_73__98_, chained_data_delayed_73__97_, chained_data_delayed_73__96_, chained_data_delayed_73__95_, chained_data_delayed_73__94_, chained_data_delayed_73__93_, chained_data_delayed_73__92_, chained_data_delayed_73__91_, chained_data_delayed_73__90_, chained_data_delayed_73__89_, chained_data_delayed_73__88_, chained_data_delayed_73__87_, chained_data_delayed_73__86_, chained_data_delayed_73__85_, chained_data_delayed_73__84_, chained_data_delayed_73__83_, chained_data_delayed_73__82_, chained_data_delayed_73__81_, chained_data_delayed_73__80_, chained_data_delayed_73__79_, chained_data_delayed_73__78_, chained_data_delayed_73__77_, chained_data_delayed_73__76_, chained_data_delayed_73__75_, chained_data_delayed_73__74_, chained_data_delayed_73__73_, chained_data_delayed_73__72_, chained_data_delayed_73__71_, chained_data_delayed_73__70_, chained_data_delayed_73__69_, chained_data_delayed_73__68_, chained_data_delayed_73__67_, chained_data_delayed_73__66_, chained_data_delayed_73__65_, chained_data_delayed_73__64_, chained_data_delayed_73__63_, chained_data_delayed_73__62_, chained_data_delayed_73__61_, chained_data_delayed_73__60_, chained_data_delayed_73__59_, chained_data_delayed_73__58_, chained_data_delayed_73__57_, chained_data_delayed_73__56_, chained_data_delayed_73__55_, chained_data_delayed_73__54_, chained_data_delayed_73__53_, chained_data_delayed_73__52_, chained_data_delayed_73__51_, chained_data_delayed_73__50_, chained_data_delayed_73__49_, chained_data_delayed_73__48_, chained_data_delayed_73__47_, chained_data_delayed_73__46_, chained_data_delayed_73__45_, chained_data_delayed_73__44_, chained_data_delayed_73__43_, chained_data_delayed_73__42_, chained_data_delayed_73__41_, chained_data_delayed_73__40_, chained_data_delayed_73__39_, chained_data_delayed_73__38_, chained_data_delayed_73__37_, chained_data_delayed_73__36_, chained_data_delayed_73__35_, chained_data_delayed_73__34_, chained_data_delayed_73__33_, chained_data_delayed_73__32_, chained_data_delayed_73__31_, chained_data_delayed_73__30_, chained_data_delayed_73__29_, chained_data_delayed_73__28_, chained_data_delayed_73__27_, chained_data_delayed_73__26_, chained_data_delayed_73__25_, chained_data_delayed_73__24_, chained_data_delayed_73__23_, chained_data_delayed_73__22_, chained_data_delayed_73__21_, chained_data_delayed_73__20_, chained_data_delayed_73__19_, chained_data_delayed_73__18_, chained_data_delayed_73__17_, chained_data_delayed_73__16_, chained_data_delayed_73__15_, chained_data_delayed_73__14_, chained_data_delayed_73__13_, chained_data_delayed_73__12_, chained_data_delayed_73__11_, chained_data_delayed_73__10_, chained_data_delayed_73__9_, chained_data_delayed_73__8_, chained_data_delayed_73__7_, chained_data_delayed_73__6_, chained_data_delayed_73__5_, chained_data_delayed_73__4_, chained_data_delayed_73__3_, chained_data_delayed_73__2_, chained_data_delayed_73__1_, chained_data_delayed_73__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_74__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_73__127_, chained_data_delayed_73__126_, chained_data_delayed_73__125_, chained_data_delayed_73__124_, chained_data_delayed_73__123_, chained_data_delayed_73__122_, chained_data_delayed_73__121_, chained_data_delayed_73__120_, chained_data_delayed_73__119_, chained_data_delayed_73__118_, chained_data_delayed_73__117_, chained_data_delayed_73__116_, chained_data_delayed_73__115_, chained_data_delayed_73__114_, chained_data_delayed_73__113_, chained_data_delayed_73__112_, chained_data_delayed_73__111_, chained_data_delayed_73__110_, chained_data_delayed_73__109_, chained_data_delayed_73__108_, chained_data_delayed_73__107_, chained_data_delayed_73__106_, chained_data_delayed_73__105_, chained_data_delayed_73__104_, chained_data_delayed_73__103_, chained_data_delayed_73__102_, chained_data_delayed_73__101_, chained_data_delayed_73__100_, chained_data_delayed_73__99_, chained_data_delayed_73__98_, chained_data_delayed_73__97_, chained_data_delayed_73__96_, chained_data_delayed_73__95_, chained_data_delayed_73__94_, chained_data_delayed_73__93_, chained_data_delayed_73__92_, chained_data_delayed_73__91_, chained_data_delayed_73__90_, chained_data_delayed_73__89_, chained_data_delayed_73__88_, chained_data_delayed_73__87_, chained_data_delayed_73__86_, chained_data_delayed_73__85_, chained_data_delayed_73__84_, chained_data_delayed_73__83_, chained_data_delayed_73__82_, chained_data_delayed_73__81_, chained_data_delayed_73__80_, chained_data_delayed_73__79_, chained_data_delayed_73__78_, chained_data_delayed_73__77_, chained_data_delayed_73__76_, chained_data_delayed_73__75_, chained_data_delayed_73__74_, chained_data_delayed_73__73_, chained_data_delayed_73__72_, chained_data_delayed_73__71_, chained_data_delayed_73__70_, chained_data_delayed_73__69_, chained_data_delayed_73__68_, chained_data_delayed_73__67_, chained_data_delayed_73__66_, chained_data_delayed_73__65_, chained_data_delayed_73__64_, chained_data_delayed_73__63_, chained_data_delayed_73__62_, chained_data_delayed_73__61_, chained_data_delayed_73__60_, chained_data_delayed_73__59_, chained_data_delayed_73__58_, chained_data_delayed_73__57_, chained_data_delayed_73__56_, chained_data_delayed_73__55_, chained_data_delayed_73__54_, chained_data_delayed_73__53_, chained_data_delayed_73__52_, chained_data_delayed_73__51_, chained_data_delayed_73__50_, chained_data_delayed_73__49_, chained_data_delayed_73__48_, chained_data_delayed_73__47_, chained_data_delayed_73__46_, chained_data_delayed_73__45_, chained_data_delayed_73__44_, chained_data_delayed_73__43_, chained_data_delayed_73__42_, chained_data_delayed_73__41_, chained_data_delayed_73__40_, chained_data_delayed_73__39_, chained_data_delayed_73__38_, chained_data_delayed_73__37_, chained_data_delayed_73__36_, chained_data_delayed_73__35_, chained_data_delayed_73__34_, chained_data_delayed_73__33_, chained_data_delayed_73__32_, chained_data_delayed_73__31_, chained_data_delayed_73__30_, chained_data_delayed_73__29_, chained_data_delayed_73__28_, chained_data_delayed_73__27_, chained_data_delayed_73__26_, chained_data_delayed_73__25_, chained_data_delayed_73__24_, chained_data_delayed_73__23_, chained_data_delayed_73__22_, chained_data_delayed_73__21_, chained_data_delayed_73__20_, chained_data_delayed_73__19_, chained_data_delayed_73__18_, chained_data_delayed_73__17_, chained_data_delayed_73__16_, chained_data_delayed_73__15_, chained_data_delayed_73__14_, chained_data_delayed_73__13_, chained_data_delayed_73__12_, chained_data_delayed_73__11_, chained_data_delayed_73__10_, chained_data_delayed_73__9_, chained_data_delayed_73__8_, chained_data_delayed_73__7_, chained_data_delayed_73__6_, chained_data_delayed_73__5_, chained_data_delayed_73__4_, chained_data_delayed_73__3_, chained_data_delayed_73__2_, chained_data_delayed_73__1_, chained_data_delayed_73__0_ }),
    .data_o({ chained_data_delayed_74__127_, chained_data_delayed_74__126_, chained_data_delayed_74__125_, chained_data_delayed_74__124_, chained_data_delayed_74__123_, chained_data_delayed_74__122_, chained_data_delayed_74__121_, chained_data_delayed_74__120_, chained_data_delayed_74__119_, chained_data_delayed_74__118_, chained_data_delayed_74__117_, chained_data_delayed_74__116_, chained_data_delayed_74__115_, chained_data_delayed_74__114_, chained_data_delayed_74__113_, chained_data_delayed_74__112_, chained_data_delayed_74__111_, chained_data_delayed_74__110_, chained_data_delayed_74__109_, chained_data_delayed_74__108_, chained_data_delayed_74__107_, chained_data_delayed_74__106_, chained_data_delayed_74__105_, chained_data_delayed_74__104_, chained_data_delayed_74__103_, chained_data_delayed_74__102_, chained_data_delayed_74__101_, chained_data_delayed_74__100_, chained_data_delayed_74__99_, chained_data_delayed_74__98_, chained_data_delayed_74__97_, chained_data_delayed_74__96_, chained_data_delayed_74__95_, chained_data_delayed_74__94_, chained_data_delayed_74__93_, chained_data_delayed_74__92_, chained_data_delayed_74__91_, chained_data_delayed_74__90_, chained_data_delayed_74__89_, chained_data_delayed_74__88_, chained_data_delayed_74__87_, chained_data_delayed_74__86_, chained_data_delayed_74__85_, chained_data_delayed_74__84_, chained_data_delayed_74__83_, chained_data_delayed_74__82_, chained_data_delayed_74__81_, chained_data_delayed_74__80_, chained_data_delayed_74__79_, chained_data_delayed_74__78_, chained_data_delayed_74__77_, chained_data_delayed_74__76_, chained_data_delayed_74__75_, chained_data_delayed_74__74_, chained_data_delayed_74__73_, chained_data_delayed_74__72_, chained_data_delayed_74__71_, chained_data_delayed_74__70_, chained_data_delayed_74__69_, chained_data_delayed_74__68_, chained_data_delayed_74__67_, chained_data_delayed_74__66_, chained_data_delayed_74__65_, chained_data_delayed_74__64_, chained_data_delayed_74__63_, chained_data_delayed_74__62_, chained_data_delayed_74__61_, chained_data_delayed_74__60_, chained_data_delayed_74__59_, chained_data_delayed_74__58_, chained_data_delayed_74__57_, chained_data_delayed_74__56_, chained_data_delayed_74__55_, chained_data_delayed_74__54_, chained_data_delayed_74__53_, chained_data_delayed_74__52_, chained_data_delayed_74__51_, chained_data_delayed_74__50_, chained_data_delayed_74__49_, chained_data_delayed_74__48_, chained_data_delayed_74__47_, chained_data_delayed_74__46_, chained_data_delayed_74__45_, chained_data_delayed_74__44_, chained_data_delayed_74__43_, chained_data_delayed_74__42_, chained_data_delayed_74__41_, chained_data_delayed_74__40_, chained_data_delayed_74__39_, chained_data_delayed_74__38_, chained_data_delayed_74__37_, chained_data_delayed_74__36_, chained_data_delayed_74__35_, chained_data_delayed_74__34_, chained_data_delayed_74__33_, chained_data_delayed_74__32_, chained_data_delayed_74__31_, chained_data_delayed_74__30_, chained_data_delayed_74__29_, chained_data_delayed_74__28_, chained_data_delayed_74__27_, chained_data_delayed_74__26_, chained_data_delayed_74__25_, chained_data_delayed_74__24_, chained_data_delayed_74__23_, chained_data_delayed_74__22_, chained_data_delayed_74__21_, chained_data_delayed_74__20_, chained_data_delayed_74__19_, chained_data_delayed_74__18_, chained_data_delayed_74__17_, chained_data_delayed_74__16_, chained_data_delayed_74__15_, chained_data_delayed_74__14_, chained_data_delayed_74__13_, chained_data_delayed_74__12_, chained_data_delayed_74__11_, chained_data_delayed_74__10_, chained_data_delayed_74__9_, chained_data_delayed_74__8_, chained_data_delayed_74__7_, chained_data_delayed_74__6_, chained_data_delayed_74__5_, chained_data_delayed_74__4_, chained_data_delayed_74__3_, chained_data_delayed_74__2_, chained_data_delayed_74__1_, chained_data_delayed_74__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_75__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_74__127_, chained_data_delayed_74__126_, chained_data_delayed_74__125_, chained_data_delayed_74__124_, chained_data_delayed_74__123_, chained_data_delayed_74__122_, chained_data_delayed_74__121_, chained_data_delayed_74__120_, chained_data_delayed_74__119_, chained_data_delayed_74__118_, chained_data_delayed_74__117_, chained_data_delayed_74__116_, chained_data_delayed_74__115_, chained_data_delayed_74__114_, chained_data_delayed_74__113_, chained_data_delayed_74__112_, chained_data_delayed_74__111_, chained_data_delayed_74__110_, chained_data_delayed_74__109_, chained_data_delayed_74__108_, chained_data_delayed_74__107_, chained_data_delayed_74__106_, chained_data_delayed_74__105_, chained_data_delayed_74__104_, chained_data_delayed_74__103_, chained_data_delayed_74__102_, chained_data_delayed_74__101_, chained_data_delayed_74__100_, chained_data_delayed_74__99_, chained_data_delayed_74__98_, chained_data_delayed_74__97_, chained_data_delayed_74__96_, chained_data_delayed_74__95_, chained_data_delayed_74__94_, chained_data_delayed_74__93_, chained_data_delayed_74__92_, chained_data_delayed_74__91_, chained_data_delayed_74__90_, chained_data_delayed_74__89_, chained_data_delayed_74__88_, chained_data_delayed_74__87_, chained_data_delayed_74__86_, chained_data_delayed_74__85_, chained_data_delayed_74__84_, chained_data_delayed_74__83_, chained_data_delayed_74__82_, chained_data_delayed_74__81_, chained_data_delayed_74__80_, chained_data_delayed_74__79_, chained_data_delayed_74__78_, chained_data_delayed_74__77_, chained_data_delayed_74__76_, chained_data_delayed_74__75_, chained_data_delayed_74__74_, chained_data_delayed_74__73_, chained_data_delayed_74__72_, chained_data_delayed_74__71_, chained_data_delayed_74__70_, chained_data_delayed_74__69_, chained_data_delayed_74__68_, chained_data_delayed_74__67_, chained_data_delayed_74__66_, chained_data_delayed_74__65_, chained_data_delayed_74__64_, chained_data_delayed_74__63_, chained_data_delayed_74__62_, chained_data_delayed_74__61_, chained_data_delayed_74__60_, chained_data_delayed_74__59_, chained_data_delayed_74__58_, chained_data_delayed_74__57_, chained_data_delayed_74__56_, chained_data_delayed_74__55_, chained_data_delayed_74__54_, chained_data_delayed_74__53_, chained_data_delayed_74__52_, chained_data_delayed_74__51_, chained_data_delayed_74__50_, chained_data_delayed_74__49_, chained_data_delayed_74__48_, chained_data_delayed_74__47_, chained_data_delayed_74__46_, chained_data_delayed_74__45_, chained_data_delayed_74__44_, chained_data_delayed_74__43_, chained_data_delayed_74__42_, chained_data_delayed_74__41_, chained_data_delayed_74__40_, chained_data_delayed_74__39_, chained_data_delayed_74__38_, chained_data_delayed_74__37_, chained_data_delayed_74__36_, chained_data_delayed_74__35_, chained_data_delayed_74__34_, chained_data_delayed_74__33_, chained_data_delayed_74__32_, chained_data_delayed_74__31_, chained_data_delayed_74__30_, chained_data_delayed_74__29_, chained_data_delayed_74__28_, chained_data_delayed_74__27_, chained_data_delayed_74__26_, chained_data_delayed_74__25_, chained_data_delayed_74__24_, chained_data_delayed_74__23_, chained_data_delayed_74__22_, chained_data_delayed_74__21_, chained_data_delayed_74__20_, chained_data_delayed_74__19_, chained_data_delayed_74__18_, chained_data_delayed_74__17_, chained_data_delayed_74__16_, chained_data_delayed_74__15_, chained_data_delayed_74__14_, chained_data_delayed_74__13_, chained_data_delayed_74__12_, chained_data_delayed_74__11_, chained_data_delayed_74__10_, chained_data_delayed_74__9_, chained_data_delayed_74__8_, chained_data_delayed_74__7_, chained_data_delayed_74__6_, chained_data_delayed_74__5_, chained_data_delayed_74__4_, chained_data_delayed_74__3_, chained_data_delayed_74__2_, chained_data_delayed_74__1_, chained_data_delayed_74__0_ }),
    .data_o({ chained_data_delayed_75__127_, chained_data_delayed_75__126_, chained_data_delayed_75__125_, chained_data_delayed_75__124_, chained_data_delayed_75__123_, chained_data_delayed_75__122_, chained_data_delayed_75__121_, chained_data_delayed_75__120_, chained_data_delayed_75__119_, chained_data_delayed_75__118_, chained_data_delayed_75__117_, chained_data_delayed_75__116_, chained_data_delayed_75__115_, chained_data_delayed_75__114_, chained_data_delayed_75__113_, chained_data_delayed_75__112_, chained_data_delayed_75__111_, chained_data_delayed_75__110_, chained_data_delayed_75__109_, chained_data_delayed_75__108_, chained_data_delayed_75__107_, chained_data_delayed_75__106_, chained_data_delayed_75__105_, chained_data_delayed_75__104_, chained_data_delayed_75__103_, chained_data_delayed_75__102_, chained_data_delayed_75__101_, chained_data_delayed_75__100_, chained_data_delayed_75__99_, chained_data_delayed_75__98_, chained_data_delayed_75__97_, chained_data_delayed_75__96_, chained_data_delayed_75__95_, chained_data_delayed_75__94_, chained_data_delayed_75__93_, chained_data_delayed_75__92_, chained_data_delayed_75__91_, chained_data_delayed_75__90_, chained_data_delayed_75__89_, chained_data_delayed_75__88_, chained_data_delayed_75__87_, chained_data_delayed_75__86_, chained_data_delayed_75__85_, chained_data_delayed_75__84_, chained_data_delayed_75__83_, chained_data_delayed_75__82_, chained_data_delayed_75__81_, chained_data_delayed_75__80_, chained_data_delayed_75__79_, chained_data_delayed_75__78_, chained_data_delayed_75__77_, chained_data_delayed_75__76_, chained_data_delayed_75__75_, chained_data_delayed_75__74_, chained_data_delayed_75__73_, chained_data_delayed_75__72_, chained_data_delayed_75__71_, chained_data_delayed_75__70_, chained_data_delayed_75__69_, chained_data_delayed_75__68_, chained_data_delayed_75__67_, chained_data_delayed_75__66_, chained_data_delayed_75__65_, chained_data_delayed_75__64_, chained_data_delayed_75__63_, chained_data_delayed_75__62_, chained_data_delayed_75__61_, chained_data_delayed_75__60_, chained_data_delayed_75__59_, chained_data_delayed_75__58_, chained_data_delayed_75__57_, chained_data_delayed_75__56_, chained_data_delayed_75__55_, chained_data_delayed_75__54_, chained_data_delayed_75__53_, chained_data_delayed_75__52_, chained_data_delayed_75__51_, chained_data_delayed_75__50_, chained_data_delayed_75__49_, chained_data_delayed_75__48_, chained_data_delayed_75__47_, chained_data_delayed_75__46_, chained_data_delayed_75__45_, chained_data_delayed_75__44_, chained_data_delayed_75__43_, chained_data_delayed_75__42_, chained_data_delayed_75__41_, chained_data_delayed_75__40_, chained_data_delayed_75__39_, chained_data_delayed_75__38_, chained_data_delayed_75__37_, chained_data_delayed_75__36_, chained_data_delayed_75__35_, chained_data_delayed_75__34_, chained_data_delayed_75__33_, chained_data_delayed_75__32_, chained_data_delayed_75__31_, chained_data_delayed_75__30_, chained_data_delayed_75__29_, chained_data_delayed_75__28_, chained_data_delayed_75__27_, chained_data_delayed_75__26_, chained_data_delayed_75__25_, chained_data_delayed_75__24_, chained_data_delayed_75__23_, chained_data_delayed_75__22_, chained_data_delayed_75__21_, chained_data_delayed_75__20_, chained_data_delayed_75__19_, chained_data_delayed_75__18_, chained_data_delayed_75__17_, chained_data_delayed_75__16_, chained_data_delayed_75__15_, chained_data_delayed_75__14_, chained_data_delayed_75__13_, chained_data_delayed_75__12_, chained_data_delayed_75__11_, chained_data_delayed_75__10_, chained_data_delayed_75__9_, chained_data_delayed_75__8_, chained_data_delayed_75__7_, chained_data_delayed_75__6_, chained_data_delayed_75__5_, chained_data_delayed_75__4_, chained_data_delayed_75__3_, chained_data_delayed_75__2_, chained_data_delayed_75__1_, chained_data_delayed_75__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_76__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_75__127_, chained_data_delayed_75__126_, chained_data_delayed_75__125_, chained_data_delayed_75__124_, chained_data_delayed_75__123_, chained_data_delayed_75__122_, chained_data_delayed_75__121_, chained_data_delayed_75__120_, chained_data_delayed_75__119_, chained_data_delayed_75__118_, chained_data_delayed_75__117_, chained_data_delayed_75__116_, chained_data_delayed_75__115_, chained_data_delayed_75__114_, chained_data_delayed_75__113_, chained_data_delayed_75__112_, chained_data_delayed_75__111_, chained_data_delayed_75__110_, chained_data_delayed_75__109_, chained_data_delayed_75__108_, chained_data_delayed_75__107_, chained_data_delayed_75__106_, chained_data_delayed_75__105_, chained_data_delayed_75__104_, chained_data_delayed_75__103_, chained_data_delayed_75__102_, chained_data_delayed_75__101_, chained_data_delayed_75__100_, chained_data_delayed_75__99_, chained_data_delayed_75__98_, chained_data_delayed_75__97_, chained_data_delayed_75__96_, chained_data_delayed_75__95_, chained_data_delayed_75__94_, chained_data_delayed_75__93_, chained_data_delayed_75__92_, chained_data_delayed_75__91_, chained_data_delayed_75__90_, chained_data_delayed_75__89_, chained_data_delayed_75__88_, chained_data_delayed_75__87_, chained_data_delayed_75__86_, chained_data_delayed_75__85_, chained_data_delayed_75__84_, chained_data_delayed_75__83_, chained_data_delayed_75__82_, chained_data_delayed_75__81_, chained_data_delayed_75__80_, chained_data_delayed_75__79_, chained_data_delayed_75__78_, chained_data_delayed_75__77_, chained_data_delayed_75__76_, chained_data_delayed_75__75_, chained_data_delayed_75__74_, chained_data_delayed_75__73_, chained_data_delayed_75__72_, chained_data_delayed_75__71_, chained_data_delayed_75__70_, chained_data_delayed_75__69_, chained_data_delayed_75__68_, chained_data_delayed_75__67_, chained_data_delayed_75__66_, chained_data_delayed_75__65_, chained_data_delayed_75__64_, chained_data_delayed_75__63_, chained_data_delayed_75__62_, chained_data_delayed_75__61_, chained_data_delayed_75__60_, chained_data_delayed_75__59_, chained_data_delayed_75__58_, chained_data_delayed_75__57_, chained_data_delayed_75__56_, chained_data_delayed_75__55_, chained_data_delayed_75__54_, chained_data_delayed_75__53_, chained_data_delayed_75__52_, chained_data_delayed_75__51_, chained_data_delayed_75__50_, chained_data_delayed_75__49_, chained_data_delayed_75__48_, chained_data_delayed_75__47_, chained_data_delayed_75__46_, chained_data_delayed_75__45_, chained_data_delayed_75__44_, chained_data_delayed_75__43_, chained_data_delayed_75__42_, chained_data_delayed_75__41_, chained_data_delayed_75__40_, chained_data_delayed_75__39_, chained_data_delayed_75__38_, chained_data_delayed_75__37_, chained_data_delayed_75__36_, chained_data_delayed_75__35_, chained_data_delayed_75__34_, chained_data_delayed_75__33_, chained_data_delayed_75__32_, chained_data_delayed_75__31_, chained_data_delayed_75__30_, chained_data_delayed_75__29_, chained_data_delayed_75__28_, chained_data_delayed_75__27_, chained_data_delayed_75__26_, chained_data_delayed_75__25_, chained_data_delayed_75__24_, chained_data_delayed_75__23_, chained_data_delayed_75__22_, chained_data_delayed_75__21_, chained_data_delayed_75__20_, chained_data_delayed_75__19_, chained_data_delayed_75__18_, chained_data_delayed_75__17_, chained_data_delayed_75__16_, chained_data_delayed_75__15_, chained_data_delayed_75__14_, chained_data_delayed_75__13_, chained_data_delayed_75__12_, chained_data_delayed_75__11_, chained_data_delayed_75__10_, chained_data_delayed_75__9_, chained_data_delayed_75__8_, chained_data_delayed_75__7_, chained_data_delayed_75__6_, chained_data_delayed_75__5_, chained_data_delayed_75__4_, chained_data_delayed_75__3_, chained_data_delayed_75__2_, chained_data_delayed_75__1_, chained_data_delayed_75__0_ }),
    .data_o({ chained_data_delayed_76__127_, chained_data_delayed_76__126_, chained_data_delayed_76__125_, chained_data_delayed_76__124_, chained_data_delayed_76__123_, chained_data_delayed_76__122_, chained_data_delayed_76__121_, chained_data_delayed_76__120_, chained_data_delayed_76__119_, chained_data_delayed_76__118_, chained_data_delayed_76__117_, chained_data_delayed_76__116_, chained_data_delayed_76__115_, chained_data_delayed_76__114_, chained_data_delayed_76__113_, chained_data_delayed_76__112_, chained_data_delayed_76__111_, chained_data_delayed_76__110_, chained_data_delayed_76__109_, chained_data_delayed_76__108_, chained_data_delayed_76__107_, chained_data_delayed_76__106_, chained_data_delayed_76__105_, chained_data_delayed_76__104_, chained_data_delayed_76__103_, chained_data_delayed_76__102_, chained_data_delayed_76__101_, chained_data_delayed_76__100_, chained_data_delayed_76__99_, chained_data_delayed_76__98_, chained_data_delayed_76__97_, chained_data_delayed_76__96_, chained_data_delayed_76__95_, chained_data_delayed_76__94_, chained_data_delayed_76__93_, chained_data_delayed_76__92_, chained_data_delayed_76__91_, chained_data_delayed_76__90_, chained_data_delayed_76__89_, chained_data_delayed_76__88_, chained_data_delayed_76__87_, chained_data_delayed_76__86_, chained_data_delayed_76__85_, chained_data_delayed_76__84_, chained_data_delayed_76__83_, chained_data_delayed_76__82_, chained_data_delayed_76__81_, chained_data_delayed_76__80_, chained_data_delayed_76__79_, chained_data_delayed_76__78_, chained_data_delayed_76__77_, chained_data_delayed_76__76_, chained_data_delayed_76__75_, chained_data_delayed_76__74_, chained_data_delayed_76__73_, chained_data_delayed_76__72_, chained_data_delayed_76__71_, chained_data_delayed_76__70_, chained_data_delayed_76__69_, chained_data_delayed_76__68_, chained_data_delayed_76__67_, chained_data_delayed_76__66_, chained_data_delayed_76__65_, chained_data_delayed_76__64_, chained_data_delayed_76__63_, chained_data_delayed_76__62_, chained_data_delayed_76__61_, chained_data_delayed_76__60_, chained_data_delayed_76__59_, chained_data_delayed_76__58_, chained_data_delayed_76__57_, chained_data_delayed_76__56_, chained_data_delayed_76__55_, chained_data_delayed_76__54_, chained_data_delayed_76__53_, chained_data_delayed_76__52_, chained_data_delayed_76__51_, chained_data_delayed_76__50_, chained_data_delayed_76__49_, chained_data_delayed_76__48_, chained_data_delayed_76__47_, chained_data_delayed_76__46_, chained_data_delayed_76__45_, chained_data_delayed_76__44_, chained_data_delayed_76__43_, chained_data_delayed_76__42_, chained_data_delayed_76__41_, chained_data_delayed_76__40_, chained_data_delayed_76__39_, chained_data_delayed_76__38_, chained_data_delayed_76__37_, chained_data_delayed_76__36_, chained_data_delayed_76__35_, chained_data_delayed_76__34_, chained_data_delayed_76__33_, chained_data_delayed_76__32_, chained_data_delayed_76__31_, chained_data_delayed_76__30_, chained_data_delayed_76__29_, chained_data_delayed_76__28_, chained_data_delayed_76__27_, chained_data_delayed_76__26_, chained_data_delayed_76__25_, chained_data_delayed_76__24_, chained_data_delayed_76__23_, chained_data_delayed_76__22_, chained_data_delayed_76__21_, chained_data_delayed_76__20_, chained_data_delayed_76__19_, chained_data_delayed_76__18_, chained_data_delayed_76__17_, chained_data_delayed_76__16_, chained_data_delayed_76__15_, chained_data_delayed_76__14_, chained_data_delayed_76__13_, chained_data_delayed_76__12_, chained_data_delayed_76__11_, chained_data_delayed_76__10_, chained_data_delayed_76__9_, chained_data_delayed_76__8_, chained_data_delayed_76__7_, chained_data_delayed_76__6_, chained_data_delayed_76__5_, chained_data_delayed_76__4_, chained_data_delayed_76__3_, chained_data_delayed_76__2_, chained_data_delayed_76__1_, chained_data_delayed_76__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_77__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_76__127_, chained_data_delayed_76__126_, chained_data_delayed_76__125_, chained_data_delayed_76__124_, chained_data_delayed_76__123_, chained_data_delayed_76__122_, chained_data_delayed_76__121_, chained_data_delayed_76__120_, chained_data_delayed_76__119_, chained_data_delayed_76__118_, chained_data_delayed_76__117_, chained_data_delayed_76__116_, chained_data_delayed_76__115_, chained_data_delayed_76__114_, chained_data_delayed_76__113_, chained_data_delayed_76__112_, chained_data_delayed_76__111_, chained_data_delayed_76__110_, chained_data_delayed_76__109_, chained_data_delayed_76__108_, chained_data_delayed_76__107_, chained_data_delayed_76__106_, chained_data_delayed_76__105_, chained_data_delayed_76__104_, chained_data_delayed_76__103_, chained_data_delayed_76__102_, chained_data_delayed_76__101_, chained_data_delayed_76__100_, chained_data_delayed_76__99_, chained_data_delayed_76__98_, chained_data_delayed_76__97_, chained_data_delayed_76__96_, chained_data_delayed_76__95_, chained_data_delayed_76__94_, chained_data_delayed_76__93_, chained_data_delayed_76__92_, chained_data_delayed_76__91_, chained_data_delayed_76__90_, chained_data_delayed_76__89_, chained_data_delayed_76__88_, chained_data_delayed_76__87_, chained_data_delayed_76__86_, chained_data_delayed_76__85_, chained_data_delayed_76__84_, chained_data_delayed_76__83_, chained_data_delayed_76__82_, chained_data_delayed_76__81_, chained_data_delayed_76__80_, chained_data_delayed_76__79_, chained_data_delayed_76__78_, chained_data_delayed_76__77_, chained_data_delayed_76__76_, chained_data_delayed_76__75_, chained_data_delayed_76__74_, chained_data_delayed_76__73_, chained_data_delayed_76__72_, chained_data_delayed_76__71_, chained_data_delayed_76__70_, chained_data_delayed_76__69_, chained_data_delayed_76__68_, chained_data_delayed_76__67_, chained_data_delayed_76__66_, chained_data_delayed_76__65_, chained_data_delayed_76__64_, chained_data_delayed_76__63_, chained_data_delayed_76__62_, chained_data_delayed_76__61_, chained_data_delayed_76__60_, chained_data_delayed_76__59_, chained_data_delayed_76__58_, chained_data_delayed_76__57_, chained_data_delayed_76__56_, chained_data_delayed_76__55_, chained_data_delayed_76__54_, chained_data_delayed_76__53_, chained_data_delayed_76__52_, chained_data_delayed_76__51_, chained_data_delayed_76__50_, chained_data_delayed_76__49_, chained_data_delayed_76__48_, chained_data_delayed_76__47_, chained_data_delayed_76__46_, chained_data_delayed_76__45_, chained_data_delayed_76__44_, chained_data_delayed_76__43_, chained_data_delayed_76__42_, chained_data_delayed_76__41_, chained_data_delayed_76__40_, chained_data_delayed_76__39_, chained_data_delayed_76__38_, chained_data_delayed_76__37_, chained_data_delayed_76__36_, chained_data_delayed_76__35_, chained_data_delayed_76__34_, chained_data_delayed_76__33_, chained_data_delayed_76__32_, chained_data_delayed_76__31_, chained_data_delayed_76__30_, chained_data_delayed_76__29_, chained_data_delayed_76__28_, chained_data_delayed_76__27_, chained_data_delayed_76__26_, chained_data_delayed_76__25_, chained_data_delayed_76__24_, chained_data_delayed_76__23_, chained_data_delayed_76__22_, chained_data_delayed_76__21_, chained_data_delayed_76__20_, chained_data_delayed_76__19_, chained_data_delayed_76__18_, chained_data_delayed_76__17_, chained_data_delayed_76__16_, chained_data_delayed_76__15_, chained_data_delayed_76__14_, chained_data_delayed_76__13_, chained_data_delayed_76__12_, chained_data_delayed_76__11_, chained_data_delayed_76__10_, chained_data_delayed_76__9_, chained_data_delayed_76__8_, chained_data_delayed_76__7_, chained_data_delayed_76__6_, chained_data_delayed_76__5_, chained_data_delayed_76__4_, chained_data_delayed_76__3_, chained_data_delayed_76__2_, chained_data_delayed_76__1_, chained_data_delayed_76__0_ }),
    .data_o({ chained_data_delayed_77__127_, chained_data_delayed_77__126_, chained_data_delayed_77__125_, chained_data_delayed_77__124_, chained_data_delayed_77__123_, chained_data_delayed_77__122_, chained_data_delayed_77__121_, chained_data_delayed_77__120_, chained_data_delayed_77__119_, chained_data_delayed_77__118_, chained_data_delayed_77__117_, chained_data_delayed_77__116_, chained_data_delayed_77__115_, chained_data_delayed_77__114_, chained_data_delayed_77__113_, chained_data_delayed_77__112_, chained_data_delayed_77__111_, chained_data_delayed_77__110_, chained_data_delayed_77__109_, chained_data_delayed_77__108_, chained_data_delayed_77__107_, chained_data_delayed_77__106_, chained_data_delayed_77__105_, chained_data_delayed_77__104_, chained_data_delayed_77__103_, chained_data_delayed_77__102_, chained_data_delayed_77__101_, chained_data_delayed_77__100_, chained_data_delayed_77__99_, chained_data_delayed_77__98_, chained_data_delayed_77__97_, chained_data_delayed_77__96_, chained_data_delayed_77__95_, chained_data_delayed_77__94_, chained_data_delayed_77__93_, chained_data_delayed_77__92_, chained_data_delayed_77__91_, chained_data_delayed_77__90_, chained_data_delayed_77__89_, chained_data_delayed_77__88_, chained_data_delayed_77__87_, chained_data_delayed_77__86_, chained_data_delayed_77__85_, chained_data_delayed_77__84_, chained_data_delayed_77__83_, chained_data_delayed_77__82_, chained_data_delayed_77__81_, chained_data_delayed_77__80_, chained_data_delayed_77__79_, chained_data_delayed_77__78_, chained_data_delayed_77__77_, chained_data_delayed_77__76_, chained_data_delayed_77__75_, chained_data_delayed_77__74_, chained_data_delayed_77__73_, chained_data_delayed_77__72_, chained_data_delayed_77__71_, chained_data_delayed_77__70_, chained_data_delayed_77__69_, chained_data_delayed_77__68_, chained_data_delayed_77__67_, chained_data_delayed_77__66_, chained_data_delayed_77__65_, chained_data_delayed_77__64_, chained_data_delayed_77__63_, chained_data_delayed_77__62_, chained_data_delayed_77__61_, chained_data_delayed_77__60_, chained_data_delayed_77__59_, chained_data_delayed_77__58_, chained_data_delayed_77__57_, chained_data_delayed_77__56_, chained_data_delayed_77__55_, chained_data_delayed_77__54_, chained_data_delayed_77__53_, chained_data_delayed_77__52_, chained_data_delayed_77__51_, chained_data_delayed_77__50_, chained_data_delayed_77__49_, chained_data_delayed_77__48_, chained_data_delayed_77__47_, chained_data_delayed_77__46_, chained_data_delayed_77__45_, chained_data_delayed_77__44_, chained_data_delayed_77__43_, chained_data_delayed_77__42_, chained_data_delayed_77__41_, chained_data_delayed_77__40_, chained_data_delayed_77__39_, chained_data_delayed_77__38_, chained_data_delayed_77__37_, chained_data_delayed_77__36_, chained_data_delayed_77__35_, chained_data_delayed_77__34_, chained_data_delayed_77__33_, chained_data_delayed_77__32_, chained_data_delayed_77__31_, chained_data_delayed_77__30_, chained_data_delayed_77__29_, chained_data_delayed_77__28_, chained_data_delayed_77__27_, chained_data_delayed_77__26_, chained_data_delayed_77__25_, chained_data_delayed_77__24_, chained_data_delayed_77__23_, chained_data_delayed_77__22_, chained_data_delayed_77__21_, chained_data_delayed_77__20_, chained_data_delayed_77__19_, chained_data_delayed_77__18_, chained_data_delayed_77__17_, chained_data_delayed_77__16_, chained_data_delayed_77__15_, chained_data_delayed_77__14_, chained_data_delayed_77__13_, chained_data_delayed_77__12_, chained_data_delayed_77__11_, chained_data_delayed_77__10_, chained_data_delayed_77__9_, chained_data_delayed_77__8_, chained_data_delayed_77__7_, chained_data_delayed_77__6_, chained_data_delayed_77__5_, chained_data_delayed_77__4_, chained_data_delayed_77__3_, chained_data_delayed_77__2_, chained_data_delayed_77__1_, chained_data_delayed_77__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_78__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_77__127_, chained_data_delayed_77__126_, chained_data_delayed_77__125_, chained_data_delayed_77__124_, chained_data_delayed_77__123_, chained_data_delayed_77__122_, chained_data_delayed_77__121_, chained_data_delayed_77__120_, chained_data_delayed_77__119_, chained_data_delayed_77__118_, chained_data_delayed_77__117_, chained_data_delayed_77__116_, chained_data_delayed_77__115_, chained_data_delayed_77__114_, chained_data_delayed_77__113_, chained_data_delayed_77__112_, chained_data_delayed_77__111_, chained_data_delayed_77__110_, chained_data_delayed_77__109_, chained_data_delayed_77__108_, chained_data_delayed_77__107_, chained_data_delayed_77__106_, chained_data_delayed_77__105_, chained_data_delayed_77__104_, chained_data_delayed_77__103_, chained_data_delayed_77__102_, chained_data_delayed_77__101_, chained_data_delayed_77__100_, chained_data_delayed_77__99_, chained_data_delayed_77__98_, chained_data_delayed_77__97_, chained_data_delayed_77__96_, chained_data_delayed_77__95_, chained_data_delayed_77__94_, chained_data_delayed_77__93_, chained_data_delayed_77__92_, chained_data_delayed_77__91_, chained_data_delayed_77__90_, chained_data_delayed_77__89_, chained_data_delayed_77__88_, chained_data_delayed_77__87_, chained_data_delayed_77__86_, chained_data_delayed_77__85_, chained_data_delayed_77__84_, chained_data_delayed_77__83_, chained_data_delayed_77__82_, chained_data_delayed_77__81_, chained_data_delayed_77__80_, chained_data_delayed_77__79_, chained_data_delayed_77__78_, chained_data_delayed_77__77_, chained_data_delayed_77__76_, chained_data_delayed_77__75_, chained_data_delayed_77__74_, chained_data_delayed_77__73_, chained_data_delayed_77__72_, chained_data_delayed_77__71_, chained_data_delayed_77__70_, chained_data_delayed_77__69_, chained_data_delayed_77__68_, chained_data_delayed_77__67_, chained_data_delayed_77__66_, chained_data_delayed_77__65_, chained_data_delayed_77__64_, chained_data_delayed_77__63_, chained_data_delayed_77__62_, chained_data_delayed_77__61_, chained_data_delayed_77__60_, chained_data_delayed_77__59_, chained_data_delayed_77__58_, chained_data_delayed_77__57_, chained_data_delayed_77__56_, chained_data_delayed_77__55_, chained_data_delayed_77__54_, chained_data_delayed_77__53_, chained_data_delayed_77__52_, chained_data_delayed_77__51_, chained_data_delayed_77__50_, chained_data_delayed_77__49_, chained_data_delayed_77__48_, chained_data_delayed_77__47_, chained_data_delayed_77__46_, chained_data_delayed_77__45_, chained_data_delayed_77__44_, chained_data_delayed_77__43_, chained_data_delayed_77__42_, chained_data_delayed_77__41_, chained_data_delayed_77__40_, chained_data_delayed_77__39_, chained_data_delayed_77__38_, chained_data_delayed_77__37_, chained_data_delayed_77__36_, chained_data_delayed_77__35_, chained_data_delayed_77__34_, chained_data_delayed_77__33_, chained_data_delayed_77__32_, chained_data_delayed_77__31_, chained_data_delayed_77__30_, chained_data_delayed_77__29_, chained_data_delayed_77__28_, chained_data_delayed_77__27_, chained_data_delayed_77__26_, chained_data_delayed_77__25_, chained_data_delayed_77__24_, chained_data_delayed_77__23_, chained_data_delayed_77__22_, chained_data_delayed_77__21_, chained_data_delayed_77__20_, chained_data_delayed_77__19_, chained_data_delayed_77__18_, chained_data_delayed_77__17_, chained_data_delayed_77__16_, chained_data_delayed_77__15_, chained_data_delayed_77__14_, chained_data_delayed_77__13_, chained_data_delayed_77__12_, chained_data_delayed_77__11_, chained_data_delayed_77__10_, chained_data_delayed_77__9_, chained_data_delayed_77__8_, chained_data_delayed_77__7_, chained_data_delayed_77__6_, chained_data_delayed_77__5_, chained_data_delayed_77__4_, chained_data_delayed_77__3_, chained_data_delayed_77__2_, chained_data_delayed_77__1_, chained_data_delayed_77__0_ }),
    .data_o({ chained_data_delayed_78__127_, chained_data_delayed_78__126_, chained_data_delayed_78__125_, chained_data_delayed_78__124_, chained_data_delayed_78__123_, chained_data_delayed_78__122_, chained_data_delayed_78__121_, chained_data_delayed_78__120_, chained_data_delayed_78__119_, chained_data_delayed_78__118_, chained_data_delayed_78__117_, chained_data_delayed_78__116_, chained_data_delayed_78__115_, chained_data_delayed_78__114_, chained_data_delayed_78__113_, chained_data_delayed_78__112_, chained_data_delayed_78__111_, chained_data_delayed_78__110_, chained_data_delayed_78__109_, chained_data_delayed_78__108_, chained_data_delayed_78__107_, chained_data_delayed_78__106_, chained_data_delayed_78__105_, chained_data_delayed_78__104_, chained_data_delayed_78__103_, chained_data_delayed_78__102_, chained_data_delayed_78__101_, chained_data_delayed_78__100_, chained_data_delayed_78__99_, chained_data_delayed_78__98_, chained_data_delayed_78__97_, chained_data_delayed_78__96_, chained_data_delayed_78__95_, chained_data_delayed_78__94_, chained_data_delayed_78__93_, chained_data_delayed_78__92_, chained_data_delayed_78__91_, chained_data_delayed_78__90_, chained_data_delayed_78__89_, chained_data_delayed_78__88_, chained_data_delayed_78__87_, chained_data_delayed_78__86_, chained_data_delayed_78__85_, chained_data_delayed_78__84_, chained_data_delayed_78__83_, chained_data_delayed_78__82_, chained_data_delayed_78__81_, chained_data_delayed_78__80_, chained_data_delayed_78__79_, chained_data_delayed_78__78_, chained_data_delayed_78__77_, chained_data_delayed_78__76_, chained_data_delayed_78__75_, chained_data_delayed_78__74_, chained_data_delayed_78__73_, chained_data_delayed_78__72_, chained_data_delayed_78__71_, chained_data_delayed_78__70_, chained_data_delayed_78__69_, chained_data_delayed_78__68_, chained_data_delayed_78__67_, chained_data_delayed_78__66_, chained_data_delayed_78__65_, chained_data_delayed_78__64_, chained_data_delayed_78__63_, chained_data_delayed_78__62_, chained_data_delayed_78__61_, chained_data_delayed_78__60_, chained_data_delayed_78__59_, chained_data_delayed_78__58_, chained_data_delayed_78__57_, chained_data_delayed_78__56_, chained_data_delayed_78__55_, chained_data_delayed_78__54_, chained_data_delayed_78__53_, chained_data_delayed_78__52_, chained_data_delayed_78__51_, chained_data_delayed_78__50_, chained_data_delayed_78__49_, chained_data_delayed_78__48_, chained_data_delayed_78__47_, chained_data_delayed_78__46_, chained_data_delayed_78__45_, chained_data_delayed_78__44_, chained_data_delayed_78__43_, chained_data_delayed_78__42_, chained_data_delayed_78__41_, chained_data_delayed_78__40_, chained_data_delayed_78__39_, chained_data_delayed_78__38_, chained_data_delayed_78__37_, chained_data_delayed_78__36_, chained_data_delayed_78__35_, chained_data_delayed_78__34_, chained_data_delayed_78__33_, chained_data_delayed_78__32_, chained_data_delayed_78__31_, chained_data_delayed_78__30_, chained_data_delayed_78__29_, chained_data_delayed_78__28_, chained_data_delayed_78__27_, chained_data_delayed_78__26_, chained_data_delayed_78__25_, chained_data_delayed_78__24_, chained_data_delayed_78__23_, chained_data_delayed_78__22_, chained_data_delayed_78__21_, chained_data_delayed_78__20_, chained_data_delayed_78__19_, chained_data_delayed_78__18_, chained_data_delayed_78__17_, chained_data_delayed_78__16_, chained_data_delayed_78__15_, chained_data_delayed_78__14_, chained_data_delayed_78__13_, chained_data_delayed_78__12_, chained_data_delayed_78__11_, chained_data_delayed_78__10_, chained_data_delayed_78__9_, chained_data_delayed_78__8_, chained_data_delayed_78__7_, chained_data_delayed_78__6_, chained_data_delayed_78__5_, chained_data_delayed_78__4_, chained_data_delayed_78__3_, chained_data_delayed_78__2_, chained_data_delayed_78__1_, chained_data_delayed_78__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_79__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_78__127_, chained_data_delayed_78__126_, chained_data_delayed_78__125_, chained_data_delayed_78__124_, chained_data_delayed_78__123_, chained_data_delayed_78__122_, chained_data_delayed_78__121_, chained_data_delayed_78__120_, chained_data_delayed_78__119_, chained_data_delayed_78__118_, chained_data_delayed_78__117_, chained_data_delayed_78__116_, chained_data_delayed_78__115_, chained_data_delayed_78__114_, chained_data_delayed_78__113_, chained_data_delayed_78__112_, chained_data_delayed_78__111_, chained_data_delayed_78__110_, chained_data_delayed_78__109_, chained_data_delayed_78__108_, chained_data_delayed_78__107_, chained_data_delayed_78__106_, chained_data_delayed_78__105_, chained_data_delayed_78__104_, chained_data_delayed_78__103_, chained_data_delayed_78__102_, chained_data_delayed_78__101_, chained_data_delayed_78__100_, chained_data_delayed_78__99_, chained_data_delayed_78__98_, chained_data_delayed_78__97_, chained_data_delayed_78__96_, chained_data_delayed_78__95_, chained_data_delayed_78__94_, chained_data_delayed_78__93_, chained_data_delayed_78__92_, chained_data_delayed_78__91_, chained_data_delayed_78__90_, chained_data_delayed_78__89_, chained_data_delayed_78__88_, chained_data_delayed_78__87_, chained_data_delayed_78__86_, chained_data_delayed_78__85_, chained_data_delayed_78__84_, chained_data_delayed_78__83_, chained_data_delayed_78__82_, chained_data_delayed_78__81_, chained_data_delayed_78__80_, chained_data_delayed_78__79_, chained_data_delayed_78__78_, chained_data_delayed_78__77_, chained_data_delayed_78__76_, chained_data_delayed_78__75_, chained_data_delayed_78__74_, chained_data_delayed_78__73_, chained_data_delayed_78__72_, chained_data_delayed_78__71_, chained_data_delayed_78__70_, chained_data_delayed_78__69_, chained_data_delayed_78__68_, chained_data_delayed_78__67_, chained_data_delayed_78__66_, chained_data_delayed_78__65_, chained_data_delayed_78__64_, chained_data_delayed_78__63_, chained_data_delayed_78__62_, chained_data_delayed_78__61_, chained_data_delayed_78__60_, chained_data_delayed_78__59_, chained_data_delayed_78__58_, chained_data_delayed_78__57_, chained_data_delayed_78__56_, chained_data_delayed_78__55_, chained_data_delayed_78__54_, chained_data_delayed_78__53_, chained_data_delayed_78__52_, chained_data_delayed_78__51_, chained_data_delayed_78__50_, chained_data_delayed_78__49_, chained_data_delayed_78__48_, chained_data_delayed_78__47_, chained_data_delayed_78__46_, chained_data_delayed_78__45_, chained_data_delayed_78__44_, chained_data_delayed_78__43_, chained_data_delayed_78__42_, chained_data_delayed_78__41_, chained_data_delayed_78__40_, chained_data_delayed_78__39_, chained_data_delayed_78__38_, chained_data_delayed_78__37_, chained_data_delayed_78__36_, chained_data_delayed_78__35_, chained_data_delayed_78__34_, chained_data_delayed_78__33_, chained_data_delayed_78__32_, chained_data_delayed_78__31_, chained_data_delayed_78__30_, chained_data_delayed_78__29_, chained_data_delayed_78__28_, chained_data_delayed_78__27_, chained_data_delayed_78__26_, chained_data_delayed_78__25_, chained_data_delayed_78__24_, chained_data_delayed_78__23_, chained_data_delayed_78__22_, chained_data_delayed_78__21_, chained_data_delayed_78__20_, chained_data_delayed_78__19_, chained_data_delayed_78__18_, chained_data_delayed_78__17_, chained_data_delayed_78__16_, chained_data_delayed_78__15_, chained_data_delayed_78__14_, chained_data_delayed_78__13_, chained_data_delayed_78__12_, chained_data_delayed_78__11_, chained_data_delayed_78__10_, chained_data_delayed_78__9_, chained_data_delayed_78__8_, chained_data_delayed_78__7_, chained_data_delayed_78__6_, chained_data_delayed_78__5_, chained_data_delayed_78__4_, chained_data_delayed_78__3_, chained_data_delayed_78__2_, chained_data_delayed_78__1_, chained_data_delayed_78__0_ }),
    .data_o({ chained_data_delayed_79__127_, chained_data_delayed_79__126_, chained_data_delayed_79__125_, chained_data_delayed_79__124_, chained_data_delayed_79__123_, chained_data_delayed_79__122_, chained_data_delayed_79__121_, chained_data_delayed_79__120_, chained_data_delayed_79__119_, chained_data_delayed_79__118_, chained_data_delayed_79__117_, chained_data_delayed_79__116_, chained_data_delayed_79__115_, chained_data_delayed_79__114_, chained_data_delayed_79__113_, chained_data_delayed_79__112_, chained_data_delayed_79__111_, chained_data_delayed_79__110_, chained_data_delayed_79__109_, chained_data_delayed_79__108_, chained_data_delayed_79__107_, chained_data_delayed_79__106_, chained_data_delayed_79__105_, chained_data_delayed_79__104_, chained_data_delayed_79__103_, chained_data_delayed_79__102_, chained_data_delayed_79__101_, chained_data_delayed_79__100_, chained_data_delayed_79__99_, chained_data_delayed_79__98_, chained_data_delayed_79__97_, chained_data_delayed_79__96_, chained_data_delayed_79__95_, chained_data_delayed_79__94_, chained_data_delayed_79__93_, chained_data_delayed_79__92_, chained_data_delayed_79__91_, chained_data_delayed_79__90_, chained_data_delayed_79__89_, chained_data_delayed_79__88_, chained_data_delayed_79__87_, chained_data_delayed_79__86_, chained_data_delayed_79__85_, chained_data_delayed_79__84_, chained_data_delayed_79__83_, chained_data_delayed_79__82_, chained_data_delayed_79__81_, chained_data_delayed_79__80_, chained_data_delayed_79__79_, chained_data_delayed_79__78_, chained_data_delayed_79__77_, chained_data_delayed_79__76_, chained_data_delayed_79__75_, chained_data_delayed_79__74_, chained_data_delayed_79__73_, chained_data_delayed_79__72_, chained_data_delayed_79__71_, chained_data_delayed_79__70_, chained_data_delayed_79__69_, chained_data_delayed_79__68_, chained_data_delayed_79__67_, chained_data_delayed_79__66_, chained_data_delayed_79__65_, chained_data_delayed_79__64_, chained_data_delayed_79__63_, chained_data_delayed_79__62_, chained_data_delayed_79__61_, chained_data_delayed_79__60_, chained_data_delayed_79__59_, chained_data_delayed_79__58_, chained_data_delayed_79__57_, chained_data_delayed_79__56_, chained_data_delayed_79__55_, chained_data_delayed_79__54_, chained_data_delayed_79__53_, chained_data_delayed_79__52_, chained_data_delayed_79__51_, chained_data_delayed_79__50_, chained_data_delayed_79__49_, chained_data_delayed_79__48_, chained_data_delayed_79__47_, chained_data_delayed_79__46_, chained_data_delayed_79__45_, chained_data_delayed_79__44_, chained_data_delayed_79__43_, chained_data_delayed_79__42_, chained_data_delayed_79__41_, chained_data_delayed_79__40_, chained_data_delayed_79__39_, chained_data_delayed_79__38_, chained_data_delayed_79__37_, chained_data_delayed_79__36_, chained_data_delayed_79__35_, chained_data_delayed_79__34_, chained_data_delayed_79__33_, chained_data_delayed_79__32_, chained_data_delayed_79__31_, chained_data_delayed_79__30_, chained_data_delayed_79__29_, chained_data_delayed_79__28_, chained_data_delayed_79__27_, chained_data_delayed_79__26_, chained_data_delayed_79__25_, chained_data_delayed_79__24_, chained_data_delayed_79__23_, chained_data_delayed_79__22_, chained_data_delayed_79__21_, chained_data_delayed_79__20_, chained_data_delayed_79__19_, chained_data_delayed_79__18_, chained_data_delayed_79__17_, chained_data_delayed_79__16_, chained_data_delayed_79__15_, chained_data_delayed_79__14_, chained_data_delayed_79__13_, chained_data_delayed_79__12_, chained_data_delayed_79__11_, chained_data_delayed_79__10_, chained_data_delayed_79__9_, chained_data_delayed_79__8_, chained_data_delayed_79__7_, chained_data_delayed_79__6_, chained_data_delayed_79__5_, chained_data_delayed_79__4_, chained_data_delayed_79__3_, chained_data_delayed_79__2_, chained_data_delayed_79__1_, chained_data_delayed_79__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_80__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_79__127_, chained_data_delayed_79__126_, chained_data_delayed_79__125_, chained_data_delayed_79__124_, chained_data_delayed_79__123_, chained_data_delayed_79__122_, chained_data_delayed_79__121_, chained_data_delayed_79__120_, chained_data_delayed_79__119_, chained_data_delayed_79__118_, chained_data_delayed_79__117_, chained_data_delayed_79__116_, chained_data_delayed_79__115_, chained_data_delayed_79__114_, chained_data_delayed_79__113_, chained_data_delayed_79__112_, chained_data_delayed_79__111_, chained_data_delayed_79__110_, chained_data_delayed_79__109_, chained_data_delayed_79__108_, chained_data_delayed_79__107_, chained_data_delayed_79__106_, chained_data_delayed_79__105_, chained_data_delayed_79__104_, chained_data_delayed_79__103_, chained_data_delayed_79__102_, chained_data_delayed_79__101_, chained_data_delayed_79__100_, chained_data_delayed_79__99_, chained_data_delayed_79__98_, chained_data_delayed_79__97_, chained_data_delayed_79__96_, chained_data_delayed_79__95_, chained_data_delayed_79__94_, chained_data_delayed_79__93_, chained_data_delayed_79__92_, chained_data_delayed_79__91_, chained_data_delayed_79__90_, chained_data_delayed_79__89_, chained_data_delayed_79__88_, chained_data_delayed_79__87_, chained_data_delayed_79__86_, chained_data_delayed_79__85_, chained_data_delayed_79__84_, chained_data_delayed_79__83_, chained_data_delayed_79__82_, chained_data_delayed_79__81_, chained_data_delayed_79__80_, chained_data_delayed_79__79_, chained_data_delayed_79__78_, chained_data_delayed_79__77_, chained_data_delayed_79__76_, chained_data_delayed_79__75_, chained_data_delayed_79__74_, chained_data_delayed_79__73_, chained_data_delayed_79__72_, chained_data_delayed_79__71_, chained_data_delayed_79__70_, chained_data_delayed_79__69_, chained_data_delayed_79__68_, chained_data_delayed_79__67_, chained_data_delayed_79__66_, chained_data_delayed_79__65_, chained_data_delayed_79__64_, chained_data_delayed_79__63_, chained_data_delayed_79__62_, chained_data_delayed_79__61_, chained_data_delayed_79__60_, chained_data_delayed_79__59_, chained_data_delayed_79__58_, chained_data_delayed_79__57_, chained_data_delayed_79__56_, chained_data_delayed_79__55_, chained_data_delayed_79__54_, chained_data_delayed_79__53_, chained_data_delayed_79__52_, chained_data_delayed_79__51_, chained_data_delayed_79__50_, chained_data_delayed_79__49_, chained_data_delayed_79__48_, chained_data_delayed_79__47_, chained_data_delayed_79__46_, chained_data_delayed_79__45_, chained_data_delayed_79__44_, chained_data_delayed_79__43_, chained_data_delayed_79__42_, chained_data_delayed_79__41_, chained_data_delayed_79__40_, chained_data_delayed_79__39_, chained_data_delayed_79__38_, chained_data_delayed_79__37_, chained_data_delayed_79__36_, chained_data_delayed_79__35_, chained_data_delayed_79__34_, chained_data_delayed_79__33_, chained_data_delayed_79__32_, chained_data_delayed_79__31_, chained_data_delayed_79__30_, chained_data_delayed_79__29_, chained_data_delayed_79__28_, chained_data_delayed_79__27_, chained_data_delayed_79__26_, chained_data_delayed_79__25_, chained_data_delayed_79__24_, chained_data_delayed_79__23_, chained_data_delayed_79__22_, chained_data_delayed_79__21_, chained_data_delayed_79__20_, chained_data_delayed_79__19_, chained_data_delayed_79__18_, chained_data_delayed_79__17_, chained_data_delayed_79__16_, chained_data_delayed_79__15_, chained_data_delayed_79__14_, chained_data_delayed_79__13_, chained_data_delayed_79__12_, chained_data_delayed_79__11_, chained_data_delayed_79__10_, chained_data_delayed_79__9_, chained_data_delayed_79__8_, chained_data_delayed_79__7_, chained_data_delayed_79__6_, chained_data_delayed_79__5_, chained_data_delayed_79__4_, chained_data_delayed_79__3_, chained_data_delayed_79__2_, chained_data_delayed_79__1_, chained_data_delayed_79__0_ }),
    .data_o({ chained_data_delayed_80__127_, chained_data_delayed_80__126_, chained_data_delayed_80__125_, chained_data_delayed_80__124_, chained_data_delayed_80__123_, chained_data_delayed_80__122_, chained_data_delayed_80__121_, chained_data_delayed_80__120_, chained_data_delayed_80__119_, chained_data_delayed_80__118_, chained_data_delayed_80__117_, chained_data_delayed_80__116_, chained_data_delayed_80__115_, chained_data_delayed_80__114_, chained_data_delayed_80__113_, chained_data_delayed_80__112_, chained_data_delayed_80__111_, chained_data_delayed_80__110_, chained_data_delayed_80__109_, chained_data_delayed_80__108_, chained_data_delayed_80__107_, chained_data_delayed_80__106_, chained_data_delayed_80__105_, chained_data_delayed_80__104_, chained_data_delayed_80__103_, chained_data_delayed_80__102_, chained_data_delayed_80__101_, chained_data_delayed_80__100_, chained_data_delayed_80__99_, chained_data_delayed_80__98_, chained_data_delayed_80__97_, chained_data_delayed_80__96_, chained_data_delayed_80__95_, chained_data_delayed_80__94_, chained_data_delayed_80__93_, chained_data_delayed_80__92_, chained_data_delayed_80__91_, chained_data_delayed_80__90_, chained_data_delayed_80__89_, chained_data_delayed_80__88_, chained_data_delayed_80__87_, chained_data_delayed_80__86_, chained_data_delayed_80__85_, chained_data_delayed_80__84_, chained_data_delayed_80__83_, chained_data_delayed_80__82_, chained_data_delayed_80__81_, chained_data_delayed_80__80_, chained_data_delayed_80__79_, chained_data_delayed_80__78_, chained_data_delayed_80__77_, chained_data_delayed_80__76_, chained_data_delayed_80__75_, chained_data_delayed_80__74_, chained_data_delayed_80__73_, chained_data_delayed_80__72_, chained_data_delayed_80__71_, chained_data_delayed_80__70_, chained_data_delayed_80__69_, chained_data_delayed_80__68_, chained_data_delayed_80__67_, chained_data_delayed_80__66_, chained_data_delayed_80__65_, chained_data_delayed_80__64_, chained_data_delayed_80__63_, chained_data_delayed_80__62_, chained_data_delayed_80__61_, chained_data_delayed_80__60_, chained_data_delayed_80__59_, chained_data_delayed_80__58_, chained_data_delayed_80__57_, chained_data_delayed_80__56_, chained_data_delayed_80__55_, chained_data_delayed_80__54_, chained_data_delayed_80__53_, chained_data_delayed_80__52_, chained_data_delayed_80__51_, chained_data_delayed_80__50_, chained_data_delayed_80__49_, chained_data_delayed_80__48_, chained_data_delayed_80__47_, chained_data_delayed_80__46_, chained_data_delayed_80__45_, chained_data_delayed_80__44_, chained_data_delayed_80__43_, chained_data_delayed_80__42_, chained_data_delayed_80__41_, chained_data_delayed_80__40_, chained_data_delayed_80__39_, chained_data_delayed_80__38_, chained_data_delayed_80__37_, chained_data_delayed_80__36_, chained_data_delayed_80__35_, chained_data_delayed_80__34_, chained_data_delayed_80__33_, chained_data_delayed_80__32_, chained_data_delayed_80__31_, chained_data_delayed_80__30_, chained_data_delayed_80__29_, chained_data_delayed_80__28_, chained_data_delayed_80__27_, chained_data_delayed_80__26_, chained_data_delayed_80__25_, chained_data_delayed_80__24_, chained_data_delayed_80__23_, chained_data_delayed_80__22_, chained_data_delayed_80__21_, chained_data_delayed_80__20_, chained_data_delayed_80__19_, chained_data_delayed_80__18_, chained_data_delayed_80__17_, chained_data_delayed_80__16_, chained_data_delayed_80__15_, chained_data_delayed_80__14_, chained_data_delayed_80__13_, chained_data_delayed_80__12_, chained_data_delayed_80__11_, chained_data_delayed_80__10_, chained_data_delayed_80__9_, chained_data_delayed_80__8_, chained_data_delayed_80__7_, chained_data_delayed_80__6_, chained_data_delayed_80__5_, chained_data_delayed_80__4_, chained_data_delayed_80__3_, chained_data_delayed_80__2_, chained_data_delayed_80__1_, chained_data_delayed_80__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_81__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_80__127_, chained_data_delayed_80__126_, chained_data_delayed_80__125_, chained_data_delayed_80__124_, chained_data_delayed_80__123_, chained_data_delayed_80__122_, chained_data_delayed_80__121_, chained_data_delayed_80__120_, chained_data_delayed_80__119_, chained_data_delayed_80__118_, chained_data_delayed_80__117_, chained_data_delayed_80__116_, chained_data_delayed_80__115_, chained_data_delayed_80__114_, chained_data_delayed_80__113_, chained_data_delayed_80__112_, chained_data_delayed_80__111_, chained_data_delayed_80__110_, chained_data_delayed_80__109_, chained_data_delayed_80__108_, chained_data_delayed_80__107_, chained_data_delayed_80__106_, chained_data_delayed_80__105_, chained_data_delayed_80__104_, chained_data_delayed_80__103_, chained_data_delayed_80__102_, chained_data_delayed_80__101_, chained_data_delayed_80__100_, chained_data_delayed_80__99_, chained_data_delayed_80__98_, chained_data_delayed_80__97_, chained_data_delayed_80__96_, chained_data_delayed_80__95_, chained_data_delayed_80__94_, chained_data_delayed_80__93_, chained_data_delayed_80__92_, chained_data_delayed_80__91_, chained_data_delayed_80__90_, chained_data_delayed_80__89_, chained_data_delayed_80__88_, chained_data_delayed_80__87_, chained_data_delayed_80__86_, chained_data_delayed_80__85_, chained_data_delayed_80__84_, chained_data_delayed_80__83_, chained_data_delayed_80__82_, chained_data_delayed_80__81_, chained_data_delayed_80__80_, chained_data_delayed_80__79_, chained_data_delayed_80__78_, chained_data_delayed_80__77_, chained_data_delayed_80__76_, chained_data_delayed_80__75_, chained_data_delayed_80__74_, chained_data_delayed_80__73_, chained_data_delayed_80__72_, chained_data_delayed_80__71_, chained_data_delayed_80__70_, chained_data_delayed_80__69_, chained_data_delayed_80__68_, chained_data_delayed_80__67_, chained_data_delayed_80__66_, chained_data_delayed_80__65_, chained_data_delayed_80__64_, chained_data_delayed_80__63_, chained_data_delayed_80__62_, chained_data_delayed_80__61_, chained_data_delayed_80__60_, chained_data_delayed_80__59_, chained_data_delayed_80__58_, chained_data_delayed_80__57_, chained_data_delayed_80__56_, chained_data_delayed_80__55_, chained_data_delayed_80__54_, chained_data_delayed_80__53_, chained_data_delayed_80__52_, chained_data_delayed_80__51_, chained_data_delayed_80__50_, chained_data_delayed_80__49_, chained_data_delayed_80__48_, chained_data_delayed_80__47_, chained_data_delayed_80__46_, chained_data_delayed_80__45_, chained_data_delayed_80__44_, chained_data_delayed_80__43_, chained_data_delayed_80__42_, chained_data_delayed_80__41_, chained_data_delayed_80__40_, chained_data_delayed_80__39_, chained_data_delayed_80__38_, chained_data_delayed_80__37_, chained_data_delayed_80__36_, chained_data_delayed_80__35_, chained_data_delayed_80__34_, chained_data_delayed_80__33_, chained_data_delayed_80__32_, chained_data_delayed_80__31_, chained_data_delayed_80__30_, chained_data_delayed_80__29_, chained_data_delayed_80__28_, chained_data_delayed_80__27_, chained_data_delayed_80__26_, chained_data_delayed_80__25_, chained_data_delayed_80__24_, chained_data_delayed_80__23_, chained_data_delayed_80__22_, chained_data_delayed_80__21_, chained_data_delayed_80__20_, chained_data_delayed_80__19_, chained_data_delayed_80__18_, chained_data_delayed_80__17_, chained_data_delayed_80__16_, chained_data_delayed_80__15_, chained_data_delayed_80__14_, chained_data_delayed_80__13_, chained_data_delayed_80__12_, chained_data_delayed_80__11_, chained_data_delayed_80__10_, chained_data_delayed_80__9_, chained_data_delayed_80__8_, chained_data_delayed_80__7_, chained_data_delayed_80__6_, chained_data_delayed_80__5_, chained_data_delayed_80__4_, chained_data_delayed_80__3_, chained_data_delayed_80__2_, chained_data_delayed_80__1_, chained_data_delayed_80__0_ }),
    .data_o({ chained_data_delayed_81__127_, chained_data_delayed_81__126_, chained_data_delayed_81__125_, chained_data_delayed_81__124_, chained_data_delayed_81__123_, chained_data_delayed_81__122_, chained_data_delayed_81__121_, chained_data_delayed_81__120_, chained_data_delayed_81__119_, chained_data_delayed_81__118_, chained_data_delayed_81__117_, chained_data_delayed_81__116_, chained_data_delayed_81__115_, chained_data_delayed_81__114_, chained_data_delayed_81__113_, chained_data_delayed_81__112_, chained_data_delayed_81__111_, chained_data_delayed_81__110_, chained_data_delayed_81__109_, chained_data_delayed_81__108_, chained_data_delayed_81__107_, chained_data_delayed_81__106_, chained_data_delayed_81__105_, chained_data_delayed_81__104_, chained_data_delayed_81__103_, chained_data_delayed_81__102_, chained_data_delayed_81__101_, chained_data_delayed_81__100_, chained_data_delayed_81__99_, chained_data_delayed_81__98_, chained_data_delayed_81__97_, chained_data_delayed_81__96_, chained_data_delayed_81__95_, chained_data_delayed_81__94_, chained_data_delayed_81__93_, chained_data_delayed_81__92_, chained_data_delayed_81__91_, chained_data_delayed_81__90_, chained_data_delayed_81__89_, chained_data_delayed_81__88_, chained_data_delayed_81__87_, chained_data_delayed_81__86_, chained_data_delayed_81__85_, chained_data_delayed_81__84_, chained_data_delayed_81__83_, chained_data_delayed_81__82_, chained_data_delayed_81__81_, chained_data_delayed_81__80_, chained_data_delayed_81__79_, chained_data_delayed_81__78_, chained_data_delayed_81__77_, chained_data_delayed_81__76_, chained_data_delayed_81__75_, chained_data_delayed_81__74_, chained_data_delayed_81__73_, chained_data_delayed_81__72_, chained_data_delayed_81__71_, chained_data_delayed_81__70_, chained_data_delayed_81__69_, chained_data_delayed_81__68_, chained_data_delayed_81__67_, chained_data_delayed_81__66_, chained_data_delayed_81__65_, chained_data_delayed_81__64_, chained_data_delayed_81__63_, chained_data_delayed_81__62_, chained_data_delayed_81__61_, chained_data_delayed_81__60_, chained_data_delayed_81__59_, chained_data_delayed_81__58_, chained_data_delayed_81__57_, chained_data_delayed_81__56_, chained_data_delayed_81__55_, chained_data_delayed_81__54_, chained_data_delayed_81__53_, chained_data_delayed_81__52_, chained_data_delayed_81__51_, chained_data_delayed_81__50_, chained_data_delayed_81__49_, chained_data_delayed_81__48_, chained_data_delayed_81__47_, chained_data_delayed_81__46_, chained_data_delayed_81__45_, chained_data_delayed_81__44_, chained_data_delayed_81__43_, chained_data_delayed_81__42_, chained_data_delayed_81__41_, chained_data_delayed_81__40_, chained_data_delayed_81__39_, chained_data_delayed_81__38_, chained_data_delayed_81__37_, chained_data_delayed_81__36_, chained_data_delayed_81__35_, chained_data_delayed_81__34_, chained_data_delayed_81__33_, chained_data_delayed_81__32_, chained_data_delayed_81__31_, chained_data_delayed_81__30_, chained_data_delayed_81__29_, chained_data_delayed_81__28_, chained_data_delayed_81__27_, chained_data_delayed_81__26_, chained_data_delayed_81__25_, chained_data_delayed_81__24_, chained_data_delayed_81__23_, chained_data_delayed_81__22_, chained_data_delayed_81__21_, chained_data_delayed_81__20_, chained_data_delayed_81__19_, chained_data_delayed_81__18_, chained_data_delayed_81__17_, chained_data_delayed_81__16_, chained_data_delayed_81__15_, chained_data_delayed_81__14_, chained_data_delayed_81__13_, chained_data_delayed_81__12_, chained_data_delayed_81__11_, chained_data_delayed_81__10_, chained_data_delayed_81__9_, chained_data_delayed_81__8_, chained_data_delayed_81__7_, chained_data_delayed_81__6_, chained_data_delayed_81__5_, chained_data_delayed_81__4_, chained_data_delayed_81__3_, chained_data_delayed_81__2_, chained_data_delayed_81__1_, chained_data_delayed_81__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_82__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_81__127_, chained_data_delayed_81__126_, chained_data_delayed_81__125_, chained_data_delayed_81__124_, chained_data_delayed_81__123_, chained_data_delayed_81__122_, chained_data_delayed_81__121_, chained_data_delayed_81__120_, chained_data_delayed_81__119_, chained_data_delayed_81__118_, chained_data_delayed_81__117_, chained_data_delayed_81__116_, chained_data_delayed_81__115_, chained_data_delayed_81__114_, chained_data_delayed_81__113_, chained_data_delayed_81__112_, chained_data_delayed_81__111_, chained_data_delayed_81__110_, chained_data_delayed_81__109_, chained_data_delayed_81__108_, chained_data_delayed_81__107_, chained_data_delayed_81__106_, chained_data_delayed_81__105_, chained_data_delayed_81__104_, chained_data_delayed_81__103_, chained_data_delayed_81__102_, chained_data_delayed_81__101_, chained_data_delayed_81__100_, chained_data_delayed_81__99_, chained_data_delayed_81__98_, chained_data_delayed_81__97_, chained_data_delayed_81__96_, chained_data_delayed_81__95_, chained_data_delayed_81__94_, chained_data_delayed_81__93_, chained_data_delayed_81__92_, chained_data_delayed_81__91_, chained_data_delayed_81__90_, chained_data_delayed_81__89_, chained_data_delayed_81__88_, chained_data_delayed_81__87_, chained_data_delayed_81__86_, chained_data_delayed_81__85_, chained_data_delayed_81__84_, chained_data_delayed_81__83_, chained_data_delayed_81__82_, chained_data_delayed_81__81_, chained_data_delayed_81__80_, chained_data_delayed_81__79_, chained_data_delayed_81__78_, chained_data_delayed_81__77_, chained_data_delayed_81__76_, chained_data_delayed_81__75_, chained_data_delayed_81__74_, chained_data_delayed_81__73_, chained_data_delayed_81__72_, chained_data_delayed_81__71_, chained_data_delayed_81__70_, chained_data_delayed_81__69_, chained_data_delayed_81__68_, chained_data_delayed_81__67_, chained_data_delayed_81__66_, chained_data_delayed_81__65_, chained_data_delayed_81__64_, chained_data_delayed_81__63_, chained_data_delayed_81__62_, chained_data_delayed_81__61_, chained_data_delayed_81__60_, chained_data_delayed_81__59_, chained_data_delayed_81__58_, chained_data_delayed_81__57_, chained_data_delayed_81__56_, chained_data_delayed_81__55_, chained_data_delayed_81__54_, chained_data_delayed_81__53_, chained_data_delayed_81__52_, chained_data_delayed_81__51_, chained_data_delayed_81__50_, chained_data_delayed_81__49_, chained_data_delayed_81__48_, chained_data_delayed_81__47_, chained_data_delayed_81__46_, chained_data_delayed_81__45_, chained_data_delayed_81__44_, chained_data_delayed_81__43_, chained_data_delayed_81__42_, chained_data_delayed_81__41_, chained_data_delayed_81__40_, chained_data_delayed_81__39_, chained_data_delayed_81__38_, chained_data_delayed_81__37_, chained_data_delayed_81__36_, chained_data_delayed_81__35_, chained_data_delayed_81__34_, chained_data_delayed_81__33_, chained_data_delayed_81__32_, chained_data_delayed_81__31_, chained_data_delayed_81__30_, chained_data_delayed_81__29_, chained_data_delayed_81__28_, chained_data_delayed_81__27_, chained_data_delayed_81__26_, chained_data_delayed_81__25_, chained_data_delayed_81__24_, chained_data_delayed_81__23_, chained_data_delayed_81__22_, chained_data_delayed_81__21_, chained_data_delayed_81__20_, chained_data_delayed_81__19_, chained_data_delayed_81__18_, chained_data_delayed_81__17_, chained_data_delayed_81__16_, chained_data_delayed_81__15_, chained_data_delayed_81__14_, chained_data_delayed_81__13_, chained_data_delayed_81__12_, chained_data_delayed_81__11_, chained_data_delayed_81__10_, chained_data_delayed_81__9_, chained_data_delayed_81__8_, chained_data_delayed_81__7_, chained_data_delayed_81__6_, chained_data_delayed_81__5_, chained_data_delayed_81__4_, chained_data_delayed_81__3_, chained_data_delayed_81__2_, chained_data_delayed_81__1_, chained_data_delayed_81__0_ }),
    .data_o({ chained_data_delayed_82__127_, chained_data_delayed_82__126_, chained_data_delayed_82__125_, chained_data_delayed_82__124_, chained_data_delayed_82__123_, chained_data_delayed_82__122_, chained_data_delayed_82__121_, chained_data_delayed_82__120_, chained_data_delayed_82__119_, chained_data_delayed_82__118_, chained_data_delayed_82__117_, chained_data_delayed_82__116_, chained_data_delayed_82__115_, chained_data_delayed_82__114_, chained_data_delayed_82__113_, chained_data_delayed_82__112_, chained_data_delayed_82__111_, chained_data_delayed_82__110_, chained_data_delayed_82__109_, chained_data_delayed_82__108_, chained_data_delayed_82__107_, chained_data_delayed_82__106_, chained_data_delayed_82__105_, chained_data_delayed_82__104_, chained_data_delayed_82__103_, chained_data_delayed_82__102_, chained_data_delayed_82__101_, chained_data_delayed_82__100_, chained_data_delayed_82__99_, chained_data_delayed_82__98_, chained_data_delayed_82__97_, chained_data_delayed_82__96_, chained_data_delayed_82__95_, chained_data_delayed_82__94_, chained_data_delayed_82__93_, chained_data_delayed_82__92_, chained_data_delayed_82__91_, chained_data_delayed_82__90_, chained_data_delayed_82__89_, chained_data_delayed_82__88_, chained_data_delayed_82__87_, chained_data_delayed_82__86_, chained_data_delayed_82__85_, chained_data_delayed_82__84_, chained_data_delayed_82__83_, chained_data_delayed_82__82_, chained_data_delayed_82__81_, chained_data_delayed_82__80_, chained_data_delayed_82__79_, chained_data_delayed_82__78_, chained_data_delayed_82__77_, chained_data_delayed_82__76_, chained_data_delayed_82__75_, chained_data_delayed_82__74_, chained_data_delayed_82__73_, chained_data_delayed_82__72_, chained_data_delayed_82__71_, chained_data_delayed_82__70_, chained_data_delayed_82__69_, chained_data_delayed_82__68_, chained_data_delayed_82__67_, chained_data_delayed_82__66_, chained_data_delayed_82__65_, chained_data_delayed_82__64_, chained_data_delayed_82__63_, chained_data_delayed_82__62_, chained_data_delayed_82__61_, chained_data_delayed_82__60_, chained_data_delayed_82__59_, chained_data_delayed_82__58_, chained_data_delayed_82__57_, chained_data_delayed_82__56_, chained_data_delayed_82__55_, chained_data_delayed_82__54_, chained_data_delayed_82__53_, chained_data_delayed_82__52_, chained_data_delayed_82__51_, chained_data_delayed_82__50_, chained_data_delayed_82__49_, chained_data_delayed_82__48_, chained_data_delayed_82__47_, chained_data_delayed_82__46_, chained_data_delayed_82__45_, chained_data_delayed_82__44_, chained_data_delayed_82__43_, chained_data_delayed_82__42_, chained_data_delayed_82__41_, chained_data_delayed_82__40_, chained_data_delayed_82__39_, chained_data_delayed_82__38_, chained_data_delayed_82__37_, chained_data_delayed_82__36_, chained_data_delayed_82__35_, chained_data_delayed_82__34_, chained_data_delayed_82__33_, chained_data_delayed_82__32_, chained_data_delayed_82__31_, chained_data_delayed_82__30_, chained_data_delayed_82__29_, chained_data_delayed_82__28_, chained_data_delayed_82__27_, chained_data_delayed_82__26_, chained_data_delayed_82__25_, chained_data_delayed_82__24_, chained_data_delayed_82__23_, chained_data_delayed_82__22_, chained_data_delayed_82__21_, chained_data_delayed_82__20_, chained_data_delayed_82__19_, chained_data_delayed_82__18_, chained_data_delayed_82__17_, chained_data_delayed_82__16_, chained_data_delayed_82__15_, chained_data_delayed_82__14_, chained_data_delayed_82__13_, chained_data_delayed_82__12_, chained_data_delayed_82__11_, chained_data_delayed_82__10_, chained_data_delayed_82__9_, chained_data_delayed_82__8_, chained_data_delayed_82__7_, chained_data_delayed_82__6_, chained_data_delayed_82__5_, chained_data_delayed_82__4_, chained_data_delayed_82__3_, chained_data_delayed_82__2_, chained_data_delayed_82__1_, chained_data_delayed_82__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_83__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_82__127_, chained_data_delayed_82__126_, chained_data_delayed_82__125_, chained_data_delayed_82__124_, chained_data_delayed_82__123_, chained_data_delayed_82__122_, chained_data_delayed_82__121_, chained_data_delayed_82__120_, chained_data_delayed_82__119_, chained_data_delayed_82__118_, chained_data_delayed_82__117_, chained_data_delayed_82__116_, chained_data_delayed_82__115_, chained_data_delayed_82__114_, chained_data_delayed_82__113_, chained_data_delayed_82__112_, chained_data_delayed_82__111_, chained_data_delayed_82__110_, chained_data_delayed_82__109_, chained_data_delayed_82__108_, chained_data_delayed_82__107_, chained_data_delayed_82__106_, chained_data_delayed_82__105_, chained_data_delayed_82__104_, chained_data_delayed_82__103_, chained_data_delayed_82__102_, chained_data_delayed_82__101_, chained_data_delayed_82__100_, chained_data_delayed_82__99_, chained_data_delayed_82__98_, chained_data_delayed_82__97_, chained_data_delayed_82__96_, chained_data_delayed_82__95_, chained_data_delayed_82__94_, chained_data_delayed_82__93_, chained_data_delayed_82__92_, chained_data_delayed_82__91_, chained_data_delayed_82__90_, chained_data_delayed_82__89_, chained_data_delayed_82__88_, chained_data_delayed_82__87_, chained_data_delayed_82__86_, chained_data_delayed_82__85_, chained_data_delayed_82__84_, chained_data_delayed_82__83_, chained_data_delayed_82__82_, chained_data_delayed_82__81_, chained_data_delayed_82__80_, chained_data_delayed_82__79_, chained_data_delayed_82__78_, chained_data_delayed_82__77_, chained_data_delayed_82__76_, chained_data_delayed_82__75_, chained_data_delayed_82__74_, chained_data_delayed_82__73_, chained_data_delayed_82__72_, chained_data_delayed_82__71_, chained_data_delayed_82__70_, chained_data_delayed_82__69_, chained_data_delayed_82__68_, chained_data_delayed_82__67_, chained_data_delayed_82__66_, chained_data_delayed_82__65_, chained_data_delayed_82__64_, chained_data_delayed_82__63_, chained_data_delayed_82__62_, chained_data_delayed_82__61_, chained_data_delayed_82__60_, chained_data_delayed_82__59_, chained_data_delayed_82__58_, chained_data_delayed_82__57_, chained_data_delayed_82__56_, chained_data_delayed_82__55_, chained_data_delayed_82__54_, chained_data_delayed_82__53_, chained_data_delayed_82__52_, chained_data_delayed_82__51_, chained_data_delayed_82__50_, chained_data_delayed_82__49_, chained_data_delayed_82__48_, chained_data_delayed_82__47_, chained_data_delayed_82__46_, chained_data_delayed_82__45_, chained_data_delayed_82__44_, chained_data_delayed_82__43_, chained_data_delayed_82__42_, chained_data_delayed_82__41_, chained_data_delayed_82__40_, chained_data_delayed_82__39_, chained_data_delayed_82__38_, chained_data_delayed_82__37_, chained_data_delayed_82__36_, chained_data_delayed_82__35_, chained_data_delayed_82__34_, chained_data_delayed_82__33_, chained_data_delayed_82__32_, chained_data_delayed_82__31_, chained_data_delayed_82__30_, chained_data_delayed_82__29_, chained_data_delayed_82__28_, chained_data_delayed_82__27_, chained_data_delayed_82__26_, chained_data_delayed_82__25_, chained_data_delayed_82__24_, chained_data_delayed_82__23_, chained_data_delayed_82__22_, chained_data_delayed_82__21_, chained_data_delayed_82__20_, chained_data_delayed_82__19_, chained_data_delayed_82__18_, chained_data_delayed_82__17_, chained_data_delayed_82__16_, chained_data_delayed_82__15_, chained_data_delayed_82__14_, chained_data_delayed_82__13_, chained_data_delayed_82__12_, chained_data_delayed_82__11_, chained_data_delayed_82__10_, chained_data_delayed_82__9_, chained_data_delayed_82__8_, chained_data_delayed_82__7_, chained_data_delayed_82__6_, chained_data_delayed_82__5_, chained_data_delayed_82__4_, chained_data_delayed_82__3_, chained_data_delayed_82__2_, chained_data_delayed_82__1_, chained_data_delayed_82__0_ }),
    .data_o({ chained_data_delayed_83__127_, chained_data_delayed_83__126_, chained_data_delayed_83__125_, chained_data_delayed_83__124_, chained_data_delayed_83__123_, chained_data_delayed_83__122_, chained_data_delayed_83__121_, chained_data_delayed_83__120_, chained_data_delayed_83__119_, chained_data_delayed_83__118_, chained_data_delayed_83__117_, chained_data_delayed_83__116_, chained_data_delayed_83__115_, chained_data_delayed_83__114_, chained_data_delayed_83__113_, chained_data_delayed_83__112_, chained_data_delayed_83__111_, chained_data_delayed_83__110_, chained_data_delayed_83__109_, chained_data_delayed_83__108_, chained_data_delayed_83__107_, chained_data_delayed_83__106_, chained_data_delayed_83__105_, chained_data_delayed_83__104_, chained_data_delayed_83__103_, chained_data_delayed_83__102_, chained_data_delayed_83__101_, chained_data_delayed_83__100_, chained_data_delayed_83__99_, chained_data_delayed_83__98_, chained_data_delayed_83__97_, chained_data_delayed_83__96_, chained_data_delayed_83__95_, chained_data_delayed_83__94_, chained_data_delayed_83__93_, chained_data_delayed_83__92_, chained_data_delayed_83__91_, chained_data_delayed_83__90_, chained_data_delayed_83__89_, chained_data_delayed_83__88_, chained_data_delayed_83__87_, chained_data_delayed_83__86_, chained_data_delayed_83__85_, chained_data_delayed_83__84_, chained_data_delayed_83__83_, chained_data_delayed_83__82_, chained_data_delayed_83__81_, chained_data_delayed_83__80_, chained_data_delayed_83__79_, chained_data_delayed_83__78_, chained_data_delayed_83__77_, chained_data_delayed_83__76_, chained_data_delayed_83__75_, chained_data_delayed_83__74_, chained_data_delayed_83__73_, chained_data_delayed_83__72_, chained_data_delayed_83__71_, chained_data_delayed_83__70_, chained_data_delayed_83__69_, chained_data_delayed_83__68_, chained_data_delayed_83__67_, chained_data_delayed_83__66_, chained_data_delayed_83__65_, chained_data_delayed_83__64_, chained_data_delayed_83__63_, chained_data_delayed_83__62_, chained_data_delayed_83__61_, chained_data_delayed_83__60_, chained_data_delayed_83__59_, chained_data_delayed_83__58_, chained_data_delayed_83__57_, chained_data_delayed_83__56_, chained_data_delayed_83__55_, chained_data_delayed_83__54_, chained_data_delayed_83__53_, chained_data_delayed_83__52_, chained_data_delayed_83__51_, chained_data_delayed_83__50_, chained_data_delayed_83__49_, chained_data_delayed_83__48_, chained_data_delayed_83__47_, chained_data_delayed_83__46_, chained_data_delayed_83__45_, chained_data_delayed_83__44_, chained_data_delayed_83__43_, chained_data_delayed_83__42_, chained_data_delayed_83__41_, chained_data_delayed_83__40_, chained_data_delayed_83__39_, chained_data_delayed_83__38_, chained_data_delayed_83__37_, chained_data_delayed_83__36_, chained_data_delayed_83__35_, chained_data_delayed_83__34_, chained_data_delayed_83__33_, chained_data_delayed_83__32_, chained_data_delayed_83__31_, chained_data_delayed_83__30_, chained_data_delayed_83__29_, chained_data_delayed_83__28_, chained_data_delayed_83__27_, chained_data_delayed_83__26_, chained_data_delayed_83__25_, chained_data_delayed_83__24_, chained_data_delayed_83__23_, chained_data_delayed_83__22_, chained_data_delayed_83__21_, chained_data_delayed_83__20_, chained_data_delayed_83__19_, chained_data_delayed_83__18_, chained_data_delayed_83__17_, chained_data_delayed_83__16_, chained_data_delayed_83__15_, chained_data_delayed_83__14_, chained_data_delayed_83__13_, chained_data_delayed_83__12_, chained_data_delayed_83__11_, chained_data_delayed_83__10_, chained_data_delayed_83__9_, chained_data_delayed_83__8_, chained_data_delayed_83__7_, chained_data_delayed_83__6_, chained_data_delayed_83__5_, chained_data_delayed_83__4_, chained_data_delayed_83__3_, chained_data_delayed_83__2_, chained_data_delayed_83__1_, chained_data_delayed_83__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_84__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_83__127_, chained_data_delayed_83__126_, chained_data_delayed_83__125_, chained_data_delayed_83__124_, chained_data_delayed_83__123_, chained_data_delayed_83__122_, chained_data_delayed_83__121_, chained_data_delayed_83__120_, chained_data_delayed_83__119_, chained_data_delayed_83__118_, chained_data_delayed_83__117_, chained_data_delayed_83__116_, chained_data_delayed_83__115_, chained_data_delayed_83__114_, chained_data_delayed_83__113_, chained_data_delayed_83__112_, chained_data_delayed_83__111_, chained_data_delayed_83__110_, chained_data_delayed_83__109_, chained_data_delayed_83__108_, chained_data_delayed_83__107_, chained_data_delayed_83__106_, chained_data_delayed_83__105_, chained_data_delayed_83__104_, chained_data_delayed_83__103_, chained_data_delayed_83__102_, chained_data_delayed_83__101_, chained_data_delayed_83__100_, chained_data_delayed_83__99_, chained_data_delayed_83__98_, chained_data_delayed_83__97_, chained_data_delayed_83__96_, chained_data_delayed_83__95_, chained_data_delayed_83__94_, chained_data_delayed_83__93_, chained_data_delayed_83__92_, chained_data_delayed_83__91_, chained_data_delayed_83__90_, chained_data_delayed_83__89_, chained_data_delayed_83__88_, chained_data_delayed_83__87_, chained_data_delayed_83__86_, chained_data_delayed_83__85_, chained_data_delayed_83__84_, chained_data_delayed_83__83_, chained_data_delayed_83__82_, chained_data_delayed_83__81_, chained_data_delayed_83__80_, chained_data_delayed_83__79_, chained_data_delayed_83__78_, chained_data_delayed_83__77_, chained_data_delayed_83__76_, chained_data_delayed_83__75_, chained_data_delayed_83__74_, chained_data_delayed_83__73_, chained_data_delayed_83__72_, chained_data_delayed_83__71_, chained_data_delayed_83__70_, chained_data_delayed_83__69_, chained_data_delayed_83__68_, chained_data_delayed_83__67_, chained_data_delayed_83__66_, chained_data_delayed_83__65_, chained_data_delayed_83__64_, chained_data_delayed_83__63_, chained_data_delayed_83__62_, chained_data_delayed_83__61_, chained_data_delayed_83__60_, chained_data_delayed_83__59_, chained_data_delayed_83__58_, chained_data_delayed_83__57_, chained_data_delayed_83__56_, chained_data_delayed_83__55_, chained_data_delayed_83__54_, chained_data_delayed_83__53_, chained_data_delayed_83__52_, chained_data_delayed_83__51_, chained_data_delayed_83__50_, chained_data_delayed_83__49_, chained_data_delayed_83__48_, chained_data_delayed_83__47_, chained_data_delayed_83__46_, chained_data_delayed_83__45_, chained_data_delayed_83__44_, chained_data_delayed_83__43_, chained_data_delayed_83__42_, chained_data_delayed_83__41_, chained_data_delayed_83__40_, chained_data_delayed_83__39_, chained_data_delayed_83__38_, chained_data_delayed_83__37_, chained_data_delayed_83__36_, chained_data_delayed_83__35_, chained_data_delayed_83__34_, chained_data_delayed_83__33_, chained_data_delayed_83__32_, chained_data_delayed_83__31_, chained_data_delayed_83__30_, chained_data_delayed_83__29_, chained_data_delayed_83__28_, chained_data_delayed_83__27_, chained_data_delayed_83__26_, chained_data_delayed_83__25_, chained_data_delayed_83__24_, chained_data_delayed_83__23_, chained_data_delayed_83__22_, chained_data_delayed_83__21_, chained_data_delayed_83__20_, chained_data_delayed_83__19_, chained_data_delayed_83__18_, chained_data_delayed_83__17_, chained_data_delayed_83__16_, chained_data_delayed_83__15_, chained_data_delayed_83__14_, chained_data_delayed_83__13_, chained_data_delayed_83__12_, chained_data_delayed_83__11_, chained_data_delayed_83__10_, chained_data_delayed_83__9_, chained_data_delayed_83__8_, chained_data_delayed_83__7_, chained_data_delayed_83__6_, chained_data_delayed_83__5_, chained_data_delayed_83__4_, chained_data_delayed_83__3_, chained_data_delayed_83__2_, chained_data_delayed_83__1_, chained_data_delayed_83__0_ }),
    .data_o({ chained_data_delayed_84__127_, chained_data_delayed_84__126_, chained_data_delayed_84__125_, chained_data_delayed_84__124_, chained_data_delayed_84__123_, chained_data_delayed_84__122_, chained_data_delayed_84__121_, chained_data_delayed_84__120_, chained_data_delayed_84__119_, chained_data_delayed_84__118_, chained_data_delayed_84__117_, chained_data_delayed_84__116_, chained_data_delayed_84__115_, chained_data_delayed_84__114_, chained_data_delayed_84__113_, chained_data_delayed_84__112_, chained_data_delayed_84__111_, chained_data_delayed_84__110_, chained_data_delayed_84__109_, chained_data_delayed_84__108_, chained_data_delayed_84__107_, chained_data_delayed_84__106_, chained_data_delayed_84__105_, chained_data_delayed_84__104_, chained_data_delayed_84__103_, chained_data_delayed_84__102_, chained_data_delayed_84__101_, chained_data_delayed_84__100_, chained_data_delayed_84__99_, chained_data_delayed_84__98_, chained_data_delayed_84__97_, chained_data_delayed_84__96_, chained_data_delayed_84__95_, chained_data_delayed_84__94_, chained_data_delayed_84__93_, chained_data_delayed_84__92_, chained_data_delayed_84__91_, chained_data_delayed_84__90_, chained_data_delayed_84__89_, chained_data_delayed_84__88_, chained_data_delayed_84__87_, chained_data_delayed_84__86_, chained_data_delayed_84__85_, chained_data_delayed_84__84_, chained_data_delayed_84__83_, chained_data_delayed_84__82_, chained_data_delayed_84__81_, chained_data_delayed_84__80_, chained_data_delayed_84__79_, chained_data_delayed_84__78_, chained_data_delayed_84__77_, chained_data_delayed_84__76_, chained_data_delayed_84__75_, chained_data_delayed_84__74_, chained_data_delayed_84__73_, chained_data_delayed_84__72_, chained_data_delayed_84__71_, chained_data_delayed_84__70_, chained_data_delayed_84__69_, chained_data_delayed_84__68_, chained_data_delayed_84__67_, chained_data_delayed_84__66_, chained_data_delayed_84__65_, chained_data_delayed_84__64_, chained_data_delayed_84__63_, chained_data_delayed_84__62_, chained_data_delayed_84__61_, chained_data_delayed_84__60_, chained_data_delayed_84__59_, chained_data_delayed_84__58_, chained_data_delayed_84__57_, chained_data_delayed_84__56_, chained_data_delayed_84__55_, chained_data_delayed_84__54_, chained_data_delayed_84__53_, chained_data_delayed_84__52_, chained_data_delayed_84__51_, chained_data_delayed_84__50_, chained_data_delayed_84__49_, chained_data_delayed_84__48_, chained_data_delayed_84__47_, chained_data_delayed_84__46_, chained_data_delayed_84__45_, chained_data_delayed_84__44_, chained_data_delayed_84__43_, chained_data_delayed_84__42_, chained_data_delayed_84__41_, chained_data_delayed_84__40_, chained_data_delayed_84__39_, chained_data_delayed_84__38_, chained_data_delayed_84__37_, chained_data_delayed_84__36_, chained_data_delayed_84__35_, chained_data_delayed_84__34_, chained_data_delayed_84__33_, chained_data_delayed_84__32_, chained_data_delayed_84__31_, chained_data_delayed_84__30_, chained_data_delayed_84__29_, chained_data_delayed_84__28_, chained_data_delayed_84__27_, chained_data_delayed_84__26_, chained_data_delayed_84__25_, chained_data_delayed_84__24_, chained_data_delayed_84__23_, chained_data_delayed_84__22_, chained_data_delayed_84__21_, chained_data_delayed_84__20_, chained_data_delayed_84__19_, chained_data_delayed_84__18_, chained_data_delayed_84__17_, chained_data_delayed_84__16_, chained_data_delayed_84__15_, chained_data_delayed_84__14_, chained_data_delayed_84__13_, chained_data_delayed_84__12_, chained_data_delayed_84__11_, chained_data_delayed_84__10_, chained_data_delayed_84__9_, chained_data_delayed_84__8_, chained_data_delayed_84__7_, chained_data_delayed_84__6_, chained_data_delayed_84__5_, chained_data_delayed_84__4_, chained_data_delayed_84__3_, chained_data_delayed_84__2_, chained_data_delayed_84__1_, chained_data_delayed_84__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_85__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_84__127_, chained_data_delayed_84__126_, chained_data_delayed_84__125_, chained_data_delayed_84__124_, chained_data_delayed_84__123_, chained_data_delayed_84__122_, chained_data_delayed_84__121_, chained_data_delayed_84__120_, chained_data_delayed_84__119_, chained_data_delayed_84__118_, chained_data_delayed_84__117_, chained_data_delayed_84__116_, chained_data_delayed_84__115_, chained_data_delayed_84__114_, chained_data_delayed_84__113_, chained_data_delayed_84__112_, chained_data_delayed_84__111_, chained_data_delayed_84__110_, chained_data_delayed_84__109_, chained_data_delayed_84__108_, chained_data_delayed_84__107_, chained_data_delayed_84__106_, chained_data_delayed_84__105_, chained_data_delayed_84__104_, chained_data_delayed_84__103_, chained_data_delayed_84__102_, chained_data_delayed_84__101_, chained_data_delayed_84__100_, chained_data_delayed_84__99_, chained_data_delayed_84__98_, chained_data_delayed_84__97_, chained_data_delayed_84__96_, chained_data_delayed_84__95_, chained_data_delayed_84__94_, chained_data_delayed_84__93_, chained_data_delayed_84__92_, chained_data_delayed_84__91_, chained_data_delayed_84__90_, chained_data_delayed_84__89_, chained_data_delayed_84__88_, chained_data_delayed_84__87_, chained_data_delayed_84__86_, chained_data_delayed_84__85_, chained_data_delayed_84__84_, chained_data_delayed_84__83_, chained_data_delayed_84__82_, chained_data_delayed_84__81_, chained_data_delayed_84__80_, chained_data_delayed_84__79_, chained_data_delayed_84__78_, chained_data_delayed_84__77_, chained_data_delayed_84__76_, chained_data_delayed_84__75_, chained_data_delayed_84__74_, chained_data_delayed_84__73_, chained_data_delayed_84__72_, chained_data_delayed_84__71_, chained_data_delayed_84__70_, chained_data_delayed_84__69_, chained_data_delayed_84__68_, chained_data_delayed_84__67_, chained_data_delayed_84__66_, chained_data_delayed_84__65_, chained_data_delayed_84__64_, chained_data_delayed_84__63_, chained_data_delayed_84__62_, chained_data_delayed_84__61_, chained_data_delayed_84__60_, chained_data_delayed_84__59_, chained_data_delayed_84__58_, chained_data_delayed_84__57_, chained_data_delayed_84__56_, chained_data_delayed_84__55_, chained_data_delayed_84__54_, chained_data_delayed_84__53_, chained_data_delayed_84__52_, chained_data_delayed_84__51_, chained_data_delayed_84__50_, chained_data_delayed_84__49_, chained_data_delayed_84__48_, chained_data_delayed_84__47_, chained_data_delayed_84__46_, chained_data_delayed_84__45_, chained_data_delayed_84__44_, chained_data_delayed_84__43_, chained_data_delayed_84__42_, chained_data_delayed_84__41_, chained_data_delayed_84__40_, chained_data_delayed_84__39_, chained_data_delayed_84__38_, chained_data_delayed_84__37_, chained_data_delayed_84__36_, chained_data_delayed_84__35_, chained_data_delayed_84__34_, chained_data_delayed_84__33_, chained_data_delayed_84__32_, chained_data_delayed_84__31_, chained_data_delayed_84__30_, chained_data_delayed_84__29_, chained_data_delayed_84__28_, chained_data_delayed_84__27_, chained_data_delayed_84__26_, chained_data_delayed_84__25_, chained_data_delayed_84__24_, chained_data_delayed_84__23_, chained_data_delayed_84__22_, chained_data_delayed_84__21_, chained_data_delayed_84__20_, chained_data_delayed_84__19_, chained_data_delayed_84__18_, chained_data_delayed_84__17_, chained_data_delayed_84__16_, chained_data_delayed_84__15_, chained_data_delayed_84__14_, chained_data_delayed_84__13_, chained_data_delayed_84__12_, chained_data_delayed_84__11_, chained_data_delayed_84__10_, chained_data_delayed_84__9_, chained_data_delayed_84__8_, chained_data_delayed_84__7_, chained_data_delayed_84__6_, chained_data_delayed_84__5_, chained_data_delayed_84__4_, chained_data_delayed_84__3_, chained_data_delayed_84__2_, chained_data_delayed_84__1_, chained_data_delayed_84__0_ }),
    .data_o({ chained_data_delayed_85__127_, chained_data_delayed_85__126_, chained_data_delayed_85__125_, chained_data_delayed_85__124_, chained_data_delayed_85__123_, chained_data_delayed_85__122_, chained_data_delayed_85__121_, chained_data_delayed_85__120_, chained_data_delayed_85__119_, chained_data_delayed_85__118_, chained_data_delayed_85__117_, chained_data_delayed_85__116_, chained_data_delayed_85__115_, chained_data_delayed_85__114_, chained_data_delayed_85__113_, chained_data_delayed_85__112_, chained_data_delayed_85__111_, chained_data_delayed_85__110_, chained_data_delayed_85__109_, chained_data_delayed_85__108_, chained_data_delayed_85__107_, chained_data_delayed_85__106_, chained_data_delayed_85__105_, chained_data_delayed_85__104_, chained_data_delayed_85__103_, chained_data_delayed_85__102_, chained_data_delayed_85__101_, chained_data_delayed_85__100_, chained_data_delayed_85__99_, chained_data_delayed_85__98_, chained_data_delayed_85__97_, chained_data_delayed_85__96_, chained_data_delayed_85__95_, chained_data_delayed_85__94_, chained_data_delayed_85__93_, chained_data_delayed_85__92_, chained_data_delayed_85__91_, chained_data_delayed_85__90_, chained_data_delayed_85__89_, chained_data_delayed_85__88_, chained_data_delayed_85__87_, chained_data_delayed_85__86_, chained_data_delayed_85__85_, chained_data_delayed_85__84_, chained_data_delayed_85__83_, chained_data_delayed_85__82_, chained_data_delayed_85__81_, chained_data_delayed_85__80_, chained_data_delayed_85__79_, chained_data_delayed_85__78_, chained_data_delayed_85__77_, chained_data_delayed_85__76_, chained_data_delayed_85__75_, chained_data_delayed_85__74_, chained_data_delayed_85__73_, chained_data_delayed_85__72_, chained_data_delayed_85__71_, chained_data_delayed_85__70_, chained_data_delayed_85__69_, chained_data_delayed_85__68_, chained_data_delayed_85__67_, chained_data_delayed_85__66_, chained_data_delayed_85__65_, chained_data_delayed_85__64_, chained_data_delayed_85__63_, chained_data_delayed_85__62_, chained_data_delayed_85__61_, chained_data_delayed_85__60_, chained_data_delayed_85__59_, chained_data_delayed_85__58_, chained_data_delayed_85__57_, chained_data_delayed_85__56_, chained_data_delayed_85__55_, chained_data_delayed_85__54_, chained_data_delayed_85__53_, chained_data_delayed_85__52_, chained_data_delayed_85__51_, chained_data_delayed_85__50_, chained_data_delayed_85__49_, chained_data_delayed_85__48_, chained_data_delayed_85__47_, chained_data_delayed_85__46_, chained_data_delayed_85__45_, chained_data_delayed_85__44_, chained_data_delayed_85__43_, chained_data_delayed_85__42_, chained_data_delayed_85__41_, chained_data_delayed_85__40_, chained_data_delayed_85__39_, chained_data_delayed_85__38_, chained_data_delayed_85__37_, chained_data_delayed_85__36_, chained_data_delayed_85__35_, chained_data_delayed_85__34_, chained_data_delayed_85__33_, chained_data_delayed_85__32_, chained_data_delayed_85__31_, chained_data_delayed_85__30_, chained_data_delayed_85__29_, chained_data_delayed_85__28_, chained_data_delayed_85__27_, chained_data_delayed_85__26_, chained_data_delayed_85__25_, chained_data_delayed_85__24_, chained_data_delayed_85__23_, chained_data_delayed_85__22_, chained_data_delayed_85__21_, chained_data_delayed_85__20_, chained_data_delayed_85__19_, chained_data_delayed_85__18_, chained_data_delayed_85__17_, chained_data_delayed_85__16_, chained_data_delayed_85__15_, chained_data_delayed_85__14_, chained_data_delayed_85__13_, chained_data_delayed_85__12_, chained_data_delayed_85__11_, chained_data_delayed_85__10_, chained_data_delayed_85__9_, chained_data_delayed_85__8_, chained_data_delayed_85__7_, chained_data_delayed_85__6_, chained_data_delayed_85__5_, chained_data_delayed_85__4_, chained_data_delayed_85__3_, chained_data_delayed_85__2_, chained_data_delayed_85__1_, chained_data_delayed_85__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_86__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_85__127_, chained_data_delayed_85__126_, chained_data_delayed_85__125_, chained_data_delayed_85__124_, chained_data_delayed_85__123_, chained_data_delayed_85__122_, chained_data_delayed_85__121_, chained_data_delayed_85__120_, chained_data_delayed_85__119_, chained_data_delayed_85__118_, chained_data_delayed_85__117_, chained_data_delayed_85__116_, chained_data_delayed_85__115_, chained_data_delayed_85__114_, chained_data_delayed_85__113_, chained_data_delayed_85__112_, chained_data_delayed_85__111_, chained_data_delayed_85__110_, chained_data_delayed_85__109_, chained_data_delayed_85__108_, chained_data_delayed_85__107_, chained_data_delayed_85__106_, chained_data_delayed_85__105_, chained_data_delayed_85__104_, chained_data_delayed_85__103_, chained_data_delayed_85__102_, chained_data_delayed_85__101_, chained_data_delayed_85__100_, chained_data_delayed_85__99_, chained_data_delayed_85__98_, chained_data_delayed_85__97_, chained_data_delayed_85__96_, chained_data_delayed_85__95_, chained_data_delayed_85__94_, chained_data_delayed_85__93_, chained_data_delayed_85__92_, chained_data_delayed_85__91_, chained_data_delayed_85__90_, chained_data_delayed_85__89_, chained_data_delayed_85__88_, chained_data_delayed_85__87_, chained_data_delayed_85__86_, chained_data_delayed_85__85_, chained_data_delayed_85__84_, chained_data_delayed_85__83_, chained_data_delayed_85__82_, chained_data_delayed_85__81_, chained_data_delayed_85__80_, chained_data_delayed_85__79_, chained_data_delayed_85__78_, chained_data_delayed_85__77_, chained_data_delayed_85__76_, chained_data_delayed_85__75_, chained_data_delayed_85__74_, chained_data_delayed_85__73_, chained_data_delayed_85__72_, chained_data_delayed_85__71_, chained_data_delayed_85__70_, chained_data_delayed_85__69_, chained_data_delayed_85__68_, chained_data_delayed_85__67_, chained_data_delayed_85__66_, chained_data_delayed_85__65_, chained_data_delayed_85__64_, chained_data_delayed_85__63_, chained_data_delayed_85__62_, chained_data_delayed_85__61_, chained_data_delayed_85__60_, chained_data_delayed_85__59_, chained_data_delayed_85__58_, chained_data_delayed_85__57_, chained_data_delayed_85__56_, chained_data_delayed_85__55_, chained_data_delayed_85__54_, chained_data_delayed_85__53_, chained_data_delayed_85__52_, chained_data_delayed_85__51_, chained_data_delayed_85__50_, chained_data_delayed_85__49_, chained_data_delayed_85__48_, chained_data_delayed_85__47_, chained_data_delayed_85__46_, chained_data_delayed_85__45_, chained_data_delayed_85__44_, chained_data_delayed_85__43_, chained_data_delayed_85__42_, chained_data_delayed_85__41_, chained_data_delayed_85__40_, chained_data_delayed_85__39_, chained_data_delayed_85__38_, chained_data_delayed_85__37_, chained_data_delayed_85__36_, chained_data_delayed_85__35_, chained_data_delayed_85__34_, chained_data_delayed_85__33_, chained_data_delayed_85__32_, chained_data_delayed_85__31_, chained_data_delayed_85__30_, chained_data_delayed_85__29_, chained_data_delayed_85__28_, chained_data_delayed_85__27_, chained_data_delayed_85__26_, chained_data_delayed_85__25_, chained_data_delayed_85__24_, chained_data_delayed_85__23_, chained_data_delayed_85__22_, chained_data_delayed_85__21_, chained_data_delayed_85__20_, chained_data_delayed_85__19_, chained_data_delayed_85__18_, chained_data_delayed_85__17_, chained_data_delayed_85__16_, chained_data_delayed_85__15_, chained_data_delayed_85__14_, chained_data_delayed_85__13_, chained_data_delayed_85__12_, chained_data_delayed_85__11_, chained_data_delayed_85__10_, chained_data_delayed_85__9_, chained_data_delayed_85__8_, chained_data_delayed_85__7_, chained_data_delayed_85__6_, chained_data_delayed_85__5_, chained_data_delayed_85__4_, chained_data_delayed_85__3_, chained_data_delayed_85__2_, chained_data_delayed_85__1_, chained_data_delayed_85__0_ }),
    .data_o({ chained_data_delayed_86__127_, chained_data_delayed_86__126_, chained_data_delayed_86__125_, chained_data_delayed_86__124_, chained_data_delayed_86__123_, chained_data_delayed_86__122_, chained_data_delayed_86__121_, chained_data_delayed_86__120_, chained_data_delayed_86__119_, chained_data_delayed_86__118_, chained_data_delayed_86__117_, chained_data_delayed_86__116_, chained_data_delayed_86__115_, chained_data_delayed_86__114_, chained_data_delayed_86__113_, chained_data_delayed_86__112_, chained_data_delayed_86__111_, chained_data_delayed_86__110_, chained_data_delayed_86__109_, chained_data_delayed_86__108_, chained_data_delayed_86__107_, chained_data_delayed_86__106_, chained_data_delayed_86__105_, chained_data_delayed_86__104_, chained_data_delayed_86__103_, chained_data_delayed_86__102_, chained_data_delayed_86__101_, chained_data_delayed_86__100_, chained_data_delayed_86__99_, chained_data_delayed_86__98_, chained_data_delayed_86__97_, chained_data_delayed_86__96_, chained_data_delayed_86__95_, chained_data_delayed_86__94_, chained_data_delayed_86__93_, chained_data_delayed_86__92_, chained_data_delayed_86__91_, chained_data_delayed_86__90_, chained_data_delayed_86__89_, chained_data_delayed_86__88_, chained_data_delayed_86__87_, chained_data_delayed_86__86_, chained_data_delayed_86__85_, chained_data_delayed_86__84_, chained_data_delayed_86__83_, chained_data_delayed_86__82_, chained_data_delayed_86__81_, chained_data_delayed_86__80_, chained_data_delayed_86__79_, chained_data_delayed_86__78_, chained_data_delayed_86__77_, chained_data_delayed_86__76_, chained_data_delayed_86__75_, chained_data_delayed_86__74_, chained_data_delayed_86__73_, chained_data_delayed_86__72_, chained_data_delayed_86__71_, chained_data_delayed_86__70_, chained_data_delayed_86__69_, chained_data_delayed_86__68_, chained_data_delayed_86__67_, chained_data_delayed_86__66_, chained_data_delayed_86__65_, chained_data_delayed_86__64_, chained_data_delayed_86__63_, chained_data_delayed_86__62_, chained_data_delayed_86__61_, chained_data_delayed_86__60_, chained_data_delayed_86__59_, chained_data_delayed_86__58_, chained_data_delayed_86__57_, chained_data_delayed_86__56_, chained_data_delayed_86__55_, chained_data_delayed_86__54_, chained_data_delayed_86__53_, chained_data_delayed_86__52_, chained_data_delayed_86__51_, chained_data_delayed_86__50_, chained_data_delayed_86__49_, chained_data_delayed_86__48_, chained_data_delayed_86__47_, chained_data_delayed_86__46_, chained_data_delayed_86__45_, chained_data_delayed_86__44_, chained_data_delayed_86__43_, chained_data_delayed_86__42_, chained_data_delayed_86__41_, chained_data_delayed_86__40_, chained_data_delayed_86__39_, chained_data_delayed_86__38_, chained_data_delayed_86__37_, chained_data_delayed_86__36_, chained_data_delayed_86__35_, chained_data_delayed_86__34_, chained_data_delayed_86__33_, chained_data_delayed_86__32_, chained_data_delayed_86__31_, chained_data_delayed_86__30_, chained_data_delayed_86__29_, chained_data_delayed_86__28_, chained_data_delayed_86__27_, chained_data_delayed_86__26_, chained_data_delayed_86__25_, chained_data_delayed_86__24_, chained_data_delayed_86__23_, chained_data_delayed_86__22_, chained_data_delayed_86__21_, chained_data_delayed_86__20_, chained_data_delayed_86__19_, chained_data_delayed_86__18_, chained_data_delayed_86__17_, chained_data_delayed_86__16_, chained_data_delayed_86__15_, chained_data_delayed_86__14_, chained_data_delayed_86__13_, chained_data_delayed_86__12_, chained_data_delayed_86__11_, chained_data_delayed_86__10_, chained_data_delayed_86__9_, chained_data_delayed_86__8_, chained_data_delayed_86__7_, chained_data_delayed_86__6_, chained_data_delayed_86__5_, chained_data_delayed_86__4_, chained_data_delayed_86__3_, chained_data_delayed_86__2_, chained_data_delayed_86__1_, chained_data_delayed_86__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_87__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_86__127_, chained_data_delayed_86__126_, chained_data_delayed_86__125_, chained_data_delayed_86__124_, chained_data_delayed_86__123_, chained_data_delayed_86__122_, chained_data_delayed_86__121_, chained_data_delayed_86__120_, chained_data_delayed_86__119_, chained_data_delayed_86__118_, chained_data_delayed_86__117_, chained_data_delayed_86__116_, chained_data_delayed_86__115_, chained_data_delayed_86__114_, chained_data_delayed_86__113_, chained_data_delayed_86__112_, chained_data_delayed_86__111_, chained_data_delayed_86__110_, chained_data_delayed_86__109_, chained_data_delayed_86__108_, chained_data_delayed_86__107_, chained_data_delayed_86__106_, chained_data_delayed_86__105_, chained_data_delayed_86__104_, chained_data_delayed_86__103_, chained_data_delayed_86__102_, chained_data_delayed_86__101_, chained_data_delayed_86__100_, chained_data_delayed_86__99_, chained_data_delayed_86__98_, chained_data_delayed_86__97_, chained_data_delayed_86__96_, chained_data_delayed_86__95_, chained_data_delayed_86__94_, chained_data_delayed_86__93_, chained_data_delayed_86__92_, chained_data_delayed_86__91_, chained_data_delayed_86__90_, chained_data_delayed_86__89_, chained_data_delayed_86__88_, chained_data_delayed_86__87_, chained_data_delayed_86__86_, chained_data_delayed_86__85_, chained_data_delayed_86__84_, chained_data_delayed_86__83_, chained_data_delayed_86__82_, chained_data_delayed_86__81_, chained_data_delayed_86__80_, chained_data_delayed_86__79_, chained_data_delayed_86__78_, chained_data_delayed_86__77_, chained_data_delayed_86__76_, chained_data_delayed_86__75_, chained_data_delayed_86__74_, chained_data_delayed_86__73_, chained_data_delayed_86__72_, chained_data_delayed_86__71_, chained_data_delayed_86__70_, chained_data_delayed_86__69_, chained_data_delayed_86__68_, chained_data_delayed_86__67_, chained_data_delayed_86__66_, chained_data_delayed_86__65_, chained_data_delayed_86__64_, chained_data_delayed_86__63_, chained_data_delayed_86__62_, chained_data_delayed_86__61_, chained_data_delayed_86__60_, chained_data_delayed_86__59_, chained_data_delayed_86__58_, chained_data_delayed_86__57_, chained_data_delayed_86__56_, chained_data_delayed_86__55_, chained_data_delayed_86__54_, chained_data_delayed_86__53_, chained_data_delayed_86__52_, chained_data_delayed_86__51_, chained_data_delayed_86__50_, chained_data_delayed_86__49_, chained_data_delayed_86__48_, chained_data_delayed_86__47_, chained_data_delayed_86__46_, chained_data_delayed_86__45_, chained_data_delayed_86__44_, chained_data_delayed_86__43_, chained_data_delayed_86__42_, chained_data_delayed_86__41_, chained_data_delayed_86__40_, chained_data_delayed_86__39_, chained_data_delayed_86__38_, chained_data_delayed_86__37_, chained_data_delayed_86__36_, chained_data_delayed_86__35_, chained_data_delayed_86__34_, chained_data_delayed_86__33_, chained_data_delayed_86__32_, chained_data_delayed_86__31_, chained_data_delayed_86__30_, chained_data_delayed_86__29_, chained_data_delayed_86__28_, chained_data_delayed_86__27_, chained_data_delayed_86__26_, chained_data_delayed_86__25_, chained_data_delayed_86__24_, chained_data_delayed_86__23_, chained_data_delayed_86__22_, chained_data_delayed_86__21_, chained_data_delayed_86__20_, chained_data_delayed_86__19_, chained_data_delayed_86__18_, chained_data_delayed_86__17_, chained_data_delayed_86__16_, chained_data_delayed_86__15_, chained_data_delayed_86__14_, chained_data_delayed_86__13_, chained_data_delayed_86__12_, chained_data_delayed_86__11_, chained_data_delayed_86__10_, chained_data_delayed_86__9_, chained_data_delayed_86__8_, chained_data_delayed_86__7_, chained_data_delayed_86__6_, chained_data_delayed_86__5_, chained_data_delayed_86__4_, chained_data_delayed_86__3_, chained_data_delayed_86__2_, chained_data_delayed_86__1_, chained_data_delayed_86__0_ }),
    .data_o({ chained_data_delayed_87__127_, chained_data_delayed_87__126_, chained_data_delayed_87__125_, chained_data_delayed_87__124_, chained_data_delayed_87__123_, chained_data_delayed_87__122_, chained_data_delayed_87__121_, chained_data_delayed_87__120_, chained_data_delayed_87__119_, chained_data_delayed_87__118_, chained_data_delayed_87__117_, chained_data_delayed_87__116_, chained_data_delayed_87__115_, chained_data_delayed_87__114_, chained_data_delayed_87__113_, chained_data_delayed_87__112_, chained_data_delayed_87__111_, chained_data_delayed_87__110_, chained_data_delayed_87__109_, chained_data_delayed_87__108_, chained_data_delayed_87__107_, chained_data_delayed_87__106_, chained_data_delayed_87__105_, chained_data_delayed_87__104_, chained_data_delayed_87__103_, chained_data_delayed_87__102_, chained_data_delayed_87__101_, chained_data_delayed_87__100_, chained_data_delayed_87__99_, chained_data_delayed_87__98_, chained_data_delayed_87__97_, chained_data_delayed_87__96_, chained_data_delayed_87__95_, chained_data_delayed_87__94_, chained_data_delayed_87__93_, chained_data_delayed_87__92_, chained_data_delayed_87__91_, chained_data_delayed_87__90_, chained_data_delayed_87__89_, chained_data_delayed_87__88_, chained_data_delayed_87__87_, chained_data_delayed_87__86_, chained_data_delayed_87__85_, chained_data_delayed_87__84_, chained_data_delayed_87__83_, chained_data_delayed_87__82_, chained_data_delayed_87__81_, chained_data_delayed_87__80_, chained_data_delayed_87__79_, chained_data_delayed_87__78_, chained_data_delayed_87__77_, chained_data_delayed_87__76_, chained_data_delayed_87__75_, chained_data_delayed_87__74_, chained_data_delayed_87__73_, chained_data_delayed_87__72_, chained_data_delayed_87__71_, chained_data_delayed_87__70_, chained_data_delayed_87__69_, chained_data_delayed_87__68_, chained_data_delayed_87__67_, chained_data_delayed_87__66_, chained_data_delayed_87__65_, chained_data_delayed_87__64_, chained_data_delayed_87__63_, chained_data_delayed_87__62_, chained_data_delayed_87__61_, chained_data_delayed_87__60_, chained_data_delayed_87__59_, chained_data_delayed_87__58_, chained_data_delayed_87__57_, chained_data_delayed_87__56_, chained_data_delayed_87__55_, chained_data_delayed_87__54_, chained_data_delayed_87__53_, chained_data_delayed_87__52_, chained_data_delayed_87__51_, chained_data_delayed_87__50_, chained_data_delayed_87__49_, chained_data_delayed_87__48_, chained_data_delayed_87__47_, chained_data_delayed_87__46_, chained_data_delayed_87__45_, chained_data_delayed_87__44_, chained_data_delayed_87__43_, chained_data_delayed_87__42_, chained_data_delayed_87__41_, chained_data_delayed_87__40_, chained_data_delayed_87__39_, chained_data_delayed_87__38_, chained_data_delayed_87__37_, chained_data_delayed_87__36_, chained_data_delayed_87__35_, chained_data_delayed_87__34_, chained_data_delayed_87__33_, chained_data_delayed_87__32_, chained_data_delayed_87__31_, chained_data_delayed_87__30_, chained_data_delayed_87__29_, chained_data_delayed_87__28_, chained_data_delayed_87__27_, chained_data_delayed_87__26_, chained_data_delayed_87__25_, chained_data_delayed_87__24_, chained_data_delayed_87__23_, chained_data_delayed_87__22_, chained_data_delayed_87__21_, chained_data_delayed_87__20_, chained_data_delayed_87__19_, chained_data_delayed_87__18_, chained_data_delayed_87__17_, chained_data_delayed_87__16_, chained_data_delayed_87__15_, chained_data_delayed_87__14_, chained_data_delayed_87__13_, chained_data_delayed_87__12_, chained_data_delayed_87__11_, chained_data_delayed_87__10_, chained_data_delayed_87__9_, chained_data_delayed_87__8_, chained_data_delayed_87__7_, chained_data_delayed_87__6_, chained_data_delayed_87__5_, chained_data_delayed_87__4_, chained_data_delayed_87__3_, chained_data_delayed_87__2_, chained_data_delayed_87__1_, chained_data_delayed_87__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_88__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_87__127_, chained_data_delayed_87__126_, chained_data_delayed_87__125_, chained_data_delayed_87__124_, chained_data_delayed_87__123_, chained_data_delayed_87__122_, chained_data_delayed_87__121_, chained_data_delayed_87__120_, chained_data_delayed_87__119_, chained_data_delayed_87__118_, chained_data_delayed_87__117_, chained_data_delayed_87__116_, chained_data_delayed_87__115_, chained_data_delayed_87__114_, chained_data_delayed_87__113_, chained_data_delayed_87__112_, chained_data_delayed_87__111_, chained_data_delayed_87__110_, chained_data_delayed_87__109_, chained_data_delayed_87__108_, chained_data_delayed_87__107_, chained_data_delayed_87__106_, chained_data_delayed_87__105_, chained_data_delayed_87__104_, chained_data_delayed_87__103_, chained_data_delayed_87__102_, chained_data_delayed_87__101_, chained_data_delayed_87__100_, chained_data_delayed_87__99_, chained_data_delayed_87__98_, chained_data_delayed_87__97_, chained_data_delayed_87__96_, chained_data_delayed_87__95_, chained_data_delayed_87__94_, chained_data_delayed_87__93_, chained_data_delayed_87__92_, chained_data_delayed_87__91_, chained_data_delayed_87__90_, chained_data_delayed_87__89_, chained_data_delayed_87__88_, chained_data_delayed_87__87_, chained_data_delayed_87__86_, chained_data_delayed_87__85_, chained_data_delayed_87__84_, chained_data_delayed_87__83_, chained_data_delayed_87__82_, chained_data_delayed_87__81_, chained_data_delayed_87__80_, chained_data_delayed_87__79_, chained_data_delayed_87__78_, chained_data_delayed_87__77_, chained_data_delayed_87__76_, chained_data_delayed_87__75_, chained_data_delayed_87__74_, chained_data_delayed_87__73_, chained_data_delayed_87__72_, chained_data_delayed_87__71_, chained_data_delayed_87__70_, chained_data_delayed_87__69_, chained_data_delayed_87__68_, chained_data_delayed_87__67_, chained_data_delayed_87__66_, chained_data_delayed_87__65_, chained_data_delayed_87__64_, chained_data_delayed_87__63_, chained_data_delayed_87__62_, chained_data_delayed_87__61_, chained_data_delayed_87__60_, chained_data_delayed_87__59_, chained_data_delayed_87__58_, chained_data_delayed_87__57_, chained_data_delayed_87__56_, chained_data_delayed_87__55_, chained_data_delayed_87__54_, chained_data_delayed_87__53_, chained_data_delayed_87__52_, chained_data_delayed_87__51_, chained_data_delayed_87__50_, chained_data_delayed_87__49_, chained_data_delayed_87__48_, chained_data_delayed_87__47_, chained_data_delayed_87__46_, chained_data_delayed_87__45_, chained_data_delayed_87__44_, chained_data_delayed_87__43_, chained_data_delayed_87__42_, chained_data_delayed_87__41_, chained_data_delayed_87__40_, chained_data_delayed_87__39_, chained_data_delayed_87__38_, chained_data_delayed_87__37_, chained_data_delayed_87__36_, chained_data_delayed_87__35_, chained_data_delayed_87__34_, chained_data_delayed_87__33_, chained_data_delayed_87__32_, chained_data_delayed_87__31_, chained_data_delayed_87__30_, chained_data_delayed_87__29_, chained_data_delayed_87__28_, chained_data_delayed_87__27_, chained_data_delayed_87__26_, chained_data_delayed_87__25_, chained_data_delayed_87__24_, chained_data_delayed_87__23_, chained_data_delayed_87__22_, chained_data_delayed_87__21_, chained_data_delayed_87__20_, chained_data_delayed_87__19_, chained_data_delayed_87__18_, chained_data_delayed_87__17_, chained_data_delayed_87__16_, chained_data_delayed_87__15_, chained_data_delayed_87__14_, chained_data_delayed_87__13_, chained_data_delayed_87__12_, chained_data_delayed_87__11_, chained_data_delayed_87__10_, chained_data_delayed_87__9_, chained_data_delayed_87__8_, chained_data_delayed_87__7_, chained_data_delayed_87__6_, chained_data_delayed_87__5_, chained_data_delayed_87__4_, chained_data_delayed_87__3_, chained_data_delayed_87__2_, chained_data_delayed_87__1_, chained_data_delayed_87__0_ }),
    .data_o({ chained_data_delayed_88__127_, chained_data_delayed_88__126_, chained_data_delayed_88__125_, chained_data_delayed_88__124_, chained_data_delayed_88__123_, chained_data_delayed_88__122_, chained_data_delayed_88__121_, chained_data_delayed_88__120_, chained_data_delayed_88__119_, chained_data_delayed_88__118_, chained_data_delayed_88__117_, chained_data_delayed_88__116_, chained_data_delayed_88__115_, chained_data_delayed_88__114_, chained_data_delayed_88__113_, chained_data_delayed_88__112_, chained_data_delayed_88__111_, chained_data_delayed_88__110_, chained_data_delayed_88__109_, chained_data_delayed_88__108_, chained_data_delayed_88__107_, chained_data_delayed_88__106_, chained_data_delayed_88__105_, chained_data_delayed_88__104_, chained_data_delayed_88__103_, chained_data_delayed_88__102_, chained_data_delayed_88__101_, chained_data_delayed_88__100_, chained_data_delayed_88__99_, chained_data_delayed_88__98_, chained_data_delayed_88__97_, chained_data_delayed_88__96_, chained_data_delayed_88__95_, chained_data_delayed_88__94_, chained_data_delayed_88__93_, chained_data_delayed_88__92_, chained_data_delayed_88__91_, chained_data_delayed_88__90_, chained_data_delayed_88__89_, chained_data_delayed_88__88_, chained_data_delayed_88__87_, chained_data_delayed_88__86_, chained_data_delayed_88__85_, chained_data_delayed_88__84_, chained_data_delayed_88__83_, chained_data_delayed_88__82_, chained_data_delayed_88__81_, chained_data_delayed_88__80_, chained_data_delayed_88__79_, chained_data_delayed_88__78_, chained_data_delayed_88__77_, chained_data_delayed_88__76_, chained_data_delayed_88__75_, chained_data_delayed_88__74_, chained_data_delayed_88__73_, chained_data_delayed_88__72_, chained_data_delayed_88__71_, chained_data_delayed_88__70_, chained_data_delayed_88__69_, chained_data_delayed_88__68_, chained_data_delayed_88__67_, chained_data_delayed_88__66_, chained_data_delayed_88__65_, chained_data_delayed_88__64_, chained_data_delayed_88__63_, chained_data_delayed_88__62_, chained_data_delayed_88__61_, chained_data_delayed_88__60_, chained_data_delayed_88__59_, chained_data_delayed_88__58_, chained_data_delayed_88__57_, chained_data_delayed_88__56_, chained_data_delayed_88__55_, chained_data_delayed_88__54_, chained_data_delayed_88__53_, chained_data_delayed_88__52_, chained_data_delayed_88__51_, chained_data_delayed_88__50_, chained_data_delayed_88__49_, chained_data_delayed_88__48_, chained_data_delayed_88__47_, chained_data_delayed_88__46_, chained_data_delayed_88__45_, chained_data_delayed_88__44_, chained_data_delayed_88__43_, chained_data_delayed_88__42_, chained_data_delayed_88__41_, chained_data_delayed_88__40_, chained_data_delayed_88__39_, chained_data_delayed_88__38_, chained_data_delayed_88__37_, chained_data_delayed_88__36_, chained_data_delayed_88__35_, chained_data_delayed_88__34_, chained_data_delayed_88__33_, chained_data_delayed_88__32_, chained_data_delayed_88__31_, chained_data_delayed_88__30_, chained_data_delayed_88__29_, chained_data_delayed_88__28_, chained_data_delayed_88__27_, chained_data_delayed_88__26_, chained_data_delayed_88__25_, chained_data_delayed_88__24_, chained_data_delayed_88__23_, chained_data_delayed_88__22_, chained_data_delayed_88__21_, chained_data_delayed_88__20_, chained_data_delayed_88__19_, chained_data_delayed_88__18_, chained_data_delayed_88__17_, chained_data_delayed_88__16_, chained_data_delayed_88__15_, chained_data_delayed_88__14_, chained_data_delayed_88__13_, chained_data_delayed_88__12_, chained_data_delayed_88__11_, chained_data_delayed_88__10_, chained_data_delayed_88__9_, chained_data_delayed_88__8_, chained_data_delayed_88__7_, chained_data_delayed_88__6_, chained_data_delayed_88__5_, chained_data_delayed_88__4_, chained_data_delayed_88__3_, chained_data_delayed_88__2_, chained_data_delayed_88__1_, chained_data_delayed_88__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_89__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_88__127_, chained_data_delayed_88__126_, chained_data_delayed_88__125_, chained_data_delayed_88__124_, chained_data_delayed_88__123_, chained_data_delayed_88__122_, chained_data_delayed_88__121_, chained_data_delayed_88__120_, chained_data_delayed_88__119_, chained_data_delayed_88__118_, chained_data_delayed_88__117_, chained_data_delayed_88__116_, chained_data_delayed_88__115_, chained_data_delayed_88__114_, chained_data_delayed_88__113_, chained_data_delayed_88__112_, chained_data_delayed_88__111_, chained_data_delayed_88__110_, chained_data_delayed_88__109_, chained_data_delayed_88__108_, chained_data_delayed_88__107_, chained_data_delayed_88__106_, chained_data_delayed_88__105_, chained_data_delayed_88__104_, chained_data_delayed_88__103_, chained_data_delayed_88__102_, chained_data_delayed_88__101_, chained_data_delayed_88__100_, chained_data_delayed_88__99_, chained_data_delayed_88__98_, chained_data_delayed_88__97_, chained_data_delayed_88__96_, chained_data_delayed_88__95_, chained_data_delayed_88__94_, chained_data_delayed_88__93_, chained_data_delayed_88__92_, chained_data_delayed_88__91_, chained_data_delayed_88__90_, chained_data_delayed_88__89_, chained_data_delayed_88__88_, chained_data_delayed_88__87_, chained_data_delayed_88__86_, chained_data_delayed_88__85_, chained_data_delayed_88__84_, chained_data_delayed_88__83_, chained_data_delayed_88__82_, chained_data_delayed_88__81_, chained_data_delayed_88__80_, chained_data_delayed_88__79_, chained_data_delayed_88__78_, chained_data_delayed_88__77_, chained_data_delayed_88__76_, chained_data_delayed_88__75_, chained_data_delayed_88__74_, chained_data_delayed_88__73_, chained_data_delayed_88__72_, chained_data_delayed_88__71_, chained_data_delayed_88__70_, chained_data_delayed_88__69_, chained_data_delayed_88__68_, chained_data_delayed_88__67_, chained_data_delayed_88__66_, chained_data_delayed_88__65_, chained_data_delayed_88__64_, chained_data_delayed_88__63_, chained_data_delayed_88__62_, chained_data_delayed_88__61_, chained_data_delayed_88__60_, chained_data_delayed_88__59_, chained_data_delayed_88__58_, chained_data_delayed_88__57_, chained_data_delayed_88__56_, chained_data_delayed_88__55_, chained_data_delayed_88__54_, chained_data_delayed_88__53_, chained_data_delayed_88__52_, chained_data_delayed_88__51_, chained_data_delayed_88__50_, chained_data_delayed_88__49_, chained_data_delayed_88__48_, chained_data_delayed_88__47_, chained_data_delayed_88__46_, chained_data_delayed_88__45_, chained_data_delayed_88__44_, chained_data_delayed_88__43_, chained_data_delayed_88__42_, chained_data_delayed_88__41_, chained_data_delayed_88__40_, chained_data_delayed_88__39_, chained_data_delayed_88__38_, chained_data_delayed_88__37_, chained_data_delayed_88__36_, chained_data_delayed_88__35_, chained_data_delayed_88__34_, chained_data_delayed_88__33_, chained_data_delayed_88__32_, chained_data_delayed_88__31_, chained_data_delayed_88__30_, chained_data_delayed_88__29_, chained_data_delayed_88__28_, chained_data_delayed_88__27_, chained_data_delayed_88__26_, chained_data_delayed_88__25_, chained_data_delayed_88__24_, chained_data_delayed_88__23_, chained_data_delayed_88__22_, chained_data_delayed_88__21_, chained_data_delayed_88__20_, chained_data_delayed_88__19_, chained_data_delayed_88__18_, chained_data_delayed_88__17_, chained_data_delayed_88__16_, chained_data_delayed_88__15_, chained_data_delayed_88__14_, chained_data_delayed_88__13_, chained_data_delayed_88__12_, chained_data_delayed_88__11_, chained_data_delayed_88__10_, chained_data_delayed_88__9_, chained_data_delayed_88__8_, chained_data_delayed_88__7_, chained_data_delayed_88__6_, chained_data_delayed_88__5_, chained_data_delayed_88__4_, chained_data_delayed_88__3_, chained_data_delayed_88__2_, chained_data_delayed_88__1_, chained_data_delayed_88__0_ }),
    .data_o({ chained_data_delayed_89__127_, chained_data_delayed_89__126_, chained_data_delayed_89__125_, chained_data_delayed_89__124_, chained_data_delayed_89__123_, chained_data_delayed_89__122_, chained_data_delayed_89__121_, chained_data_delayed_89__120_, chained_data_delayed_89__119_, chained_data_delayed_89__118_, chained_data_delayed_89__117_, chained_data_delayed_89__116_, chained_data_delayed_89__115_, chained_data_delayed_89__114_, chained_data_delayed_89__113_, chained_data_delayed_89__112_, chained_data_delayed_89__111_, chained_data_delayed_89__110_, chained_data_delayed_89__109_, chained_data_delayed_89__108_, chained_data_delayed_89__107_, chained_data_delayed_89__106_, chained_data_delayed_89__105_, chained_data_delayed_89__104_, chained_data_delayed_89__103_, chained_data_delayed_89__102_, chained_data_delayed_89__101_, chained_data_delayed_89__100_, chained_data_delayed_89__99_, chained_data_delayed_89__98_, chained_data_delayed_89__97_, chained_data_delayed_89__96_, chained_data_delayed_89__95_, chained_data_delayed_89__94_, chained_data_delayed_89__93_, chained_data_delayed_89__92_, chained_data_delayed_89__91_, chained_data_delayed_89__90_, chained_data_delayed_89__89_, chained_data_delayed_89__88_, chained_data_delayed_89__87_, chained_data_delayed_89__86_, chained_data_delayed_89__85_, chained_data_delayed_89__84_, chained_data_delayed_89__83_, chained_data_delayed_89__82_, chained_data_delayed_89__81_, chained_data_delayed_89__80_, chained_data_delayed_89__79_, chained_data_delayed_89__78_, chained_data_delayed_89__77_, chained_data_delayed_89__76_, chained_data_delayed_89__75_, chained_data_delayed_89__74_, chained_data_delayed_89__73_, chained_data_delayed_89__72_, chained_data_delayed_89__71_, chained_data_delayed_89__70_, chained_data_delayed_89__69_, chained_data_delayed_89__68_, chained_data_delayed_89__67_, chained_data_delayed_89__66_, chained_data_delayed_89__65_, chained_data_delayed_89__64_, chained_data_delayed_89__63_, chained_data_delayed_89__62_, chained_data_delayed_89__61_, chained_data_delayed_89__60_, chained_data_delayed_89__59_, chained_data_delayed_89__58_, chained_data_delayed_89__57_, chained_data_delayed_89__56_, chained_data_delayed_89__55_, chained_data_delayed_89__54_, chained_data_delayed_89__53_, chained_data_delayed_89__52_, chained_data_delayed_89__51_, chained_data_delayed_89__50_, chained_data_delayed_89__49_, chained_data_delayed_89__48_, chained_data_delayed_89__47_, chained_data_delayed_89__46_, chained_data_delayed_89__45_, chained_data_delayed_89__44_, chained_data_delayed_89__43_, chained_data_delayed_89__42_, chained_data_delayed_89__41_, chained_data_delayed_89__40_, chained_data_delayed_89__39_, chained_data_delayed_89__38_, chained_data_delayed_89__37_, chained_data_delayed_89__36_, chained_data_delayed_89__35_, chained_data_delayed_89__34_, chained_data_delayed_89__33_, chained_data_delayed_89__32_, chained_data_delayed_89__31_, chained_data_delayed_89__30_, chained_data_delayed_89__29_, chained_data_delayed_89__28_, chained_data_delayed_89__27_, chained_data_delayed_89__26_, chained_data_delayed_89__25_, chained_data_delayed_89__24_, chained_data_delayed_89__23_, chained_data_delayed_89__22_, chained_data_delayed_89__21_, chained_data_delayed_89__20_, chained_data_delayed_89__19_, chained_data_delayed_89__18_, chained_data_delayed_89__17_, chained_data_delayed_89__16_, chained_data_delayed_89__15_, chained_data_delayed_89__14_, chained_data_delayed_89__13_, chained_data_delayed_89__12_, chained_data_delayed_89__11_, chained_data_delayed_89__10_, chained_data_delayed_89__9_, chained_data_delayed_89__8_, chained_data_delayed_89__7_, chained_data_delayed_89__6_, chained_data_delayed_89__5_, chained_data_delayed_89__4_, chained_data_delayed_89__3_, chained_data_delayed_89__2_, chained_data_delayed_89__1_, chained_data_delayed_89__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_90__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_89__127_, chained_data_delayed_89__126_, chained_data_delayed_89__125_, chained_data_delayed_89__124_, chained_data_delayed_89__123_, chained_data_delayed_89__122_, chained_data_delayed_89__121_, chained_data_delayed_89__120_, chained_data_delayed_89__119_, chained_data_delayed_89__118_, chained_data_delayed_89__117_, chained_data_delayed_89__116_, chained_data_delayed_89__115_, chained_data_delayed_89__114_, chained_data_delayed_89__113_, chained_data_delayed_89__112_, chained_data_delayed_89__111_, chained_data_delayed_89__110_, chained_data_delayed_89__109_, chained_data_delayed_89__108_, chained_data_delayed_89__107_, chained_data_delayed_89__106_, chained_data_delayed_89__105_, chained_data_delayed_89__104_, chained_data_delayed_89__103_, chained_data_delayed_89__102_, chained_data_delayed_89__101_, chained_data_delayed_89__100_, chained_data_delayed_89__99_, chained_data_delayed_89__98_, chained_data_delayed_89__97_, chained_data_delayed_89__96_, chained_data_delayed_89__95_, chained_data_delayed_89__94_, chained_data_delayed_89__93_, chained_data_delayed_89__92_, chained_data_delayed_89__91_, chained_data_delayed_89__90_, chained_data_delayed_89__89_, chained_data_delayed_89__88_, chained_data_delayed_89__87_, chained_data_delayed_89__86_, chained_data_delayed_89__85_, chained_data_delayed_89__84_, chained_data_delayed_89__83_, chained_data_delayed_89__82_, chained_data_delayed_89__81_, chained_data_delayed_89__80_, chained_data_delayed_89__79_, chained_data_delayed_89__78_, chained_data_delayed_89__77_, chained_data_delayed_89__76_, chained_data_delayed_89__75_, chained_data_delayed_89__74_, chained_data_delayed_89__73_, chained_data_delayed_89__72_, chained_data_delayed_89__71_, chained_data_delayed_89__70_, chained_data_delayed_89__69_, chained_data_delayed_89__68_, chained_data_delayed_89__67_, chained_data_delayed_89__66_, chained_data_delayed_89__65_, chained_data_delayed_89__64_, chained_data_delayed_89__63_, chained_data_delayed_89__62_, chained_data_delayed_89__61_, chained_data_delayed_89__60_, chained_data_delayed_89__59_, chained_data_delayed_89__58_, chained_data_delayed_89__57_, chained_data_delayed_89__56_, chained_data_delayed_89__55_, chained_data_delayed_89__54_, chained_data_delayed_89__53_, chained_data_delayed_89__52_, chained_data_delayed_89__51_, chained_data_delayed_89__50_, chained_data_delayed_89__49_, chained_data_delayed_89__48_, chained_data_delayed_89__47_, chained_data_delayed_89__46_, chained_data_delayed_89__45_, chained_data_delayed_89__44_, chained_data_delayed_89__43_, chained_data_delayed_89__42_, chained_data_delayed_89__41_, chained_data_delayed_89__40_, chained_data_delayed_89__39_, chained_data_delayed_89__38_, chained_data_delayed_89__37_, chained_data_delayed_89__36_, chained_data_delayed_89__35_, chained_data_delayed_89__34_, chained_data_delayed_89__33_, chained_data_delayed_89__32_, chained_data_delayed_89__31_, chained_data_delayed_89__30_, chained_data_delayed_89__29_, chained_data_delayed_89__28_, chained_data_delayed_89__27_, chained_data_delayed_89__26_, chained_data_delayed_89__25_, chained_data_delayed_89__24_, chained_data_delayed_89__23_, chained_data_delayed_89__22_, chained_data_delayed_89__21_, chained_data_delayed_89__20_, chained_data_delayed_89__19_, chained_data_delayed_89__18_, chained_data_delayed_89__17_, chained_data_delayed_89__16_, chained_data_delayed_89__15_, chained_data_delayed_89__14_, chained_data_delayed_89__13_, chained_data_delayed_89__12_, chained_data_delayed_89__11_, chained_data_delayed_89__10_, chained_data_delayed_89__9_, chained_data_delayed_89__8_, chained_data_delayed_89__7_, chained_data_delayed_89__6_, chained_data_delayed_89__5_, chained_data_delayed_89__4_, chained_data_delayed_89__3_, chained_data_delayed_89__2_, chained_data_delayed_89__1_, chained_data_delayed_89__0_ }),
    .data_o({ chained_data_delayed_90__127_, chained_data_delayed_90__126_, chained_data_delayed_90__125_, chained_data_delayed_90__124_, chained_data_delayed_90__123_, chained_data_delayed_90__122_, chained_data_delayed_90__121_, chained_data_delayed_90__120_, chained_data_delayed_90__119_, chained_data_delayed_90__118_, chained_data_delayed_90__117_, chained_data_delayed_90__116_, chained_data_delayed_90__115_, chained_data_delayed_90__114_, chained_data_delayed_90__113_, chained_data_delayed_90__112_, chained_data_delayed_90__111_, chained_data_delayed_90__110_, chained_data_delayed_90__109_, chained_data_delayed_90__108_, chained_data_delayed_90__107_, chained_data_delayed_90__106_, chained_data_delayed_90__105_, chained_data_delayed_90__104_, chained_data_delayed_90__103_, chained_data_delayed_90__102_, chained_data_delayed_90__101_, chained_data_delayed_90__100_, chained_data_delayed_90__99_, chained_data_delayed_90__98_, chained_data_delayed_90__97_, chained_data_delayed_90__96_, chained_data_delayed_90__95_, chained_data_delayed_90__94_, chained_data_delayed_90__93_, chained_data_delayed_90__92_, chained_data_delayed_90__91_, chained_data_delayed_90__90_, chained_data_delayed_90__89_, chained_data_delayed_90__88_, chained_data_delayed_90__87_, chained_data_delayed_90__86_, chained_data_delayed_90__85_, chained_data_delayed_90__84_, chained_data_delayed_90__83_, chained_data_delayed_90__82_, chained_data_delayed_90__81_, chained_data_delayed_90__80_, chained_data_delayed_90__79_, chained_data_delayed_90__78_, chained_data_delayed_90__77_, chained_data_delayed_90__76_, chained_data_delayed_90__75_, chained_data_delayed_90__74_, chained_data_delayed_90__73_, chained_data_delayed_90__72_, chained_data_delayed_90__71_, chained_data_delayed_90__70_, chained_data_delayed_90__69_, chained_data_delayed_90__68_, chained_data_delayed_90__67_, chained_data_delayed_90__66_, chained_data_delayed_90__65_, chained_data_delayed_90__64_, chained_data_delayed_90__63_, chained_data_delayed_90__62_, chained_data_delayed_90__61_, chained_data_delayed_90__60_, chained_data_delayed_90__59_, chained_data_delayed_90__58_, chained_data_delayed_90__57_, chained_data_delayed_90__56_, chained_data_delayed_90__55_, chained_data_delayed_90__54_, chained_data_delayed_90__53_, chained_data_delayed_90__52_, chained_data_delayed_90__51_, chained_data_delayed_90__50_, chained_data_delayed_90__49_, chained_data_delayed_90__48_, chained_data_delayed_90__47_, chained_data_delayed_90__46_, chained_data_delayed_90__45_, chained_data_delayed_90__44_, chained_data_delayed_90__43_, chained_data_delayed_90__42_, chained_data_delayed_90__41_, chained_data_delayed_90__40_, chained_data_delayed_90__39_, chained_data_delayed_90__38_, chained_data_delayed_90__37_, chained_data_delayed_90__36_, chained_data_delayed_90__35_, chained_data_delayed_90__34_, chained_data_delayed_90__33_, chained_data_delayed_90__32_, chained_data_delayed_90__31_, chained_data_delayed_90__30_, chained_data_delayed_90__29_, chained_data_delayed_90__28_, chained_data_delayed_90__27_, chained_data_delayed_90__26_, chained_data_delayed_90__25_, chained_data_delayed_90__24_, chained_data_delayed_90__23_, chained_data_delayed_90__22_, chained_data_delayed_90__21_, chained_data_delayed_90__20_, chained_data_delayed_90__19_, chained_data_delayed_90__18_, chained_data_delayed_90__17_, chained_data_delayed_90__16_, chained_data_delayed_90__15_, chained_data_delayed_90__14_, chained_data_delayed_90__13_, chained_data_delayed_90__12_, chained_data_delayed_90__11_, chained_data_delayed_90__10_, chained_data_delayed_90__9_, chained_data_delayed_90__8_, chained_data_delayed_90__7_, chained_data_delayed_90__6_, chained_data_delayed_90__5_, chained_data_delayed_90__4_, chained_data_delayed_90__3_, chained_data_delayed_90__2_, chained_data_delayed_90__1_, chained_data_delayed_90__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_91__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_90__127_, chained_data_delayed_90__126_, chained_data_delayed_90__125_, chained_data_delayed_90__124_, chained_data_delayed_90__123_, chained_data_delayed_90__122_, chained_data_delayed_90__121_, chained_data_delayed_90__120_, chained_data_delayed_90__119_, chained_data_delayed_90__118_, chained_data_delayed_90__117_, chained_data_delayed_90__116_, chained_data_delayed_90__115_, chained_data_delayed_90__114_, chained_data_delayed_90__113_, chained_data_delayed_90__112_, chained_data_delayed_90__111_, chained_data_delayed_90__110_, chained_data_delayed_90__109_, chained_data_delayed_90__108_, chained_data_delayed_90__107_, chained_data_delayed_90__106_, chained_data_delayed_90__105_, chained_data_delayed_90__104_, chained_data_delayed_90__103_, chained_data_delayed_90__102_, chained_data_delayed_90__101_, chained_data_delayed_90__100_, chained_data_delayed_90__99_, chained_data_delayed_90__98_, chained_data_delayed_90__97_, chained_data_delayed_90__96_, chained_data_delayed_90__95_, chained_data_delayed_90__94_, chained_data_delayed_90__93_, chained_data_delayed_90__92_, chained_data_delayed_90__91_, chained_data_delayed_90__90_, chained_data_delayed_90__89_, chained_data_delayed_90__88_, chained_data_delayed_90__87_, chained_data_delayed_90__86_, chained_data_delayed_90__85_, chained_data_delayed_90__84_, chained_data_delayed_90__83_, chained_data_delayed_90__82_, chained_data_delayed_90__81_, chained_data_delayed_90__80_, chained_data_delayed_90__79_, chained_data_delayed_90__78_, chained_data_delayed_90__77_, chained_data_delayed_90__76_, chained_data_delayed_90__75_, chained_data_delayed_90__74_, chained_data_delayed_90__73_, chained_data_delayed_90__72_, chained_data_delayed_90__71_, chained_data_delayed_90__70_, chained_data_delayed_90__69_, chained_data_delayed_90__68_, chained_data_delayed_90__67_, chained_data_delayed_90__66_, chained_data_delayed_90__65_, chained_data_delayed_90__64_, chained_data_delayed_90__63_, chained_data_delayed_90__62_, chained_data_delayed_90__61_, chained_data_delayed_90__60_, chained_data_delayed_90__59_, chained_data_delayed_90__58_, chained_data_delayed_90__57_, chained_data_delayed_90__56_, chained_data_delayed_90__55_, chained_data_delayed_90__54_, chained_data_delayed_90__53_, chained_data_delayed_90__52_, chained_data_delayed_90__51_, chained_data_delayed_90__50_, chained_data_delayed_90__49_, chained_data_delayed_90__48_, chained_data_delayed_90__47_, chained_data_delayed_90__46_, chained_data_delayed_90__45_, chained_data_delayed_90__44_, chained_data_delayed_90__43_, chained_data_delayed_90__42_, chained_data_delayed_90__41_, chained_data_delayed_90__40_, chained_data_delayed_90__39_, chained_data_delayed_90__38_, chained_data_delayed_90__37_, chained_data_delayed_90__36_, chained_data_delayed_90__35_, chained_data_delayed_90__34_, chained_data_delayed_90__33_, chained_data_delayed_90__32_, chained_data_delayed_90__31_, chained_data_delayed_90__30_, chained_data_delayed_90__29_, chained_data_delayed_90__28_, chained_data_delayed_90__27_, chained_data_delayed_90__26_, chained_data_delayed_90__25_, chained_data_delayed_90__24_, chained_data_delayed_90__23_, chained_data_delayed_90__22_, chained_data_delayed_90__21_, chained_data_delayed_90__20_, chained_data_delayed_90__19_, chained_data_delayed_90__18_, chained_data_delayed_90__17_, chained_data_delayed_90__16_, chained_data_delayed_90__15_, chained_data_delayed_90__14_, chained_data_delayed_90__13_, chained_data_delayed_90__12_, chained_data_delayed_90__11_, chained_data_delayed_90__10_, chained_data_delayed_90__9_, chained_data_delayed_90__8_, chained_data_delayed_90__7_, chained_data_delayed_90__6_, chained_data_delayed_90__5_, chained_data_delayed_90__4_, chained_data_delayed_90__3_, chained_data_delayed_90__2_, chained_data_delayed_90__1_, chained_data_delayed_90__0_ }),
    .data_o({ chained_data_delayed_91__127_, chained_data_delayed_91__126_, chained_data_delayed_91__125_, chained_data_delayed_91__124_, chained_data_delayed_91__123_, chained_data_delayed_91__122_, chained_data_delayed_91__121_, chained_data_delayed_91__120_, chained_data_delayed_91__119_, chained_data_delayed_91__118_, chained_data_delayed_91__117_, chained_data_delayed_91__116_, chained_data_delayed_91__115_, chained_data_delayed_91__114_, chained_data_delayed_91__113_, chained_data_delayed_91__112_, chained_data_delayed_91__111_, chained_data_delayed_91__110_, chained_data_delayed_91__109_, chained_data_delayed_91__108_, chained_data_delayed_91__107_, chained_data_delayed_91__106_, chained_data_delayed_91__105_, chained_data_delayed_91__104_, chained_data_delayed_91__103_, chained_data_delayed_91__102_, chained_data_delayed_91__101_, chained_data_delayed_91__100_, chained_data_delayed_91__99_, chained_data_delayed_91__98_, chained_data_delayed_91__97_, chained_data_delayed_91__96_, chained_data_delayed_91__95_, chained_data_delayed_91__94_, chained_data_delayed_91__93_, chained_data_delayed_91__92_, chained_data_delayed_91__91_, chained_data_delayed_91__90_, chained_data_delayed_91__89_, chained_data_delayed_91__88_, chained_data_delayed_91__87_, chained_data_delayed_91__86_, chained_data_delayed_91__85_, chained_data_delayed_91__84_, chained_data_delayed_91__83_, chained_data_delayed_91__82_, chained_data_delayed_91__81_, chained_data_delayed_91__80_, chained_data_delayed_91__79_, chained_data_delayed_91__78_, chained_data_delayed_91__77_, chained_data_delayed_91__76_, chained_data_delayed_91__75_, chained_data_delayed_91__74_, chained_data_delayed_91__73_, chained_data_delayed_91__72_, chained_data_delayed_91__71_, chained_data_delayed_91__70_, chained_data_delayed_91__69_, chained_data_delayed_91__68_, chained_data_delayed_91__67_, chained_data_delayed_91__66_, chained_data_delayed_91__65_, chained_data_delayed_91__64_, chained_data_delayed_91__63_, chained_data_delayed_91__62_, chained_data_delayed_91__61_, chained_data_delayed_91__60_, chained_data_delayed_91__59_, chained_data_delayed_91__58_, chained_data_delayed_91__57_, chained_data_delayed_91__56_, chained_data_delayed_91__55_, chained_data_delayed_91__54_, chained_data_delayed_91__53_, chained_data_delayed_91__52_, chained_data_delayed_91__51_, chained_data_delayed_91__50_, chained_data_delayed_91__49_, chained_data_delayed_91__48_, chained_data_delayed_91__47_, chained_data_delayed_91__46_, chained_data_delayed_91__45_, chained_data_delayed_91__44_, chained_data_delayed_91__43_, chained_data_delayed_91__42_, chained_data_delayed_91__41_, chained_data_delayed_91__40_, chained_data_delayed_91__39_, chained_data_delayed_91__38_, chained_data_delayed_91__37_, chained_data_delayed_91__36_, chained_data_delayed_91__35_, chained_data_delayed_91__34_, chained_data_delayed_91__33_, chained_data_delayed_91__32_, chained_data_delayed_91__31_, chained_data_delayed_91__30_, chained_data_delayed_91__29_, chained_data_delayed_91__28_, chained_data_delayed_91__27_, chained_data_delayed_91__26_, chained_data_delayed_91__25_, chained_data_delayed_91__24_, chained_data_delayed_91__23_, chained_data_delayed_91__22_, chained_data_delayed_91__21_, chained_data_delayed_91__20_, chained_data_delayed_91__19_, chained_data_delayed_91__18_, chained_data_delayed_91__17_, chained_data_delayed_91__16_, chained_data_delayed_91__15_, chained_data_delayed_91__14_, chained_data_delayed_91__13_, chained_data_delayed_91__12_, chained_data_delayed_91__11_, chained_data_delayed_91__10_, chained_data_delayed_91__9_, chained_data_delayed_91__8_, chained_data_delayed_91__7_, chained_data_delayed_91__6_, chained_data_delayed_91__5_, chained_data_delayed_91__4_, chained_data_delayed_91__3_, chained_data_delayed_91__2_, chained_data_delayed_91__1_, chained_data_delayed_91__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_92__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_91__127_, chained_data_delayed_91__126_, chained_data_delayed_91__125_, chained_data_delayed_91__124_, chained_data_delayed_91__123_, chained_data_delayed_91__122_, chained_data_delayed_91__121_, chained_data_delayed_91__120_, chained_data_delayed_91__119_, chained_data_delayed_91__118_, chained_data_delayed_91__117_, chained_data_delayed_91__116_, chained_data_delayed_91__115_, chained_data_delayed_91__114_, chained_data_delayed_91__113_, chained_data_delayed_91__112_, chained_data_delayed_91__111_, chained_data_delayed_91__110_, chained_data_delayed_91__109_, chained_data_delayed_91__108_, chained_data_delayed_91__107_, chained_data_delayed_91__106_, chained_data_delayed_91__105_, chained_data_delayed_91__104_, chained_data_delayed_91__103_, chained_data_delayed_91__102_, chained_data_delayed_91__101_, chained_data_delayed_91__100_, chained_data_delayed_91__99_, chained_data_delayed_91__98_, chained_data_delayed_91__97_, chained_data_delayed_91__96_, chained_data_delayed_91__95_, chained_data_delayed_91__94_, chained_data_delayed_91__93_, chained_data_delayed_91__92_, chained_data_delayed_91__91_, chained_data_delayed_91__90_, chained_data_delayed_91__89_, chained_data_delayed_91__88_, chained_data_delayed_91__87_, chained_data_delayed_91__86_, chained_data_delayed_91__85_, chained_data_delayed_91__84_, chained_data_delayed_91__83_, chained_data_delayed_91__82_, chained_data_delayed_91__81_, chained_data_delayed_91__80_, chained_data_delayed_91__79_, chained_data_delayed_91__78_, chained_data_delayed_91__77_, chained_data_delayed_91__76_, chained_data_delayed_91__75_, chained_data_delayed_91__74_, chained_data_delayed_91__73_, chained_data_delayed_91__72_, chained_data_delayed_91__71_, chained_data_delayed_91__70_, chained_data_delayed_91__69_, chained_data_delayed_91__68_, chained_data_delayed_91__67_, chained_data_delayed_91__66_, chained_data_delayed_91__65_, chained_data_delayed_91__64_, chained_data_delayed_91__63_, chained_data_delayed_91__62_, chained_data_delayed_91__61_, chained_data_delayed_91__60_, chained_data_delayed_91__59_, chained_data_delayed_91__58_, chained_data_delayed_91__57_, chained_data_delayed_91__56_, chained_data_delayed_91__55_, chained_data_delayed_91__54_, chained_data_delayed_91__53_, chained_data_delayed_91__52_, chained_data_delayed_91__51_, chained_data_delayed_91__50_, chained_data_delayed_91__49_, chained_data_delayed_91__48_, chained_data_delayed_91__47_, chained_data_delayed_91__46_, chained_data_delayed_91__45_, chained_data_delayed_91__44_, chained_data_delayed_91__43_, chained_data_delayed_91__42_, chained_data_delayed_91__41_, chained_data_delayed_91__40_, chained_data_delayed_91__39_, chained_data_delayed_91__38_, chained_data_delayed_91__37_, chained_data_delayed_91__36_, chained_data_delayed_91__35_, chained_data_delayed_91__34_, chained_data_delayed_91__33_, chained_data_delayed_91__32_, chained_data_delayed_91__31_, chained_data_delayed_91__30_, chained_data_delayed_91__29_, chained_data_delayed_91__28_, chained_data_delayed_91__27_, chained_data_delayed_91__26_, chained_data_delayed_91__25_, chained_data_delayed_91__24_, chained_data_delayed_91__23_, chained_data_delayed_91__22_, chained_data_delayed_91__21_, chained_data_delayed_91__20_, chained_data_delayed_91__19_, chained_data_delayed_91__18_, chained_data_delayed_91__17_, chained_data_delayed_91__16_, chained_data_delayed_91__15_, chained_data_delayed_91__14_, chained_data_delayed_91__13_, chained_data_delayed_91__12_, chained_data_delayed_91__11_, chained_data_delayed_91__10_, chained_data_delayed_91__9_, chained_data_delayed_91__8_, chained_data_delayed_91__7_, chained_data_delayed_91__6_, chained_data_delayed_91__5_, chained_data_delayed_91__4_, chained_data_delayed_91__3_, chained_data_delayed_91__2_, chained_data_delayed_91__1_, chained_data_delayed_91__0_ }),
    .data_o({ chained_data_delayed_92__127_, chained_data_delayed_92__126_, chained_data_delayed_92__125_, chained_data_delayed_92__124_, chained_data_delayed_92__123_, chained_data_delayed_92__122_, chained_data_delayed_92__121_, chained_data_delayed_92__120_, chained_data_delayed_92__119_, chained_data_delayed_92__118_, chained_data_delayed_92__117_, chained_data_delayed_92__116_, chained_data_delayed_92__115_, chained_data_delayed_92__114_, chained_data_delayed_92__113_, chained_data_delayed_92__112_, chained_data_delayed_92__111_, chained_data_delayed_92__110_, chained_data_delayed_92__109_, chained_data_delayed_92__108_, chained_data_delayed_92__107_, chained_data_delayed_92__106_, chained_data_delayed_92__105_, chained_data_delayed_92__104_, chained_data_delayed_92__103_, chained_data_delayed_92__102_, chained_data_delayed_92__101_, chained_data_delayed_92__100_, chained_data_delayed_92__99_, chained_data_delayed_92__98_, chained_data_delayed_92__97_, chained_data_delayed_92__96_, chained_data_delayed_92__95_, chained_data_delayed_92__94_, chained_data_delayed_92__93_, chained_data_delayed_92__92_, chained_data_delayed_92__91_, chained_data_delayed_92__90_, chained_data_delayed_92__89_, chained_data_delayed_92__88_, chained_data_delayed_92__87_, chained_data_delayed_92__86_, chained_data_delayed_92__85_, chained_data_delayed_92__84_, chained_data_delayed_92__83_, chained_data_delayed_92__82_, chained_data_delayed_92__81_, chained_data_delayed_92__80_, chained_data_delayed_92__79_, chained_data_delayed_92__78_, chained_data_delayed_92__77_, chained_data_delayed_92__76_, chained_data_delayed_92__75_, chained_data_delayed_92__74_, chained_data_delayed_92__73_, chained_data_delayed_92__72_, chained_data_delayed_92__71_, chained_data_delayed_92__70_, chained_data_delayed_92__69_, chained_data_delayed_92__68_, chained_data_delayed_92__67_, chained_data_delayed_92__66_, chained_data_delayed_92__65_, chained_data_delayed_92__64_, chained_data_delayed_92__63_, chained_data_delayed_92__62_, chained_data_delayed_92__61_, chained_data_delayed_92__60_, chained_data_delayed_92__59_, chained_data_delayed_92__58_, chained_data_delayed_92__57_, chained_data_delayed_92__56_, chained_data_delayed_92__55_, chained_data_delayed_92__54_, chained_data_delayed_92__53_, chained_data_delayed_92__52_, chained_data_delayed_92__51_, chained_data_delayed_92__50_, chained_data_delayed_92__49_, chained_data_delayed_92__48_, chained_data_delayed_92__47_, chained_data_delayed_92__46_, chained_data_delayed_92__45_, chained_data_delayed_92__44_, chained_data_delayed_92__43_, chained_data_delayed_92__42_, chained_data_delayed_92__41_, chained_data_delayed_92__40_, chained_data_delayed_92__39_, chained_data_delayed_92__38_, chained_data_delayed_92__37_, chained_data_delayed_92__36_, chained_data_delayed_92__35_, chained_data_delayed_92__34_, chained_data_delayed_92__33_, chained_data_delayed_92__32_, chained_data_delayed_92__31_, chained_data_delayed_92__30_, chained_data_delayed_92__29_, chained_data_delayed_92__28_, chained_data_delayed_92__27_, chained_data_delayed_92__26_, chained_data_delayed_92__25_, chained_data_delayed_92__24_, chained_data_delayed_92__23_, chained_data_delayed_92__22_, chained_data_delayed_92__21_, chained_data_delayed_92__20_, chained_data_delayed_92__19_, chained_data_delayed_92__18_, chained_data_delayed_92__17_, chained_data_delayed_92__16_, chained_data_delayed_92__15_, chained_data_delayed_92__14_, chained_data_delayed_92__13_, chained_data_delayed_92__12_, chained_data_delayed_92__11_, chained_data_delayed_92__10_, chained_data_delayed_92__9_, chained_data_delayed_92__8_, chained_data_delayed_92__7_, chained_data_delayed_92__6_, chained_data_delayed_92__5_, chained_data_delayed_92__4_, chained_data_delayed_92__3_, chained_data_delayed_92__2_, chained_data_delayed_92__1_, chained_data_delayed_92__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_93__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_92__127_, chained_data_delayed_92__126_, chained_data_delayed_92__125_, chained_data_delayed_92__124_, chained_data_delayed_92__123_, chained_data_delayed_92__122_, chained_data_delayed_92__121_, chained_data_delayed_92__120_, chained_data_delayed_92__119_, chained_data_delayed_92__118_, chained_data_delayed_92__117_, chained_data_delayed_92__116_, chained_data_delayed_92__115_, chained_data_delayed_92__114_, chained_data_delayed_92__113_, chained_data_delayed_92__112_, chained_data_delayed_92__111_, chained_data_delayed_92__110_, chained_data_delayed_92__109_, chained_data_delayed_92__108_, chained_data_delayed_92__107_, chained_data_delayed_92__106_, chained_data_delayed_92__105_, chained_data_delayed_92__104_, chained_data_delayed_92__103_, chained_data_delayed_92__102_, chained_data_delayed_92__101_, chained_data_delayed_92__100_, chained_data_delayed_92__99_, chained_data_delayed_92__98_, chained_data_delayed_92__97_, chained_data_delayed_92__96_, chained_data_delayed_92__95_, chained_data_delayed_92__94_, chained_data_delayed_92__93_, chained_data_delayed_92__92_, chained_data_delayed_92__91_, chained_data_delayed_92__90_, chained_data_delayed_92__89_, chained_data_delayed_92__88_, chained_data_delayed_92__87_, chained_data_delayed_92__86_, chained_data_delayed_92__85_, chained_data_delayed_92__84_, chained_data_delayed_92__83_, chained_data_delayed_92__82_, chained_data_delayed_92__81_, chained_data_delayed_92__80_, chained_data_delayed_92__79_, chained_data_delayed_92__78_, chained_data_delayed_92__77_, chained_data_delayed_92__76_, chained_data_delayed_92__75_, chained_data_delayed_92__74_, chained_data_delayed_92__73_, chained_data_delayed_92__72_, chained_data_delayed_92__71_, chained_data_delayed_92__70_, chained_data_delayed_92__69_, chained_data_delayed_92__68_, chained_data_delayed_92__67_, chained_data_delayed_92__66_, chained_data_delayed_92__65_, chained_data_delayed_92__64_, chained_data_delayed_92__63_, chained_data_delayed_92__62_, chained_data_delayed_92__61_, chained_data_delayed_92__60_, chained_data_delayed_92__59_, chained_data_delayed_92__58_, chained_data_delayed_92__57_, chained_data_delayed_92__56_, chained_data_delayed_92__55_, chained_data_delayed_92__54_, chained_data_delayed_92__53_, chained_data_delayed_92__52_, chained_data_delayed_92__51_, chained_data_delayed_92__50_, chained_data_delayed_92__49_, chained_data_delayed_92__48_, chained_data_delayed_92__47_, chained_data_delayed_92__46_, chained_data_delayed_92__45_, chained_data_delayed_92__44_, chained_data_delayed_92__43_, chained_data_delayed_92__42_, chained_data_delayed_92__41_, chained_data_delayed_92__40_, chained_data_delayed_92__39_, chained_data_delayed_92__38_, chained_data_delayed_92__37_, chained_data_delayed_92__36_, chained_data_delayed_92__35_, chained_data_delayed_92__34_, chained_data_delayed_92__33_, chained_data_delayed_92__32_, chained_data_delayed_92__31_, chained_data_delayed_92__30_, chained_data_delayed_92__29_, chained_data_delayed_92__28_, chained_data_delayed_92__27_, chained_data_delayed_92__26_, chained_data_delayed_92__25_, chained_data_delayed_92__24_, chained_data_delayed_92__23_, chained_data_delayed_92__22_, chained_data_delayed_92__21_, chained_data_delayed_92__20_, chained_data_delayed_92__19_, chained_data_delayed_92__18_, chained_data_delayed_92__17_, chained_data_delayed_92__16_, chained_data_delayed_92__15_, chained_data_delayed_92__14_, chained_data_delayed_92__13_, chained_data_delayed_92__12_, chained_data_delayed_92__11_, chained_data_delayed_92__10_, chained_data_delayed_92__9_, chained_data_delayed_92__8_, chained_data_delayed_92__7_, chained_data_delayed_92__6_, chained_data_delayed_92__5_, chained_data_delayed_92__4_, chained_data_delayed_92__3_, chained_data_delayed_92__2_, chained_data_delayed_92__1_, chained_data_delayed_92__0_ }),
    .data_o({ chained_data_delayed_93__127_, chained_data_delayed_93__126_, chained_data_delayed_93__125_, chained_data_delayed_93__124_, chained_data_delayed_93__123_, chained_data_delayed_93__122_, chained_data_delayed_93__121_, chained_data_delayed_93__120_, chained_data_delayed_93__119_, chained_data_delayed_93__118_, chained_data_delayed_93__117_, chained_data_delayed_93__116_, chained_data_delayed_93__115_, chained_data_delayed_93__114_, chained_data_delayed_93__113_, chained_data_delayed_93__112_, chained_data_delayed_93__111_, chained_data_delayed_93__110_, chained_data_delayed_93__109_, chained_data_delayed_93__108_, chained_data_delayed_93__107_, chained_data_delayed_93__106_, chained_data_delayed_93__105_, chained_data_delayed_93__104_, chained_data_delayed_93__103_, chained_data_delayed_93__102_, chained_data_delayed_93__101_, chained_data_delayed_93__100_, chained_data_delayed_93__99_, chained_data_delayed_93__98_, chained_data_delayed_93__97_, chained_data_delayed_93__96_, chained_data_delayed_93__95_, chained_data_delayed_93__94_, chained_data_delayed_93__93_, chained_data_delayed_93__92_, chained_data_delayed_93__91_, chained_data_delayed_93__90_, chained_data_delayed_93__89_, chained_data_delayed_93__88_, chained_data_delayed_93__87_, chained_data_delayed_93__86_, chained_data_delayed_93__85_, chained_data_delayed_93__84_, chained_data_delayed_93__83_, chained_data_delayed_93__82_, chained_data_delayed_93__81_, chained_data_delayed_93__80_, chained_data_delayed_93__79_, chained_data_delayed_93__78_, chained_data_delayed_93__77_, chained_data_delayed_93__76_, chained_data_delayed_93__75_, chained_data_delayed_93__74_, chained_data_delayed_93__73_, chained_data_delayed_93__72_, chained_data_delayed_93__71_, chained_data_delayed_93__70_, chained_data_delayed_93__69_, chained_data_delayed_93__68_, chained_data_delayed_93__67_, chained_data_delayed_93__66_, chained_data_delayed_93__65_, chained_data_delayed_93__64_, chained_data_delayed_93__63_, chained_data_delayed_93__62_, chained_data_delayed_93__61_, chained_data_delayed_93__60_, chained_data_delayed_93__59_, chained_data_delayed_93__58_, chained_data_delayed_93__57_, chained_data_delayed_93__56_, chained_data_delayed_93__55_, chained_data_delayed_93__54_, chained_data_delayed_93__53_, chained_data_delayed_93__52_, chained_data_delayed_93__51_, chained_data_delayed_93__50_, chained_data_delayed_93__49_, chained_data_delayed_93__48_, chained_data_delayed_93__47_, chained_data_delayed_93__46_, chained_data_delayed_93__45_, chained_data_delayed_93__44_, chained_data_delayed_93__43_, chained_data_delayed_93__42_, chained_data_delayed_93__41_, chained_data_delayed_93__40_, chained_data_delayed_93__39_, chained_data_delayed_93__38_, chained_data_delayed_93__37_, chained_data_delayed_93__36_, chained_data_delayed_93__35_, chained_data_delayed_93__34_, chained_data_delayed_93__33_, chained_data_delayed_93__32_, chained_data_delayed_93__31_, chained_data_delayed_93__30_, chained_data_delayed_93__29_, chained_data_delayed_93__28_, chained_data_delayed_93__27_, chained_data_delayed_93__26_, chained_data_delayed_93__25_, chained_data_delayed_93__24_, chained_data_delayed_93__23_, chained_data_delayed_93__22_, chained_data_delayed_93__21_, chained_data_delayed_93__20_, chained_data_delayed_93__19_, chained_data_delayed_93__18_, chained_data_delayed_93__17_, chained_data_delayed_93__16_, chained_data_delayed_93__15_, chained_data_delayed_93__14_, chained_data_delayed_93__13_, chained_data_delayed_93__12_, chained_data_delayed_93__11_, chained_data_delayed_93__10_, chained_data_delayed_93__9_, chained_data_delayed_93__8_, chained_data_delayed_93__7_, chained_data_delayed_93__6_, chained_data_delayed_93__5_, chained_data_delayed_93__4_, chained_data_delayed_93__3_, chained_data_delayed_93__2_, chained_data_delayed_93__1_, chained_data_delayed_93__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_94__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_93__127_, chained_data_delayed_93__126_, chained_data_delayed_93__125_, chained_data_delayed_93__124_, chained_data_delayed_93__123_, chained_data_delayed_93__122_, chained_data_delayed_93__121_, chained_data_delayed_93__120_, chained_data_delayed_93__119_, chained_data_delayed_93__118_, chained_data_delayed_93__117_, chained_data_delayed_93__116_, chained_data_delayed_93__115_, chained_data_delayed_93__114_, chained_data_delayed_93__113_, chained_data_delayed_93__112_, chained_data_delayed_93__111_, chained_data_delayed_93__110_, chained_data_delayed_93__109_, chained_data_delayed_93__108_, chained_data_delayed_93__107_, chained_data_delayed_93__106_, chained_data_delayed_93__105_, chained_data_delayed_93__104_, chained_data_delayed_93__103_, chained_data_delayed_93__102_, chained_data_delayed_93__101_, chained_data_delayed_93__100_, chained_data_delayed_93__99_, chained_data_delayed_93__98_, chained_data_delayed_93__97_, chained_data_delayed_93__96_, chained_data_delayed_93__95_, chained_data_delayed_93__94_, chained_data_delayed_93__93_, chained_data_delayed_93__92_, chained_data_delayed_93__91_, chained_data_delayed_93__90_, chained_data_delayed_93__89_, chained_data_delayed_93__88_, chained_data_delayed_93__87_, chained_data_delayed_93__86_, chained_data_delayed_93__85_, chained_data_delayed_93__84_, chained_data_delayed_93__83_, chained_data_delayed_93__82_, chained_data_delayed_93__81_, chained_data_delayed_93__80_, chained_data_delayed_93__79_, chained_data_delayed_93__78_, chained_data_delayed_93__77_, chained_data_delayed_93__76_, chained_data_delayed_93__75_, chained_data_delayed_93__74_, chained_data_delayed_93__73_, chained_data_delayed_93__72_, chained_data_delayed_93__71_, chained_data_delayed_93__70_, chained_data_delayed_93__69_, chained_data_delayed_93__68_, chained_data_delayed_93__67_, chained_data_delayed_93__66_, chained_data_delayed_93__65_, chained_data_delayed_93__64_, chained_data_delayed_93__63_, chained_data_delayed_93__62_, chained_data_delayed_93__61_, chained_data_delayed_93__60_, chained_data_delayed_93__59_, chained_data_delayed_93__58_, chained_data_delayed_93__57_, chained_data_delayed_93__56_, chained_data_delayed_93__55_, chained_data_delayed_93__54_, chained_data_delayed_93__53_, chained_data_delayed_93__52_, chained_data_delayed_93__51_, chained_data_delayed_93__50_, chained_data_delayed_93__49_, chained_data_delayed_93__48_, chained_data_delayed_93__47_, chained_data_delayed_93__46_, chained_data_delayed_93__45_, chained_data_delayed_93__44_, chained_data_delayed_93__43_, chained_data_delayed_93__42_, chained_data_delayed_93__41_, chained_data_delayed_93__40_, chained_data_delayed_93__39_, chained_data_delayed_93__38_, chained_data_delayed_93__37_, chained_data_delayed_93__36_, chained_data_delayed_93__35_, chained_data_delayed_93__34_, chained_data_delayed_93__33_, chained_data_delayed_93__32_, chained_data_delayed_93__31_, chained_data_delayed_93__30_, chained_data_delayed_93__29_, chained_data_delayed_93__28_, chained_data_delayed_93__27_, chained_data_delayed_93__26_, chained_data_delayed_93__25_, chained_data_delayed_93__24_, chained_data_delayed_93__23_, chained_data_delayed_93__22_, chained_data_delayed_93__21_, chained_data_delayed_93__20_, chained_data_delayed_93__19_, chained_data_delayed_93__18_, chained_data_delayed_93__17_, chained_data_delayed_93__16_, chained_data_delayed_93__15_, chained_data_delayed_93__14_, chained_data_delayed_93__13_, chained_data_delayed_93__12_, chained_data_delayed_93__11_, chained_data_delayed_93__10_, chained_data_delayed_93__9_, chained_data_delayed_93__8_, chained_data_delayed_93__7_, chained_data_delayed_93__6_, chained_data_delayed_93__5_, chained_data_delayed_93__4_, chained_data_delayed_93__3_, chained_data_delayed_93__2_, chained_data_delayed_93__1_, chained_data_delayed_93__0_ }),
    .data_o({ chained_data_delayed_94__127_, chained_data_delayed_94__126_, chained_data_delayed_94__125_, chained_data_delayed_94__124_, chained_data_delayed_94__123_, chained_data_delayed_94__122_, chained_data_delayed_94__121_, chained_data_delayed_94__120_, chained_data_delayed_94__119_, chained_data_delayed_94__118_, chained_data_delayed_94__117_, chained_data_delayed_94__116_, chained_data_delayed_94__115_, chained_data_delayed_94__114_, chained_data_delayed_94__113_, chained_data_delayed_94__112_, chained_data_delayed_94__111_, chained_data_delayed_94__110_, chained_data_delayed_94__109_, chained_data_delayed_94__108_, chained_data_delayed_94__107_, chained_data_delayed_94__106_, chained_data_delayed_94__105_, chained_data_delayed_94__104_, chained_data_delayed_94__103_, chained_data_delayed_94__102_, chained_data_delayed_94__101_, chained_data_delayed_94__100_, chained_data_delayed_94__99_, chained_data_delayed_94__98_, chained_data_delayed_94__97_, chained_data_delayed_94__96_, chained_data_delayed_94__95_, chained_data_delayed_94__94_, chained_data_delayed_94__93_, chained_data_delayed_94__92_, chained_data_delayed_94__91_, chained_data_delayed_94__90_, chained_data_delayed_94__89_, chained_data_delayed_94__88_, chained_data_delayed_94__87_, chained_data_delayed_94__86_, chained_data_delayed_94__85_, chained_data_delayed_94__84_, chained_data_delayed_94__83_, chained_data_delayed_94__82_, chained_data_delayed_94__81_, chained_data_delayed_94__80_, chained_data_delayed_94__79_, chained_data_delayed_94__78_, chained_data_delayed_94__77_, chained_data_delayed_94__76_, chained_data_delayed_94__75_, chained_data_delayed_94__74_, chained_data_delayed_94__73_, chained_data_delayed_94__72_, chained_data_delayed_94__71_, chained_data_delayed_94__70_, chained_data_delayed_94__69_, chained_data_delayed_94__68_, chained_data_delayed_94__67_, chained_data_delayed_94__66_, chained_data_delayed_94__65_, chained_data_delayed_94__64_, chained_data_delayed_94__63_, chained_data_delayed_94__62_, chained_data_delayed_94__61_, chained_data_delayed_94__60_, chained_data_delayed_94__59_, chained_data_delayed_94__58_, chained_data_delayed_94__57_, chained_data_delayed_94__56_, chained_data_delayed_94__55_, chained_data_delayed_94__54_, chained_data_delayed_94__53_, chained_data_delayed_94__52_, chained_data_delayed_94__51_, chained_data_delayed_94__50_, chained_data_delayed_94__49_, chained_data_delayed_94__48_, chained_data_delayed_94__47_, chained_data_delayed_94__46_, chained_data_delayed_94__45_, chained_data_delayed_94__44_, chained_data_delayed_94__43_, chained_data_delayed_94__42_, chained_data_delayed_94__41_, chained_data_delayed_94__40_, chained_data_delayed_94__39_, chained_data_delayed_94__38_, chained_data_delayed_94__37_, chained_data_delayed_94__36_, chained_data_delayed_94__35_, chained_data_delayed_94__34_, chained_data_delayed_94__33_, chained_data_delayed_94__32_, chained_data_delayed_94__31_, chained_data_delayed_94__30_, chained_data_delayed_94__29_, chained_data_delayed_94__28_, chained_data_delayed_94__27_, chained_data_delayed_94__26_, chained_data_delayed_94__25_, chained_data_delayed_94__24_, chained_data_delayed_94__23_, chained_data_delayed_94__22_, chained_data_delayed_94__21_, chained_data_delayed_94__20_, chained_data_delayed_94__19_, chained_data_delayed_94__18_, chained_data_delayed_94__17_, chained_data_delayed_94__16_, chained_data_delayed_94__15_, chained_data_delayed_94__14_, chained_data_delayed_94__13_, chained_data_delayed_94__12_, chained_data_delayed_94__11_, chained_data_delayed_94__10_, chained_data_delayed_94__9_, chained_data_delayed_94__8_, chained_data_delayed_94__7_, chained_data_delayed_94__6_, chained_data_delayed_94__5_, chained_data_delayed_94__4_, chained_data_delayed_94__3_, chained_data_delayed_94__2_, chained_data_delayed_94__1_, chained_data_delayed_94__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_95__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_94__127_, chained_data_delayed_94__126_, chained_data_delayed_94__125_, chained_data_delayed_94__124_, chained_data_delayed_94__123_, chained_data_delayed_94__122_, chained_data_delayed_94__121_, chained_data_delayed_94__120_, chained_data_delayed_94__119_, chained_data_delayed_94__118_, chained_data_delayed_94__117_, chained_data_delayed_94__116_, chained_data_delayed_94__115_, chained_data_delayed_94__114_, chained_data_delayed_94__113_, chained_data_delayed_94__112_, chained_data_delayed_94__111_, chained_data_delayed_94__110_, chained_data_delayed_94__109_, chained_data_delayed_94__108_, chained_data_delayed_94__107_, chained_data_delayed_94__106_, chained_data_delayed_94__105_, chained_data_delayed_94__104_, chained_data_delayed_94__103_, chained_data_delayed_94__102_, chained_data_delayed_94__101_, chained_data_delayed_94__100_, chained_data_delayed_94__99_, chained_data_delayed_94__98_, chained_data_delayed_94__97_, chained_data_delayed_94__96_, chained_data_delayed_94__95_, chained_data_delayed_94__94_, chained_data_delayed_94__93_, chained_data_delayed_94__92_, chained_data_delayed_94__91_, chained_data_delayed_94__90_, chained_data_delayed_94__89_, chained_data_delayed_94__88_, chained_data_delayed_94__87_, chained_data_delayed_94__86_, chained_data_delayed_94__85_, chained_data_delayed_94__84_, chained_data_delayed_94__83_, chained_data_delayed_94__82_, chained_data_delayed_94__81_, chained_data_delayed_94__80_, chained_data_delayed_94__79_, chained_data_delayed_94__78_, chained_data_delayed_94__77_, chained_data_delayed_94__76_, chained_data_delayed_94__75_, chained_data_delayed_94__74_, chained_data_delayed_94__73_, chained_data_delayed_94__72_, chained_data_delayed_94__71_, chained_data_delayed_94__70_, chained_data_delayed_94__69_, chained_data_delayed_94__68_, chained_data_delayed_94__67_, chained_data_delayed_94__66_, chained_data_delayed_94__65_, chained_data_delayed_94__64_, chained_data_delayed_94__63_, chained_data_delayed_94__62_, chained_data_delayed_94__61_, chained_data_delayed_94__60_, chained_data_delayed_94__59_, chained_data_delayed_94__58_, chained_data_delayed_94__57_, chained_data_delayed_94__56_, chained_data_delayed_94__55_, chained_data_delayed_94__54_, chained_data_delayed_94__53_, chained_data_delayed_94__52_, chained_data_delayed_94__51_, chained_data_delayed_94__50_, chained_data_delayed_94__49_, chained_data_delayed_94__48_, chained_data_delayed_94__47_, chained_data_delayed_94__46_, chained_data_delayed_94__45_, chained_data_delayed_94__44_, chained_data_delayed_94__43_, chained_data_delayed_94__42_, chained_data_delayed_94__41_, chained_data_delayed_94__40_, chained_data_delayed_94__39_, chained_data_delayed_94__38_, chained_data_delayed_94__37_, chained_data_delayed_94__36_, chained_data_delayed_94__35_, chained_data_delayed_94__34_, chained_data_delayed_94__33_, chained_data_delayed_94__32_, chained_data_delayed_94__31_, chained_data_delayed_94__30_, chained_data_delayed_94__29_, chained_data_delayed_94__28_, chained_data_delayed_94__27_, chained_data_delayed_94__26_, chained_data_delayed_94__25_, chained_data_delayed_94__24_, chained_data_delayed_94__23_, chained_data_delayed_94__22_, chained_data_delayed_94__21_, chained_data_delayed_94__20_, chained_data_delayed_94__19_, chained_data_delayed_94__18_, chained_data_delayed_94__17_, chained_data_delayed_94__16_, chained_data_delayed_94__15_, chained_data_delayed_94__14_, chained_data_delayed_94__13_, chained_data_delayed_94__12_, chained_data_delayed_94__11_, chained_data_delayed_94__10_, chained_data_delayed_94__9_, chained_data_delayed_94__8_, chained_data_delayed_94__7_, chained_data_delayed_94__6_, chained_data_delayed_94__5_, chained_data_delayed_94__4_, chained_data_delayed_94__3_, chained_data_delayed_94__2_, chained_data_delayed_94__1_, chained_data_delayed_94__0_ }),
    .data_o({ chained_data_delayed_95__127_, chained_data_delayed_95__126_, chained_data_delayed_95__125_, chained_data_delayed_95__124_, chained_data_delayed_95__123_, chained_data_delayed_95__122_, chained_data_delayed_95__121_, chained_data_delayed_95__120_, chained_data_delayed_95__119_, chained_data_delayed_95__118_, chained_data_delayed_95__117_, chained_data_delayed_95__116_, chained_data_delayed_95__115_, chained_data_delayed_95__114_, chained_data_delayed_95__113_, chained_data_delayed_95__112_, chained_data_delayed_95__111_, chained_data_delayed_95__110_, chained_data_delayed_95__109_, chained_data_delayed_95__108_, chained_data_delayed_95__107_, chained_data_delayed_95__106_, chained_data_delayed_95__105_, chained_data_delayed_95__104_, chained_data_delayed_95__103_, chained_data_delayed_95__102_, chained_data_delayed_95__101_, chained_data_delayed_95__100_, chained_data_delayed_95__99_, chained_data_delayed_95__98_, chained_data_delayed_95__97_, chained_data_delayed_95__96_, chained_data_delayed_95__95_, chained_data_delayed_95__94_, chained_data_delayed_95__93_, chained_data_delayed_95__92_, chained_data_delayed_95__91_, chained_data_delayed_95__90_, chained_data_delayed_95__89_, chained_data_delayed_95__88_, chained_data_delayed_95__87_, chained_data_delayed_95__86_, chained_data_delayed_95__85_, chained_data_delayed_95__84_, chained_data_delayed_95__83_, chained_data_delayed_95__82_, chained_data_delayed_95__81_, chained_data_delayed_95__80_, chained_data_delayed_95__79_, chained_data_delayed_95__78_, chained_data_delayed_95__77_, chained_data_delayed_95__76_, chained_data_delayed_95__75_, chained_data_delayed_95__74_, chained_data_delayed_95__73_, chained_data_delayed_95__72_, chained_data_delayed_95__71_, chained_data_delayed_95__70_, chained_data_delayed_95__69_, chained_data_delayed_95__68_, chained_data_delayed_95__67_, chained_data_delayed_95__66_, chained_data_delayed_95__65_, chained_data_delayed_95__64_, chained_data_delayed_95__63_, chained_data_delayed_95__62_, chained_data_delayed_95__61_, chained_data_delayed_95__60_, chained_data_delayed_95__59_, chained_data_delayed_95__58_, chained_data_delayed_95__57_, chained_data_delayed_95__56_, chained_data_delayed_95__55_, chained_data_delayed_95__54_, chained_data_delayed_95__53_, chained_data_delayed_95__52_, chained_data_delayed_95__51_, chained_data_delayed_95__50_, chained_data_delayed_95__49_, chained_data_delayed_95__48_, chained_data_delayed_95__47_, chained_data_delayed_95__46_, chained_data_delayed_95__45_, chained_data_delayed_95__44_, chained_data_delayed_95__43_, chained_data_delayed_95__42_, chained_data_delayed_95__41_, chained_data_delayed_95__40_, chained_data_delayed_95__39_, chained_data_delayed_95__38_, chained_data_delayed_95__37_, chained_data_delayed_95__36_, chained_data_delayed_95__35_, chained_data_delayed_95__34_, chained_data_delayed_95__33_, chained_data_delayed_95__32_, chained_data_delayed_95__31_, chained_data_delayed_95__30_, chained_data_delayed_95__29_, chained_data_delayed_95__28_, chained_data_delayed_95__27_, chained_data_delayed_95__26_, chained_data_delayed_95__25_, chained_data_delayed_95__24_, chained_data_delayed_95__23_, chained_data_delayed_95__22_, chained_data_delayed_95__21_, chained_data_delayed_95__20_, chained_data_delayed_95__19_, chained_data_delayed_95__18_, chained_data_delayed_95__17_, chained_data_delayed_95__16_, chained_data_delayed_95__15_, chained_data_delayed_95__14_, chained_data_delayed_95__13_, chained_data_delayed_95__12_, chained_data_delayed_95__11_, chained_data_delayed_95__10_, chained_data_delayed_95__9_, chained_data_delayed_95__8_, chained_data_delayed_95__7_, chained_data_delayed_95__6_, chained_data_delayed_95__5_, chained_data_delayed_95__4_, chained_data_delayed_95__3_, chained_data_delayed_95__2_, chained_data_delayed_95__1_, chained_data_delayed_95__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_96__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_95__127_, chained_data_delayed_95__126_, chained_data_delayed_95__125_, chained_data_delayed_95__124_, chained_data_delayed_95__123_, chained_data_delayed_95__122_, chained_data_delayed_95__121_, chained_data_delayed_95__120_, chained_data_delayed_95__119_, chained_data_delayed_95__118_, chained_data_delayed_95__117_, chained_data_delayed_95__116_, chained_data_delayed_95__115_, chained_data_delayed_95__114_, chained_data_delayed_95__113_, chained_data_delayed_95__112_, chained_data_delayed_95__111_, chained_data_delayed_95__110_, chained_data_delayed_95__109_, chained_data_delayed_95__108_, chained_data_delayed_95__107_, chained_data_delayed_95__106_, chained_data_delayed_95__105_, chained_data_delayed_95__104_, chained_data_delayed_95__103_, chained_data_delayed_95__102_, chained_data_delayed_95__101_, chained_data_delayed_95__100_, chained_data_delayed_95__99_, chained_data_delayed_95__98_, chained_data_delayed_95__97_, chained_data_delayed_95__96_, chained_data_delayed_95__95_, chained_data_delayed_95__94_, chained_data_delayed_95__93_, chained_data_delayed_95__92_, chained_data_delayed_95__91_, chained_data_delayed_95__90_, chained_data_delayed_95__89_, chained_data_delayed_95__88_, chained_data_delayed_95__87_, chained_data_delayed_95__86_, chained_data_delayed_95__85_, chained_data_delayed_95__84_, chained_data_delayed_95__83_, chained_data_delayed_95__82_, chained_data_delayed_95__81_, chained_data_delayed_95__80_, chained_data_delayed_95__79_, chained_data_delayed_95__78_, chained_data_delayed_95__77_, chained_data_delayed_95__76_, chained_data_delayed_95__75_, chained_data_delayed_95__74_, chained_data_delayed_95__73_, chained_data_delayed_95__72_, chained_data_delayed_95__71_, chained_data_delayed_95__70_, chained_data_delayed_95__69_, chained_data_delayed_95__68_, chained_data_delayed_95__67_, chained_data_delayed_95__66_, chained_data_delayed_95__65_, chained_data_delayed_95__64_, chained_data_delayed_95__63_, chained_data_delayed_95__62_, chained_data_delayed_95__61_, chained_data_delayed_95__60_, chained_data_delayed_95__59_, chained_data_delayed_95__58_, chained_data_delayed_95__57_, chained_data_delayed_95__56_, chained_data_delayed_95__55_, chained_data_delayed_95__54_, chained_data_delayed_95__53_, chained_data_delayed_95__52_, chained_data_delayed_95__51_, chained_data_delayed_95__50_, chained_data_delayed_95__49_, chained_data_delayed_95__48_, chained_data_delayed_95__47_, chained_data_delayed_95__46_, chained_data_delayed_95__45_, chained_data_delayed_95__44_, chained_data_delayed_95__43_, chained_data_delayed_95__42_, chained_data_delayed_95__41_, chained_data_delayed_95__40_, chained_data_delayed_95__39_, chained_data_delayed_95__38_, chained_data_delayed_95__37_, chained_data_delayed_95__36_, chained_data_delayed_95__35_, chained_data_delayed_95__34_, chained_data_delayed_95__33_, chained_data_delayed_95__32_, chained_data_delayed_95__31_, chained_data_delayed_95__30_, chained_data_delayed_95__29_, chained_data_delayed_95__28_, chained_data_delayed_95__27_, chained_data_delayed_95__26_, chained_data_delayed_95__25_, chained_data_delayed_95__24_, chained_data_delayed_95__23_, chained_data_delayed_95__22_, chained_data_delayed_95__21_, chained_data_delayed_95__20_, chained_data_delayed_95__19_, chained_data_delayed_95__18_, chained_data_delayed_95__17_, chained_data_delayed_95__16_, chained_data_delayed_95__15_, chained_data_delayed_95__14_, chained_data_delayed_95__13_, chained_data_delayed_95__12_, chained_data_delayed_95__11_, chained_data_delayed_95__10_, chained_data_delayed_95__9_, chained_data_delayed_95__8_, chained_data_delayed_95__7_, chained_data_delayed_95__6_, chained_data_delayed_95__5_, chained_data_delayed_95__4_, chained_data_delayed_95__3_, chained_data_delayed_95__2_, chained_data_delayed_95__1_, chained_data_delayed_95__0_ }),
    .data_o({ chained_data_delayed_96__127_, chained_data_delayed_96__126_, chained_data_delayed_96__125_, chained_data_delayed_96__124_, chained_data_delayed_96__123_, chained_data_delayed_96__122_, chained_data_delayed_96__121_, chained_data_delayed_96__120_, chained_data_delayed_96__119_, chained_data_delayed_96__118_, chained_data_delayed_96__117_, chained_data_delayed_96__116_, chained_data_delayed_96__115_, chained_data_delayed_96__114_, chained_data_delayed_96__113_, chained_data_delayed_96__112_, chained_data_delayed_96__111_, chained_data_delayed_96__110_, chained_data_delayed_96__109_, chained_data_delayed_96__108_, chained_data_delayed_96__107_, chained_data_delayed_96__106_, chained_data_delayed_96__105_, chained_data_delayed_96__104_, chained_data_delayed_96__103_, chained_data_delayed_96__102_, chained_data_delayed_96__101_, chained_data_delayed_96__100_, chained_data_delayed_96__99_, chained_data_delayed_96__98_, chained_data_delayed_96__97_, chained_data_delayed_96__96_, chained_data_delayed_96__95_, chained_data_delayed_96__94_, chained_data_delayed_96__93_, chained_data_delayed_96__92_, chained_data_delayed_96__91_, chained_data_delayed_96__90_, chained_data_delayed_96__89_, chained_data_delayed_96__88_, chained_data_delayed_96__87_, chained_data_delayed_96__86_, chained_data_delayed_96__85_, chained_data_delayed_96__84_, chained_data_delayed_96__83_, chained_data_delayed_96__82_, chained_data_delayed_96__81_, chained_data_delayed_96__80_, chained_data_delayed_96__79_, chained_data_delayed_96__78_, chained_data_delayed_96__77_, chained_data_delayed_96__76_, chained_data_delayed_96__75_, chained_data_delayed_96__74_, chained_data_delayed_96__73_, chained_data_delayed_96__72_, chained_data_delayed_96__71_, chained_data_delayed_96__70_, chained_data_delayed_96__69_, chained_data_delayed_96__68_, chained_data_delayed_96__67_, chained_data_delayed_96__66_, chained_data_delayed_96__65_, chained_data_delayed_96__64_, chained_data_delayed_96__63_, chained_data_delayed_96__62_, chained_data_delayed_96__61_, chained_data_delayed_96__60_, chained_data_delayed_96__59_, chained_data_delayed_96__58_, chained_data_delayed_96__57_, chained_data_delayed_96__56_, chained_data_delayed_96__55_, chained_data_delayed_96__54_, chained_data_delayed_96__53_, chained_data_delayed_96__52_, chained_data_delayed_96__51_, chained_data_delayed_96__50_, chained_data_delayed_96__49_, chained_data_delayed_96__48_, chained_data_delayed_96__47_, chained_data_delayed_96__46_, chained_data_delayed_96__45_, chained_data_delayed_96__44_, chained_data_delayed_96__43_, chained_data_delayed_96__42_, chained_data_delayed_96__41_, chained_data_delayed_96__40_, chained_data_delayed_96__39_, chained_data_delayed_96__38_, chained_data_delayed_96__37_, chained_data_delayed_96__36_, chained_data_delayed_96__35_, chained_data_delayed_96__34_, chained_data_delayed_96__33_, chained_data_delayed_96__32_, chained_data_delayed_96__31_, chained_data_delayed_96__30_, chained_data_delayed_96__29_, chained_data_delayed_96__28_, chained_data_delayed_96__27_, chained_data_delayed_96__26_, chained_data_delayed_96__25_, chained_data_delayed_96__24_, chained_data_delayed_96__23_, chained_data_delayed_96__22_, chained_data_delayed_96__21_, chained_data_delayed_96__20_, chained_data_delayed_96__19_, chained_data_delayed_96__18_, chained_data_delayed_96__17_, chained_data_delayed_96__16_, chained_data_delayed_96__15_, chained_data_delayed_96__14_, chained_data_delayed_96__13_, chained_data_delayed_96__12_, chained_data_delayed_96__11_, chained_data_delayed_96__10_, chained_data_delayed_96__9_, chained_data_delayed_96__8_, chained_data_delayed_96__7_, chained_data_delayed_96__6_, chained_data_delayed_96__5_, chained_data_delayed_96__4_, chained_data_delayed_96__3_, chained_data_delayed_96__2_, chained_data_delayed_96__1_, chained_data_delayed_96__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_97__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_96__127_, chained_data_delayed_96__126_, chained_data_delayed_96__125_, chained_data_delayed_96__124_, chained_data_delayed_96__123_, chained_data_delayed_96__122_, chained_data_delayed_96__121_, chained_data_delayed_96__120_, chained_data_delayed_96__119_, chained_data_delayed_96__118_, chained_data_delayed_96__117_, chained_data_delayed_96__116_, chained_data_delayed_96__115_, chained_data_delayed_96__114_, chained_data_delayed_96__113_, chained_data_delayed_96__112_, chained_data_delayed_96__111_, chained_data_delayed_96__110_, chained_data_delayed_96__109_, chained_data_delayed_96__108_, chained_data_delayed_96__107_, chained_data_delayed_96__106_, chained_data_delayed_96__105_, chained_data_delayed_96__104_, chained_data_delayed_96__103_, chained_data_delayed_96__102_, chained_data_delayed_96__101_, chained_data_delayed_96__100_, chained_data_delayed_96__99_, chained_data_delayed_96__98_, chained_data_delayed_96__97_, chained_data_delayed_96__96_, chained_data_delayed_96__95_, chained_data_delayed_96__94_, chained_data_delayed_96__93_, chained_data_delayed_96__92_, chained_data_delayed_96__91_, chained_data_delayed_96__90_, chained_data_delayed_96__89_, chained_data_delayed_96__88_, chained_data_delayed_96__87_, chained_data_delayed_96__86_, chained_data_delayed_96__85_, chained_data_delayed_96__84_, chained_data_delayed_96__83_, chained_data_delayed_96__82_, chained_data_delayed_96__81_, chained_data_delayed_96__80_, chained_data_delayed_96__79_, chained_data_delayed_96__78_, chained_data_delayed_96__77_, chained_data_delayed_96__76_, chained_data_delayed_96__75_, chained_data_delayed_96__74_, chained_data_delayed_96__73_, chained_data_delayed_96__72_, chained_data_delayed_96__71_, chained_data_delayed_96__70_, chained_data_delayed_96__69_, chained_data_delayed_96__68_, chained_data_delayed_96__67_, chained_data_delayed_96__66_, chained_data_delayed_96__65_, chained_data_delayed_96__64_, chained_data_delayed_96__63_, chained_data_delayed_96__62_, chained_data_delayed_96__61_, chained_data_delayed_96__60_, chained_data_delayed_96__59_, chained_data_delayed_96__58_, chained_data_delayed_96__57_, chained_data_delayed_96__56_, chained_data_delayed_96__55_, chained_data_delayed_96__54_, chained_data_delayed_96__53_, chained_data_delayed_96__52_, chained_data_delayed_96__51_, chained_data_delayed_96__50_, chained_data_delayed_96__49_, chained_data_delayed_96__48_, chained_data_delayed_96__47_, chained_data_delayed_96__46_, chained_data_delayed_96__45_, chained_data_delayed_96__44_, chained_data_delayed_96__43_, chained_data_delayed_96__42_, chained_data_delayed_96__41_, chained_data_delayed_96__40_, chained_data_delayed_96__39_, chained_data_delayed_96__38_, chained_data_delayed_96__37_, chained_data_delayed_96__36_, chained_data_delayed_96__35_, chained_data_delayed_96__34_, chained_data_delayed_96__33_, chained_data_delayed_96__32_, chained_data_delayed_96__31_, chained_data_delayed_96__30_, chained_data_delayed_96__29_, chained_data_delayed_96__28_, chained_data_delayed_96__27_, chained_data_delayed_96__26_, chained_data_delayed_96__25_, chained_data_delayed_96__24_, chained_data_delayed_96__23_, chained_data_delayed_96__22_, chained_data_delayed_96__21_, chained_data_delayed_96__20_, chained_data_delayed_96__19_, chained_data_delayed_96__18_, chained_data_delayed_96__17_, chained_data_delayed_96__16_, chained_data_delayed_96__15_, chained_data_delayed_96__14_, chained_data_delayed_96__13_, chained_data_delayed_96__12_, chained_data_delayed_96__11_, chained_data_delayed_96__10_, chained_data_delayed_96__9_, chained_data_delayed_96__8_, chained_data_delayed_96__7_, chained_data_delayed_96__6_, chained_data_delayed_96__5_, chained_data_delayed_96__4_, chained_data_delayed_96__3_, chained_data_delayed_96__2_, chained_data_delayed_96__1_, chained_data_delayed_96__0_ }),
    .data_o({ chained_data_delayed_97__127_, chained_data_delayed_97__126_, chained_data_delayed_97__125_, chained_data_delayed_97__124_, chained_data_delayed_97__123_, chained_data_delayed_97__122_, chained_data_delayed_97__121_, chained_data_delayed_97__120_, chained_data_delayed_97__119_, chained_data_delayed_97__118_, chained_data_delayed_97__117_, chained_data_delayed_97__116_, chained_data_delayed_97__115_, chained_data_delayed_97__114_, chained_data_delayed_97__113_, chained_data_delayed_97__112_, chained_data_delayed_97__111_, chained_data_delayed_97__110_, chained_data_delayed_97__109_, chained_data_delayed_97__108_, chained_data_delayed_97__107_, chained_data_delayed_97__106_, chained_data_delayed_97__105_, chained_data_delayed_97__104_, chained_data_delayed_97__103_, chained_data_delayed_97__102_, chained_data_delayed_97__101_, chained_data_delayed_97__100_, chained_data_delayed_97__99_, chained_data_delayed_97__98_, chained_data_delayed_97__97_, chained_data_delayed_97__96_, chained_data_delayed_97__95_, chained_data_delayed_97__94_, chained_data_delayed_97__93_, chained_data_delayed_97__92_, chained_data_delayed_97__91_, chained_data_delayed_97__90_, chained_data_delayed_97__89_, chained_data_delayed_97__88_, chained_data_delayed_97__87_, chained_data_delayed_97__86_, chained_data_delayed_97__85_, chained_data_delayed_97__84_, chained_data_delayed_97__83_, chained_data_delayed_97__82_, chained_data_delayed_97__81_, chained_data_delayed_97__80_, chained_data_delayed_97__79_, chained_data_delayed_97__78_, chained_data_delayed_97__77_, chained_data_delayed_97__76_, chained_data_delayed_97__75_, chained_data_delayed_97__74_, chained_data_delayed_97__73_, chained_data_delayed_97__72_, chained_data_delayed_97__71_, chained_data_delayed_97__70_, chained_data_delayed_97__69_, chained_data_delayed_97__68_, chained_data_delayed_97__67_, chained_data_delayed_97__66_, chained_data_delayed_97__65_, chained_data_delayed_97__64_, chained_data_delayed_97__63_, chained_data_delayed_97__62_, chained_data_delayed_97__61_, chained_data_delayed_97__60_, chained_data_delayed_97__59_, chained_data_delayed_97__58_, chained_data_delayed_97__57_, chained_data_delayed_97__56_, chained_data_delayed_97__55_, chained_data_delayed_97__54_, chained_data_delayed_97__53_, chained_data_delayed_97__52_, chained_data_delayed_97__51_, chained_data_delayed_97__50_, chained_data_delayed_97__49_, chained_data_delayed_97__48_, chained_data_delayed_97__47_, chained_data_delayed_97__46_, chained_data_delayed_97__45_, chained_data_delayed_97__44_, chained_data_delayed_97__43_, chained_data_delayed_97__42_, chained_data_delayed_97__41_, chained_data_delayed_97__40_, chained_data_delayed_97__39_, chained_data_delayed_97__38_, chained_data_delayed_97__37_, chained_data_delayed_97__36_, chained_data_delayed_97__35_, chained_data_delayed_97__34_, chained_data_delayed_97__33_, chained_data_delayed_97__32_, chained_data_delayed_97__31_, chained_data_delayed_97__30_, chained_data_delayed_97__29_, chained_data_delayed_97__28_, chained_data_delayed_97__27_, chained_data_delayed_97__26_, chained_data_delayed_97__25_, chained_data_delayed_97__24_, chained_data_delayed_97__23_, chained_data_delayed_97__22_, chained_data_delayed_97__21_, chained_data_delayed_97__20_, chained_data_delayed_97__19_, chained_data_delayed_97__18_, chained_data_delayed_97__17_, chained_data_delayed_97__16_, chained_data_delayed_97__15_, chained_data_delayed_97__14_, chained_data_delayed_97__13_, chained_data_delayed_97__12_, chained_data_delayed_97__11_, chained_data_delayed_97__10_, chained_data_delayed_97__9_, chained_data_delayed_97__8_, chained_data_delayed_97__7_, chained_data_delayed_97__6_, chained_data_delayed_97__5_, chained_data_delayed_97__4_, chained_data_delayed_97__3_, chained_data_delayed_97__2_, chained_data_delayed_97__1_, chained_data_delayed_97__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_98__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_97__127_, chained_data_delayed_97__126_, chained_data_delayed_97__125_, chained_data_delayed_97__124_, chained_data_delayed_97__123_, chained_data_delayed_97__122_, chained_data_delayed_97__121_, chained_data_delayed_97__120_, chained_data_delayed_97__119_, chained_data_delayed_97__118_, chained_data_delayed_97__117_, chained_data_delayed_97__116_, chained_data_delayed_97__115_, chained_data_delayed_97__114_, chained_data_delayed_97__113_, chained_data_delayed_97__112_, chained_data_delayed_97__111_, chained_data_delayed_97__110_, chained_data_delayed_97__109_, chained_data_delayed_97__108_, chained_data_delayed_97__107_, chained_data_delayed_97__106_, chained_data_delayed_97__105_, chained_data_delayed_97__104_, chained_data_delayed_97__103_, chained_data_delayed_97__102_, chained_data_delayed_97__101_, chained_data_delayed_97__100_, chained_data_delayed_97__99_, chained_data_delayed_97__98_, chained_data_delayed_97__97_, chained_data_delayed_97__96_, chained_data_delayed_97__95_, chained_data_delayed_97__94_, chained_data_delayed_97__93_, chained_data_delayed_97__92_, chained_data_delayed_97__91_, chained_data_delayed_97__90_, chained_data_delayed_97__89_, chained_data_delayed_97__88_, chained_data_delayed_97__87_, chained_data_delayed_97__86_, chained_data_delayed_97__85_, chained_data_delayed_97__84_, chained_data_delayed_97__83_, chained_data_delayed_97__82_, chained_data_delayed_97__81_, chained_data_delayed_97__80_, chained_data_delayed_97__79_, chained_data_delayed_97__78_, chained_data_delayed_97__77_, chained_data_delayed_97__76_, chained_data_delayed_97__75_, chained_data_delayed_97__74_, chained_data_delayed_97__73_, chained_data_delayed_97__72_, chained_data_delayed_97__71_, chained_data_delayed_97__70_, chained_data_delayed_97__69_, chained_data_delayed_97__68_, chained_data_delayed_97__67_, chained_data_delayed_97__66_, chained_data_delayed_97__65_, chained_data_delayed_97__64_, chained_data_delayed_97__63_, chained_data_delayed_97__62_, chained_data_delayed_97__61_, chained_data_delayed_97__60_, chained_data_delayed_97__59_, chained_data_delayed_97__58_, chained_data_delayed_97__57_, chained_data_delayed_97__56_, chained_data_delayed_97__55_, chained_data_delayed_97__54_, chained_data_delayed_97__53_, chained_data_delayed_97__52_, chained_data_delayed_97__51_, chained_data_delayed_97__50_, chained_data_delayed_97__49_, chained_data_delayed_97__48_, chained_data_delayed_97__47_, chained_data_delayed_97__46_, chained_data_delayed_97__45_, chained_data_delayed_97__44_, chained_data_delayed_97__43_, chained_data_delayed_97__42_, chained_data_delayed_97__41_, chained_data_delayed_97__40_, chained_data_delayed_97__39_, chained_data_delayed_97__38_, chained_data_delayed_97__37_, chained_data_delayed_97__36_, chained_data_delayed_97__35_, chained_data_delayed_97__34_, chained_data_delayed_97__33_, chained_data_delayed_97__32_, chained_data_delayed_97__31_, chained_data_delayed_97__30_, chained_data_delayed_97__29_, chained_data_delayed_97__28_, chained_data_delayed_97__27_, chained_data_delayed_97__26_, chained_data_delayed_97__25_, chained_data_delayed_97__24_, chained_data_delayed_97__23_, chained_data_delayed_97__22_, chained_data_delayed_97__21_, chained_data_delayed_97__20_, chained_data_delayed_97__19_, chained_data_delayed_97__18_, chained_data_delayed_97__17_, chained_data_delayed_97__16_, chained_data_delayed_97__15_, chained_data_delayed_97__14_, chained_data_delayed_97__13_, chained_data_delayed_97__12_, chained_data_delayed_97__11_, chained_data_delayed_97__10_, chained_data_delayed_97__9_, chained_data_delayed_97__8_, chained_data_delayed_97__7_, chained_data_delayed_97__6_, chained_data_delayed_97__5_, chained_data_delayed_97__4_, chained_data_delayed_97__3_, chained_data_delayed_97__2_, chained_data_delayed_97__1_, chained_data_delayed_97__0_ }),
    .data_o({ chained_data_delayed_98__127_, chained_data_delayed_98__126_, chained_data_delayed_98__125_, chained_data_delayed_98__124_, chained_data_delayed_98__123_, chained_data_delayed_98__122_, chained_data_delayed_98__121_, chained_data_delayed_98__120_, chained_data_delayed_98__119_, chained_data_delayed_98__118_, chained_data_delayed_98__117_, chained_data_delayed_98__116_, chained_data_delayed_98__115_, chained_data_delayed_98__114_, chained_data_delayed_98__113_, chained_data_delayed_98__112_, chained_data_delayed_98__111_, chained_data_delayed_98__110_, chained_data_delayed_98__109_, chained_data_delayed_98__108_, chained_data_delayed_98__107_, chained_data_delayed_98__106_, chained_data_delayed_98__105_, chained_data_delayed_98__104_, chained_data_delayed_98__103_, chained_data_delayed_98__102_, chained_data_delayed_98__101_, chained_data_delayed_98__100_, chained_data_delayed_98__99_, chained_data_delayed_98__98_, chained_data_delayed_98__97_, chained_data_delayed_98__96_, chained_data_delayed_98__95_, chained_data_delayed_98__94_, chained_data_delayed_98__93_, chained_data_delayed_98__92_, chained_data_delayed_98__91_, chained_data_delayed_98__90_, chained_data_delayed_98__89_, chained_data_delayed_98__88_, chained_data_delayed_98__87_, chained_data_delayed_98__86_, chained_data_delayed_98__85_, chained_data_delayed_98__84_, chained_data_delayed_98__83_, chained_data_delayed_98__82_, chained_data_delayed_98__81_, chained_data_delayed_98__80_, chained_data_delayed_98__79_, chained_data_delayed_98__78_, chained_data_delayed_98__77_, chained_data_delayed_98__76_, chained_data_delayed_98__75_, chained_data_delayed_98__74_, chained_data_delayed_98__73_, chained_data_delayed_98__72_, chained_data_delayed_98__71_, chained_data_delayed_98__70_, chained_data_delayed_98__69_, chained_data_delayed_98__68_, chained_data_delayed_98__67_, chained_data_delayed_98__66_, chained_data_delayed_98__65_, chained_data_delayed_98__64_, chained_data_delayed_98__63_, chained_data_delayed_98__62_, chained_data_delayed_98__61_, chained_data_delayed_98__60_, chained_data_delayed_98__59_, chained_data_delayed_98__58_, chained_data_delayed_98__57_, chained_data_delayed_98__56_, chained_data_delayed_98__55_, chained_data_delayed_98__54_, chained_data_delayed_98__53_, chained_data_delayed_98__52_, chained_data_delayed_98__51_, chained_data_delayed_98__50_, chained_data_delayed_98__49_, chained_data_delayed_98__48_, chained_data_delayed_98__47_, chained_data_delayed_98__46_, chained_data_delayed_98__45_, chained_data_delayed_98__44_, chained_data_delayed_98__43_, chained_data_delayed_98__42_, chained_data_delayed_98__41_, chained_data_delayed_98__40_, chained_data_delayed_98__39_, chained_data_delayed_98__38_, chained_data_delayed_98__37_, chained_data_delayed_98__36_, chained_data_delayed_98__35_, chained_data_delayed_98__34_, chained_data_delayed_98__33_, chained_data_delayed_98__32_, chained_data_delayed_98__31_, chained_data_delayed_98__30_, chained_data_delayed_98__29_, chained_data_delayed_98__28_, chained_data_delayed_98__27_, chained_data_delayed_98__26_, chained_data_delayed_98__25_, chained_data_delayed_98__24_, chained_data_delayed_98__23_, chained_data_delayed_98__22_, chained_data_delayed_98__21_, chained_data_delayed_98__20_, chained_data_delayed_98__19_, chained_data_delayed_98__18_, chained_data_delayed_98__17_, chained_data_delayed_98__16_, chained_data_delayed_98__15_, chained_data_delayed_98__14_, chained_data_delayed_98__13_, chained_data_delayed_98__12_, chained_data_delayed_98__11_, chained_data_delayed_98__10_, chained_data_delayed_98__9_, chained_data_delayed_98__8_, chained_data_delayed_98__7_, chained_data_delayed_98__6_, chained_data_delayed_98__5_, chained_data_delayed_98__4_, chained_data_delayed_98__3_, chained_data_delayed_98__2_, chained_data_delayed_98__1_, chained_data_delayed_98__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_99__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_98__127_, chained_data_delayed_98__126_, chained_data_delayed_98__125_, chained_data_delayed_98__124_, chained_data_delayed_98__123_, chained_data_delayed_98__122_, chained_data_delayed_98__121_, chained_data_delayed_98__120_, chained_data_delayed_98__119_, chained_data_delayed_98__118_, chained_data_delayed_98__117_, chained_data_delayed_98__116_, chained_data_delayed_98__115_, chained_data_delayed_98__114_, chained_data_delayed_98__113_, chained_data_delayed_98__112_, chained_data_delayed_98__111_, chained_data_delayed_98__110_, chained_data_delayed_98__109_, chained_data_delayed_98__108_, chained_data_delayed_98__107_, chained_data_delayed_98__106_, chained_data_delayed_98__105_, chained_data_delayed_98__104_, chained_data_delayed_98__103_, chained_data_delayed_98__102_, chained_data_delayed_98__101_, chained_data_delayed_98__100_, chained_data_delayed_98__99_, chained_data_delayed_98__98_, chained_data_delayed_98__97_, chained_data_delayed_98__96_, chained_data_delayed_98__95_, chained_data_delayed_98__94_, chained_data_delayed_98__93_, chained_data_delayed_98__92_, chained_data_delayed_98__91_, chained_data_delayed_98__90_, chained_data_delayed_98__89_, chained_data_delayed_98__88_, chained_data_delayed_98__87_, chained_data_delayed_98__86_, chained_data_delayed_98__85_, chained_data_delayed_98__84_, chained_data_delayed_98__83_, chained_data_delayed_98__82_, chained_data_delayed_98__81_, chained_data_delayed_98__80_, chained_data_delayed_98__79_, chained_data_delayed_98__78_, chained_data_delayed_98__77_, chained_data_delayed_98__76_, chained_data_delayed_98__75_, chained_data_delayed_98__74_, chained_data_delayed_98__73_, chained_data_delayed_98__72_, chained_data_delayed_98__71_, chained_data_delayed_98__70_, chained_data_delayed_98__69_, chained_data_delayed_98__68_, chained_data_delayed_98__67_, chained_data_delayed_98__66_, chained_data_delayed_98__65_, chained_data_delayed_98__64_, chained_data_delayed_98__63_, chained_data_delayed_98__62_, chained_data_delayed_98__61_, chained_data_delayed_98__60_, chained_data_delayed_98__59_, chained_data_delayed_98__58_, chained_data_delayed_98__57_, chained_data_delayed_98__56_, chained_data_delayed_98__55_, chained_data_delayed_98__54_, chained_data_delayed_98__53_, chained_data_delayed_98__52_, chained_data_delayed_98__51_, chained_data_delayed_98__50_, chained_data_delayed_98__49_, chained_data_delayed_98__48_, chained_data_delayed_98__47_, chained_data_delayed_98__46_, chained_data_delayed_98__45_, chained_data_delayed_98__44_, chained_data_delayed_98__43_, chained_data_delayed_98__42_, chained_data_delayed_98__41_, chained_data_delayed_98__40_, chained_data_delayed_98__39_, chained_data_delayed_98__38_, chained_data_delayed_98__37_, chained_data_delayed_98__36_, chained_data_delayed_98__35_, chained_data_delayed_98__34_, chained_data_delayed_98__33_, chained_data_delayed_98__32_, chained_data_delayed_98__31_, chained_data_delayed_98__30_, chained_data_delayed_98__29_, chained_data_delayed_98__28_, chained_data_delayed_98__27_, chained_data_delayed_98__26_, chained_data_delayed_98__25_, chained_data_delayed_98__24_, chained_data_delayed_98__23_, chained_data_delayed_98__22_, chained_data_delayed_98__21_, chained_data_delayed_98__20_, chained_data_delayed_98__19_, chained_data_delayed_98__18_, chained_data_delayed_98__17_, chained_data_delayed_98__16_, chained_data_delayed_98__15_, chained_data_delayed_98__14_, chained_data_delayed_98__13_, chained_data_delayed_98__12_, chained_data_delayed_98__11_, chained_data_delayed_98__10_, chained_data_delayed_98__9_, chained_data_delayed_98__8_, chained_data_delayed_98__7_, chained_data_delayed_98__6_, chained_data_delayed_98__5_, chained_data_delayed_98__4_, chained_data_delayed_98__3_, chained_data_delayed_98__2_, chained_data_delayed_98__1_, chained_data_delayed_98__0_ }),
    .data_o({ chained_data_delayed_99__127_, chained_data_delayed_99__126_, chained_data_delayed_99__125_, chained_data_delayed_99__124_, chained_data_delayed_99__123_, chained_data_delayed_99__122_, chained_data_delayed_99__121_, chained_data_delayed_99__120_, chained_data_delayed_99__119_, chained_data_delayed_99__118_, chained_data_delayed_99__117_, chained_data_delayed_99__116_, chained_data_delayed_99__115_, chained_data_delayed_99__114_, chained_data_delayed_99__113_, chained_data_delayed_99__112_, chained_data_delayed_99__111_, chained_data_delayed_99__110_, chained_data_delayed_99__109_, chained_data_delayed_99__108_, chained_data_delayed_99__107_, chained_data_delayed_99__106_, chained_data_delayed_99__105_, chained_data_delayed_99__104_, chained_data_delayed_99__103_, chained_data_delayed_99__102_, chained_data_delayed_99__101_, chained_data_delayed_99__100_, chained_data_delayed_99__99_, chained_data_delayed_99__98_, chained_data_delayed_99__97_, chained_data_delayed_99__96_, chained_data_delayed_99__95_, chained_data_delayed_99__94_, chained_data_delayed_99__93_, chained_data_delayed_99__92_, chained_data_delayed_99__91_, chained_data_delayed_99__90_, chained_data_delayed_99__89_, chained_data_delayed_99__88_, chained_data_delayed_99__87_, chained_data_delayed_99__86_, chained_data_delayed_99__85_, chained_data_delayed_99__84_, chained_data_delayed_99__83_, chained_data_delayed_99__82_, chained_data_delayed_99__81_, chained_data_delayed_99__80_, chained_data_delayed_99__79_, chained_data_delayed_99__78_, chained_data_delayed_99__77_, chained_data_delayed_99__76_, chained_data_delayed_99__75_, chained_data_delayed_99__74_, chained_data_delayed_99__73_, chained_data_delayed_99__72_, chained_data_delayed_99__71_, chained_data_delayed_99__70_, chained_data_delayed_99__69_, chained_data_delayed_99__68_, chained_data_delayed_99__67_, chained_data_delayed_99__66_, chained_data_delayed_99__65_, chained_data_delayed_99__64_, chained_data_delayed_99__63_, chained_data_delayed_99__62_, chained_data_delayed_99__61_, chained_data_delayed_99__60_, chained_data_delayed_99__59_, chained_data_delayed_99__58_, chained_data_delayed_99__57_, chained_data_delayed_99__56_, chained_data_delayed_99__55_, chained_data_delayed_99__54_, chained_data_delayed_99__53_, chained_data_delayed_99__52_, chained_data_delayed_99__51_, chained_data_delayed_99__50_, chained_data_delayed_99__49_, chained_data_delayed_99__48_, chained_data_delayed_99__47_, chained_data_delayed_99__46_, chained_data_delayed_99__45_, chained_data_delayed_99__44_, chained_data_delayed_99__43_, chained_data_delayed_99__42_, chained_data_delayed_99__41_, chained_data_delayed_99__40_, chained_data_delayed_99__39_, chained_data_delayed_99__38_, chained_data_delayed_99__37_, chained_data_delayed_99__36_, chained_data_delayed_99__35_, chained_data_delayed_99__34_, chained_data_delayed_99__33_, chained_data_delayed_99__32_, chained_data_delayed_99__31_, chained_data_delayed_99__30_, chained_data_delayed_99__29_, chained_data_delayed_99__28_, chained_data_delayed_99__27_, chained_data_delayed_99__26_, chained_data_delayed_99__25_, chained_data_delayed_99__24_, chained_data_delayed_99__23_, chained_data_delayed_99__22_, chained_data_delayed_99__21_, chained_data_delayed_99__20_, chained_data_delayed_99__19_, chained_data_delayed_99__18_, chained_data_delayed_99__17_, chained_data_delayed_99__16_, chained_data_delayed_99__15_, chained_data_delayed_99__14_, chained_data_delayed_99__13_, chained_data_delayed_99__12_, chained_data_delayed_99__11_, chained_data_delayed_99__10_, chained_data_delayed_99__9_, chained_data_delayed_99__8_, chained_data_delayed_99__7_, chained_data_delayed_99__6_, chained_data_delayed_99__5_, chained_data_delayed_99__4_, chained_data_delayed_99__3_, chained_data_delayed_99__2_, chained_data_delayed_99__1_, chained_data_delayed_99__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_100__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_99__127_, chained_data_delayed_99__126_, chained_data_delayed_99__125_, chained_data_delayed_99__124_, chained_data_delayed_99__123_, chained_data_delayed_99__122_, chained_data_delayed_99__121_, chained_data_delayed_99__120_, chained_data_delayed_99__119_, chained_data_delayed_99__118_, chained_data_delayed_99__117_, chained_data_delayed_99__116_, chained_data_delayed_99__115_, chained_data_delayed_99__114_, chained_data_delayed_99__113_, chained_data_delayed_99__112_, chained_data_delayed_99__111_, chained_data_delayed_99__110_, chained_data_delayed_99__109_, chained_data_delayed_99__108_, chained_data_delayed_99__107_, chained_data_delayed_99__106_, chained_data_delayed_99__105_, chained_data_delayed_99__104_, chained_data_delayed_99__103_, chained_data_delayed_99__102_, chained_data_delayed_99__101_, chained_data_delayed_99__100_, chained_data_delayed_99__99_, chained_data_delayed_99__98_, chained_data_delayed_99__97_, chained_data_delayed_99__96_, chained_data_delayed_99__95_, chained_data_delayed_99__94_, chained_data_delayed_99__93_, chained_data_delayed_99__92_, chained_data_delayed_99__91_, chained_data_delayed_99__90_, chained_data_delayed_99__89_, chained_data_delayed_99__88_, chained_data_delayed_99__87_, chained_data_delayed_99__86_, chained_data_delayed_99__85_, chained_data_delayed_99__84_, chained_data_delayed_99__83_, chained_data_delayed_99__82_, chained_data_delayed_99__81_, chained_data_delayed_99__80_, chained_data_delayed_99__79_, chained_data_delayed_99__78_, chained_data_delayed_99__77_, chained_data_delayed_99__76_, chained_data_delayed_99__75_, chained_data_delayed_99__74_, chained_data_delayed_99__73_, chained_data_delayed_99__72_, chained_data_delayed_99__71_, chained_data_delayed_99__70_, chained_data_delayed_99__69_, chained_data_delayed_99__68_, chained_data_delayed_99__67_, chained_data_delayed_99__66_, chained_data_delayed_99__65_, chained_data_delayed_99__64_, chained_data_delayed_99__63_, chained_data_delayed_99__62_, chained_data_delayed_99__61_, chained_data_delayed_99__60_, chained_data_delayed_99__59_, chained_data_delayed_99__58_, chained_data_delayed_99__57_, chained_data_delayed_99__56_, chained_data_delayed_99__55_, chained_data_delayed_99__54_, chained_data_delayed_99__53_, chained_data_delayed_99__52_, chained_data_delayed_99__51_, chained_data_delayed_99__50_, chained_data_delayed_99__49_, chained_data_delayed_99__48_, chained_data_delayed_99__47_, chained_data_delayed_99__46_, chained_data_delayed_99__45_, chained_data_delayed_99__44_, chained_data_delayed_99__43_, chained_data_delayed_99__42_, chained_data_delayed_99__41_, chained_data_delayed_99__40_, chained_data_delayed_99__39_, chained_data_delayed_99__38_, chained_data_delayed_99__37_, chained_data_delayed_99__36_, chained_data_delayed_99__35_, chained_data_delayed_99__34_, chained_data_delayed_99__33_, chained_data_delayed_99__32_, chained_data_delayed_99__31_, chained_data_delayed_99__30_, chained_data_delayed_99__29_, chained_data_delayed_99__28_, chained_data_delayed_99__27_, chained_data_delayed_99__26_, chained_data_delayed_99__25_, chained_data_delayed_99__24_, chained_data_delayed_99__23_, chained_data_delayed_99__22_, chained_data_delayed_99__21_, chained_data_delayed_99__20_, chained_data_delayed_99__19_, chained_data_delayed_99__18_, chained_data_delayed_99__17_, chained_data_delayed_99__16_, chained_data_delayed_99__15_, chained_data_delayed_99__14_, chained_data_delayed_99__13_, chained_data_delayed_99__12_, chained_data_delayed_99__11_, chained_data_delayed_99__10_, chained_data_delayed_99__9_, chained_data_delayed_99__8_, chained_data_delayed_99__7_, chained_data_delayed_99__6_, chained_data_delayed_99__5_, chained_data_delayed_99__4_, chained_data_delayed_99__3_, chained_data_delayed_99__2_, chained_data_delayed_99__1_, chained_data_delayed_99__0_ }),
    .data_o({ chained_data_delayed_100__127_, chained_data_delayed_100__126_, chained_data_delayed_100__125_, chained_data_delayed_100__124_, chained_data_delayed_100__123_, chained_data_delayed_100__122_, chained_data_delayed_100__121_, chained_data_delayed_100__120_, chained_data_delayed_100__119_, chained_data_delayed_100__118_, chained_data_delayed_100__117_, chained_data_delayed_100__116_, chained_data_delayed_100__115_, chained_data_delayed_100__114_, chained_data_delayed_100__113_, chained_data_delayed_100__112_, chained_data_delayed_100__111_, chained_data_delayed_100__110_, chained_data_delayed_100__109_, chained_data_delayed_100__108_, chained_data_delayed_100__107_, chained_data_delayed_100__106_, chained_data_delayed_100__105_, chained_data_delayed_100__104_, chained_data_delayed_100__103_, chained_data_delayed_100__102_, chained_data_delayed_100__101_, chained_data_delayed_100__100_, chained_data_delayed_100__99_, chained_data_delayed_100__98_, chained_data_delayed_100__97_, chained_data_delayed_100__96_, chained_data_delayed_100__95_, chained_data_delayed_100__94_, chained_data_delayed_100__93_, chained_data_delayed_100__92_, chained_data_delayed_100__91_, chained_data_delayed_100__90_, chained_data_delayed_100__89_, chained_data_delayed_100__88_, chained_data_delayed_100__87_, chained_data_delayed_100__86_, chained_data_delayed_100__85_, chained_data_delayed_100__84_, chained_data_delayed_100__83_, chained_data_delayed_100__82_, chained_data_delayed_100__81_, chained_data_delayed_100__80_, chained_data_delayed_100__79_, chained_data_delayed_100__78_, chained_data_delayed_100__77_, chained_data_delayed_100__76_, chained_data_delayed_100__75_, chained_data_delayed_100__74_, chained_data_delayed_100__73_, chained_data_delayed_100__72_, chained_data_delayed_100__71_, chained_data_delayed_100__70_, chained_data_delayed_100__69_, chained_data_delayed_100__68_, chained_data_delayed_100__67_, chained_data_delayed_100__66_, chained_data_delayed_100__65_, chained_data_delayed_100__64_, chained_data_delayed_100__63_, chained_data_delayed_100__62_, chained_data_delayed_100__61_, chained_data_delayed_100__60_, chained_data_delayed_100__59_, chained_data_delayed_100__58_, chained_data_delayed_100__57_, chained_data_delayed_100__56_, chained_data_delayed_100__55_, chained_data_delayed_100__54_, chained_data_delayed_100__53_, chained_data_delayed_100__52_, chained_data_delayed_100__51_, chained_data_delayed_100__50_, chained_data_delayed_100__49_, chained_data_delayed_100__48_, chained_data_delayed_100__47_, chained_data_delayed_100__46_, chained_data_delayed_100__45_, chained_data_delayed_100__44_, chained_data_delayed_100__43_, chained_data_delayed_100__42_, chained_data_delayed_100__41_, chained_data_delayed_100__40_, chained_data_delayed_100__39_, chained_data_delayed_100__38_, chained_data_delayed_100__37_, chained_data_delayed_100__36_, chained_data_delayed_100__35_, chained_data_delayed_100__34_, chained_data_delayed_100__33_, chained_data_delayed_100__32_, chained_data_delayed_100__31_, chained_data_delayed_100__30_, chained_data_delayed_100__29_, chained_data_delayed_100__28_, chained_data_delayed_100__27_, chained_data_delayed_100__26_, chained_data_delayed_100__25_, chained_data_delayed_100__24_, chained_data_delayed_100__23_, chained_data_delayed_100__22_, chained_data_delayed_100__21_, chained_data_delayed_100__20_, chained_data_delayed_100__19_, chained_data_delayed_100__18_, chained_data_delayed_100__17_, chained_data_delayed_100__16_, chained_data_delayed_100__15_, chained_data_delayed_100__14_, chained_data_delayed_100__13_, chained_data_delayed_100__12_, chained_data_delayed_100__11_, chained_data_delayed_100__10_, chained_data_delayed_100__9_, chained_data_delayed_100__8_, chained_data_delayed_100__7_, chained_data_delayed_100__6_, chained_data_delayed_100__5_, chained_data_delayed_100__4_, chained_data_delayed_100__3_, chained_data_delayed_100__2_, chained_data_delayed_100__1_, chained_data_delayed_100__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_101__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_100__127_, chained_data_delayed_100__126_, chained_data_delayed_100__125_, chained_data_delayed_100__124_, chained_data_delayed_100__123_, chained_data_delayed_100__122_, chained_data_delayed_100__121_, chained_data_delayed_100__120_, chained_data_delayed_100__119_, chained_data_delayed_100__118_, chained_data_delayed_100__117_, chained_data_delayed_100__116_, chained_data_delayed_100__115_, chained_data_delayed_100__114_, chained_data_delayed_100__113_, chained_data_delayed_100__112_, chained_data_delayed_100__111_, chained_data_delayed_100__110_, chained_data_delayed_100__109_, chained_data_delayed_100__108_, chained_data_delayed_100__107_, chained_data_delayed_100__106_, chained_data_delayed_100__105_, chained_data_delayed_100__104_, chained_data_delayed_100__103_, chained_data_delayed_100__102_, chained_data_delayed_100__101_, chained_data_delayed_100__100_, chained_data_delayed_100__99_, chained_data_delayed_100__98_, chained_data_delayed_100__97_, chained_data_delayed_100__96_, chained_data_delayed_100__95_, chained_data_delayed_100__94_, chained_data_delayed_100__93_, chained_data_delayed_100__92_, chained_data_delayed_100__91_, chained_data_delayed_100__90_, chained_data_delayed_100__89_, chained_data_delayed_100__88_, chained_data_delayed_100__87_, chained_data_delayed_100__86_, chained_data_delayed_100__85_, chained_data_delayed_100__84_, chained_data_delayed_100__83_, chained_data_delayed_100__82_, chained_data_delayed_100__81_, chained_data_delayed_100__80_, chained_data_delayed_100__79_, chained_data_delayed_100__78_, chained_data_delayed_100__77_, chained_data_delayed_100__76_, chained_data_delayed_100__75_, chained_data_delayed_100__74_, chained_data_delayed_100__73_, chained_data_delayed_100__72_, chained_data_delayed_100__71_, chained_data_delayed_100__70_, chained_data_delayed_100__69_, chained_data_delayed_100__68_, chained_data_delayed_100__67_, chained_data_delayed_100__66_, chained_data_delayed_100__65_, chained_data_delayed_100__64_, chained_data_delayed_100__63_, chained_data_delayed_100__62_, chained_data_delayed_100__61_, chained_data_delayed_100__60_, chained_data_delayed_100__59_, chained_data_delayed_100__58_, chained_data_delayed_100__57_, chained_data_delayed_100__56_, chained_data_delayed_100__55_, chained_data_delayed_100__54_, chained_data_delayed_100__53_, chained_data_delayed_100__52_, chained_data_delayed_100__51_, chained_data_delayed_100__50_, chained_data_delayed_100__49_, chained_data_delayed_100__48_, chained_data_delayed_100__47_, chained_data_delayed_100__46_, chained_data_delayed_100__45_, chained_data_delayed_100__44_, chained_data_delayed_100__43_, chained_data_delayed_100__42_, chained_data_delayed_100__41_, chained_data_delayed_100__40_, chained_data_delayed_100__39_, chained_data_delayed_100__38_, chained_data_delayed_100__37_, chained_data_delayed_100__36_, chained_data_delayed_100__35_, chained_data_delayed_100__34_, chained_data_delayed_100__33_, chained_data_delayed_100__32_, chained_data_delayed_100__31_, chained_data_delayed_100__30_, chained_data_delayed_100__29_, chained_data_delayed_100__28_, chained_data_delayed_100__27_, chained_data_delayed_100__26_, chained_data_delayed_100__25_, chained_data_delayed_100__24_, chained_data_delayed_100__23_, chained_data_delayed_100__22_, chained_data_delayed_100__21_, chained_data_delayed_100__20_, chained_data_delayed_100__19_, chained_data_delayed_100__18_, chained_data_delayed_100__17_, chained_data_delayed_100__16_, chained_data_delayed_100__15_, chained_data_delayed_100__14_, chained_data_delayed_100__13_, chained_data_delayed_100__12_, chained_data_delayed_100__11_, chained_data_delayed_100__10_, chained_data_delayed_100__9_, chained_data_delayed_100__8_, chained_data_delayed_100__7_, chained_data_delayed_100__6_, chained_data_delayed_100__5_, chained_data_delayed_100__4_, chained_data_delayed_100__3_, chained_data_delayed_100__2_, chained_data_delayed_100__1_, chained_data_delayed_100__0_ }),
    .data_o({ chained_data_delayed_101__127_, chained_data_delayed_101__126_, chained_data_delayed_101__125_, chained_data_delayed_101__124_, chained_data_delayed_101__123_, chained_data_delayed_101__122_, chained_data_delayed_101__121_, chained_data_delayed_101__120_, chained_data_delayed_101__119_, chained_data_delayed_101__118_, chained_data_delayed_101__117_, chained_data_delayed_101__116_, chained_data_delayed_101__115_, chained_data_delayed_101__114_, chained_data_delayed_101__113_, chained_data_delayed_101__112_, chained_data_delayed_101__111_, chained_data_delayed_101__110_, chained_data_delayed_101__109_, chained_data_delayed_101__108_, chained_data_delayed_101__107_, chained_data_delayed_101__106_, chained_data_delayed_101__105_, chained_data_delayed_101__104_, chained_data_delayed_101__103_, chained_data_delayed_101__102_, chained_data_delayed_101__101_, chained_data_delayed_101__100_, chained_data_delayed_101__99_, chained_data_delayed_101__98_, chained_data_delayed_101__97_, chained_data_delayed_101__96_, chained_data_delayed_101__95_, chained_data_delayed_101__94_, chained_data_delayed_101__93_, chained_data_delayed_101__92_, chained_data_delayed_101__91_, chained_data_delayed_101__90_, chained_data_delayed_101__89_, chained_data_delayed_101__88_, chained_data_delayed_101__87_, chained_data_delayed_101__86_, chained_data_delayed_101__85_, chained_data_delayed_101__84_, chained_data_delayed_101__83_, chained_data_delayed_101__82_, chained_data_delayed_101__81_, chained_data_delayed_101__80_, chained_data_delayed_101__79_, chained_data_delayed_101__78_, chained_data_delayed_101__77_, chained_data_delayed_101__76_, chained_data_delayed_101__75_, chained_data_delayed_101__74_, chained_data_delayed_101__73_, chained_data_delayed_101__72_, chained_data_delayed_101__71_, chained_data_delayed_101__70_, chained_data_delayed_101__69_, chained_data_delayed_101__68_, chained_data_delayed_101__67_, chained_data_delayed_101__66_, chained_data_delayed_101__65_, chained_data_delayed_101__64_, chained_data_delayed_101__63_, chained_data_delayed_101__62_, chained_data_delayed_101__61_, chained_data_delayed_101__60_, chained_data_delayed_101__59_, chained_data_delayed_101__58_, chained_data_delayed_101__57_, chained_data_delayed_101__56_, chained_data_delayed_101__55_, chained_data_delayed_101__54_, chained_data_delayed_101__53_, chained_data_delayed_101__52_, chained_data_delayed_101__51_, chained_data_delayed_101__50_, chained_data_delayed_101__49_, chained_data_delayed_101__48_, chained_data_delayed_101__47_, chained_data_delayed_101__46_, chained_data_delayed_101__45_, chained_data_delayed_101__44_, chained_data_delayed_101__43_, chained_data_delayed_101__42_, chained_data_delayed_101__41_, chained_data_delayed_101__40_, chained_data_delayed_101__39_, chained_data_delayed_101__38_, chained_data_delayed_101__37_, chained_data_delayed_101__36_, chained_data_delayed_101__35_, chained_data_delayed_101__34_, chained_data_delayed_101__33_, chained_data_delayed_101__32_, chained_data_delayed_101__31_, chained_data_delayed_101__30_, chained_data_delayed_101__29_, chained_data_delayed_101__28_, chained_data_delayed_101__27_, chained_data_delayed_101__26_, chained_data_delayed_101__25_, chained_data_delayed_101__24_, chained_data_delayed_101__23_, chained_data_delayed_101__22_, chained_data_delayed_101__21_, chained_data_delayed_101__20_, chained_data_delayed_101__19_, chained_data_delayed_101__18_, chained_data_delayed_101__17_, chained_data_delayed_101__16_, chained_data_delayed_101__15_, chained_data_delayed_101__14_, chained_data_delayed_101__13_, chained_data_delayed_101__12_, chained_data_delayed_101__11_, chained_data_delayed_101__10_, chained_data_delayed_101__9_, chained_data_delayed_101__8_, chained_data_delayed_101__7_, chained_data_delayed_101__6_, chained_data_delayed_101__5_, chained_data_delayed_101__4_, chained_data_delayed_101__3_, chained_data_delayed_101__2_, chained_data_delayed_101__1_, chained_data_delayed_101__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_102__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_101__127_, chained_data_delayed_101__126_, chained_data_delayed_101__125_, chained_data_delayed_101__124_, chained_data_delayed_101__123_, chained_data_delayed_101__122_, chained_data_delayed_101__121_, chained_data_delayed_101__120_, chained_data_delayed_101__119_, chained_data_delayed_101__118_, chained_data_delayed_101__117_, chained_data_delayed_101__116_, chained_data_delayed_101__115_, chained_data_delayed_101__114_, chained_data_delayed_101__113_, chained_data_delayed_101__112_, chained_data_delayed_101__111_, chained_data_delayed_101__110_, chained_data_delayed_101__109_, chained_data_delayed_101__108_, chained_data_delayed_101__107_, chained_data_delayed_101__106_, chained_data_delayed_101__105_, chained_data_delayed_101__104_, chained_data_delayed_101__103_, chained_data_delayed_101__102_, chained_data_delayed_101__101_, chained_data_delayed_101__100_, chained_data_delayed_101__99_, chained_data_delayed_101__98_, chained_data_delayed_101__97_, chained_data_delayed_101__96_, chained_data_delayed_101__95_, chained_data_delayed_101__94_, chained_data_delayed_101__93_, chained_data_delayed_101__92_, chained_data_delayed_101__91_, chained_data_delayed_101__90_, chained_data_delayed_101__89_, chained_data_delayed_101__88_, chained_data_delayed_101__87_, chained_data_delayed_101__86_, chained_data_delayed_101__85_, chained_data_delayed_101__84_, chained_data_delayed_101__83_, chained_data_delayed_101__82_, chained_data_delayed_101__81_, chained_data_delayed_101__80_, chained_data_delayed_101__79_, chained_data_delayed_101__78_, chained_data_delayed_101__77_, chained_data_delayed_101__76_, chained_data_delayed_101__75_, chained_data_delayed_101__74_, chained_data_delayed_101__73_, chained_data_delayed_101__72_, chained_data_delayed_101__71_, chained_data_delayed_101__70_, chained_data_delayed_101__69_, chained_data_delayed_101__68_, chained_data_delayed_101__67_, chained_data_delayed_101__66_, chained_data_delayed_101__65_, chained_data_delayed_101__64_, chained_data_delayed_101__63_, chained_data_delayed_101__62_, chained_data_delayed_101__61_, chained_data_delayed_101__60_, chained_data_delayed_101__59_, chained_data_delayed_101__58_, chained_data_delayed_101__57_, chained_data_delayed_101__56_, chained_data_delayed_101__55_, chained_data_delayed_101__54_, chained_data_delayed_101__53_, chained_data_delayed_101__52_, chained_data_delayed_101__51_, chained_data_delayed_101__50_, chained_data_delayed_101__49_, chained_data_delayed_101__48_, chained_data_delayed_101__47_, chained_data_delayed_101__46_, chained_data_delayed_101__45_, chained_data_delayed_101__44_, chained_data_delayed_101__43_, chained_data_delayed_101__42_, chained_data_delayed_101__41_, chained_data_delayed_101__40_, chained_data_delayed_101__39_, chained_data_delayed_101__38_, chained_data_delayed_101__37_, chained_data_delayed_101__36_, chained_data_delayed_101__35_, chained_data_delayed_101__34_, chained_data_delayed_101__33_, chained_data_delayed_101__32_, chained_data_delayed_101__31_, chained_data_delayed_101__30_, chained_data_delayed_101__29_, chained_data_delayed_101__28_, chained_data_delayed_101__27_, chained_data_delayed_101__26_, chained_data_delayed_101__25_, chained_data_delayed_101__24_, chained_data_delayed_101__23_, chained_data_delayed_101__22_, chained_data_delayed_101__21_, chained_data_delayed_101__20_, chained_data_delayed_101__19_, chained_data_delayed_101__18_, chained_data_delayed_101__17_, chained_data_delayed_101__16_, chained_data_delayed_101__15_, chained_data_delayed_101__14_, chained_data_delayed_101__13_, chained_data_delayed_101__12_, chained_data_delayed_101__11_, chained_data_delayed_101__10_, chained_data_delayed_101__9_, chained_data_delayed_101__8_, chained_data_delayed_101__7_, chained_data_delayed_101__6_, chained_data_delayed_101__5_, chained_data_delayed_101__4_, chained_data_delayed_101__3_, chained_data_delayed_101__2_, chained_data_delayed_101__1_, chained_data_delayed_101__0_ }),
    .data_o({ chained_data_delayed_102__127_, chained_data_delayed_102__126_, chained_data_delayed_102__125_, chained_data_delayed_102__124_, chained_data_delayed_102__123_, chained_data_delayed_102__122_, chained_data_delayed_102__121_, chained_data_delayed_102__120_, chained_data_delayed_102__119_, chained_data_delayed_102__118_, chained_data_delayed_102__117_, chained_data_delayed_102__116_, chained_data_delayed_102__115_, chained_data_delayed_102__114_, chained_data_delayed_102__113_, chained_data_delayed_102__112_, chained_data_delayed_102__111_, chained_data_delayed_102__110_, chained_data_delayed_102__109_, chained_data_delayed_102__108_, chained_data_delayed_102__107_, chained_data_delayed_102__106_, chained_data_delayed_102__105_, chained_data_delayed_102__104_, chained_data_delayed_102__103_, chained_data_delayed_102__102_, chained_data_delayed_102__101_, chained_data_delayed_102__100_, chained_data_delayed_102__99_, chained_data_delayed_102__98_, chained_data_delayed_102__97_, chained_data_delayed_102__96_, chained_data_delayed_102__95_, chained_data_delayed_102__94_, chained_data_delayed_102__93_, chained_data_delayed_102__92_, chained_data_delayed_102__91_, chained_data_delayed_102__90_, chained_data_delayed_102__89_, chained_data_delayed_102__88_, chained_data_delayed_102__87_, chained_data_delayed_102__86_, chained_data_delayed_102__85_, chained_data_delayed_102__84_, chained_data_delayed_102__83_, chained_data_delayed_102__82_, chained_data_delayed_102__81_, chained_data_delayed_102__80_, chained_data_delayed_102__79_, chained_data_delayed_102__78_, chained_data_delayed_102__77_, chained_data_delayed_102__76_, chained_data_delayed_102__75_, chained_data_delayed_102__74_, chained_data_delayed_102__73_, chained_data_delayed_102__72_, chained_data_delayed_102__71_, chained_data_delayed_102__70_, chained_data_delayed_102__69_, chained_data_delayed_102__68_, chained_data_delayed_102__67_, chained_data_delayed_102__66_, chained_data_delayed_102__65_, chained_data_delayed_102__64_, chained_data_delayed_102__63_, chained_data_delayed_102__62_, chained_data_delayed_102__61_, chained_data_delayed_102__60_, chained_data_delayed_102__59_, chained_data_delayed_102__58_, chained_data_delayed_102__57_, chained_data_delayed_102__56_, chained_data_delayed_102__55_, chained_data_delayed_102__54_, chained_data_delayed_102__53_, chained_data_delayed_102__52_, chained_data_delayed_102__51_, chained_data_delayed_102__50_, chained_data_delayed_102__49_, chained_data_delayed_102__48_, chained_data_delayed_102__47_, chained_data_delayed_102__46_, chained_data_delayed_102__45_, chained_data_delayed_102__44_, chained_data_delayed_102__43_, chained_data_delayed_102__42_, chained_data_delayed_102__41_, chained_data_delayed_102__40_, chained_data_delayed_102__39_, chained_data_delayed_102__38_, chained_data_delayed_102__37_, chained_data_delayed_102__36_, chained_data_delayed_102__35_, chained_data_delayed_102__34_, chained_data_delayed_102__33_, chained_data_delayed_102__32_, chained_data_delayed_102__31_, chained_data_delayed_102__30_, chained_data_delayed_102__29_, chained_data_delayed_102__28_, chained_data_delayed_102__27_, chained_data_delayed_102__26_, chained_data_delayed_102__25_, chained_data_delayed_102__24_, chained_data_delayed_102__23_, chained_data_delayed_102__22_, chained_data_delayed_102__21_, chained_data_delayed_102__20_, chained_data_delayed_102__19_, chained_data_delayed_102__18_, chained_data_delayed_102__17_, chained_data_delayed_102__16_, chained_data_delayed_102__15_, chained_data_delayed_102__14_, chained_data_delayed_102__13_, chained_data_delayed_102__12_, chained_data_delayed_102__11_, chained_data_delayed_102__10_, chained_data_delayed_102__9_, chained_data_delayed_102__8_, chained_data_delayed_102__7_, chained_data_delayed_102__6_, chained_data_delayed_102__5_, chained_data_delayed_102__4_, chained_data_delayed_102__3_, chained_data_delayed_102__2_, chained_data_delayed_102__1_, chained_data_delayed_102__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_103__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_102__127_, chained_data_delayed_102__126_, chained_data_delayed_102__125_, chained_data_delayed_102__124_, chained_data_delayed_102__123_, chained_data_delayed_102__122_, chained_data_delayed_102__121_, chained_data_delayed_102__120_, chained_data_delayed_102__119_, chained_data_delayed_102__118_, chained_data_delayed_102__117_, chained_data_delayed_102__116_, chained_data_delayed_102__115_, chained_data_delayed_102__114_, chained_data_delayed_102__113_, chained_data_delayed_102__112_, chained_data_delayed_102__111_, chained_data_delayed_102__110_, chained_data_delayed_102__109_, chained_data_delayed_102__108_, chained_data_delayed_102__107_, chained_data_delayed_102__106_, chained_data_delayed_102__105_, chained_data_delayed_102__104_, chained_data_delayed_102__103_, chained_data_delayed_102__102_, chained_data_delayed_102__101_, chained_data_delayed_102__100_, chained_data_delayed_102__99_, chained_data_delayed_102__98_, chained_data_delayed_102__97_, chained_data_delayed_102__96_, chained_data_delayed_102__95_, chained_data_delayed_102__94_, chained_data_delayed_102__93_, chained_data_delayed_102__92_, chained_data_delayed_102__91_, chained_data_delayed_102__90_, chained_data_delayed_102__89_, chained_data_delayed_102__88_, chained_data_delayed_102__87_, chained_data_delayed_102__86_, chained_data_delayed_102__85_, chained_data_delayed_102__84_, chained_data_delayed_102__83_, chained_data_delayed_102__82_, chained_data_delayed_102__81_, chained_data_delayed_102__80_, chained_data_delayed_102__79_, chained_data_delayed_102__78_, chained_data_delayed_102__77_, chained_data_delayed_102__76_, chained_data_delayed_102__75_, chained_data_delayed_102__74_, chained_data_delayed_102__73_, chained_data_delayed_102__72_, chained_data_delayed_102__71_, chained_data_delayed_102__70_, chained_data_delayed_102__69_, chained_data_delayed_102__68_, chained_data_delayed_102__67_, chained_data_delayed_102__66_, chained_data_delayed_102__65_, chained_data_delayed_102__64_, chained_data_delayed_102__63_, chained_data_delayed_102__62_, chained_data_delayed_102__61_, chained_data_delayed_102__60_, chained_data_delayed_102__59_, chained_data_delayed_102__58_, chained_data_delayed_102__57_, chained_data_delayed_102__56_, chained_data_delayed_102__55_, chained_data_delayed_102__54_, chained_data_delayed_102__53_, chained_data_delayed_102__52_, chained_data_delayed_102__51_, chained_data_delayed_102__50_, chained_data_delayed_102__49_, chained_data_delayed_102__48_, chained_data_delayed_102__47_, chained_data_delayed_102__46_, chained_data_delayed_102__45_, chained_data_delayed_102__44_, chained_data_delayed_102__43_, chained_data_delayed_102__42_, chained_data_delayed_102__41_, chained_data_delayed_102__40_, chained_data_delayed_102__39_, chained_data_delayed_102__38_, chained_data_delayed_102__37_, chained_data_delayed_102__36_, chained_data_delayed_102__35_, chained_data_delayed_102__34_, chained_data_delayed_102__33_, chained_data_delayed_102__32_, chained_data_delayed_102__31_, chained_data_delayed_102__30_, chained_data_delayed_102__29_, chained_data_delayed_102__28_, chained_data_delayed_102__27_, chained_data_delayed_102__26_, chained_data_delayed_102__25_, chained_data_delayed_102__24_, chained_data_delayed_102__23_, chained_data_delayed_102__22_, chained_data_delayed_102__21_, chained_data_delayed_102__20_, chained_data_delayed_102__19_, chained_data_delayed_102__18_, chained_data_delayed_102__17_, chained_data_delayed_102__16_, chained_data_delayed_102__15_, chained_data_delayed_102__14_, chained_data_delayed_102__13_, chained_data_delayed_102__12_, chained_data_delayed_102__11_, chained_data_delayed_102__10_, chained_data_delayed_102__9_, chained_data_delayed_102__8_, chained_data_delayed_102__7_, chained_data_delayed_102__6_, chained_data_delayed_102__5_, chained_data_delayed_102__4_, chained_data_delayed_102__3_, chained_data_delayed_102__2_, chained_data_delayed_102__1_, chained_data_delayed_102__0_ }),
    .data_o({ chained_data_delayed_103__127_, chained_data_delayed_103__126_, chained_data_delayed_103__125_, chained_data_delayed_103__124_, chained_data_delayed_103__123_, chained_data_delayed_103__122_, chained_data_delayed_103__121_, chained_data_delayed_103__120_, chained_data_delayed_103__119_, chained_data_delayed_103__118_, chained_data_delayed_103__117_, chained_data_delayed_103__116_, chained_data_delayed_103__115_, chained_data_delayed_103__114_, chained_data_delayed_103__113_, chained_data_delayed_103__112_, chained_data_delayed_103__111_, chained_data_delayed_103__110_, chained_data_delayed_103__109_, chained_data_delayed_103__108_, chained_data_delayed_103__107_, chained_data_delayed_103__106_, chained_data_delayed_103__105_, chained_data_delayed_103__104_, chained_data_delayed_103__103_, chained_data_delayed_103__102_, chained_data_delayed_103__101_, chained_data_delayed_103__100_, chained_data_delayed_103__99_, chained_data_delayed_103__98_, chained_data_delayed_103__97_, chained_data_delayed_103__96_, chained_data_delayed_103__95_, chained_data_delayed_103__94_, chained_data_delayed_103__93_, chained_data_delayed_103__92_, chained_data_delayed_103__91_, chained_data_delayed_103__90_, chained_data_delayed_103__89_, chained_data_delayed_103__88_, chained_data_delayed_103__87_, chained_data_delayed_103__86_, chained_data_delayed_103__85_, chained_data_delayed_103__84_, chained_data_delayed_103__83_, chained_data_delayed_103__82_, chained_data_delayed_103__81_, chained_data_delayed_103__80_, chained_data_delayed_103__79_, chained_data_delayed_103__78_, chained_data_delayed_103__77_, chained_data_delayed_103__76_, chained_data_delayed_103__75_, chained_data_delayed_103__74_, chained_data_delayed_103__73_, chained_data_delayed_103__72_, chained_data_delayed_103__71_, chained_data_delayed_103__70_, chained_data_delayed_103__69_, chained_data_delayed_103__68_, chained_data_delayed_103__67_, chained_data_delayed_103__66_, chained_data_delayed_103__65_, chained_data_delayed_103__64_, chained_data_delayed_103__63_, chained_data_delayed_103__62_, chained_data_delayed_103__61_, chained_data_delayed_103__60_, chained_data_delayed_103__59_, chained_data_delayed_103__58_, chained_data_delayed_103__57_, chained_data_delayed_103__56_, chained_data_delayed_103__55_, chained_data_delayed_103__54_, chained_data_delayed_103__53_, chained_data_delayed_103__52_, chained_data_delayed_103__51_, chained_data_delayed_103__50_, chained_data_delayed_103__49_, chained_data_delayed_103__48_, chained_data_delayed_103__47_, chained_data_delayed_103__46_, chained_data_delayed_103__45_, chained_data_delayed_103__44_, chained_data_delayed_103__43_, chained_data_delayed_103__42_, chained_data_delayed_103__41_, chained_data_delayed_103__40_, chained_data_delayed_103__39_, chained_data_delayed_103__38_, chained_data_delayed_103__37_, chained_data_delayed_103__36_, chained_data_delayed_103__35_, chained_data_delayed_103__34_, chained_data_delayed_103__33_, chained_data_delayed_103__32_, chained_data_delayed_103__31_, chained_data_delayed_103__30_, chained_data_delayed_103__29_, chained_data_delayed_103__28_, chained_data_delayed_103__27_, chained_data_delayed_103__26_, chained_data_delayed_103__25_, chained_data_delayed_103__24_, chained_data_delayed_103__23_, chained_data_delayed_103__22_, chained_data_delayed_103__21_, chained_data_delayed_103__20_, chained_data_delayed_103__19_, chained_data_delayed_103__18_, chained_data_delayed_103__17_, chained_data_delayed_103__16_, chained_data_delayed_103__15_, chained_data_delayed_103__14_, chained_data_delayed_103__13_, chained_data_delayed_103__12_, chained_data_delayed_103__11_, chained_data_delayed_103__10_, chained_data_delayed_103__9_, chained_data_delayed_103__8_, chained_data_delayed_103__7_, chained_data_delayed_103__6_, chained_data_delayed_103__5_, chained_data_delayed_103__4_, chained_data_delayed_103__3_, chained_data_delayed_103__2_, chained_data_delayed_103__1_, chained_data_delayed_103__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_104__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_103__127_, chained_data_delayed_103__126_, chained_data_delayed_103__125_, chained_data_delayed_103__124_, chained_data_delayed_103__123_, chained_data_delayed_103__122_, chained_data_delayed_103__121_, chained_data_delayed_103__120_, chained_data_delayed_103__119_, chained_data_delayed_103__118_, chained_data_delayed_103__117_, chained_data_delayed_103__116_, chained_data_delayed_103__115_, chained_data_delayed_103__114_, chained_data_delayed_103__113_, chained_data_delayed_103__112_, chained_data_delayed_103__111_, chained_data_delayed_103__110_, chained_data_delayed_103__109_, chained_data_delayed_103__108_, chained_data_delayed_103__107_, chained_data_delayed_103__106_, chained_data_delayed_103__105_, chained_data_delayed_103__104_, chained_data_delayed_103__103_, chained_data_delayed_103__102_, chained_data_delayed_103__101_, chained_data_delayed_103__100_, chained_data_delayed_103__99_, chained_data_delayed_103__98_, chained_data_delayed_103__97_, chained_data_delayed_103__96_, chained_data_delayed_103__95_, chained_data_delayed_103__94_, chained_data_delayed_103__93_, chained_data_delayed_103__92_, chained_data_delayed_103__91_, chained_data_delayed_103__90_, chained_data_delayed_103__89_, chained_data_delayed_103__88_, chained_data_delayed_103__87_, chained_data_delayed_103__86_, chained_data_delayed_103__85_, chained_data_delayed_103__84_, chained_data_delayed_103__83_, chained_data_delayed_103__82_, chained_data_delayed_103__81_, chained_data_delayed_103__80_, chained_data_delayed_103__79_, chained_data_delayed_103__78_, chained_data_delayed_103__77_, chained_data_delayed_103__76_, chained_data_delayed_103__75_, chained_data_delayed_103__74_, chained_data_delayed_103__73_, chained_data_delayed_103__72_, chained_data_delayed_103__71_, chained_data_delayed_103__70_, chained_data_delayed_103__69_, chained_data_delayed_103__68_, chained_data_delayed_103__67_, chained_data_delayed_103__66_, chained_data_delayed_103__65_, chained_data_delayed_103__64_, chained_data_delayed_103__63_, chained_data_delayed_103__62_, chained_data_delayed_103__61_, chained_data_delayed_103__60_, chained_data_delayed_103__59_, chained_data_delayed_103__58_, chained_data_delayed_103__57_, chained_data_delayed_103__56_, chained_data_delayed_103__55_, chained_data_delayed_103__54_, chained_data_delayed_103__53_, chained_data_delayed_103__52_, chained_data_delayed_103__51_, chained_data_delayed_103__50_, chained_data_delayed_103__49_, chained_data_delayed_103__48_, chained_data_delayed_103__47_, chained_data_delayed_103__46_, chained_data_delayed_103__45_, chained_data_delayed_103__44_, chained_data_delayed_103__43_, chained_data_delayed_103__42_, chained_data_delayed_103__41_, chained_data_delayed_103__40_, chained_data_delayed_103__39_, chained_data_delayed_103__38_, chained_data_delayed_103__37_, chained_data_delayed_103__36_, chained_data_delayed_103__35_, chained_data_delayed_103__34_, chained_data_delayed_103__33_, chained_data_delayed_103__32_, chained_data_delayed_103__31_, chained_data_delayed_103__30_, chained_data_delayed_103__29_, chained_data_delayed_103__28_, chained_data_delayed_103__27_, chained_data_delayed_103__26_, chained_data_delayed_103__25_, chained_data_delayed_103__24_, chained_data_delayed_103__23_, chained_data_delayed_103__22_, chained_data_delayed_103__21_, chained_data_delayed_103__20_, chained_data_delayed_103__19_, chained_data_delayed_103__18_, chained_data_delayed_103__17_, chained_data_delayed_103__16_, chained_data_delayed_103__15_, chained_data_delayed_103__14_, chained_data_delayed_103__13_, chained_data_delayed_103__12_, chained_data_delayed_103__11_, chained_data_delayed_103__10_, chained_data_delayed_103__9_, chained_data_delayed_103__8_, chained_data_delayed_103__7_, chained_data_delayed_103__6_, chained_data_delayed_103__5_, chained_data_delayed_103__4_, chained_data_delayed_103__3_, chained_data_delayed_103__2_, chained_data_delayed_103__1_, chained_data_delayed_103__0_ }),
    .data_o({ chained_data_delayed_104__127_, chained_data_delayed_104__126_, chained_data_delayed_104__125_, chained_data_delayed_104__124_, chained_data_delayed_104__123_, chained_data_delayed_104__122_, chained_data_delayed_104__121_, chained_data_delayed_104__120_, chained_data_delayed_104__119_, chained_data_delayed_104__118_, chained_data_delayed_104__117_, chained_data_delayed_104__116_, chained_data_delayed_104__115_, chained_data_delayed_104__114_, chained_data_delayed_104__113_, chained_data_delayed_104__112_, chained_data_delayed_104__111_, chained_data_delayed_104__110_, chained_data_delayed_104__109_, chained_data_delayed_104__108_, chained_data_delayed_104__107_, chained_data_delayed_104__106_, chained_data_delayed_104__105_, chained_data_delayed_104__104_, chained_data_delayed_104__103_, chained_data_delayed_104__102_, chained_data_delayed_104__101_, chained_data_delayed_104__100_, chained_data_delayed_104__99_, chained_data_delayed_104__98_, chained_data_delayed_104__97_, chained_data_delayed_104__96_, chained_data_delayed_104__95_, chained_data_delayed_104__94_, chained_data_delayed_104__93_, chained_data_delayed_104__92_, chained_data_delayed_104__91_, chained_data_delayed_104__90_, chained_data_delayed_104__89_, chained_data_delayed_104__88_, chained_data_delayed_104__87_, chained_data_delayed_104__86_, chained_data_delayed_104__85_, chained_data_delayed_104__84_, chained_data_delayed_104__83_, chained_data_delayed_104__82_, chained_data_delayed_104__81_, chained_data_delayed_104__80_, chained_data_delayed_104__79_, chained_data_delayed_104__78_, chained_data_delayed_104__77_, chained_data_delayed_104__76_, chained_data_delayed_104__75_, chained_data_delayed_104__74_, chained_data_delayed_104__73_, chained_data_delayed_104__72_, chained_data_delayed_104__71_, chained_data_delayed_104__70_, chained_data_delayed_104__69_, chained_data_delayed_104__68_, chained_data_delayed_104__67_, chained_data_delayed_104__66_, chained_data_delayed_104__65_, chained_data_delayed_104__64_, chained_data_delayed_104__63_, chained_data_delayed_104__62_, chained_data_delayed_104__61_, chained_data_delayed_104__60_, chained_data_delayed_104__59_, chained_data_delayed_104__58_, chained_data_delayed_104__57_, chained_data_delayed_104__56_, chained_data_delayed_104__55_, chained_data_delayed_104__54_, chained_data_delayed_104__53_, chained_data_delayed_104__52_, chained_data_delayed_104__51_, chained_data_delayed_104__50_, chained_data_delayed_104__49_, chained_data_delayed_104__48_, chained_data_delayed_104__47_, chained_data_delayed_104__46_, chained_data_delayed_104__45_, chained_data_delayed_104__44_, chained_data_delayed_104__43_, chained_data_delayed_104__42_, chained_data_delayed_104__41_, chained_data_delayed_104__40_, chained_data_delayed_104__39_, chained_data_delayed_104__38_, chained_data_delayed_104__37_, chained_data_delayed_104__36_, chained_data_delayed_104__35_, chained_data_delayed_104__34_, chained_data_delayed_104__33_, chained_data_delayed_104__32_, chained_data_delayed_104__31_, chained_data_delayed_104__30_, chained_data_delayed_104__29_, chained_data_delayed_104__28_, chained_data_delayed_104__27_, chained_data_delayed_104__26_, chained_data_delayed_104__25_, chained_data_delayed_104__24_, chained_data_delayed_104__23_, chained_data_delayed_104__22_, chained_data_delayed_104__21_, chained_data_delayed_104__20_, chained_data_delayed_104__19_, chained_data_delayed_104__18_, chained_data_delayed_104__17_, chained_data_delayed_104__16_, chained_data_delayed_104__15_, chained_data_delayed_104__14_, chained_data_delayed_104__13_, chained_data_delayed_104__12_, chained_data_delayed_104__11_, chained_data_delayed_104__10_, chained_data_delayed_104__9_, chained_data_delayed_104__8_, chained_data_delayed_104__7_, chained_data_delayed_104__6_, chained_data_delayed_104__5_, chained_data_delayed_104__4_, chained_data_delayed_104__3_, chained_data_delayed_104__2_, chained_data_delayed_104__1_, chained_data_delayed_104__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_105__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_104__127_, chained_data_delayed_104__126_, chained_data_delayed_104__125_, chained_data_delayed_104__124_, chained_data_delayed_104__123_, chained_data_delayed_104__122_, chained_data_delayed_104__121_, chained_data_delayed_104__120_, chained_data_delayed_104__119_, chained_data_delayed_104__118_, chained_data_delayed_104__117_, chained_data_delayed_104__116_, chained_data_delayed_104__115_, chained_data_delayed_104__114_, chained_data_delayed_104__113_, chained_data_delayed_104__112_, chained_data_delayed_104__111_, chained_data_delayed_104__110_, chained_data_delayed_104__109_, chained_data_delayed_104__108_, chained_data_delayed_104__107_, chained_data_delayed_104__106_, chained_data_delayed_104__105_, chained_data_delayed_104__104_, chained_data_delayed_104__103_, chained_data_delayed_104__102_, chained_data_delayed_104__101_, chained_data_delayed_104__100_, chained_data_delayed_104__99_, chained_data_delayed_104__98_, chained_data_delayed_104__97_, chained_data_delayed_104__96_, chained_data_delayed_104__95_, chained_data_delayed_104__94_, chained_data_delayed_104__93_, chained_data_delayed_104__92_, chained_data_delayed_104__91_, chained_data_delayed_104__90_, chained_data_delayed_104__89_, chained_data_delayed_104__88_, chained_data_delayed_104__87_, chained_data_delayed_104__86_, chained_data_delayed_104__85_, chained_data_delayed_104__84_, chained_data_delayed_104__83_, chained_data_delayed_104__82_, chained_data_delayed_104__81_, chained_data_delayed_104__80_, chained_data_delayed_104__79_, chained_data_delayed_104__78_, chained_data_delayed_104__77_, chained_data_delayed_104__76_, chained_data_delayed_104__75_, chained_data_delayed_104__74_, chained_data_delayed_104__73_, chained_data_delayed_104__72_, chained_data_delayed_104__71_, chained_data_delayed_104__70_, chained_data_delayed_104__69_, chained_data_delayed_104__68_, chained_data_delayed_104__67_, chained_data_delayed_104__66_, chained_data_delayed_104__65_, chained_data_delayed_104__64_, chained_data_delayed_104__63_, chained_data_delayed_104__62_, chained_data_delayed_104__61_, chained_data_delayed_104__60_, chained_data_delayed_104__59_, chained_data_delayed_104__58_, chained_data_delayed_104__57_, chained_data_delayed_104__56_, chained_data_delayed_104__55_, chained_data_delayed_104__54_, chained_data_delayed_104__53_, chained_data_delayed_104__52_, chained_data_delayed_104__51_, chained_data_delayed_104__50_, chained_data_delayed_104__49_, chained_data_delayed_104__48_, chained_data_delayed_104__47_, chained_data_delayed_104__46_, chained_data_delayed_104__45_, chained_data_delayed_104__44_, chained_data_delayed_104__43_, chained_data_delayed_104__42_, chained_data_delayed_104__41_, chained_data_delayed_104__40_, chained_data_delayed_104__39_, chained_data_delayed_104__38_, chained_data_delayed_104__37_, chained_data_delayed_104__36_, chained_data_delayed_104__35_, chained_data_delayed_104__34_, chained_data_delayed_104__33_, chained_data_delayed_104__32_, chained_data_delayed_104__31_, chained_data_delayed_104__30_, chained_data_delayed_104__29_, chained_data_delayed_104__28_, chained_data_delayed_104__27_, chained_data_delayed_104__26_, chained_data_delayed_104__25_, chained_data_delayed_104__24_, chained_data_delayed_104__23_, chained_data_delayed_104__22_, chained_data_delayed_104__21_, chained_data_delayed_104__20_, chained_data_delayed_104__19_, chained_data_delayed_104__18_, chained_data_delayed_104__17_, chained_data_delayed_104__16_, chained_data_delayed_104__15_, chained_data_delayed_104__14_, chained_data_delayed_104__13_, chained_data_delayed_104__12_, chained_data_delayed_104__11_, chained_data_delayed_104__10_, chained_data_delayed_104__9_, chained_data_delayed_104__8_, chained_data_delayed_104__7_, chained_data_delayed_104__6_, chained_data_delayed_104__5_, chained_data_delayed_104__4_, chained_data_delayed_104__3_, chained_data_delayed_104__2_, chained_data_delayed_104__1_, chained_data_delayed_104__0_ }),
    .data_o({ chained_data_delayed_105__127_, chained_data_delayed_105__126_, chained_data_delayed_105__125_, chained_data_delayed_105__124_, chained_data_delayed_105__123_, chained_data_delayed_105__122_, chained_data_delayed_105__121_, chained_data_delayed_105__120_, chained_data_delayed_105__119_, chained_data_delayed_105__118_, chained_data_delayed_105__117_, chained_data_delayed_105__116_, chained_data_delayed_105__115_, chained_data_delayed_105__114_, chained_data_delayed_105__113_, chained_data_delayed_105__112_, chained_data_delayed_105__111_, chained_data_delayed_105__110_, chained_data_delayed_105__109_, chained_data_delayed_105__108_, chained_data_delayed_105__107_, chained_data_delayed_105__106_, chained_data_delayed_105__105_, chained_data_delayed_105__104_, chained_data_delayed_105__103_, chained_data_delayed_105__102_, chained_data_delayed_105__101_, chained_data_delayed_105__100_, chained_data_delayed_105__99_, chained_data_delayed_105__98_, chained_data_delayed_105__97_, chained_data_delayed_105__96_, chained_data_delayed_105__95_, chained_data_delayed_105__94_, chained_data_delayed_105__93_, chained_data_delayed_105__92_, chained_data_delayed_105__91_, chained_data_delayed_105__90_, chained_data_delayed_105__89_, chained_data_delayed_105__88_, chained_data_delayed_105__87_, chained_data_delayed_105__86_, chained_data_delayed_105__85_, chained_data_delayed_105__84_, chained_data_delayed_105__83_, chained_data_delayed_105__82_, chained_data_delayed_105__81_, chained_data_delayed_105__80_, chained_data_delayed_105__79_, chained_data_delayed_105__78_, chained_data_delayed_105__77_, chained_data_delayed_105__76_, chained_data_delayed_105__75_, chained_data_delayed_105__74_, chained_data_delayed_105__73_, chained_data_delayed_105__72_, chained_data_delayed_105__71_, chained_data_delayed_105__70_, chained_data_delayed_105__69_, chained_data_delayed_105__68_, chained_data_delayed_105__67_, chained_data_delayed_105__66_, chained_data_delayed_105__65_, chained_data_delayed_105__64_, chained_data_delayed_105__63_, chained_data_delayed_105__62_, chained_data_delayed_105__61_, chained_data_delayed_105__60_, chained_data_delayed_105__59_, chained_data_delayed_105__58_, chained_data_delayed_105__57_, chained_data_delayed_105__56_, chained_data_delayed_105__55_, chained_data_delayed_105__54_, chained_data_delayed_105__53_, chained_data_delayed_105__52_, chained_data_delayed_105__51_, chained_data_delayed_105__50_, chained_data_delayed_105__49_, chained_data_delayed_105__48_, chained_data_delayed_105__47_, chained_data_delayed_105__46_, chained_data_delayed_105__45_, chained_data_delayed_105__44_, chained_data_delayed_105__43_, chained_data_delayed_105__42_, chained_data_delayed_105__41_, chained_data_delayed_105__40_, chained_data_delayed_105__39_, chained_data_delayed_105__38_, chained_data_delayed_105__37_, chained_data_delayed_105__36_, chained_data_delayed_105__35_, chained_data_delayed_105__34_, chained_data_delayed_105__33_, chained_data_delayed_105__32_, chained_data_delayed_105__31_, chained_data_delayed_105__30_, chained_data_delayed_105__29_, chained_data_delayed_105__28_, chained_data_delayed_105__27_, chained_data_delayed_105__26_, chained_data_delayed_105__25_, chained_data_delayed_105__24_, chained_data_delayed_105__23_, chained_data_delayed_105__22_, chained_data_delayed_105__21_, chained_data_delayed_105__20_, chained_data_delayed_105__19_, chained_data_delayed_105__18_, chained_data_delayed_105__17_, chained_data_delayed_105__16_, chained_data_delayed_105__15_, chained_data_delayed_105__14_, chained_data_delayed_105__13_, chained_data_delayed_105__12_, chained_data_delayed_105__11_, chained_data_delayed_105__10_, chained_data_delayed_105__9_, chained_data_delayed_105__8_, chained_data_delayed_105__7_, chained_data_delayed_105__6_, chained_data_delayed_105__5_, chained_data_delayed_105__4_, chained_data_delayed_105__3_, chained_data_delayed_105__2_, chained_data_delayed_105__1_, chained_data_delayed_105__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_106__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_105__127_, chained_data_delayed_105__126_, chained_data_delayed_105__125_, chained_data_delayed_105__124_, chained_data_delayed_105__123_, chained_data_delayed_105__122_, chained_data_delayed_105__121_, chained_data_delayed_105__120_, chained_data_delayed_105__119_, chained_data_delayed_105__118_, chained_data_delayed_105__117_, chained_data_delayed_105__116_, chained_data_delayed_105__115_, chained_data_delayed_105__114_, chained_data_delayed_105__113_, chained_data_delayed_105__112_, chained_data_delayed_105__111_, chained_data_delayed_105__110_, chained_data_delayed_105__109_, chained_data_delayed_105__108_, chained_data_delayed_105__107_, chained_data_delayed_105__106_, chained_data_delayed_105__105_, chained_data_delayed_105__104_, chained_data_delayed_105__103_, chained_data_delayed_105__102_, chained_data_delayed_105__101_, chained_data_delayed_105__100_, chained_data_delayed_105__99_, chained_data_delayed_105__98_, chained_data_delayed_105__97_, chained_data_delayed_105__96_, chained_data_delayed_105__95_, chained_data_delayed_105__94_, chained_data_delayed_105__93_, chained_data_delayed_105__92_, chained_data_delayed_105__91_, chained_data_delayed_105__90_, chained_data_delayed_105__89_, chained_data_delayed_105__88_, chained_data_delayed_105__87_, chained_data_delayed_105__86_, chained_data_delayed_105__85_, chained_data_delayed_105__84_, chained_data_delayed_105__83_, chained_data_delayed_105__82_, chained_data_delayed_105__81_, chained_data_delayed_105__80_, chained_data_delayed_105__79_, chained_data_delayed_105__78_, chained_data_delayed_105__77_, chained_data_delayed_105__76_, chained_data_delayed_105__75_, chained_data_delayed_105__74_, chained_data_delayed_105__73_, chained_data_delayed_105__72_, chained_data_delayed_105__71_, chained_data_delayed_105__70_, chained_data_delayed_105__69_, chained_data_delayed_105__68_, chained_data_delayed_105__67_, chained_data_delayed_105__66_, chained_data_delayed_105__65_, chained_data_delayed_105__64_, chained_data_delayed_105__63_, chained_data_delayed_105__62_, chained_data_delayed_105__61_, chained_data_delayed_105__60_, chained_data_delayed_105__59_, chained_data_delayed_105__58_, chained_data_delayed_105__57_, chained_data_delayed_105__56_, chained_data_delayed_105__55_, chained_data_delayed_105__54_, chained_data_delayed_105__53_, chained_data_delayed_105__52_, chained_data_delayed_105__51_, chained_data_delayed_105__50_, chained_data_delayed_105__49_, chained_data_delayed_105__48_, chained_data_delayed_105__47_, chained_data_delayed_105__46_, chained_data_delayed_105__45_, chained_data_delayed_105__44_, chained_data_delayed_105__43_, chained_data_delayed_105__42_, chained_data_delayed_105__41_, chained_data_delayed_105__40_, chained_data_delayed_105__39_, chained_data_delayed_105__38_, chained_data_delayed_105__37_, chained_data_delayed_105__36_, chained_data_delayed_105__35_, chained_data_delayed_105__34_, chained_data_delayed_105__33_, chained_data_delayed_105__32_, chained_data_delayed_105__31_, chained_data_delayed_105__30_, chained_data_delayed_105__29_, chained_data_delayed_105__28_, chained_data_delayed_105__27_, chained_data_delayed_105__26_, chained_data_delayed_105__25_, chained_data_delayed_105__24_, chained_data_delayed_105__23_, chained_data_delayed_105__22_, chained_data_delayed_105__21_, chained_data_delayed_105__20_, chained_data_delayed_105__19_, chained_data_delayed_105__18_, chained_data_delayed_105__17_, chained_data_delayed_105__16_, chained_data_delayed_105__15_, chained_data_delayed_105__14_, chained_data_delayed_105__13_, chained_data_delayed_105__12_, chained_data_delayed_105__11_, chained_data_delayed_105__10_, chained_data_delayed_105__9_, chained_data_delayed_105__8_, chained_data_delayed_105__7_, chained_data_delayed_105__6_, chained_data_delayed_105__5_, chained_data_delayed_105__4_, chained_data_delayed_105__3_, chained_data_delayed_105__2_, chained_data_delayed_105__1_, chained_data_delayed_105__0_ }),
    .data_o({ chained_data_delayed_106__127_, chained_data_delayed_106__126_, chained_data_delayed_106__125_, chained_data_delayed_106__124_, chained_data_delayed_106__123_, chained_data_delayed_106__122_, chained_data_delayed_106__121_, chained_data_delayed_106__120_, chained_data_delayed_106__119_, chained_data_delayed_106__118_, chained_data_delayed_106__117_, chained_data_delayed_106__116_, chained_data_delayed_106__115_, chained_data_delayed_106__114_, chained_data_delayed_106__113_, chained_data_delayed_106__112_, chained_data_delayed_106__111_, chained_data_delayed_106__110_, chained_data_delayed_106__109_, chained_data_delayed_106__108_, chained_data_delayed_106__107_, chained_data_delayed_106__106_, chained_data_delayed_106__105_, chained_data_delayed_106__104_, chained_data_delayed_106__103_, chained_data_delayed_106__102_, chained_data_delayed_106__101_, chained_data_delayed_106__100_, chained_data_delayed_106__99_, chained_data_delayed_106__98_, chained_data_delayed_106__97_, chained_data_delayed_106__96_, chained_data_delayed_106__95_, chained_data_delayed_106__94_, chained_data_delayed_106__93_, chained_data_delayed_106__92_, chained_data_delayed_106__91_, chained_data_delayed_106__90_, chained_data_delayed_106__89_, chained_data_delayed_106__88_, chained_data_delayed_106__87_, chained_data_delayed_106__86_, chained_data_delayed_106__85_, chained_data_delayed_106__84_, chained_data_delayed_106__83_, chained_data_delayed_106__82_, chained_data_delayed_106__81_, chained_data_delayed_106__80_, chained_data_delayed_106__79_, chained_data_delayed_106__78_, chained_data_delayed_106__77_, chained_data_delayed_106__76_, chained_data_delayed_106__75_, chained_data_delayed_106__74_, chained_data_delayed_106__73_, chained_data_delayed_106__72_, chained_data_delayed_106__71_, chained_data_delayed_106__70_, chained_data_delayed_106__69_, chained_data_delayed_106__68_, chained_data_delayed_106__67_, chained_data_delayed_106__66_, chained_data_delayed_106__65_, chained_data_delayed_106__64_, chained_data_delayed_106__63_, chained_data_delayed_106__62_, chained_data_delayed_106__61_, chained_data_delayed_106__60_, chained_data_delayed_106__59_, chained_data_delayed_106__58_, chained_data_delayed_106__57_, chained_data_delayed_106__56_, chained_data_delayed_106__55_, chained_data_delayed_106__54_, chained_data_delayed_106__53_, chained_data_delayed_106__52_, chained_data_delayed_106__51_, chained_data_delayed_106__50_, chained_data_delayed_106__49_, chained_data_delayed_106__48_, chained_data_delayed_106__47_, chained_data_delayed_106__46_, chained_data_delayed_106__45_, chained_data_delayed_106__44_, chained_data_delayed_106__43_, chained_data_delayed_106__42_, chained_data_delayed_106__41_, chained_data_delayed_106__40_, chained_data_delayed_106__39_, chained_data_delayed_106__38_, chained_data_delayed_106__37_, chained_data_delayed_106__36_, chained_data_delayed_106__35_, chained_data_delayed_106__34_, chained_data_delayed_106__33_, chained_data_delayed_106__32_, chained_data_delayed_106__31_, chained_data_delayed_106__30_, chained_data_delayed_106__29_, chained_data_delayed_106__28_, chained_data_delayed_106__27_, chained_data_delayed_106__26_, chained_data_delayed_106__25_, chained_data_delayed_106__24_, chained_data_delayed_106__23_, chained_data_delayed_106__22_, chained_data_delayed_106__21_, chained_data_delayed_106__20_, chained_data_delayed_106__19_, chained_data_delayed_106__18_, chained_data_delayed_106__17_, chained_data_delayed_106__16_, chained_data_delayed_106__15_, chained_data_delayed_106__14_, chained_data_delayed_106__13_, chained_data_delayed_106__12_, chained_data_delayed_106__11_, chained_data_delayed_106__10_, chained_data_delayed_106__9_, chained_data_delayed_106__8_, chained_data_delayed_106__7_, chained_data_delayed_106__6_, chained_data_delayed_106__5_, chained_data_delayed_106__4_, chained_data_delayed_106__3_, chained_data_delayed_106__2_, chained_data_delayed_106__1_, chained_data_delayed_106__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_107__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_106__127_, chained_data_delayed_106__126_, chained_data_delayed_106__125_, chained_data_delayed_106__124_, chained_data_delayed_106__123_, chained_data_delayed_106__122_, chained_data_delayed_106__121_, chained_data_delayed_106__120_, chained_data_delayed_106__119_, chained_data_delayed_106__118_, chained_data_delayed_106__117_, chained_data_delayed_106__116_, chained_data_delayed_106__115_, chained_data_delayed_106__114_, chained_data_delayed_106__113_, chained_data_delayed_106__112_, chained_data_delayed_106__111_, chained_data_delayed_106__110_, chained_data_delayed_106__109_, chained_data_delayed_106__108_, chained_data_delayed_106__107_, chained_data_delayed_106__106_, chained_data_delayed_106__105_, chained_data_delayed_106__104_, chained_data_delayed_106__103_, chained_data_delayed_106__102_, chained_data_delayed_106__101_, chained_data_delayed_106__100_, chained_data_delayed_106__99_, chained_data_delayed_106__98_, chained_data_delayed_106__97_, chained_data_delayed_106__96_, chained_data_delayed_106__95_, chained_data_delayed_106__94_, chained_data_delayed_106__93_, chained_data_delayed_106__92_, chained_data_delayed_106__91_, chained_data_delayed_106__90_, chained_data_delayed_106__89_, chained_data_delayed_106__88_, chained_data_delayed_106__87_, chained_data_delayed_106__86_, chained_data_delayed_106__85_, chained_data_delayed_106__84_, chained_data_delayed_106__83_, chained_data_delayed_106__82_, chained_data_delayed_106__81_, chained_data_delayed_106__80_, chained_data_delayed_106__79_, chained_data_delayed_106__78_, chained_data_delayed_106__77_, chained_data_delayed_106__76_, chained_data_delayed_106__75_, chained_data_delayed_106__74_, chained_data_delayed_106__73_, chained_data_delayed_106__72_, chained_data_delayed_106__71_, chained_data_delayed_106__70_, chained_data_delayed_106__69_, chained_data_delayed_106__68_, chained_data_delayed_106__67_, chained_data_delayed_106__66_, chained_data_delayed_106__65_, chained_data_delayed_106__64_, chained_data_delayed_106__63_, chained_data_delayed_106__62_, chained_data_delayed_106__61_, chained_data_delayed_106__60_, chained_data_delayed_106__59_, chained_data_delayed_106__58_, chained_data_delayed_106__57_, chained_data_delayed_106__56_, chained_data_delayed_106__55_, chained_data_delayed_106__54_, chained_data_delayed_106__53_, chained_data_delayed_106__52_, chained_data_delayed_106__51_, chained_data_delayed_106__50_, chained_data_delayed_106__49_, chained_data_delayed_106__48_, chained_data_delayed_106__47_, chained_data_delayed_106__46_, chained_data_delayed_106__45_, chained_data_delayed_106__44_, chained_data_delayed_106__43_, chained_data_delayed_106__42_, chained_data_delayed_106__41_, chained_data_delayed_106__40_, chained_data_delayed_106__39_, chained_data_delayed_106__38_, chained_data_delayed_106__37_, chained_data_delayed_106__36_, chained_data_delayed_106__35_, chained_data_delayed_106__34_, chained_data_delayed_106__33_, chained_data_delayed_106__32_, chained_data_delayed_106__31_, chained_data_delayed_106__30_, chained_data_delayed_106__29_, chained_data_delayed_106__28_, chained_data_delayed_106__27_, chained_data_delayed_106__26_, chained_data_delayed_106__25_, chained_data_delayed_106__24_, chained_data_delayed_106__23_, chained_data_delayed_106__22_, chained_data_delayed_106__21_, chained_data_delayed_106__20_, chained_data_delayed_106__19_, chained_data_delayed_106__18_, chained_data_delayed_106__17_, chained_data_delayed_106__16_, chained_data_delayed_106__15_, chained_data_delayed_106__14_, chained_data_delayed_106__13_, chained_data_delayed_106__12_, chained_data_delayed_106__11_, chained_data_delayed_106__10_, chained_data_delayed_106__9_, chained_data_delayed_106__8_, chained_data_delayed_106__7_, chained_data_delayed_106__6_, chained_data_delayed_106__5_, chained_data_delayed_106__4_, chained_data_delayed_106__3_, chained_data_delayed_106__2_, chained_data_delayed_106__1_, chained_data_delayed_106__0_ }),
    .data_o({ chained_data_delayed_107__127_, chained_data_delayed_107__126_, chained_data_delayed_107__125_, chained_data_delayed_107__124_, chained_data_delayed_107__123_, chained_data_delayed_107__122_, chained_data_delayed_107__121_, chained_data_delayed_107__120_, chained_data_delayed_107__119_, chained_data_delayed_107__118_, chained_data_delayed_107__117_, chained_data_delayed_107__116_, chained_data_delayed_107__115_, chained_data_delayed_107__114_, chained_data_delayed_107__113_, chained_data_delayed_107__112_, chained_data_delayed_107__111_, chained_data_delayed_107__110_, chained_data_delayed_107__109_, chained_data_delayed_107__108_, chained_data_delayed_107__107_, chained_data_delayed_107__106_, chained_data_delayed_107__105_, chained_data_delayed_107__104_, chained_data_delayed_107__103_, chained_data_delayed_107__102_, chained_data_delayed_107__101_, chained_data_delayed_107__100_, chained_data_delayed_107__99_, chained_data_delayed_107__98_, chained_data_delayed_107__97_, chained_data_delayed_107__96_, chained_data_delayed_107__95_, chained_data_delayed_107__94_, chained_data_delayed_107__93_, chained_data_delayed_107__92_, chained_data_delayed_107__91_, chained_data_delayed_107__90_, chained_data_delayed_107__89_, chained_data_delayed_107__88_, chained_data_delayed_107__87_, chained_data_delayed_107__86_, chained_data_delayed_107__85_, chained_data_delayed_107__84_, chained_data_delayed_107__83_, chained_data_delayed_107__82_, chained_data_delayed_107__81_, chained_data_delayed_107__80_, chained_data_delayed_107__79_, chained_data_delayed_107__78_, chained_data_delayed_107__77_, chained_data_delayed_107__76_, chained_data_delayed_107__75_, chained_data_delayed_107__74_, chained_data_delayed_107__73_, chained_data_delayed_107__72_, chained_data_delayed_107__71_, chained_data_delayed_107__70_, chained_data_delayed_107__69_, chained_data_delayed_107__68_, chained_data_delayed_107__67_, chained_data_delayed_107__66_, chained_data_delayed_107__65_, chained_data_delayed_107__64_, chained_data_delayed_107__63_, chained_data_delayed_107__62_, chained_data_delayed_107__61_, chained_data_delayed_107__60_, chained_data_delayed_107__59_, chained_data_delayed_107__58_, chained_data_delayed_107__57_, chained_data_delayed_107__56_, chained_data_delayed_107__55_, chained_data_delayed_107__54_, chained_data_delayed_107__53_, chained_data_delayed_107__52_, chained_data_delayed_107__51_, chained_data_delayed_107__50_, chained_data_delayed_107__49_, chained_data_delayed_107__48_, chained_data_delayed_107__47_, chained_data_delayed_107__46_, chained_data_delayed_107__45_, chained_data_delayed_107__44_, chained_data_delayed_107__43_, chained_data_delayed_107__42_, chained_data_delayed_107__41_, chained_data_delayed_107__40_, chained_data_delayed_107__39_, chained_data_delayed_107__38_, chained_data_delayed_107__37_, chained_data_delayed_107__36_, chained_data_delayed_107__35_, chained_data_delayed_107__34_, chained_data_delayed_107__33_, chained_data_delayed_107__32_, chained_data_delayed_107__31_, chained_data_delayed_107__30_, chained_data_delayed_107__29_, chained_data_delayed_107__28_, chained_data_delayed_107__27_, chained_data_delayed_107__26_, chained_data_delayed_107__25_, chained_data_delayed_107__24_, chained_data_delayed_107__23_, chained_data_delayed_107__22_, chained_data_delayed_107__21_, chained_data_delayed_107__20_, chained_data_delayed_107__19_, chained_data_delayed_107__18_, chained_data_delayed_107__17_, chained_data_delayed_107__16_, chained_data_delayed_107__15_, chained_data_delayed_107__14_, chained_data_delayed_107__13_, chained_data_delayed_107__12_, chained_data_delayed_107__11_, chained_data_delayed_107__10_, chained_data_delayed_107__9_, chained_data_delayed_107__8_, chained_data_delayed_107__7_, chained_data_delayed_107__6_, chained_data_delayed_107__5_, chained_data_delayed_107__4_, chained_data_delayed_107__3_, chained_data_delayed_107__2_, chained_data_delayed_107__1_, chained_data_delayed_107__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_108__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_107__127_, chained_data_delayed_107__126_, chained_data_delayed_107__125_, chained_data_delayed_107__124_, chained_data_delayed_107__123_, chained_data_delayed_107__122_, chained_data_delayed_107__121_, chained_data_delayed_107__120_, chained_data_delayed_107__119_, chained_data_delayed_107__118_, chained_data_delayed_107__117_, chained_data_delayed_107__116_, chained_data_delayed_107__115_, chained_data_delayed_107__114_, chained_data_delayed_107__113_, chained_data_delayed_107__112_, chained_data_delayed_107__111_, chained_data_delayed_107__110_, chained_data_delayed_107__109_, chained_data_delayed_107__108_, chained_data_delayed_107__107_, chained_data_delayed_107__106_, chained_data_delayed_107__105_, chained_data_delayed_107__104_, chained_data_delayed_107__103_, chained_data_delayed_107__102_, chained_data_delayed_107__101_, chained_data_delayed_107__100_, chained_data_delayed_107__99_, chained_data_delayed_107__98_, chained_data_delayed_107__97_, chained_data_delayed_107__96_, chained_data_delayed_107__95_, chained_data_delayed_107__94_, chained_data_delayed_107__93_, chained_data_delayed_107__92_, chained_data_delayed_107__91_, chained_data_delayed_107__90_, chained_data_delayed_107__89_, chained_data_delayed_107__88_, chained_data_delayed_107__87_, chained_data_delayed_107__86_, chained_data_delayed_107__85_, chained_data_delayed_107__84_, chained_data_delayed_107__83_, chained_data_delayed_107__82_, chained_data_delayed_107__81_, chained_data_delayed_107__80_, chained_data_delayed_107__79_, chained_data_delayed_107__78_, chained_data_delayed_107__77_, chained_data_delayed_107__76_, chained_data_delayed_107__75_, chained_data_delayed_107__74_, chained_data_delayed_107__73_, chained_data_delayed_107__72_, chained_data_delayed_107__71_, chained_data_delayed_107__70_, chained_data_delayed_107__69_, chained_data_delayed_107__68_, chained_data_delayed_107__67_, chained_data_delayed_107__66_, chained_data_delayed_107__65_, chained_data_delayed_107__64_, chained_data_delayed_107__63_, chained_data_delayed_107__62_, chained_data_delayed_107__61_, chained_data_delayed_107__60_, chained_data_delayed_107__59_, chained_data_delayed_107__58_, chained_data_delayed_107__57_, chained_data_delayed_107__56_, chained_data_delayed_107__55_, chained_data_delayed_107__54_, chained_data_delayed_107__53_, chained_data_delayed_107__52_, chained_data_delayed_107__51_, chained_data_delayed_107__50_, chained_data_delayed_107__49_, chained_data_delayed_107__48_, chained_data_delayed_107__47_, chained_data_delayed_107__46_, chained_data_delayed_107__45_, chained_data_delayed_107__44_, chained_data_delayed_107__43_, chained_data_delayed_107__42_, chained_data_delayed_107__41_, chained_data_delayed_107__40_, chained_data_delayed_107__39_, chained_data_delayed_107__38_, chained_data_delayed_107__37_, chained_data_delayed_107__36_, chained_data_delayed_107__35_, chained_data_delayed_107__34_, chained_data_delayed_107__33_, chained_data_delayed_107__32_, chained_data_delayed_107__31_, chained_data_delayed_107__30_, chained_data_delayed_107__29_, chained_data_delayed_107__28_, chained_data_delayed_107__27_, chained_data_delayed_107__26_, chained_data_delayed_107__25_, chained_data_delayed_107__24_, chained_data_delayed_107__23_, chained_data_delayed_107__22_, chained_data_delayed_107__21_, chained_data_delayed_107__20_, chained_data_delayed_107__19_, chained_data_delayed_107__18_, chained_data_delayed_107__17_, chained_data_delayed_107__16_, chained_data_delayed_107__15_, chained_data_delayed_107__14_, chained_data_delayed_107__13_, chained_data_delayed_107__12_, chained_data_delayed_107__11_, chained_data_delayed_107__10_, chained_data_delayed_107__9_, chained_data_delayed_107__8_, chained_data_delayed_107__7_, chained_data_delayed_107__6_, chained_data_delayed_107__5_, chained_data_delayed_107__4_, chained_data_delayed_107__3_, chained_data_delayed_107__2_, chained_data_delayed_107__1_, chained_data_delayed_107__0_ }),
    .data_o({ chained_data_delayed_108__127_, chained_data_delayed_108__126_, chained_data_delayed_108__125_, chained_data_delayed_108__124_, chained_data_delayed_108__123_, chained_data_delayed_108__122_, chained_data_delayed_108__121_, chained_data_delayed_108__120_, chained_data_delayed_108__119_, chained_data_delayed_108__118_, chained_data_delayed_108__117_, chained_data_delayed_108__116_, chained_data_delayed_108__115_, chained_data_delayed_108__114_, chained_data_delayed_108__113_, chained_data_delayed_108__112_, chained_data_delayed_108__111_, chained_data_delayed_108__110_, chained_data_delayed_108__109_, chained_data_delayed_108__108_, chained_data_delayed_108__107_, chained_data_delayed_108__106_, chained_data_delayed_108__105_, chained_data_delayed_108__104_, chained_data_delayed_108__103_, chained_data_delayed_108__102_, chained_data_delayed_108__101_, chained_data_delayed_108__100_, chained_data_delayed_108__99_, chained_data_delayed_108__98_, chained_data_delayed_108__97_, chained_data_delayed_108__96_, chained_data_delayed_108__95_, chained_data_delayed_108__94_, chained_data_delayed_108__93_, chained_data_delayed_108__92_, chained_data_delayed_108__91_, chained_data_delayed_108__90_, chained_data_delayed_108__89_, chained_data_delayed_108__88_, chained_data_delayed_108__87_, chained_data_delayed_108__86_, chained_data_delayed_108__85_, chained_data_delayed_108__84_, chained_data_delayed_108__83_, chained_data_delayed_108__82_, chained_data_delayed_108__81_, chained_data_delayed_108__80_, chained_data_delayed_108__79_, chained_data_delayed_108__78_, chained_data_delayed_108__77_, chained_data_delayed_108__76_, chained_data_delayed_108__75_, chained_data_delayed_108__74_, chained_data_delayed_108__73_, chained_data_delayed_108__72_, chained_data_delayed_108__71_, chained_data_delayed_108__70_, chained_data_delayed_108__69_, chained_data_delayed_108__68_, chained_data_delayed_108__67_, chained_data_delayed_108__66_, chained_data_delayed_108__65_, chained_data_delayed_108__64_, chained_data_delayed_108__63_, chained_data_delayed_108__62_, chained_data_delayed_108__61_, chained_data_delayed_108__60_, chained_data_delayed_108__59_, chained_data_delayed_108__58_, chained_data_delayed_108__57_, chained_data_delayed_108__56_, chained_data_delayed_108__55_, chained_data_delayed_108__54_, chained_data_delayed_108__53_, chained_data_delayed_108__52_, chained_data_delayed_108__51_, chained_data_delayed_108__50_, chained_data_delayed_108__49_, chained_data_delayed_108__48_, chained_data_delayed_108__47_, chained_data_delayed_108__46_, chained_data_delayed_108__45_, chained_data_delayed_108__44_, chained_data_delayed_108__43_, chained_data_delayed_108__42_, chained_data_delayed_108__41_, chained_data_delayed_108__40_, chained_data_delayed_108__39_, chained_data_delayed_108__38_, chained_data_delayed_108__37_, chained_data_delayed_108__36_, chained_data_delayed_108__35_, chained_data_delayed_108__34_, chained_data_delayed_108__33_, chained_data_delayed_108__32_, chained_data_delayed_108__31_, chained_data_delayed_108__30_, chained_data_delayed_108__29_, chained_data_delayed_108__28_, chained_data_delayed_108__27_, chained_data_delayed_108__26_, chained_data_delayed_108__25_, chained_data_delayed_108__24_, chained_data_delayed_108__23_, chained_data_delayed_108__22_, chained_data_delayed_108__21_, chained_data_delayed_108__20_, chained_data_delayed_108__19_, chained_data_delayed_108__18_, chained_data_delayed_108__17_, chained_data_delayed_108__16_, chained_data_delayed_108__15_, chained_data_delayed_108__14_, chained_data_delayed_108__13_, chained_data_delayed_108__12_, chained_data_delayed_108__11_, chained_data_delayed_108__10_, chained_data_delayed_108__9_, chained_data_delayed_108__8_, chained_data_delayed_108__7_, chained_data_delayed_108__6_, chained_data_delayed_108__5_, chained_data_delayed_108__4_, chained_data_delayed_108__3_, chained_data_delayed_108__2_, chained_data_delayed_108__1_, chained_data_delayed_108__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_109__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_108__127_, chained_data_delayed_108__126_, chained_data_delayed_108__125_, chained_data_delayed_108__124_, chained_data_delayed_108__123_, chained_data_delayed_108__122_, chained_data_delayed_108__121_, chained_data_delayed_108__120_, chained_data_delayed_108__119_, chained_data_delayed_108__118_, chained_data_delayed_108__117_, chained_data_delayed_108__116_, chained_data_delayed_108__115_, chained_data_delayed_108__114_, chained_data_delayed_108__113_, chained_data_delayed_108__112_, chained_data_delayed_108__111_, chained_data_delayed_108__110_, chained_data_delayed_108__109_, chained_data_delayed_108__108_, chained_data_delayed_108__107_, chained_data_delayed_108__106_, chained_data_delayed_108__105_, chained_data_delayed_108__104_, chained_data_delayed_108__103_, chained_data_delayed_108__102_, chained_data_delayed_108__101_, chained_data_delayed_108__100_, chained_data_delayed_108__99_, chained_data_delayed_108__98_, chained_data_delayed_108__97_, chained_data_delayed_108__96_, chained_data_delayed_108__95_, chained_data_delayed_108__94_, chained_data_delayed_108__93_, chained_data_delayed_108__92_, chained_data_delayed_108__91_, chained_data_delayed_108__90_, chained_data_delayed_108__89_, chained_data_delayed_108__88_, chained_data_delayed_108__87_, chained_data_delayed_108__86_, chained_data_delayed_108__85_, chained_data_delayed_108__84_, chained_data_delayed_108__83_, chained_data_delayed_108__82_, chained_data_delayed_108__81_, chained_data_delayed_108__80_, chained_data_delayed_108__79_, chained_data_delayed_108__78_, chained_data_delayed_108__77_, chained_data_delayed_108__76_, chained_data_delayed_108__75_, chained_data_delayed_108__74_, chained_data_delayed_108__73_, chained_data_delayed_108__72_, chained_data_delayed_108__71_, chained_data_delayed_108__70_, chained_data_delayed_108__69_, chained_data_delayed_108__68_, chained_data_delayed_108__67_, chained_data_delayed_108__66_, chained_data_delayed_108__65_, chained_data_delayed_108__64_, chained_data_delayed_108__63_, chained_data_delayed_108__62_, chained_data_delayed_108__61_, chained_data_delayed_108__60_, chained_data_delayed_108__59_, chained_data_delayed_108__58_, chained_data_delayed_108__57_, chained_data_delayed_108__56_, chained_data_delayed_108__55_, chained_data_delayed_108__54_, chained_data_delayed_108__53_, chained_data_delayed_108__52_, chained_data_delayed_108__51_, chained_data_delayed_108__50_, chained_data_delayed_108__49_, chained_data_delayed_108__48_, chained_data_delayed_108__47_, chained_data_delayed_108__46_, chained_data_delayed_108__45_, chained_data_delayed_108__44_, chained_data_delayed_108__43_, chained_data_delayed_108__42_, chained_data_delayed_108__41_, chained_data_delayed_108__40_, chained_data_delayed_108__39_, chained_data_delayed_108__38_, chained_data_delayed_108__37_, chained_data_delayed_108__36_, chained_data_delayed_108__35_, chained_data_delayed_108__34_, chained_data_delayed_108__33_, chained_data_delayed_108__32_, chained_data_delayed_108__31_, chained_data_delayed_108__30_, chained_data_delayed_108__29_, chained_data_delayed_108__28_, chained_data_delayed_108__27_, chained_data_delayed_108__26_, chained_data_delayed_108__25_, chained_data_delayed_108__24_, chained_data_delayed_108__23_, chained_data_delayed_108__22_, chained_data_delayed_108__21_, chained_data_delayed_108__20_, chained_data_delayed_108__19_, chained_data_delayed_108__18_, chained_data_delayed_108__17_, chained_data_delayed_108__16_, chained_data_delayed_108__15_, chained_data_delayed_108__14_, chained_data_delayed_108__13_, chained_data_delayed_108__12_, chained_data_delayed_108__11_, chained_data_delayed_108__10_, chained_data_delayed_108__9_, chained_data_delayed_108__8_, chained_data_delayed_108__7_, chained_data_delayed_108__6_, chained_data_delayed_108__5_, chained_data_delayed_108__4_, chained_data_delayed_108__3_, chained_data_delayed_108__2_, chained_data_delayed_108__1_, chained_data_delayed_108__0_ }),
    .data_o({ chained_data_delayed_109__127_, chained_data_delayed_109__126_, chained_data_delayed_109__125_, chained_data_delayed_109__124_, chained_data_delayed_109__123_, chained_data_delayed_109__122_, chained_data_delayed_109__121_, chained_data_delayed_109__120_, chained_data_delayed_109__119_, chained_data_delayed_109__118_, chained_data_delayed_109__117_, chained_data_delayed_109__116_, chained_data_delayed_109__115_, chained_data_delayed_109__114_, chained_data_delayed_109__113_, chained_data_delayed_109__112_, chained_data_delayed_109__111_, chained_data_delayed_109__110_, chained_data_delayed_109__109_, chained_data_delayed_109__108_, chained_data_delayed_109__107_, chained_data_delayed_109__106_, chained_data_delayed_109__105_, chained_data_delayed_109__104_, chained_data_delayed_109__103_, chained_data_delayed_109__102_, chained_data_delayed_109__101_, chained_data_delayed_109__100_, chained_data_delayed_109__99_, chained_data_delayed_109__98_, chained_data_delayed_109__97_, chained_data_delayed_109__96_, chained_data_delayed_109__95_, chained_data_delayed_109__94_, chained_data_delayed_109__93_, chained_data_delayed_109__92_, chained_data_delayed_109__91_, chained_data_delayed_109__90_, chained_data_delayed_109__89_, chained_data_delayed_109__88_, chained_data_delayed_109__87_, chained_data_delayed_109__86_, chained_data_delayed_109__85_, chained_data_delayed_109__84_, chained_data_delayed_109__83_, chained_data_delayed_109__82_, chained_data_delayed_109__81_, chained_data_delayed_109__80_, chained_data_delayed_109__79_, chained_data_delayed_109__78_, chained_data_delayed_109__77_, chained_data_delayed_109__76_, chained_data_delayed_109__75_, chained_data_delayed_109__74_, chained_data_delayed_109__73_, chained_data_delayed_109__72_, chained_data_delayed_109__71_, chained_data_delayed_109__70_, chained_data_delayed_109__69_, chained_data_delayed_109__68_, chained_data_delayed_109__67_, chained_data_delayed_109__66_, chained_data_delayed_109__65_, chained_data_delayed_109__64_, chained_data_delayed_109__63_, chained_data_delayed_109__62_, chained_data_delayed_109__61_, chained_data_delayed_109__60_, chained_data_delayed_109__59_, chained_data_delayed_109__58_, chained_data_delayed_109__57_, chained_data_delayed_109__56_, chained_data_delayed_109__55_, chained_data_delayed_109__54_, chained_data_delayed_109__53_, chained_data_delayed_109__52_, chained_data_delayed_109__51_, chained_data_delayed_109__50_, chained_data_delayed_109__49_, chained_data_delayed_109__48_, chained_data_delayed_109__47_, chained_data_delayed_109__46_, chained_data_delayed_109__45_, chained_data_delayed_109__44_, chained_data_delayed_109__43_, chained_data_delayed_109__42_, chained_data_delayed_109__41_, chained_data_delayed_109__40_, chained_data_delayed_109__39_, chained_data_delayed_109__38_, chained_data_delayed_109__37_, chained_data_delayed_109__36_, chained_data_delayed_109__35_, chained_data_delayed_109__34_, chained_data_delayed_109__33_, chained_data_delayed_109__32_, chained_data_delayed_109__31_, chained_data_delayed_109__30_, chained_data_delayed_109__29_, chained_data_delayed_109__28_, chained_data_delayed_109__27_, chained_data_delayed_109__26_, chained_data_delayed_109__25_, chained_data_delayed_109__24_, chained_data_delayed_109__23_, chained_data_delayed_109__22_, chained_data_delayed_109__21_, chained_data_delayed_109__20_, chained_data_delayed_109__19_, chained_data_delayed_109__18_, chained_data_delayed_109__17_, chained_data_delayed_109__16_, chained_data_delayed_109__15_, chained_data_delayed_109__14_, chained_data_delayed_109__13_, chained_data_delayed_109__12_, chained_data_delayed_109__11_, chained_data_delayed_109__10_, chained_data_delayed_109__9_, chained_data_delayed_109__8_, chained_data_delayed_109__7_, chained_data_delayed_109__6_, chained_data_delayed_109__5_, chained_data_delayed_109__4_, chained_data_delayed_109__3_, chained_data_delayed_109__2_, chained_data_delayed_109__1_, chained_data_delayed_109__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_110__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_109__127_, chained_data_delayed_109__126_, chained_data_delayed_109__125_, chained_data_delayed_109__124_, chained_data_delayed_109__123_, chained_data_delayed_109__122_, chained_data_delayed_109__121_, chained_data_delayed_109__120_, chained_data_delayed_109__119_, chained_data_delayed_109__118_, chained_data_delayed_109__117_, chained_data_delayed_109__116_, chained_data_delayed_109__115_, chained_data_delayed_109__114_, chained_data_delayed_109__113_, chained_data_delayed_109__112_, chained_data_delayed_109__111_, chained_data_delayed_109__110_, chained_data_delayed_109__109_, chained_data_delayed_109__108_, chained_data_delayed_109__107_, chained_data_delayed_109__106_, chained_data_delayed_109__105_, chained_data_delayed_109__104_, chained_data_delayed_109__103_, chained_data_delayed_109__102_, chained_data_delayed_109__101_, chained_data_delayed_109__100_, chained_data_delayed_109__99_, chained_data_delayed_109__98_, chained_data_delayed_109__97_, chained_data_delayed_109__96_, chained_data_delayed_109__95_, chained_data_delayed_109__94_, chained_data_delayed_109__93_, chained_data_delayed_109__92_, chained_data_delayed_109__91_, chained_data_delayed_109__90_, chained_data_delayed_109__89_, chained_data_delayed_109__88_, chained_data_delayed_109__87_, chained_data_delayed_109__86_, chained_data_delayed_109__85_, chained_data_delayed_109__84_, chained_data_delayed_109__83_, chained_data_delayed_109__82_, chained_data_delayed_109__81_, chained_data_delayed_109__80_, chained_data_delayed_109__79_, chained_data_delayed_109__78_, chained_data_delayed_109__77_, chained_data_delayed_109__76_, chained_data_delayed_109__75_, chained_data_delayed_109__74_, chained_data_delayed_109__73_, chained_data_delayed_109__72_, chained_data_delayed_109__71_, chained_data_delayed_109__70_, chained_data_delayed_109__69_, chained_data_delayed_109__68_, chained_data_delayed_109__67_, chained_data_delayed_109__66_, chained_data_delayed_109__65_, chained_data_delayed_109__64_, chained_data_delayed_109__63_, chained_data_delayed_109__62_, chained_data_delayed_109__61_, chained_data_delayed_109__60_, chained_data_delayed_109__59_, chained_data_delayed_109__58_, chained_data_delayed_109__57_, chained_data_delayed_109__56_, chained_data_delayed_109__55_, chained_data_delayed_109__54_, chained_data_delayed_109__53_, chained_data_delayed_109__52_, chained_data_delayed_109__51_, chained_data_delayed_109__50_, chained_data_delayed_109__49_, chained_data_delayed_109__48_, chained_data_delayed_109__47_, chained_data_delayed_109__46_, chained_data_delayed_109__45_, chained_data_delayed_109__44_, chained_data_delayed_109__43_, chained_data_delayed_109__42_, chained_data_delayed_109__41_, chained_data_delayed_109__40_, chained_data_delayed_109__39_, chained_data_delayed_109__38_, chained_data_delayed_109__37_, chained_data_delayed_109__36_, chained_data_delayed_109__35_, chained_data_delayed_109__34_, chained_data_delayed_109__33_, chained_data_delayed_109__32_, chained_data_delayed_109__31_, chained_data_delayed_109__30_, chained_data_delayed_109__29_, chained_data_delayed_109__28_, chained_data_delayed_109__27_, chained_data_delayed_109__26_, chained_data_delayed_109__25_, chained_data_delayed_109__24_, chained_data_delayed_109__23_, chained_data_delayed_109__22_, chained_data_delayed_109__21_, chained_data_delayed_109__20_, chained_data_delayed_109__19_, chained_data_delayed_109__18_, chained_data_delayed_109__17_, chained_data_delayed_109__16_, chained_data_delayed_109__15_, chained_data_delayed_109__14_, chained_data_delayed_109__13_, chained_data_delayed_109__12_, chained_data_delayed_109__11_, chained_data_delayed_109__10_, chained_data_delayed_109__9_, chained_data_delayed_109__8_, chained_data_delayed_109__7_, chained_data_delayed_109__6_, chained_data_delayed_109__5_, chained_data_delayed_109__4_, chained_data_delayed_109__3_, chained_data_delayed_109__2_, chained_data_delayed_109__1_, chained_data_delayed_109__0_ }),
    .data_o({ chained_data_delayed_110__127_, chained_data_delayed_110__126_, chained_data_delayed_110__125_, chained_data_delayed_110__124_, chained_data_delayed_110__123_, chained_data_delayed_110__122_, chained_data_delayed_110__121_, chained_data_delayed_110__120_, chained_data_delayed_110__119_, chained_data_delayed_110__118_, chained_data_delayed_110__117_, chained_data_delayed_110__116_, chained_data_delayed_110__115_, chained_data_delayed_110__114_, chained_data_delayed_110__113_, chained_data_delayed_110__112_, chained_data_delayed_110__111_, chained_data_delayed_110__110_, chained_data_delayed_110__109_, chained_data_delayed_110__108_, chained_data_delayed_110__107_, chained_data_delayed_110__106_, chained_data_delayed_110__105_, chained_data_delayed_110__104_, chained_data_delayed_110__103_, chained_data_delayed_110__102_, chained_data_delayed_110__101_, chained_data_delayed_110__100_, chained_data_delayed_110__99_, chained_data_delayed_110__98_, chained_data_delayed_110__97_, chained_data_delayed_110__96_, chained_data_delayed_110__95_, chained_data_delayed_110__94_, chained_data_delayed_110__93_, chained_data_delayed_110__92_, chained_data_delayed_110__91_, chained_data_delayed_110__90_, chained_data_delayed_110__89_, chained_data_delayed_110__88_, chained_data_delayed_110__87_, chained_data_delayed_110__86_, chained_data_delayed_110__85_, chained_data_delayed_110__84_, chained_data_delayed_110__83_, chained_data_delayed_110__82_, chained_data_delayed_110__81_, chained_data_delayed_110__80_, chained_data_delayed_110__79_, chained_data_delayed_110__78_, chained_data_delayed_110__77_, chained_data_delayed_110__76_, chained_data_delayed_110__75_, chained_data_delayed_110__74_, chained_data_delayed_110__73_, chained_data_delayed_110__72_, chained_data_delayed_110__71_, chained_data_delayed_110__70_, chained_data_delayed_110__69_, chained_data_delayed_110__68_, chained_data_delayed_110__67_, chained_data_delayed_110__66_, chained_data_delayed_110__65_, chained_data_delayed_110__64_, chained_data_delayed_110__63_, chained_data_delayed_110__62_, chained_data_delayed_110__61_, chained_data_delayed_110__60_, chained_data_delayed_110__59_, chained_data_delayed_110__58_, chained_data_delayed_110__57_, chained_data_delayed_110__56_, chained_data_delayed_110__55_, chained_data_delayed_110__54_, chained_data_delayed_110__53_, chained_data_delayed_110__52_, chained_data_delayed_110__51_, chained_data_delayed_110__50_, chained_data_delayed_110__49_, chained_data_delayed_110__48_, chained_data_delayed_110__47_, chained_data_delayed_110__46_, chained_data_delayed_110__45_, chained_data_delayed_110__44_, chained_data_delayed_110__43_, chained_data_delayed_110__42_, chained_data_delayed_110__41_, chained_data_delayed_110__40_, chained_data_delayed_110__39_, chained_data_delayed_110__38_, chained_data_delayed_110__37_, chained_data_delayed_110__36_, chained_data_delayed_110__35_, chained_data_delayed_110__34_, chained_data_delayed_110__33_, chained_data_delayed_110__32_, chained_data_delayed_110__31_, chained_data_delayed_110__30_, chained_data_delayed_110__29_, chained_data_delayed_110__28_, chained_data_delayed_110__27_, chained_data_delayed_110__26_, chained_data_delayed_110__25_, chained_data_delayed_110__24_, chained_data_delayed_110__23_, chained_data_delayed_110__22_, chained_data_delayed_110__21_, chained_data_delayed_110__20_, chained_data_delayed_110__19_, chained_data_delayed_110__18_, chained_data_delayed_110__17_, chained_data_delayed_110__16_, chained_data_delayed_110__15_, chained_data_delayed_110__14_, chained_data_delayed_110__13_, chained_data_delayed_110__12_, chained_data_delayed_110__11_, chained_data_delayed_110__10_, chained_data_delayed_110__9_, chained_data_delayed_110__8_, chained_data_delayed_110__7_, chained_data_delayed_110__6_, chained_data_delayed_110__5_, chained_data_delayed_110__4_, chained_data_delayed_110__3_, chained_data_delayed_110__2_, chained_data_delayed_110__1_, chained_data_delayed_110__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_111__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_110__127_, chained_data_delayed_110__126_, chained_data_delayed_110__125_, chained_data_delayed_110__124_, chained_data_delayed_110__123_, chained_data_delayed_110__122_, chained_data_delayed_110__121_, chained_data_delayed_110__120_, chained_data_delayed_110__119_, chained_data_delayed_110__118_, chained_data_delayed_110__117_, chained_data_delayed_110__116_, chained_data_delayed_110__115_, chained_data_delayed_110__114_, chained_data_delayed_110__113_, chained_data_delayed_110__112_, chained_data_delayed_110__111_, chained_data_delayed_110__110_, chained_data_delayed_110__109_, chained_data_delayed_110__108_, chained_data_delayed_110__107_, chained_data_delayed_110__106_, chained_data_delayed_110__105_, chained_data_delayed_110__104_, chained_data_delayed_110__103_, chained_data_delayed_110__102_, chained_data_delayed_110__101_, chained_data_delayed_110__100_, chained_data_delayed_110__99_, chained_data_delayed_110__98_, chained_data_delayed_110__97_, chained_data_delayed_110__96_, chained_data_delayed_110__95_, chained_data_delayed_110__94_, chained_data_delayed_110__93_, chained_data_delayed_110__92_, chained_data_delayed_110__91_, chained_data_delayed_110__90_, chained_data_delayed_110__89_, chained_data_delayed_110__88_, chained_data_delayed_110__87_, chained_data_delayed_110__86_, chained_data_delayed_110__85_, chained_data_delayed_110__84_, chained_data_delayed_110__83_, chained_data_delayed_110__82_, chained_data_delayed_110__81_, chained_data_delayed_110__80_, chained_data_delayed_110__79_, chained_data_delayed_110__78_, chained_data_delayed_110__77_, chained_data_delayed_110__76_, chained_data_delayed_110__75_, chained_data_delayed_110__74_, chained_data_delayed_110__73_, chained_data_delayed_110__72_, chained_data_delayed_110__71_, chained_data_delayed_110__70_, chained_data_delayed_110__69_, chained_data_delayed_110__68_, chained_data_delayed_110__67_, chained_data_delayed_110__66_, chained_data_delayed_110__65_, chained_data_delayed_110__64_, chained_data_delayed_110__63_, chained_data_delayed_110__62_, chained_data_delayed_110__61_, chained_data_delayed_110__60_, chained_data_delayed_110__59_, chained_data_delayed_110__58_, chained_data_delayed_110__57_, chained_data_delayed_110__56_, chained_data_delayed_110__55_, chained_data_delayed_110__54_, chained_data_delayed_110__53_, chained_data_delayed_110__52_, chained_data_delayed_110__51_, chained_data_delayed_110__50_, chained_data_delayed_110__49_, chained_data_delayed_110__48_, chained_data_delayed_110__47_, chained_data_delayed_110__46_, chained_data_delayed_110__45_, chained_data_delayed_110__44_, chained_data_delayed_110__43_, chained_data_delayed_110__42_, chained_data_delayed_110__41_, chained_data_delayed_110__40_, chained_data_delayed_110__39_, chained_data_delayed_110__38_, chained_data_delayed_110__37_, chained_data_delayed_110__36_, chained_data_delayed_110__35_, chained_data_delayed_110__34_, chained_data_delayed_110__33_, chained_data_delayed_110__32_, chained_data_delayed_110__31_, chained_data_delayed_110__30_, chained_data_delayed_110__29_, chained_data_delayed_110__28_, chained_data_delayed_110__27_, chained_data_delayed_110__26_, chained_data_delayed_110__25_, chained_data_delayed_110__24_, chained_data_delayed_110__23_, chained_data_delayed_110__22_, chained_data_delayed_110__21_, chained_data_delayed_110__20_, chained_data_delayed_110__19_, chained_data_delayed_110__18_, chained_data_delayed_110__17_, chained_data_delayed_110__16_, chained_data_delayed_110__15_, chained_data_delayed_110__14_, chained_data_delayed_110__13_, chained_data_delayed_110__12_, chained_data_delayed_110__11_, chained_data_delayed_110__10_, chained_data_delayed_110__9_, chained_data_delayed_110__8_, chained_data_delayed_110__7_, chained_data_delayed_110__6_, chained_data_delayed_110__5_, chained_data_delayed_110__4_, chained_data_delayed_110__3_, chained_data_delayed_110__2_, chained_data_delayed_110__1_, chained_data_delayed_110__0_ }),
    .data_o({ chained_data_delayed_111__127_, chained_data_delayed_111__126_, chained_data_delayed_111__125_, chained_data_delayed_111__124_, chained_data_delayed_111__123_, chained_data_delayed_111__122_, chained_data_delayed_111__121_, chained_data_delayed_111__120_, chained_data_delayed_111__119_, chained_data_delayed_111__118_, chained_data_delayed_111__117_, chained_data_delayed_111__116_, chained_data_delayed_111__115_, chained_data_delayed_111__114_, chained_data_delayed_111__113_, chained_data_delayed_111__112_, chained_data_delayed_111__111_, chained_data_delayed_111__110_, chained_data_delayed_111__109_, chained_data_delayed_111__108_, chained_data_delayed_111__107_, chained_data_delayed_111__106_, chained_data_delayed_111__105_, chained_data_delayed_111__104_, chained_data_delayed_111__103_, chained_data_delayed_111__102_, chained_data_delayed_111__101_, chained_data_delayed_111__100_, chained_data_delayed_111__99_, chained_data_delayed_111__98_, chained_data_delayed_111__97_, chained_data_delayed_111__96_, chained_data_delayed_111__95_, chained_data_delayed_111__94_, chained_data_delayed_111__93_, chained_data_delayed_111__92_, chained_data_delayed_111__91_, chained_data_delayed_111__90_, chained_data_delayed_111__89_, chained_data_delayed_111__88_, chained_data_delayed_111__87_, chained_data_delayed_111__86_, chained_data_delayed_111__85_, chained_data_delayed_111__84_, chained_data_delayed_111__83_, chained_data_delayed_111__82_, chained_data_delayed_111__81_, chained_data_delayed_111__80_, chained_data_delayed_111__79_, chained_data_delayed_111__78_, chained_data_delayed_111__77_, chained_data_delayed_111__76_, chained_data_delayed_111__75_, chained_data_delayed_111__74_, chained_data_delayed_111__73_, chained_data_delayed_111__72_, chained_data_delayed_111__71_, chained_data_delayed_111__70_, chained_data_delayed_111__69_, chained_data_delayed_111__68_, chained_data_delayed_111__67_, chained_data_delayed_111__66_, chained_data_delayed_111__65_, chained_data_delayed_111__64_, chained_data_delayed_111__63_, chained_data_delayed_111__62_, chained_data_delayed_111__61_, chained_data_delayed_111__60_, chained_data_delayed_111__59_, chained_data_delayed_111__58_, chained_data_delayed_111__57_, chained_data_delayed_111__56_, chained_data_delayed_111__55_, chained_data_delayed_111__54_, chained_data_delayed_111__53_, chained_data_delayed_111__52_, chained_data_delayed_111__51_, chained_data_delayed_111__50_, chained_data_delayed_111__49_, chained_data_delayed_111__48_, chained_data_delayed_111__47_, chained_data_delayed_111__46_, chained_data_delayed_111__45_, chained_data_delayed_111__44_, chained_data_delayed_111__43_, chained_data_delayed_111__42_, chained_data_delayed_111__41_, chained_data_delayed_111__40_, chained_data_delayed_111__39_, chained_data_delayed_111__38_, chained_data_delayed_111__37_, chained_data_delayed_111__36_, chained_data_delayed_111__35_, chained_data_delayed_111__34_, chained_data_delayed_111__33_, chained_data_delayed_111__32_, chained_data_delayed_111__31_, chained_data_delayed_111__30_, chained_data_delayed_111__29_, chained_data_delayed_111__28_, chained_data_delayed_111__27_, chained_data_delayed_111__26_, chained_data_delayed_111__25_, chained_data_delayed_111__24_, chained_data_delayed_111__23_, chained_data_delayed_111__22_, chained_data_delayed_111__21_, chained_data_delayed_111__20_, chained_data_delayed_111__19_, chained_data_delayed_111__18_, chained_data_delayed_111__17_, chained_data_delayed_111__16_, chained_data_delayed_111__15_, chained_data_delayed_111__14_, chained_data_delayed_111__13_, chained_data_delayed_111__12_, chained_data_delayed_111__11_, chained_data_delayed_111__10_, chained_data_delayed_111__9_, chained_data_delayed_111__8_, chained_data_delayed_111__7_, chained_data_delayed_111__6_, chained_data_delayed_111__5_, chained_data_delayed_111__4_, chained_data_delayed_111__3_, chained_data_delayed_111__2_, chained_data_delayed_111__1_, chained_data_delayed_111__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_112__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_111__127_, chained_data_delayed_111__126_, chained_data_delayed_111__125_, chained_data_delayed_111__124_, chained_data_delayed_111__123_, chained_data_delayed_111__122_, chained_data_delayed_111__121_, chained_data_delayed_111__120_, chained_data_delayed_111__119_, chained_data_delayed_111__118_, chained_data_delayed_111__117_, chained_data_delayed_111__116_, chained_data_delayed_111__115_, chained_data_delayed_111__114_, chained_data_delayed_111__113_, chained_data_delayed_111__112_, chained_data_delayed_111__111_, chained_data_delayed_111__110_, chained_data_delayed_111__109_, chained_data_delayed_111__108_, chained_data_delayed_111__107_, chained_data_delayed_111__106_, chained_data_delayed_111__105_, chained_data_delayed_111__104_, chained_data_delayed_111__103_, chained_data_delayed_111__102_, chained_data_delayed_111__101_, chained_data_delayed_111__100_, chained_data_delayed_111__99_, chained_data_delayed_111__98_, chained_data_delayed_111__97_, chained_data_delayed_111__96_, chained_data_delayed_111__95_, chained_data_delayed_111__94_, chained_data_delayed_111__93_, chained_data_delayed_111__92_, chained_data_delayed_111__91_, chained_data_delayed_111__90_, chained_data_delayed_111__89_, chained_data_delayed_111__88_, chained_data_delayed_111__87_, chained_data_delayed_111__86_, chained_data_delayed_111__85_, chained_data_delayed_111__84_, chained_data_delayed_111__83_, chained_data_delayed_111__82_, chained_data_delayed_111__81_, chained_data_delayed_111__80_, chained_data_delayed_111__79_, chained_data_delayed_111__78_, chained_data_delayed_111__77_, chained_data_delayed_111__76_, chained_data_delayed_111__75_, chained_data_delayed_111__74_, chained_data_delayed_111__73_, chained_data_delayed_111__72_, chained_data_delayed_111__71_, chained_data_delayed_111__70_, chained_data_delayed_111__69_, chained_data_delayed_111__68_, chained_data_delayed_111__67_, chained_data_delayed_111__66_, chained_data_delayed_111__65_, chained_data_delayed_111__64_, chained_data_delayed_111__63_, chained_data_delayed_111__62_, chained_data_delayed_111__61_, chained_data_delayed_111__60_, chained_data_delayed_111__59_, chained_data_delayed_111__58_, chained_data_delayed_111__57_, chained_data_delayed_111__56_, chained_data_delayed_111__55_, chained_data_delayed_111__54_, chained_data_delayed_111__53_, chained_data_delayed_111__52_, chained_data_delayed_111__51_, chained_data_delayed_111__50_, chained_data_delayed_111__49_, chained_data_delayed_111__48_, chained_data_delayed_111__47_, chained_data_delayed_111__46_, chained_data_delayed_111__45_, chained_data_delayed_111__44_, chained_data_delayed_111__43_, chained_data_delayed_111__42_, chained_data_delayed_111__41_, chained_data_delayed_111__40_, chained_data_delayed_111__39_, chained_data_delayed_111__38_, chained_data_delayed_111__37_, chained_data_delayed_111__36_, chained_data_delayed_111__35_, chained_data_delayed_111__34_, chained_data_delayed_111__33_, chained_data_delayed_111__32_, chained_data_delayed_111__31_, chained_data_delayed_111__30_, chained_data_delayed_111__29_, chained_data_delayed_111__28_, chained_data_delayed_111__27_, chained_data_delayed_111__26_, chained_data_delayed_111__25_, chained_data_delayed_111__24_, chained_data_delayed_111__23_, chained_data_delayed_111__22_, chained_data_delayed_111__21_, chained_data_delayed_111__20_, chained_data_delayed_111__19_, chained_data_delayed_111__18_, chained_data_delayed_111__17_, chained_data_delayed_111__16_, chained_data_delayed_111__15_, chained_data_delayed_111__14_, chained_data_delayed_111__13_, chained_data_delayed_111__12_, chained_data_delayed_111__11_, chained_data_delayed_111__10_, chained_data_delayed_111__9_, chained_data_delayed_111__8_, chained_data_delayed_111__7_, chained_data_delayed_111__6_, chained_data_delayed_111__5_, chained_data_delayed_111__4_, chained_data_delayed_111__3_, chained_data_delayed_111__2_, chained_data_delayed_111__1_, chained_data_delayed_111__0_ }),
    .data_o({ chained_data_delayed_112__127_, chained_data_delayed_112__126_, chained_data_delayed_112__125_, chained_data_delayed_112__124_, chained_data_delayed_112__123_, chained_data_delayed_112__122_, chained_data_delayed_112__121_, chained_data_delayed_112__120_, chained_data_delayed_112__119_, chained_data_delayed_112__118_, chained_data_delayed_112__117_, chained_data_delayed_112__116_, chained_data_delayed_112__115_, chained_data_delayed_112__114_, chained_data_delayed_112__113_, chained_data_delayed_112__112_, chained_data_delayed_112__111_, chained_data_delayed_112__110_, chained_data_delayed_112__109_, chained_data_delayed_112__108_, chained_data_delayed_112__107_, chained_data_delayed_112__106_, chained_data_delayed_112__105_, chained_data_delayed_112__104_, chained_data_delayed_112__103_, chained_data_delayed_112__102_, chained_data_delayed_112__101_, chained_data_delayed_112__100_, chained_data_delayed_112__99_, chained_data_delayed_112__98_, chained_data_delayed_112__97_, chained_data_delayed_112__96_, chained_data_delayed_112__95_, chained_data_delayed_112__94_, chained_data_delayed_112__93_, chained_data_delayed_112__92_, chained_data_delayed_112__91_, chained_data_delayed_112__90_, chained_data_delayed_112__89_, chained_data_delayed_112__88_, chained_data_delayed_112__87_, chained_data_delayed_112__86_, chained_data_delayed_112__85_, chained_data_delayed_112__84_, chained_data_delayed_112__83_, chained_data_delayed_112__82_, chained_data_delayed_112__81_, chained_data_delayed_112__80_, chained_data_delayed_112__79_, chained_data_delayed_112__78_, chained_data_delayed_112__77_, chained_data_delayed_112__76_, chained_data_delayed_112__75_, chained_data_delayed_112__74_, chained_data_delayed_112__73_, chained_data_delayed_112__72_, chained_data_delayed_112__71_, chained_data_delayed_112__70_, chained_data_delayed_112__69_, chained_data_delayed_112__68_, chained_data_delayed_112__67_, chained_data_delayed_112__66_, chained_data_delayed_112__65_, chained_data_delayed_112__64_, chained_data_delayed_112__63_, chained_data_delayed_112__62_, chained_data_delayed_112__61_, chained_data_delayed_112__60_, chained_data_delayed_112__59_, chained_data_delayed_112__58_, chained_data_delayed_112__57_, chained_data_delayed_112__56_, chained_data_delayed_112__55_, chained_data_delayed_112__54_, chained_data_delayed_112__53_, chained_data_delayed_112__52_, chained_data_delayed_112__51_, chained_data_delayed_112__50_, chained_data_delayed_112__49_, chained_data_delayed_112__48_, chained_data_delayed_112__47_, chained_data_delayed_112__46_, chained_data_delayed_112__45_, chained_data_delayed_112__44_, chained_data_delayed_112__43_, chained_data_delayed_112__42_, chained_data_delayed_112__41_, chained_data_delayed_112__40_, chained_data_delayed_112__39_, chained_data_delayed_112__38_, chained_data_delayed_112__37_, chained_data_delayed_112__36_, chained_data_delayed_112__35_, chained_data_delayed_112__34_, chained_data_delayed_112__33_, chained_data_delayed_112__32_, chained_data_delayed_112__31_, chained_data_delayed_112__30_, chained_data_delayed_112__29_, chained_data_delayed_112__28_, chained_data_delayed_112__27_, chained_data_delayed_112__26_, chained_data_delayed_112__25_, chained_data_delayed_112__24_, chained_data_delayed_112__23_, chained_data_delayed_112__22_, chained_data_delayed_112__21_, chained_data_delayed_112__20_, chained_data_delayed_112__19_, chained_data_delayed_112__18_, chained_data_delayed_112__17_, chained_data_delayed_112__16_, chained_data_delayed_112__15_, chained_data_delayed_112__14_, chained_data_delayed_112__13_, chained_data_delayed_112__12_, chained_data_delayed_112__11_, chained_data_delayed_112__10_, chained_data_delayed_112__9_, chained_data_delayed_112__8_, chained_data_delayed_112__7_, chained_data_delayed_112__6_, chained_data_delayed_112__5_, chained_data_delayed_112__4_, chained_data_delayed_112__3_, chained_data_delayed_112__2_, chained_data_delayed_112__1_, chained_data_delayed_112__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_113__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_112__127_, chained_data_delayed_112__126_, chained_data_delayed_112__125_, chained_data_delayed_112__124_, chained_data_delayed_112__123_, chained_data_delayed_112__122_, chained_data_delayed_112__121_, chained_data_delayed_112__120_, chained_data_delayed_112__119_, chained_data_delayed_112__118_, chained_data_delayed_112__117_, chained_data_delayed_112__116_, chained_data_delayed_112__115_, chained_data_delayed_112__114_, chained_data_delayed_112__113_, chained_data_delayed_112__112_, chained_data_delayed_112__111_, chained_data_delayed_112__110_, chained_data_delayed_112__109_, chained_data_delayed_112__108_, chained_data_delayed_112__107_, chained_data_delayed_112__106_, chained_data_delayed_112__105_, chained_data_delayed_112__104_, chained_data_delayed_112__103_, chained_data_delayed_112__102_, chained_data_delayed_112__101_, chained_data_delayed_112__100_, chained_data_delayed_112__99_, chained_data_delayed_112__98_, chained_data_delayed_112__97_, chained_data_delayed_112__96_, chained_data_delayed_112__95_, chained_data_delayed_112__94_, chained_data_delayed_112__93_, chained_data_delayed_112__92_, chained_data_delayed_112__91_, chained_data_delayed_112__90_, chained_data_delayed_112__89_, chained_data_delayed_112__88_, chained_data_delayed_112__87_, chained_data_delayed_112__86_, chained_data_delayed_112__85_, chained_data_delayed_112__84_, chained_data_delayed_112__83_, chained_data_delayed_112__82_, chained_data_delayed_112__81_, chained_data_delayed_112__80_, chained_data_delayed_112__79_, chained_data_delayed_112__78_, chained_data_delayed_112__77_, chained_data_delayed_112__76_, chained_data_delayed_112__75_, chained_data_delayed_112__74_, chained_data_delayed_112__73_, chained_data_delayed_112__72_, chained_data_delayed_112__71_, chained_data_delayed_112__70_, chained_data_delayed_112__69_, chained_data_delayed_112__68_, chained_data_delayed_112__67_, chained_data_delayed_112__66_, chained_data_delayed_112__65_, chained_data_delayed_112__64_, chained_data_delayed_112__63_, chained_data_delayed_112__62_, chained_data_delayed_112__61_, chained_data_delayed_112__60_, chained_data_delayed_112__59_, chained_data_delayed_112__58_, chained_data_delayed_112__57_, chained_data_delayed_112__56_, chained_data_delayed_112__55_, chained_data_delayed_112__54_, chained_data_delayed_112__53_, chained_data_delayed_112__52_, chained_data_delayed_112__51_, chained_data_delayed_112__50_, chained_data_delayed_112__49_, chained_data_delayed_112__48_, chained_data_delayed_112__47_, chained_data_delayed_112__46_, chained_data_delayed_112__45_, chained_data_delayed_112__44_, chained_data_delayed_112__43_, chained_data_delayed_112__42_, chained_data_delayed_112__41_, chained_data_delayed_112__40_, chained_data_delayed_112__39_, chained_data_delayed_112__38_, chained_data_delayed_112__37_, chained_data_delayed_112__36_, chained_data_delayed_112__35_, chained_data_delayed_112__34_, chained_data_delayed_112__33_, chained_data_delayed_112__32_, chained_data_delayed_112__31_, chained_data_delayed_112__30_, chained_data_delayed_112__29_, chained_data_delayed_112__28_, chained_data_delayed_112__27_, chained_data_delayed_112__26_, chained_data_delayed_112__25_, chained_data_delayed_112__24_, chained_data_delayed_112__23_, chained_data_delayed_112__22_, chained_data_delayed_112__21_, chained_data_delayed_112__20_, chained_data_delayed_112__19_, chained_data_delayed_112__18_, chained_data_delayed_112__17_, chained_data_delayed_112__16_, chained_data_delayed_112__15_, chained_data_delayed_112__14_, chained_data_delayed_112__13_, chained_data_delayed_112__12_, chained_data_delayed_112__11_, chained_data_delayed_112__10_, chained_data_delayed_112__9_, chained_data_delayed_112__8_, chained_data_delayed_112__7_, chained_data_delayed_112__6_, chained_data_delayed_112__5_, chained_data_delayed_112__4_, chained_data_delayed_112__3_, chained_data_delayed_112__2_, chained_data_delayed_112__1_, chained_data_delayed_112__0_ }),
    .data_o({ chained_data_delayed_113__127_, chained_data_delayed_113__126_, chained_data_delayed_113__125_, chained_data_delayed_113__124_, chained_data_delayed_113__123_, chained_data_delayed_113__122_, chained_data_delayed_113__121_, chained_data_delayed_113__120_, chained_data_delayed_113__119_, chained_data_delayed_113__118_, chained_data_delayed_113__117_, chained_data_delayed_113__116_, chained_data_delayed_113__115_, chained_data_delayed_113__114_, chained_data_delayed_113__113_, chained_data_delayed_113__112_, chained_data_delayed_113__111_, chained_data_delayed_113__110_, chained_data_delayed_113__109_, chained_data_delayed_113__108_, chained_data_delayed_113__107_, chained_data_delayed_113__106_, chained_data_delayed_113__105_, chained_data_delayed_113__104_, chained_data_delayed_113__103_, chained_data_delayed_113__102_, chained_data_delayed_113__101_, chained_data_delayed_113__100_, chained_data_delayed_113__99_, chained_data_delayed_113__98_, chained_data_delayed_113__97_, chained_data_delayed_113__96_, chained_data_delayed_113__95_, chained_data_delayed_113__94_, chained_data_delayed_113__93_, chained_data_delayed_113__92_, chained_data_delayed_113__91_, chained_data_delayed_113__90_, chained_data_delayed_113__89_, chained_data_delayed_113__88_, chained_data_delayed_113__87_, chained_data_delayed_113__86_, chained_data_delayed_113__85_, chained_data_delayed_113__84_, chained_data_delayed_113__83_, chained_data_delayed_113__82_, chained_data_delayed_113__81_, chained_data_delayed_113__80_, chained_data_delayed_113__79_, chained_data_delayed_113__78_, chained_data_delayed_113__77_, chained_data_delayed_113__76_, chained_data_delayed_113__75_, chained_data_delayed_113__74_, chained_data_delayed_113__73_, chained_data_delayed_113__72_, chained_data_delayed_113__71_, chained_data_delayed_113__70_, chained_data_delayed_113__69_, chained_data_delayed_113__68_, chained_data_delayed_113__67_, chained_data_delayed_113__66_, chained_data_delayed_113__65_, chained_data_delayed_113__64_, chained_data_delayed_113__63_, chained_data_delayed_113__62_, chained_data_delayed_113__61_, chained_data_delayed_113__60_, chained_data_delayed_113__59_, chained_data_delayed_113__58_, chained_data_delayed_113__57_, chained_data_delayed_113__56_, chained_data_delayed_113__55_, chained_data_delayed_113__54_, chained_data_delayed_113__53_, chained_data_delayed_113__52_, chained_data_delayed_113__51_, chained_data_delayed_113__50_, chained_data_delayed_113__49_, chained_data_delayed_113__48_, chained_data_delayed_113__47_, chained_data_delayed_113__46_, chained_data_delayed_113__45_, chained_data_delayed_113__44_, chained_data_delayed_113__43_, chained_data_delayed_113__42_, chained_data_delayed_113__41_, chained_data_delayed_113__40_, chained_data_delayed_113__39_, chained_data_delayed_113__38_, chained_data_delayed_113__37_, chained_data_delayed_113__36_, chained_data_delayed_113__35_, chained_data_delayed_113__34_, chained_data_delayed_113__33_, chained_data_delayed_113__32_, chained_data_delayed_113__31_, chained_data_delayed_113__30_, chained_data_delayed_113__29_, chained_data_delayed_113__28_, chained_data_delayed_113__27_, chained_data_delayed_113__26_, chained_data_delayed_113__25_, chained_data_delayed_113__24_, chained_data_delayed_113__23_, chained_data_delayed_113__22_, chained_data_delayed_113__21_, chained_data_delayed_113__20_, chained_data_delayed_113__19_, chained_data_delayed_113__18_, chained_data_delayed_113__17_, chained_data_delayed_113__16_, chained_data_delayed_113__15_, chained_data_delayed_113__14_, chained_data_delayed_113__13_, chained_data_delayed_113__12_, chained_data_delayed_113__11_, chained_data_delayed_113__10_, chained_data_delayed_113__9_, chained_data_delayed_113__8_, chained_data_delayed_113__7_, chained_data_delayed_113__6_, chained_data_delayed_113__5_, chained_data_delayed_113__4_, chained_data_delayed_113__3_, chained_data_delayed_113__2_, chained_data_delayed_113__1_, chained_data_delayed_113__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_114__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_113__127_, chained_data_delayed_113__126_, chained_data_delayed_113__125_, chained_data_delayed_113__124_, chained_data_delayed_113__123_, chained_data_delayed_113__122_, chained_data_delayed_113__121_, chained_data_delayed_113__120_, chained_data_delayed_113__119_, chained_data_delayed_113__118_, chained_data_delayed_113__117_, chained_data_delayed_113__116_, chained_data_delayed_113__115_, chained_data_delayed_113__114_, chained_data_delayed_113__113_, chained_data_delayed_113__112_, chained_data_delayed_113__111_, chained_data_delayed_113__110_, chained_data_delayed_113__109_, chained_data_delayed_113__108_, chained_data_delayed_113__107_, chained_data_delayed_113__106_, chained_data_delayed_113__105_, chained_data_delayed_113__104_, chained_data_delayed_113__103_, chained_data_delayed_113__102_, chained_data_delayed_113__101_, chained_data_delayed_113__100_, chained_data_delayed_113__99_, chained_data_delayed_113__98_, chained_data_delayed_113__97_, chained_data_delayed_113__96_, chained_data_delayed_113__95_, chained_data_delayed_113__94_, chained_data_delayed_113__93_, chained_data_delayed_113__92_, chained_data_delayed_113__91_, chained_data_delayed_113__90_, chained_data_delayed_113__89_, chained_data_delayed_113__88_, chained_data_delayed_113__87_, chained_data_delayed_113__86_, chained_data_delayed_113__85_, chained_data_delayed_113__84_, chained_data_delayed_113__83_, chained_data_delayed_113__82_, chained_data_delayed_113__81_, chained_data_delayed_113__80_, chained_data_delayed_113__79_, chained_data_delayed_113__78_, chained_data_delayed_113__77_, chained_data_delayed_113__76_, chained_data_delayed_113__75_, chained_data_delayed_113__74_, chained_data_delayed_113__73_, chained_data_delayed_113__72_, chained_data_delayed_113__71_, chained_data_delayed_113__70_, chained_data_delayed_113__69_, chained_data_delayed_113__68_, chained_data_delayed_113__67_, chained_data_delayed_113__66_, chained_data_delayed_113__65_, chained_data_delayed_113__64_, chained_data_delayed_113__63_, chained_data_delayed_113__62_, chained_data_delayed_113__61_, chained_data_delayed_113__60_, chained_data_delayed_113__59_, chained_data_delayed_113__58_, chained_data_delayed_113__57_, chained_data_delayed_113__56_, chained_data_delayed_113__55_, chained_data_delayed_113__54_, chained_data_delayed_113__53_, chained_data_delayed_113__52_, chained_data_delayed_113__51_, chained_data_delayed_113__50_, chained_data_delayed_113__49_, chained_data_delayed_113__48_, chained_data_delayed_113__47_, chained_data_delayed_113__46_, chained_data_delayed_113__45_, chained_data_delayed_113__44_, chained_data_delayed_113__43_, chained_data_delayed_113__42_, chained_data_delayed_113__41_, chained_data_delayed_113__40_, chained_data_delayed_113__39_, chained_data_delayed_113__38_, chained_data_delayed_113__37_, chained_data_delayed_113__36_, chained_data_delayed_113__35_, chained_data_delayed_113__34_, chained_data_delayed_113__33_, chained_data_delayed_113__32_, chained_data_delayed_113__31_, chained_data_delayed_113__30_, chained_data_delayed_113__29_, chained_data_delayed_113__28_, chained_data_delayed_113__27_, chained_data_delayed_113__26_, chained_data_delayed_113__25_, chained_data_delayed_113__24_, chained_data_delayed_113__23_, chained_data_delayed_113__22_, chained_data_delayed_113__21_, chained_data_delayed_113__20_, chained_data_delayed_113__19_, chained_data_delayed_113__18_, chained_data_delayed_113__17_, chained_data_delayed_113__16_, chained_data_delayed_113__15_, chained_data_delayed_113__14_, chained_data_delayed_113__13_, chained_data_delayed_113__12_, chained_data_delayed_113__11_, chained_data_delayed_113__10_, chained_data_delayed_113__9_, chained_data_delayed_113__8_, chained_data_delayed_113__7_, chained_data_delayed_113__6_, chained_data_delayed_113__5_, chained_data_delayed_113__4_, chained_data_delayed_113__3_, chained_data_delayed_113__2_, chained_data_delayed_113__1_, chained_data_delayed_113__0_ }),
    .data_o({ chained_data_delayed_114__127_, chained_data_delayed_114__126_, chained_data_delayed_114__125_, chained_data_delayed_114__124_, chained_data_delayed_114__123_, chained_data_delayed_114__122_, chained_data_delayed_114__121_, chained_data_delayed_114__120_, chained_data_delayed_114__119_, chained_data_delayed_114__118_, chained_data_delayed_114__117_, chained_data_delayed_114__116_, chained_data_delayed_114__115_, chained_data_delayed_114__114_, chained_data_delayed_114__113_, chained_data_delayed_114__112_, chained_data_delayed_114__111_, chained_data_delayed_114__110_, chained_data_delayed_114__109_, chained_data_delayed_114__108_, chained_data_delayed_114__107_, chained_data_delayed_114__106_, chained_data_delayed_114__105_, chained_data_delayed_114__104_, chained_data_delayed_114__103_, chained_data_delayed_114__102_, chained_data_delayed_114__101_, chained_data_delayed_114__100_, chained_data_delayed_114__99_, chained_data_delayed_114__98_, chained_data_delayed_114__97_, chained_data_delayed_114__96_, chained_data_delayed_114__95_, chained_data_delayed_114__94_, chained_data_delayed_114__93_, chained_data_delayed_114__92_, chained_data_delayed_114__91_, chained_data_delayed_114__90_, chained_data_delayed_114__89_, chained_data_delayed_114__88_, chained_data_delayed_114__87_, chained_data_delayed_114__86_, chained_data_delayed_114__85_, chained_data_delayed_114__84_, chained_data_delayed_114__83_, chained_data_delayed_114__82_, chained_data_delayed_114__81_, chained_data_delayed_114__80_, chained_data_delayed_114__79_, chained_data_delayed_114__78_, chained_data_delayed_114__77_, chained_data_delayed_114__76_, chained_data_delayed_114__75_, chained_data_delayed_114__74_, chained_data_delayed_114__73_, chained_data_delayed_114__72_, chained_data_delayed_114__71_, chained_data_delayed_114__70_, chained_data_delayed_114__69_, chained_data_delayed_114__68_, chained_data_delayed_114__67_, chained_data_delayed_114__66_, chained_data_delayed_114__65_, chained_data_delayed_114__64_, chained_data_delayed_114__63_, chained_data_delayed_114__62_, chained_data_delayed_114__61_, chained_data_delayed_114__60_, chained_data_delayed_114__59_, chained_data_delayed_114__58_, chained_data_delayed_114__57_, chained_data_delayed_114__56_, chained_data_delayed_114__55_, chained_data_delayed_114__54_, chained_data_delayed_114__53_, chained_data_delayed_114__52_, chained_data_delayed_114__51_, chained_data_delayed_114__50_, chained_data_delayed_114__49_, chained_data_delayed_114__48_, chained_data_delayed_114__47_, chained_data_delayed_114__46_, chained_data_delayed_114__45_, chained_data_delayed_114__44_, chained_data_delayed_114__43_, chained_data_delayed_114__42_, chained_data_delayed_114__41_, chained_data_delayed_114__40_, chained_data_delayed_114__39_, chained_data_delayed_114__38_, chained_data_delayed_114__37_, chained_data_delayed_114__36_, chained_data_delayed_114__35_, chained_data_delayed_114__34_, chained_data_delayed_114__33_, chained_data_delayed_114__32_, chained_data_delayed_114__31_, chained_data_delayed_114__30_, chained_data_delayed_114__29_, chained_data_delayed_114__28_, chained_data_delayed_114__27_, chained_data_delayed_114__26_, chained_data_delayed_114__25_, chained_data_delayed_114__24_, chained_data_delayed_114__23_, chained_data_delayed_114__22_, chained_data_delayed_114__21_, chained_data_delayed_114__20_, chained_data_delayed_114__19_, chained_data_delayed_114__18_, chained_data_delayed_114__17_, chained_data_delayed_114__16_, chained_data_delayed_114__15_, chained_data_delayed_114__14_, chained_data_delayed_114__13_, chained_data_delayed_114__12_, chained_data_delayed_114__11_, chained_data_delayed_114__10_, chained_data_delayed_114__9_, chained_data_delayed_114__8_, chained_data_delayed_114__7_, chained_data_delayed_114__6_, chained_data_delayed_114__5_, chained_data_delayed_114__4_, chained_data_delayed_114__3_, chained_data_delayed_114__2_, chained_data_delayed_114__1_, chained_data_delayed_114__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_115__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_114__127_, chained_data_delayed_114__126_, chained_data_delayed_114__125_, chained_data_delayed_114__124_, chained_data_delayed_114__123_, chained_data_delayed_114__122_, chained_data_delayed_114__121_, chained_data_delayed_114__120_, chained_data_delayed_114__119_, chained_data_delayed_114__118_, chained_data_delayed_114__117_, chained_data_delayed_114__116_, chained_data_delayed_114__115_, chained_data_delayed_114__114_, chained_data_delayed_114__113_, chained_data_delayed_114__112_, chained_data_delayed_114__111_, chained_data_delayed_114__110_, chained_data_delayed_114__109_, chained_data_delayed_114__108_, chained_data_delayed_114__107_, chained_data_delayed_114__106_, chained_data_delayed_114__105_, chained_data_delayed_114__104_, chained_data_delayed_114__103_, chained_data_delayed_114__102_, chained_data_delayed_114__101_, chained_data_delayed_114__100_, chained_data_delayed_114__99_, chained_data_delayed_114__98_, chained_data_delayed_114__97_, chained_data_delayed_114__96_, chained_data_delayed_114__95_, chained_data_delayed_114__94_, chained_data_delayed_114__93_, chained_data_delayed_114__92_, chained_data_delayed_114__91_, chained_data_delayed_114__90_, chained_data_delayed_114__89_, chained_data_delayed_114__88_, chained_data_delayed_114__87_, chained_data_delayed_114__86_, chained_data_delayed_114__85_, chained_data_delayed_114__84_, chained_data_delayed_114__83_, chained_data_delayed_114__82_, chained_data_delayed_114__81_, chained_data_delayed_114__80_, chained_data_delayed_114__79_, chained_data_delayed_114__78_, chained_data_delayed_114__77_, chained_data_delayed_114__76_, chained_data_delayed_114__75_, chained_data_delayed_114__74_, chained_data_delayed_114__73_, chained_data_delayed_114__72_, chained_data_delayed_114__71_, chained_data_delayed_114__70_, chained_data_delayed_114__69_, chained_data_delayed_114__68_, chained_data_delayed_114__67_, chained_data_delayed_114__66_, chained_data_delayed_114__65_, chained_data_delayed_114__64_, chained_data_delayed_114__63_, chained_data_delayed_114__62_, chained_data_delayed_114__61_, chained_data_delayed_114__60_, chained_data_delayed_114__59_, chained_data_delayed_114__58_, chained_data_delayed_114__57_, chained_data_delayed_114__56_, chained_data_delayed_114__55_, chained_data_delayed_114__54_, chained_data_delayed_114__53_, chained_data_delayed_114__52_, chained_data_delayed_114__51_, chained_data_delayed_114__50_, chained_data_delayed_114__49_, chained_data_delayed_114__48_, chained_data_delayed_114__47_, chained_data_delayed_114__46_, chained_data_delayed_114__45_, chained_data_delayed_114__44_, chained_data_delayed_114__43_, chained_data_delayed_114__42_, chained_data_delayed_114__41_, chained_data_delayed_114__40_, chained_data_delayed_114__39_, chained_data_delayed_114__38_, chained_data_delayed_114__37_, chained_data_delayed_114__36_, chained_data_delayed_114__35_, chained_data_delayed_114__34_, chained_data_delayed_114__33_, chained_data_delayed_114__32_, chained_data_delayed_114__31_, chained_data_delayed_114__30_, chained_data_delayed_114__29_, chained_data_delayed_114__28_, chained_data_delayed_114__27_, chained_data_delayed_114__26_, chained_data_delayed_114__25_, chained_data_delayed_114__24_, chained_data_delayed_114__23_, chained_data_delayed_114__22_, chained_data_delayed_114__21_, chained_data_delayed_114__20_, chained_data_delayed_114__19_, chained_data_delayed_114__18_, chained_data_delayed_114__17_, chained_data_delayed_114__16_, chained_data_delayed_114__15_, chained_data_delayed_114__14_, chained_data_delayed_114__13_, chained_data_delayed_114__12_, chained_data_delayed_114__11_, chained_data_delayed_114__10_, chained_data_delayed_114__9_, chained_data_delayed_114__8_, chained_data_delayed_114__7_, chained_data_delayed_114__6_, chained_data_delayed_114__5_, chained_data_delayed_114__4_, chained_data_delayed_114__3_, chained_data_delayed_114__2_, chained_data_delayed_114__1_, chained_data_delayed_114__0_ }),
    .data_o({ chained_data_delayed_115__127_, chained_data_delayed_115__126_, chained_data_delayed_115__125_, chained_data_delayed_115__124_, chained_data_delayed_115__123_, chained_data_delayed_115__122_, chained_data_delayed_115__121_, chained_data_delayed_115__120_, chained_data_delayed_115__119_, chained_data_delayed_115__118_, chained_data_delayed_115__117_, chained_data_delayed_115__116_, chained_data_delayed_115__115_, chained_data_delayed_115__114_, chained_data_delayed_115__113_, chained_data_delayed_115__112_, chained_data_delayed_115__111_, chained_data_delayed_115__110_, chained_data_delayed_115__109_, chained_data_delayed_115__108_, chained_data_delayed_115__107_, chained_data_delayed_115__106_, chained_data_delayed_115__105_, chained_data_delayed_115__104_, chained_data_delayed_115__103_, chained_data_delayed_115__102_, chained_data_delayed_115__101_, chained_data_delayed_115__100_, chained_data_delayed_115__99_, chained_data_delayed_115__98_, chained_data_delayed_115__97_, chained_data_delayed_115__96_, chained_data_delayed_115__95_, chained_data_delayed_115__94_, chained_data_delayed_115__93_, chained_data_delayed_115__92_, chained_data_delayed_115__91_, chained_data_delayed_115__90_, chained_data_delayed_115__89_, chained_data_delayed_115__88_, chained_data_delayed_115__87_, chained_data_delayed_115__86_, chained_data_delayed_115__85_, chained_data_delayed_115__84_, chained_data_delayed_115__83_, chained_data_delayed_115__82_, chained_data_delayed_115__81_, chained_data_delayed_115__80_, chained_data_delayed_115__79_, chained_data_delayed_115__78_, chained_data_delayed_115__77_, chained_data_delayed_115__76_, chained_data_delayed_115__75_, chained_data_delayed_115__74_, chained_data_delayed_115__73_, chained_data_delayed_115__72_, chained_data_delayed_115__71_, chained_data_delayed_115__70_, chained_data_delayed_115__69_, chained_data_delayed_115__68_, chained_data_delayed_115__67_, chained_data_delayed_115__66_, chained_data_delayed_115__65_, chained_data_delayed_115__64_, chained_data_delayed_115__63_, chained_data_delayed_115__62_, chained_data_delayed_115__61_, chained_data_delayed_115__60_, chained_data_delayed_115__59_, chained_data_delayed_115__58_, chained_data_delayed_115__57_, chained_data_delayed_115__56_, chained_data_delayed_115__55_, chained_data_delayed_115__54_, chained_data_delayed_115__53_, chained_data_delayed_115__52_, chained_data_delayed_115__51_, chained_data_delayed_115__50_, chained_data_delayed_115__49_, chained_data_delayed_115__48_, chained_data_delayed_115__47_, chained_data_delayed_115__46_, chained_data_delayed_115__45_, chained_data_delayed_115__44_, chained_data_delayed_115__43_, chained_data_delayed_115__42_, chained_data_delayed_115__41_, chained_data_delayed_115__40_, chained_data_delayed_115__39_, chained_data_delayed_115__38_, chained_data_delayed_115__37_, chained_data_delayed_115__36_, chained_data_delayed_115__35_, chained_data_delayed_115__34_, chained_data_delayed_115__33_, chained_data_delayed_115__32_, chained_data_delayed_115__31_, chained_data_delayed_115__30_, chained_data_delayed_115__29_, chained_data_delayed_115__28_, chained_data_delayed_115__27_, chained_data_delayed_115__26_, chained_data_delayed_115__25_, chained_data_delayed_115__24_, chained_data_delayed_115__23_, chained_data_delayed_115__22_, chained_data_delayed_115__21_, chained_data_delayed_115__20_, chained_data_delayed_115__19_, chained_data_delayed_115__18_, chained_data_delayed_115__17_, chained_data_delayed_115__16_, chained_data_delayed_115__15_, chained_data_delayed_115__14_, chained_data_delayed_115__13_, chained_data_delayed_115__12_, chained_data_delayed_115__11_, chained_data_delayed_115__10_, chained_data_delayed_115__9_, chained_data_delayed_115__8_, chained_data_delayed_115__7_, chained_data_delayed_115__6_, chained_data_delayed_115__5_, chained_data_delayed_115__4_, chained_data_delayed_115__3_, chained_data_delayed_115__2_, chained_data_delayed_115__1_, chained_data_delayed_115__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_116__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_115__127_, chained_data_delayed_115__126_, chained_data_delayed_115__125_, chained_data_delayed_115__124_, chained_data_delayed_115__123_, chained_data_delayed_115__122_, chained_data_delayed_115__121_, chained_data_delayed_115__120_, chained_data_delayed_115__119_, chained_data_delayed_115__118_, chained_data_delayed_115__117_, chained_data_delayed_115__116_, chained_data_delayed_115__115_, chained_data_delayed_115__114_, chained_data_delayed_115__113_, chained_data_delayed_115__112_, chained_data_delayed_115__111_, chained_data_delayed_115__110_, chained_data_delayed_115__109_, chained_data_delayed_115__108_, chained_data_delayed_115__107_, chained_data_delayed_115__106_, chained_data_delayed_115__105_, chained_data_delayed_115__104_, chained_data_delayed_115__103_, chained_data_delayed_115__102_, chained_data_delayed_115__101_, chained_data_delayed_115__100_, chained_data_delayed_115__99_, chained_data_delayed_115__98_, chained_data_delayed_115__97_, chained_data_delayed_115__96_, chained_data_delayed_115__95_, chained_data_delayed_115__94_, chained_data_delayed_115__93_, chained_data_delayed_115__92_, chained_data_delayed_115__91_, chained_data_delayed_115__90_, chained_data_delayed_115__89_, chained_data_delayed_115__88_, chained_data_delayed_115__87_, chained_data_delayed_115__86_, chained_data_delayed_115__85_, chained_data_delayed_115__84_, chained_data_delayed_115__83_, chained_data_delayed_115__82_, chained_data_delayed_115__81_, chained_data_delayed_115__80_, chained_data_delayed_115__79_, chained_data_delayed_115__78_, chained_data_delayed_115__77_, chained_data_delayed_115__76_, chained_data_delayed_115__75_, chained_data_delayed_115__74_, chained_data_delayed_115__73_, chained_data_delayed_115__72_, chained_data_delayed_115__71_, chained_data_delayed_115__70_, chained_data_delayed_115__69_, chained_data_delayed_115__68_, chained_data_delayed_115__67_, chained_data_delayed_115__66_, chained_data_delayed_115__65_, chained_data_delayed_115__64_, chained_data_delayed_115__63_, chained_data_delayed_115__62_, chained_data_delayed_115__61_, chained_data_delayed_115__60_, chained_data_delayed_115__59_, chained_data_delayed_115__58_, chained_data_delayed_115__57_, chained_data_delayed_115__56_, chained_data_delayed_115__55_, chained_data_delayed_115__54_, chained_data_delayed_115__53_, chained_data_delayed_115__52_, chained_data_delayed_115__51_, chained_data_delayed_115__50_, chained_data_delayed_115__49_, chained_data_delayed_115__48_, chained_data_delayed_115__47_, chained_data_delayed_115__46_, chained_data_delayed_115__45_, chained_data_delayed_115__44_, chained_data_delayed_115__43_, chained_data_delayed_115__42_, chained_data_delayed_115__41_, chained_data_delayed_115__40_, chained_data_delayed_115__39_, chained_data_delayed_115__38_, chained_data_delayed_115__37_, chained_data_delayed_115__36_, chained_data_delayed_115__35_, chained_data_delayed_115__34_, chained_data_delayed_115__33_, chained_data_delayed_115__32_, chained_data_delayed_115__31_, chained_data_delayed_115__30_, chained_data_delayed_115__29_, chained_data_delayed_115__28_, chained_data_delayed_115__27_, chained_data_delayed_115__26_, chained_data_delayed_115__25_, chained_data_delayed_115__24_, chained_data_delayed_115__23_, chained_data_delayed_115__22_, chained_data_delayed_115__21_, chained_data_delayed_115__20_, chained_data_delayed_115__19_, chained_data_delayed_115__18_, chained_data_delayed_115__17_, chained_data_delayed_115__16_, chained_data_delayed_115__15_, chained_data_delayed_115__14_, chained_data_delayed_115__13_, chained_data_delayed_115__12_, chained_data_delayed_115__11_, chained_data_delayed_115__10_, chained_data_delayed_115__9_, chained_data_delayed_115__8_, chained_data_delayed_115__7_, chained_data_delayed_115__6_, chained_data_delayed_115__5_, chained_data_delayed_115__4_, chained_data_delayed_115__3_, chained_data_delayed_115__2_, chained_data_delayed_115__1_, chained_data_delayed_115__0_ }),
    .data_o({ chained_data_delayed_116__127_, chained_data_delayed_116__126_, chained_data_delayed_116__125_, chained_data_delayed_116__124_, chained_data_delayed_116__123_, chained_data_delayed_116__122_, chained_data_delayed_116__121_, chained_data_delayed_116__120_, chained_data_delayed_116__119_, chained_data_delayed_116__118_, chained_data_delayed_116__117_, chained_data_delayed_116__116_, chained_data_delayed_116__115_, chained_data_delayed_116__114_, chained_data_delayed_116__113_, chained_data_delayed_116__112_, chained_data_delayed_116__111_, chained_data_delayed_116__110_, chained_data_delayed_116__109_, chained_data_delayed_116__108_, chained_data_delayed_116__107_, chained_data_delayed_116__106_, chained_data_delayed_116__105_, chained_data_delayed_116__104_, chained_data_delayed_116__103_, chained_data_delayed_116__102_, chained_data_delayed_116__101_, chained_data_delayed_116__100_, chained_data_delayed_116__99_, chained_data_delayed_116__98_, chained_data_delayed_116__97_, chained_data_delayed_116__96_, chained_data_delayed_116__95_, chained_data_delayed_116__94_, chained_data_delayed_116__93_, chained_data_delayed_116__92_, chained_data_delayed_116__91_, chained_data_delayed_116__90_, chained_data_delayed_116__89_, chained_data_delayed_116__88_, chained_data_delayed_116__87_, chained_data_delayed_116__86_, chained_data_delayed_116__85_, chained_data_delayed_116__84_, chained_data_delayed_116__83_, chained_data_delayed_116__82_, chained_data_delayed_116__81_, chained_data_delayed_116__80_, chained_data_delayed_116__79_, chained_data_delayed_116__78_, chained_data_delayed_116__77_, chained_data_delayed_116__76_, chained_data_delayed_116__75_, chained_data_delayed_116__74_, chained_data_delayed_116__73_, chained_data_delayed_116__72_, chained_data_delayed_116__71_, chained_data_delayed_116__70_, chained_data_delayed_116__69_, chained_data_delayed_116__68_, chained_data_delayed_116__67_, chained_data_delayed_116__66_, chained_data_delayed_116__65_, chained_data_delayed_116__64_, chained_data_delayed_116__63_, chained_data_delayed_116__62_, chained_data_delayed_116__61_, chained_data_delayed_116__60_, chained_data_delayed_116__59_, chained_data_delayed_116__58_, chained_data_delayed_116__57_, chained_data_delayed_116__56_, chained_data_delayed_116__55_, chained_data_delayed_116__54_, chained_data_delayed_116__53_, chained_data_delayed_116__52_, chained_data_delayed_116__51_, chained_data_delayed_116__50_, chained_data_delayed_116__49_, chained_data_delayed_116__48_, chained_data_delayed_116__47_, chained_data_delayed_116__46_, chained_data_delayed_116__45_, chained_data_delayed_116__44_, chained_data_delayed_116__43_, chained_data_delayed_116__42_, chained_data_delayed_116__41_, chained_data_delayed_116__40_, chained_data_delayed_116__39_, chained_data_delayed_116__38_, chained_data_delayed_116__37_, chained_data_delayed_116__36_, chained_data_delayed_116__35_, chained_data_delayed_116__34_, chained_data_delayed_116__33_, chained_data_delayed_116__32_, chained_data_delayed_116__31_, chained_data_delayed_116__30_, chained_data_delayed_116__29_, chained_data_delayed_116__28_, chained_data_delayed_116__27_, chained_data_delayed_116__26_, chained_data_delayed_116__25_, chained_data_delayed_116__24_, chained_data_delayed_116__23_, chained_data_delayed_116__22_, chained_data_delayed_116__21_, chained_data_delayed_116__20_, chained_data_delayed_116__19_, chained_data_delayed_116__18_, chained_data_delayed_116__17_, chained_data_delayed_116__16_, chained_data_delayed_116__15_, chained_data_delayed_116__14_, chained_data_delayed_116__13_, chained_data_delayed_116__12_, chained_data_delayed_116__11_, chained_data_delayed_116__10_, chained_data_delayed_116__9_, chained_data_delayed_116__8_, chained_data_delayed_116__7_, chained_data_delayed_116__6_, chained_data_delayed_116__5_, chained_data_delayed_116__4_, chained_data_delayed_116__3_, chained_data_delayed_116__2_, chained_data_delayed_116__1_, chained_data_delayed_116__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_117__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_116__127_, chained_data_delayed_116__126_, chained_data_delayed_116__125_, chained_data_delayed_116__124_, chained_data_delayed_116__123_, chained_data_delayed_116__122_, chained_data_delayed_116__121_, chained_data_delayed_116__120_, chained_data_delayed_116__119_, chained_data_delayed_116__118_, chained_data_delayed_116__117_, chained_data_delayed_116__116_, chained_data_delayed_116__115_, chained_data_delayed_116__114_, chained_data_delayed_116__113_, chained_data_delayed_116__112_, chained_data_delayed_116__111_, chained_data_delayed_116__110_, chained_data_delayed_116__109_, chained_data_delayed_116__108_, chained_data_delayed_116__107_, chained_data_delayed_116__106_, chained_data_delayed_116__105_, chained_data_delayed_116__104_, chained_data_delayed_116__103_, chained_data_delayed_116__102_, chained_data_delayed_116__101_, chained_data_delayed_116__100_, chained_data_delayed_116__99_, chained_data_delayed_116__98_, chained_data_delayed_116__97_, chained_data_delayed_116__96_, chained_data_delayed_116__95_, chained_data_delayed_116__94_, chained_data_delayed_116__93_, chained_data_delayed_116__92_, chained_data_delayed_116__91_, chained_data_delayed_116__90_, chained_data_delayed_116__89_, chained_data_delayed_116__88_, chained_data_delayed_116__87_, chained_data_delayed_116__86_, chained_data_delayed_116__85_, chained_data_delayed_116__84_, chained_data_delayed_116__83_, chained_data_delayed_116__82_, chained_data_delayed_116__81_, chained_data_delayed_116__80_, chained_data_delayed_116__79_, chained_data_delayed_116__78_, chained_data_delayed_116__77_, chained_data_delayed_116__76_, chained_data_delayed_116__75_, chained_data_delayed_116__74_, chained_data_delayed_116__73_, chained_data_delayed_116__72_, chained_data_delayed_116__71_, chained_data_delayed_116__70_, chained_data_delayed_116__69_, chained_data_delayed_116__68_, chained_data_delayed_116__67_, chained_data_delayed_116__66_, chained_data_delayed_116__65_, chained_data_delayed_116__64_, chained_data_delayed_116__63_, chained_data_delayed_116__62_, chained_data_delayed_116__61_, chained_data_delayed_116__60_, chained_data_delayed_116__59_, chained_data_delayed_116__58_, chained_data_delayed_116__57_, chained_data_delayed_116__56_, chained_data_delayed_116__55_, chained_data_delayed_116__54_, chained_data_delayed_116__53_, chained_data_delayed_116__52_, chained_data_delayed_116__51_, chained_data_delayed_116__50_, chained_data_delayed_116__49_, chained_data_delayed_116__48_, chained_data_delayed_116__47_, chained_data_delayed_116__46_, chained_data_delayed_116__45_, chained_data_delayed_116__44_, chained_data_delayed_116__43_, chained_data_delayed_116__42_, chained_data_delayed_116__41_, chained_data_delayed_116__40_, chained_data_delayed_116__39_, chained_data_delayed_116__38_, chained_data_delayed_116__37_, chained_data_delayed_116__36_, chained_data_delayed_116__35_, chained_data_delayed_116__34_, chained_data_delayed_116__33_, chained_data_delayed_116__32_, chained_data_delayed_116__31_, chained_data_delayed_116__30_, chained_data_delayed_116__29_, chained_data_delayed_116__28_, chained_data_delayed_116__27_, chained_data_delayed_116__26_, chained_data_delayed_116__25_, chained_data_delayed_116__24_, chained_data_delayed_116__23_, chained_data_delayed_116__22_, chained_data_delayed_116__21_, chained_data_delayed_116__20_, chained_data_delayed_116__19_, chained_data_delayed_116__18_, chained_data_delayed_116__17_, chained_data_delayed_116__16_, chained_data_delayed_116__15_, chained_data_delayed_116__14_, chained_data_delayed_116__13_, chained_data_delayed_116__12_, chained_data_delayed_116__11_, chained_data_delayed_116__10_, chained_data_delayed_116__9_, chained_data_delayed_116__8_, chained_data_delayed_116__7_, chained_data_delayed_116__6_, chained_data_delayed_116__5_, chained_data_delayed_116__4_, chained_data_delayed_116__3_, chained_data_delayed_116__2_, chained_data_delayed_116__1_, chained_data_delayed_116__0_ }),
    .data_o({ chained_data_delayed_117__127_, chained_data_delayed_117__126_, chained_data_delayed_117__125_, chained_data_delayed_117__124_, chained_data_delayed_117__123_, chained_data_delayed_117__122_, chained_data_delayed_117__121_, chained_data_delayed_117__120_, chained_data_delayed_117__119_, chained_data_delayed_117__118_, chained_data_delayed_117__117_, chained_data_delayed_117__116_, chained_data_delayed_117__115_, chained_data_delayed_117__114_, chained_data_delayed_117__113_, chained_data_delayed_117__112_, chained_data_delayed_117__111_, chained_data_delayed_117__110_, chained_data_delayed_117__109_, chained_data_delayed_117__108_, chained_data_delayed_117__107_, chained_data_delayed_117__106_, chained_data_delayed_117__105_, chained_data_delayed_117__104_, chained_data_delayed_117__103_, chained_data_delayed_117__102_, chained_data_delayed_117__101_, chained_data_delayed_117__100_, chained_data_delayed_117__99_, chained_data_delayed_117__98_, chained_data_delayed_117__97_, chained_data_delayed_117__96_, chained_data_delayed_117__95_, chained_data_delayed_117__94_, chained_data_delayed_117__93_, chained_data_delayed_117__92_, chained_data_delayed_117__91_, chained_data_delayed_117__90_, chained_data_delayed_117__89_, chained_data_delayed_117__88_, chained_data_delayed_117__87_, chained_data_delayed_117__86_, chained_data_delayed_117__85_, chained_data_delayed_117__84_, chained_data_delayed_117__83_, chained_data_delayed_117__82_, chained_data_delayed_117__81_, chained_data_delayed_117__80_, chained_data_delayed_117__79_, chained_data_delayed_117__78_, chained_data_delayed_117__77_, chained_data_delayed_117__76_, chained_data_delayed_117__75_, chained_data_delayed_117__74_, chained_data_delayed_117__73_, chained_data_delayed_117__72_, chained_data_delayed_117__71_, chained_data_delayed_117__70_, chained_data_delayed_117__69_, chained_data_delayed_117__68_, chained_data_delayed_117__67_, chained_data_delayed_117__66_, chained_data_delayed_117__65_, chained_data_delayed_117__64_, chained_data_delayed_117__63_, chained_data_delayed_117__62_, chained_data_delayed_117__61_, chained_data_delayed_117__60_, chained_data_delayed_117__59_, chained_data_delayed_117__58_, chained_data_delayed_117__57_, chained_data_delayed_117__56_, chained_data_delayed_117__55_, chained_data_delayed_117__54_, chained_data_delayed_117__53_, chained_data_delayed_117__52_, chained_data_delayed_117__51_, chained_data_delayed_117__50_, chained_data_delayed_117__49_, chained_data_delayed_117__48_, chained_data_delayed_117__47_, chained_data_delayed_117__46_, chained_data_delayed_117__45_, chained_data_delayed_117__44_, chained_data_delayed_117__43_, chained_data_delayed_117__42_, chained_data_delayed_117__41_, chained_data_delayed_117__40_, chained_data_delayed_117__39_, chained_data_delayed_117__38_, chained_data_delayed_117__37_, chained_data_delayed_117__36_, chained_data_delayed_117__35_, chained_data_delayed_117__34_, chained_data_delayed_117__33_, chained_data_delayed_117__32_, chained_data_delayed_117__31_, chained_data_delayed_117__30_, chained_data_delayed_117__29_, chained_data_delayed_117__28_, chained_data_delayed_117__27_, chained_data_delayed_117__26_, chained_data_delayed_117__25_, chained_data_delayed_117__24_, chained_data_delayed_117__23_, chained_data_delayed_117__22_, chained_data_delayed_117__21_, chained_data_delayed_117__20_, chained_data_delayed_117__19_, chained_data_delayed_117__18_, chained_data_delayed_117__17_, chained_data_delayed_117__16_, chained_data_delayed_117__15_, chained_data_delayed_117__14_, chained_data_delayed_117__13_, chained_data_delayed_117__12_, chained_data_delayed_117__11_, chained_data_delayed_117__10_, chained_data_delayed_117__9_, chained_data_delayed_117__8_, chained_data_delayed_117__7_, chained_data_delayed_117__6_, chained_data_delayed_117__5_, chained_data_delayed_117__4_, chained_data_delayed_117__3_, chained_data_delayed_117__2_, chained_data_delayed_117__1_, chained_data_delayed_117__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_118__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_117__127_, chained_data_delayed_117__126_, chained_data_delayed_117__125_, chained_data_delayed_117__124_, chained_data_delayed_117__123_, chained_data_delayed_117__122_, chained_data_delayed_117__121_, chained_data_delayed_117__120_, chained_data_delayed_117__119_, chained_data_delayed_117__118_, chained_data_delayed_117__117_, chained_data_delayed_117__116_, chained_data_delayed_117__115_, chained_data_delayed_117__114_, chained_data_delayed_117__113_, chained_data_delayed_117__112_, chained_data_delayed_117__111_, chained_data_delayed_117__110_, chained_data_delayed_117__109_, chained_data_delayed_117__108_, chained_data_delayed_117__107_, chained_data_delayed_117__106_, chained_data_delayed_117__105_, chained_data_delayed_117__104_, chained_data_delayed_117__103_, chained_data_delayed_117__102_, chained_data_delayed_117__101_, chained_data_delayed_117__100_, chained_data_delayed_117__99_, chained_data_delayed_117__98_, chained_data_delayed_117__97_, chained_data_delayed_117__96_, chained_data_delayed_117__95_, chained_data_delayed_117__94_, chained_data_delayed_117__93_, chained_data_delayed_117__92_, chained_data_delayed_117__91_, chained_data_delayed_117__90_, chained_data_delayed_117__89_, chained_data_delayed_117__88_, chained_data_delayed_117__87_, chained_data_delayed_117__86_, chained_data_delayed_117__85_, chained_data_delayed_117__84_, chained_data_delayed_117__83_, chained_data_delayed_117__82_, chained_data_delayed_117__81_, chained_data_delayed_117__80_, chained_data_delayed_117__79_, chained_data_delayed_117__78_, chained_data_delayed_117__77_, chained_data_delayed_117__76_, chained_data_delayed_117__75_, chained_data_delayed_117__74_, chained_data_delayed_117__73_, chained_data_delayed_117__72_, chained_data_delayed_117__71_, chained_data_delayed_117__70_, chained_data_delayed_117__69_, chained_data_delayed_117__68_, chained_data_delayed_117__67_, chained_data_delayed_117__66_, chained_data_delayed_117__65_, chained_data_delayed_117__64_, chained_data_delayed_117__63_, chained_data_delayed_117__62_, chained_data_delayed_117__61_, chained_data_delayed_117__60_, chained_data_delayed_117__59_, chained_data_delayed_117__58_, chained_data_delayed_117__57_, chained_data_delayed_117__56_, chained_data_delayed_117__55_, chained_data_delayed_117__54_, chained_data_delayed_117__53_, chained_data_delayed_117__52_, chained_data_delayed_117__51_, chained_data_delayed_117__50_, chained_data_delayed_117__49_, chained_data_delayed_117__48_, chained_data_delayed_117__47_, chained_data_delayed_117__46_, chained_data_delayed_117__45_, chained_data_delayed_117__44_, chained_data_delayed_117__43_, chained_data_delayed_117__42_, chained_data_delayed_117__41_, chained_data_delayed_117__40_, chained_data_delayed_117__39_, chained_data_delayed_117__38_, chained_data_delayed_117__37_, chained_data_delayed_117__36_, chained_data_delayed_117__35_, chained_data_delayed_117__34_, chained_data_delayed_117__33_, chained_data_delayed_117__32_, chained_data_delayed_117__31_, chained_data_delayed_117__30_, chained_data_delayed_117__29_, chained_data_delayed_117__28_, chained_data_delayed_117__27_, chained_data_delayed_117__26_, chained_data_delayed_117__25_, chained_data_delayed_117__24_, chained_data_delayed_117__23_, chained_data_delayed_117__22_, chained_data_delayed_117__21_, chained_data_delayed_117__20_, chained_data_delayed_117__19_, chained_data_delayed_117__18_, chained_data_delayed_117__17_, chained_data_delayed_117__16_, chained_data_delayed_117__15_, chained_data_delayed_117__14_, chained_data_delayed_117__13_, chained_data_delayed_117__12_, chained_data_delayed_117__11_, chained_data_delayed_117__10_, chained_data_delayed_117__9_, chained_data_delayed_117__8_, chained_data_delayed_117__7_, chained_data_delayed_117__6_, chained_data_delayed_117__5_, chained_data_delayed_117__4_, chained_data_delayed_117__3_, chained_data_delayed_117__2_, chained_data_delayed_117__1_, chained_data_delayed_117__0_ }),
    .data_o({ chained_data_delayed_118__127_, chained_data_delayed_118__126_, chained_data_delayed_118__125_, chained_data_delayed_118__124_, chained_data_delayed_118__123_, chained_data_delayed_118__122_, chained_data_delayed_118__121_, chained_data_delayed_118__120_, chained_data_delayed_118__119_, chained_data_delayed_118__118_, chained_data_delayed_118__117_, chained_data_delayed_118__116_, chained_data_delayed_118__115_, chained_data_delayed_118__114_, chained_data_delayed_118__113_, chained_data_delayed_118__112_, chained_data_delayed_118__111_, chained_data_delayed_118__110_, chained_data_delayed_118__109_, chained_data_delayed_118__108_, chained_data_delayed_118__107_, chained_data_delayed_118__106_, chained_data_delayed_118__105_, chained_data_delayed_118__104_, chained_data_delayed_118__103_, chained_data_delayed_118__102_, chained_data_delayed_118__101_, chained_data_delayed_118__100_, chained_data_delayed_118__99_, chained_data_delayed_118__98_, chained_data_delayed_118__97_, chained_data_delayed_118__96_, chained_data_delayed_118__95_, chained_data_delayed_118__94_, chained_data_delayed_118__93_, chained_data_delayed_118__92_, chained_data_delayed_118__91_, chained_data_delayed_118__90_, chained_data_delayed_118__89_, chained_data_delayed_118__88_, chained_data_delayed_118__87_, chained_data_delayed_118__86_, chained_data_delayed_118__85_, chained_data_delayed_118__84_, chained_data_delayed_118__83_, chained_data_delayed_118__82_, chained_data_delayed_118__81_, chained_data_delayed_118__80_, chained_data_delayed_118__79_, chained_data_delayed_118__78_, chained_data_delayed_118__77_, chained_data_delayed_118__76_, chained_data_delayed_118__75_, chained_data_delayed_118__74_, chained_data_delayed_118__73_, chained_data_delayed_118__72_, chained_data_delayed_118__71_, chained_data_delayed_118__70_, chained_data_delayed_118__69_, chained_data_delayed_118__68_, chained_data_delayed_118__67_, chained_data_delayed_118__66_, chained_data_delayed_118__65_, chained_data_delayed_118__64_, chained_data_delayed_118__63_, chained_data_delayed_118__62_, chained_data_delayed_118__61_, chained_data_delayed_118__60_, chained_data_delayed_118__59_, chained_data_delayed_118__58_, chained_data_delayed_118__57_, chained_data_delayed_118__56_, chained_data_delayed_118__55_, chained_data_delayed_118__54_, chained_data_delayed_118__53_, chained_data_delayed_118__52_, chained_data_delayed_118__51_, chained_data_delayed_118__50_, chained_data_delayed_118__49_, chained_data_delayed_118__48_, chained_data_delayed_118__47_, chained_data_delayed_118__46_, chained_data_delayed_118__45_, chained_data_delayed_118__44_, chained_data_delayed_118__43_, chained_data_delayed_118__42_, chained_data_delayed_118__41_, chained_data_delayed_118__40_, chained_data_delayed_118__39_, chained_data_delayed_118__38_, chained_data_delayed_118__37_, chained_data_delayed_118__36_, chained_data_delayed_118__35_, chained_data_delayed_118__34_, chained_data_delayed_118__33_, chained_data_delayed_118__32_, chained_data_delayed_118__31_, chained_data_delayed_118__30_, chained_data_delayed_118__29_, chained_data_delayed_118__28_, chained_data_delayed_118__27_, chained_data_delayed_118__26_, chained_data_delayed_118__25_, chained_data_delayed_118__24_, chained_data_delayed_118__23_, chained_data_delayed_118__22_, chained_data_delayed_118__21_, chained_data_delayed_118__20_, chained_data_delayed_118__19_, chained_data_delayed_118__18_, chained_data_delayed_118__17_, chained_data_delayed_118__16_, chained_data_delayed_118__15_, chained_data_delayed_118__14_, chained_data_delayed_118__13_, chained_data_delayed_118__12_, chained_data_delayed_118__11_, chained_data_delayed_118__10_, chained_data_delayed_118__9_, chained_data_delayed_118__8_, chained_data_delayed_118__7_, chained_data_delayed_118__6_, chained_data_delayed_118__5_, chained_data_delayed_118__4_, chained_data_delayed_118__3_, chained_data_delayed_118__2_, chained_data_delayed_118__1_, chained_data_delayed_118__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_119__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_118__127_, chained_data_delayed_118__126_, chained_data_delayed_118__125_, chained_data_delayed_118__124_, chained_data_delayed_118__123_, chained_data_delayed_118__122_, chained_data_delayed_118__121_, chained_data_delayed_118__120_, chained_data_delayed_118__119_, chained_data_delayed_118__118_, chained_data_delayed_118__117_, chained_data_delayed_118__116_, chained_data_delayed_118__115_, chained_data_delayed_118__114_, chained_data_delayed_118__113_, chained_data_delayed_118__112_, chained_data_delayed_118__111_, chained_data_delayed_118__110_, chained_data_delayed_118__109_, chained_data_delayed_118__108_, chained_data_delayed_118__107_, chained_data_delayed_118__106_, chained_data_delayed_118__105_, chained_data_delayed_118__104_, chained_data_delayed_118__103_, chained_data_delayed_118__102_, chained_data_delayed_118__101_, chained_data_delayed_118__100_, chained_data_delayed_118__99_, chained_data_delayed_118__98_, chained_data_delayed_118__97_, chained_data_delayed_118__96_, chained_data_delayed_118__95_, chained_data_delayed_118__94_, chained_data_delayed_118__93_, chained_data_delayed_118__92_, chained_data_delayed_118__91_, chained_data_delayed_118__90_, chained_data_delayed_118__89_, chained_data_delayed_118__88_, chained_data_delayed_118__87_, chained_data_delayed_118__86_, chained_data_delayed_118__85_, chained_data_delayed_118__84_, chained_data_delayed_118__83_, chained_data_delayed_118__82_, chained_data_delayed_118__81_, chained_data_delayed_118__80_, chained_data_delayed_118__79_, chained_data_delayed_118__78_, chained_data_delayed_118__77_, chained_data_delayed_118__76_, chained_data_delayed_118__75_, chained_data_delayed_118__74_, chained_data_delayed_118__73_, chained_data_delayed_118__72_, chained_data_delayed_118__71_, chained_data_delayed_118__70_, chained_data_delayed_118__69_, chained_data_delayed_118__68_, chained_data_delayed_118__67_, chained_data_delayed_118__66_, chained_data_delayed_118__65_, chained_data_delayed_118__64_, chained_data_delayed_118__63_, chained_data_delayed_118__62_, chained_data_delayed_118__61_, chained_data_delayed_118__60_, chained_data_delayed_118__59_, chained_data_delayed_118__58_, chained_data_delayed_118__57_, chained_data_delayed_118__56_, chained_data_delayed_118__55_, chained_data_delayed_118__54_, chained_data_delayed_118__53_, chained_data_delayed_118__52_, chained_data_delayed_118__51_, chained_data_delayed_118__50_, chained_data_delayed_118__49_, chained_data_delayed_118__48_, chained_data_delayed_118__47_, chained_data_delayed_118__46_, chained_data_delayed_118__45_, chained_data_delayed_118__44_, chained_data_delayed_118__43_, chained_data_delayed_118__42_, chained_data_delayed_118__41_, chained_data_delayed_118__40_, chained_data_delayed_118__39_, chained_data_delayed_118__38_, chained_data_delayed_118__37_, chained_data_delayed_118__36_, chained_data_delayed_118__35_, chained_data_delayed_118__34_, chained_data_delayed_118__33_, chained_data_delayed_118__32_, chained_data_delayed_118__31_, chained_data_delayed_118__30_, chained_data_delayed_118__29_, chained_data_delayed_118__28_, chained_data_delayed_118__27_, chained_data_delayed_118__26_, chained_data_delayed_118__25_, chained_data_delayed_118__24_, chained_data_delayed_118__23_, chained_data_delayed_118__22_, chained_data_delayed_118__21_, chained_data_delayed_118__20_, chained_data_delayed_118__19_, chained_data_delayed_118__18_, chained_data_delayed_118__17_, chained_data_delayed_118__16_, chained_data_delayed_118__15_, chained_data_delayed_118__14_, chained_data_delayed_118__13_, chained_data_delayed_118__12_, chained_data_delayed_118__11_, chained_data_delayed_118__10_, chained_data_delayed_118__9_, chained_data_delayed_118__8_, chained_data_delayed_118__7_, chained_data_delayed_118__6_, chained_data_delayed_118__5_, chained_data_delayed_118__4_, chained_data_delayed_118__3_, chained_data_delayed_118__2_, chained_data_delayed_118__1_, chained_data_delayed_118__0_ }),
    .data_o({ chained_data_delayed_119__127_, chained_data_delayed_119__126_, chained_data_delayed_119__125_, chained_data_delayed_119__124_, chained_data_delayed_119__123_, chained_data_delayed_119__122_, chained_data_delayed_119__121_, chained_data_delayed_119__120_, chained_data_delayed_119__119_, chained_data_delayed_119__118_, chained_data_delayed_119__117_, chained_data_delayed_119__116_, chained_data_delayed_119__115_, chained_data_delayed_119__114_, chained_data_delayed_119__113_, chained_data_delayed_119__112_, chained_data_delayed_119__111_, chained_data_delayed_119__110_, chained_data_delayed_119__109_, chained_data_delayed_119__108_, chained_data_delayed_119__107_, chained_data_delayed_119__106_, chained_data_delayed_119__105_, chained_data_delayed_119__104_, chained_data_delayed_119__103_, chained_data_delayed_119__102_, chained_data_delayed_119__101_, chained_data_delayed_119__100_, chained_data_delayed_119__99_, chained_data_delayed_119__98_, chained_data_delayed_119__97_, chained_data_delayed_119__96_, chained_data_delayed_119__95_, chained_data_delayed_119__94_, chained_data_delayed_119__93_, chained_data_delayed_119__92_, chained_data_delayed_119__91_, chained_data_delayed_119__90_, chained_data_delayed_119__89_, chained_data_delayed_119__88_, chained_data_delayed_119__87_, chained_data_delayed_119__86_, chained_data_delayed_119__85_, chained_data_delayed_119__84_, chained_data_delayed_119__83_, chained_data_delayed_119__82_, chained_data_delayed_119__81_, chained_data_delayed_119__80_, chained_data_delayed_119__79_, chained_data_delayed_119__78_, chained_data_delayed_119__77_, chained_data_delayed_119__76_, chained_data_delayed_119__75_, chained_data_delayed_119__74_, chained_data_delayed_119__73_, chained_data_delayed_119__72_, chained_data_delayed_119__71_, chained_data_delayed_119__70_, chained_data_delayed_119__69_, chained_data_delayed_119__68_, chained_data_delayed_119__67_, chained_data_delayed_119__66_, chained_data_delayed_119__65_, chained_data_delayed_119__64_, chained_data_delayed_119__63_, chained_data_delayed_119__62_, chained_data_delayed_119__61_, chained_data_delayed_119__60_, chained_data_delayed_119__59_, chained_data_delayed_119__58_, chained_data_delayed_119__57_, chained_data_delayed_119__56_, chained_data_delayed_119__55_, chained_data_delayed_119__54_, chained_data_delayed_119__53_, chained_data_delayed_119__52_, chained_data_delayed_119__51_, chained_data_delayed_119__50_, chained_data_delayed_119__49_, chained_data_delayed_119__48_, chained_data_delayed_119__47_, chained_data_delayed_119__46_, chained_data_delayed_119__45_, chained_data_delayed_119__44_, chained_data_delayed_119__43_, chained_data_delayed_119__42_, chained_data_delayed_119__41_, chained_data_delayed_119__40_, chained_data_delayed_119__39_, chained_data_delayed_119__38_, chained_data_delayed_119__37_, chained_data_delayed_119__36_, chained_data_delayed_119__35_, chained_data_delayed_119__34_, chained_data_delayed_119__33_, chained_data_delayed_119__32_, chained_data_delayed_119__31_, chained_data_delayed_119__30_, chained_data_delayed_119__29_, chained_data_delayed_119__28_, chained_data_delayed_119__27_, chained_data_delayed_119__26_, chained_data_delayed_119__25_, chained_data_delayed_119__24_, chained_data_delayed_119__23_, chained_data_delayed_119__22_, chained_data_delayed_119__21_, chained_data_delayed_119__20_, chained_data_delayed_119__19_, chained_data_delayed_119__18_, chained_data_delayed_119__17_, chained_data_delayed_119__16_, chained_data_delayed_119__15_, chained_data_delayed_119__14_, chained_data_delayed_119__13_, chained_data_delayed_119__12_, chained_data_delayed_119__11_, chained_data_delayed_119__10_, chained_data_delayed_119__9_, chained_data_delayed_119__8_, chained_data_delayed_119__7_, chained_data_delayed_119__6_, chained_data_delayed_119__5_, chained_data_delayed_119__4_, chained_data_delayed_119__3_, chained_data_delayed_119__2_, chained_data_delayed_119__1_, chained_data_delayed_119__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_120__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_119__127_, chained_data_delayed_119__126_, chained_data_delayed_119__125_, chained_data_delayed_119__124_, chained_data_delayed_119__123_, chained_data_delayed_119__122_, chained_data_delayed_119__121_, chained_data_delayed_119__120_, chained_data_delayed_119__119_, chained_data_delayed_119__118_, chained_data_delayed_119__117_, chained_data_delayed_119__116_, chained_data_delayed_119__115_, chained_data_delayed_119__114_, chained_data_delayed_119__113_, chained_data_delayed_119__112_, chained_data_delayed_119__111_, chained_data_delayed_119__110_, chained_data_delayed_119__109_, chained_data_delayed_119__108_, chained_data_delayed_119__107_, chained_data_delayed_119__106_, chained_data_delayed_119__105_, chained_data_delayed_119__104_, chained_data_delayed_119__103_, chained_data_delayed_119__102_, chained_data_delayed_119__101_, chained_data_delayed_119__100_, chained_data_delayed_119__99_, chained_data_delayed_119__98_, chained_data_delayed_119__97_, chained_data_delayed_119__96_, chained_data_delayed_119__95_, chained_data_delayed_119__94_, chained_data_delayed_119__93_, chained_data_delayed_119__92_, chained_data_delayed_119__91_, chained_data_delayed_119__90_, chained_data_delayed_119__89_, chained_data_delayed_119__88_, chained_data_delayed_119__87_, chained_data_delayed_119__86_, chained_data_delayed_119__85_, chained_data_delayed_119__84_, chained_data_delayed_119__83_, chained_data_delayed_119__82_, chained_data_delayed_119__81_, chained_data_delayed_119__80_, chained_data_delayed_119__79_, chained_data_delayed_119__78_, chained_data_delayed_119__77_, chained_data_delayed_119__76_, chained_data_delayed_119__75_, chained_data_delayed_119__74_, chained_data_delayed_119__73_, chained_data_delayed_119__72_, chained_data_delayed_119__71_, chained_data_delayed_119__70_, chained_data_delayed_119__69_, chained_data_delayed_119__68_, chained_data_delayed_119__67_, chained_data_delayed_119__66_, chained_data_delayed_119__65_, chained_data_delayed_119__64_, chained_data_delayed_119__63_, chained_data_delayed_119__62_, chained_data_delayed_119__61_, chained_data_delayed_119__60_, chained_data_delayed_119__59_, chained_data_delayed_119__58_, chained_data_delayed_119__57_, chained_data_delayed_119__56_, chained_data_delayed_119__55_, chained_data_delayed_119__54_, chained_data_delayed_119__53_, chained_data_delayed_119__52_, chained_data_delayed_119__51_, chained_data_delayed_119__50_, chained_data_delayed_119__49_, chained_data_delayed_119__48_, chained_data_delayed_119__47_, chained_data_delayed_119__46_, chained_data_delayed_119__45_, chained_data_delayed_119__44_, chained_data_delayed_119__43_, chained_data_delayed_119__42_, chained_data_delayed_119__41_, chained_data_delayed_119__40_, chained_data_delayed_119__39_, chained_data_delayed_119__38_, chained_data_delayed_119__37_, chained_data_delayed_119__36_, chained_data_delayed_119__35_, chained_data_delayed_119__34_, chained_data_delayed_119__33_, chained_data_delayed_119__32_, chained_data_delayed_119__31_, chained_data_delayed_119__30_, chained_data_delayed_119__29_, chained_data_delayed_119__28_, chained_data_delayed_119__27_, chained_data_delayed_119__26_, chained_data_delayed_119__25_, chained_data_delayed_119__24_, chained_data_delayed_119__23_, chained_data_delayed_119__22_, chained_data_delayed_119__21_, chained_data_delayed_119__20_, chained_data_delayed_119__19_, chained_data_delayed_119__18_, chained_data_delayed_119__17_, chained_data_delayed_119__16_, chained_data_delayed_119__15_, chained_data_delayed_119__14_, chained_data_delayed_119__13_, chained_data_delayed_119__12_, chained_data_delayed_119__11_, chained_data_delayed_119__10_, chained_data_delayed_119__9_, chained_data_delayed_119__8_, chained_data_delayed_119__7_, chained_data_delayed_119__6_, chained_data_delayed_119__5_, chained_data_delayed_119__4_, chained_data_delayed_119__3_, chained_data_delayed_119__2_, chained_data_delayed_119__1_, chained_data_delayed_119__0_ }),
    .data_o({ chained_data_delayed_120__127_, chained_data_delayed_120__126_, chained_data_delayed_120__125_, chained_data_delayed_120__124_, chained_data_delayed_120__123_, chained_data_delayed_120__122_, chained_data_delayed_120__121_, chained_data_delayed_120__120_, chained_data_delayed_120__119_, chained_data_delayed_120__118_, chained_data_delayed_120__117_, chained_data_delayed_120__116_, chained_data_delayed_120__115_, chained_data_delayed_120__114_, chained_data_delayed_120__113_, chained_data_delayed_120__112_, chained_data_delayed_120__111_, chained_data_delayed_120__110_, chained_data_delayed_120__109_, chained_data_delayed_120__108_, chained_data_delayed_120__107_, chained_data_delayed_120__106_, chained_data_delayed_120__105_, chained_data_delayed_120__104_, chained_data_delayed_120__103_, chained_data_delayed_120__102_, chained_data_delayed_120__101_, chained_data_delayed_120__100_, chained_data_delayed_120__99_, chained_data_delayed_120__98_, chained_data_delayed_120__97_, chained_data_delayed_120__96_, chained_data_delayed_120__95_, chained_data_delayed_120__94_, chained_data_delayed_120__93_, chained_data_delayed_120__92_, chained_data_delayed_120__91_, chained_data_delayed_120__90_, chained_data_delayed_120__89_, chained_data_delayed_120__88_, chained_data_delayed_120__87_, chained_data_delayed_120__86_, chained_data_delayed_120__85_, chained_data_delayed_120__84_, chained_data_delayed_120__83_, chained_data_delayed_120__82_, chained_data_delayed_120__81_, chained_data_delayed_120__80_, chained_data_delayed_120__79_, chained_data_delayed_120__78_, chained_data_delayed_120__77_, chained_data_delayed_120__76_, chained_data_delayed_120__75_, chained_data_delayed_120__74_, chained_data_delayed_120__73_, chained_data_delayed_120__72_, chained_data_delayed_120__71_, chained_data_delayed_120__70_, chained_data_delayed_120__69_, chained_data_delayed_120__68_, chained_data_delayed_120__67_, chained_data_delayed_120__66_, chained_data_delayed_120__65_, chained_data_delayed_120__64_, chained_data_delayed_120__63_, chained_data_delayed_120__62_, chained_data_delayed_120__61_, chained_data_delayed_120__60_, chained_data_delayed_120__59_, chained_data_delayed_120__58_, chained_data_delayed_120__57_, chained_data_delayed_120__56_, chained_data_delayed_120__55_, chained_data_delayed_120__54_, chained_data_delayed_120__53_, chained_data_delayed_120__52_, chained_data_delayed_120__51_, chained_data_delayed_120__50_, chained_data_delayed_120__49_, chained_data_delayed_120__48_, chained_data_delayed_120__47_, chained_data_delayed_120__46_, chained_data_delayed_120__45_, chained_data_delayed_120__44_, chained_data_delayed_120__43_, chained_data_delayed_120__42_, chained_data_delayed_120__41_, chained_data_delayed_120__40_, chained_data_delayed_120__39_, chained_data_delayed_120__38_, chained_data_delayed_120__37_, chained_data_delayed_120__36_, chained_data_delayed_120__35_, chained_data_delayed_120__34_, chained_data_delayed_120__33_, chained_data_delayed_120__32_, chained_data_delayed_120__31_, chained_data_delayed_120__30_, chained_data_delayed_120__29_, chained_data_delayed_120__28_, chained_data_delayed_120__27_, chained_data_delayed_120__26_, chained_data_delayed_120__25_, chained_data_delayed_120__24_, chained_data_delayed_120__23_, chained_data_delayed_120__22_, chained_data_delayed_120__21_, chained_data_delayed_120__20_, chained_data_delayed_120__19_, chained_data_delayed_120__18_, chained_data_delayed_120__17_, chained_data_delayed_120__16_, chained_data_delayed_120__15_, chained_data_delayed_120__14_, chained_data_delayed_120__13_, chained_data_delayed_120__12_, chained_data_delayed_120__11_, chained_data_delayed_120__10_, chained_data_delayed_120__9_, chained_data_delayed_120__8_, chained_data_delayed_120__7_, chained_data_delayed_120__6_, chained_data_delayed_120__5_, chained_data_delayed_120__4_, chained_data_delayed_120__3_, chained_data_delayed_120__2_, chained_data_delayed_120__1_, chained_data_delayed_120__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_121__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_120__127_, chained_data_delayed_120__126_, chained_data_delayed_120__125_, chained_data_delayed_120__124_, chained_data_delayed_120__123_, chained_data_delayed_120__122_, chained_data_delayed_120__121_, chained_data_delayed_120__120_, chained_data_delayed_120__119_, chained_data_delayed_120__118_, chained_data_delayed_120__117_, chained_data_delayed_120__116_, chained_data_delayed_120__115_, chained_data_delayed_120__114_, chained_data_delayed_120__113_, chained_data_delayed_120__112_, chained_data_delayed_120__111_, chained_data_delayed_120__110_, chained_data_delayed_120__109_, chained_data_delayed_120__108_, chained_data_delayed_120__107_, chained_data_delayed_120__106_, chained_data_delayed_120__105_, chained_data_delayed_120__104_, chained_data_delayed_120__103_, chained_data_delayed_120__102_, chained_data_delayed_120__101_, chained_data_delayed_120__100_, chained_data_delayed_120__99_, chained_data_delayed_120__98_, chained_data_delayed_120__97_, chained_data_delayed_120__96_, chained_data_delayed_120__95_, chained_data_delayed_120__94_, chained_data_delayed_120__93_, chained_data_delayed_120__92_, chained_data_delayed_120__91_, chained_data_delayed_120__90_, chained_data_delayed_120__89_, chained_data_delayed_120__88_, chained_data_delayed_120__87_, chained_data_delayed_120__86_, chained_data_delayed_120__85_, chained_data_delayed_120__84_, chained_data_delayed_120__83_, chained_data_delayed_120__82_, chained_data_delayed_120__81_, chained_data_delayed_120__80_, chained_data_delayed_120__79_, chained_data_delayed_120__78_, chained_data_delayed_120__77_, chained_data_delayed_120__76_, chained_data_delayed_120__75_, chained_data_delayed_120__74_, chained_data_delayed_120__73_, chained_data_delayed_120__72_, chained_data_delayed_120__71_, chained_data_delayed_120__70_, chained_data_delayed_120__69_, chained_data_delayed_120__68_, chained_data_delayed_120__67_, chained_data_delayed_120__66_, chained_data_delayed_120__65_, chained_data_delayed_120__64_, chained_data_delayed_120__63_, chained_data_delayed_120__62_, chained_data_delayed_120__61_, chained_data_delayed_120__60_, chained_data_delayed_120__59_, chained_data_delayed_120__58_, chained_data_delayed_120__57_, chained_data_delayed_120__56_, chained_data_delayed_120__55_, chained_data_delayed_120__54_, chained_data_delayed_120__53_, chained_data_delayed_120__52_, chained_data_delayed_120__51_, chained_data_delayed_120__50_, chained_data_delayed_120__49_, chained_data_delayed_120__48_, chained_data_delayed_120__47_, chained_data_delayed_120__46_, chained_data_delayed_120__45_, chained_data_delayed_120__44_, chained_data_delayed_120__43_, chained_data_delayed_120__42_, chained_data_delayed_120__41_, chained_data_delayed_120__40_, chained_data_delayed_120__39_, chained_data_delayed_120__38_, chained_data_delayed_120__37_, chained_data_delayed_120__36_, chained_data_delayed_120__35_, chained_data_delayed_120__34_, chained_data_delayed_120__33_, chained_data_delayed_120__32_, chained_data_delayed_120__31_, chained_data_delayed_120__30_, chained_data_delayed_120__29_, chained_data_delayed_120__28_, chained_data_delayed_120__27_, chained_data_delayed_120__26_, chained_data_delayed_120__25_, chained_data_delayed_120__24_, chained_data_delayed_120__23_, chained_data_delayed_120__22_, chained_data_delayed_120__21_, chained_data_delayed_120__20_, chained_data_delayed_120__19_, chained_data_delayed_120__18_, chained_data_delayed_120__17_, chained_data_delayed_120__16_, chained_data_delayed_120__15_, chained_data_delayed_120__14_, chained_data_delayed_120__13_, chained_data_delayed_120__12_, chained_data_delayed_120__11_, chained_data_delayed_120__10_, chained_data_delayed_120__9_, chained_data_delayed_120__8_, chained_data_delayed_120__7_, chained_data_delayed_120__6_, chained_data_delayed_120__5_, chained_data_delayed_120__4_, chained_data_delayed_120__3_, chained_data_delayed_120__2_, chained_data_delayed_120__1_, chained_data_delayed_120__0_ }),
    .data_o({ chained_data_delayed_121__127_, chained_data_delayed_121__126_, chained_data_delayed_121__125_, chained_data_delayed_121__124_, chained_data_delayed_121__123_, chained_data_delayed_121__122_, chained_data_delayed_121__121_, chained_data_delayed_121__120_, chained_data_delayed_121__119_, chained_data_delayed_121__118_, chained_data_delayed_121__117_, chained_data_delayed_121__116_, chained_data_delayed_121__115_, chained_data_delayed_121__114_, chained_data_delayed_121__113_, chained_data_delayed_121__112_, chained_data_delayed_121__111_, chained_data_delayed_121__110_, chained_data_delayed_121__109_, chained_data_delayed_121__108_, chained_data_delayed_121__107_, chained_data_delayed_121__106_, chained_data_delayed_121__105_, chained_data_delayed_121__104_, chained_data_delayed_121__103_, chained_data_delayed_121__102_, chained_data_delayed_121__101_, chained_data_delayed_121__100_, chained_data_delayed_121__99_, chained_data_delayed_121__98_, chained_data_delayed_121__97_, chained_data_delayed_121__96_, chained_data_delayed_121__95_, chained_data_delayed_121__94_, chained_data_delayed_121__93_, chained_data_delayed_121__92_, chained_data_delayed_121__91_, chained_data_delayed_121__90_, chained_data_delayed_121__89_, chained_data_delayed_121__88_, chained_data_delayed_121__87_, chained_data_delayed_121__86_, chained_data_delayed_121__85_, chained_data_delayed_121__84_, chained_data_delayed_121__83_, chained_data_delayed_121__82_, chained_data_delayed_121__81_, chained_data_delayed_121__80_, chained_data_delayed_121__79_, chained_data_delayed_121__78_, chained_data_delayed_121__77_, chained_data_delayed_121__76_, chained_data_delayed_121__75_, chained_data_delayed_121__74_, chained_data_delayed_121__73_, chained_data_delayed_121__72_, chained_data_delayed_121__71_, chained_data_delayed_121__70_, chained_data_delayed_121__69_, chained_data_delayed_121__68_, chained_data_delayed_121__67_, chained_data_delayed_121__66_, chained_data_delayed_121__65_, chained_data_delayed_121__64_, chained_data_delayed_121__63_, chained_data_delayed_121__62_, chained_data_delayed_121__61_, chained_data_delayed_121__60_, chained_data_delayed_121__59_, chained_data_delayed_121__58_, chained_data_delayed_121__57_, chained_data_delayed_121__56_, chained_data_delayed_121__55_, chained_data_delayed_121__54_, chained_data_delayed_121__53_, chained_data_delayed_121__52_, chained_data_delayed_121__51_, chained_data_delayed_121__50_, chained_data_delayed_121__49_, chained_data_delayed_121__48_, chained_data_delayed_121__47_, chained_data_delayed_121__46_, chained_data_delayed_121__45_, chained_data_delayed_121__44_, chained_data_delayed_121__43_, chained_data_delayed_121__42_, chained_data_delayed_121__41_, chained_data_delayed_121__40_, chained_data_delayed_121__39_, chained_data_delayed_121__38_, chained_data_delayed_121__37_, chained_data_delayed_121__36_, chained_data_delayed_121__35_, chained_data_delayed_121__34_, chained_data_delayed_121__33_, chained_data_delayed_121__32_, chained_data_delayed_121__31_, chained_data_delayed_121__30_, chained_data_delayed_121__29_, chained_data_delayed_121__28_, chained_data_delayed_121__27_, chained_data_delayed_121__26_, chained_data_delayed_121__25_, chained_data_delayed_121__24_, chained_data_delayed_121__23_, chained_data_delayed_121__22_, chained_data_delayed_121__21_, chained_data_delayed_121__20_, chained_data_delayed_121__19_, chained_data_delayed_121__18_, chained_data_delayed_121__17_, chained_data_delayed_121__16_, chained_data_delayed_121__15_, chained_data_delayed_121__14_, chained_data_delayed_121__13_, chained_data_delayed_121__12_, chained_data_delayed_121__11_, chained_data_delayed_121__10_, chained_data_delayed_121__9_, chained_data_delayed_121__8_, chained_data_delayed_121__7_, chained_data_delayed_121__6_, chained_data_delayed_121__5_, chained_data_delayed_121__4_, chained_data_delayed_121__3_, chained_data_delayed_121__2_, chained_data_delayed_121__1_, chained_data_delayed_121__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_122__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_121__127_, chained_data_delayed_121__126_, chained_data_delayed_121__125_, chained_data_delayed_121__124_, chained_data_delayed_121__123_, chained_data_delayed_121__122_, chained_data_delayed_121__121_, chained_data_delayed_121__120_, chained_data_delayed_121__119_, chained_data_delayed_121__118_, chained_data_delayed_121__117_, chained_data_delayed_121__116_, chained_data_delayed_121__115_, chained_data_delayed_121__114_, chained_data_delayed_121__113_, chained_data_delayed_121__112_, chained_data_delayed_121__111_, chained_data_delayed_121__110_, chained_data_delayed_121__109_, chained_data_delayed_121__108_, chained_data_delayed_121__107_, chained_data_delayed_121__106_, chained_data_delayed_121__105_, chained_data_delayed_121__104_, chained_data_delayed_121__103_, chained_data_delayed_121__102_, chained_data_delayed_121__101_, chained_data_delayed_121__100_, chained_data_delayed_121__99_, chained_data_delayed_121__98_, chained_data_delayed_121__97_, chained_data_delayed_121__96_, chained_data_delayed_121__95_, chained_data_delayed_121__94_, chained_data_delayed_121__93_, chained_data_delayed_121__92_, chained_data_delayed_121__91_, chained_data_delayed_121__90_, chained_data_delayed_121__89_, chained_data_delayed_121__88_, chained_data_delayed_121__87_, chained_data_delayed_121__86_, chained_data_delayed_121__85_, chained_data_delayed_121__84_, chained_data_delayed_121__83_, chained_data_delayed_121__82_, chained_data_delayed_121__81_, chained_data_delayed_121__80_, chained_data_delayed_121__79_, chained_data_delayed_121__78_, chained_data_delayed_121__77_, chained_data_delayed_121__76_, chained_data_delayed_121__75_, chained_data_delayed_121__74_, chained_data_delayed_121__73_, chained_data_delayed_121__72_, chained_data_delayed_121__71_, chained_data_delayed_121__70_, chained_data_delayed_121__69_, chained_data_delayed_121__68_, chained_data_delayed_121__67_, chained_data_delayed_121__66_, chained_data_delayed_121__65_, chained_data_delayed_121__64_, chained_data_delayed_121__63_, chained_data_delayed_121__62_, chained_data_delayed_121__61_, chained_data_delayed_121__60_, chained_data_delayed_121__59_, chained_data_delayed_121__58_, chained_data_delayed_121__57_, chained_data_delayed_121__56_, chained_data_delayed_121__55_, chained_data_delayed_121__54_, chained_data_delayed_121__53_, chained_data_delayed_121__52_, chained_data_delayed_121__51_, chained_data_delayed_121__50_, chained_data_delayed_121__49_, chained_data_delayed_121__48_, chained_data_delayed_121__47_, chained_data_delayed_121__46_, chained_data_delayed_121__45_, chained_data_delayed_121__44_, chained_data_delayed_121__43_, chained_data_delayed_121__42_, chained_data_delayed_121__41_, chained_data_delayed_121__40_, chained_data_delayed_121__39_, chained_data_delayed_121__38_, chained_data_delayed_121__37_, chained_data_delayed_121__36_, chained_data_delayed_121__35_, chained_data_delayed_121__34_, chained_data_delayed_121__33_, chained_data_delayed_121__32_, chained_data_delayed_121__31_, chained_data_delayed_121__30_, chained_data_delayed_121__29_, chained_data_delayed_121__28_, chained_data_delayed_121__27_, chained_data_delayed_121__26_, chained_data_delayed_121__25_, chained_data_delayed_121__24_, chained_data_delayed_121__23_, chained_data_delayed_121__22_, chained_data_delayed_121__21_, chained_data_delayed_121__20_, chained_data_delayed_121__19_, chained_data_delayed_121__18_, chained_data_delayed_121__17_, chained_data_delayed_121__16_, chained_data_delayed_121__15_, chained_data_delayed_121__14_, chained_data_delayed_121__13_, chained_data_delayed_121__12_, chained_data_delayed_121__11_, chained_data_delayed_121__10_, chained_data_delayed_121__9_, chained_data_delayed_121__8_, chained_data_delayed_121__7_, chained_data_delayed_121__6_, chained_data_delayed_121__5_, chained_data_delayed_121__4_, chained_data_delayed_121__3_, chained_data_delayed_121__2_, chained_data_delayed_121__1_, chained_data_delayed_121__0_ }),
    .data_o({ chained_data_delayed_122__127_, chained_data_delayed_122__126_, chained_data_delayed_122__125_, chained_data_delayed_122__124_, chained_data_delayed_122__123_, chained_data_delayed_122__122_, chained_data_delayed_122__121_, chained_data_delayed_122__120_, chained_data_delayed_122__119_, chained_data_delayed_122__118_, chained_data_delayed_122__117_, chained_data_delayed_122__116_, chained_data_delayed_122__115_, chained_data_delayed_122__114_, chained_data_delayed_122__113_, chained_data_delayed_122__112_, chained_data_delayed_122__111_, chained_data_delayed_122__110_, chained_data_delayed_122__109_, chained_data_delayed_122__108_, chained_data_delayed_122__107_, chained_data_delayed_122__106_, chained_data_delayed_122__105_, chained_data_delayed_122__104_, chained_data_delayed_122__103_, chained_data_delayed_122__102_, chained_data_delayed_122__101_, chained_data_delayed_122__100_, chained_data_delayed_122__99_, chained_data_delayed_122__98_, chained_data_delayed_122__97_, chained_data_delayed_122__96_, chained_data_delayed_122__95_, chained_data_delayed_122__94_, chained_data_delayed_122__93_, chained_data_delayed_122__92_, chained_data_delayed_122__91_, chained_data_delayed_122__90_, chained_data_delayed_122__89_, chained_data_delayed_122__88_, chained_data_delayed_122__87_, chained_data_delayed_122__86_, chained_data_delayed_122__85_, chained_data_delayed_122__84_, chained_data_delayed_122__83_, chained_data_delayed_122__82_, chained_data_delayed_122__81_, chained_data_delayed_122__80_, chained_data_delayed_122__79_, chained_data_delayed_122__78_, chained_data_delayed_122__77_, chained_data_delayed_122__76_, chained_data_delayed_122__75_, chained_data_delayed_122__74_, chained_data_delayed_122__73_, chained_data_delayed_122__72_, chained_data_delayed_122__71_, chained_data_delayed_122__70_, chained_data_delayed_122__69_, chained_data_delayed_122__68_, chained_data_delayed_122__67_, chained_data_delayed_122__66_, chained_data_delayed_122__65_, chained_data_delayed_122__64_, chained_data_delayed_122__63_, chained_data_delayed_122__62_, chained_data_delayed_122__61_, chained_data_delayed_122__60_, chained_data_delayed_122__59_, chained_data_delayed_122__58_, chained_data_delayed_122__57_, chained_data_delayed_122__56_, chained_data_delayed_122__55_, chained_data_delayed_122__54_, chained_data_delayed_122__53_, chained_data_delayed_122__52_, chained_data_delayed_122__51_, chained_data_delayed_122__50_, chained_data_delayed_122__49_, chained_data_delayed_122__48_, chained_data_delayed_122__47_, chained_data_delayed_122__46_, chained_data_delayed_122__45_, chained_data_delayed_122__44_, chained_data_delayed_122__43_, chained_data_delayed_122__42_, chained_data_delayed_122__41_, chained_data_delayed_122__40_, chained_data_delayed_122__39_, chained_data_delayed_122__38_, chained_data_delayed_122__37_, chained_data_delayed_122__36_, chained_data_delayed_122__35_, chained_data_delayed_122__34_, chained_data_delayed_122__33_, chained_data_delayed_122__32_, chained_data_delayed_122__31_, chained_data_delayed_122__30_, chained_data_delayed_122__29_, chained_data_delayed_122__28_, chained_data_delayed_122__27_, chained_data_delayed_122__26_, chained_data_delayed_122__25_, chained_data_delayed_122__24_, chained_data_delayed_122__23_, chained_data_delayed_122__22_, chained_data_delayed_122__21_, chained_data_delayed_122__20_, chained_data_delayed_122__19_, chained_data_delayed_122__18_, chained_data_delayed_122__17_, chained_data_delayed_122__16_, chained_data_delayed_122__15_, chained_data_delayed_122__14_, chained_data_delayed_122__13_, chained_data_delayed_122__12_, chained_data_delayed_122__11_, chained_data_delayed_122__10_, chained_data_delayed_122__9_, chained_data_delayed_122__8_, chained_data_delayed_122__7_, chained_data_delayed_122__6_, chained_data_delayed_122__5_, chained_data_delayed_122__4_, chained_data_delayed_122__3_, chained_data_delayed_122__2_, chained_data_delayed_122__1_, chained_data_delayed_122__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_123__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_122__127_, chained_data_delayed_122__126_, chained_data_delayed_122__125_, chained_data_delayed_122__124_, chained_data_delayed_122__123_, chained_data_delayed_122__122_, chained_data_delayed_122__121_, chained_data_delayed_122__120_, chained_data_delayed_122__119_, chained_data_delayed_122__118_, chained_data_delayed_122__117_, chained_data_delayed_122__116_, chained_data_delayed_122__115_, chained_data_delayed_122__114_, chained_data_delayed_122__113_, chained_data_delayed_122__112_, chained_data_delayed_122__111_, chained_data_delayed_122__110_, chained_data_delayed_122__109_, chained_data_delayed_122__108_, chained_data_delayed_122__107_, chained_data_delayed_122__106_, chained_data_delayed_122__105_, chained_data_delayed_122__104_, chained_data_delayed_122__103_, chained_data_delayed_122__102_, chained_data_delayed_122__101_, chained_data_delayed_122__100_, chained_data_delayed_122__99_, chained_data_delayed_122__98_, chained_data_delayed_122__97_, chained_data_delayed_122__96_, chained_data_delayed_122__95_, chained_data_delayed_122__94_, chained_data_delayed_122__93_, chained_data_delayed_122__92_, chained_data_delayed_122__91_, chained_data_delayed_122__90_, chained_data_delayed_122__89_, chained_data_delayed_122__88_, chained_data_delayed_122__87_, chained_data_delayed_122__86_, chained_data_delayed_122__85_, chained_data_delayed_122__84_, chained_data_delayed_122__83_, chained_data_delayed_122__82_, chained_data_delayed_122__81_, chained_data_delayed_122__80_, chained_data_delayed_122__79_, chained_data_delayed_122__78_, chained_data_delayed_122__77_, chained_data_delayed_122__76_, chained_data_delayed_122__75_, chained_data_delayed_122__74_, chained_data_delayed_122__73_, chained_data_delayed_122__72_, chained_data_delayed_122__71_, chained_data_delayed_122__70_, chained_data_delayed_122__69_, chained_data_delayed_122__68_, chained_data_delayed_122__67_, chained_data_delayed_122__66_, chained_data_delayed_122__65_, chained_data_delayed_122__64_, chained_data_delayed_122__63_, chained_data_delayed_122__62_, chained_data_delayed_122__61_, chained_data_delayed_122__60_, chained_data_delayed_122__59_, chained_data_delayed_122__58_, chained_data_delayed_122__57_, chained_data_delayed_122__56_, chained_data_delayed_122__55_, chained_data_delayed_122__54_, chained_data_delayed_122__53_, chained_data_delayed_122__52_, chained_data_delayed_122__51_, chained_data_delayed_122__50_, chained_data_delayed_122__49_, chained_data_delayed_122__48_, chained_data_delayed_122__47_, chained_data_delayed_122__46_, chained_data_delayed_122__45_, chained_data_delayed_122__44_, chained_data_delayed_122__43_, chained_data_delayed_122__42_, chained_data_delayed_122__41_, chained_data_delayed_122__40_, chained_data_delayed_122__39_, chained_data_delayed_122__38_, chained_data_delayed_122__37_, chained_data_delayed_122__36_, chained_data_delayed_122__35_, chained_data_delayed_122__34_, chained_data_delayed_122__33_, chained_data_delayed_122__32_, chained_data_delayed_122__31_, chained_data_delayed_122__30_, chained_data_delayed_122__29_, chained_data_delayed_122__28_, chained_data_delayed_122__27_, chained_data_delayed_122__26_, chained_data_delayed_122__25_, chained_data_delayed_122__24_, chained_data_delayed_122__23_, chained_data_delayed_122__22_, chained_data_delayed_122__21_, chained_data_delayed_122__20_, chained_data_delayed_122__19_, chained_data_delayed_122__18_, chained_data_delayed_122__17_, chained_data_delayed_122__16_, chained_data_delayed_122__15_, chained_data_delayed_122__14_, chained_data_delayed_122__13_, chained_data_delayed_122__12_, chained_data_delayed_122__11_, chained_data_delayed_122__10_, chained_data_delayed_122__9_, chained_data_delayed_122__8_, chained_data_delayed_122__7_, chained_data_delayed_122__6_, chained_data_delayed_122__5_, chained_data_delayed_122__4_, chained_data_delayed_122__3_, chained_data_delayed_122__2_, chained_data_delayed_122__1_, chained_data_delayed_122__0_ }),
    .data_o({ chained_data_delayed_123__127_, chained_data_delayed_123__126_, chained_data_delayed_123__125_, chained_data_delayed_123__124_, chained_data_delayed_123__123_, chained_data_delayed_123__122_, chained_data_delayed_123__121_, chained_data_delayed_123__120_, chained_data_delayed_123__119_, chained_data_delayed_123__118_, chained_data_delayed_123__117_, chained_data_delayed_123__116_, chained_data_delayed_123__115_, chained_data_delayed_123__114_, chained_data_delayed_123__113_, chained_data_delayed_123__112_, chained_data_delayed_123__111_, chained_data_delayed_123__110_, chained_data_delayed_123__109_, chained_data_delayed_123__108_, chained_data_delayed_123__107_, chained_data_delayed_123__106_, chained_data_delayed_123__105_, chained_data_delayed_123__104_, chained_data_delayed_123__103_, chained_data_delayed_123__102_, chained_data_delayed_123__101_, chained_data_delayed_123__100_, chained_data_delayed_123__99_, chained_data_delayed_123__98_, chained_data_delayed_123__97_, chained_data_delayed_123__96_, chained_data_delayed_123__95_, chained_data_delayed_123__94_, chained_data_delayed_123__93_, chained_data_delayed_123__92_, chained_data_delayed_123__91_, chained_data_delayed_123__90_, chained_data_delayed_123__89_, chained_data_delayed_123__88_, chained_data_delayed_123__87_, chained_data_delayed_123__86_, chained_data_delayed_123__85_, chained_data_delayed_123__84_, chained_data_delayed_123__83_, chained_data_delayed_123__82_, chained_data_delayed_123__81_, chained_data_delayed_123__80_, chained_data_delayed_123__79_, chained_data_delayed_123__78_, chained_data_delayed_123__77_, chained_data_delayed_123__76_, chained_data_delayed_123__75_, chained_data_delayed_123__74_, chained_data_delayed_123__73_, chained_data_delayed_123__72_, chained_data_delayed_123__71_, chained_data_delayed_123__70_, chained_data_delayed_123__69_, chained_data_delayed_123__68_, chained_data_delayed_123__67_, chained_data_delayed_123__66_, chained_data_delayed_123__65_, chained_data_delayed_123__64_, chained_data_delayed_123__63_, chained_data_delayed_123__62_, chained_data_delayed_123__61_, chained_data_delayed_123__60_, chained_data_delayed_123__59_, chained_data_delayed_123__58_, chained_data_delayed_123__57_, chained_data_delayed_123__56_, chained_data_delayed_123__55_, chained_data_delayed_123__54_, chained_data_delayed_123__53_, chained_data_delayed_123__52_, chained_data_delayed_123__51_, chained_data_delayed_123__50_, chained_data_delayed_123__49_, chained_data_delayed_123__48_, chained_data_delayed_123__47_, chained_data_delayed_123__46_, chained_data_delayed_123__45_, chained_data_delayed_123__44_, chained_data_delayed_123__43_, chained_data_delayed_123__42_, chained_data_delayed_123__41_, chained_data_delayed_123__40_, chained_data_delayed_123__39_, chained_data_delayed_123__38_, chained_data_delayed_123__37_, chained_data_delayed_123__36_, chained_data_delayed_123__35_, chained_data_delayed_123__34_, chained_data_delayed_123__33_, chained_data_delayed_123__32_, chained_data_delayed_123__31_, chained_data_delayed_123__30_, chained_data_delayed_123__29_, chained_data_delayed_123__28_, chained_data_delayed_123__27_, chained_data_delayed_123__26_, chained_data_delayed_123__25_, chained_data_delayed_123__24_, chained_data_delayed_123__23_, chained_data_delayed_123__22_, chained_data_delayed_123__21_, chained_data_delayed_123__20_, chained_data_delayed_123__19_, chained_data_delayed_123__18_, chained_data_delayed_123__17_, chained_data_delayed_123__16_, chained_data_delayed_123__15_, chained_data_delayed_123__14_, chained_data_delayed_123__13_, chained_data_delayed_123__12_, chained_data_delayed_123__11_, chained_data_delayed_123__10_, chained_data_delayed_123__9_, chained_data_delayed_123__8_, chained_data_delayed_123__7_, chained_data_delayed_123__6_, chained_data_delayed_123__5_, chained_data_delayed_123__4_, chained_data_delayed_123__3_, chained_data_delayed_123__2_, chained_data_delayed_123__1_, chained_data_delayed_123__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_124__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_123__127_, chained_data_delayed_123__126_, chained_data_delayed_123__125_, chained_data_delayed_123__124_, chained_data_delayed_123__123_, chained_data_delayed_123__122_, chained_data_delayed_123__121_, chained_data_delayed_123__120_, chained_data_delayed_123__119_, chained_data_delayed_123__118_, chained_data_delayed_123__117_, chained_data_delayed_123__116_, chained_data_delayed_123__115_, chained_data_delayed_123__114_, chained_data_delayed_123__113_, chained_data_delayed_123__112_, chained_data_delayed_123__111_, chained_data_delayed_123__110_, chained_data_delayed_123__109_, chained_data_delayed_123__108_, chained_data_delayed_123__107_, chained_data_delayed_123__106_, chained_data_delayed_123__105_, chained_data_delayed_123__104_, chained_data_delayed_123__103_, chained_data_delayed_123__102_, chained_data_delayed_123__101_, chained_data_delayed_123__100_, chained_data_delayed_123__99_, chained_data_delayed_123__98_, chained_data_delayed_123__97_, chained_data_delayed_123__96_, chained_data_delayed_123__95_, chained_data_delayed_123__94_, chained_data_delayed_123__93_, chained_data_delayed_123__92_, chained_data_delayed_123__91_, chained_data_delayed_123__90_, chained_data_delayed_123__89_, chained_data_delayed_123__88_, chained_data_delayed_123__87_, chained_data_delayed_123__86_, chained_data_delayed_123__85_, chained_data_delayed_123__84_, chained_data_delayed_123__83_, chained_data_delayed_123__82_, chained_data_delayed_123__81_, chained_data_delayed_123__80_, chained_data_delayed_123__79_, chained_data_delayed_123__78_, chained_data_delayed_123__77_, chained_data_delayed_123__76_, chained_data_delayed_123__75_, chained_data_delayed_123__74_, chained_data_delayed_123__73_, chained_data_delayed_123__72_, chained_data_delayed_123__71_, chained_data_delayed_123__70_, chained_data_delayed_123__69_, chained_data_delayed_123__68_, chained_data_delayed_123__67_, chained_data_delayed_123__66_, chained_data_delayed_123__65_, chained_data_delayed_123__64_, chained_data_delayed_123__63_, chained_data_delayed_123__62_, chained_data_delayed_123__61_, chained_data_delayed_123__60_, chained_data_delayed_123__59_, chained_data_delayed_123__58_, chained_data_delayed_123__57_, chained_data_delayed_123__56_, chained_data_delayed_123__55_, chained_data_delayed_123__54_, chained_data_delayed_123__53_, chained_data_delayed_123__52_, chained_data_delayed_123__51_, chained_data_delayed_123__50_, chained_data_delayed_123__49_, chained_data_delayed_123__48_, chained_data_delayed_123__47_, chained_data_delayed_123__46_, chained_data_delayed_123__45_, chained_data_delayed_123__44_, chained_data_delayed_123__43_, chained_data_delayed_123__42_, chained_data_delayed_123__41_, chained_data_delayed_123__40_, chained_data_delayed_123__39_, chained_data_delayed_123__38_, chained_data_delayed_123__37_, chained_data_delayed_123__36_, chained_data_delayed_123__35_, chained_data_delayed_123__34_, chained_data_delayed_123__33_, chained_data_delayed_123__32_, chained_data_delayed_123__31_, chained_data_delayed_123__30_, chained_data_delayed_123__29_, chained_data_delayed_123__28_, chained_data_delayed_123__27_, chained_data_delayed_123__26_, chained_data_delayed_123__25_, chained_data_delayed_123__24_, chained_data_delayed_123__23_, chained_data_delayed_123__22_, chained_data_delayed_123__21_, chained_data_delayed_123__20_, chained_data_delayed_123__19_, chained_data_delayed_123__18_, chained_data_delayed_123__17_, chained_data_delayed_123__16_, chained_data_delayed_123__15_, chained_data_delayed_123__14_, chained_data_delayed_123__13_, chained_data_delayed_123__12_, chained_data_delayed_123__11_, chained_data_delayed_123__10_, chained_data_delayed_123__9_, chained_data_delayed_123__8_, chained_data_delayed_123__7_, chained_data_delayed_123__6_, chained_data_delayed_123__5_, chained_data_delayed_123__4_, chained_data_delayed_123__3_, chained_data_delayed_123__2_, chained_data_delayed_123__1_, chained_data_delayed_123__0_ }),
    .data_o({ chained_data_delayed_124__127_, chained_data_delayed_124__126_, chained_data_delayed_124__125_, chained_data_delayed_124__124_, chained_data_delayed_124__123_, chained_data_delayed_124__122_, chained_data_delayed_124__121_, chained_data_delayed_124__120_, chained_data_delayed_124__119_, chained_data_delayed_124__118_, chained_data_delayed_124__117_, chained_data_delayed_124__116_, chained_data_delayed_124__115_, chained_data_delayed_124__114_, chained_data_delayed_124__113_, chained_data_delayed_124__112_, chained_data_delayed_124__111_, chained_data_delayed_124__110_, chained_data_delayed_124__109_, chained_data_delayed_124__108_, chained_data_delayed_124__107_, chained_data_delayed_124__106_, chained_data_delayed_124__105_, chained_data_delayed_124__104_, chained_data_delayed_124__103_, chained_data_delayed_124__102_, chained_data_delayed_124__101_, chained_data_delayed_124__100_, chained_data_delayed_124__99_, chained_data_delayed_124__98_, chained_data_delayed_124__97_, chained_data_delayed_124__96_, chained_data_delayed_124__95_, chained_data_delayed_124__94_, chained_data_delayed_124__93_, chained_data_delayed_124__92_, chained_data_delayed_124__91_, chained_data_delayed_124__90_, chained_data_delayed_124__89_, chained_data_delayed_124__88_, chained_data_delayed_124__87_, chained_data_delayed_124__86_, chained_data_delayed_124__85_, chained_data_delayed_124__84_, chained_data_delayed_124__83_, chained_data_delayed_124__82_, chained_data_delayed_124__81_, chained_data_delayed_124__80_, chained_data_delayed_124__79_, chained_data_delayed_124__78_, chained_data_delayed_124__77_, chained_data_delayed_124__76_, chained_data_delayed_124__75_, chained_data_delayed_124__74_, chained_data_delayed_124__73_, chained_data_delayed_124__72_, chained_data_delayed_124__71_, chained_data_delayed_124__70_, chained_data_delayed_124__69_, chained_data_delayed_124__68_, chained_data_delayed_124__67_, chained_data_delayed_124__66_, chained_data_delayed_124__65_, chained_data_delayed_124__64_, chained_data_delayed_124__63_, chained_data_delayed_124__62_, chained_data_delayed_124__61_, chained_data_delayed_124__60_, chained_data_delayed_124__59_, chained_data_delayed_124__58_, chained_data_delayed_124__57_, chained_data_delayed_124__56_, chained_data_delayed_124__55_, chained_data_delayed_124__54_, chained_data_delayed_124__53_, chained_data_delayed_124__52_, chained_data_delayed_124__51_, chained_data_delayed_124__50_, chained_data_delayed_124__49_, chained_data_delayed_124__48_, chained_data_delayed_124__47_, chained_data_delayed_124__46_, chained_data_delayed_124__45_, chained_data_delayed_124__44_, chained_data_delayed_124__43_, chained_data_delayed_124__42_, chained_data_delayed_124__41_, chained_data_delayed_124__40_, chained_data_delayed_124__39_, chained_data_delayed_124__38_, chained_data_delayed_124__37_, chained_data_delayed_124__36_, chained_data_delayed_124__35_, chained_data_delayed_124__34_, chained_data_delayed_124__33_, chained_data_delayed_124__32_, chained_data_delayed_124__31_, chained_data_delayed_124__30_, chained_data_delayed_124__29_, chained_data_delayed_124__28_, chained_data_delayed_124__27_, chained_data_delayed_124__26_, chained_data_delayed_124__25_, chained_data_delayed_124__24_, chained_data_delayed_124__23_, chained_data_delayed_124__22_, chained_data_delayed_124__21_, chained_data_delayed_124__20_, chained_data_delayed_124__19_, chained_data_delayed_124__18_, chained_data_delayed_124__17_, chained_data_delayed_124__16_, chained_data_delayed_124__15_, chained_data_delayed_124__14_, chained_data_delayed_124__13_, chained_data_delayed_124__12_, chained_data_delayed_124__11_, chained_data_delayed_124__10_, chained_data_delayed_124__9_, chained_data_delayed_124__8_, chained_data_delayed_124__7_, chained_data_delayed_124__6_, chained_data_delayed_124__5_, chained_data_delayed_124__4_, chained_data_delayed_124__3_, chained_data_delayed_124__2_, chained_data_delayed_124__1_, chained_data_delayed_124__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_125__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_124__127_, chained_data_delayed_124__126_, chained_data_delayed_124__125_, chained_data_delayed_124__124_, chained_data_delayed_124__123_, chained_data_delayed_124__122_, chained_data_delayed_124__121_, chained_data_delayed_124__120_, chained_data_delayed_124__119_, chained_data_delayed_124__118_, chained_data_delayed_124__117_, chained_data_delayed_124__116_, chained_data_delayed_124__115_, chained_data_delayed_124__114_, chained_data_delayed_124__113_, chained_data_delayed_124__112_, chained_data_delayed_124__111_, chained_data_delayed_124__110_, chained_data_delayed_124__109_, chained_data_delayed_124__108_, chained_data_delayed_124__107_, chained_data_delayed_124__106_, chained_data_delayed_124__105_, chained_data_delayed_124__104_, chained_data_delayed_124__103_, chained_data_delayed_124__102_, chained_data_delayed_124__101_, chained_data_delayed_124__100_, chained_data_delayed_124__99_, chained_data_delayed_124__98_, chained_data_delayed_124__97_, chained_data_delayed_124__96_, chained_data_delayed_124__95_, chained_data_delayed_124__94_, chained_data_delayed_124__93_, chained_data_delayed_124__92_, chained_data_delayed_124__91_, chained_data_delayed_124__90_, chained_data_delayed_124__89_, chained_data_delayed_124__88_, chained_data_delayed_124__87_, chained_data_delayed_124__86_, chained_data_delayed_124__85_, chained_data_delayed_124__84_, chained_data_delayed_124__83_, chained_data_delayed_124__82_, chained_data_delayed_124__81_, chained_data_delayed_124__80_, chained_data_delayed_124__79_, chained_data_delayed_124__78_, chained_data_delayed_124__77_, chained_data_delayed_124__76_, chained_data_delayed_124__75_, chained_data_delayed_124__74_, chained_data_delayed_124__73_, chained_data_delayed_124__72_, chained_data_delayed_124__71_, chained_data_delayed_124__70_, chained_data_delayed_124__69_, chained_data_delayed_124__68_, chained_data_delayed_124__67_, chained_data_delayed_124__66_, chained_data_delayed_124__65_, chained_data_delayed_124__64_, chained_data_delayed_124__63_, chained_data_delayed_124__62_, chained_data_delayed_124__61_, chained_data_delayed_124__60_, chained_data_delayed_124__59_, chained_data_delayed_124__58_, chained_data_delayed_124__57_, chained_data_delayed_124__56_, chained_data_delayed_124__55_, chained_data_delayed_124__54_, chained_data_delayed_124__53_, chained_data_delayed_124__52_, chained_data_delayed_124__51_, chained_data_delayed_124__50_, chained_data_delayed_124__49_, chained_data_delayed_124__48_, chained_data_delayed_124__47_, chained_data_delayed_124__46_, chained_data_delayed_124__45_, chained_data_delayed_124__44_, chained_data_delayed_124__43_, chained_data_delayed_124__42_, chained_data_delayed_124__41_, chained_data_delayed_124__40_, chained_data_delayed_124__39_, chained_data_delayed_124__38_, chained_data_delayed_124__37_, chained_data_delayed_124__36_, chained_data_delayed_124__35_, chained_data_delayed_124__34_, chained_data_delayed_124__33_, chained_data_delayed_124__32_, chained_data_delayed_124__31_, chained_data_delayed_124__30_, chained_data_delayed_124__29_, chained_data_delayed_124__28_, chained_data_delayed_124__27_, chained_data_delayed_124__26_, chained_data_delayed_124__25_, chained_data_delayed_124__24_, chained_data_delayed_124__23_, chained_data_delayed_124__22_, chained_data_delayed_124__21_, chained_data_delayed_124__20_, chained_data_delayed_124__19_, chained_data_delayed_124__18_, chained_data_delayed_124__17_, chained_data_delayed_124__16_, chained_data_delayed_124__15_, chained_data_delayed_124__14_, chained_data_delayed_124__13_, chained_data_delayed_124__12_, chained_data_delayed_124__11_, chained_data_delayed_124__10_, chained_data_delayed_124__9_, chained_data_delayed_124__8_, chained_data_delayed_124__7_, chained_data_delayed_124__6_, chained_data_delayed_124__5_, chained_data_delayed_124__4_, chained_data_delayed_124__3_, chained_data_delayed_124__2_, chained_data_delayed_124__1_, chained_data_delayed_124__0_ }),
    .data_o({ chained_data_delayed_125__127_, chained_data_delayed_125__126_, chained_data_delayed_125__125_, chained_data_delayed_125__124_, chained_data_delayed_125__123_, chained_data_delayed_125__122_, chained_data_delayed_125__121_, chained_data_delayed_125__120_, chained_data_delayed_125__119_, chained_data_delayed_125__118_, chained_data_delayed_125__117_, chained_data_delayed_125__116_, chained_data_delayed_125__115_, chained_data_delayed_125__114_, chained_data_delayed_125__113_, chained_data_delayed_125__112_, chained_data_delayed_125__111_, chained_data_delayed_125__110_, chained_data_delayed_125__109_, chained_data_delayed_125__108_, chained_data_delayed_125__107_, chained_data_delayed_125__106_, chained_data_delayed_125__105_, chained_data_delayed_125__104_, chained_data_delayed_125__103_, chained_data_delayed_125__102_, chained_data_delayed_125__101_, chained_data_delayed_125__100_, chained_data_delayed_125__99_, chained_data_delayed_125__98_, chained_data_delayed_125__97_, chained_data_delayed_125__96_, chained_data_delayed_125__95_, chained_data_delayed_125__94_, chained_data_delayed_125__93_, chained_data_delayed_125__92_, chained_data_delayed_125__91_, chained_data_delayed_125__90_, chained_data_delayed_125__89_, chained_data_delayed_125__88_, chained_data_delayed_125__87_, chained_data_delayed_125__86_, chained_data_delayed_125__85_, chained_data_delayed_125__84_, chained_data_delayed_125__83_, chained_data_delayed_125__82_, chained_data_delayed_125__81_, chained_data_delayed_125__80_, chained_data_delayed_125__79_, chained_data_delayed_125__78_, chained_data_delayed_125__77_, chained_data_delayed_125__76_, chained_data_delayed_125__75_, chained_data_delayed_125__74_, chained_data_delayed_125__73_, chained_data_delayed_125__72_, chained_data_delayed_125__71_, chained_data_delayed_125__70_, chained_data_delayed_125__69_, chained_data_delayed_125__68_, chained_data_delayed_125__67_, chained_data_delayed_125__66_, chained_data_delayed_125__65_, chained_data_delayed_125__64_, chained_data_delayed_125__63_, chained_data_delayed_125__62_, chained_data_delayed_125__61_, chained_data_delayed_125__60_, chained_data_delayed_125__59_, chained_data_delayed_125__58_, chained_data_delayed_125__57_, chained_data_delayed_125__56_, chained_data_delayed_125__55_, chained_data_delayed_125__54_, chained_data_delayed_125__53_, chained_data_delayed_125__52_, chained_data_delayed_125__51_, chained_data_delayed_125__50_, chained_data_delayed_125__49_, chained_data_delayed_125__48_, chained_data_delayed_125__47_, chained_data_delayed_125__46_, chained_data_delayed_125__45_, chained_data_delayed_125__44_, chained_data_delayed_125__43_, chained_data_delayed_125__42_, chained_data_delayed_125__41_, chained_data_delayed_125__40_, chained_data_delayed_125__39_, chained_data_delayed_125__38_, chained_data_delayed_125__37_, chained_data_delayed_125__36_, chained_data_delayed_125__35_, chained_data_delayed_125__34_, chained_data_delayed_125__33_, chained_data_delayed_125__32_, chained_data_delayed_125__31_, chained_data_delayed_125__30_, chained_data_delayed_125__29_, chained_data_delayed_125__28_, chained_data_delayed_125__27_, chained_data_delayed_125__26_, chained_data_delayed_125__25_, chained_data_delayed_125__24_, chained_data_delayed_125__23_, chained_data_delayed_125__22_, chained_data_delayed_125__21_, chained_data_delayed_125__20_, chained_data_delayed_125__19_, chained_data_delayed_125__18_, chained_data_delayed_125__17_, chained_data_delayed_125__16_, chained_data_delayed_125__15_, chained_data_delayed_125__14_, chained_data_delayed_125__13_, chained_data_delayed_125__12_, chained_data_delayed_125__11_, chained_data_delayed_125__10_, chained_data_delayed_125__9_, chained_data_delayed_125__8_, chained_data_delayed_125__7_, chained_data_delayed_125__6_, chained_data_delayed_125__5_, chained_data_delayed_125__4_, chained_data_delayed_125__3_, chained_data_delayed_125__2_, chained_data_delayed_125__1_, chained_data_delayed_125__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_126__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_125__127_, chained_data_delayed_125__126_, chained_data_delayed_125__125_, chained_data_delayed_125__124_, chained_data_delayed_125__123_, chained_data_delayed_125__122_, chained_data_delayed_125__121_, chained_data_delayed_125__120_, chained_data_delayed_125__119_, chained_data_delayed_125__118_, chained_data_delayed_125__117_, chained_data_delayed_125__116_, chained_data_delayed_125__115_, chained_data_delayed_125__114_, chained_data_delayed_125__113_, chained_data_delayed_125__112_, chained_data_delayed_125__111_, chained_data_delayed_125__110_, chained_data_delayed_125__109_, chained_data_delayed_125__108_, chained_data_delayed_125__107_, chained_data_delayed_125__106_, chained_data_delayed_125__105_, chained_data_delayed_125__104_, chained_data_delayed_125__103_, chained_data_delayed_125__102_, chained_data_delayed_125__101_, chained_data_delayed_125__100_, chained_data_delayed_125__99_, chained_data_delayed_125__98_, chained_data_delayed_125__97_, chained_data_delayed_125__96_, chained_data_delayed_125__95_, chained_data_delayed_125__94_, chained_data_delayed_125__93_, chained_data_delayed_125__92_, chained_data_delayed_125__91_, chained_data_delayed_125__90_, chained_data_delayed_125__89_, chained_data_delayed_125__88_, chained_data_delayed_125__87_, chained_data_delayed_125__86_, chained_data_delayed_125__85_, chained_data_delayed_125__84_, chained_data_delayed_125__83_, chained_data_delayed_125__82_, chained_data_delayed_125__81_, chained_data_delayed_125__80_, chained_data_delayed_125__79_, chained_data_delayed_125__78_, chained_data_delayed_125__77_, chained_data_delayed_125__76_, chained_data_delayed_125__75_, chained_data_delayed_125__74_, chained_data_delayed_125__73_, chained_data_delayed_125__72_, chained_data_delayed_125__71_, chained_data_delayed_125__70_, chained_data_delayed_125__69_, chained_data_delayed_125__68_, chained_data_delayed_125__67_, chained_data_delayed_125__66_, chained_data_delayed_125__65_, chained_data_delayed_125__64_, chained_data_delayed_125__63_, chained_data_delayed_125__62_, chained_data_delayed_125__61_, chained_data_delayed_125__60_, chained_data_delayed_125__59_, chained_data_delayed_125__58_, chained_data_delayed_125__57_, chained_data_delayed_125__56_, chained_data_delayed_125__55_, chained_data_delayed_125__54_, chained_data_delayed_125__53_, chained_data_delayed_125__52_, chained_data_delayed_125__51_, chained_data_delayed_125__50_, chained_data_delayed_125__49_, chained_data_delayed_125__48_, chained_data_delayed_125__47_, chained_data_delayed_125__46_, chained_data_delayed_125__45_, chained_data_delayed_125__44_, chained_data_delayed_125__43_, chained_data_delayed_125__42_, chained_data_delayed_125__41_, chained_data_delayed_125__40_, chained_data_delayed_125__39_, chained_data_delayed_125__38_, chained_data_delayed_125__37_, chained_data_delayed_125__36_, chained_data_delayed_125__35_, chained_data_delayed_125__34_, chained_data_delayed_125__33_, chained_data_delayed_125__32_, chained_data_delayed_125__31_, chained_data_delayed_125__30_, chained_data_delayed_125__29_, chained_data_delayed_125__28_, chained_data_delayed_125__27_, chained_data_delayed_125__26_, chained_data_delayed_125__25_, chained_data_delayed_125__24_, chained_data_delayed_125__23_, chained_data_delayed_125__22_, chained_data_delayed_125__21_, chained_data_delayed_125__20_, chained_data_delayed_125__19_, chained_data_delayed_125__18_, chained_data_delayed_125__17_, chained_data_delayed_125__16_, chained_data_delayed_125__15_, chained_data_delayed_125__14_, chained_data_delayed_125__13_, chained_data_delayed_125__12_, chained_data_delayed_125__11_, chained_data_delayed_125__10_, chained_data_delayed_125__9_, chained_data_delayed_125__8_, chained_data_delayed_125__7_, chained_data_delayed_125__6_, chained_data_delayed_125__5_, chained_data_delayed_125__4_, chained_data_delayed_125__3_, chained_data_delayed_125__2_, chained_data_delayed_125__1_, chained_data_delayed_125__0_ }),
    .data_o({ chained_data_delayed_126__127_, chained_data_delayed_126__126_, chained_data_delayed_126__125_, chained_data_delayed_126__124_, chained_data_delayed_126__123_, chained_data_delayed_126__122_, chained_data_delayed_126__121_, chained_data_delayed_126__120_, chained_data_delayed_126__119_, chained_data_delayed_126__118_, chained_data_delayed_126__117_, chained_data_delayed_126__116_, chained_data_delayed_126__115_, chained_data_delayed_126__114_, chained_data_delayed_126__113_, chained_data_delayed_126__112_, chained_data_delayed_126__111_, chained_data_delayed_126__110_, chained_data_delayed_126__109_, chained_data_delayed_126__108_, chained_data_delayed_126__107_, chained_data_delayed_126__106_, chained_data_delayed_126__105_, chained_data_delayed_126__104_, chained_data_delayed_126__103_, chained_data_delayed_126__102_, chained_data_delayed_126__101_, chained_data_delayed_126__100_, chained_data_delayed_126__99_, chained_data_delayed_126__98_, chained_data_delayed_126__97_, chained_data_delayed_126__96_, chained_data_delayed_126__95_, chained_data_delayed_126__94_, chained_data_delayed_126__93_, chained_data_delayed_126__92_, chained_data_delayed_126__91_, chained_data_delayed_126__90_, chained_data_delayed_126__89_, chained_data_delayed_126__88_, chained_data_delayed_126__87_, chained_data_delayed_126__86_, chained_data_delayed_126__85_, chained_data_delayed_126__84_, chained_data_delayed_126__83_, chained_data_delayed_126__82_, chained_data_delayed_126__81_, chained_data_delayed_126__80_, chained_data_delayed_126__79_, chained_data_delayed_126__78_, chained_data_delayed_126__77_, chained_data_delayed_126__76_, chained_data_delayed_126__75_, chained_data_delayed_126__74_, chained_data_delayed_126__73_, chained_data_delayed_126__72_, chained_data_delayed_126__71_, chained_data_delayed_126__70_, chained_data_delayed_126__69_, chained_data_delayed_126__68_, chained_data_delayed_126__67_, chained_data_delayed_126__66_, chained_data_delayed_126__65_, chained_data_delayed_126__64_, chained_data_delayed_126__63_, chained_data_delayed_126__62_, chained_data_delayed_126__61_, chained_data_delayed_126__60_, chained_data_delayed_126__59_, chained_data_delayed_126__58_, chained_data_delayed_126__57_, chained_data_delayed_126__56_, chained_data_delayed_126__55_, chained_data_delayed_126__54_, chained_data_delayed_126__53_, chained_data_delayed_126__52_, chained_data_delayed_126__51_, chained_data_delayed_126__50_, chained_data_delayed_126__49_, chained_data_delayed_126__48_, chained_data_delayed_126__47_, chained_data_delayed_126__46_, chained_data_delayed_126__45_, chained_data_delayed_126__44_, chained_data_delayed_126__43_, chained_data_delayed_126__42_, chained_data_delayed_126__41_, chained_data_delayed_126__40_, chained_data_delayed_126__39_, chained_data_delayed_126__38_, chained_data_delayed_126__37_, chained_data_delayed_126__36_, chained_data_delayed_126__35_, chained_data_delayed_126__34_, chained_data_delayed_126__33_, chained_data_delayed_126__32_, chained_data_delayed_126__31_, chained_data_delayed_126__30_, chained_data_delayed_126__29_, chained_data_delayed_126__28_, chained_data_delayed_126__27_, chained_data_delayed_126__26_, chained_data_delayed_126__25_, chained_data_delayed_126__24_, chained_data_delayed_126__23_, chained_data_delayed_126__22_, chained_data_delayed_126__21_, chained_data_delayed_126__20_, chained_data_delayed_126__19_, chained_data_delayed_126__18_, chained_data_delayed_126__17_, chained_data_delayed_126__16_, chained_data_delayed_126__15_, chained_data_delayed_126__14_, chained_data_delayed_126__13_, chained_data_delayed_126__12_, chained_data_delayed_126__11_, chained_data_delayed_126__10_, chained_data_delayed_126__9_, chained_data_delayed_126__8_, chained_data_delayed_126__7_, chained_data_delayed_126__6_, chained_data_delayed_126__5_, chained_data_delayed_126__4_, chained_data_delayed_126__3_, chained_data_delayed_126__2_, chained_data_delayed_126__1_, chained_data_delayed_126__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_127__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_126__127_, chained_data_delayed_126__126_, chained_data_delayed_126__125_, chained_data_delayed_126__124_, chained_data_delayed_126__123_, chained_data_delayed_126__122_, chained_data_delayed_126__121_, chained_data_delayed_126__120_, chained_data_delayed_126__119_, chained_data_delayed_126__118_, chained_data_delayed_126__117_, chained_data_delayed_126__116_, chained_data_delayed_126__115_, chained_data_delayed_126__114_, chained_data_delayed_126__113_, chained_data_delayed_126__112_, chained_data_delayed_126__111_, chained_data_delayed_126__110_, chained_data_delayed_126__109_, chained_data_delayed_126__108_, chained_data_delayed_126__107_, chained_data_delayed_126__106_, chained_data_delayed_126__105_, chained_data_delayed_126__104_, chained_data_delayed_126__103_, chained_data_delayed_126__102_, chained_data_delayed_126__101_, chained_data_delayed_126__100_, chained_data_delayed_126__99_, chained_data_delayed_126__98_, chained_data_delayed_126__97_, chained_data_delayed_126__96_, chained_data_delayed_126__95_, chained_data_delayed_126__94_, chained_data_delayed_126__93_, chained_data_delayed_126__92_, chained_data_delayed_126__91_, chained_data_delayed_126__90_, chained_data_delayed_126__89_, chained_data_delayed_126__88_, chained_data_delayed_126__87_, chained_data_delayed_126__86_, chained_data_delayed_126__85_, chained_data_delayed_126__84_, chained_data_delayed_126__83_, chained_data_delayed_126__82_, chained_data_delayed_126__81_, chained_data_delayed_126__80_, chained_data_delayed_126__79_, chained_data_delayed_126__78_, chained_data_delayed_126__77_, chained_data_delayed_126__76_, chained_data_delayed_126__75_, chained_data_delayed_126__74_, chained_data_delayed_126__73_, chained_data_delayed_126__72_, chained_data_delayed_126__71_, chained_data_delayed_126__70_, chained_data_delayed_126__69_, chained_data_delayed_126__68_, chained_data_delayed_126__67_, chained_data_delayed_126__66_, chained_data_delayed_126__65_, chained_data_delayed_126__64_, chained_data_delayed_126__63_, chained_data_delayed_126__62_, chained_data_delayed_126__61_, chained_data_delayed_126__60_, chained_data_delayed_126__59_, chained_data_delayed_126__58_, chained_data_delayed_126__57_, chained_data_delayed_126__56_, chained_data_delayed_126__55_, chained_data_delayed_126__54_, chained_data_delayed_126__53_, chained_data_delayed_126__52_, chained_data_delayed_126__51_, chained_data_delayed_126__50_, chained_data_delayed_126__49_, chained_data_delayed_126__48_, chained_data_delayed_126__47_, chained_data_delayed_126__46_, chained_data_delayed_126__45_, chained_data_delayed_126__44_, chained_data_delayed_126__43_, chained_data_delayed_126__42_, chained_data_delayed_126__41_, chained_data_delayed_126__40_, chained_data_delayed_126__39_, chained_data_delayed_126__38_, chained_data_delayed_126__37_, chained_data_delayed_126__36_, chained_data_delayed_126__35_, chained_data_delayed_126__34_, chained_data_delayed_126__33_, chained_data_delayed_126__32_, chained_data_delayed_126__31_, chained_data_delayed_126__30_, chained_data_delayed_126__29_, chained_data_delayed_126__28_, chained_data_delayed_126__27_, chained_data_delayed_126__26_, chained_data_delayed_126__25_, chained_data_delayed_126__24_, chained_data_delayed_126__23_, chained_data_delayed_126__22_, chained_data_delayed_126__21_, chained_data_delayed_126__20_, chained_data_delayed_126__19_, chained_data_delayed_126__18_, chained_data_delayed_126__17_, chained_data_delayed_126__16_, chained_data_delayed_126__15_, chained_data_delayed_126__14_, chained_data_delayed_126__13_, chained_data_delayed_126__12_, chained_data_delayed_126__11_, chained_data_delayed_126__10_, chained_data_delayed_126__9_, chained_data_delayed_126__8_, chained_data_delayed_126__7_, chained_data_delayed_126__6_, chained_data_delayed_126__5_, chained_data_delayed_126__4_, chained_data_delayed_126__3_, chained_data_delayed_126__2_, chained_data_delayed_126__1_, chained_data_delayed_126__0_ }),
    .data_o({ chained_data_delayed_127__127_, chained_data_delayed_127__126_, chained_data_delayed_127__125_, chained_data_delayed_127__124_, chained_data_delayed_127__123_, chained_data_delayed_127__122_, chained_data_delayed_127__121_, chained_data_delayed_127__120_, chained_data_delayed_127__119_, chained_data_delayed_127__118_, chained_data_delayed_127__117_, chained_data_delayed_127__116_, chained_data_delayed_127__115_, chained_data_delayed_127__114_, chained_data_delayed_127__113_, chained_data_delayed_127__112_, chained_data_delayed_127__111_, chained_data_delayed_127__110_, chained_data_delayed_127__109_, chained_data_delayed_127__108_, chained_data_delayed_127__107_, chained_data_delayed_127__106_, chained_data_delayed_127__105_, chained_data_delayed_127__104_, chained_data_delayed_127__103_, chained_data_delayed_127__102_, chained_data_delayed_127__101_, chained_data_delayed_127__100_, chained_data_delayed_127__99_, chained_data_delayed_127__98_, chained_data_delayed_127__97_, chained_data_delayed_127__96_, chained_data_delayed_127__95_, chained_data_delayed_127__94_, chained_data_delayed_127__93_, chained_data_delayed_127__92_, chained_data_delayed_127__91_, chained_data_delayed_127__90_, chained_data_delayed_127__89_, chained_data_delayed_127__88_, chained_data_delayed_127__87_, chained_data_delayed_127__86_, chained_data_delayed_127__85_, chained_data_delayed_127__84_, chained_data_delayed_127__83_, chained_data_delayed_127__82_, chained_data_delayed_127__81_, chained_data_delayed_127__80_, chained_data_delayed_127__79_, chained_data_delayed_127__78_, chained_data_delayed_127__77_, chained_data_delayed_127__76_, chained_data_delayed_127__75_, chained_data_delayed_127__74_, chained_data_delayed_127__73_, chained_data_delayed_127__72_, chained_data_delayed_127__71_, chained_data_delayed_127__70_, chained_data_delayed_127__69_, chained_data_delayed_127__68_, chained_data_delayed_127__67_, chained_data_delayed_127__66_, chained_data_delayed_127__65_, chained_data_delayed_127__64_, chained_data_delayed_127__63_, chained_data_delayed_127__62_, chained_data_delayed_127__61_, chained_data_delayed_127__60_, chained_data_delayed_127__59_, chained_data_delayed_127__58_, chained_data_delayed_127__57_, chained_data_delayed_127__56_, chained_data_delayed_127__55_, chained_data_delayed_127__54_, chained_data_delayed_127__53_, chained_data_delayed_127__52_, chained_data_delayed_127__51_, chained_data_delayed_127__50_, chained_data_delayed_127__49_, chained_data_delayed_127__48_, chained_data_delayed_127__47_, chained_data_delayed_127__46_, chained_data_delayed_127__45_, chained_data_delayed_127__44_, chained_data_delayed_127__43_, chained_data_delayed_127__42_, chained_data_delayed_127__41_, chained_data_delayed_127__40_, chained_data_delayed_127__39_, chained_data_delayed_127__38_, chained_data_delayed_127__37_, chained_data_delayed_127__36_, chained_data_delayed_127__35_, chained_data_delayed_127__34_, chained_data_delayed_127__33_, chained_data_delayed_127__32_, chained_data_delayed_127__31_, chained_data_delayed_127__30_, chained_data_delayed_127__29_, chained_data_delayed_127__28_, chained_data_delayed_127__27_, chained_data_delayed_127__26_, chained_data_delayed_127__25_, chained_data_delayed_127__24_, chained_data_delayed_127__23_, chained_data_delayed_127__22_, chained_data_delayed_127__21_, chained_data_delayed_127__20_, chained_data_delayed_127__19_, chained_data_delayed_127__18_, chained_data_delayed_127__17_, chained_data_delayed_127__16_, chained_data_delayed_127__15_, chained_data_delayed_127__14_, chained_data_delayed_127__13_, chained_data_delayed_127__12_, chained_data_delayed_127__11_, chained_data_delayed_127__10_, chained_data_delayed_127__9_, chained_data_delayed_127__8_, chained_data_delayed_127__7_, chained_data_delayed_127__6_, chained_data_delayed_127__5_, chained_data_delayed_127__4_, chained_data_delayed_127__3_, chained_data_delayed_127__2_, chained_data_delayed_127__1_, chained_data_delayed_127__0_ })
  );


  bsg_dff_width_p128
  chained_genblk1_128__ch_reg
  (
    .clk_i(clk_i),
    .data_i({ chained_data_delayed_127__127_, chained_data_delayed_127__126_, chained_data_delayed_127__125_, chained_data_delayed_127__124_, chained_data_delayed_127__123_, chained_data_delayed_127__122_, chained_data_delayed_127__121_, chained_data_delayed_127__120_, chained_data_delayed_127__119_, chained_data_delayed_127__118_, chained_data_delayed_127__117_, chained_data_delayed_127__116_, chained_data_delayed_127__115_, chained_data_delayed_127__114_, chained_data_delayed_127__113_, chained_data_delayed_127__112_, chained_data_delayed_127__111_, chained_data_delayed_127__110_, chained_data_delayed_127__109_, chained_data_delayed_127__108_, chained_data_delayed_127__107_, chained_data_delayed_127__106_, chained_data_delayed_127__105_, chained_data_delayed_127__104_, chained_data_delayed_127__103_, chained_data_delayed_127__102_, chained_data_delayed_127__101_, chained_data_delayed_127__100_, chained_data_delayed_127__99_, chained_data_delayed_127__98_, chained_data_delayed_127__97_, chained_data_delayed_127__96_, chained_data_delayed_127__95_, chained_data_delayed_127__94_, chained_data_delayed_127__93_, chained_data_delayed_127__92_, chained_data_delayed_127__91_, chained_data_delayed_127__90_, chained_data_delayed_127__89_, chained_data_delayed_127__88_, chained_data_delayed_127__87_, chained_data_delayed_127__86_, chained_data_delayed_127__85_, chained_data_delayed_127__84_, chained_data_delayed_127__83_, chained_data_delayed_127__82_, chained_data_delayed_127__81_, chained_data_delayed_127__80_, chained_data_delayed_127__79_, chained_data_delayed_127__78_, chained_data_delayed_127__77_, chained_data_delayed_127__76_, chained_data_delayed_127__75_, chained_data_delayed_127__74_, chained_data_delayed_127__73_, chained_data_delayed_127__72_, chained_data_delayed_127__71_, chained_data_delayed_127__70_, chained_data_delayed_127__69_, chained_data_delayed_127__68_, chained_data_delayed_127__67_, chained_data_delayed_127__66_, chained_data_delayed_127__65_, chained_data_delayed_127__64_, chained_data_delayed_127__63_, chained_data_delayed_127__62_, chained_data_delayed_127__61_, chained_data_delayed_127__60_, chained_data_delayed_127__59_, chained_data_delayed_127__58_, chained_data_delayed_127__57_, chained_data_delayed_127__56_, chained_data_delayed_127__55_, chained_data_delayed_127__54_, chained_data_delayed_127__53_, chained_data_delayed_127__52_, chained_data_delayed_127__51_, chained_data_delayed_127__50_, chained_data_delayed_127__49_, chained_data_delayed_127__48_, chained_data_delayed_127__47_, chained_data_delayed_127__46_, chained_data_delayed_127__45_, chained_data_delayed_127__44_, chained_data_delayed_127__43_, chained_data_delayed_127__42_, chained_data_delayed_127__41_, chained_data_delayed_127__40_, chained_data_delayed_127__39_, chained_data_delayed_127__38_, chained_data_delayed_127__37_, chained_data_delayed_127__36_, chained_data_delayed_127__35_, chained_data_delayed_127__34_, chained_data_delayed_127__33_, chained_data_delayed_127__32_, chained_data_delayed_127__31_, chained_data_delayed_127__30_, chained_data_delayed_127__29_, chained_data_delayed_127__28_, chained_data_delayed_127__27_, chained_data_delayed_127__26_, chained_data_delayed_127__25_, chained_data_delayed_127__24_, chained_data_delayed_127__23_, chained_data_delayed_127__22_, chained_data_delayed_127__21_, chained_data_delayed_127__20_, chained_data_delayed_127__19_, chained_data_delayed_127__18_, chained_data_delayed_127__17_, chained_data_delayed_127__16_, chained_data_delayed_127__15_, chained_data_delayed_127__14_, chained_data_delayed_127__13_, chained_data_delayed_127__12_, chained_data_delayed_127__11_, chained_data_delayed_127__10_, chained_data_delayed_127__9_, chained_data_delayed_127__8_, chained_data_delayed_127__7_, chained_data_delayed_127__6_, chained_data_delayed_127__5_, chained_data_delayed_127__4_, chained_data_delayed_127__3_, chained_data_delayed_127__2_, chained_data_delayed_127__1_, chained_data_delayed_127__0_ }),
    .data_o(data_o)
  );


endmodule

