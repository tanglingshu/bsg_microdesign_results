

module top
(
  i,
  o
);

  input [639:0] i;
  output [9:0] o;

  bsg_reduce_segmented
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_reduce_segmented
(
  i,
  o
);

  input [639:0] i;
  output [9:0] o;
  wire [9:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619;
  assign o[0] = N61 | i[0];
  assign N61 = N60 | i[1];
  assign N60 = N59 | i[2];
  assign N59 = N58 | i[3];
  assign N58 = N57 | i[4];
  assign N57 = N56 | i[5];
  assign N56 = N55 | i[6];
  assign N55 = N54 | i[7];
  assign N54 = N53 | i[8];
  assign N53 = N52 | i[9];
  assign N52 = N51 | i[10];
  assign N51 = N50 | i[11];
  assign N50 = N49 | i[12];
  assign N49 = N48 | i[13];
  assign N48 = N47 | i[14];
  assign N47 = N46 | i[15];
  assign N46 = N45 | i[16];
  assign N45 = N44 | i[17];
  assign N44 = N43 | i[18];
  assign N43 = N42 | i[19];
  assign N42 = N41 | i[20];
  assign N41 = N40 | i[21];
  assign N40 = N39 | i[22];
  assign N39 = N38 | i[23];
  assign N38 = N37 | i[24];
  assign N37 = N36 | i[25];
  assign N36 = N35 | i[26];
  assign N35 = N34 | i[27];
  assign N34 = N33 | i[28];
  assign N33 = N32 | i[29];
  assign N32 = N31 | i[30];
  assign N31 = N30 | i[31];
  assign N30 = N29 | i[32];
  assign N29 = N28 | i[33];
  assign N28 = N27 | i[34];
  assign N27 = N26 | i[35];
  assign N26 = N25 | i[36];
  assign N25 = N24 | i[37];
  assign N24 = N23 | i[38];
  assign N23 = N22 | i[39];
  assign N22 = N21 | i[40];
  assign N21 = N20 | i[41];
  assign N20 = N19 | i[42];
  assign N19 = N18 | i[43];
  assign N18 = N17 | i[44];
  assign N17 = N16 | i[45];
  assign N16 = N15 | i[46];
  assign N15 = N14 | i[47];
  assign N14 = N13 | i[48];
  assign N13 = N12 | i[49];
  assign N12 = N11 | i[50];
  assign N11 = N10 | i[51];
  assign N10 = N9 | i[52];
  assign N9 = N8 | i[53];
  assign N8 = N7 | i[54];
  assign N7 = N6 | i[55];
  assign N6 = N5 | i[56];
  assign N5 = N4 | i[57];
  assign N4 = N3 | i[58];
  assign N3 = N2 | i[59];
  assign N2 = N1 | i[60];
  assign N1 = N0 | i[61];
  assign N0 = i[63] | i[62];
  assign o[1] = N123 | i[64];
  assign N123 = N122 | i[65];
  assign N122 = N121 | i[66];
  assign N121 = N120 | i[67];
  assign N120 = N119 | i[68];
  assign N119 = N118 | i[69];
  assign N118 = N117 | i[70];
  assign N117 = N116 | i[71];
  assign N116 = N115 | i[72];
  assign N115 = N114 | i[73];
  assign N114 = N113 | i[74];
  assign N113 = N112 | i[75];
  assign N112 = N111 | i[76];
  assign N111 = N110 | i[77];
  assign N110 = N109 | i[78];
  assign N109 = N108 | i[79];
  assign N108 = N107 | i[80];
  assign N107 = N106 | i[81];
  assign N106 = N105 | i[82];
  assign N105 = N104 | i[83];
  assign N104 = N103 | i[84];
  assign N103 = N102 | i[85];
  assign N102 = N101 | i[86];
  assign N101 = N100 | i[87];
  assign N100 = N99 | i[88];
  assign N99 = N98 | i[89];
  assign N98 = N97 | i[90];
  assign N97 = N96 | i[91];
  assign N96 = N95 | i[92];
  assign N95 = N94 | i[93];
  assign N94 = N93 | i[94];
  assign N93 = N92 | i[95];
  assign N92 = N91 | i[96];
  assign N91 = N90 | i[97];
  assign N90 = N89 | i[98];
  assign N89 = N88 | i[99];
  assign N88 = N87 | i[100];
  assign N87 = N86 | i[101];
  assign N86 = N85 | i[102];
  assign N85 = N84 | i[103];
  assign N84 = N83 | i[104];
  assign N83 = N82 | i[105];
  assign N82 = N81 | i[106];
  assign N81 = N80 | i[107];
  assign N80 = N79 | i[108];
  assign N79 = N78 | i[109];
  assign N78 = N77 | i[110];
  assign N77 = N76 | i[111];
  assign N76 = N75 | i[112];
  assign N75 = N74 | i[113];
  assign N74 = N73 | i[114];
  assign N73 = N72 | i[115];
  assign N72 = N71 | i[116];
  assign N71 = N70 | i[117];
  assign N70 = N69 | i[118];
  assign N69 = N68 | i[119];
  assign N68 = N67 | i[120];
  assign N67 = N66 | i[121];
  assign N66 = N65 | i[122];
  assign N65 = N64 | i[123];
  assign N64 = N63 | i[124];
  assign N63 = N62 | i[125];
  assign N62 = i[127] | i[126];
  assign o[2] = N185 | i[128];
  assign N185 = N184 | i[129];
  assign N184 = N183 | i[130];
  assign N183 = N182 | i[131];
  assign N182 = N181 | i[132];
  assign N181 = N180 | i[133];
  assign N180 = N179 | i[134];
  assign N179 = N178 | i[135];
  assign N178 = N177 | i[136];
  assign N177 = N176 | i[137];
  assign N176 = N175 | i[138];
  assign N175 = N174 | i[139];
  assign N174 = N173 | i[140];
  assign N173 = N172 | i[141];
  assign N172 = N171 | i[142];
  assign N171 = N170 | i[143];
  assign N170 = N169 | i[144];
  assign N169 = N168 | i[145];
  assign N168 = N167 | i[146];
  assign N167 = N166 | i[147];
  assign N166 = N165 | i[148];
  assign N165 = N164 | i[149];
  assign N164 = N163 | i[150];
  assign N163 = N162 | i[151];
  assign N162 = N161 | i[152];
  assign N161 = N160 | i[153];
  assign N160 = N159 | i[154];
  assign N159 = N158 | i[155];
  assign N158 = N157 | i[156];
  assign N157 = N156 | i[157];
  assign N156 = N155 | i[158];
  assign N155 = N154 | i[159];
  assign N154 = N153 | i[160];
  assign N153 = N152 | i[161];
  assign N152 = N151 | i[162];
  assign N151 = N150 | i[163];
  assign N150 = N149 | i[164];
  assign N149 = N148 | i[165];
  assign N148 = N147 | i[166];
  assign N147 = N146 | i[167];
  assign N146 = N145 | i[168];
  assign N145 = N144 | i[169];
  assign N144 = N143 | i[170];
  assign N143 = N142 | i[171];
  assign N142 = N141 | i[172];
  assign N141 = N140 | i[173];
  assign N140 = N139 | i[174];
  assign N139 = N138 | i[175];
  assign N138 = N137 | i[176];
  assign N137 = N136 | i[177];
  assign N136 = N135 | i[178];
  assign N135 = N134 | i[179];
  assign N134 = N133 | i[180];
  assign N133 = N132 | i[181];
  assign N132 = N131 | i[182];
  assign N131 = N130 | i[183];
  assign N130 = N129 | i[184];
  assign N129 = N128 | i[185];
  assign N128 = N127 | i[186];
  assign N127 = N126 | i[187];
  assign N126 = N125 | i[188];
  assign N125 = N124 | i[189];
  assign N124 = i[191] | i[190];
  assign o[3] = N247 | i[192];
  assign N247 = N246 | i[193];
  assign N246 = N245 | i[194];
  assign N245 = N244 | i[195];
  assign N244 = N243 | i[196];
  assign N243 = N242 | i[197];
  assign N242 = N241 | i[198];
  assign N241 = N240 | i[199];
  assign N240 = N239 | i[200];
  assign N239 = N238 | i[201];
  assign N238 = N237 | i[202];
  assign N237 = N236 | i[203];
  assign N236 = N235 | i[204];
  assign N235 = N234 | i[205];
  assign N234 = N233 | i[206];
  assign N233 = N232 | i[207];
  assign N232 = N231 | i[208];
  assign N231 = N230 | i[209];
  assign N230 = N229 | i[210];
  assign N229 = N228 | i[211];
  assign N228 = N227 | i[212];
  assign N227 = N226 | i[213];
  assign N226 = N225 | i[214];
  assign N225 = N224 | i[215];
  assign N224 = N223 | i[216];
  assign N223 = N222 | i[217];
  assign N222 = N221 | i[218];
  assign N221 = N220 | i[219];
  assign N220 = N219 | i[220];
  assign N219 = N218 | i[221];
  assign N218 = N217 | i[222];
  assign N217 = N216 | i[223];
  assign N216 = N215 | i[224];
  assign N215 = N214 | i[225];
  assign N214 = N213 | i[226];
  assign N213 = N212 | i[227];
  assign N212 = N211 | i[228];
  assign N211 = N210 | i[229];
  assign N210 = N209 | i[230];
  assign N209 = N208 | i[231];
  assign N208 = N207 | i[232];
  assign N207 = N206 | i[233];
  assign N206 = N205 | i[234];
  assign N205 = N204 | i[235];
  assign N204 = N203 | i[236];
  assign N203 = N202 | i[237];
  assign N202 = N201 | i[238];
  assign N201 = N200 | i[239];
  assign N200 = N199 | i[240];
  assign N199 = N198 | i[241];
  assign N198 = N197 | i[242];
  assign N197 = N196 | i[243];
  assign N196 = N195 | i[244];
  assign N195 = N194 | i[245];
  assign N194 = N193 | i[246];
  assign N193 = N192 | i[247];
  assign N192 = N191 | i[248];
  assign N191 = N190 | i[249];
  assign N190 = N189 | i[250];
  assign N189 = N188 | i[251];
  assign N188 = N187 | i[252];
  assign N187 = N186 | i[253];
  assign N186 = i[255] | i[254];
  assign o[4] = N309 | i[256];
  assign N309 = N308 | i[257];
  assign N308 = N307 | i[258];
  assign N307 = N306 | i[259];
  assign N306 = N305 | i[260];
  assign N305 = N304 | i[261];
  assign N304 = N303 | i[262];
  assign N303 = N302 | i[263];
  assign N302 = N301 | i[264];
  assign N301 = N300 | i[265];
  assign N300 = N299 | i[266];
  assign N299 = N298 | i[267];
  assign N298 = N297 | i[268];
  assign N297 = N296 | i[269];
  assign N296 = N295 | i[270];
  assign N295 = N294 | i[271];
  assign N294 = N293 | i[272];
  assign N293 = N292 | i[273];
  assign N292 = N291 | i[274];
  assign N291 = N290 | i[275];
  assign N290 = N289 | i[276];
  assign N289 = N288 | i[277];
  assign N288 = N287 | i[278];
  assign N287 = N286 | i[279];
  assign N286 = N285 | i[280];
  assign N285 = N284 | i[281];
  assign N284 = N283 | i[282];
  assign N283 = N282 | i[283];
  assign N282 = N281 | i[284];
  assign N281 = N280 | i[285];
  assign N280 = N279 | i[286];
  assign N279 = N278 | i[287];
  assign N278 = N277 | i[288];
  assign N277 = N276 | i[289];
  assign N276 = N275 | i[290];
  assign N275 = N274 | i[291];
  assign N274 = N273 | i[292];
  assign N273 = N272 | i[293];
  assign N272 = N271 | i[294];
  assign N271 = N270 | i[295];
  assign N270 = N269 | i[296];
  assign N269 = N268 | i[297];
  assign N268 = N267 | i[298];
  assign N267 = N266 | i[299];
  assign N266 = N265 | i[300];
  assign N265 = N264 | i[301];
  assign N264 = N263 | i[302];
  assign N263 = N262 | i[303];
  assign N262 = N261 | i[304];
  assign N261 = N260 | i[305];
  assign N260 = N259 | i[306];
  assign N259 = N258 | i[307];
  assign N258 = N257 | i[308];
  assign N257 = N256 | i[309];
  assign N256 = N255 | i[310];
  assign N255 = N254 | i[311];
  assign N254 = N253 | i[312];
  assign N253 = N252 | i[313];
  assign N252 = N251 | i[314];
  assign N251 = N250 | i[315];
  assign N250 = N249 | i[316];
  assign N249 = N248 | i[317];
  assign N248 = i[319] | i[318];
  assign o[5] = N371 | i[320];
  assign N371 = N370 | i[321];
  assign N370 = N369 | i[322];
  assign N369 = N368 | i[323];
  assign N368 = N367 | i[324];
  assign N367 = N366 | i[325];
  assign N366 = N365 | i[326];
  assign N365 = N364 | i[327];
  assign N364 = N363 | i[328];
  assign N363 = N362 | i[329];
  assign N362 = N361 | i[330];
  assign N361 = N360 | i[331];
  assign N360 = N359 | i[332];
  assign N359 = N358 | i[333];
  assign N358 = N357 | i[334];
  assign N357 = N356 | i[335];
  assign N356 = N355 | i[336];
  assign N355 = N354 | i[337];
  assign N354 = N353 | i[338];
  assign N353 = N352 | i[339];
  assign N352 = N351 | i[340];
  assign N351 = N350 | i[341];
  assign N350 = N349 | i[342];
  assign N349 = N348 | i[343];
  assign N348 = N347 | i[344];
  assign N347 = N346 | i[345];
  assign N346 = N345 | i[346];
  assign N345 = N344 | i[347];
  assign N344 = N343 | i[348];
  assign N343 = N342 | i[349];
  assign N342 = N341 | i[350];
  assign N341 = N340 | i[351];
  assign N340 = N339 | i[352];
  assign N339 = N338 | i[353];
  assign N338 = N337 | i[354];
  assign N337 = N336 | i[355];
  assign N336 = N335 | i[356];
  assign N335 = N334 | i[357];
  assign N334 = N333 | i[358];
  assign N333 = N332 | i[359];
  assign N332 = N331 | i[360];
  assign N331 = N330 | i[361];
  assign N330 = N329 | i[362];
  assign N329 = N328 | i[363];
  assign N328 = N327 | i[364];
  assign N327 = N326 | i[365];
  assign N326 = N325 | i[366];
  assign N325 = N324 | i[367];
  assign N324 = N323 | i[368];
  assign N323 = N322 | i[369];
  assign N322 = N321 | i[370];
  assign N321 = N320 | i[371];
  assign N320 = N319 | i[372];
  assign N319 = N318 | i[373];
  assign N318 = N317 | i[374];
  assign N317 = N316 | i[375];
  assign N316 = N315 | i[376];
  assign N315 = N314 | i[377];
  assign N314 = N313 | i[378];
  assign N313 = N312 | i[379];
  assign N312 = N311 | i[380];
  assign N311 = N310 | i[381];
  assign N310 = i[383] | i[382];
  assign o[6] = N433 | i[384];
  assign N433 = N432 | i[385];
  assign N432 = N431 | i[386];
  assign N431 = N430 | i[387];
  assign N430 = N429 | i[388];
  assign N429 = N428 | i[389];
  assign N428 = N427 | i[390];
  assign N427 = N426 | i[391];
  assign N426 = N425 | i[392];
  assign N425 = N424 | i[393];
  assign N424 = N423 | i[394];
  assign N423 = N422 | i[395];
  assign N422 = N421 | i[396];
  assign N421 = N420 | i[397];
  assign N420 = N419 | i[398];
  assign N419 = N418 | i[399];
  assign N418 = N417 | i[400];
  assign N417 = N416 | i[401];
  assign N416 = N415 | i[402];
  assign N415 = N414 | i[403];
  assign N414 = N413 | i[404];
  assign N413 = N412 | i[405];
  assign N412 = N411 | i[406];
  assign N411 = N410 | i[407];
  assign N410 = N409 | i[408];
  assign N409 = N408 | i[409];
  assign N408 = N407 | i[410];
  assign N407 = N406 | i[411];
  assign N406 = N405 | i[412];
  assign N405 = N404 | i[413];
  assign N404 = N403 | i[414];
  assign N403 = N402 | i[415];
  assign N402 = N401 | i[416];
  assign N401 = N400 | i[417];
  assign N400 = N399 | i[418];
  assign N399 = N398 | i[419];
  assign N398 = N397 | i[420];
  assign N397 = N396 | i[421];
  assign N396 = N395 | i[422];
  assign N395 = N394 | i[423];
  assign N394 = N393 | i[424];
  assign N393 = N392 | i[425];
  assign N392 = N391 | i[426];
  assign N391 = N390 | i[427];
  assign N390 = N389 | i[428];
  assign N389 = N388 | i[429];
  assign N388 = N387 | i[430];
  assign N387 = N386 | i[431];
  assign N386 = N385 | i[432];
  assign N385 = N384 | i[433];
  assign N384 = N383 | i[434];
  assign N383 = N382 | i[435];
  assign N382 = N381 | i[436];
  assign N381 = N380 | i[437];
  assign N380 = N379 | i[438];
  assign N379 = N378 | i[439];
  assign N378 = N377 | i[440];
  assign N377 = N376 | i[441];
  assign N376 = N375 | i[442];
  assign N375 = N374 | i[443];
  assign N374 = N373 | i[444];
  assign N373 = N372 | i[445];
  assign N372 = i[447] | i[446];
  assign o[7] = N495 | i[448];
  assign N495 = N494 | i[449];
  assign N494 = N493 | i[450];
  assign N493 = N492 | i[451];
  assign N492 = N491 | i[452];
  assign N491 = N490 | i[453];
  assign N490 = N489 | i[454];
  assign N489 = N488 | i[455];
  assign N488 = N487 | i[456];
  assign N487 = N486 | i[457];
  assign N486 = N485 | i[458];
  assign N485 = N484 | i[459];
  assign N484 = N483 | i[460];
  assign N483 = N482 | i[461];
  assign N482 = N481 | i[462];
  assign N481 = N480 | i[463];
  assign N480 = N479 | i[464];
  assign N479 = N478 | i[465];
  assign N478 = N477 | i[466];
  assign N477 = N476 | i[467];
  assign N476 = N475 | i[468];
  assign N475 = N474 | i[469];
  assign N474 = N473 | i[470];
  assign N473 = N472 | i[471];
  assign N472 = N471 | i[472];
  assign N471 = N470 | i[473];
  assign N470 = N469 | i[474];
  assign N469 = N468 | i[475];
  assign N468 = N467 | i[476];
  assign N467 = N466 | i[477];
  assign N466 = N465 | i[478];
  assign N465 = N464 | i[479];
  assign N464 = N463 | i[480];
  assign N463 = N462 | i[481];
  assign N462 = N461 | i[482];
  assign N461 = N460 | i[483];
  assign N460 = N459 | i[484];
  assign N459 = N458 | i[485];
  assign N458 = N457 | i[486];
  assign N457 = N456 | i[487];
  assign N456 = N455 | i[488];
  assign N455 = N454 | i[489];
  assign N454 = N453 | i[490];
  assign N453 = N452 | i[491];
  assign N452 = N451 | i[492];
  assign N451 = N450 | i[493];
  assign N450 = N449 | i[494];
  assign N449 = N448 | i[495];
  assign N448 = N447 | i[496];
  assign N447 = N446 | i[497];
  assign N446 = N445 | i[498];
  assign N445 = N444 | i[499];
  assign N444 = N443 | i[500];
  assign N443 = N442 | i[501];
  assign N442 = N441 | i[502];
  assign N441 = N440 | i[503];
  assign N440 = N439 | i[504];
  assign N439 = N438 | i[505];
  assign N438 = N437 | i[506];
  assign N437 = N436 | i[507];
  assign N436 = N435 | i[508];
  assign N435 = N434 | i[509];
  assign N434 = i[511] | i[510];
  assign o[8] = N557 | i[512];
  assign N557 = N556 | i[513];
  assign N556 = N555 | i[514];
  assign N555 = N554 | i[515];
  assign N554 = N553 | i[516];
  assign N553 = N552 | i[517];
  assign N552 = N551 | i[518];
  assign N551 = N550 | i[519];
  assign N550 = N549 | i[520];
  assign N549 = N548 | i[521];
  assign N548 = N547 | i[522];
  assign N547 = N546 | i[523];
  assign N546 = N545 | i[524];
  assign N545 = N544 | i[525];
  assign N544 = N543 | i[526];
  assign N543 = N542 | i[527];
  assign N542 = N541 | i[528];
  assign N541 = N540 | i[529];
  assign N540 = N539 | i[530];
  assign N539 = N538 | i[531];
  assign N538 = N537 | i[532];
  assign N537 = N536 | i[533];
  assign N536 = N535 | i[534];
  assign N535 = N534 | i[535];
  assign N534 = N533 | i[536];
  assign N533 = N532 | i[537];
  assign N532 = N531 | i[538];
  assign N531 = N530 | i[539];
  assign N530 = N529 | i[540];
  assign N529 = N528 | i[541];
  assign N528 = N527 | i[542];
  assign N527 = N526 | i[543];
  assign N526 = N525 | i[544];
  assign N525 = N524 | i[545];
  assign N524 = N523 | i[546];
  assign N523 = N522 | i[547];
  assign N522 = N521 | i[548];
  assign N521 = N520 | i[549];
  assign N520 = N519 | i[550];
  assign N519 = N518 | i[551];
  assign N518 = N517 | i[552];
  assign N517 = N516 | i[553];
  assign N516 = N515 | i[554];
  assign N515 = N514 | i[555];
  assign N514 = N513 | i[556];
  assign N513 = N512 | i[557];
  assign N512 = N511 | i[558];
  assign N511 = N510 | i[559];
  assign N510 = N509 | i[560];
  assign N509 = N508 | i[561];
  assign N508 = N507 | i[562];
  assign N507 = N506 | i[563];
  assign N506 = N505 | i[564];
  assign N505 = N504 | i[565];
  assign N504 = N503 | i[566];
  assign N503 = N502 | i[567];
  assign N502 = N501 | i[568];
  assign N501 = N500 | i[569];
  assign N500 = N499 | i[570];
  assign N499 = N498 | i[571];
  assign N498 = N497 | i[572];
  assign N497 = N496 | i[573];
  assign N496 = i[575] | i[574];
  assign o[9] = N619 | i[576];
  assign N619 = N618 | i[577];
  assign N618 = N617 | i[578];
  assign N617 = N616 | i[579];
  assign N616 = N615 | i[580];
  assign N615 = N614 | i[581];
  assign N614 = N613 | i[582];
  assign N613 = N612 | i[583];
  assign N612 = N611 | i[584];
  assign N611 = N610 | i[585];
  assign N610 = N609 | i[586];
  assign N609 = N608 | i[587];
  assign N608 = N607 | i[588];
  assign N607 = N606 | i[589];
  assign N606 = N605 | i[590];
  assign N605 = N604 | i[591];
  assign N604 = N603 | i[592];
  assign N603 = N602 | i[593];
  assign N602 = N601 | i[594];
  assign N601 = N600 | i[595];
  assign N600 = N599 | i[596];
  assign N599 = N598 | i[597];
  assign N598 = N597 | i[598];
  assign N597 = N596 | i[599];
  assign N596 = N595 | i[600];
  assign N595 = N594 | i[601];
  assign N594 = N593 | i[602];
  assign N593 = N592 | i[603];
  assign N592 = N591 | i[604];
  assign N591 = N590 | i[605];
  assign N590 = N589 | i[606];
  assign N589 = N588 | i[607];
  assign N588 = N587 | i[608];
  assign N587 = N586 | i[609];
  assign N586 = N585 | i[610];
  assign N585 = N584 | i[611];
  assign N584 = N583 | i[612];
  assign N583 = N582 | i[613];
  assign N582 = N581 | i[614];
  assign N581 = N580 | i[615];
  assign N580 = N579 | i[616];
  assign N579 = N578 | i[617];
  assign N578 = N577 | i[618];
  assign N577 = N576 | i[619];
  assign N576 = N575 | i[620];
  assign N575 = N574 | i[621];
  assign N574 = N573 | i[622];
  assign N573 = N572 | i[623];
  assign N572 = N571 | i[624];
  assign N571 = N570 | i[625];
  assign N570 = N569 | i[626];
  assign N569 = N568 | i[627];
  assign N568 = N567 | i[628];
  assign N567 = N566 | i[629];
  assign N566 = N565 | i[630];
  assign N565 = N564 | i[631];
  assign N564 = N563 | i[632];
  assign N563 = N562 | i[633];
  assign N562 = N561 | i[634];
  assign N561 = N560 | i[635];
  assign N560 = N559 | i[636];
  assign N559 = N558 | i[637];
  assign N558 = i[639] | i[638];

endmodule

