

module top
(
  i,
  o
);

  input [2559:0] i;
  output [19:0] o;

  bsg_reduce_segmented
  wrapper
  (
    .i(i),
    .o(o)
  );


endmodule



module bsg_reduce_segmented
(
  i,
  o
);

  input [2559:0] i;
  output [19:0] o;
  wire [19:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,
  N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,
  N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
  N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,
  N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,
  N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,
  N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,
  N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,
  N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,
  N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,
  N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,
  N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,
  N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,
  N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,
  N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,
  N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,
  N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539;
  assign o[0] = ~N126;
  assign N126 = N125 | i[0];
  assign N125 = N124 | i[1];
  assign N124 = N123 | i[2];
  assign N123 = N122 | i[3];
  assign N122 = N121 | i[4];
  assign N121 = N120 | i[5];
  assign N120 = N119 | i[6];
  assign N119 = N118 | i[7];
  assign N118 = N117 | i[8];
  assign N117 = N116 | i[9];
  assign N116 = N115 | i[10];
  assign N115 = N114 | i[11];
  assign N114 = N113 | i[12];
  assign N113 = N112 | i[13];
  assign N112 = N111 | i[14];
  assign N111 = N110 | i[15];
  assign N110 = N109 | i[16];
  assign N109 = N108 | i[17];
  assign N108 = N107 | i[18];
  assign N107 = N106 | i[19];
  assign N106 = N105 | i[20];
  assign N105 = N104 | i[21];
  assign N104 = N103 | i[22];
  assign N103 = N102 | i[23];
  assign N102 = N101 | i[24];
  assign N101 = N100 | i[25];
  assign N100 = N99 | i[26];
  assign N99 = N98 | i[27];
  assign N98 = N97 | i[28];
  assign N97 = N96 | i[29];
  assign N96 = N95 | i[30];
  assign N95 = N94 | i[31];
  assign N94 = N93 | i[32];
  assign N93 = N92 | i[33];
  assign N92 = N91 | i[34];
  assign N91 = N90 | i[35];
  assign N90 = N89 | i[36];
  assign N89 = N88 | i[37];
  assign N88 = N87 | i[38];
  assign N87 = N86 | i[39];
  assign N86 = N85 | i[40];
  assign N85 = N84 | i[41];
  assign N84 = N83 | i[42];
  assign N83 = N82 | i[43];
  assign N82 = N81 | i[44];
  assign N81 = N80 | i[45];
  assign N80 = N79 | i[46];
  assign N79 = N78 | i[47];
  assign N78 = N77 | i[48];
  assign N77 = N76 | i[49];
  assign N76 = N75 | i[50];
  assign N75 = N74 | i[51];
  assign N74 = N73 | i[52];
  assign N73 = N72 | i[53];
  assign N72 = N71 | i[54];
  assign N71 = N70 | i[55];
  assign N70 = N69 | i[56];
  assign N69 = N68 | i[57];
  assign N68 = N67 | i[58];
  assign N67 = N66 | i[59];
  assign N66 = N65 | i[60];
  assign N65 = N64 | i[61];
  assign N64 = N63 | i[62];
  assign N63 = N62 | i[63];
  assign N62 = N61 | i[64];
  assign N61 = N60 | i[65];
  assign N60 = N59 | i[66];
  assign N59 = N58 | i[67];
  assign N58 = N57 | i[68];
  assign N57 = N56 | i[69];
  assign N56 = N55 | i[70];
  assign N55 = N54 | i[71];
  assign N54 = N53 | i[72];
  assign N53 = N52 | i[73];
  assign N52 = N51 | i[74];
  assign N51 = N50 | i[75];
  assign N50 = N49 | i[76];
  assign N49 = N48 | i[77];
  assign N48 = N47 | i[78];
  assign N47 = N46 | i[79];
  assign N46 = N45 | i[80];
  assign N45 = N44 | i[81];
  assign N44 = N43 | i[82];
  assign N43 = N42 | i[83];
  assign N42 = N41 | i[84];
  assign N41 = N40 | i[85];
  assign N40 = N39 | i[86];
  assign N39 = N38 | i[87];
  assign N38 = N37 | i[88];
  assign N37 = N36 | i[89];
  assign N36 = N35 | i[90];
  assign N35 = N34 | i[91];
  assign N34 = N33 | i[92];
  assign N33 = N32 | i[93];
  assign N32 = N31 | i[94];
  assign N31 = N30 | i[95];
  assign N30 = N29 | i[96];
  assign N29 = N28 | i[97];
  assign N28 = N27 | i[98];
  assign N27 = N26 | i[99];
  assign N26 = N25 | i[100];
  assign N25 = N24 | i[101];
  assign N24 = N23 | i[102];
  assign N23 = N22 | i[103];
  assign N22 = N21 | i[104];
  assign N21 = N20 | i[105];
  assign N20 = N19 | i[106];
  assign N19 = N18 | i[107];
  assign N18 = N17 | i[108];
  assign N17 = N16 | i[109];
  assign N16 = N15 | i[110];
  assign N15 = N14 | i[111];
  assign N14 = N13 | i[112];
  assign N13 = N12 | i[113];
  assign N12 = N11 | i[114];
  assign N11 = N10 | i[115];
  assign N10 = N9 | i[116];
  assign N9 = N8 | i[117];
  assign N8 = N7 | i[118];
  assign N7 = N6 | i[119];
  assign N6 = N5 | i[120];
  assign N5 = N4 | i[121];
  assign N4 = N3 | i[122];
  assign N3 = N2 | i[123];
  assign N2 = N1 | i[124];
  assign N1 = N0 | i[125];
  assign N0 = i[127] | i[126];
  assign o[1] = ~N253;
  assign N253 = N252 | i[128];
  assign N252 = N251 | i[129];
  assign N251 = N250 | i[130];
  assign N250 = N249 | i[131];
  assign N249 = N248 | i[132];
  assign N248 = N247 | i[133];
  assign N247 = N246 | i[134];
  assign N246 = N245 | i[135];
  assign N245 = N244 | i[136];
  assign N244 = N243 | i[137];
  assign N243 = N242 | i[138];
  assign N242 = N241 | i[139];
  assign N241 = N240 | i[140];
  assign N240 = N239 | i[141];
  assign N239 = N238 | i[142];
  assign N238 = N237 | i[143];
  assign N237 = N236 | i[144];
  assign N236 = N235 | i[145];
  assign N235 = N234 | i[146];
  assign N234 = N233 | i[147];
  assign N233 = N232 | i[148];
  assign N232 = N231 | i[149];
  assign N231 = N230 | i[150];
  assign N230 = N229 | i[151];
  assign N229 = N228 | i[152];
  assign N228 = N227 | i[153];
  assign N227 = N226 | i[154];
  assign N226 = N225 | i[155];
  assign N225 = N224 | i[156];
  assign N224 = N223 | i[157];
  assign N223 = N222 | i[158];
  assign N222 = N221 | i[159];
  assign N221 = N220 | i[160];
  assign N220 = N219 | i[161];
  assign N219 = N218 | i[162];
  assign N218 = N217 | i[163];
  assign N217 = N216 | i[164];
  assign N216 = N215 | i[165];
  assign N215 = N214 | i[166];
  assign N214 = N213 | i[167];
  assign N213 = N212 | i[168];
  assign N212 = N211 | i[169];
  assign N211 = N210 | i[170];
  assign N210 = N209 | i[171];
  assign N209 = N208 | i[172];
  assign N208 = N207 | i[173];
  assign N207 = N206 | i[174];
  assign N206 = N205 | i[175];
  assign N205 = N204 | i[176];
  assign N204 = N203 | i[177];
  assign N203 = N202 | i[178];
  assign N202 = N201 | i[179];
  assign N201 = N200 | i[180];
  assign N200 = N199 | i[181];
  assign N199 = N198 | i[182];
  assign N198 = N197 | i[183];
  assign N197 = N196 | i[184];
  assign N196 = N195 | i[185];
  assign N195 = N194 | i[186];
  assign N194 = N193 | i[187];
  assign N193 = N192 | i[188];
  assign N192 = N191 | i[189];
  assign N191 = N190 | i[190];
  assign N190 = N189 | i[191];
  assign N189 = N188 | i[192];
  assign N188 = N187 | i[193];
  assign N187 = N186 | i[194];
  assign N186 = N185 | i[195];
  assign N185 = N184 | i[196];
  assign N184 = N183 | i[197];
  assign N183 = N182 | i[198];
  assign N182 = N181 | i[199];
  assign N181 = N180 | i[200];
  assign N180 = N179 | i[201];
  assign N179 = N178 | i[202];
  assign N178 = N177 | i[203];
  assign N177 = N176 | i[204];
  assign N176 = N175 | i[205];
  assign N175 = N174 | i[206];
  assign N174 = N173 | i[207];
  assign N173 = N172 | i[208];
  assign N172 = N171 | i[209];
  assign N171 = N170 | i[210];
  assign N170 = N169 | i[211];
  assign N169 = N168 | i[212];
  assign N168 = N167 | i[213];
  assign N167 = N166 | i[214];
  assign N166 = N165 | i[215];
  assign N165 = N164 | i[216];
  assign N164 = N163 | i[217];
  assign N163 = N162 | i[218];
  assign N162 = N161 | i[219];
  assign N161 = N160 | i[220];
  assign N160 = N159 | i[221];
  assign N159 = N158 | i[222];
  assign N158 = N157 | i[223];
  assign N157 = N156 | i[224];
  assign N156 = N155 | i[225];
  assign N155 = N154 | i[226];
  assign N154 = N153 | i[227];
  assign N153 = N152 | i[228];
  assign N152 = N151 | i[229];
  assign N151 = N150 | i[230];
  assign N150 = N149 | i[231];
  assign N149 = N148 | i[232];
  assign N148 = N147 | i[233];
  assign N147 = N146 | i[234];
  assign N146 = N145 | i[235];
  assign N145 = N144 | i[236];
  assign N144 = N143 | i[237];
  assign N143 = N142 | i[238];
  assign N142 = N141 | i[239];
  assign N141 = N140 | i[240];
  assign N140 = N139 | i[241];
  assign N139 = N138 | i[242];
  assign N138 = N137 | i[243];
  assign N137 = N136 | i[244];
  assign N136 = N135 | i[245];
  assign N135 = N134 | i[246];
  assign N134 = N133 | i[247];
  assign N133 = N132 | i[248];
  assign N132 = N131 | i[249];
  assign N131 = N130 | i[250];
  assign N130 = N129 | i[251];
  assign N129 = N128 | i[252];
  assign N128 = N127 | i[253];
  assign N127 = i[255] | i[254];
  assign o[2] = ~N380;
  assign N380 = N379 | i[256];
  assign N379 = N378 | i[257];
  assign N378 = N377 | i[258];
  assign N377 = N376 | i[259];
  assign N376 = N375 | i[260];
  assign N375 = N374 | i[261];
  assign N374 = N373 | i[262];
  assign N373 = N372 | i[263];
  assign N372 = N371 | i[264];
  assign N371 = N370 | i[265];
  assign N370 = N369 | i[266];
  assign N369 = N368 | i[267];
  assign N368 = N367 | i[268];
  assign N367 = N366 | i[269];
  assign N366 = N365 | i[270];
  assign N365 = N364 | i[271];
  assign N364 = N363 | i[272];
  assign N363 = N362 | i[273];
  assign N362 = N361 | i[274];
  assign N361 = N360 | i[275];
  assign N360 = N359 | i[276];
  assign N359 = N358 | i[277];
  assign N358 = N357 | i[278];
  assign N357 = N356 | i[279];
  assign N356 = N355 | i[280];
  assign N355 = N354 | i[281];
  assign N354 = N353 | i[282];
  assign N353 = N352 | i[283];
  assign N352 = N351 | i[284];
  assign N351 = N350 | i[285];
  assign N350 = N349 | i[286];
  assign N349 = N348 | i[287];
  assign N348 = N347 | i[288];
  assign N347 = N346 | i[289];
  assign N346 = N345 | i[290];
  assign N345 = N344 | i[291];
  assign N344 = N343 | i[292];
  assign N343 = N342 | i[293];
  assign N342 = N341 | i[294];
  assign N341 = N340 | i[295];
  assign N340 = N339 | i[296];
  assign N339 = N338 | i[297];
  assign N338 = N337 | i[298];
  assign N337 = N336 | i[299];
  assign N336 = N335 | i[300];
  assign N335 = N334 | i[301];
  assign N334 = N333 | i[302];
  assign N333 = N332 | i[303];
  assign N332 = N331 | i[304];
  assign N331 = N330 | i[305];
  assign N330 = N329 | i[306];
  assign N329 = N328 | i[307];
  assign N328 = N327 | i[308];
  assign N327 = N326 | i[309];
  assign N326 = N325 | i[310];
  assign N325 = N324 | i[311];
  assign N324 = N323 | i[312];
  assign N323 = N322 | i[313];
  assign N322 = N321 | i[314];
  assign N321 = N320 | i[315];
  assign N320 = N319 | i[316];
  assign N319 = N318 | i[317];
  assign N318 = N317 | i[318];
  assign N317 = N316 | i[319];
  assign N316 = N315 | i[320];
  assign N315 = N314 | i[321];
  assign N314 = N313 | i[322];
  assign N313 = N312 | i[323];
  assign N312 = N311 | i[324];
  assign N311 = N310 | i[325];
  assign N310 = N309 | i[326];
  assign N309 = N308 | i[327];
  assign N308 = N307 | i[328];
  assign N307 = N306 | i[329];
  assign N306 = N305 | i[330];
  assign N305 = N304 | i[331];
  assign N304 = N303 | i[332];
  assign N303 = N302 | i[333];
  assign N302 = N301 | i[334];
  assign N301 = N300 | i[335];
  assign N300 = N299 | i[336];
  assign N299 = N298 | i[337];
  assign N298 = N297 | i[338];
  assign N297 = N296 | i[339];
  assign N296 = N295 | i[340];
  assign N295 = N294 | i[341];
  assign N294 = N293 | i[342];
  assign N293 = N292 | i[343];
  assign N292 = N291 | i[344];
  assign N291 = N290 | i[345];
  assign N290 = N289 | i[346];
  assign N289 = N288 | i[347];
  assign N288 = N287 | i[348];
  assign N287 = N286 | i[349];
  assign N286 = N285 | i[350];
  assign N285 = N284 | i[351];
  assign N284 = N283 | i[352];
  assign N283 = N282 | i[353];
  assign N282 = N281 | i[354];
  assign N281 = N280 | i[355];
  assign N280 = N279 | i[356];
  assign N279 = N278 | i[357];
  assign N278 = N277 | i[358];
  assign N277 = N276 | i[359];
  assign N276 = N275 | i[360];
  assign N275 = N274 | i[361];
  assign N274 = N273 | i[362];
  assign N273 = N272 | i[363];
  assign N272 = N271 | i[364];
  assign N271 = N270 | i[365];
  assign N270 = N269 | i[366];
  assign N269 = N268 | i[367];
  assign N268 = N267 | i[368];
  assign N267 = N266 | i[369];
  assign N266 = N265 | i[370];
  assign N265 = N264 | i[371];
  assign N264 = N263 | i[372];
  assign N263 = N262 | i[373];
  assign N262 = N261 | i[374];
  assign N261 = N260 | i[375];
  assign N260 = N259 | i[376];
  assign N259 = N258 | i[377];
  assign N258 = N257 | i[378];
  assign N257 = N256 | i[379];
  assign N256 = N255 | i[380];
  assign N255 = N254 | i[381];
  assign N254 = i[383] | i[382];
  assign o[3] = ~N507;
  assign N507 = N506 | i[384];
  assign N506 = N505 | i[385];
  assign N505 = N504 | i[386];
  assign N504 = N503 | i[387];
  assign N503 = N502 | i[388];
  assign N502 = N501 | i[389];
  assign N501 = N500 | i[390];
  assign N500 = N499 | i[391];
  assign N499 = N498 | i[392];
  assign N498 = N497 | i[393];
  assign N497 = N496 | i[394];
  assign N496 = N495 | i[395];
  assign N495 = N494 | i[396];
  assign N494 = N493 | i[397];
  assign N493 = N492 | i[398];
  assign N492 = N491 | i[399];
  assign N491 = N490 | i[400];
  assign N490 = N489 | i[401];
  assign N489 = N488 | i[402];
  assign N488 = N487 | i[403];
  assign N487 = N486 | i[404];
  assign N486 = N485 | i[405];
  assign N485 = N484 | i[406];
  assign N484 = N483 | i[407];
  assign N483 = N482 | i[408];
  assign N482 = N481 | i[409];
  assign N481 = N480 | i[410];
  assign N480 = N479 | i[411];
  assign N479 = N478 | i[412];
  assign N478 = N477 | i[413];
  assign N477 = N476 | i[414];
  assign N476 = N475 | i[415];
  assign N475 = N474 | i[416];
  assign N474 = N473 | i[417];
  assign N473 = N472 | i[418];
  assign N472 = N471 | i[419];
  assign N471 = N470 | i[420];
  assign N470 = N469 | i[421];
  assign N469 = N468 | i[422];
  assign N468 = N467 | i[423];
  assign N467 = N466 | i[424];
  assign N466 = N465 | i[425];
  assign N465 = N464 | i[426];
  assign N464 = N463 | i[427];
  assign N463 = N462 | i[428];
  assign N462 = N461 | i[429];
  assign N461 = N460 | i[430];
  assign N460 = N459 | i[431];
  assign N459 = N458 | i[432];
  assign N458 = N457 | i[433];
  assign N457 = N456 | i[434];
  assign N456 = N455 | i[435];
  assign N455 = N454 | i[436];
  assign N454 = N453 | i[437];
  assign N453 = N452 | i[438];
  assign N452 = N451 | i[439];
  assign N451 = N450 | i[440];
  assign N450 = N449 | i[441];
  assign N449 = N448 | i[442];
  assign N448 = N447 | i[443];
  assign N447 = N446 | i[444];
  assign N446 = N445 | i[445];
  assign N445 = N444 | i[446];
  assign N444 = N443 | i[447];
  assign N443 = N442 | i[448];
  assign N442 = N441 | i[449];
  assign N441 = N440 | i[450];
  assign N440 = N439 | i[451];
  assign N439 = N438 | i[452];
  assign N438 = N437 | i[453];
  assign N437 = N436 | i[454];
  assign N436 = N435 | i[455];
  assign N435 = N434 | i[456];
  assign N434 = N433 | i[457];
  assign N433 = N432 | i[458];
  assign N432 = N431 | i[459];
  assign N431 = N430 | i[460];
  assign N430 = N429 | i[461];
  assign N429 = N428 | i[462];
  assign N428 = N427 | i[463];
  assign N427 = N426 | i[464];
  assign N426 = N425 | i[465];
  assign N425 = N424 | i[466];
  assign N424 = N423 | i[467];
  assign N423 = N422 | i[468];
  assign N422 = N421 | i[469];
  assign N421 = N420 | i[470];
  assign N420 = N419 | i[471];
  assign N419 = N418 | i[472];
  assign N418 = N417 | i[473];
  assign N417 = N416 | i[474];
  assign N416 = N415 | i[475];
  assign N415 = N414 | i[476];
  assign N414 = N413 | i[477];
  assign N413 = N412 | i[478];
  assign N412 = N411 | i[479];
  assign N411 = N410 | i[480];
  assign N410 = N409 | i[481];
  assign N409 = N408 | i[482];
  assign N408 = N407 | i[483];
  assign N407 = N406 | i[484];
  assign N406 = N405 | i[485];
  assign N405 = N404 | i[486];
  assign N404 = N403 | i[487];
  assign N403 = N402 | i[488];
  assign N402 = N401 | i[489];
  assign N401 = N400 | i[490];
  assign N400 = N399 | i[491];
  assign N399 = N398 | i[492];
  assign N398 = N397 | i[493];
  assign N397 = N396 | i[494];
  assign N396 = N395 | i[495];
  assign N395 = N394 | i[496];
  assign N394 = N393 | i[497];
  assign N393 = N392 | i[498];
  assign N392 = N391 | i[499];
  assign N391 = N390 | i[500];
  assign N390 = N389 | i[501];
  assign N389 = N388 | i[502];
  assign N388 = N387 | i[503];
  assign N387 = N386 | i[504];
  assign N386 = N385 | i[505];
  assign N385 = N384 | i[506];
  assign N384 = N383 | i[507];
  assign N383 = N382 | i[508];
  assign N382 = N381 | i[509];
  assign N381 = i[511] | i[510];
  assign o[4] = ~N634;
  assign N634 = N633 | i[512];
  assign N633 = N632 | i[513];
  assign N632 = N631 | i[514];
  assign N631 = N630 | i[515];
  assign N630 = N629 | i[516];
  assign N629 = N628 | i[517];
  assign N628 = N627 | i[518];
  assign N627 = N626 | i[519];
  assign N626 = N625 | i[520];
  assign N625 = N624 | i[521];
  assign N624 = N623 | i[522];
  assign N623 = N622 | i[523];
  assign N622 = N621 | i[524];
  assign N621 = N620 | i[525];
  assign N620 = N619 | i[526];
  assign N619 = N618 | i[527];
  assign N618 = N617 | i[528];
  assign N617 = N616 | i[529];
  assign N616 = N615 | i[530];
  assign N615 = N614 | i[531];
  assign N614 = N613 | i[532];
  assign N613 = N612 | i[533];
  assign N612 = N611 | i[534];
  assign N611 = N610 | i[535];
  assign N610 = N609 | i[536];
  assign N609 = N608 | i[537];
  assign N608 = N607 | i[538];
  assign N607 = N606 | i[539];
  assign N606 = N605 | i[540];
  assign N605 = N604 | i[541];
  assign N604 = N603 | i[542];
  assign N603 = N602 | i[543];
  assign N602 = N601 | i[544];
  assign N601 = N600 | i[545];
  assign N600 = N599 | i[546];
  assign N599 = N598 | i[547];
  assign N598 = N597 | i[548];
  assign N597 = N596 | i[549];
  assign N596 = N595 | i[550];
  assign N595 = N594 | i[551];
  assign N594 = N593 | i[552];
  assign N593 = N592 | i[553];
  assign N592 = N591 | i[554];
  assign N591 = N590 | i[555];
  assign N590 = N589 | i[556];
  assign N589 = N588 | i[557];
  assign N588 = N587 | i[558];
  assign N587 = N586 | i[559];
  assign N586 = N585 | i[560];
  assign N585 = N584 | i[561];
  assign N584 = N583 | i[562];
  assign N583 = N582 | i[563];
  assign N582 = N581 | i[564];
  assign N581 = N580 | i[565];
  assign N580 = N579 | i[566];
  assign N579 = N578 | i[567];
  assign N578 = N577 | i[568];
  assign N577 = N576 | i[569];
  assign N576 = N575 | i[570];
  assign N575 = N574 | i[571];
  assign N574 = N573 | i[572];
  assign N573 = N572 | i[573];
  assign N572 = N571 | i[574];
  assign N571 = N570 | i[575];
  assign N570 = N569 | i[576];
  assign N569 = N568 | i[577];
  assign N568 = N567 | i[578];
  assign N567 = N566 | i[579];
  assign N566 = N565 | i[580];
  assign N565 = N564 | i[581];
  assign N564 = N563 | i[582];
  assign N563 = N562 | i[583];
  assign N562 = N561 | i[584];
  assign N561 = N560 | i[585];
  assign N560 = N559 | i[586];
  assign N559 = N558 | i[587];
  assign N558 = N557 | i[588];
  assign N557 = N556 | i[589];
  assign N556 = N555 | i[590];
  assign N555 = N554 | i[591];
  assign N554 = N553 | i[592];
  assign N553 = N552 | i[593];
  assign N552 = N551 | i[594];
  assign N551 = N550 | i[595];
  assign N550 = N549 | i[596];
  assign N549 = N548 | i[597];
  assign N548 = N547 | i[598];
  assign N547 = N546 | i[599];
  assign N546 = N545 | i[600];
  assign N545 = N544 | i[601];
  assign N544 = N543 | i[602];
  assign N543 = N542 | i[603];
  assign N542 = N541 | i[604];
  assign N541 = N540 | i[605];
  assign N540 = N539 | i[606];
  assign N539 = N538 | i[607];
  assign N538 = N537 | i[608];
  assign N537 = N536 | i[609];
  assign N536 = N535 | i[610];
  assign N535 = N534 | i[611];
  assign N534 = N533 | i[612];
  assign N533 = N532 | i[613];
  assign N532 = N531 | i[614];
  assign N531 = N530 | i[615];
  assign N530 = N529 | i[616];
  assign N529 = N528 | i[617];
  assign N528 = N527 | i[618];
  assign N527 = N526 | i[619];
  assign N526 = N525 | i[620];
  assign N525 = N524 | i[621];
  assign N524 = N523 | i[622];
  assign N523 = N522 | i[623];
  assign N522 = N521 | i[624];
  assign N521 = N520 | i[625];
  assign N520 = N519 | i[626];
  assign N519 = N518 | i[627];
  assign N518 = N517 | i[628];
  assign N517 = N516 | i[629];
  assign N516 = N515 | i[630];
  assign N515 = N514 | i[631];
  assign N514 = N513 | i[632];
  assign N513 = N512 | i[633];
  assign N512 = N511 | i[634];
  assign N511 = N510 | i[635];
  assign N510 = N509 | i[636];
  assign N509 = N508 | i[637];
  assign N508 = i[639] | i[638];
  assign o[5] = ~N761;
  assign N761 = N760 | i[640];
  assign N760 = N759 | i[641];
  assign N759 = N758 | i[642];
  assign N758 = N757 | i[643];
  assign N757 = N756 | i[644];
  assign N756 = N755 | i[645];
  assign N755 = N754 | i[646];
  assign N754 = N753 | i[647];
  assign N753 = N752 | i[648];
  assign N752 = N751 | i[649];
  assign N751 = N750 | i[650];
  assign N750 = N749 | i[651];
  assign N749 = N748 | i[652];
  assign N748 = N747 | i[653];
  assign N747 = N746 | i[654];
  assign N746 = N745 | i[655];
  assign N745 = N744 | i[656];
  assign N744 = N743 | i[657];
  assign N743 = N742 | i[658];
  assign N742 = N741 | i[659];
  assign N741 = N740 | i[660];
  assign N740 = N739 | i[661];
  assign N739 = N738 | i[662];
  assign N738 = N737 | i[663];
  assign N737 = N736 | i[664];
  assign N736 = N735 | i[665];
  assign N735 = N734 | i[666];
  assign N734 = N733 | i[667];
  assign N733 = N732 | i[668];
  assign N732 = N731 | i[669];
  assign N731 = N730 | i[670];
  assign N730 = N729 | i[671];
  assign N729 = N728 | i[672];
  assign N728 = N727 | i[673];
  assign N727 = N726 | i[674];
  assign N726 = N725 | i[675];
  assign N725 = N724 | i[676];
  assign N724 = N723 | i[677];
  assign N723 = N722 | i[678];
  assign N722 = N721 | i[679];
  assign N721 = N720 | i[680];
  assign N720 = N719 | i[681];
  assign N719 = N718 | i[682];
  assign N718 = N717 | i[683];
  assign N717 = N716 | i[684];
  assign N716 = N715 | i[685];
  assign N715 = N714 | i[686];
  assign N714 = N713 | i[687];
  assign N713 = N712 | i[688];
  assign N712 = N711 | i[689];
  assign N711 = N710 | i[690];
  assign N710 = N709 | i[691];
  assign N709 = N708 | i[692];
  assign N708 = N707 | i[693];
  assign N707 = N706 | i[694];
  assign N706 = N705 | i[695];
  assign N705 = N704 | i[696];
  assign N704 = N703 | i[697];
  assign N703 = N702 | i[698];
  assign N702 = N701 | i[699];
  assign N701 = N700 | i[700];
  assign N700 = N699 | i[701];
  assign N699 = N698 | i[702];
  assign N698 = N697 | i[703];
  assign N697 = N696 | i[704];
  assign N696 = N695 | i[705];
  assign N695 = N694 | i[706];
  assign N694 = N693 | i[707];
  assign N693 = N692 | i[708];
  assign N692 = N691 | i[709];
  assign N691 = N690 | i[710];
  assign N690 = N689 | i[711];
  assign N689 = N688 | i[712];
  assign N688 = N687 | i[713];
  assign N687 = N686 | i[714];
  assign N686 = N685 | i[715];
  assign N685 = N684 | i[716];
  assign N684 = N683 | i[717];
  assign N683 = N682 | i[718];
  assign N682 = N681 | i[719];
  assign N681 = N680 | i[720];
  assign N680 = N679 | i[721];
  assign N679 = N678 | i[722];
  assign N678 = N677 | i[723];
  assign N677 = N676 | i[724];
  assign N676 = N675 | i[725];
  assign N675 = N674 | i[726];
  assign N674 = N673 | i[727];
  assign N673 = N672 | i[728];
  assign N672 = N671 | i[729];
  assign N671 = N670 | i[730];
  assign N670 = N669 | i[731];
  assign N669 = N668 | i[732];
  assign N668 = N667 | i[733];
  assign N667 = N666 | i[734];
  assign N666 = N665 | i[735];
  assign N665 = N664 | i[736];
  assign N664 = N663 | i[737];
  assign N663 = N662 | i[738];
  assign N662 = N661 | i[739];
  assign N661 = N660 | i[740];
  assign N660 = N659 | i[741];
  assign N659 = N658 | i[742];
  assign N658 = N657 | i[743];
  assign N657 = N656 | i[744];
  assign N656 = N655 | i[745];
  assign N655 = N654 | i[746];
  assign N654 = N653 | i[747];
  assign N653 = N652 | i[748];
  assign N652 = N651 | i[749];
  assign N651 = N650 | i[750];
  assign N650 = N649 | i[751];
  assign N649 = N648 | i[752];
  assign N648 = N647 | i[753];
  assign N647 = N646 | i[754];
  assign N646 = N645 | i[755];
  assign N645 = N644 | i[756];
  assign N644 = N643 | i[757];
  assign N643 = N642 | i[758];
  assign N642 = N641 | i[759];
  assign N641 = N640 | i[760];
  assign N640 = N639 | i[761];
  assign N639 = N638 | i[762];
  assign N638 = N637 | i[763];
  assign N637 = N636 | i[764];
  assign N636 = N635 | i[765];
  assign N635 = i[767] | i[766];
  assign o[6] = ~N888;
  assign N888 = N887 | i[768];
  assign N887 = N886 | i[769];
  assign N886 = N885 | i[770];
  assign N885 = N884 | i[771];
  assign N884 = N883 | i[772];
  assign N883 = N882 | i[773];
  assign N882 = N881 | i[774];
  assign N881 = N880 | i[775];
  assign N880 = N879 | i[776];
  assign N879 = N878 | i[777];
  assign N878 = N877 | i[778];
  assign N877 = N876 | i[779];
  assign N876 = N875 | i[780];
  assign N875 = N874 | i[781];
  assign N874 = N873 | i[782];
  assign N873 = N872 | i[783];
  assign N872 = N871 | i[784];
  assign N871 = N870 | i[785];
  assign N870 = N869 | i[786];
  assign N869 = N868 | i[787];
  assign N868 = N867 | i[788];
  assign N867 = N866 | i[789];
  assign N866 = N865 | i[790];
  assign N865 = N864 | i[791];
  assign N864 = N863 | i[792];
  assign N863 = N862 | i[793];
  assign N862 = N861 | i[794];
  assign N861 = N860 | i[795];
  assign N860 = N859 | i[796];
  assign N859 = N858 | i[797];
  assign N858 = N857 | i[798];
  assign N857 = N856 | i[799];
  assign N856 = N855 | i[800];
  assign N855 = N854 | i[801];
  assign N854 = N853 | i[802];
  assign N853 = N852 | i[803];
  assign N852 = N851 | i[804];
  assign N851 = N850 | i[805];
  assign N850 = N849 | i[806];
  assign N849 = N848 | i[807];
  assign N848 = N847 | i[808];
  assign N847 = N846 | i[809];
  assign N846 = N845 | i[810];
  assign N845 = N844 | i[811];
  assign N844 = N843 | i[812];
  assign N843 = N842 | i[813];
  assign N842 = N841 | i[814];
  assign N841 = N840 | i[815];
  assign N840 = N839 | i[816];
  assign N839 = N838 | i[817];
  assign N838 = N837 | i[818];
  assign N837 = N836 | i[819];
  assign N836 = N835 | i[820];
  assign N835 = N834 | i[821];
  assign N834 = N833 | i[822];
  assign N833 = N832 | i[823];
  assign N832 = N831 | i[824];
  assign N831 = N830 | i[825];
  assign N830 = N829 | i[826];
  assign N829 = N828 | i[827];
  assign N828 = N827 | i[828];
  assign N827 = N826 | i[829];
  assign N826 = N825 | i[830];
  assign N825 = N824 | i[831];
  assign N824 = N823 | i[832];
  assign N823 = N822 | i[833];
  assign N822 = N821 | i[834];
  assign N821 = N820 | i[835];
  assign N820 = N819 | i[836];
  assign N819 = N818 | i[837];
  assign N818 = N817 | i[838];
  assign N817 = N816 | i[839];
  assign N816 = N815 | i[840];
  assign N815 = N814 | i[841];
  assign N814 = N813 | i[842];
  assign N813 = N812 | i[843];
  assign N812 = N811 | i[844];
  assign N811 = N810 | i[845];
  assign N810 = N809 | i[846];
  assign N809 = N808 | i[847];
  assign N808 = N807 | i[848];
  assign N807 = N806 | i[849];
  assign N806 = N805 | i[850];
  assign N805 = N804 | i[851];
  assign N804 = N803 | i[852];
  assign N803 = N802 | i[853];
  assign N802 = N801 | i[854];
  assign N801 = N800 | i[855];
  assign N800 = N799 | i[856];
  assign N799 = N798 | i[857];
  assign N798 = N797 | i[858];
  assign N797 = N796 | i[859];
  assign N796 = N795 | i[860];
  assign N795 = N794 | i[861];
  assign N794 = N793 | i[862];
  assign N793 = N792 | i[863];
  assign N792 = N791 | i[864];
  assign N791 = N790 | i[865];
  assign N790 = N789 | i[866];
  assign N789 = N788 | i[867];
  assign N788 = N787 | i[868];
  assign N787 = N786 | i[869];
  assign N786 = N785 | i[870];
  assign N785 = N784 | i[871];
  assign N784 = N783 | i[872];
  assign N783 = N782 | i[873];
  assign N782 = N781 | i[874];
  assign N781 = N780 | i[875];
  assign N780 = N779 | i[876];
  assign N779 = N778 | i[877];
  assign N778 = N777 | i[878];
  assign N777 = N776 | i[879];
  assign N776 = N775 | i[880];
  assign N775 = N774 | i[881];
  assign N774 = N773 | i[882];
  assign N773 = N772 | i[883];
  assign N772 = N771 | i[884];
  assign N771 = N770 | i[885];
  assign N770 = N769 | i[886];
  assign N769 = N768 | i[887];
  assign N768 = N767 | i[888];
  assign N767 = N766 | i[889];
  assign N766 = N765 | i[890];
  assign N765 = N764 | i[891];
  assign N764 = N763 | i[892];
  assign N763 = N762 | i[893];
  assign N762 = i[895] | i[894];
  assign o[7] = ~N1015;
  assign N1015 = N1014 | i[896];
  assign N1014 = N1013 | i[897];
  assign N1013 = N1012 | i[898];
  assign N1012 = N1011 | i[899];
  assign N1011 = N1010 | i[900];
  assign N1010 = N1009 | i[901];
  assign N1009 = N1008 | i[902];
  assign N1008 = N1007 | i[903];
  assign N1007 = N1006 | i[904];
  assign N1006 = N1005 | i[905];
  assign N1005 = N1004 | i[906];
  assign N1004 = N1003 | i[907];
  assign N1003 = N1002 | i[908];
  assign N1002 = N1001 | i[909];
  assign N1001 = N1000 | i[910];
  assign N1000 = N999 | i[911];
  assign N999 = N998 | i[912];
  assign N998 = N997 | i[913];
  assign N997 = N996 | i[914];
  assign N996 = N995 | i[915];
  assign N995 = N994 | i[916];
  assign N994 = N993 | i[917];
  assign N993 = N992 | i[918];
  assign N992 = N991 | i[919];
  assign N991 = N990 | i[920];
  assign N990 = N989 | i[921];
  assign N989 = N988 | i[922];
  assign N988 = N987 | i[923];
  assign N987 = N986 | i[924];
  assign N986 = N985 | i[925];
  assign N985 = N984 | i[926];
  assign N984 = N983 | i[927];
  assign N983 = N982 | i[928];
  assign N982 = N981 | i[929];
  assign N981 = N980 | i[930];
  assign N980 = N979 | i[931];
  assign N979 = N978 | i[932];
  assign N978 = N977 | i[933];
  assign N977 = N976 | i[934];
  assign N976 = N975 | i[935];
  assign N975 = N974 | i[936];
  assign N974 = N973 | i[937];
  assign N973 = N972 | i[938];
  assign N972 = N971 | i[939];
  assign N971 = N970 | i[940];
  assign N970 = N969 | i[941];
  assign N969 = N968 | i[942];
  assign N968 = N967 | i[943];
  assign N967 = N966 | i[944];
  assign N966 = N965 | i[945];
  assign N965 = N964 | i[946];
  assign N964 = N963 | i[947];
  assign N963 = N962 | i[948];
  assign N962 = N961 | i[949];
  assign N961 = N960 | i[950];
  assign N960 = N959 | i[951];
  assign N959 = N958 | i[952];
  assign N958 = N957 | i[953];
  assign N957 = N956 | i[954];
  assign N956 = N955 | i[955];
  assign N955 = N954 | i[956];
  assign N954 = N953 | i[957];
  assign N953 = N952 | i[958];
  assign N952 = N951 | i[959];
  assign N951 = N950 | i[960];
  assign N950 = N949 | i[961];
  assign N949 = N948 | i[962];
  assign N948 = N947 | i[963];
  assign N947 = N946 | i[964];
  assign N946 = N945 | i[965];
  assign N945 = N944 | i[966];
  assign N944 = N943 | i[967];
  assign N943 = N942 | i[968];
  assign N942 = N941 | i[969];
  assign N941 = N940 | i[970];
  assign N940 = N939 | i[971];
  assign N939 = N938 | i[972];
  assign N938 = N937 | i[973];
  assign N937 = N936 | i[974];
  assign N936 = N935 | i[975];
  assign N935 = N934 | i[976];
  assign N934 = N933 | i[977];
  assign N933 = N932 | i[978];
  assign N932 = N931 | i[979];
  assign N931 = N930 | i[980];
  assign N930 = N929 | i[981];
  assign N929 = N928 | i[982];
  assign N928 = N927 | i[983];
  assign N927 = N926 | i[984];
  assign N926 = N925 | i[985];
  assign N925 = N924 | i[986];
  assign N924 = N923 | i[987];
  assign N923 = N922 | i[988];
  assign N922 = N921 | i[989];
  assign N921 = N920 | i[990];
  assign N920 = N919 | i[991];
  assign N919 = N918 | i[992];
  assign N918 = N917 | i[993];
  assign N917 = N916 | i[994];
  assign N916 = N915 | i[995];
  assign N915 = N914 | i[996];
  assign N914 = N913 | i[997];
  assign N913 = N912 | i[998];
  assign N912 = N911 | i[999];
  assign N911 = N910 | i[1000];
  assign N910 = N909 | i[1001];
  assign N909 = N908 | i[1002];
  assign N908 = N907 | i[1003];
  assign N907 = N906 | i[1004];
  assign N906 = N905 | i[1005];
  assign N905 = N904 | i[1006];
  assign N904 = N903 | i[1007];
  assign N903 = N902 | i[1008];
  assign N902 = N901 | i[1009];
  assign N901 = N900 | i[1010];
  assign N900 = N899 | i[1011];
  assign N899 = N898 | i[1012];
  assign N898 = N897 | i[1013];
  assign N897 = N896 | i[1014];
  assign N896 = N895 | i[1015];
  assign N895 = N894 | i[1016];
  assign N894 = N893 | i[1017];
  assign N893 = N892 | i[1018];
  assign N892 = N891 | i[1019];
  assign N891 = N890 | i[1020];
  assign N890 = N889 | i[1021];
  assign N889 = i[1023] | i[1022];
  assign o[8] = ~N1142;
  assign N1142 = N1141 | i[1024];
  assign N1141 = N1140 | i[1025];
  assign N1140 = N1139 | i[1026];
  assign N1139 = N1138 | i[1027];
  assign N1138 = N1137 | i[1028];
  assign N1137 = N1136 | i[1029];
  assign N1136 = N1135 | i[1030];
  assign N1135 = N1134 | i[1031];
  assign N1134 = N1133 | i[1032];
  assign N1133 = N1132 | i[1033];
  assign N1132 = N1131 | i[1034];
  assign N1131 = N1130 | i[1035];
  assign N1130 = N1129 | i[1036];
  assign N1129 = N1128 | i[1037];
  assign N1128 = N1127 | i[1038];
  assign N1127 = N1126 | i[1039];
  assign N1126 = N1125 | i[1040];
  assign N1125 = N1124 | i[1041];
  assign N1124 = N1123 | i[1042];
  assign N1123 = N1122 | i[1043];
  assign N1122 = N1121 | i[1044];
  assign N1121 = N1120 | i[1045];
  assign N1120 = N1119 | i[1046];
  assign N1119 = N1118 | i[1047];
  assign N1118 = N1117 | i[1048];
  assign N1117 = N1116 | i[1049];
  assign N1116 = N1115 | i[1050];
  assign N1115 = N1114 | i[1051];
  assign N1114 = N1113 | i[1052];
  assign N1113 = N1112 | i[1053];
  assign N1112 = N1111 | i[1054];
  assign N1111 = N1110 | i[1055];
  assign N1110 = N1109 | i[1056];
  assign N1109 = N1108 | i[1057];
  assign N1108 = N1107 | i[1058];
  assign N1107 = N1106 | i[1059];
  assign N1106 = N1105 | i[1060];
  assign N1105 = N1104 | i[1061];
  assign N1104 = N1103 | i[1062];
  assign N1103 = N1102 | i[1063];
  assign N1102 = N1101 | i[1064];
  assign N1101 = N1100 | i[1065];
  assign N1100 = N1099 | i[1066];
  assign N1099 = N1098 | i[1067];
  assign N1098 = N1097 | i[1068];
  assign N1097 = N1096 | i[1069];
  assign N1096 = N1095 | i[1070];
  assign N1095 = N1094 | i[1071];
  assign N1094 = N1093 | i[1072];
  assign N1093 = N1092 | i[1073];
  assign N1092 = N1091 | i[1074];
  assign N1091 = N1090 | i[1075];
  assign N1090 = N1089 | i[1076];
  assign N1089 = N1088 | i[1077];
  assign N1088 = N1087 | i[1078];
  assign N1087 = N1086 | i[1079];
  assign N1086 = N1085 | i[1080];
  assign N1085 = N1084 | i[1081];
  assign N1084 = N1083 | i[1082];
  assign N1083 = N1082 | i[1083];
  assign N1082 = N1081 | i[1084];
  assign N1081 = N1080 | i[1085];
  assign N1080 = N1079 | i[1086];
  assign N1079 = N1078 | i[1087];
  assign N1078 = N1077 | i[1088];
  assign N1077 = N1076 | i[1089];
  assign N1076 = N1075 | i[1090];
  assign N1075 = N1074 | i[1091];
  assign N1074 = N1073 | i[1092];
  assign N1073 = N1072 | i[1093];
  assign N1072 = N1071 | i[1094];
  assign N1071 = N1070 | i[1095];
  assign N1070 = N1069 | i[1096];
  assign N1069 = N1068 | i[1097];
  assign N1068 = N1067 | i[1098];
  assign N1067 = N1066 | i[1099];
  assign N1066 = N1065 | i[1100];
  assign N1065 = N1064 | i[1101];
  assign N1064 = N1063 | i[1102];
  assign N1063 = N1062 | i[1103];
  assign N1062 = N1061 | i[1104];
  assign N1061 = N1060 | i[1105];
  assign N1060 = N1059 | i[1106];
  assign N1059 = N1058 | i[1107];
  assign N1058 = N1057 | i[1108];
  assign N1057 = N1056 | i[1109];
  assign N1056 = N1055 | i[1110];
  assign N1055 = N1054 | i[1111];
  assign N1054 = N1053 | i[1112];
  assign N1053 = N1052 | i[1113];
  assign N1052 = N1051 | i[1114];
  assign N1051 = N1050 | i[1115];
  assign N1050 = N1049 | i[1116];
  assign N1049 = N1048 | i[1117];
  assign N1048 = N1047 | i[1118];
  assign N1047 = N1046 | i[1119];
  assign N1046 = N1045 | i[1120];
  assign N1045 = N1044 | i[1121];
  assign N1044 = N1043 | i[1122];
  assign N1043 = N1042 | i[1123];
  assign N1042 = N1041 | i[1124];
  assign N1041 = N1040 | i[1125];
  assign N1040 = N1039 | i[1126];
  assign N1039 = N1038 | i[1127];
  assign N1038 = N1037 | i[1128];
  assign N1037 = N1036 | i[1129];
  assign N1036 = N1035 | i[1130];
  assign N1035 = N1034 | i[1131];
  assign N1034 = N1033 | i[1132];
  assign N1033 = N1032 | i[1133];
  assign N1032 = N1031 | i[1134];
  assign N1031 = N1030 | i[1135];
  assign N1030 = N1029 | i[1136];
  assign N1029 = N1028 | i[1137];
  assign N1028 = N1027 | i[1138];
  assign N1027 = N1026 | i[1139];
  assign N1026 = N1025 | i[1140];
  assign N1025 = N1024 | i[1141];
  assign N1024 = N1023 | i[1142];
  assign N1023 = N1022 | i[1143];
  assign N1022 = N1021 | i[1144];
  assign N1021 = N1020 | i[1145];
  assign N1020 = N1019 | i[1146];
  assign N1019 = N1018 | i[1147];
  assign N1018 = N1017 | i[1148];
  assign N1017 = N1016 | i[1149];
  assign N1016 = i[1151] | i[1150];
  assign o[9] = ~N1269;
  assign N1269 = N1268 | i[1152];
  assign N1268 = N1267 | i[1153];
  assign N1267 = N1266 | i[1154];
  assign N1266 = N1265 | i[1155];
  assign N1265 = N1264 | i[1156];
  assign N1264 = N1263 | i[1157];
  assign N1263 = N1262 | i[1158];
  assign N1262 = N1261 | i[1159];
  assign N1261 = N1260 | i[1160];
  assign N1260 = N1259 | i[1161];
  assign N1259 = N1258 | i[1162];
  assign N1258 = N1257 | i[1163];
  assign N1257 = N1256 | i[1164];
  assign N1256 = N1255 | i[1165];
  assign N1255 = N1254 | i[1166];
  assign N1254 = N1253 | i[1167];
  assign N1253 = N1252 | i[1168];
  assign N1252 = N1251 | i[1169];
  assign N1251 = N1250 | i[1170];
  assign N1250 = N1249 | i[1171];
  assign N1249 = N1248 | i[1172];
  assign N1248 = N1247 | i[1173];
  assign N1247 = N1246 | i[1174];
  assign N1246 = N1245 | i[1175];
  assign N1245 = N1244 | i[1176];
  assign N1244 = N1243 | i[1177];
  assign N1243 = N1242 | i[1178];
  assign N1242 = N1241 | i[1179];
  assign N1241 = N1240 | i[1180];
  assign N1240 = N1239 | i[1181];
  assign N1239 = N1238 | i[1182];
  assign N1238 = N1237 | i[1183];
  assign N1237 = N1236 | i[1184];
  assign N1236 = N1235 | i[1185];
  assign N1235 = N1234 | i[1186];
  assign N1234 = N1233 | i[1187];
  assign N1233 = N1232 | i[1188];
  assign N1232 = N1231 | i[1189];
  assign N1231 = N1230 | i[1190];
  assign N1230 = N1229 | i[1191];
  assign N1229 = N1228 | i[1192];
  assign N1228 = N1227 | i[1193];
  assign N1227 = N1226 | i[1194];
  assign N1226 = N1225 | i[1195];
  assign N1225 = N1224 | i[1196];
  assign N1224 = N1223 | i[1197];
  assign N1223 = N1222 | i[1198];
  assign N1222 = N1221 | i[1199];
  assign N1221 = N1220 | i[1200];
  assign N1220 = N1219 | i[1201];
  assign N1219 = N1218 | i[1202];
  assign N1218 = N1217 | i[1203];
  assign N1217 = N1216 | i[1204];
  assign N1216 = N1215 | i[1205];
  assign N1215 = N1214 | i[1206];
  assign N1214 = N1213 | i[1207];
  assign N1213 = N1212 | i[1208];
  assign N1212 = N1211 | i[1209];
  assign N1211 = N1210 | i[1210];
  assign N1210 = N1209 | i[1211];
  assign N1209 = N1208 | i[1212];
  assign N1208 = N1207 | i[1213];
  assign N1207 = N1206 | i[1214];
  assign N1206 = N1205 | i[1215];
  assign N1205 = N1204 | i[1216];
  assign N1204 = N1203 | i[1217];
  assign N1203 = N1202 | i[1218];
  assign N1202 = N1201 | i[1219];
  assign N1201 = N1200 | i[1220];
  assign N1200 = N1199 | i[1221];
  assign N1199 = N1198 | i[1222];
  assign N1198 = N1197 | i[1223];
  assign N1197 = N1196 | i[1224];
  assign N1196 = N1195 | i[1225];
  assign N1195 = N1194 | i[1226];
  assign N1194 = N1193 | i[1227];
  assign N1193 = N1192 | i[1228];
  assign N1192 = N1191 | i[1229];
  assign N1191 = N1190 | i[1230];
  assign N1190 = N1189 | i[1231];
  assign N1189 = N1188 | i[1232];
  assign N1188 = N1187 | i[1233];
  assign N1187 = N1186 | i[1234];
  assign N1186 = N1185 | i[1235];
  assign N1185 = N1184 | i[1236];
  assign N1184 = N1183 | i[1237];
  assign N1183 = N1182 | i[1238];
  assign N1182 = N1181 | i[1239];
  assign N1181 = N1180 | i[1240];
  assign N1180 = N1179 | i[1241];
  assign N1179 = N1178 | i[1242];
  assign N1178 = N1177 | i[1243];
  assign N1177 = N1176 | i[1244];
  assign N1176 = N1175 | i[1245];
  assign N1175 = N1174 | i[1246];
  assign N1174 = N1173 | i[1247];
  assign N1173 = N1172 | i[1248];
  assign N1172 = N1171 | i[1249];
  assign N1171 = N1170 | i[1250];
  assign N1170 = N1169 | i[1251];
  assign N1169 = N1168 | i[1252];
  assign N1168 = N1167 | i[1253];
  assign N1167 = N1166 | i[1254];
  assign N1166 = N1165 | i[1255];
  assign N1165 = N1164 | i[1256];
  assign N1164 = N1163 | i[1257];
  assign N1163 = N1162 | i[1258];
  assign N1162 = N1161 | i[1259];
  assign N1161 = N1160 | i[1260];
  assign N1160 = N1159 | i[1261];
  assign N1159 = N1158 | i[1262];
  assign N1158 = N1157 | i[1263];
  assign N1157 = N1156 | i[1264];
  assign N1156 = N1155 | i[1265];
  assign N1155 = N1154 | i[1266];
  assign N1154 = N1153 | i[1267];
  assign N1153 = N1152 | i[1268];
  assign N1152 = N1151 | i[1269];
  assign N1151 = N1150 | i[1270];
  assign N1150 = N1149 | i[1271];
  assign N1149 = N1148 | i[1272];
  assign N1148 = N1147 | i[1273];
  assign N1147 = N1146 | i[1274];
  assign N1146 = N1145 | i[1275];
  assign N1145 = N1144 | i[1276];
  assign N1144 = N1143 | i[1277];
  assign N1143 = i[1279] | i[1278];
  assign o[10] = ~N1396;
  assign N1396 = N1395 | i[1280];
  assign N1395 = N1394 | i[1281];
  assign N1394 = N1393 | i[1282];
  assign N1393 = N1392 | i[1283];
  assign N1392 = N1391 | i[1284];
  assign N1391 = N1390 | i[1285];
  assign N1390 = N1389 | i[1286];
  assign N1389 = N1388 | i[1287];
  assign N1388 = N1387 | i[1288];
  assign N1387 = N1386 | i[1289];
  assign N1386 = N1385 | i[1290];
  assign N1385 = N1384 | i[1291];
  assign N1384 = N1383 | i[1292];
  assign N1383 = N1382 | i[1293];
  assign N1382 = N1381 | i[1294];
  assign N1381 = N1380 | i[1295];
  assign N1380 = N1379 | i[1296];
  assign N1379 = N1378 | i[1297];
  assign N1378 = N1377 | i[1298];
  assign N1377 = N1376 | i[1299];
  assign N1376 = N1375 | i[1300];
  assign N1375 = N1374 | i[1301];
  assign N1374 = N1373 | i[1302];
  assign N1373 = N1372 | i[1303];
  assign N1372 = N1371 | i[1304];
  assign N1371 = N1370 | i[1305];
  assign N1370 = N1369 | i[1306];
  assign N1369 = N1368 | i[1307];
  assign N1368 = N1367 | i[1308];
  assign N1367 = N1366 | i[1309];
  assign N1366 = N1365 | i[1310];
  assign N1365 = N1364 | i[1311];
  assign N1364 = N1363 | i[1312];
  assign N1363 = N1362 | i[1313];
  assign N1362 = N1361 | i[1314];
  assign N1361 = N1360 | i[1315];
  assign N1360 = N1359 | i[1316];
  assign N1359 = N1358 | i[1317];
  assign N1358 = N1357 | i[1318];
  assign N1357 = N1356 | i[1319];
  assign N1356 = N1355 | i[1320];
  assign N1355 = N1354 | i[1321];
  assign N1354 = N1353 | i[1322];
  assign N1353 = N1352 | i[1323];
  assign N1352 = N1351 | i[1324];
  assign N1351 = N1350 | i[1325];
  assign N1350 = N1349 | i[1326];
  assign N1349 = N1348 | i[1327];
  assign N1348 = N1347 | i[1328];
  assign N1347 = N1346 | i[1329];
  assign N1346 = N1345 | i[1330];
  assign N1345 = N1344 | i[1331];
  assign N1344 = N1343 | i[1332];
  assign N1343 = N1342 | i[1333];
  assign N1342 = N1341 | i[1334];
  assign N1341 = N1340 | i[1335];
  assign N1340 = N1339 | i[1336];
  assign N1339 = N1338 | i[1337];
  assign N1338 = N1337 | i[1338];
  assign N1337 = N1336 | i[1339];
  assign N1336 = N1335 | i[1340];
  assign N1335 = N1334 | i[1341];
  assign N1334 = N1333 | i[1342];
  assign N1333 = N1332 | i[1343];
  assign N1332 = N1331 | i[1344];
  assign N1331 = N1330 | i[1345];
  assign N1330 = N1329 | i[1346];
  assign N1329 = N1328 | i[1347];
  assign N1328 = N1327 | i[1348];
  assign N1327 = N1326 | i[1349];
  assign N1326 = N1325 | i[1350];
  assign N1325 = N1324 | i[1351];
  assign N1324 = N1323 | i[1352];
  assign N1323 = N1322 | i[1353];
  assign N1322 = N1321 | i[1354];
  assign N1321 = N1320 | i[1355];
  assign N1320 = N1319 | i[1356];
  assign N1319 = N1318 | i[1357];
  assign N1318 = N1317 | i[1358];
  assign N1317 = N1316 | i[1359];
  assign N1316 = N1315 | i[1360];
  assign N1315 = N1314 | i[1361];
  assign N1314 = N1313 | i[1362];
  assign N1313 = N1312 | i[1363];
  assign N1312 = N1311 | i[1364];
  assign N1311 = N1310 | i[1365];
  assign N1310 = N1309 | i[1366];
  assign N1309 = N1308 | i[1367];
  assign N1308 = N1307 | i[1368];
  assign N1307 = N1306 | i[1369];
  assign N1306 = N1305 | i[1370];
  assign N1305 = N1304 | i[1371];
  assign N1304 = N1303 | i[1372];
  assign N1303 = N1302 | i[1373];
  assign N1302 = N1301 | i[1374];
  assign N1301 = N1300 | i[1375];
  assign N1300 = N1299 | i[1376];
  assign N1299 = N1298 | i[1377];
  assign N1298 = N1297 | i[1378];
  assign N1297 = N1296 | i[1379];
  assign N1296 = N1295 | i[1380];
  assign N1295 = N1294 | i[1381];
  assign N1294 = N1293 | i[1382];
  assign N1293 = N1292 | i[1383];
  assign N1292 = N1291 | i[1384];
  assign N1291 = N1290 | i[1385];
  assign N1290 = N1289 | i[1386];
  assign N1289 = N1288 | i[1387];
  assign N1288 = N1287 | i[1388];
  assign N1287 = N1286 | i[1389];
  assign N1286 = N1285 | i[1390];
  assign N1285 = N1284 | i[1391];
  assign N1284 = N1283 | i[1392];
  assign N1283 = N1282 | i[1393];
  assign N1282 = N1281 | i[1394];
  assign N1281 = N1280 | i[1395];
  assign N1280 = N1279 | i[1396];
  assign N1279 = N1278 | i[1397];
  assign N1278 = N1277 | i[1398];
  assign N1277 = N1276 | i[1399];
  assign N1276 = N1275 | i[1400];
  assign N1275 = N1274 | i[1401];
  assign N1274 = N1273 | i[1402];
  assign N1273 = N1272 | i[1403];
  assign N1272 = N1271 | i[1404];
  assign N1271 = N1270 | i[1405];
  assign N1270 = i[1407] | i[1406];
  assign o[11] = ~N1523;
  assign N1523 = N1522 | i[1408];
  assign N1522 = N1521 | i[1409];
  assign N1521 = N1520 | i[1410];
  assign N1520 = N1519 | i[1411];
  assign N1519 = N1518 | i[1412];
  assign N1518 = N1517 | i[1413];
  assign N1517 = N1516 | i[1414];
  assign N1516 = N1515 | i[1415];
  assign N1515 = N1514 | i[1416];
  assign N1514 = N1513 | i[1417];
  assign N1513 = N1512 | i[1418];
  assign N1512 = N1511 | i[1419];
  assign N1511 = N1510 | i[1420];
  assign N1510 = N1509 | i[1421];
  assign N1509 = N1508 | i[1422];
  assign N1508 = N1507 | i[1423];
  assign N1507 = N1506 | i[1424];
  assign N1506 = N1505 | i[1425];
  assign N1505 = N1504 | i[1426];
  assign N1504 = N1503 | i[1427];
  assign N1503 = N1502 | i[1428];
  assign N1502 = N1501 | i[1429];
  assign N1501 = N1500 | i[1430];
  assign N1500 = N1499 | i[1431];
  assign N1499 = N1498 | i[1432];
  assign N1498 = N1497 | i[1433];
  assign N1497 = N1496 | i[1434];
  assign N1496 = N1495 | i[1435];
  assign N1495 = N1494 | i[1436];
  assign N1494 = N1493 | i[1437];
  assign N1493 = N1492 | i[1438];
  assign N1492 = N1491 | i[1439];
  assign N1491 = N1490 | i[1440];
  assign N1490 = N1489 | i[1441];
  assign N1489 = N1488 | i[1442];
  assign N1488 = N1487 | i[1443];
  assign N1487 = N1486 | i[1444];
  assign N1486 = N1485 | i[1445];
  assign N1485 = N1484 | i[1446];
  assign N1484 = N1483 | i[1447];
  assign N1483 = N1482 | i[1448];
  assign N1482 = N1481 | i[1449];
  assign N1481 = N1480 | i[1450];
  assign N1480 = N1479 | i[1451];
  assign N1479 = N1478 | i[1452];
  assign N1478 = N1477 | i[1453];
  assign N1477 = N1476 | i[1454];
  assign N1476 = N1475 | i[1455];
  assign N1475 = N1474 | i[1456];
  assign N1474 = N1473 | i[1457];
  assign N1473 = N1472 | i[1458];
  assign N1472 = N1471 | i[1459];
  assign N1471 = N1470 | i[1460];
  assign N1470 = N1469 | i[1461];
  assign N1469 = N1468 | i[1462];
  assign N1468 = N1467 | i[1463];
  assign N1467 = N1466 | i[1464];
  assign N1466 = N1465 | i[1465];
  assign N1465 = N1464 | i[1466];
  assign N1464 = N1463 | i[1467];
  assign N1463 = N1462 | i[1468];
  assign N1462 = N1461 | i[1469];
  assign N1461 = N1460 | i[1470];
  assign N1460 = N1459 | i[1471];
  assign N1459 = N1458 | i[1472];
  assign N1458 = N1457 | i[1473];
  assign N1457 = N1456 | i[1474];
  assign N1456 = N1455 | i[1475];
  assign N1455 = N1454 | i[1476];
  assign N1454 = N1453 | i[1477];
  assign N1453 = N1452 | i[1478];
  assign N1452 = N1451 | i[1479];
  assign N1451 = N1450 | i[1480];
  assign N1450 = N1449 | i[1481];
  assign N1449 = N1448 | i[1482];
  assign N1448 = N1447 | i[1483];
  assign N1447 = N1446 | i[1484];
  assign N1446 = N1445 | i[1485];
  assign N1445 = N1444 | i[1486];
  assign N1444 = N1443 | i[1487];
  assign N1443 = N1442 | i[1488];
  assign N1442 = N1441 | i[1489];
  assign N1441 = N1440 | i[1490];
  assign N1440 = N1439 | i[1491];
  assign N1439 = N1438 | i[1492];
  assign N1438 = N1437 | i[1493];
  assign N1437 = N1436 | i[1494];
  assign N1436 = N1435 | i[1495];
  assign N1435 = N1434 | i[1496];
  assign N1434 = N1433 | i[1497];
  assign N1433 = N1432 | i[1498];
  assign N1432 = N1431 | i[1499];
  assign N1431 = N1430 | i[1500];
  assign N1430 = N1429 | i[1501];
  assign N1429 = N1428 | i[1502];
  assign N1428 = N1427 | i[1503];
  assign N1427 = N1426 | i[1504];
  assign N1426 = N1425 | i[1505];
  assign N1425 = N1424 | i[1506];
  assign N1424 = N1423 | i[1507];
  assign N1423 = N1422 | i[1508];
  assign N1422 = N1421 | i[1509];
  assign N1421 = N1420 | i[1510];
  assign N1420 = N1419 | i[1511];
  assign N1419 = N1418 | i[1512];
  assign N1418 = N1417 | i[1513];
  assign N1417 = N1416 | i[1514];
  assign N1416 = N1415 | i[1515];
  assign N1415 = N1414 | i[1516];
  assign N1414 = N1413 | i[1517];
  assign N1413 = N1412 | i[1518];
  assign N1412 = N1411 | i[1519];
  assign N1411 = N1410 | i[1520];
  assign N1410 = N1409 | i[1521];
  assign N1409 = N1408 | i[1522];
  assign N1408 = N1407 | i[1523];
  assign N1407 = N1406 | i[1524];
  assign N1406 = N1405 | i[1525];
  assign N1405 = N1404 | i[1526];
  assign N1404 = N1403 | i[1527];
  assign N1403 = N1402 | i[1528];
  assign N1402 = N1401 | i[1529];
  assign N1401 = N1400 | i[1530];
  assign N1400 = N1399 | i[1531];
  assign N1399 = N1398 | i[1532];
  assign N1398 = N1397 | i[1533];
  assign N1397 = i[1535] | i[1534];
  assign o[12] = ~N1650;
  assign N1650 = N1649 | i[1536];
  assign N1649 = N1648 | i[1537];
  assign N1648 = N1647 | i[1538];
  assign N1647 = N1646 | i[1539];
  assign N1646 = N1645 | i[1540];
  assign N1645 = N1644 | i[1541];
  assign N1644 = N1643 | i[1542];
  assign N1643 = N1642 | i[1543];
  assign N1642 = N1641 | i[1544];
  assign N1641 = N1640 | i[1545];
  assign N1640 = N1639 | i[1546];
  assign N1639 = N1638 | i[1547];
  assign N1638 = N1637 | i[1548];
  assign N1637 = N1636 | i[1549];
  assign N1636 = N1635 | i[1550];
  assign N1635 = N1634 | i[1551];
  assign N1634 = N1633 | i[1552];
  assign N1633 = N1632 | i[1553];
  assign N1632 = N1631 | i[1554];
  assign N1631 = N1630 | i[1555];
  assign N1630 = N1629 | i[1556];
  assign N1629 = N1628 | i[1557];
  assign N1628 = N1627 | i[1558];
  assign N1627 = N1626 | i[1559];
  assign N1626 = N1625 | i[1560];
  assign N1625 = N1624 | i[1561];
  assign N1624 = N1623 | i[1562];
  assign N1623 = N1622 | i[1563];
  assign N1622 = N1621 | i[1564];
  assign N1621 = N1620 | i[1565];
  assign N1620 = N1619 | i[1566];
  assign N1619 = N1618 | i[1567];
  assign N1618 = N1617 | i[1568];
  assign N1617 = N1616 | i[1569];
  assign N1616 = N1615 | i[1570];
  assign N1615 = N1614 | i[1571];
  assign N1614 = N1613 | i[1572];
  assign N1613 = N1612 | i[1573];
  assign N1612 = N1611 | i[1574];
  assign N1611 = N1610 | i[1575];
  assign N1610 = N1609 | i[1576];
  assign N1609 = N1608 | i[1577];
  assign N1608 = N1607 | i[1578];
  assign N1607 = N1606 | i[1579];
  assign N1606 = N1605 | i[1580];
  assign N1605 = N1604 | i[1581];
  assign N1604 = N1603 | i[1582];
  assign N1603 = N1602 | i[1583];
  assign N1602 = N1601 | i[1584];
  assign N1601 = N1600 | i[1585];
  assign N1600 = N1599 | i[1586];
  assign N1599 = N1598 | i[1587];
  assign N1598 = N1597 | i[1588];
  assign N1597 = N1596 | i[1589];
  assign N1596 = N1595 | i[1590];
  assign N1595 = N1594 | i[1591];
  assign N1594 = N1593 | i[1592];
  assign N1593 = N1592 | i[1593];
  assign N1592 = N1591 | i[1594];
  assign N1591 = N1590 | i[1595];
  assign N1590 = N1589 | i[1596];
  assign N1589 = N1588 | i[1597];
  assign N1588 = N1587 | i[1598];
  assign N1587 = N1586 | i[1599];
  assign N1586 = N1585 | i[1600];
  assign N1585 = N1584 | i[1601];
  assign N1584 = N1583 | i[1602];
  assign N1583 = N1582 | i[1603];
  assign N1582 = N1581 | i[1604];
  assign N1581 = N1580 | i[1605];
  assign N1580 = N1579 | i[1606];
  assign N1579 = N1578 | i[1607];
  assign N1578 = N1577 | i[1608];
  assign N1577 = N1576 | i[1609];
  assign N1576 = N1575 | i[1610];
  assign N1575 = N1574 | i[1611];
  assign N1574 = N1573 | i[1612];
  assign N1573 = N1572 | i[1613];
  assign N1572 = N1571 | i[1614];
  assign N1571 = N1570 | i[1615];
  assign N1570 = N1569 | i[1616];
  assign N1569 = N1568 | i[1617];
  assign N1568 = N1567 | i[1618];
  assign N1567 = N1566 | i[1619];
  assign N1566 = N1565 | i[1620];
  assign N1565 = N1564 | i[1621];
  assign N1564 = N1563 | i[1622];
  assign N1563 = N1562 | i[1623];
  assign N1562 = N1561 | i[1624];
  assign N1561 = N1560 | i[1625];
  assign N1560 = N1559 | i[1626];
  assign N1559 = N1558 | i[1627];
  assign N1558 = N1557 | i[1628];
  assign N1557 = N1556 | i[1629];
  assign N1556 = N1555 | i[1630];
  assign N1555 = N1554 | i[1631];
  assign N1554 = N1553 | i[1632];
  assign N1553 = N1552 | i[1633];
  assign N1552 = N1551 | i[1634];
  assign N1551 = N1550 | i[1635];
  assign N1550 = N1549 | i[1636];
  assign N1549 = N1548 | i[1637];
  assign N1548 = N1547 | i[1638];
  assign N1547 = N1546 | i[1639];
  assign N1546 = N1545 | i[1640];
  assign N1545 = N1544 | i[1641];
  assign N1544 = N1543 | i[1642];
  assign N1543 = N1542 | i[1643];
  assign N1542 = N1541 | i[1644];
  assign N1541 = N1540 | i[1645];
  assign N1540 = N1539 | i[1646];
  assign N1539 = N1538 | i[1647];
  assign N1538 = N1537 | i[1648];
  assign N1537 = N1536 | i[1649];
  assign N1536 = N1535 | i[1650];
  assign N1535 = N1534 | i[1651];
  assign N1534 = N1533 | i[1652];
  assign N1533 = N1532 | i[1653];
  assign N1532 = N1531 | i[1654];
  assign N1531 = N1530 | i[1655];
  assign N1530 = N1529 | i[1656];
  assign N1529 = N1528 | i[1657];
  assign N1528 = N1527 | i[1658];
  assign N1527 = N1526 | i[1659];
  assign N1526 = N1525 | i[1660];
  assign N1525 = N1524 | i[1661];
  assign N1524 = i[1663] | i[1662];
  assign o[13] = ~N1777;
  assign N1777 = N1776 | i[1664];
  assign N1776 = N1775 | i[1665];
  assign N1775 = N1774 | i[1666];
  assign N1774 = N1773 | i[1667];
  assign N1773 = N1772 | i[1668];
  assign N1772 = N1771 | i[1669];
  assign N1771 = N1770 | i[1670];
  assign N1770 = N1769 | i[1671];
  assign N1769 = N1768 | i[1672];
  assign N1768 = N1767 | i[1673];
  assign N1767 = N1766 | i[1674];
  assign N1766 = N1765 | i[1675];
  assign N1765 = N1764 | i[1676];
  assign N1764 = N1763 | i[1677];
  assign N1763 = N1762 | i[1678];
  assign N1762 = N1761 | i[1679];
  assign N1761 = N1760 | i[1680];
  assign N1760 = N1759 | i[1681];
  assign N1759 = N1758 | i[1682];
  assign N1758 = N1757 | i[1683];
  assign N1757 = N1756 | i[1684];
  assign N1756 = N1755 | i[1685];
  assign N1755 = N1754 | i[1686];
  assign N1754 = N1753 | i[1687];
  assign N1753 = N1752 | i[1688];
  assign N1752 = N1751 | i[1689];
  assign N1751 = N1750 | i[1690];
  assign N1750 = N1749 | i[1691];
  assign N1749 = N1748 | i[1692];
  assign N1748 = N1747 | i[1693];
  assign N1747 = N1746 | i[1694];
  assign N1746 = N1745 | i[1695];
  assign N1745 = N1744 | i[1696];
  assign N1744 = N1743 | i[1697];
  assign N1743 = N1742 | i[1698];
  assign N1742 = N1741 | i[1699];
  assign N1741 = N1740 | i[1700];
  assign N1740 = N1739 | i[1701];
  assign N1739 = N1738 | i[1702];
  assign N1738 = N1737 | i[1703];
  assign N1737 = N1736 | i[1704];
  assign N1736 = N1735 | i[1705];
  assign N1735 = N1734 | i[1706];
  assign N1734 = N1733 | i[1707];
  assign N1733 = N1732 | i[1708];
  assign N1732 = N1731 | i[1709];
  assign N1731 = N1730 | i[1710];
  assign N1730 = N1729 | i[1711];
  assign N1729 = N1728 | i[1712];
  assign N1728 = N1727 | i[1713];
  assign N1727 = N1726 | i[1714];
  assign N1726 = N1725 | i[1715];
  assign N1725 = N1724 | i[1716];
  assign N1724 = N1723 | i[1717];
  assign N1723 = N1722 | i[1718];
  assign N1722 = N1721 | i[1719];
  assign N1721 = N1720 | i[1720];
  assign N1720 = N1719 | i[1721];
  assign N1719 = N1718 | i[1722];
  assign N1718 = N1717 | i[1723];
  assign N1717 = N1716 | i[1724];
  assign N1716 = N1715 | i[1725];
  assign N1715 = N1714 | i[1726];
  assign N1714 = N1713 | i[1727];
  assign N1713 = N1712 | i[1728];
  assign N1712 = N1711 | i[1729];
  assign N1711 = N1710 | i[1730];
  assign N1710 = N1709 | i[1731];
  assign N1709 = N1708 | i[1732];
  assign N1708 = N1707 | i[1733];
  assign N1707 = N1706 | i[1734];
  assign N1706 = N1705 | i[1735];
  assign N1705 = N1704 | i[1736];
  assign N1704 = N1703 | i[1737];
  assign N1703 = N1702 | i[1738];
  assign N1702 = N1701 | i[1739];
  assign N1701 = N1700 | i[1740];
  assign N1700 = N1699 | i[1741];
  assign N1699 = N1698 | i[1742];
  assign N1698 = N1697 | i[1743];
  assign N1697 = N1696 | i[1744];
  assign N1696 = N1695 | i[1745];
  assign N1695 = N1694 | i[1746];
  assign N1694 = N1693 | i[1747];
  assign N1693 = N1692 | i[1748];
  assign N1692 = N1691 | i[1749];
  assign N1691 = N1690 | i[1750];
  assign N1690 = N1689 | i[1751];
  assign N1689 = N1688 | i[1752];
  assign N1688 = N1687 | i[1753];
  assign N1687 = N1686 | i[1754];
  assign N1686 = N1685 | i[1755];
  assign N1685 = N1684 | i[1756];
  assign N1684 = N1683 | i[1757];
  assign N1683 = N1682 | i[1758];
  assign N1682 = N1681 | i[1759];
  assign N1681 = N1680 | i[1760];
  assign N1680 = N1679 | i[1761];
  assign N1679 = N1678 | i[1762];
  assign N1678 = N1677 | i[1763];
  assign N1677 = N1676 | i[1764];
  assign N1676 = N1675 | i[1765];
  assign N1675 = N1674 | i[1766];
  assign N1674 = N1673 | i[1767];
  assign N1673 = N1672 | i[1768];
  assign N1672 = N1671 | i[1769];
  assign N1671 = N1670 | i[1770];
  assign N1670 = N1669 | i[1771];
  assign N1669 = N1668 | i[1772];
  assign N1668 = N1667 | i[1773];
  assign N1667 = N1666 | i[1774];
  assign N1666 = N1665 | i[1775];
  assign N1665 = N1664 | i[1776];
  assign N1664 = N1663 | i[1777];
  assign N1663 = N1662 | i[1778];
  assign N1662 = N1661 | i[1779];
  assign N1661 = N1660 | i[1780];
  assign N1660 = N1659 | i[1781];
  assign N1659 = N1658 | i[1782];
  assign N1658 = N1657 | i[1783];
  assign N1657 = N1656 | i[1784];
  assign N1656 = N1655 | i[1785];
  assign N1655 = N1654 | i[1786];
  assign N1654 = N1653 | i[1787];
  assign N1653 = N1652 | i[1788];
  assign N1652 = N1651 | i[1789];
  assign N1651 = i[1791] | i[1790];
  assign o[14] = ~N1904;
  assign N1904 = N1903 | i[1792];
  assign N1903 = N1902 | i[1793];
  assign N1902 = N1901 | i[1794];
  assign N1901 = N1900 | i[1795];
  assign N1900 = N1899 | i[1796];
  assign N1899 = N1898 | i[1797];
  assign N1898 = N1897 | i[1798];
  assign N1897 = N1896 | i[1799];
  assign N1896 = N1895 | i[1800];
  assign N1895 = N1894 | i[1801];
  assign N1894 = N1893 | i[1802];
  assign N1893 = N1892 | i[1803];
  assign N1892 = N1891 | i[1804];
  assign N1891 = N1890 | i[1805];
  assign N1890 = N1889 | i[1806];
  assign N1889 = N1888 | i[1807];
  assign N1888 = N1887 | i[1808];
  assign N1887 = N1886 | i[1809];
  assign N1886 = N1885 | i[1810];
  assign N1885 = N1884 | i[1811];
  assign N1884 = N1883 | i[1812];
  assign N1883 = N1882 | i[1813];
  assign N1882 = N1881 | i[1814];
  assign N1881 = N1880 | i[1815];
  assign N1880 = N1879 | i[1816];
  assign N1879 = N1878 | i[1817];
  assign N1878 = N1877 | i[1818];
  assign N1877 = N1876 | i[1819];
  assign N1876 = N1875 | i[1820];
  assign N1875 = N1874 | i[1821];
  assign N1874 = N1873 | i[1822];
  assign N1873 = N1872 | i[1823];
  assign N1872 = N1871 | i[1824];
  assign N1871 = N1870 | i[1825];
  assign N1870 = N1869 | i[1826];
  assign N1869 = N1868 | i[1827];
  assign N1868 = N1867 | i[1828];
  assign N1867 = N1866 | i[1829];
  assign N1866 = N1865 | i[1830];
  assign N1865 = N1864 | i[1831];
  assign N1864 = N1863 | i[1832];
  assign N1863 = N1862 | i[1833];
  assign N1862 = N1861 | i[1834];
  assign N1861 = N1860 | i[1835];
  assign N1860 = N1859 | i[1836];
  assign N1859 = N1858 | i[1837];
  assign N1858 = N1857 | i[1838];
  assign N1857 = N1856 | i[1839];
  assign N1856 = N1855 | i[1840];
  assign N1855 = N1854 | i[1841];
  assign N1854 = N1853 | i[1842];
  assign N1853 = N1852 | i[1843];
  assign N1852 = N1851 | i[1844];
  assign N1851 = N1850 | i[1845];
  assign N1850 = N1849 | i[1846];
  assign N1849 = N1848 | i[1847];
  assign N1848 = N1847 | i[1848];
  assign N1847 = N1846 | i[1849];
  assign N1846 = N1845 | i[1850];
  assign N1845 = N1844 | i[1851];
  assign N1844 = N1843 | i[1852];
  assign N1843 = N1842 | i[1853];
  assign N1842 = N1841 | i[1854];
  assign N1841 = N1840 | i[1855];
  assign N1840 = N1839 | i[1856];
  assign N1839 = N1838 | i[1857];
  assign N1838 = N1837 | i[1858];
  assign N1837 = N1836 | i[1859];
  assign N1836 = N1835 | i[1860];
  assign N1835 = N1834 | i[1861];
  assign N1834 = N1833 | i[1862];
  assign N1833 = N1832 | i[1863];
  assign N1832 = N1831 | i[1864];
  assign N1831 = N1830 | i[1865];
  assign N1830 = N1829 | i[1866];
  assign N1829 = N1828 | i[1867];
  assign N1828 = N1827 | i[1868];
  assign N1827 = N1826 | i[1869];
  assign N1826 = N1825 | i[1870];
  assign N1825 = N1824 | i[1871];
  assign N1824 = N1823 | i[1872];
  assign N1823 = N1822 | i[1873];
  assign N1822 = N1821 | i[1874];
  assign N1821 = N1820 | i[1875];
  assign N1820 = N1819 | i[1876];
  assign N1819 = N1818 | i[1877];
  assign N1818 = N1817 | i[1878];
  assign N1817 = N1816 | i[1879];
  assign N1816 = N1815 | i[1880];
  assign N1815 = N1814 | i[1881];
  assign N1814 = N1813 | i[1882];
  assign N1813 = N1812 | i[1883];
  assign N1812 = N1811 | i[1884];
  assign N1811 = N1810 | i[1885];
  assign N1810 = N1809 | i[1886];
  assign N1809 = N1808 | i[1887];
  assign N1808 = N1807 | i[1888];
  assign N1807 = N1806 | i[1889];
  assign N1806 = N1805 | i[1890];
  assign N1805 = N1804 | i[1891];
  assign N1804 = N1803 | i[1892];
  assign N1803 = N1802 | i[1893];
  assign N1802 = N1801 | i[1894];
  assign N1801 = N1800 | i[1895];
  assign N1800 = N1799 | i[1896];
  assign N1799 = N1798 | i[1897];
  assign N1798 = N1797 | i[1898];
  assign N1797 = N1796 | i[1899];
  assign N1796 = N1795 | i[1900];
  assign N1795 = N1794 | i[1901];
  assign N1794 = N1793 | i[1902];
  assign N1793 = N1792 | i[1903];
  assign N1792 = N1791 | i[1904];
  assign N1791 = N1790 | i[1905];
  assign N1790 = N1789 | i[1906];
  assign N1789 = N1788 | i[1907];
  assign N1788 = N1787 | i[1908];
  assign N1787 = N1786 | i[1909];
  assign N1786 = N1785 | i[1910];
  assign N1785 = N1784 | i[1911];
  assign N1784 = N1783 | i[1912];
  assign N1783 = N1782 | i[1913];
  assign N1782 = N1781 | i[1914];
  assign N1781 = N1780 | i[1915];
  assign N1780 = N1779 | i[1916];
  assign N1779 = N1778 | i[1917];
  assign N1778 = i[1919] | i[1918];
  assign o[15] = ~N2031;
  assign N2031 = N2030 | i[1920];
  assign N2030 = N2029 | i[1921];
  assign N2029 = N2028 | i[1922];
  assign N2028 = N2027 | i[1923];
  assign N2027 = N2026 | i[1924];
  assign N2026 = N2025 | i[1925];
  assign N2025 = N2024 | i[1926];
  assign N2024 = N2023 | i[1927];
  assign N2023 = N2022 | i[1928];
  assign N2022 = N2021 | i[1929];
  assign N2021 = N2020 | i[1930];
  assign N2020 = N2019 | i[1931];
  assign N2019 = N2018 | i[1932];
  assign N2018 = N2017 | i[1933];
  assign N2017 = N2016 | i[1934];
  assign N2016 = N2015 | i[1935];
  assign N2015 = N2014 | i[1936];
  assign N2014 = N2013 | i[1937];
  assign N2013 = N2012 | i[1938];
  assign N2012 = N2011 | i[1939];
  assign N2011 = N2010 | i[1940];
  assign N2010 = N2009 | i[1941];
  assign N2009 = N2008 | i[1942];
  assign N2008 = N2007 | i[1943];
  assign N2007 = N2006 | i[1944];
  assign N2006 = N2005 | i[1945];
  assign N2005 = N2004 | i[1946];
  assign N2004 = N2003 | i[1947];
  assign N2003 = N2002 | i[1948];
  assign N2002 = N2001 | i[1949];
  assign N2001 = N2000 | i[1950];
  assign N2000 = N1999 | i[1951];
  assign N1999 = N1998 | i[1952];
  assign N1998 = N1997 | i[1953];
  assign N1997 = N1996 | i[1954];
  assign N1996 = N1995 | i[1955];
  assign N1995 = N1994 | i[1956];
  assign N1994 = N1993 | i[1957];
  assign N1993 = N1992 | i[1958];
  assign N1992 = N1991 | i[1959];
  assign N1991 = N1990 | i[1960];
  assign N1990 = N1989 | i[1961];
  assign N1989 = N1988 | i[1962];
  assign N1988 = N1987 | i[1963];
  assign N1987 = N1986 | i[1964];
  assign N1986 = N1985 | i[1965];
  assign N1985 = N1984 | i[1966];
  assign N1984 = N1983 | i[1967];
  assign N1983 = N1982 | i[1968];
  assign N1982 = N1981 | i[1969];
  assign N1981 = N1980 | i[1970];
  assign N1980 = N1979 | i[1971];
  assign N1979 = N1978 | i[1972];
  assign N1978 = N1977 | i[1973];
  assign N1977 = N1976 | i[1974];
  assign N1976 = N1975 | i[1975];
  assign N1975 = N1974 | i[1976];
  assign N1974 = N1973 | i[1977];
  assign N1973 = N1972 | i[1978];
  assign N1972 = N1971 | i[1979];
  assign N1971 = N1970 | i[1980];
  assign N1970 = N1969 | i[1981];
  assign N1969 = N1968 | i[1982];
  assign N1968 = N1967 | i[1983];
  assign N1967 = N1966 | i[1984];
  assign N1966 = N1965 | i[1985];
  assign N1965 = N1964 | i[1986];
  assign N1964 = N1963 | i[1987];
  assign N1963 = N1962 | i[1988];
  assign N1962 = N1961 | i[1989];
  assign N1961 = N1960 | i[1990];
  assign N1960 = N1959 | i[1991];
  assign N1959 = N1958 | i[1992];
  assign N1958 = N1957 | i[1993];
  assign N1957 = N1956 | i[1994];
  assign N1956 = N1955 | i[1995];
  assign N1955 = N1954 | i[1996];
  assign N1954 = N1953 | i[1997];
  assign N1953 = N1952 | i[1998];
  assign N1952 = N1951 | i[1999];
  assign N1951 = N1950 | i[2000];
  assign N1950 = N1949 | i[2001];
  assign N1949 = N1948 | i[2002];
  assign N1948 = N1947 | i[2003];
  assign N1947 = N1946 | i[2004];
  assign N1946 = N1945 | i[2005];
  assign N1945 = N1944 | i[2006];
  assign N1944 = N1943 | i[2007];
  assign N1943 = N1942 | i[2008];
  assign N1942 = N1941 | i[2009];
  assign N1941 = N1940 | i[2010];
  assign N1940 = N1939 | i[2011];
  assign N1939 = N1938 | i[2012];
  assign N1938 = N1937 | i[2013];
  assign N1937 = N1936 | i[2014];
  assign N1936 = N1935 | i[2015];
  assign N1935 = N1934 | i[2016];
  assign N1934 = N1933 | i[2017];
  assign N1933 = N1932 | i[2018];
  assign N1932 = N1931 | i[2019];
  assign N1931 = N1930 | i[2020];
  assign N1930 = N1929 | i[2021];
  assign N1929 = N1928 | i[2022];
  assign N1928 = N1927 | i[2023];
  assign N1927 = N1926 | i[2024];
  assign N1926 = N1925 | i[2025];
  assign N1925 = N1924 | i[2026];
  assign N1924 = N1923 | i[2027];
  assign N1923 = N1922 | i[2028];
  assign N1922 = N1921 | i[2029];
  assign N1921 = N1920 | i[2030];
  assign N1920 = N1919 | i[2031];
  assign N1919 = N1918 | i[2032];
  assign N1918 = N1917 | i[2033];
  assign N1917 = N1916 | i[2034];
  assign N1916 = N1915 | i[2035];
  assign N1915 = N1914 | i[2036];
  assign N1914 = N1913 | i[2037];
  assign N1913 = N1912 | i[2038];
  assign N1912 = N1911 | i[2039];
  assign N1911 = N1910 | i[2040];
  assign N1910 = N1909 | i[2041];
  assign N1909 = N1908 | i[2042];
  assign N1908 = N1907 | i[2043];
  assign N1907 = N1906 | i[2044];
  assign N1906 = N1905 | i[2045];
  assign N1905 = i[2047] | i[2046];
  assign o[16] = ~N2158;
  assign N2158 = N2157 | i[2048];
  assign N2157 = N2156 | i[2049];
  assign N2156 = N2155 | i[2050];
  assign N2155 = N2154 | i[2051];
  assign N2154 = N2153 | i[2052];
  assign N2153 = N2152 | i[2053];
  assign N2152 = N2151 | i[2054];
  assign N2151 = N2150 | i[2055];
  assign N2150 = N2149 | i[2056];
  assign N2149 = N2148 | i[2057];
  assign N2148 = N2147 | i[2058];
  assign N2147 = N2146 | i[2059];
  assign N2146 = N2145 | i[2060];
  assign N2145 = N2144 | i[2061];
  assign N2144 = N2143 | i[2062];
  assign N2143 = N2142 | i[2063];
  assign N2142 = N2141 | i[2064];
  assign N2141 = N2140 | i[2065];
  assign N2140 = N2139 | i[2066];
  assign N2139 = N2138 | i[2067];
  assign N2138 = N2137 | i[2068];
  assign N2137 = N2136 | i[2069];
  assign N2136 = N2135 | i[2070];
  assign N2135 = N2134 | i[2071];
  assign N2134 = N2133 | i[2072];
  assign N2133 = N2132 | i[2073];
  assign N2132 = N2131 | i[2074];
  assign N2131 = N2130 | i[2075];
  assign N2130 = N2129 | i[2076];
  assign N2129 = N2128 | i[2077];
  assign N2128 = N2127 | i[2078];
  assign N2127 = N2126 | i[2079];
  assign N2126 = N2125 | i[2080];
  assign N2125 = N2124 | i[2081];
  assign N2124 = N2123 | i[2082];
  assign N2123 = N2122 | i[2083];
  assign N2122 = N2121 | i[2084];
  assign N2121 = N2120 | i[2085];
  assign N2120 = N2119 | i[2086];
  assign N2119 = N2118 | i[2087];
  assign N2118 = N2117 | i[2088];
  assign N2117 = N2116 | i[2089];
  assign N2116 = N2115 | i[2090];
  assign N2115 = N2114 | i[2091];
  assign N2114 = N2113 | i[2092];
  assign N2113 = N2112 | i[2093];
  assign N2112 = N2111 | i[2094];
  assign N2111 = N2110 | i[2095];
  assign N2110 = N2109 | i[2096];
  assign N2109 = N2108 | i[2097];
  assign N2108 = N2107 | i[2098];
  assign N2107 = N2106 | i[2099];
  assign N2106 = N2105 | i[2100];
  assign N2105 = N2104 | i[2101];
  assign N2104 = N2103 | i[2102];
  assign N2103 = N2102 | i[2103];
  assign N2102 = N2101 | i[2104];
  assign N2101 = N2100 | i[2105];
  assign N2100 = N2099 | i[2106];
  assign N2099 = N2098 | i[2107];
  assign N2098 = N2097 | i[2108];
  assign N2097 = N2096 | i[2109];
  assign N2096 = N2095 | i[2110];
  assign N2095 = N2094 | i[2111];
  assign N2094 = N2093 | i[2112];
  assign N2093 = N2092 | i[2113];
  assign N2092 = N2091 | i[2114];
  assign N2091 = N2090 | i[2115];
  assign N2090 = N2089 | i[2116];
  assign N2089 = N2088 | i[2117];
  assign N2088 = N2087 | i[2118];
  assign N2087 = N2086 | i[2119];
  assign N2086 = N2085 | i[2120];
  assign N2085 = N2084 | i[2121];
  assign N2084 = N2083 | i[2122];
  assign N2083 = N2082 | i[2123];
  assign N2082 = N2081 | i[2124];
  assign N2081 = N2080 | i[2125];
  assign N2080 = N2079 | i[2126];
  assign N2079 = N2078 | i[2127];
  assign N2078 = N2077 | i[2128];
  assign N2077 = N2076 | i[2129];
  assign N2076 = N2075 | i[2130];
  assign N2075 = N2074 | i[2131];
  assign N2074 = N2073 | i[2132];
  assign N2073 = N2072 | i[2133];
  assign N2072 = N2071 | i[2134];
  assign N2071 = N2070 | i[2135];
  assign N2070 = N2069 | i[2136];
  assign N2069 = N2068 | i[2137];
  assign N2068 = N2067 | i[2138];
  assign N2067 = N2066 | i[2139];
  assign N2066 = N2065 | i[2140];
  assign N2065 = N2064 | i[2141];
  assign N2064 = N2063 | i[2142];
  assign N2063 = N2062 | i[2143];
  assign N2062 = N2061 | i[2144];
  assign N2061 = N2060 | i[2145];
  assign N2060 = N2059 | i[2146];
  assign N2059 = N2058 | i[2147];
  assign N2058 = N2057 | i[2148];
  assign N2057 = N2056 | i[2149];
  assign N2056 = N2055 | i[2150];
  assign N2055 = N2054 | i[2151];
  assign N2054 = N2053 | i[2152];
  assign N2053 = N2052 | i[2153];
  assign N2052 = N2051 | i[2154];
  assign N2051 = N2050 | i[2155];
  assign N2050 = N2049 | i[2156];
  assign N2049 = N2048 | i[2157];
  assign N2048 = N2047 | i[2158];
  assign N2047 = N2046 | i[2159];
  assign N2046 = N2045 | i[2160];
  assign N2045 = N2044 | i[2161];
  assign N2044 = N2043 | i[2162];
  assign N2043 = N2042 | i[2163];
  assign N2042 = N2041 | i[2164];
  assign N2041 = N2040 | i[2165];
  assign N2040 = N2039 | i[2166];
  assign N2039 = N2038 | i[2167];
  assign N2038 = N2037 | i[2168];
  assign N2037 = N2036 | i[2169];
  assign N2036 = N2035 | i[2170];
  assign N2035 = N2034 | i[2171];
  assign N2034 = N2033 | i[2172];
  assign N2033 = N2032 | i[2173];
  assign N2032 = i[2175] | i[2174];
  assign o[17] = ~N2285;
  assign N2285 = N2284 | i[2176];
  assign N2284 = N2283 | i[2177];
  assign N2283 = N2282 | i[2178];
  assign N2282 = N2281 | i[2179];
  assign N2281 = N2280 | i[2180];
  assign N2280 = N2279 | i[2181];
  assign N2279 = N2278 | i[2182];
  assign N2278 = N2277 | i[2183];
  assign N2277 = N2276 | i[2184];
  assign N2276 = N2275 | i[2185];
  assign N2275 = N2274 | i[2186];
  assign N2274 = N2273 | i[2187];
  assign N2273 = N2272 | i[2188];
  assign N2272 = N2271 | i[2189];
  assign N2271 = N2270 | i[2190];
  assign N2270 = N2269 | i[2191];
  assign N2269 = N2268 | i[2192];
  assign N2268 = N2267 | i[2193];
  assign N2267 = N2266 | i[2194];
  assign N2266 = N2265 | i[2195];
  assign N2265 = N2264 | i[2196];
  assign N2264 = N2263 | i[2197];
  assign N2263 = N2262 | i[2198];
  assign N2262 = N2261 | i[2199];
  assign N2261 = N2260 | i[2200];
  assign N2260 = N2259 | i[2201];
  assign N2259 = N2258 | i[2202];
  assign N2258 = N2257 | i[2203];
  assign N2257 = N2256 | i[2204];
  assign N2256 = N2255 | i[2205];
  assign N2255 = N2254 | i[2206];
  assign N2254 = N2253 | i[2207];
  assign N2253 = N2252 | i[2208];
  assign N2252 = N2251 | i[2209];
  assign N2251 = N2250 | i[2210];
  assign N2250 = N2249 | i[2211];
  assign N2249 = N2248 | i[2212];
  assign N2248 = N2247 | i[2213];
  assign N2247 = N2246 | i[2214];
  assign N2246 = N2245 | i[2215];
  assign N2245 = N2244 | i[2216];
  assign N2244 = N2243 | i[2217];
  assign N2243 = N2242 | i[2218];
  assign N2242 = N2241 | i[2219];
  assign N2241 = N2240 | i[2220];
  assign N2240 = N2239 | i[2221];
  assign N2239 = N2238 | i[2222];
  assign N2238 = N2237 | i[2223];
  assign N2237 = N2236 | i[2224];
  assign N2236 = N2235 | i[2225];
  assign N2235 = N2234 | i[2226];
  assign N2234 = N2233 | i[2227];
  assign N2233 = N2232 | i[2228];
  assign N2232 = N2231 | i[2229];
  assign N2231 = N2230 | i[2230];
  assign N2230 = N2229 | i[2231];
  assign N2229 = N2228 | i[2232];
  assign N2228 = N2227 | i[2233];
  assign N2227 = N2226 | i[2234];
  assign N2226 = N2225 | i[2235];
  assign N2225 = N2224 | i[2236];
  assign N2224 = N2223 | i[2237];
  assign N2223 = N2222 | i[2238];
  assign N2222 = N2221 | i[2239];
  assign N2221 = N2220 | i[2240];
  assign N2220 = N2219 | i[2241];
  assign N2219 = N2218 | i[2242];
  assign N2218 = N2217 | i[2243];
  assign N2217 = N2216 | i[2244];
  assign N2216 = N2215 | i[2245];
  assign N2215 = N2214 | i[2246];
  assign N2214 = N2213 | i[2247];
  assign N2213 = N2212 | i[2248];
  assign N2212 = N2211 | i[2249];
  assign N2211 = N2210 | i[2250];
  assign N2210 = N2209 | i[2251];
  assign N2209 = N2208 | i[2252];
  assign N2208 = N2207 | i[2253];
  assign N2207 = N2206 | i[2254];
  assign N2206 = N2205 | i[2255];
  assign N2205 = N2204 | i[2256];
  assign N2204 = N2203 | i[2257];
  assign N2203 = N2202 | i[2258];
  assign N2202 = N2201 | i[2259];
  assign N2201 = N2200 | i[2260];
  assign N2200 = N2199 | i[2261];
  assign N2199 = N2198 | i[2262];
  assign N2198 = N2197 | i[2263];
  assign N2197 = N2196 | i[2264];
  assign N2196 = N2195 | i[2265];
  assign N2195 = N2194 | i[2266];
  assign N2194 = N2193 | i[2267];
  assign N2193 = N2192 | i[2268];
  assign N2192 = N2191 | i[2269];
  assign N2191 = N2190 | i[2270];
  assign N2190 = N2189 | i[2271];
  assign N2189 = N2188 | i[2272];
  assign N2188 = N2187 | i[2273];
  assign N2187 = N2186 | i[2274];
  assign N2186 = N2185 | i[2275];
  assign N2185 = N2184 | i[2276];
  assign N2184 = N2183 | i[2277];
  assign N2183 = N2182 | i[2278];
  assign N2182 = N2181 | i[2279];
  assign N2181 = N2180 | i[2280];
  assign N2180 = N2179 | i[2281];
  assign N2179 = N2178 | i[2282];
  assign N2178 = N2177 | i[2283];
  assign N2177 = N2176 | i[2284];
  assign N2176 = N2175 | i[2285];
  assign N2175 = N2174 | i[2286];
  assign N2174 = N2173 | i[2287];
  assign N2173 = N2172 | i[2288];
  assign N2172 = N2171 | i[2289];
  assign N2171 = N2170 | i[2290];
  assign N2170 = N2169 | i[2291];
  assign N2169 = N2168 | i[2292];
  assign N2168 = N2167 | i[2293];
  assign N2167 = N2166 | i[2294];
  assign N2166 = N2165 | i[2295];
  assign N2165 = N2164 | i[2296];
  assign N2164 = N2163 | i[2297];
  assign N2163 = N2162 | i[2298];
  assign N2162 = N2161 | i[2299];
  assign N2161 = N2160 | i[2300];
  assign N2160 = N2159 | i[2301];
  assign N2159 = i[2303] | i[2302];
  assign o[18] = ~N2412;
  assign N2412 = N2411 | i[2304];
  assign N2411 = N2410 | i[2305];
  assign N2410 = N2409 | i[2306];
  assign N2409 = N2408 | i[2307];
  assign N2408 = N2407 | i[2308];
  assign N2407 = N2406 | i[2309];
  assign N2406 = N2405 | i[2310];
  assign N2405 = N2404 | i[2311];
  assign N2404 = N2403 | i[2312];
  assign N2403 = N2402 | i[2313];
  assign N2402 = N2401 | i[2314];
  assign N2401 = N2400 | i[2315];
  assign N2400 = N2399 | i[2316];
  assign N2399 = N2398 | i[2317];
  assign N2398 = N2397 | i[2318];
  assign N2397 = N2396 | i[2319];
  assign N2396 = N2395 | i[2320];
  assign N2395 = N2394 | i[2321];
  assign N2394 = N2393 | i[2322];
  assign N2393 = N2392 | i[2323];
  assign N2392 = N2391 | i[2324];
  assign N2391 = N2390 | i[2325];
  assign N2390 = N2389 | i[2326];
  assign N2389 = N2388 | i[2327];
  assign N2388 = N2387 | i[2328];
  assign N2387 = N2386 | i[2329];
  assign N2386 = N2385 | i[2330];
  assign N2385 = N2384 | i[2331];
  assign N2384 = N2383 | i[2332];
  assign N2383 = N2382 | i[2333];
  assign N2382 = N2381 | i[2334];
  assign N2381 = N2380 | i[2335];
  assign N2380 = N2379 | i[2336];
  assign N2379 = N2378 | i[2337];
  assign N2378 = N2377 | i[2338];
  assign N2377 = N2376 | i[2339];
  assign N2376 = N2375 | i[2340];
  assign N2375 = N2374 | i[2341];
  assign N2374 = N2373 | i[2342];
  assign N2373 = N2372 | i[2343];
  assign N2372 = N2371 | i[2344];
  assign N2371 = N2370 | i[2345];
  assign N2370 = N2369 | i[2346];
  assign N2369 = N2368 | i[2347];
  assign N2368 = N2367 | i[2348];
  assign N2367 = N2366 | i[2349];
  assign N2366 = N2365 | i[2350];
  assign N2365 = N2364 | i[2351];
  assign N2364 = N2363 | i[2352];
  assign N2363 = N2362 | i[2353];
  assign N2362 = N2361 | i[2354];
  assign N2361 = N2360 | i[2355];
  assign N2360 = N2359 | i[2356];
  assign N2359 = N2358 | i[2357];
  assign N2358 = N2357 | i[2358];
  assign N2357 = N2356 | i[2359];
  assign N2356 = N2355 | i[2360];
  assign N2355 = N2354 | i[2361];
  assign N2354 = N2353 | i[2362];
  assign N2353 = N2352 | i[2363];
  assign N2352 = N2351 | i[2364];
  assign N2351 = N2350 | i[2365];
  assign N2350 = N2349 | i[2366];
  assign N2349 = N2348 | i[2367];
  assign N2348 = N2347 | i[2368];
  assign N2347 = N2346 | i[2369];
  assign N2346 = N2345 | i[2370];
  assign N2345 = N2344 | i[2371];
  assign N2344 = N2343 | i[2372];
  assign N2343 = N2342 | i[2373];
  assign N2342 = N2341 | i[2374];
  assign N2341 = N2340 | i[2375];
  assign N2340 = N2339 | i[2376];
  assign N2339 = N2338 | i[2377];
  assign N2338 = N2337 | i[2378];
  assign N2337 = N2336 | i[2379];
  assign N2336 = N2335 | i[2380];
  assign N2335 = N2334 | i[2381];
  assign N2334 = N2333 | i[2382];
  assign N2333 = N2332 | i[2383];
  assign N2332 = N2331 | i[2384];
  assign N2331 = N2330 | i[2385];
  assign N2330 = N2329 | i[2386];
  assign N2329 = N2328 | i[2387];
  assign N2328 = N2327 | i[2388];
  assign N2327 = N2326 | i[2389];
  assign N2326 = N2325 | i[2390];
  assign N2325 = N2324 | i[2391];
  assign N2324 = N2323 | i[2392];
  assign N2323 = N2322 | i[2393];
  assign N2322 = N2321 | i[2394];
  assign N2321 = N2320 | i[2395];
  assign N2320 = N2319 | i[2396];
  assign N2319 = N2318 | i[2397];
  assign N2318 = N2317 | i[2398];
  assign N2317 = N2316 | i[2399];
  assign N2316 = N2315 | i[2400];
  assign N2315 = N2314 | i[2401];
  assign N2314 = N2313 | i[2402];
  assign N2313 = N2312 | i[2403];
  assign N2312 = N2311 | i[2404];
  assign N2311 = N2310 | i[2405];
  assign N2310 = N2309 | i[2406];
  assign N2309 = N2308 | i[2407];
  assign N2308 = N2307 | i[2408];
  assign N2307 = N2306 | i[2409];
  assign N2306 = N2305 | i[2410];
  assign N2305 = N2304 | i[2411];
  assign N2304 = N2303 | i[2412];
  assign N2303 = N2302 | i[2413];
  assign N2302 = N2301 | i[2414];
  assign N2301 = N2300 | i[2415];
  assign N2300 = N2299 | i[2416];
  assign N2299 = N2298 | i[2417];
  assign N2298 = N2297 | i[2418];
  assign N2297 = N2296 | i[2419];
  assign N2296 = N2295 | i[2420];
  assign N2295 = N2294 | i[2421];
  assign N2294 = N2293 | i[2422];
  assign N2293 = N2292 | i[2423];
  assign N2292 = N2291 | i[2424];
  assign N2291 = N2290 | i[2425];
  assign N2290 = N2289 | i[2426];
  assign N2289 = N2288 | i[2427];
  assign N2288 = N2287 | i[2428];
  assign N2287 = N2286 | i[2429];
  assign N2286 = i[2431] | i[2430];
  assign o[19] = ~N2539;
  assign N2539 = N2538 | i[2432];
  assign N2538 = N2537 | i[2433];
  assign N2537 = N2536 | i[2434];
  assign N2536 = N2535 | i[2435];
  assign N2535 = N2534 | i[2436];
  assign N2534 = N2533 | i[2437];
  assign N2533 = N2532 | i[2438];
  assign N2532 = N2531 | i[2439];
  assign N2531 = N2530 | i[2440];
  assign N2530 = N2529 | i[2441];
  assign N2529 = N2528 | i[2442];
  assign N2528 = N2527 | i[2443];
  assign N2527 = N2526 | i[2444];
  assign N2526 = N2525 | i[2445];
  assign N2525 = N2524 | i[2446];
  assign N2524 = N2523 | i[2447];
  assign N2523 = N2522 | i[2448];
  assign N2522 = N2521 | i[2449];
  assign N2521 = N2520 | i[2450];
  assign N2520 = N2519 | i[2451];
  assign N2519 = N2518 | i[2452];
  assign N2518 = N2517 | i[2453];
  assign N2517 = N2516 | i[2454];
  assign N2516 = N2515 | i[2455];
  assign N2515 = N2514 | i[2456];
  assign N2514 = N2513 | i[2457];
  assign N2513 = N2512 | i[2458];
  assign N2512 = N2511 | i[2459];
  assign N2511 = N2510 | i[2460];
  assign N2510 = N2509 | i[2461];
  assign N2509 = N2508 | i[2462];
  assign N2508 = N2507 | i[2463];
  assign N2507 = N2506 | i[2464];
  assign N2506 = N2505 | i[2465];
  assign N2505 = N2504 | i[2466];
  assign N2504 = N2503 | i[2467];
  assign N2503 = N2502 | i[2468];
  assign N2502 = N2501 | i[2469];
  assign N2501 = N2500 | i[2470];
  assign N2500 = N2499 | i[2471];
  assign N2499 = N2498 | i[2472];
  assign N2498 = N2497 | i[2473];
  assign N2497 = N2496 | i[2474];
  assign N2496 = N2495 | i[2475];
  assign N2495 = N2494 | i[2476];
  assign N2494 = N2493 | i[2477];
  assign N2493 = N2492 | i[2478];
  assign N2492 = N2491 | i[2479];
  assign N2491 = N2490 | i[2480];
  assign N2490 = N2489 | i[2481];
  assign N2489 = N2488 | i[2482];
  assign N2488 = N2487 | i[2483];
  assign N2487 = N2486 | i[2484];
  assign N2486 = N2485 | i[2485];
  assign N2485 = N2484 | i[2486];
  assign N2484 = N2483 | i[2487];
  assign N2483 = N2482 | i[2488];
  assign N2482 = N2481 | i[2489];
  assign N2481 = N2480 | i[2490];
  assign N2480 = N2479 | i[2491];
  assign N2479 = N2478 | i[2492];
  assign N2478 = N2477 | i[2493];
  assign N2477 = N2476 | i[2494];
  assign N2476 = N2475 | i[2495];
  assign N2475 = N2474 | i[2496];
  assign N2474 = N2473 | i[2497];
  assign N2473 = N2472 | i[2498];
  assign N2472 = N2471 | i[2499];
  assign N2471 = N2470 | i[2500];
  assign N2470 = N2469 | i[2501];
  assign N2469 = N2468 | i[2502];
  assign N2468 = N2467 | i[2503];
  assign N2467 = N2466 | i[2504];
  assign N2466 = N2465 | i[2505];
  assign N2465 = N2464 | i[2506];
  assign N2464 = N2463 | i[2507];
  assign N2463 = N2462 | i[2508];
  assign N2462 = N2461 | i[2509];
  assign N2461 = N2460 | i[2510];
  assign N2460 = N2459 | i[2511];
  assign N2459 = N2458 | i[2512];
  assign N2458 = N2457 | i[2513];
  assign N2457 = N2456 | i[2514];
  assign N2456 = N2455 | i[2515];
  assign N2455 = N2454 | i[2516];
  assign N2454 = N2453 | i[2517];
  assign N2453 = N2452 | i[2518];
  assign N2452 = N2451 | i[2519];
  assign N2451 = N2450 | i[2520];
  assign N2450 = N2449 | i[2521];
  assign N2449 = N2448 | i[2522];
  assign N2448 = N2447 | i[2523];
  assign N2447 = N2446 | i[2524];
  assign N2446 = N2445 | i[2525];
  assign N2445 = N2444 | i[2526];
  assign N2444 = N2443 | i[2527];
  assign N2443 = N2442 | i[2528];
  assign N2442 = N2441 | i[2529];
  assign N2441 = N2440 | i[2530];
  assign N2440 = N2439 | i[2531];
  assign N2439 = N2438 | i[2532];
  assign N2438 = N2437 | i[2533];
  assign N2437 = N2436 | i[2534];
  assign N2436 = N2435 | i[2535];
  assign N2435 = N2434 | i[2536];
  assign N2434 = N2433 | i[2537];
  assign N2433 = N2432 | i[2538];
  assign N2432 = N2431 | i[2539];
  assign N2431 = N2430 | i[2540];
  assign N2430 = N2429 | i[2541];
  assign N2429 = N2428 | i[2542];
  assign N2428 = N2427 | i[2543];
  assign N2427 = N2426 | i[2544];
  assign N2426 = N2425 | i[2545];
  assign N2425 = N2424 | i[2546];
  assign N2424 = N2423 | i[2547];
  assign N2423 = N2422 | i[2548];
  assign N2422 = N2421 | i[2549];
  assign N2421 = N2420 | i[2550];
  assign N2420 = N2419 | i[2551];
  assign N2419 = N2418 | i[2552];
  assign N2418 = N2417 | i[2553];
  assign N2417 = N2416 | i[2554];
  assign N2416 = N2415 | i[2555];
  assign N2415 = N2414 | i[2556];
  assign N2414 = N2413 | i[2557];
  assign N2413 = i[2559] | i[2558];

endmodule

