

module top
(
  binary_i,
  gray_o
);

  input [127:0] binary_i;
  output [127:0] gray_o;

  bsg_binary_plus_one_to_gray
  wrapper
  (
    .binary_i(binary_i),
    .gray_o(gray_o)
  );


endmodule



module bsg_scan_width_p128_and_p1_lo_to_hi_p1
(
  i,
  o
);

  input [127:0] i;
  output [127:0] o;
  wire [127:0] o;
  wire t_3__127_,t_3__126_,t_3__125_,t_3__124_,t_3__123_,t_3__122_,t_3__121_,t_3__120_,
  t_3__119_,t_3__118_,t_3__117_,t_3__116_,t_3__115_,t_3__114_,t_3__113_,t_3__112_,
  t_3__111_,t_3__110_,t_3__109_,t_3__108_,t_3__107_,t_3__106_,t_3__105_,t_3__104_,
  t_3__103_,t_3__102_,t_3__101_,t_3__100_,t_3__99_,t_3__98_,t_3__97_,t_3__96_,
  t_3__95_,t_3__94_,t_3__93_,t_3__92_,t_3__91_,t_3__90_,t_3__89_,t_3__88_,t_3__87_,
  t_3__86_,t_3__85_,t_3__84_,t_3__83_,t_3__82_,t_3__81_,t_3__80_,t_3__79_,t_3__78_,
  t_3__77_,t_3__76_,t_3__75_,t_3__74_,t_3__73_,t_3__72_,t_3__71_,t_3__70_,t_3__69_,
  t_3__68_,t_3__67_,t_3__66_,t_3__65_,t_3__64_,t_3__63_,t_3__62_,t_3__61_,t_3__60_,
  t_3__59_,t_3__58_,t_3__57_,t_3__56_,t_3__55_,t_3__54_,t_3__53_,t_3__52_,
  t_3__51_,t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,t_3__45_,t_3__44_,t_3__43_,
  t_3__42_,t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,t_3__36_,t_3__35_,t_3__34_,
  t_3__33_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,t_3__26_,t_3__25_,
  t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,t_3__17_,t_3__16_,
  t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,
  t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_2__127_,t_2__126_,t_2__125_,
  t_2__124_,t_2__123_,t_2__122_,t_2__121_,t_2__120_,t_2__119_,t_2__118_,t_2__117_,
  t_2__116_,t_2__115_,t_2__114_,t_2__113_,t_2__112_,t_2__111_,t_2__110_,t_2__109_,
  t_2__108_,t_2__107_,t_2__106_,t_2__105_,t_2__104_,t_2__103_,t_2__102_,t_2__101_,
  t_2__100_,t_2__99_,t_2__98_,t_2__97_,t_2__96_,t_2__95_,t_2__94_,t_2__93_,
  t_2__92_,t_2__91_,t_2__90_,t_2__89_,t_2__88_,t_2__87_,t_2__86_,t_2__85_,t_2__84_,
  t_2__83_,t_2__82_,t_2__81_,t_2__80_,t_2__79_,t_2__78_,t_2__77_,t_2__76_,t_2__75_,
  t_2__74_,t_2__73_,t_2__72_,t_2__71_,t_2__70_,t_2__69_,t_2__68_,t_2__67_,t_2__66_,
  t_2__65_,t_2__64_,t_2__63_,t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,t_2__57_,
  t_2__56_,t_2__55_,t_2__54_,t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,t_2__48_,
  t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,t_2__39_,
  t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,t_2__30_,
  t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,
  t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,
  t_2__2_,t_2__1_,t_2__0_,t_1__127_,t_1__126_,t_1__125_,t_1__124_,t_1__123_,t_1__122_,
  t_1__121_,t_1__120_,t_1__119_,t_1__118_,t_1__117_,t_1__116_,t_1__115_,t_1__114_,
  t_1__113_,t_1__112_,t_1__111_,t_1__110_,t_1__109_,t_1__108_,t_1__107_,t_1__106_,
  t_1__105_,t_1__104_,t_1__103_,t_1__102_,t_1__101_,t_1__100_,t_1__99_,t_1__98_,
  t_1__97_,t_1__96_,t_1__95_,t_1__94_,t_1__93_,t_1__92_,t_1__91_,t_1__90_,t_1__89_,
  t_1__88_,t_1__87_,t_1__86_,t_1__85_,t_1__84_,t_1__83_,t_1__82_,t_1__81_,t_1__80_,
  t_1__79_,t_1__78_,t_1__77_,t_1__76_,t_1__75_,t_1__74_,t_1__73_,t_1__72_,
  t_1__71_,t_1__70_,t_1__69_,t_1__68_,t_1__67_,t_1__66_,t_1__65_,t_1__64_,t_1__63_,
  t_1__62_,t_1__61_,t_1__60_,t_1__59_,t_1__58_,t_1__57_,t_1__56_,t_1__55_,t_1__54_,
  t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,t_1__48_,t_1__47_,t_1__46_,t_1__45_,
  t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,t_1__39_,t_1__38_,t_1__37_,t_1__36_,
  t_1__35_,t_1__34_,t_1__33_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,t_1__27_,
  t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,t_1__18_,
  t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,t_1__9_,
  t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_,t_6__127_,
  t_6__126_,t_6__125_,t_6__124_,t_6__123_,t_6__122_,t_6__121_,t_6__120_,t_6__119_,
  t_6__118_,t_6__117_,t_6__116_,t_6__115_,t_6__114_,t_6__113_,t_6__112_,t_6__111_,
  t_6__110_,t_6__109_,t_6__108_,t_6__107_,t_6__106_,t_6__105_,t_6__104_,t_6__103_,
  t_6__102_,t_6__101_,t_6__100_,t_6__99_,t_6__98_,t_6__97_,t_6__96_,t_6__95_,
  t_6__94_,t_6__93_,t_6__92_,t_6__91_,t_6__90_,t_6__89_,t_6__88_,t_6__87_,t_6__86_,
  t_6__85_,t_6__84_,t_6__83_,t_6__82_,t_6__81_,t_6__80_,t_6__79_,t_6__78_,t_6__77_,
  t_6__76_,t_6__75_,t_6__74_,t_6__73_,t_6__72_,t_6__71_,t_6__70_,t_6__69_,t_6__68_,
  t_6__67_,t_6__66_,t_6__65_,t_6__64_,t_6__63_,t_6__62_,t_6__61_,t_6__60_,t_6__59_,
  t_6__58_,t_6__57_,t_6__56_,t_6__55_,t_6__54_,t_6__53_,t_6__52_,t_6__51_,t_6__50_,
  t_6__49_,t_6__48_,t_6__47_,t_6__46_,t_6__45_,t_6__44_,t_6__43_,t_6__42_,
  t_6__41_,t_6__40_,t_6__39_,t_6__38_,t_6__37_,t_6__36_,t_6__35_,t_6__34_,t_6__33_,
  t_6__32_,t_6__31_,t_6__30_,t_6__29_,t_6__28_,t_6__27_,t_6__26_,t_6__25_,t_6__24_,
  t_6__23_,t_6__22_,t_6__21_,t_6__20_,t_6__19_,t_6__18_,t_6__17_,t_6__16_,t_6__15_,
  t_6__14_,t_6__13_,t_6__12_,t_6__11_,t_6__10_,t_6__9_,t_6__8_,t_6__7_,t_6__6_,t_6__5_,
  t_6__4_,t_6__3_,t_6__2_,t_6__1_,t_6__0_,t_5__127_,t_5__126_,t_5__125_,t_5__124_,
  t_5__123_,t_5__122_,t_5__121_,t_5__120_,t_5__119_,t_5__118_,t_5__117_,t_5__116_,
  t_5__115_,t_5__114_,t_5__113_,t_5__112_,t_5__111_,t_5__110_,t_5__109_,t_5__108_,
  t_5__107_,t_5__106_,t_5__105_,t_5__104_,t_5__103_,t_5__102_,t_5__101_,t_5__100_,
  t_5__99_,t_5__98_,t_5__97_,t_5__96_,t_5__95_,t_5__94_,t_5__93_,t_5__92_,
  t_5__91_,t_5__90_,t_5__89_,t_5__88_,t_5__87_,t_5__86_,t_5__85_,t_5__84_,t_5__83_,
  t_5__82_,t_5__81_,t_5__80_,t_5__79_,t_5__78_,t_5__77_,t_5__76_,t_5__75_,t_5__74_,
  t_5__73_,t_5__72_,t_5__71_,t_5__70_,t_5__69_,t_5__68_,t_5__67_,t_5__66_,t_5__65_,
  t_5__64_,t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,t_5__58_,t_5__57_,t_5__56_,
  t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,
  t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,
  t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,
  t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,
  t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,
  t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,
  t_5__1_,t_5__0_,t_4__127_,t_4__126_,t_4__125_,t_4__124_,t_4__123_,t_4__122_,t_4__121_,
  t_4__120_,t_4__119_,t_4__118_,t_4__117_,t_4__116_,t_4__115_,t_4__114_,t_4__113_,
  t_4__112_,t_4__111_,t_4__110_,t_4__109_,t_4__108_,t_4__107_,t_4__106_,t_4__105_,
  t_4__104_,t_4__103_,t_4__102_,t_4__101_,t_4__100_,t_4__99_,t_4__98_,t_4__97_,
  t_4__96_,t_4__95_,t_4__94_,t_4__93_,t_4__92_,t_4__91_,t_4__90_,t_4__89_,t_4__88_,
  t_4__87_,t_4__86_,t_4__85_,t_4__84_,t_4__83_,t_4__82_,t_4__81_,t_4__80_,t_4__79_,
  t_4__78_,t_4__77_,t_4__76_,t_4__75_,t_4__74_,t_4__73_,t_4__72_,t_4__71_,t_4__70_,
  t_4__69_,t_4__68_,t_4__67_,t_4__66_,t_4__65_,t_4__64_,t_4__63_,t_4__62_,
  t_4__61_,t_4__60_,t_4__59_,t_4__58_,t_4__57_,t_4__56_,t_4__55_,t_4__54_,t_4__53_,
  t_4__52_,t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,
  t_4__43_,t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,
  t_4__34_,t_4__33_,t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,
  t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,
  t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,
  t_4__7_,t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_;
  assign t_1__127_ = i[0] & 1'b1;
  assign t_1__126_ = i[1] & i[0];
  assign t_1__125_ = i[2] & i[1];
  assign t_1__124_ = i[3] & i[2];
  assign t_1__123_ = i[4] & i[3];
  assign t_1__122_ = i[5] & i[4];
  assign t_1__121_ = i[6] & i[5];
  assign t_1__120_ = i[7] & i[6];
  assign t_1__119_ = i[8] & i[7];
  assign t_1__118_ = i[9] & i[8];
  assign t_1__117_ = i[10] & i[9];
  assign t_1__116_ = i[11] & i[10];
  assign t_1__115_ = i[12] & i[11];
  assign t_1__114_ = i[13] & i[12];
  assign t_1__113_ = i[14] & i[13];
  assign t_1__112_ = i[15] & i[14];
  assign t_1__111_ = i[16] & i[15];
  assign t_1__110_ = i[17] & i[16];
  assign t_1__109_ = i[18] & i[17];
  assign t_1__108_ = i[19] & i[18];
  assign t_1__107_ = i[20] & i[19];
  assign t_1__106_ = i[21] & i[20];
  assign t_1__105_ = i[22] & i[21];
  assign t_1__104_ = i[23] & i[22];
  assign t_1__103_ = i[24] & i[23];
  assign t_1__102_ = i[25] & i[24];
  assign t_1__101_ = i[26] & i[25];
  assign t_1__100_ = i[27] & i[26];
  assign t_1__99_ = i[28] & i[27];
  assign t_1__98_ = i[29] & i[28];
  assign t_1__97_ = i[30] & i[29];
  assign t_1__96_ = i[31] & i[30];
  assign t_1__95_ = i[32] & i[31];
  assign t_1__94_ = i[33] & i[32];
  assign t_1__93_ = i[34] & i[33];
  assign t_1__92_ = i[35] & i[34];
  assign t_1__91_ = i[36] & i[35];
  assign t_1__90_ = i[37] & i[36];
  assign t_1__89_ = i[38] & i[37];
  assign t_1__88_ = i[39] & i[38];
  assign t_1__87_ = i[40] & i[39];
  assign t_1__86_ = i[41] & i[40];
  assign t_1__85_ = i[42] & i[41];
  assign t_1__84_ = i[43] & i[42];
  assign t_1__83_ = i[44] & i[43];
  assign t_1__82_ = i[45] & i[44];
  assign t_1__81_ = i[46] & i[45];
  assign t_1__80_ = i[47] & i[46];
  assign t_1__79_ = i[48] & i[47];
  assign t_1__78_ = i[49] & i[48];
  assign t_1__77_ = i[50] & i[49];
  assign t_1__76_ = i[51] & i[50];
  assign t_1__75_ = i[52] & i[51];
  assign t_1__74_ = i[53] & i[52];
  assign t_1__73_ = i[54] & i[53];
  assign t_1__72_ = i[55] & i[54];
  assign t_1__71_ = i[56] & i[55];
  assign t_1__70_ = i[57] & i[56];
  assign t_1__69_ = i[58] & i[57];
  assign t_1__68_ = i[59] & i[58];
  assign t_1__67_ = i[60] & i[59];
  assign t_1__66_ = i[61] & i[60];
  assign t_1__65_ = i[62] & i[61];
  assign t_1__64_ = i[63] & i[62];
  assign t_1__63_ = i[64] & i[63];
  assign t_1__62_ = i[65] & i[64];
  assign t_1__61_ = i[66] & i[65];
  assign t_1__60_ = i[67] & i[66];
  assign t_1__59_ = i[68] & i[67];
  assign t_1__58_ = i[69] & i[68];
  assign t_1__57_ = i[70] & i[69];
  assign t_1__56_ = i[71] & i[70];
  assign t_1__55_ = i[72] & i[71];
  assign t_1__54_ = i[73] & i[72];
  assign t_1__53_ = i[74] & i[73];
  assign t_1__52_ = i[75] & i[74];
  assign t_1__51_ = i[76] & i[75];
  assign t_1__50_ = i[77] & i[76];
  assign t_1__49_ = i[78] & i[77];
  assign t_1__48_ = i[79] & i[78];
  assign t_1__47_ = i[80] & i[79];
  assign t_1__46_ = i[81] & i[80];
  assign t_1__45_ = i[82] & i[81];
  assign t_1__44_ = i[83] & i[82];
  assign t_1__43_ = i[84] & i[83];
  assign t_1__42_ = i[85] & i[84];
  assign t_1__41_ = i[86] & i[85];
  assign t_1__40_ = i[87] & i[86];
  assign t_1__39_ = i[88] & i[87];
  assign t_1__38_ = i[89] & i[88];
  assign t_1__37_ = i[90] & i[89];
  assign t_1__36_ = i[91] & i[90];
  assign t_1__35_ = i[92] & i[91];
  assign t_1__34_ = i[93] & i[92];
  assign t_1__33_ = i[94] & i[93];
  assign t_1__32_ = i[95] & i[94];
  assign t_1__31_ = i[96] & i[95];
  assign t_1__30_ = i[97] & i[96];
  assign t_1__29_ = i[98] & i[97];
  assign t_1__28_ = i[99] & i[98];
  assign t_1__27_ = i[100] & i[99];
  assign t_1__26_ = i[101] & i[100];
  assign t_1__25_ = i[102] & i[101];
  assign t_1__24_ = i[103] & i[102];
  assign t_1__23_ = i[104] & i[103];
  assign t_1__22_ = i[105] & i[104];
  assign t_1__21_ = i[106] & i[105];
  assign t_1__20_ = i[107] & i[106];
  assign t_1__19_ = i[108] & i[107];
  assign t_1__18_ = i[109] & i[108];
  assign t_1__17_ = i[110] & i[109];
  assign t_1__16_ = i[111] & i[110];
  assign t_1__15_ = i[112] & i[111];
  assign t_1__14_ = i[113] & i[112];
  assign t_1__13_ = i[114] & i[113];
  assign t_1__12_ = i[115] & i[114];
  assign t_1__11_ = i[116] & i[115];
  assign t_1__10_ = i[117] & i[116];
  assign t_1__9_ = i[118] & i[117];
  assign t_1__8_ = i[119] & i[118];
  assign t_1__7_ = i[120] & i[119];
  assign t_1__6_ = i[121] & i[120];
  assign t_1__5_ = i[122] & i[121];
  assign t_1__4_ = i[123] & i[122];
  assign t_1__3_ = i[124] & i[123];
  assign t_1__2_ = i[125] & i[124];
  assign t_1__1_ = i[126] & i[125];
  assign t_1__0_ = i[127] & i[126];
  assign t_2__127_ = t_1__127_ & 1'b1;
  assign t_2__126_ = t_1__126_ & 1'b1;
  assign t_2__125_ = t_1__125_ & t_1__127_;
  assign t_2__124_ = t_1__124_ & t_1__126_;
  assign t_2__123_ = t_1__123_ & t_1__125_;
  assign t_2__122_ = t_1__122_ & t_1__124_;
  assign t_2__121_ = t_1__121_ & t_1__123_;
  assign t_2__120_ = t_1__120_ & t_1__122_;
  assign t_2__119_ = t_1__119_ & t_1__121_;
  assign t_2__118_ = t_1__118_ & t_1__120_;
  assign t_2__117_ = t_1__117_ & t_1__119_;
  assign t_2__116_ = t_1__116_ & t_1__118_;
  assign t_2__115_ = t_1__115_ & t_1__117_;
  assign t_2__114_ = t_1__114_ & t_1__116_;
  assign t_2__113_ = t_1__113_ & t_1__115_;
  assign t_2__112_ = t_1__112_ & t_1__114_;
  assign t_2__111_ = t_1__111_ & t_1__113_;
  assign t_2__110_ = t_1__110_ & t_1__112_;
  assign t_2__109_ = t_1__109_ & t_1__111_;
  assign t_2__108_ = t_1__108_ & t_1__110_;
  assign t_2__107_ = t_1__107_ & t_1__109_;
  assign t_2__106_ = t_1__106_ & t_1__108_;
  assign t_2__105_ = t_1__105_ & t_1__107_;
  assign t_2__104_ = t_1__104_ & t_1__106_;
  assign t_2__103_ = t_1__103_ & t_1__105_;
  assign t_2__102_ = t_1__102_ & t_1__104_;
  assign t_2__101_ = t_1__101_ & t_1__103_;
  assign t_2__100_ = t_1__100_ & t_1__102_;
  assign t_2__99_ = t_1__99_ & t_1__101_;
  assign t_2__98_ = t_1__98_ & t_1__100_;
  assign t_2__97_ = t_1__97_ & t_1__99_;
  assign t_2__96_ = t_1__96_ & t_1__98_;
  assign t_2__95_ = t_1__95_ & t_1__97_;
  assign t_2__94_ = t_1__94_ & t_1__96_;
  assign t_2__93_ = t_1__93_ & t_1__95_;
  assign t_2__92_ = t_1__92_ & t_1__94_;
  assign t_2__91_ = t_1__91_ & t_1__93_;
  assign t_2__90_ = t_1__90_ & t_1__92_;
  assign t_2__89_ = t_1__89_ & t_1__91_;
  assign t_2__88_ = t_1__88_ & t_1__90_;
  assign t_2__87_ = t_1__87_ & t_1__89_;
  assign t_2__86_ = t_1__86_ & t_1__88_;
  assign t_2__85_ = t_1__85_ & t_1__87_;
  assign t_2__84_ = t_1__84_ & t_1__86_;
  assign t_2__83_ = t_1__83_ & t_1__85_;
  assign t_2__82_ = t_1__82_ & t_1__84_;
  assign t_2__81_ = t_1__81_ & t_1__83_;
  assign t_2__80_ = t_1__80_ & t_1__82_;
  assign t_2__79_ = t_1__79_ & t_1__81_;
  assign t_2__78_ = t_1__78_ & t_1__80_;
  assign t_2__77_ = t_1__77_ & t_1__79_;
  assign t_2__76_ = t_1__76_ & t_1__78_;
  assign t_2__75_ = t_1__75_ & t_1__77_;
  assign t_2__74_ = t_1__74_ & t_1__76_;
  assign t_2__73_ = t_1__73_ & t_1__75_;
  assign t_2__72_ = t_1__72_ & t_1__74_;
  assign t_2__71_ = t_1__71_ & t_1__73_;
  assign t_2__70_ = t_1__70_ & t_1__72_;
  assign t_2__69_ = t_1__69_ & t_1__71_;
  assign t_2__68_ = t_1__68_ & t_1__70_;
  assign t_2__67_ = t_1__67_ & t_1__69_;
  assign t_2__66_ = t_1__66_ & t_1__68_;
  assign t_2__65_ = t_1__65_ & t_1__67_;
  assign t_2__64_ = t_1__64_ & t_1__66_;
  assign t_2__63_ = t_1__63_ & t_1__65_;
  assign t_2__62_ = t_1__62_ & t_1__64_;
  assign t_2__61_ = t_1__61_ & t_1__63_;
  assign t_2__60_ = t_1__60_ & t_1__62_;
  assign t_2__59_ = t_1__59_ & t_1__61_;
  assign t_2__58_ = t_1__58_ & t_1__60_;
  assign t_2__57_ = t_1__57_ & t_1__59_;
  assign t_2__56_ = t_1__56_ & t_1__58_;
  assign t_2__55_ = t_1__55_ & t_1__57_;
  assign t_2__54_ = t_1__54_ & t_1__56_;
  assign t_2__53_ = t_1__53_ & t_1__55_;
  assign t_2__52_ = t_1__52_ & t_1__54_;
  assign t_2__51_ = t_1__51_ & t_1__53_;
  assign t_2__50_ = t_1__50_ & t_1__52_;
  assign t_2__49_ = t_1__49_ & t_1__51_;
  assign t_2__48_ = t_1__48_ & t_1__50_;
  assign t_2__47_ = t_1__47_ & t_1__49_;
  assign t_2__46_ = t_1__46_ & t_1__48_;
  assign t_2__45_ = t_1__45_ & t_1__47_;
  assign t_2__44_ = t_1__44_ & t_1__46_;
  assign t_2__43_ = t_1__43_ & t_1__45_;
  assign t_2__42_ = t_1__42_ & t_1__44_;
  assign t_2__41_ = t_1__41_ & t_1__43_;
  assign t_2__40_ = t_1__40_ & t_1__42_;
  assign t_2__39_ = t_1__39_ & t_1__41_;
  assign t_2__38_ = t_1__38_ & t_1__40_;
  assign t_2__37_ = t_1__37_ & t_1__39_;
  assign t_2__36_ = t_1__36_ & t_1__38_;
  assign t_2__35_ = t_1__35_ & t_1__37_;
  assign t_2__34_ = t_1__34_ & t_1__36_;
  assign t_2__33_ = t_1__33_ & t_1__35_;
  assign t_2__32_ = t_1__32_ & t_1__34_;
  assign t_2__31_ = t_1__31_ & t_1__33_;
  assign t_2__30_ = t_1__30_ & t_1__32_;
  assign t_2__29_ = t_1__29_ & t_1__31_;
  assign t_2__28_ = t_1__28_ & t_1__30_;
  assign t_2__27_ = t_1__27_ & t_1__29_;
  assign t_2__26_ = t_1__26_ & t_1__28_;
  assign t_2__25_ = t_1__25_ & t_1__27_;
  assign t_2__24_ = t_1__24_ & t_1__26_;
  assign t_2__23_ = t_1__23_ & t_1__25_;
  assign t_2__22_ = t_1__22_ & t_1__24_;
  assign t_2__21_ = t_1__21_ & t_1__23_;
  assign t_2__20_ = t_1__20_ & t_1__22_;
  assign t_2__19_ = t_1__19_ & t_1__21_;
  assign t_2__18_ = t_1__18_ & t_1__20_;
  assign t_2__17_ = t_1__17_ & t_1__19_;
  assign t_2__16_ = t_1__16_ & t_1__18_;
  assign t_2__15_ = t_1__15_ & t_1__17_;
  assign t_2__14_ = t_1__14_ & t_1__16_;
  assign t_2__13_ = t_1__13_ & t_1__15_;
  assign t_2__12_ = t_1__12_ & t_1__14_;
  assign t_2__11_ = t_1__11_ & t_1__13_;
  assign t_2__10_ = t_1__10_ & t_1__12_;
  assign t_2__9_ = t_1__9_ & t_1__11_;
  assign t_2__8_ = t_1__8_ & t_1__10_;
  assign t_2__7_ = t_1__7_ & t_1__9_;
  assign t_2__6_ = t_1__6_ & t_1__8_;
  assign t_2__5_ = t_1__5_ & t_1__7_;
  assign t_2__4_ = t_1__4_ & t_1__6_;
  assign t_2__3_ = t_1__3_ & t_1__5_;
  assign t_2__2_ = t_1__2_ & t_1__4_;
  assign t_2__1_ = t_1__1_ & t_1__3_;
  assign t_2__0_ = t_1__0_ & t_1__2_;
  assign t_3__127_ = t_2__127_ & 1'b1;
  assign t_3__126_ = t_2__126_ & 1'b1;
  assign t_3__125_ = t_2__125_ & 1'b1;
  assign t_3__124_ = t_2__124_ & 1'b1;
  assign t_3__123_ = t_2__123_ & t_2__127_;
  assign t_3__122_ = t_2__122_ & t_2__126_;
  assign t_3__121_ = t_2__121_ & t_2__125_;
  assign t_3__120_ = t_2__120_ & t_2__124_;
  assign t_3__119_ = t_2__119_ & t_2__123_;
  assign t_3__118_ = t_2__118_ & t_2__122_;
  assign t_3__117_ = t_2__117_ & t_2__121_;
  assign t_3__116_ = t_2__116_ & t_2__120_;
  assign t_3__115_ = t_2__115_ & t_2__119_;
  assign t_3__114_ = t_2__114_ & t_2__118_;
  assign t_3__113_ = t_2__113_ & t_2__117_;
  assign t_3__112_ = t_2__112_ & t_2__116_;
  assign t_3__111_ = t_2__111_ & t_2__115_;
  assign t_3__110_ = t_2__110_ & t_2__114_;
  assign t_3__109_ = t_2__109_ & t_2__113_;
  assign t_3__108_ = t_2__108_ & t_2__112_;
  assign t_3__107_ = t_2__107_ & t_2__111_;
  assign t_3__106_ = t_2__106_ & t_2__110_;
  assign t_3__105_ = t_2__105_ & t_2__109_;
  assign t_3__104_ = t_2__104_ & t_2__108_;
  assign t_3__103_ = t_2__103_ & t_2__107_;
  assign t_3__102_ = t_2__102_ & t_2__106_;
  assign t_3__101_ = t_2__101_ & t_2__105_;
  assign t_3__100_ = t_2__100_ & t_2__104_;
  assign t_3__99_ = t_2__99_ & t_2__103_;
  assign t_3__98_ = t_2__98_ & t_2__102_;
  assign t_3__97_ = t_2__97_ & t_2__101_;
  assign t_3__96_ = t_2__96_ & t_2__100_;
  assign t_3__95_ = t_2__95_ & t_2__99_;
  assign t_3__94_ = t_2__94_ & t_2__98_;
  assign t_3__93_ = t_2__93_ & t_2__97_;
  assign t_3__92_ = t_2__92_ & t_2__96_;
  assign t_3__91_ = t_2__91_ & t_2__95_;
  assign t_3__90_ = t_2__90_ & t_2__94_;
  assign t_3__89_ = t_2__89_ & t_2__93_;
  assign t_3__88_ = t_2__88_ & t_2__92_;
  assign t_3__87_ = t_2__87_ & t_2__91_;
  assign t_3__86_ = t_2__86_ & t_2__90_;
  assign t_3__85_ = t_2__85_ & t_2__89_;
  assign t_3__84_ = t_2__84_ & t_2__88_;
  assign t_3__83_ = t_2__83_ & t_2__87_;
  assign t_3__82_ = t_2__82_ & t_2__86_;
  assign t_3__81_ = t_2__81_ & t_2__85_;
  assign t_3__80_ = t_2__80_ & t_2__84_;
  assign t_3__79_ = t_2__79_ & t_2__83_;
  assign t_3__78_ = t_2__78_ & t_2__82_;
  assign t_3__77_ = t_2__77_ & t_2__81_;
  assign t_3__76_ = t_2__76_ & t_2__80_;
  assign t_3__75_ = t_2__75_ & t_2__79_;
  assign t_3__74_ = t_2__74_ & t_2__78_;
  assign t_3__73_ = t_2__73_ & t_2__77_;
  assign t_3__72_ = t_2__72_ & t_2__76_;
  assign t_3__71_ = t_2__71_ & t_2__75_;
  assign t_3__70_ = t_2__70_ & t_2__74_;
  assign t_3__69_ = t_2__69_ & t_2__73_;
  assign t_3__68_ = t_2__68_ & t_2__72_;
  assign t_3__67_ = t_2__67_ & t_2__71_;
  assign t_3__66_ = t_2__66_ & t_2__70_;
  assign t_3__65_ = t_2__65_ & t_2__69_;
  assign t_3__64_ = t_2__64_ & t_2__68_;
  assign t_3__63_ = t_2__63_ & t_2__67_;
  assign t_3__62_ = t_2__62_ & t_2__66_;
  assign t_3__61_ = t_2__61_ & t_2__65_;
  assign t_3__60_ = t_2__60_ & t_2__64_;
  assign t_3__59_ = t_2__59_ & t_2__63_;
  assign t_3__58_ = t_2__58_ & t_2__62_;
  assign t_3__57_ = t_2__57_ & t_2__61_;
  assign t_3__56_ = t_2__56_ & t_2__60_;
  assign t_3__55_ = t_2__55_ & t_2__59_;
  assign t_3__54_ = t_2__54_ & t_2__58_;
  assign t_3__53_ = t_2__53_ & t_2__57_;
  assign t_3__52_ = t_2__52_ & t_2__56_;
  assign t_3__51_ = t_2__51_ & t_2__55_;
  assign t_3__50_ = t_2__50_ & t_2__54_;
  assign t_3__49_ = t_2__49_ & t_2__53_;
  assign t_3__48_ = t_2__48_ & t_2__52_;
  assign t_3__47_ = t_2__47_ & t_2__51_;
  assign t_3__46_ = t_2__46_ & t_2__50_;
  assign t_3__45_ = t_2__45_ & t_2__49_;
  assign t_3__44_ = t_2__44_ & t_2__48_;
  assign t_3__43_ = t_2__43_ & t_2__47_;
  assign t_3__42_ = t_2__42_ & t_2__46_;
  assign t_3__41_ = t_2__41_ & t_2__45_;
  assign t_3__40_ = t_2__40_ & t_2__44_;
  assign t_3__39_ = t_2__39_ & t_2__43_;
  assign t_3__38_ = t_2__38_ & t_2__42_;
  assign t_3__37_ = t_2__37_ & t_2__41_;
  assign t_3__36_ = t_2__36_ & t_2__40_;
  assign t_3__35_ = t_2__35_ & t_2__39_;
  assign t_3__34_ = t_2__34_ & t_2__38_;
  assign t_3__33_ = t_2__33_ & t_2__37_;
  assign t_3__32_ = t_2__32_ & t_2__36_;
  assign t_3__31_ = t_2__31_ & t_2__35_;
  assign t_3__30_ = t_2__30_ & t_2__34_;
  assign t_3__29_ = t_2__29_ & t_2__33_;
  assign t_3__28_ = t_2__28_ & t_2__32_;
  assign t_3__27_ = t_2__27_ & t_2__31_;
  assign t_3__26_ = t_2__26_ & t_2__30_;
  assign t_3__25_ = t_2__25_ & t_2__29_;
  assign t_3__24_ = t_2__24_ & t_2__28_;
  assign t_3__23_ = t_2__23_ & t_2__27_;
  assign t_3__22_ = t_2__22_ & t_2__26_;
  assign t_3__21_ = t_2__21_ & t_2__25_;
  assign t_3__20_ = t_2__20_ & t_2__24_;
  assign t_3__19_ = t_2__19_ & t_2__23_;
  assign t_3__18_ = t_2__18_ & t_2__22_;
  assign t_3__17_ = t_2__17_ & t_2__21_;
  assign t_3__16_ = t_2__16_ & t_2__20_;
  assign t_3__15_ = t_2__15_ & t_2__19_;
  assign t_3__14_ = t_2__14_ & t_2__18_;
  assign t_3__13_ = t_2__13_ & t_2__17_;
  assign t_3__12_ = t_2__12_ & t_2__16_;
  assign t_3__11_ = t_2__11_ & t_2__15_;
  assign t_3__10_ = t_2__10_ & t_2__14_;
  assign t_3__9_ = t_2__9_ & t_2__13_;
  assign t_3__8_ = t_2__8_ & t_2__12_;
  assign t_3__7_ = t_2__7_ & t_2__11_;
  assign t_3__6_ = t_2__6_ & t_2__10_;
  assign t_3__5_ = t_2__5_ & t_2__9_;
  assign t_3__4_ = t_2__4_ & t_2__8_;
  assign t_3__3_ = t_2__3_ & t_2__7_;
  assign t_3__2_ = t_2__2_ & t_2__6_;
  assign t_3__1_ = t_2__1_ & t_2__5_;
  assign t_3__0_ = t_2__0_ & t_2__4_;
  assign t_4__127_ = t_3__127_ & 1'b1;
  assign t_4__126_ = t_3__126_ & 1'b1;
  assign t_4__125_ = t_3__125_ & 1'b1;
  assign t_4__124_ = t_3__124_ & 1'b1;
  assign t_4__123_ = t_3__123_ & 1'b1;
  assign t_4__122_ = t_3__122_ & 1'b1;
  assign t_4__121_ = t_3__121_ & 1'b1;
  assign t_4__120_ = t_3__120_ & 1'b1;
  assign t_4__119_ = t_3__119_ & t_3__127_;
  assign t_4__118_ = t_3__118_ & t_3__126_;
  assign t_4__117_ = t_3__117_ & t_3__125_;
  assign t_4__116_ = t_3__116_ & t_3__124_;
  assign t_4__115_ = t_3__115_ & t_3__123_;
  assign t_4__114_ = t_3__114_ & t_3__122_;
  assign t_4__113_ = t_3__113_ & t_3__121_;
  assign t_4__112_ = t_3__112_ & t_3__120_;
  assign t_4__111_ = t_3__111_ & t_3__119_;
  assign t_4__110_ = t_3__110_ & t_3__118_;
  assign t_4__109_ = t_3__109_ & t_3__117_;
  assign t_4__108_ = t_3__108_ & t_3__116_;
  assign t_4__107_ = t_3__107_ & t_3__115_;
  assign t_4__106_ = t_3__106_ & t_3__114_;
  assign t_4__105_ = t_3__105_ & t_3__113_;
  assign t_4__104_ = t_3__104_ & t_3__112_;
  assign t_4__103_ = t_3__103_ & t_3__111_;
  assign t_4__102_ = t_3__102_ & t_3__110_;
  assign t_4__101_ = t_3__101_ & t_3__109_;
  assign t_4__100_ = t_3__100_ & t_3__108_;
  assign t_4__99_ = t_3__99_ & t_3__107_;
  assign t_4__98_ = t_3__98_ & t_3__106_;
  assign t_4__97_ = t_3__97_ & t_3__105_;
  assign t_4__96_ = t_3__96_ & t_3__104_;
  assign t_4__95_ = t_3__95_ & t_3__103_;
  assign t_4__94_ = t_3__94_ & t_3__102_;
  assign t_4__93_ = t_3__93_ & t_3__101_;
  assign t_4__92_ = t_3__92_ & t_3__100_;
  assign t_4__91_ = t_3__91_ & t_3__99_;
  assign t_4__90_ = t_3__90_ & t_3__98_;
  assign t_4__89_ = t_3__89_ & t_3__97_;
  assign t_4__88_ = t_3__88_ & t_3__96_;
  assign t_4__87_ = t_3__87_ & t_3__95_;
  assign t_4__86_ = t_3__86_ & t_3__94_;
  assign t_4__85_ = t_3__85_ & t_3__93_;
  assign t_4__84_ = t_3__84_ & t_3__92_;
  assign t_4__83_ = t_3__83_ & t_3__91_;
  assign t_4__82_ = t_3__82_ & t_3__90_;
  assign t_4__81_ = t_3__81_ & t_3__89_;
  assign t_4__80_ = t_3__80_ & t_3__88_;
  assign t_4__79_ = t_3__79_ & t_3__87_;
  assign t_4__78_ = t_3__78_ & t_3__86_;
  assign t_4__77_ = t_3__77_ & t_3__85_;
  assign t_4__76_ = t_3__76_ & t_3__84_;
  assign t_4__75_ = t_3__75_ & t_3__83_;
  assign t_4__74_ = t_3__74_ & t_3__82_;
  assign t_4__73_ = t_3__73_ & t_3__81_;
  assign t_4__72_ = t_3__72_ & t_3__80_;
  assign t_4__71_ = t_3__71_ & t_3__79_;
  assign t_4__70_ = t_3__70_ & t_3__78_;
  assign t_4__69_ = t_3__69_ & t_3__77_;
  assign t_4__68_ = t_3__68_ & t_3__76_;
  assign t_4__67_ = t_3__67_ & t_3__75_;
  assign t_4__66_ = t_3__66_ & t_3__74_;
  assign t_4__65_ = t_3__65_ & t_3__73_;
  assign t_4__64_ = t_3__64_ & t_3__72_;
  assign t_4__63_ = t_3__63_ & t_3__71_;
  assign t_4__62_ = t_3__62_ & t_3__70_;
  assign t_4__61_ = t_3__61_ & t_3__69_;
  assign t_4__60_ = t_3__60_ & t_3__68_;
  assign t_4__59_ = t_3__59_ & t_3__67_;
  assign t_4__58_ = t_3__58_ & t_3__66_;
  assign t_4__57_ = t_3__57_ & t_3__65_;
  assign t_4__56_ = t_3__56_ & t_3__64_;
  assign t_4__55_ = t_3__55_ & t_3__63_;
  assign t_4__54_ = t_3__54_ & t_3__62_;
  assign t_4__53_ = t_3__53_ & t_3__61_;
  assign t_4__52_ = t_3__52_ & t_3__60_;
  assign t_4__51_ = t_3__51_ & t_3__59_;
  assign t_4__50_ = t_3__50_ & t_3__58_;
  assign t_4__49_ = t_3__49_ & t_3__57_;
  assign t_4__48_ = t_3__48_ & t_3__56_;
  assign t_4__47_ = t_3__47_ & t_3__55_;
  assign t_4__46_ = t_3__46_ & t_3__54_;
  assign t_4__45_ = t_3__45_ & t_3__53_;
  assign t_4__44_ = t_3__44_ & t_3__52_;
  assign t_4__43_ = t_3__43_ & t_3__51_;
  assign t_4__42_ = t_3__42_ & t_3__50_;
  assign t_4__41_ = t_3__41_ & t_3__49_;
  assign t_4__40_ = t_3__40_ & t_3__48_;
  assign t_4__39_ = t_3__39_ & t_3__47_;
  assign t_4__38_ = t_3__38_ & t_3__46_;
  assign t_4__37_ = t_3__37_ & t_3__45_;
  assign t_4__36_ = t_3__36_ & t_3__44_;
  assign t_4__35_ = t_3__35_ & t_3__43_;
  assign t_4__34_ = t_3__34_ & t_3__42_;
  assign t_4__33_ = t_3__33_ & t_3__41_;
  assign t_4__32_ = t_3__32_ & t_3__40_;
  assign t_4__31_ = t_3__31_ & t_3__39_;
  assign t_4__30_ = t_3__30_ & t_3__38_;
  assign t_4__29_ = t_3__29_ & t_3__37_;
  assign t_4__28_ = t_3__28_ & t_3__36_;
  assign t_4__27_ = t_3__27_ & t_3__35_;
  assign t_4__26_ = t_3__26_ & t_3__34_;
  assign t_4__25_ = t_3__25_ & t_3__33_;
  assign t_4__24_ = t_3__24_ & t_3__32_;
  assign t_4__23_ = t_3__23_ & t_3__31_;
  assign t_4__22_ = t_3__22_ & t_3__30_;
  assign t_4__21_ = t_3__21_ & t_3__29_;
  assign t_4__20_ = t_3__20_ & t_3__28_;
  assign t_4__19_ = t_3__19_ & t_3__27_;
  assign t_4__18_ = t_3__18_ & t_3__26_;
  assign t_4__17_ = t_3__17_ & t_3__25_;
  assign t_4__16_ = t_3__16_ & t_3__24_;
  assign t_4__15_ = t_3__15_ & t_3__23_;
  assign t_4__14_ = t_3__14_ & t_3__22_;
  assign t_4__13_ = t_3__13_ & t_3__21_;
  assign t_4__12_ = t_3__12_ & t_3__20_;
  assign t_4__11_ = t_3__11_ & t_3__19_;
  assign t_4__10_ = t_3__10_ & t_3__18_;
  assign t_4__9_ = t_3__9_ & t_3__17_;
  assign t_4__8_ = t_3__8_ & t_3__16_;
  assign t_4__7_ = t_3__7_ & t_3__15_;
  assign t_4__6_ = t_3__6_ & t_3__14_;
  assign t_4__5_ = t_3__5_ & t_3__13_;
  assign t_4__4_ = t_3__4_ & t_3__12_;
  assign t_4__3_ = t_3__3_ & t_3__11_;
  assign t_4__2_ = t_3__2_ & t_3__10_;
  assign t_4__1_ = t_3__1_ & t_3__9_;
  assign t_4__0_ = t_3__0_ & t_3__8_;
  assign t_5__127_ = t_4__127_ & 1'b1;
  assign t_5__126_ = t_4__126_ & 1'b1;
  assign t_5__125_ = t_4__125_ & 1'b1;
  assign t_5__124_ = t_4__124_ & 1'b1;
  assign t_5__123_ = t_4__123_ & 1'b1;
  assign t_5__122_ = t_4__122_ & 1'b1;
  assign t_5__121_ = t_4__121_ & 1'b1;
  assign t_5__120_ = t_4__120_ & 1'b1;
  assign t_5__119_ = t_4__119_ & 1'b1;
  assign t_5__118_ = t_4__118_ & 1'b1;
  assign t_5__117_ = t_4__117_ & 1'b1;
  assign t_5__116_ = t_4__116_ & 1'b1;
  assign t_5__115_ = t_4__115_ & 1'b1;
  assign t_5__114_ = t_4__114_ & 1'b1;
  assign t_5__113_ = t_4__113_ & 1'b1;
  assign t_5__112_ = t_4__112_ & 1'b1;
  assign t_5__111_ = t_4__111_ & t_4__127_;
  assign t_5__110_ = t_4__110_ & t_4__126_;
  assign t_5__109_ = t_4__109_ & t_4__125_;
  assign t_5__108_ = t_4__108_ & t_4__124_;
  assign t_5__107_ = t_4__107_ & t_4__123_;
  assign t_5__106_ = t_4__106_ & t_4__122_;
  assign t_5__105_ = t_4__105_ & t_4__121_;
  assign t_5__104_ = t_4__104_ & t_4__120_;
  assign t_5__103_ = t_4__103_ & t_4__119_;
  assign t_5__102_ = t_4__102_ & t_4__118_;
  assign t_5__101_ = t_4__101_ & t_4__117_;
  assign t_5__100_ = t_4__100_ & t_4__116_;
  assign t_5__99_ = t_4__99_ & t_4__115_;
  assign t_5__98_ = t_4__98_ & t_4__114_;
  assign t_5__97_ = t_4__97_ & t_4__113_;
  assign t_5__96_ = t_4__96_ & t_4__112_;
  assign t_5__95_ = t_4__95_ & t_4__111_;
  assign t_5__94_ = t_4__94_ & t_4__110_;
  assign t_5__93_ = t_4__93_ & t_4__109_;
  assign t_5__92_ = t_4__92_ & t_4__108_;
  assign t_5__91_ = t_4__91_ & t_4__107_;
  assign t_5__90_ = t_4__90_ & t_4__106_;
  assign t_5__89_ = t_4__89_ & t_4__105_;
  assign t_5__88_ = t_4__88_ & t_4__104_;
  assign t_5__87_ = t_4__87_ & t_4__103_;
  assign t_5__86_ = t_4__86_ & t_4__102_;
  assign t_5__85_ = t_4__85_ & t_4__101_;
  assign t_5__84_ = t_4__84_ & t_4__100_;
  assign t_5__83_ = t_4__83_ & t_4__99_;
  assign t_5__82_ = t_4__82_ & t_4__98_;
  assign t_5__81_ = t_4__81_ & t_4__97_;
  assign t_5__80_ = t_4__80_ & t_4__96_;
  assign t_5__79_ = t_4__79_ & t_4__95_;
  assign t_5__78_ = t_4__78_ & t_4__94_;
  assign t_5__77_ = t_4__77_ & t_4__93_;
  assign t_5__76_ = t_4__76_ & t_4__92_;
  assign t_5__75_ = t_4__75_ & t_4__91_;
  assign t_5__74_ = t_4__74_ & t_4__90_;
  assign t_5__73_ = t_4__73_ & t_4__89_;
  assign t_5__72_ = t_4__72_ & t_4__88_;
  assign t_5__71_ = t_4__71_ & t_4__87_;
  assign t_5__70_ = t_4__70_ & t_4__86_;
  assign t_5__69_ = t_4__69_ & t_4__85_;
  assign t_5__68_ = t_4__68_ & t_4__84_;
  assign t_5__67_ = t_4__67_ & t_4__83_;
  assign t_5__66_ = t_4__66_ & t_4__82_;
  assign t_5__65_ = t_4__65_ & t_4__81_;
  assign t_5__64_ = t_4__64_ & t_4__80_;
  assign t_5__63_ = t_4__63_ & t_4__79_;
  assign t_5__62_ = t_4__62_ & t_4__78_;
  assign t_5__61_ = t_4__61_ & t_4__77_;
  assign t_5__60_ = t_4__60_ & t_4__76_;
  assign t_5__59_ = t_4__59_ & t_4__75_;
  assign t_5__58_ = t_4__58_ & t_4__74_;
  assign t_5__57_ = t_4__57_ & t_4__73_;
  assign t_5__56_ = t_4__56_ & t_4__72_;
  assign t_5__55_ = t_4__55_ & t_4__71_;
  assign t_5__54_ = t_4__54_ & t_4__70_;
  assign t_5__53_ = t_4__53_ & t_4__69_;
  assign t_5__52_ = t_4__52_ & t_4__68_;
  assign t_5__51_ = t_4__51_ & t_4__67_;
  assign t_5__50_ = t_4__50_ & t_4__66_;
  assign t_5__49_ = t_4__49_ & t_4__65_;
  assign t_5__48_ = t_4__48_ & t_4__64_;
  assign t_5__47_ = t_4__47_ & t_4__63_;
  assign t_5__46_ = t_4__46_ & t_4__62_;
  assign t_5__45_ = t_4__45_ & t_4__61_;
  assign t_5__44_ = t_4__44_ & t_4__60_;
  assign t_5__43_ = t_4__43_ & t_4__59_;
  assign t_5__42_ = t_4__42_ & t_4__58_;
  assign t_5__41_ = t_4__41_ & t_4__57_;
  assign t_5__40_ = t_4__40_ & t_4__56_;
  assign t_5__39_ = t_4__39_ & t_4__55_;
  assign t_5__38_ = t_4__38_ & t_4__54_;
  assign t_5__37_ = t_4__37_ & t_4__53_;
  assign t_5__36_ = t_4__36_ & t_4__52_;
  assign t_5__35_ = t_4__35_ & t_4__51_;
  assign t_5__34_ = t_4__34_ & t_4__50_;
  assign t_5__33_ = t_4__33_ & t_4__49_;
  assign t_5__32_ = t_4__32_ & t_4__48_;
  assign t_5__31_ = t_4__31_ & t_4__47_;
  assign t_5__30_ = t_4__30_ & t_4__46_;
  assign t_5__29_ = t_4__29_ & t_4__45_;
  assign t_5__28_ = t_4__28_ & t_4__44_;
  assign t_5__27_ = t_4__27_ & t_4__43_;
  assign t_5__26_ = t_4__26_ & t_4__42_;
  assign t_5__25_ = t_4__25_ & t_4__41_;
  assign t_5__24_ = t_4__24_ & t_4__40_;
  assign t_5__23_ = t_4__23_ & t_4__39_;
  assign t_5__22_ = t_4__22_ & t_4__38_;
  assign t_5__21_ = t_4__21_ & t_4__37_;
  assign t_5__20_ = t_4__20_ & t_4__36_;
  assign t_5__19_ = t_4__19_ & t_4__35_;
  assign t_5__18_ = t_4__18_ & t_4__34_;
  assign t_5__17_ = t_4__17_ & t_4__33_;
  assign t_5__16_ = t_4__16_ & t_4__32_;
  assign t_5__15_ = t_4__15_ & t_4__31_;
  assign t_5__14_ = t_4__14_ & t_4__30_;
  assign t_5__13_ = t_4__13_ & t_4__29_;
  assign t_5__12_ = t_4__12_ & t_4__28_;
  assign t_5__11_ = t_4__11_ & t_4__27_;
  assign t_5__10_ = t_4__10_ & t_4__26_;
  assign t_5__9_ = t_4__9_ & t_4__25_;
  assign t_5__8_ = t_4__8_ & t_4__24_;
  assign t_5__7_ = t_4__7_ & t_4__23_;
  assign t_5__6_ = t_4__6_ & t_4__22_;
  assign t_5__5_ = t_4__5_ & t_4__21_;
  assign t_5__4_ = t_4__4_ & t_4__20_;
  assign t_5__3_ = t_4__3_ & t_4__19_;
  assign t_5__2_ = t_4__2_ & t_4__18_;
  assign t_5__1_ = t_4__1_ & t_4__17_;
  assign t_5__0_ = t_4__0_ & t_4__16_;
  assign t_6__127_ = t_5__127_ & 1'b1;
  assign t_6__126_ = t_5__126_ & 1'b1;
  assign t_6__125_ = t_5__125_ & 1'b1;
  assign t_6__124_ = t_5__124_ & 1'b1;
  assign t_6__123_ = t_5__123_ & 1'b1;
  assign t_6__122_ = t_5__122_ & 1'b1;
  assign t_6__121_ = t_5__121_ & 1'b1;
  assign t_6__120_ = t_5__120_ & 1'b1;
  assign t_6__119_ = t_5__119_ & 1'b1;
  assign t_6__118_ = t_5__118_ & 1'b1;
  assign t_6__117_ = t_5__117_ & 1'b1;
  assign t_6__116_ = t_5__116_ & 1'b1;
  assign t_6__115_ = t_5__115_ & 1'b1;
  assign t_6__114_ = t_5__114_ & 1'b1;
  assign t_6__113_ = t_5__113_ & 1'b1;
  assign t_6__112_ = t_5__112_ & 1'b1;
  assign t_6__111_ = t_5__111_ & 1'b1;
  assign t_6__110_ = t_5__110_ & 1'b1;
  assign t_6__109_ = t_5__109_ & 1'b1;
  assign t_6__108_ = t_5__108_ & 1'b1;
  assign t_6__107_ = t_5__107_ & 1'b1;
  assign t_6__106_ = t_5__106_ & 1'b1;
  assign t_6__105_ = t_5__105_ & 1'b1;
  assign t_6__104_ = t_5__104_ & 1'b1;
  assign t_6__103_ = t_5__103_ & 1'b1;
  assign t_6__102_ = t_5__102_ & 1'b1;
  assign t_6__101_ = t_5__101_ & 1'b1;
  assign t_6__100_ = t_5__100_ & 1'b1;
  assign t_6__99_ = t_5__99_ & 1'b1;
  assign t_6__98_ = t_5__98_ & 1'b1;
  assign t_6__97_ = t_5__97_ & 1'b1;
  assign t_6__96_ = t_5__96_ & 1'b1;
  assign t_6__95_ = t_5__95_ & t_5__127_;
  assign t_6__94_ = t_5__94_ & t_5__126_;
  assign t_6__93_ = t_5__93_ & t_5__125_;
  assign t_6__92_ = t_5__92_ & t_5__124_;
  assign t_6__91_ = t_5__91_ & t_5__123_;
  assign t_6__90_ = t_5__90_ & t_5__122_;
  assign t_6__89_ = t_5__89_ & t_5__121_;
  assign t_6__88_ = t_5__88_ & t_5__120_;
  assign t_6__87_ = t_5__87_ & t_5__119_;
  assign t_6__86_ = t_5__86_ & t_5__118_;
  assign t_6__85_ = t_5__85_ & t_5__117_;
  assign t_6__84_ = t_5__84_ & t_5__116_;
  assign t_6__83_ = t_5__83_ & t_5__115_;
  assign t_6__82_ = t_5__82_ & t_5__114_;
  assign t_6__81_ = t_5__81_ & t_5__113_;
  assign t_6__80_ = t_5__80_ & t_5__112_;
  assign t_6__79_ = t_5__79_ & t_5__111_;
  assign t_6__78_ = t_5__78_ & t_5__110_;
  assign t_6__77_ = t_5__77_ & t_5__109_;
  assign t_6__76_ = t_5__76_ & t_5__108_;
  assign t_6__75_ = t_5__75_ & t_5__107_;
  assign t_6__74_ = t_5__74_ & t_5__106_;
  assign t_6__73_ = t_5__73_ & t_5__105_;
  assign t_6__72_ = t_5__72_ & t_5__104_;
  assign t_6__71_ = t_5__71_ & t_5__103_;
  assign t_6__70_ = t_5__70_ & t_5__102_;
  assign t_6__69_ = t_5__69_ & t_5__101_;
  assign t_6__68_ = t_5__68_ & t_5__100_;
  assign t_6__67_ = t_5__67_ & t_5__99_;
  assign t_6__66_ = t_5__66_ & t_5__98_;
  assign t_6__65_ = t_5__65_ & t_5__97_;
  assign t_6__64_ = t_5__64_ & t_5__96_;
  assign t_6__63_ = t_5__63_ & t_5__95_;
  assign t_6__62_ = t_5__62_ & t_5__94_;
  assign t_6__61_ = t_5__61_ & t_5__93_;
  assign t_6__60_ = t_5__60_ & t_5__92_;
  assign t_6__59_ = t_5__59_ & t_5__91_;
  assign t_6__58_ = t_5__58_ & t_5__90_;
  assign t_6__57_ = t_5__57_ & t_5__89_;
  assign t_6__56_ = t_5__56_ & t_5__88_;
  assign t_6__55_ = t_5__55_ & t_5__87_;
  assign t_6__54_ = t_5__54_ & t_5__86_;
  assign t_6__53_ = t_5__53_ & t_5__85_;
  assign t_6__52_ = t_5__52_ & t_5__84_;
  assign t_6__51_ = t_5__51_ & t_5__83_;
  assign t_6__50_ = t_5__50_ & t_5__82_;
  assign t_6__49_ = t_5__49_ & t_5__81_;
  assign t_6__48_ = t_5__48_ & t_5__80_;
  assign t_6__47_ = t_5__47_ & t_5__79_;
  assign t_6__46_ = t_5__46_ & t_5__78_;
  assign t_6__45_ = t_5__45_ & t_5__77_;
  assign t_6__44_ = t_5__44_ & t_5__76_;
  assign t_6__43_ = t_5__43_ & t_5__75_;
  assign t_6__42_ = t_5__42_ & t_5__74_;
  assign t_6__41_ = t_5__41_ & t_5__73_;
  assign t_6__40_ = t_5__40_ & t_5__72_;
  assign t_6__39_ = t_5__39_ & t_5__71_;
  assign t_6__38_ = t_5__38_ & t_5__70_;
  assign t_6__37_ = t_5__37_ & t_5__69_;
  assign t_6__36_ = t_5__36_ & t_5__68_;
  assign t_6__35_ = t_5__35_ & t_5__67_;
  assign t_6__34_ = t_5__34_ & t_5__66_;
  assign t_6__33_ = t_5__33_ & t_5__65_;
  assign t_6__32_ = t_5__32_ & t_5__64_;
  assign t_6__31_ = t_5__31_ & t_5__63_;
  assign t_6__30_ = t_5__30_ & t_5__62_;
  assign t_6__29_ = t_5__29_ & t_5__61_;
  assign t_6__28_ = t_5__28_ & t_5__60_;
  assign t_6__27_ = t_5__27_ & t_5__59_;
  assign t_6__26_ = t_5__26_ & t_5__58_;
  assign t_6__25_ = t_5__25_ & t_5__57_;
  assign t_6__24_ = t_5__24_ & t_5__56_;
  assign t_6__23_ = t_5__23_ & t_5__55_;
  assign t_6__22_ = t_5__22_ & t_5__54_;
  assign t_6__21_ = t_5__21_ & t_5__53_;
  assign t_6__20_ = t_5__20_ & t_5__52_;
  assign t_6__19_ = t_5__19_ & t_5__51_;
  assign t_6__18_ = t_5__18_ & t_5__50_;
  assign t_6__17_ = t_5__17_ & t_5__49_;
  assign t_6__16_ = t_5__16_ & t_5__48_;
  assign t_6__15_ = t_5__15_ & t_5__47_;
  assign t_6__14_ = t_5__14_ & t_5__46_;
  assign t_6__13_ = t_5__13_ & t_5__45_;
  assign t_6__12_ = t_5__12_ & t_5__44_;
  assign t_6__11_ = t_5__11_ & t_5__43_;
  assign t_6__10_ = t_5__10_ & t_5__42_;
  assign t_6__9_ = t_5__9_ & t_5__41_;
  assign t_6__8_ = t_5__8_ & t_5__40_;
  assign t_6__7_ = t_5__7_ & t_5__39_;
  assign t_6__6_ = t_5__6_ & t_5__38_;
  assign t_6__5_ = t_5__5_ & t_5__37_;
  assign t_6__4_ = t_5__4_ & t_5__36_;
  assign t_6__3_ = t_5__3_ & t_5__35_;
  assign t_6__2_ = t_5__2_ & t_5__34_;
  assign t_6__1_ = t_5__1_ & t_5__33_;
  assign t_6__0_ = t_5__0_ & t_5__32_;
  assign o[0] = t_6__127_ & 1'b1;
  assign o[1] = t_6__126_ & 1'b1;
  assign o[2] = t_6__125_ & 1'b1;
  assign o[3] = t_6__124_ & 1'b1;
  assign o[4] = t_6__123_ & 1'b1;
  assign o[5] = t_6__122_ & 1'b1;
  assign o[6] = t_6__121_ & 1'b1;
  assign o[7] = t_6__120_ & 1'b1;
  assign o[8] = t_6__119_ & 1'b1;
  assign o[9] = t_6__118_ & 1'b1;
  assign o[10] = t_6__117_ & 1'b1;
  assign o[11] = t_6__116_ & 1'b1;
  assign o[12] = t_6__115_ & 1'b1;
  assign o[13] = t_6__114_ & 1'b1;
  assign o[14] = t_6__113_ & 1'b1;
  assign o[15] = t_6__112_ & 1'b1;
  assign o[16] = t_6__111_ & 1'b1;
  assign o[17] = t_6__110_ & 1'b1;
  assign o[18] = t_6__109_ & 1'b1;
  assign o[19] = t_6__108_ & 1'b1;
  assign o[20] = t_6__107_ & 1'b1;
  assign o[21] = t_6__106_ & 1'b1;
  assign o[22] = t_6__105_ & 1'b1;
  assign o[23] = t_6__104_ & 1'b1;
  assign o[24] = t_6__103_ & 1'b1;
  assign o[25] = t_6__102_ & 1'b1;
  assign o[26] = t_6__101_ & 1'b1;
  assign o[27] = t_6__100_ & 1'b1;
  assign o[28] = t_6__99_ & 1'b1;
  assign o[29] = t_6__98_ & 1'b1;
  assign o[30] = t_6__97_ & 1'b1;
  assign o[31] = t_6__96_ & 1'b1;
  assign o[32] = t_6__95_ & 1'b1;
  assign o[33] = t_6__94_ & 1'b1;
  assign o[34] = t_6__93_ & 1'b1;
  assign o[35] = t_6__92_ & 1'b1;
  assign o[36] = t_6__91_ & 1'b1;
  assign o[37] = t_6__90_ & 1'b1;
  assign o[38] = t_6__89_ & 1'b1;
  assign o[39] = t_6__88_ & 1'b1;
  assign o[40] = t_6__87_ & 1'b1;
  assign o[41] = t_6__86_ & 1'b1;
  assign o[42] = t_6__85_ & 1'b1;
  assign o[43] = t_6__84_ & 1'b1;
  assign o[44] = t_6__83_ & 1'b1;
  assign o[45] = t_6__82_ & 1'b1;
  assign o[46] = t_6__81_ & 1'b1;
  assign o[47] = t_6__80_ & 1'b1;
  assign o[48] = t_6__79_ & 1'b1;
  assign o[49] = t_6__78_ & 1'b1;
  assign o[50] = t_6__77_ & 1'b1;
  assign o[51] = t_6__76_ & 1'b1;
  assign o[52] = t_6__75_ & 1'b1;
  assign o[53] = t_6__74_ & 1'b1;
  assign o[54] = t_6__73_ & 1'b1;
  assign o[55] = t_6__72_ & 1'b1;
  assign o[56] = t_6__71_ & 1'b1;
  assign o[57] = t_6__70_ & 1'b1;
  assign o[58] = t_6__69_ & 1'b1;
  assign o[59] = t_6__68_ & 1'b1;
  assign o[60] = t_6__67_ & 1'b1;
  assign o[61] = t_6__66_ & 1'b1;
  assign o[62] = t_6__65_ & 1'b1;
  assign o[63] = t_6__64_ & 1'b1;
  assign o[64] = t_6__63_ & t_6__127_;
  assign o[65] = t_6__62_ & t_6__126_;
  assign o[66] = t_6__61_ & t_6__125_;
  assign o[67] = t_6__60_ & t_6__124_;
  assign o[68] = t_6__59_ & t_6__123_;
  assign o[69] = t_6__58_ & t_6__122_;
  assign o[70] = t_6__57_ & t_6__121_;
  assign o[71] = t_6__56_ & t_6__120_;
  assign o[72] = t_6__55_ & t_6__119_;
  assign o[73] = t_6__54_ & t_6__118_;
  assign o[74] = t_6__53_ & t_6__117_;
  assign o[75] = t_6__52_ & t_6__116_;
  assign o[76] = t_6__51_ & t_6__115_;
  assign o[77] = t_6__50_ & t_6__114_;
  assign o[78] = t_6__49_ & t_6__113_;
  assign o[79] = t_6__48_ & t_6__112_;
  assign o[80] = t_6__47_ & t_6__111_;
  assign o[81] = t_6__46_ & t_6__110_;
  assign o[82] = t_6__45_ & t_6__109_;
  assign o[83] = t_6__44_ & t_6__108_;
  assign o[84] = t_6__43_ & t_6__107_;
  assign o[85] = t_6__42_ & t_6__106_;
  assign o[86] = t_6__41_ & t_6__105_;
  assign o[87] = t_6__40_ & t_6__104_;
  assign o[88] = t_6__39_ & t_6__103_;
  assign o[89] = t_6__38_ & t_6__102_;
  assign o[90] = t_6__37_ & t_6__101_;
  assign o[91] = t_6__36_ & t_6__100_;
  assign o[92] = t_6__35_ & t_6__99_;
  assign o[93] = t_6__34_ & t_6__98_;
  assign o[94] = t_6__33_ & t_6__97_;
  assign o[95] = t_6__32_ & t_6__96_;
  assign o[96] = t_6__31_ & t_6__95_;
  assign o[97] = t_6__30_ & t_6__94_;
  assign o[98] = t_6__29_ & t_6__93_;
  assign o[99] = t_6__28_ & t_6__92_;
  assign o[100] = t_6__27_ & t_6__91_;
  assign o[101] = t_6__26_ & t_6__90_;
  assign o[102] = t_6__25_ & t_6__89_;
  assign o[103] = t_6__24_ & t_6__88_;
  assign o[104] = t_6__23_ & t_6__87_;
  assign o[105] = t_6__22_ & t_6__86_;
  assign o[106] = t_6__21_ & t_6__85_;
  assign o[107] = t_6__20_ & t_6__84_;
  assign o[108] = t_6__19_ & t_6__83_;
  assign o[109] = t_6__18_ & t_6__82_;
  assign o[110] = t_6__17_ & t_6__81_;
  assign o[111] = t_6__16_ & t_6__80_;
  assign o[112] = t_6__15_ & t_6__79_;
  assign o[113] = t_6__14_ & t_6__78_;
  assign o[114] = t_6__13_ & t_6__77_;
  assign o[115] = t_6__12_ & t_6__76_;
  assign o[116] = t_6__11_ & t_6__75_;
  assign o[117] = t_6__10_ & t_6__74_;
  assign o[118] = t_6__9_ & t_6__73_;
  assign o[119] = t_6__8_ & t_6__72_;
  assign o[120] = t_6__7_ & t_6__71_;
  assign o[121] = t_6__6_ & t_6__70_;
  assign o[122] = t_6__5_ & t_6__69_;
  assign o[123] = t_6__4_ & t_6__68_;
  assign o[124] = t_6__3_ & t_6__67_;
  assign o[125] = t_6__2_ & t_6__66_;
  assign o[126] = t_6__1_ & t_6__65_;
  assign o[127] = t_6__0_ & t_6__64_;

endmodule



module bsg_binary_plus_one_to_gray
(
  binary_i,
  gray_o
);

  input [127:0] binary_i;
  output [127:0] gray_o;
  wire [127:0] gray_o,binary_scan,edge_detect;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254;

  bsg_scan_width_p128_and_p1_lo_to_hi_p1
  scan_and
  (
    .i(binary_i),
    .o(binary_scan)
  );

  assign edge_detect[127] = N0 & binary_scan[126];
  assign N0 = ~1'b0;
  assign edge_detect[126] = N1 & binary_scan[125];
  assign N1 = ~binary_scan[126];
  assign edge_detect[125] = N2 & binary_scan[124];
  assign N2 = ~binary_scan[125];
  assign edge_detect[124] = N3 & binary_scan[123];
  assign N3 = ~binary_scan[124];
  assign edge_detect[123] = N4 & binary_scan[122];
  assign N4 = ~binary_scan[123];
  assign edge_detect[122] = N5 & binary_scan[121];
  assign N5 = ~binary_scan[122];
  assign edge_detect[121] = N6 & binary_scan[120];
  assign N6 = ~binary_scan[121];
  assign edge_detect[120] = N7 & binary_scan[119];
  assign N7 = ~binary_scan[120];
  assign edge_detect[119] = N8 & binary_scan[118];
  assign N8 = ~binary_scan[119];
  assign edge_detect[118] = N9 & binary_scan[117];
  assign N9 = ~binary_scan[118];
  assign edge_detect[117] = N10 & binary_scan[116];
  assign N10 = ~binary_scan[117];
  assign edge_detect[116] = N11 & binary_scan[115];
  assign N11 = ~binary_scan[116];
  assign edge_detect[115] = N12 & binary_scan[114];
  assign N12 = ~binary_scan[115];
  assign edge_detect[114] = N13 & binary_scan[113];
  assign N13 = ~binary_scan[114];
  assign edge_detect[113] = N14 & binary_scan[112];
  assign N14 = ~binary_scan[113];
  assign edge_detect[112] = N15 & binary_scan[111];
  assign N15 = ~binary_scan[112];
  assign edge_detect[111] = N16 & binary_scan[110];
  assign N16 = ~binary_scan[111];
  assign edge_detect[110] = N17 & binary_scan[109];
  assign N17 = ~binary_scan[110];
  assign edge_detect[109] = N18 & binary_scan[108];
  assign N18 = ~binary_scan[109];
  assign edge_detect[108] = N19 & binary_scan[107];
  assign N19 = ~binary_scan[108];
  assign edge_detect[107] = N20 & binary_scan[106];
  assign N20 = ~binary_scan[107];
  assign edge_detect[106] = N21 & binary_scan[105];
  assign N21 = ~binary_scan[106];
  assign edge_detect[105] = N22 & binary_scan[104];
  assign N22 = ~binary_scan[105];
  assign edge_detect[104] = N23 & binary_scan[103];
  assign N23 = ~binary_scan[104];
  assign edge_detect[103] = N24 & binary_scan[102];
  assign N24 = ~binary_scan[103];
  assign edge_detect[102] = N25 & binary_scan[101];
  assign N25 = ~binary_scan[102];
  assign edge_detect[101] = N26 & binary_scan[100];
  assign N26 = ~binary_scan[101];
  assign edge_detect[100] = N27 & binary_scan[99];
  assign N27 = ~binary_scan[100];
  assign edge_detect[99] = N28 & binary_scan[98];
  assign N28 = ~binary_scan[99];
  assign edge_detect[98] = N29 & binary_scan[97];
  assign N29 = ~binary_scan[98];
  assign edge_detect[97] = N30 & binary_scan[96];
  assign N30 = ~binary_scan[97];
  assign edge_detect[96] = N31 & binary_scan[95];
  assign N31 = ~binary_scan[96];
  assign edge_detect[95] = N32 & binary_scan[94];
  assign N32 = ~binary_scan[95];
  assign edge_detect[94] = N33 & binary_scan[93];
  assign N33 = ~binary_scan[94];
  assign edge_detect[93] = N34 & binary_scan[92];
  assign N34 = ~binary_scan[93];
  assign edge_detect[92] = N35 & binary_scan[91];
  assign N35 = ~binary_scan[92];
  assign edge_detect[91] = N36 & binary_scan[90];
  assign N36 = ~binary_scan[91];
  assign edge_detect[90] = N37 & binary_scan[89];
  assign N37 = ~binary_scan[90];
  assign edge_detect[89] = N38 & binary_scan[88];
  assign N38 = ~binary_scan[89];
  assign edge_detect[88] = N39 & binary_scan[87];
  assign N39 = ~binary_scan[88];
  assign edge_detect[87] = N40 & binary_scan[86];
  assign N40 = ~binary_scan[87];
  assign edge_detect[86] = N41 & binary_scan[85];
  assign N41 = ~binary_scan[86];
  assign edge_detect[85] = N42 & binary_scan[84];
  assign N42 = ~binary_scan[85];
  assign edge_detect[84] = N43 & binary_scan[83];
  assign N43 = ~binary_scan[84];
  assign edge_detect[83] = N44 & binary_scan[82];
  assign N44 = ~binary_scan[83];
  assign edge_detect[82] = N45 & binary_scan[81];
  assign N45 = ~binary_scan[82];
  assign edge_detect[81] = N46 & binary_scan[80];
  assign N46 = ~binary_scan[81];
  assign edge_detect[80] = N47 & binary_scan[79];
  assign N47 = ~binary_scan[80];
  assign edge_detect[79] = N48 & binary_scan[78];
  assign N48 = ~binary_scan[79];
  assign edge_detect[78] = N49 & binary_scan[77];
  assign N49 = ~binary_scan[78];
  assign edge_detect[77] = N50 & binary_scan[76];
  assign N50 = ~binary_scan[77];
  assign edge_detect[76] = N51 & binary_scan[75];
  assign N51 = ~binary_scan[76];
  assign edge_detect[75] = N52 & binary_scan[74];
  assign N52 = ~binary_scan[75];
  assign edge_detect[74] = N53 & binary_scan[73];
  assign N53 = ~binary_scan[74];
  assign edge_detect[73] = N54 & binary_scan[72];
  assign N54 = ~binary_scan[73];
  assign edge_detect[72] = N55 & binary_scan[71];
  assign N55 = ~binary_scan[72];
  assign edge_detect[71] = N56 & binary_scan[70];
  assign N56 = ~binary_scan[71];
  assign edge_detect[70] = N57 & binary_scan[69];
  assign N57 = ~binary_scan[70];
  assign edge_detect[69] = N58 & binary_scan[68];
  assign N58 = ~binary_scan[69];
  assign edge_detect[68] = N59 & binary_scan[67];
  assign N59 = ~binary_scan[68];
  assign edge_detect[67] = N60 & binary_scan[66];
  assign N60 = ~binary_scan[67];
  assign edge_detect[66] = N61 & binary_scan[65];
  assign N61 = ~binary_scan[66];
  assign edge_detect[65] = N62 & binary_scan[64];
  assign N62 = ~binary_scan[65];
  assign edge_detect[64] = N63 & binary_scan[63];
  assign N63 = ~binary_scan[64];
  assign edge_detect[63] = N64 & binary_scan[62];
  assign N64 = ~binary_scan[63];
  assign edge_detect[62] = N65 & binary_scan[61];
  assign N65 = ~binary_scan[62];
  assign edge_detect[61] = N66 & binary_scan[60];
  assign N66 = ~binary_scan[61];
  assign edge_detect[60] = N67 & binary_scan[59];
  assign N67 = ~binary_scan[60];
  assign edge_detect[59] = N68 & binary_scan[58];
  assign N68 = ~binary_scan[59];
  assign edge_detect[58] = N69 & binary_scan[57];
  assign N69 = ~binary_scan[58];
  assign edge_detect[57] = N70 & binary_scan[56];
  assign N70 = ~binary_scan[57];
  assign edge_detect[56] = N71 & binary_scan[55];
  assign N71 = ~binary_scan[56];
  assign edge_detect[55] = N72 & binary_scan[54];
  assign N72 = ~binary_scan[55];
  assign edge_detect[54] = N73 & binary_scan[53];
  assign N73 = ~binary_scan[54];
  assign edge_detect[53] = N74 & binary_scan[52];
  assign N74 = ~binary_scan[53];
  assign edge_detect[52] = N75 & binary_scan[51];
  assign N75 = ~binary_scan[52];
  assign edge_detect[51] = N76 & binary_scan[50];
  assign N76 = ~binary_scan[51];
  assign edge_detect[50] = N77 & binary_scan[49];
  assign N77 = ~binary_scan[50];
  assign edge_detect[49] = N78 & binary_scan[48];
  assign N78 = ~binary_scan[49];
  assign edge_detect[48] = N79 & binary_scan[47];
  assign N79 = ~binary_scan[48];
  assign edge_detect[47] = N80 & binary_scan[46];
  assign N80 = ~binary_scan[47];
  assign edge_detect[46] = N81 & binary_scan[45];
  assign N81 = ~binary_scan[46];
  assign edge_detect[45] = N82 & binary_scan[44];
  assign N82 = ~binary_scan[45];
  assign edge_detect[44] = N83 & binary_scan[43];
  assign N83 = ~binary_scan[44];
  assign edge_detect[43] = N84 & binary_scan[42];
  assign N84 = ~binary_scan[43];
  assign edge_detect[42] = N85 & binary_scan[41];
  assign N85 = ~binary_scan[42];
  assign edge_detect[41] = N86 & binary_scan[40];
  assign N86 = ~binary_scan[41];
  assign edge_detect[40] = N87 & binary_scan[39];
  assign N87 = ~binary_scan[40];
  assign edge_detect[39] = N88 & binary_scan[38];
  assign N88 = ~binary_scan[39];
  assign edge_detect[38] = N89 & binary_scan[37];
  assign N89 = ~binary_scan[38];
  assign edge_detect[37] = N90 & binary_scan[36];
  assign N90 = ~binary_scan[37];
  assign edge_detect[36] = N91 & binary_scan[35];
  assign N91 = ~binary_scan[36];
  assign edge_detect[35] = N92 & binary_scan[34];
  assign N92 = ~binary_scan[35];
  assign edge_detect[34] = N93 & binary_scan[33];
  assign N93 = ~binary_scan[34];
  assign edge_detect[33] = N94 & binary_scan[32];
  assign N94 = ~binary_scan[33];
  assign edge_detect[32] = N95 & binary_scan[31];
  assign N95 = ~binary_scan[32];
  assign edge_detect[31] = N96 & binary_scan[30];
  assign N96 = ~binary_scan[31];
  assign edge_detect[30] = N97 & binary_scan[29];
  assign N97 = ~binary_scan[30];
  assign edge_detect[29] = N98 & binary_scan[28];
  assign N98 = ~binary_scan[29];
  assign edge_detect[28] = N99 & binary_scan[27];
  assign N99 = ~binary_scan[28];
  assign edge_detect[27] = N100 & binary_scan[26];
  assign N100 = ~binary_scan[27];
  assign edge_detect[26] = N101 & binary_scan[25];
  assign N101 = ~binary_scan[26];
  assign edge_detect[25] = N102 & binary_scan[24];
  assign N102 = ~binary_scan[25];
  assign edge_detect[24] = N103 & binary_scan[23];
  assign N103 = ~binary_scan[24];
  assign edge_detect[23] = N104 & binary_scan[22];
  assign N104 = ~binary_scan[23];
  assign edge_detect[22] = N105 & binary_scan[21];
  assign N105 = ~binary_scan[22];
  assign edge_detect[21] = N106 & binary_scan[20];
  assign N106 = ~binary_scan[21];
  assign edge_detect[20] = N107 & binary_scan[19];
  assign N107 = ~binary_scan[20];
  assign edge_detect[19] = N108 & binary_scan[18];
  assign N108 = ~binary_scan[19];
  assign edge_detect[18] = N109 & binary_scan[17];
  assign N109 = ~binary_scan[18];
  assign edge_detect[17] = N110 & binary_scan[16];
  assign N110 = ~binary_scan[17];
  assign edge_detect[16] = N111 & binary_scan[15];
  assign N111 = ~binary_scan[16];
  assign edge_detect[15] = N112 & binary_scan[14];
  assign N112 = ~binary_scan[15];
  assign edge_detect[14] = N113 & binary_scan[13];
  assign N113 = ~binary_scan[14];
  assign edge_detect[13] = N114 & binary_scan[12];
  assign N114 = ~binary_scan[13];
  assign edge_detect[12] = N115 & binary_scan[11];
  assign N115 = ~binary_scan[12];
  assign edge_detect[11] = N116 & binary_scan[10];
  assign N116 = ~binary_scan[11];
  assign edge_detect[10] = N117 & binary_scan[9];
  assign N117 = ~binary_scan[10];
  assign edge_detect[9] = N118 & binary_scan[8];
  assign N118 = ~binary_scan[9];
  assign edge_detect[8] = N119 & binary_scan[7];
  assign N119 = ~binary_scan[8];
  assign edge_detect[7] = N120 & binary_scan[6];
  assign N120 = ~binary_scan[7];
  assign edge_detect[6] = N121 & binary_scan[5];
  assign N121 = ~binary_scan[6];
  assign edge_detect[5] = N122 & binary_scan[4];
  assign N122 = ~binary_scan[5];
  assign edge_detect[4] = N123 & binary_scan[3];
  assign N123 = ~binary_scan[4];
  assign edge_detect[3] = N124 & binary_scan[2];
  assign N124 = ~binary_scan[3];
  assign edge_detect[2] = N125 & binary_scan[1];
  assign N125 = ~binary_scan[2];
  assign edge_detect[1] = N126 & binary_scan[0];
  assign N126 = ~binary_scan[1];
  assign edge_detect[0] = N127 & 1'b1;
  assign N127 = ~binary_scan[0];
  assign gray_o[127] = binary_i[127] ^ edge_detect[127];
  assign gray_o[126] = N128 ^ edge_detect[126];
  assign N128 = binary_i[127] ^ binary_i[126];
  assign gray_o[125] = N129 ^ edge_detect[125];
  assign N129 = binary_i[126] ^ binary_i[125];
  assign gray_o[124] = N130 ^ edge_detect[124];
  assign N130 = binary_i[125] ^ binary_i[124];
  assign gray_o[123] = N131 ^ edge_detect[123];
  assign N131 = binary_i[124] ^ binary_i[123];
  assign gray_o[122] = N132 ^ edge_detect[122];
  assign N132 = binary_i[123] ^ binary_i[122];
  assign gray_o[121] = N133 ^ edge_detect[121];
  assign N133 = binary_i[122] ^ binary_i[121];
  assign gray_o[120] = N134 ^ edge_detect[120];
  assign N134 = binary_i[121] ^ binary_i[120];
  assign gray_o[119] = N135 ^ edge_detect[119];
  assign N135 = binary_i[120] ^ binary_i[119];
  assign gray_o[118] = N136 ^ edge_detect[118];
  assign N136 = binary_i[119] ^ binary_i[118];
  assign gray_o[117] = N137 ^ edge_detect[117];
  assign N137 = binary_i[118] ^ binary_i[117];
  assign gray_o[116] = N138 ^ edge_detect[116];
  assign N138 = binary_i[117] ^ binary_i[116];
  assign gray_o[115] = N139 ^ edge_detect[115];
  assign N139 = binary_i[116] ^ binary_i[115];
  assign gray_o[114] = N140 ^ edge_detect[114];
  assign N140 = binary_i[115] ^ binary_i[114];
  assign gray_o[113] = N141 ^ edge_detect[113];
  assign N141 = binary_i[114] ^ binary_i[113];
  assign gray_o[112] = N142 ^ edge_detect[112];
  assign N142 = binary_i[113] ^ binary_i[112];
  assign gray_o[111] = N143 ^ edge_detect[111];
  assign N143 = binary_i[112] ^ binary_i[111];
  assign gray_o[110] = N144 ^ edge_detect[110];
  assign N144 = binary_i[111] ^ binary_i[110];
  assign gray_o[109] = N145 ^ edge_detect[109];
  assign N145 = binary_i[110] ^ binary_i[109];
  assign gray_o[108] = N146 ^ edge_detect[108];
  assign N146 = binary_i[109] ^ binary_i[108];
  assign gray_o[107] = N147 ^ edge_detect[107];
  assign N147 = binary_i[108] ^ binary_i[107];
  assign gray_o[106] = N148 ^ edge_detect[106];
  assign N148 = binary_i[107] ^ binary_i[106];
  assign gray_o[105] = N149 ^ edge_detect[105];
  assign N149 = binary_i[106] ^ binary_i[105];
  assign gray_o[104] = N150 ^ edge_detect[104];
  assign N150 = binary_i[105] ^ binary_i[104];
  assign gray_o[103] = N151 ^ edge_detect[103];
  assign N151 = binary_i[104] ^ binary_i[103];
  assign gray_o[102] = N152 ^ edge_detect[102];
  assign N152 = binary_i[103] ^ binary_i[102];
  assign gray_o[101] = N153 ^ edge_detect[101];
  assign N153 = binary_i[102] ^ binary_i[101];
  assign gray_o[100] = N154 ^ edge_detect[100];
  assign N154 = binary_i[101] ^ binary_i[100];
  assign gray_o[99] = N155 ^ edge_detect[99];
  assign N155 = binary_i[100] ^ binary_i[99];
  assign gray_o[98] = N156 ^ edge_detect[98];
  assign N156 = binary_i[99] ^ binary_i[98];
  assign gray_o[97] = N157 ^ edge_detect[97];
  assign N157 = binary_i[98] ^ binary_i[97];
  assign gray_o[96] = N158 ^ edge_detect[96];
  assign N158 = binary_i[97] ^ binary_i[96];
  assign gray_o[95] = N159 ^ edge_detect[95];
  assign N159 = binary_i[96] ^ binary_i[95];
  assign gray_o[94] = N160 ^ edge_detect[94];
  assign N160 = binary_i[95] ^ binary_i[94];
  assign gray_o[93] = N161 ^ edge_detect[93];
  assign N161 = binary_i[94] ^ binary_i[93];
  assign gray_o[92] = N162 ^ edge_detect[92];
  assign N162 = binary_i[93] ^ binary_i[92];
  assign gray_o[91] = N163 ^ edge_detect[91];
  assign N163 = binary_i[92] ^ binary_i[91];
  assign gray_o[90] = N164 ^ edge_detect[90];
  assign N164 = binary_i[91] ^ binary_i[90];
  assign gray_o[89] = N165 ^ edge_detect[89];
  assign N165 = binary_i[90] ^ binary_i[89];
  assign gray_o[88] = N166 ^ edge_detect[88];
  assign N166 = binary_i[89] ^ binary_i[88];
  assign gray_o[87] = N167 ^ edge_detect[87];
  assign N167 = binary_i[88] ^ binary_i[87];
  assign gray_o[86] = N168 ^ edge_detect[86];
  assign N168 = binary_i[87] ^ binary_i[86];
  assign gray_o[85] = N169 ^ edge_detect[85];
  assign N169 = binary_i[86] ^ binary_i[85];
  assign gray_o[84] = N170 ^ edge_detect[84];
  assign N170 = binary_i[85] ^ binary_i[84];
  assign gray_o[83] = N171 ^ edge_detect[83];
  assign N171 = binary_i[84] ^ binary_i[83];
  assign gray_o[82] = N172 ^ edge_detect[82];
  assign N172 = binary_i[83] ^ binary_i[82];
  assign gray_o[81] = N173 ^ edge_detect[81];
  assign N173 = binary_i[82] ^ binary_i[81];
  assign gray_o[80] = N174 ^ edge_detect[80];
  assign N174 = binary_i[81] ^ binary_i[80];
  assign gray_o[79] = N175 ^ edge_detect[79];
  assign N175 = binary_i[80] ^ binary_i[79];
  assign gray_o[78] = N176 ^ edge_detect[78];
  assign N176 = binary_i[79] ^ binary_i[78];
  assign gray_o[77] = N177 ^ edge_detect[77];
  assign N177 = binary_i[78] ^ binary_i[77];
  assign gray_o[76] = N178 ^ edge_detect[76];
  assign N178 = binary_i[77] ^ binary_i[76];
  assign gray_o[75] = N179 ^ edge_detect[75];
  assign N179 = binary_i[76] ^ binary_i[75];
  assign gray_o[74] = N180 ^ edge_detect[74];
  assign N180 = binary_i[75] ^ binary_i[74];
  assign gray_o[73] = N181 ^ edge_detect[73];
  assign N181 = binary_i[74] ^ binary_i[73];
  assign gray_o[72] = N182 ^ edge_detect[72];
  assign N182 = binary_i[73] ^ binary_i[72];
  assign gray_o[71] = N183 ^ edge_detect[71];
  assign N183 = binary_i[72] ^ binary_i[71];
  assign gray_o[70] = N184 ^ edge_detect[70];
  assign N184 = binary_i[71] ^ binary_i[70];
  assign gray_o[69] = N185 ^ edge_detect[69];
  assign N185 = binary_i[70] ^ binary_i[69];
  assign gray_o[68] = N186 ^ edge_detect[68];
  assign N186 = binary_i[69] ^ binary_i[68];
  assign gray_o[67] = N187 ^ edge_detect[67];
  assign N187 = binary_i[68] ^ binary_i[67];
  assign gray_o[66] = N188 ^ edge_detect[66];
  assign N188 = binary_i[67] ^ binary_i[66];
  assign gray_o[65] = N189 ^ edge_detect[65];
  assign N189 = binary_i[66] ^ binary_i[65];
  assign gray_o[64] = N190 ^ edge_detect[64];
  assign N190 = binary_i[65] ^ binary_i[64];
  assign gray_o[63] = N191 ^ edge_detect[63];
  assign N191 = binary_i[64] ^ binary_i[63];
  assign gray_o[62] = N192 ^ edge_detect[62];
  assign N192 = binary_i[63] ^ binary_i[62];
  assign gray_o[61] = N193 ^ edge_detect[61];
  assign N193 = binary_i[62] ^ binary_i[61];
  assign gray_o[60] = N194 ^ edge_detect[60];
  assign N194 = binary_i[61] ^ binary_i[60];
  assign gray_o[59] = N195 ^ edge_detect[59];
  assign N195 = binary_i[60] ^ binary_i[59];
  assign gray_o[58] = N196 ^ edge_detect[58];
  assign N196 = binary_i[59] ^ binary_i[58];
  assign gray_o[57] = N197 ^ edge_detect[57];
  assign N197 = binary_i[58] ^ binary_i[57];
  assign gray_o[56] = N198 ^ edge_detect[56];
  assign N198 = binary_i[57] ^ binary_i[56];
  assign gray_o[55] = N199 ^ edge_detect[55];
  assign N199 = binary_i[56] ^ binary_i[55];
  assign gray_o[54] = N200 ^ edge_detect[54];
  assign N200 = binary_i[55] ^ binary_i[54];
  assign gray_o[53] = N201 ^ edge_detect[53];
  assign N201 = binary_i[54] ^ binary_i[53];
  assign gray_o[52] = N202 ^ edge_detect[52];
  assign N202 = binary_i[53] ^ binary_i[52];
  assign gray_o[51] = N203 ^ edge_detect[51];
  assign N203 = binary_i[52] ^ binary_i[51];
  assign gray_o[50] = N204 ^ edge_detect[50];
  assign N204 = binary_i[51] ^ binary_i[50];
  assign gray_o[49] = N205 ^ edge_detect[49];
  assign N205 = binary_i[50] ^ binary_i[49];
  assign gray_o[48] = N206 ^ edge_detect[48];
  assign N206 = binary_i[49] ^ binary_i[48];
  assign gray_o[47] = N207 ^ edge_detect[47];
  assign N207 = binary_i[48] ^ binary_i[47];
  assign gray_o[46] = N208 ^ edge_detect[46];
  assign N208 = binary_i[47] ^ binary_i[46];
  assign gray_o[45] = N209 ^ edge_detect[45];
  assign N209 = binary_i[46] ^ binary_i[45];
  assign gray_o[44] = N210 ^ edge_detect[44];
  assign N210 = binary_i[45] ^ binary_i[44];
  assign gray_o[43] = N211 ^ edge_detect[43];
  assign N211 = binary_i[44] ^ binary_i[43];
  assign gray_o[42] = N212 ^ edge_detect[42];
  assign N212 = binary_i[43] ^ binary_i[42];
  assign gray_o[41] = N213 ^ edge_detect[41];
  assign N213 = binary_i[42] ^ binary_i[41];
  assign gray_o[40] = N214 ^ edge_detect[40];
  assign N214 = binary_i[41] ^ binary_i[40];
  assign gray_o[39] = N215 ^ edge_detect[39];
  assign N215 = binary_i[40] ^ binary_i[39];
  assign gray_o[38] = N216 ^ edge_detect[38];
  assign N216 = binary_i[39] ^ binary_i[38];
  assign gray_o[37] = N217 ^ edge_detect[37];
  assign N217 = binary_i[38] ^ binary_i[37];
  assign gray_o[36] = N218 ^ edge_detect[36];
  assign N218 = binary_i[37] ^ binary_i[36];
  assign gray_o[35] = N219 ^ edge_detect[35];
  assign N219 = binary_i[36] ^ binary_i[35];
  assign gray_o[34] = N220 ^ edge_detect[34];
  assign N220 = binary_i[35] ^ binary_i[34];
  assign gray_o[33] = N221 ^ edge_detect[33];
  assign N221 = binary_i[34] ^ binary_i[33];
  assign gray_o[32] = N222 ^ edge_detect[32];
  assign N222 = binary_i[33] ^ binary_i[32];
  assign gray_o[31] = N223 ^ edge_detect[31];
  assign N223 = binary_i[32] ^ binary_i[31];
  assign gray_o[30] = N224 ^ edge_detect[30];
  assign N224 = binary_i[31] ^ binary_i[30];
  assign gray_o[29] = N225 ^ edge_detect[29];
  assign N225 = binary_i[30] ^ binary_i[29];
  assign gray_o[28] = N226 ^ edge_detect[28];
  assign N226 = binary_i[29] ^ binary_i[28];
  assign gray_o[27] = N227 ^ edge_detect[27];
  assign N227 = binary_i[28] ^ binary_i[27];
  assign gray_o[26] = N228 ^ edge_detect[26];
  assign N228 = binary_i[27] ^ binary_i[26];
  assign gray_o[25] = N229 ^ edge_detect[25];
  assign N229 = binary_i[26] ^ binary_i[25];
  assign gray_o[24] = N230 ^ edge_detect[24];
  assign N230 = binary_i[25] ^ binary_i[24];
  assign gray_o[23] = N231 ^ edge_detect[23];
  assign N231 = binary_i[24] ^ binary_i[23];
  assign gray_o[22] = N232 ^ edge_detect[22];
  assign N232 = binary_i[23] ^ binary_i[22];
  assign gray_o[21] = N233 ^ edge_detect[21];
  assign N233 = binary_i[22] ^ binary_i[21];
  assign gray_o[20] = N234 ^ edge_detect[20];
  assign N234 = binary_i[21] ^ binary_i[20];
  assign gray_o[19] = N235 ^ edge_detect[19];
  assign N235 = binary_i[20] ^ binary_i[19];
  assign gray_o[18] = N236 ^ edge_detect[18];
  assign N236 = binary_i[19] ^ binary_i[18];
  assign gray_o[17] = N237 ^ edge_detect[17];
  assign N237 = binary_i[18] ^ binary_i[17];
  assign gray_o[16] = N238 ^ edge_detect[16];
  assign N238 = binary_i[17] ^ binary_i[16];
  assign gray_o[15] = N239 ^ edge_detect[15];
  assign N239 = binary_i[16] ^ binary_i[15];
  assign gray_o[14] = N240 ^ edge_detect[14];
  assign N240 = binary_i[15] ^ binary_i[14];
  assign gray_o[13] = N241 ^ edge_detect[13];
  assign N241 = binary_i[14] ^ binary_i[13];
  assign gray_o[12] = N242 ^ edge_detect[12];
  assign N242 = binary_i[13] ^ binary_i[12];
  assign gray_o[11] = N243 ^ edge_detect[11];
  assign N243 = binary_i[12] ^ binary_i[11];
  assign gray_o[10] = N244 ^ edge_detect[10];
  assign N244 = binary_i[11] ^ binary_i[10];
  assign gray_o[9] = N245 ^ edge_detect[9];
  assign N245 = binary_i[10] ^ binary_i[9];
  assign gray_o[8] = N246 ^ edge_detect[8];
  assign N246 = binary_i[9] ^ binary_i[8];
  assign gray_o[7] = N247 ^ edge_detect[7];
  assign N247 = binary_i[8] ^ binary_i[7];
  assign gray_o[6] = N248 ^ edge_detect[6];
  assign N248 = binary_i[7] ^ binary_i[6];
  assign gray_o[5] = N249 ^ edge_detect[5];
  assign N249 = binary_i[6] ^ binary_i[5];
  assign gray_o[4] = N250 ^ edge_detect[4];
  assign N250 = binary_i[5] ^ binary_i[4];
  assign gray_o[3] = N251 ^ edge_detect[3];
  assign N251 = binary_i[4] ^ binary_i[3];
  assign gray_o[2] = N252 ^ edge_detect[2];
  assign N252 = binary_i[3] ^ binary_i[2];
  assign gray_o[1] = N253 ^ edge_detect[1];
  assign N253 = binary_i[2] ^ binary_i[1];
  assign gray_o[0] = N254 ^ edge_detect[0];
  assign N254 = binary_i[1] ^ binary_i[0];

endmodule

