

module top
(
  lru_i,
  way_id_o
);

  input [30:0] lru_i;
  output [4:0] way_id_o;

  bsg_lru_pseudo_tree_encode
  wrapper
  (
    .lru_i(lru_i),
    .way_id_o(way_id_o)
  );


endmodule



module bsg_lru_pseudo_tree_encode
(
  lru_i,
  way_id_o
);

  input [30:0] lru_i;
  output [4:0] way_id_o;
  wire [4:0] way_id_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,pe_o_4__4_,pe_o_4__3_,pe_o_4__2_,pe_o_4__1_,pe_o_4__0_,pe_o_3__4_,
  pe_o_3__3_,pe_o_3__2_,pe_o_3__1_,pe_o_3__0_,pe_o_2__4_,pe_o_2__3_,pe_o_2__2_,
  pe_o_2__1_,pe_o_2__0_,pe_o_1__4_,pe_o_1__3_,pe_o_1__2_,pe_o_1__1_,pe_o_1__0_,N424,N425,
  N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,
  N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,
  N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,
  N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,pe_i_4__30_,pe_i_4__29_,
  pe_i_4__28_,pe_i_4__27_,pe_i_4__26_,pe_i_4__25_,pe_i_4__24_,pe_i_4__23_,pe_i_4__22_,
  pe_i_4__21_,pe_i_4__20_,pe_i_4__19_,pe_i_4__18_,pe_i_4__17_,pe_i_4__16_,
  pe_i_4__15_,pe_i_4__14_,pe_i_4__13_,pe_i_4__12_,pe_i_4__11_,pe_i_4__10_,pe_i_4__9_,
  pe_i_4__8_,pe_i_4__7_,pe_i_4__6_,pe_i_4__5_,pe_i_4__4_,pe_i_4__3_,pe_i_4__2_,
  pe_i_4__1_,pe_i_4__0_,pe_i_3__30_,pe_i_3__29_,pe_i_3__28_,pe_i_3__27_,pe_i_3__26_,
  pe_i_3__25_,pe_i_3__24_,pe_i_3__23_,pe_i_3__22_,pe_i_3__21_,pe_i_3__20_,pe_i_3__19_,
  pe_i_3__18_,pe_i_3__17_,pe_i_3__16_,pe_i_3__15_,pe_i_3__14_,pe_i_3__13_,pe_i_3__12_,
  pe_i_3__11_,pe_i_3__10_,pe_i_3__9_,pe_i_3__8_,pe_i_3__7_,pe_i_3__6_,pe_i_3__5_,
  pe_i_3__4_,pe_i_3__3_,pe_i_3__2_,pe_i_3__1_,pe_i_3__0_,pe_i_2__30_,pe_i_2__29_,
  pe_i_2__28_,pe_i_2__27_,pe_i_2__26_,pe_i_2__25_,pe_i_2__24_,pe_i_2__23_,
  pe_i_2__22_,pe_i_2__21_,pe_i_2__20_,pe_i_2__19_,pe_i_2__18_,pe_i_2__17_,pe_i_2__16_,
  pe_i_2__15_,pe_i_2__14_,pe_i_2__13_,pe_i_2__12_,pe_i_2__11_,pe_i_2__10_,pe_i_2__9_,
  pe_i_2__8_,pe_i_2__7_,pe_i_2__6_,pe_i_2__5_,pe_i_2__4_,pe_i_2__3_,pe_i_2__2_,
  pe_i_2__1_,pe_i_2__0_,pe_i_1__30_,pe_i_1__29_,pe_i_1__28_,pe_i_1__27_,pe_i_1__26_,
  pe_i_1__25_,pe_i_1__24_,pe_i_1__23_,pe_i_1__22_,pe_i_1__21_,pe_i_1__20_,pe_i_1__19_,
  pe_i_1__18_,pe_i_1__17_,pe_i_1__16_,pe_i_1__15_,pe_i_1__14_,pe_i_1__13_,
  pe_i_1__12_,pe_i_1__11_,pe_i_1__10_,pe_i_1__9_,pe_i_1__8_,pe_i_1__7_,pe_i_1__6_,
  pe_i_1__5_,pe_i_1__4_,pe_i_1__3_,pe_i_1__2_,pe_i_1__1_,pe_i_1__0_,N484,N485,N486,N487,
  N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,
  N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
  N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,
  N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,
  N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,
  N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
  N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,
  N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,
  N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,
  N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,
  N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,
  N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,
  N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,
  N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,
  N712,N713,N714,N715;
  wire [30:1] mask;

  bsg_priority_encode
  rof2_1__fi3_pe
  (
    .i({ pe_i_1__30_, pe_i_1__29_, pe_i_1__28_, pe_i_1__27_, pe_i_1__26_, pe_i_1__25_, pe_i_1__24_, pe_i_1__23_, pe_i_1__22_, pe_i_1__21_, pe_i_1__20_, pe_i_1__19_, pe_i_1__18_, pe_i_1__17_, pe_i_1__16_, pe_i_1__15_, pe_i_1__14_, pe_i_1__13_, pe_i_1__12_, pe_i_1__11_, pe_i_1__10_, pe_i_1__9_, pe_i_1__8_, pe_i_1__7_, pe_i_1__6_, pe_i_1__5_, pe_i_1__4_, pe_i_1__3_, pe_i_1__2_, pe_i_1__1_, pe_i_1__0_ }),
    .addr_o({ pe_o_1__4_, pe_o_1__3_, pe_o_1__2_, pe_o_1__1_, pe_o_1__0_ })
  );

  assign { N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_1__4_, pe_o_1__3_, pe_o_1__2_, pe_o_1__1_, pe_o_1__0_ };

  bsg_priority_encode
  rof2_2__fi3_pe
  (
    .i({ pe_i_2__30_, pe_i_2__29_, pe_i_2__28_, pe_i_2__27_, pe_i_2__26_, pe_i_2__25_, pe_i_2__24_, pe_i_2__23_, pe_i_2__22_, pe_i_2__21_, pe_i_2__20_, pe_i_2__19_, pe_i_2__18_, pe_i_2__17_, pe_i_2__16_, pe_i_2__15_, pe_i_2__14_, pe_i_2__13_, pe_i_2__12_, pe_i_2__11_, pe_i_2__10_, pe_i_2__9_, pe_i_2__8_, pe_i_2__7_, pe_i_2__6_, pe_i_2__5_, pe_i_2__4_, pe_i_2__3_, pe_i_2__2_, pe_i_2__1_, pe_i_2__0_ }),
    .addr_o({ pe_o_2__4_, pe_o_2__3_, pe_o_2__2_, pe_o_2__1_, pe_o_2__0_ })
  );

  assign { N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_2__4_, pe_o_2__3_, pe_o_2__2_, pe_o_2__1_, pe_o_2__0_ };

  bsg_priority_encode
  rof2_3__fi3_pe
  (
    .i({ pe_i_3__30_, pe_i_3__29_, pe_i_3__28_, pe_i_3__27_, pe_i_3__26_, pe_i_3__25_, pe_i_3__24_, pe_i_3__23_, pe_i_3__22_, pe_i_3__21_, pe_i_3__20_, pe_i_3__19_, pe_i_3__18_, pe_i_3__17_, pe_i_3__16_, pe_i_3__15_, pe_i_3__14_, pe_i_3__13_, pe_i_3__12_, pe_i_3__11_, pe_i_3__10_, pe_i_3__9_, pe_i_3__8_, pe_i_3__7_, pe_i_3__6_, pe_i_3__5_, pe_i_3__4_, pe_i_3__3_, pe_i_3__2_, pe_i_3__1_, pe_i_3__0_ }),
    .addr_o({ pe_o_3__4_, pe_o_3__3_, pe_o_3__2_, pe_o_3__1_, pe_o_3__0_ })
  );

  assign { N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670 } = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << { pe_o_3__4_, pe_o_3__3_, pe_o_3__2_, pe_o_3__1_, pe_o_3__0_ };

  bsg_priority_encode
  rof2_4__fi3_pe
  (
    .i({ pe_i_4__30_, pe_i_4__29_, pe_i_4__28_, pe_i_4__27_, pe_i_4__26_, pe_i_4__25_, pe_i_4__24_, pe_i_4__23_, pe_i_4__22_, pe_i_4__21_, pe_i_4__20_, pe_i_4__19_, pe_i_4__18_, pe_i_4__17_, pe_i_4__16_, pe_i_4__15_, pe_i_4__14_, pe_i_4__13_, pe_i_4__12_, pe_i_4__11_, pe_i_4__10_, pe_i_4__9_, pe_i_4__8_, pe_i_4__7_, pe_i_4__6_, pe_i_4__5_, pe_i_4__4_, pe_i_4__3_, pe_i_4__2_, pe_i_4__1_, pe_i_4__0_ }),
    .addr_o({ pe_o_4__4_, pe_o_4__3_, pe_o_4__2_, pe_o_4__1_, pe_o_4__0_ })
  );

  assign N484 = N0 & N1 & (N2 & N3) & N4;
  assign N0 = ~pe_o_1__4_;
  assign N1 = ~pe_o_1__3_;
  assign N2 = ~pe_o_1__2_;
  assign N3 = ~pe_o_1__0_;
  assign N4 = ~pe_o_1__1_;
  assign N485 = pe_o_1__4_ & N5 & (N6 & N7) & N8;
  assign N5 = ~pe_o_1__3_;
  assign N6 = ~pe_o_1__2_;
  assign N7 = ~pe_o_1__0_;
  assign N8 = ~pe_o_1__1_;
  assign N486 = N9 & N10 & (N11 & pe_o_1__0_) & N12;
  assign N9 = ~pe_o_1__4_;
  assign N10 = ~pe_o_1__3_;
  assign N11 = ~pe_o_1__2_;
  assign N12 = ~pe_o_1__1_;
  assign N488 = N13 & N14 & (N15 & N16) & pe_o_1__1_;
  assign N13 = ~pe_o_1__4_;
  assign N14 = ~pe_o_1__3_;
  assign N15 = ~pe_o_1__2_;
  assign N16 = ~pe_o_1__0_;
  assign N490 = N17 & N18 & (N19 & pe_o_1__0_) & pe_o_1__1_;
  assign N17 = ~pe_o_1__4_;
  assign N18 = ~pe_o_1__3_;
  assign N19 = ~pe_o_1__2_;
  assign N492 = N20 & N21 & (pe_o_1__2_ & N22) & N23;
  assign N20 = ~pe_o_1__4_;
  assign N21 = ~pe_o_1__3_;
  assign N22 = ~pe_o_1__0_;
  assign N23 = ~pe_o_1__1_;
  assign N494 = N24 & N25 & (pe_o_1__2_ & pe_o_1__0_) & N26;
  assign N24 = ~pe_o_1__4_;
  assign N25 = ~pe_o_1__3_;
  assign N26 = ~pe_o_1__1_;
  assign N496 = N27 & N28 & (pe_o_1__2_ & N29) & pe_o_1__1_;
  assign N27 = ~pe_o_1__4_;
  assign N28 = ~pe_o_1__3_;
  assign N29 = ~pe_o_1__0_;
  assign N498 = N30 & N31 & (pe_o_1__2_ & pe_o_1__0_) & pe_o_1__1_;
  assign N30 = ~pe_o_1__4_;
  assign N31 = ~pe_o_1__3_;
  assign N500 = N32 & pe_o_1__3_ & (N33 & N34) & N35;
  assign N32 = ~pe_o_1__4_;
  assign N33 = ~pe_o_1__2_;
  assign N34 = ~pe_o_1__0_;
  assign N35 = ~pe_o_1__1_;
  assign N502 = N36 & pe_o_1__3_ & (N37 & pe_o_1__0_) & N38;
  assign N36 = ~pe_o_1__4_;
  assign N37 = ~pe_o_1__2_;
  assign N38 = ~pe_o_1__1_;
  assign N504 = N39 & pe_o_1__3_ & (N40 & N41) & pe_o_1__1_;
  assign N39 = ~pe_o_1__4_;
  assign N40 = ~pe_o_1__2_;
  assign N41 = ~pe_o_1__0_;
  assign N506 = N42 & pe_o_1__3_ & (N43 & pe_o_1__0_) & pe_o_1__1_;
  assign N42 = ~pe_o_1__4_;
  assign N43 = ~pe_o_1__2_;
  assign N508 = N44 & pe_o_1__3_ & (pe_o_1__2_ & N45) & N46;
  assign N44 = ~pe_o_1__4_;
  assign N45 = ~pe_o_1__0_;
  assign N46 = ~pe_o_1__1_;
  assign N510 = N47 & pe_o_1__3_ & (pe_o_1__2_ & pe_o_1__0_) & N48;
  assign N47 = ~pe_o_1__4_;
  assign N48 = ~pe_o_1__1_;
  assign N512 = N49 & pe_o_1__3_ & (pe_o_1__2_ & N50) & pe_o_1__1_;
  assign N49 = ~pe_o_1__4_;
  assign N50 = ~pe_o_1__0_;
  assign N514 = pe_o_1__3_ & pe_o_1__2_ & (pe_o_1__0_ & pe_o_1__1_);
  assign N487 = pe_o_1__4_ & N51 & (N52 & pe_o_1__0_) & N53;
  assign N51 = ~pe_o_1__3_;
  assign N52 = ~pe_o_1__2_;
  assign N53 = ~pe_o_1__1_;
  assign N489 = pe_o_1__4_ & N54 & (N55 & N56) & pe_o_1__1_;
  assign N54 = ~pe_o_1__3_;
  assign N55 = ~pe_o_1__2_;
  assign N56 = ~pe_o_1__0_;
  assign N491 = pe_o_1__4_ & N57 & (N58 & pe_o_1__0_) & pe_o_1__1_;
  assign N57 = ~pe_o_1__3_;
  assign N58 = ~pe_o_1__2_;
  assign N493 = pe_o_1__4_ & N59 & (pe_o_1__2_ & N60) & N61;
  assign N59 = ~pe_o_1__3_;
  assign N60 = ~pe_o_1__0_;
  assign N61 = ~pe_o_1__1_;
  assign N495 = pe_o_1__4_ & N62 & (pe_o_1__2_ & pe_o_1__0_) & N63;
  assign N62 = ~pe_o_1__3_;
  assign N63 = ~pe_o_1__1_;
  assign N497 = pe_o_1__4_ & N64 & (pe_o_1__2_ & N65) & pe_o_1__1_;
  assign N64 = ~pe_o_1__3_;
  assign N65 = ~pe_o_1__0_;
  assign N499 = pe_o_1__4_ & pe_o_1__2_ & (pe_o_1__0_ & pe_o_1__1_);
  assign N501 = pe_o_1__4_ & pe_o_1__3_ & (N66 & N67) & N68;
  assign N66 = ~pe_o_1__2_;
  assign N67 = ~pe_o_1__0_;
  assign N68 = ~pe_o_1__1_;
  assign N503 = pe_o_1__4_ & pe_o_1__3_ & (N69 & pe_o_1__0_) & N70;
  assign N69 = ~pe_o_1__2_;
  assign N70 = ~pe_o_1__1_;
  assign N505 = pe_o_1__4_ & pe_o_1__3_ & (N71 & N72) & pe_o_1__1_;
  assign N71 = ~pe_o_1__2_;
  assign N72 = ~pe_o_1__0_;
  assign N507 = pe_o_1__4_ & pe_o_1__3_ & (pe_o_1__0_ & pe_o_1__1_);
  assign N509 = pe_o_1__4_ & pe_o_1__3_ & (pe_o_1__2_ & N73) & N74;
  assign N73 = ~pe_o_1__0_;
  assign N74 = ~pe_o_1__1_;
  assign N511 = pe_o_1__4_ & pe_o_1__3_ & (pe_o_1__2_ & pe_o_1__0_);
  assign N513 = pe_o_1__4_ & pe_o_1__3_ & (pe_o_1__2_ & pe_o_1__1_);
  assign N515 = N75 & N76 & (N77 & N78) & N79;
  assign N75 = ~pe_o_2__4_;
  assign N76 = ~pe_o_2__3_;
  assign N77 = ~pe_o_2__2_;
  assign N78 = ~pe_o_2__0_;
  assign N79 = ~pe_o_2__1_;
  assign N516 = pe_o_2__4_ & N80 & (N81 & N82) & N83;
  assign N80 = ~pe_o_2__3_;
  assign N81 = ~pe_o_2__2_;
  assign N82 = ~pe_o_2__0_;
  assign N83 = ~pe_o_2__1_;
  assign N517 = N84 & N85 & (N86 & pe_o_2__0_) & N87;
  assign N84 = ~pe_o_2__4_;
  assign N85 = ~pe_o_2__3_;
  assign N86 = ~pe_o_2__2_;
  assign N87 = ~pe_o_2__1_;
  assign N519 = N88 & N89 & (N90 & N91) & pe_o_2__1_;
  assign N88 = ~pe_o_2__4_;
  assign N89 = ~pe_o_2__3_;
  assign N90 = ~pe_o_2__2_;
  assign N91 = ~pe_o_2__0_;
  assign N521 = N92 & N93 & (N94 & pe_o_2__0_) & pe_o_2__1_;
  assign N92 = ~pe_o_2__4_;
  assign N93 = ~pe_o_2__3_;
  assign N94 = ~pe_o_2__2_;
  assign N523 = N95 & N96 & (pe_o_2__2_ & N97) & N98;
  assign N95 = ~pe_o_2__4_;
  assign N96 = ~pe_o_2__3_;
  assign N97 = ~pe_o_2__0_;
  assign N98 = ~pe_o_2__1_;
  assign N525 = N99 & N100 & (pe_o_2__2_ & pe_o_2__0_) & N101;
  assign N99 = ~pe_o_2__4_;
  assign N100 = ~pe_o_2__3_;
  assign N101 = ~pe_o_2__1_;
  assign N527 = N102 & N103 & (pe_o_2__2_ & N104) & pe_o_2__1_;
  assign N102 = ~pe_o_2__4_;
  assign N103 = ~pe_o_2__3_;
  assign N104 = ~pe_o_2__0_;
  assign N529 = N105 & N106 & (pe_o_2__2_ & pe_o_2__0_) & pe_o_2__1_;
  assign N105 = ~pe_o_2__4_;
  assign N106 = ~pe_o_2__3_;
  assign N531 = N107 & pe_o_2__3_ & (N108 & N109) & N110;
  assign N107 = ~pe_o_2__4_;
  assign N108 = ~pe_o_2__2_;
  assign N109 = ~pe_o_2__0_;
  assign N110 = ~pe_o_2__1_;
  assign N533 = N111 & pe_o_2__3_ & (N112 & pe_o_2__0_) & N113;
  assign N111 = ~pe_o_2__4_;
  assign N112 = ~pe_o_2__2_;
  assign N113 = ~pe_o_2__1_;
  assign N535 = N114 & pe_o_2__3_ & (N115 & N116) & pe_o_2__1_;
  assign N114 = ~pe_o_2__4_;
  assign N115 = ~pe_o_2__2_;
  assign N116 = ~pe_o_2__0_;
  assign N537 = N117 & pe_o_2__3_ & (N118 & pe_o_2__0_) & pe_o_2__1_;
  assign N117 = ~pe_o_2__4_;
  assign N118 = ~pe_o_2__2_;
  assign N539 = N119 & pe_o_2__3_ & (pe_o_2__2_ & N120) & N121;
  assign N119 = ~pe_o_2__4_;
  assign N120 = ~pe_o_2__0_;
  assign N121 = ~pe_o_2__1_;
  assign N541 = N122 & pe_o_2__3_ & (pe_o_2__2_ & pe_o_2__0_) & N123;
  assign N122 = ~pe_o_2__4_;
  assign N123 = ~pe_o_2__1_;
  assign N543 = N124 & pe_o_2__3_ & (pe_o_2__2_ & N125) & pe_o_2__1_;
  assign N124 = ~pe_o_2__4_;
  assign N125 = ~pe_o_2__0_;
  assign N545 = pe_o_2__3_ & pe_o_2__2_ & (pe_o_2__0_ & pe_o_2__1_);
  assign N518 = pe_o_2__4_ & N126 & (N127 & pe_o_2__0_) & N128;
  assign N126 = ~pe_o_2__3_;
  assign N127 = ~pe_o_2__2_;
  assign N128 = ~pe_o_2__1_;
  assign N520 = pe_o_2__4_ & N129 & (N130 & N131) & pe_o_2__1_;
  assign N129 = ~pe_o_2__3_;
  assign N130 = ~pe_o_2__2_;
  assign N131 = ~pe_o_2__0_;
  assign N522 = pe_o_2__4_ & N132 & (N133 & pe_o_2__0_) & pe_o_2__1_;
  assign N132 = ~pe_o_2__3_;
  assign N133 = ~pe_o_2__2_;
  assign N524 = pe_o_2__4_ & N134 & (pe_o_2__2_ & N135) & N136;
  assign N134 = ~pe_o_2__3_;
  assign N135 = ~pe_o_2__0_;
  assign N136 = ~pe_o_2__1_;
  assign N526 = pe_o_2__4_ & N137 & (pe_o_2__2_ & pe_o_2__0_) & N138;
  assign N137 = ~pe_o_2__3_;
  assign N138 = ~pe_o_2__1_;
  assign N528 = pe_o_2__4_ & N139 & (pe_o_2__2_ & N140) & pe_o_2__1_;
  assign N139 = ~pe_o_2__3_;
  assign N140 = ~pe_o_2__0_;
  assign N530 = pe_o_2__4_ & pe_o_2__2_ & (pe_o_2__0_ & pe_o_2__1_);
  assign N532 = pe_o_2__4_ & pe_o_2__3_ & (N141 & N142) & N143;
  assign N141 = ~pe_o_2__2_;
  assign N142 = ~pe_o_2__0_;
  assign N143 = ~pe_o_2__1_;
  assign N534 = pe_o_2__4_ & pe_o_2__3_ & (N144 & pe_o_2__0_) & N145;
  assign N144 = ~pe_o_2__2_;
  assign N145 = ~pe_o_2__1_;
  assign N536 = pe_o_2__4_ & pe_o_2__3_ & (N146 & N147) & pe_o_2__1_;
  assign N146 = ~pe_o_2__2_;
  assign N147 = ~pe_o_2__0_;
  assign N538 = pe_o_2__4_ & pe_o_2__3_ & (pe_o_2__0_ & pe_o_2__1_);
  assign N540 = pe_o_2__4_ & pe_o_2__3_ & (pe_o_2__2_ & N148) & N149;
  assign N148 = ~pe_o_2__0_;
  assign N149 = ~pe_o_2__1_;
  assign N542 = pe_o_2__4_ & pe_o_2__3_ & (pe_o_2__2_ & pe_o_2__0_);
  assign N544 = pe_o_2__4_ & pe_o_2__3_ & (pe_o_2__2_ & pe_o_2__1_);
  assign N577 = N150 & N151 & (N152 & N153) & N154;
  assign N150 = ~pe_o_3__4_;
  assign N151 = ~pe_o_3__3_;
  assign N152 = ~pe_o_3__2_;
  assign N153 = ~pe_o_3__0_;
  assign N154 = ~pe_o_3__1_;
  assign N578 = pe_o_3__4_ & N155 & (N156 & N157) & N158;
  assign N155 = ~pe_o_3__3_;
  assign N156 = ~pe_o_3__2_;
  assign N157 = ~pe_o_3__0_;
  assign N158 = ~pe_o_3__1_;
  assign N579 = N159 & N160 & (N161 & pe_o_3__0_) & N162;
  assign N159 = ~pe_o_3__4_;
  assign N160 = ~pe_o_3__3_;
  assign N161 = ~pe_o_3__2_;
  assign N162 = ~pe_o_3__1_;
  assign N581 = N163 & N164 & (N165 & N166) & pe_o_3__1_;
  assign N163 = ~pe_o_3__4_;
  assign N164 = ~pe_o_3__3_;
  assign N165 = ~pe_o_3__2_;
  assign N166 = ~pe_o_3__0_;
  assign N583 = N167 & N168 & (N169 & pe_o_3__0_) & pe_o_3__1_;
  assign N167 = ~pe_o_3__4_;
  assign N168 = ~pe_o_3__3_;
  assign N169 = ~pe_o_3__2_;
  assign N585 = N170 & N171 & (pe_o_3__2_ & N172) & N173;
  assign N170 = ~pe_o_3__4_;
  assign N171 = ~pe_o_3__3_;
  assign N172 = ~pe_o_3__0_;
  assign N173 = ~pe_o_3__1_;
  assign N587 = N174 & N175 & (pe_o_3__2_ & pe_o_3__0_) & N176;
  assign N174 = ~pe_o_3__4_;
  assign N175 = ~pe_o_3__3_;
  assign N176 = ~pe_o_3__1_;
  assign N589 = N177 & N178 & (pe_o_3__2_ & N179) & pe_o_3__1_;
  assign N177 = ~pe_o_3__4_;
  assign N178 = ~pe_o_3__3_;
  assign N179 = ~pe_o_3__0_;
  assign N591 = N180 & N181 & (pe_o_3__2_ & pe_o_3__0_) & pe_o_3__1_;
  assign N180 = ~pe_o_3__4_;
  assign N181 = ~pe_o_3__3_;
  assign N593 = N182 & pe_o_3__3_ & (N183 & N184) & N185;
  assign N182 = ~pe_o_3__4_;
  assign N183 = ~pe_o_3__2_;
  assign N184 = ~pe_o_3__0_;
  assign N185 = ~pe_o_3__1_;
  assign N595 = N186 & pe_o_3__3_ & (N187 & pe_o_3__0_) & N188;
  assign N186 = ~pe_o_3__4_;
  assign N187 = ~pe_o_3__2_;
  assign N188 = ~pe_o_3__1_;
  assign N597 = N189 & pe_o_3__3_ & (N190 & N191) & pe_o_3__1_;
  assign N189 = ~pe_o_3__4_;
  assign N190 = ~pe_o_3__2_;
  assign N191 = ~pe_o_3__0_;
  assign N599 = N192 & pe_o_3__3_ & (N193 & pe_o_3__0_) & pe_o_3__1_;
  assign N192 = ~pe_o_3__4_;
  assign N193 = ~pe_o_3__2_;
  assign N601 = N194 & pe_o_3__3_ & (pe_o_3__2_ & N195) & N196;
  assign N194 = ~pe_o_3__4_;
  assign N195 = ~pe_o_3__0_;
  assign N196 = ~pe_o_3__1_;
  assign N603 = N197 & pe_o_3__3_ & (pe_o_3__2_ & pe_o_3__0_) & N198;
  assign N197 = ~pe_o_3__4_;
  assign N198 = ~pe_o_3__1_;
  assign N605 = N199 & pe_o_3__3_ & (pe_o_3__2_ & N200) & pe_o_3__1_;
  assign N199 = ~pe_o_3__4_;
  assign N200 = ~pe_o_3__0_;
  assign N607 = pe_o_3__3_ & pe_o_3__2_ & (pe_o_3__0_ & pe_o_3__1_);
  assign N580 = pe_o_3__4_ & N201 & (N202 & pe_o_3__0_) & N203;
  assign N201 = ~pe_o_3__3_;
  assign N202 = ~pe_o_3__2_;
  assign N203 = ~pe_o_3__1_;
  assign N582 = pe_o_3__4_ & N204 & (N205 & N206) & pe_o_3__1_;
  assign N204 = ~pe_o_3__3_;
  assign N205 = ~pe_o_3__2_;
  assign N206 = ~pe_o_3__0_;
  assign N584 = pe_o_3__4_ & N207 & (N208 & pe_o_3__0_) & pe_o_3__1_;
  assign N207 = ~pe_o_3__3_;
  assign N208 = ~pe_o_3__2_;
  assign N586 = pe_o_3__4_ & N209 & (pe_o_3__2_ & N210) & N211;
  assign N209 = ~pe_o_3__3_;
  assign N210 = ~pe_o_3__0_;
  assign N211 = ~pe_o_3__1_;
  assign N588 = pe_o_3__4_ & N212 & (pe_o_3__2_ & pe_o_3__0_) & N213;
  assign N212 = ~pe_o_3__3_;
  assign N213 = ~pe_o_3__1_;
  assign N590 = pe_o_3__4_ & N214 & (pe_o_3__2_ & N215) & pe_o_3__1_;
  assign N214 = ~pe_o_3__3_;
  assign N215 = ~pe_o_3__0_;
  assign N592 = pe_o_3__4_ & pe_o_3__2_ & (pe_o_3__0_ & pe_o_3__1_);
  assign N594 = pe_o_3__4_ & pe_o_3__3_ & (N216 & N217) & N218;
  assign N216 = ~pe_o_3__2_;
  assign N217 = ~pe_o_3__0_;
  assign N218 = ~pe_o_3__1_;
  assign N596 = pe_o_3__4_ & pe_o_3__3_ & (N219 & pe_o_3__0_) & N220;
  assign N219 = ~pe_o_3__2_;
  assign N220 = ~pe_o_3__1_;
  assign N598 = pe_o_3__4_ & pe_o_3__3_ & (N221 & N222) & pe_o_3__1_;
  assign N221 = ~pe_o_3__2_;
  assign N222 = ~pe_o_3__0_;
  assign N600 = pe_o_3__4_ & pe_o_3__3_ & (pe_o_3__0_ & pe_o_3__1_);
  assign N602 = pe_o_3__4_ & pe_o_3__3_ & (pe_o_3__2_ & N223) & N224;
  assign N223 = ~pe_o_3__0_;
  assign N224 = ~pe_o_3__1_;
  assign N604 = pe_o_3__4_ & pe_o_3__3_ & (pe_o_3__2_ & pe_o_3__0_);
  assign N606 = pe_o_3__4_ & pe_o_3__3_ & (pe_o_3__2_ & pe_o_3__1_);
  assign N639 = N225 & N226 & (N227 & N228) & N229;
  assign N225 = ~pe_o_4__4_;
  assign N226 = ~pe_o_4__3_;
  assign N227 = ~pe_o_4__2_;
  assign N228 = ~pe_o_4__0_;
  assign N229 = ~pe_o_4__1_;
  assign N640 = pe_o_4__4_ & N230 & (N231 & N232) & N233;
  assign N230 = ~pe_o_4__3_;
  assign N231 = ~pe_o_4__2_;
  assign N232 = ~pe_o_4__0_;
  assign N233 = ~pe_o_4__1_;
  assign N641 = N234 & N235 & (N236 & pe_o_4__0_) & N237;
  assign N234 = ~pe_o_4__4_;
  assign N235 = ~pe_o_4__3_;
  assign N236 = ~pe_o_4__2_;
  assign N237 = ~pe_o_4__1_;
  assign N643 = N238 & N239 & (N240 & N241) & pe_o_4__1_;
  assign N238 = ~pe_o_4__4_;
  assign N239 = ~pe_o_4__3_;
  assign N240 = ~pe_o_4__2_;
  assign N241 = ~pe_o_4__0_;
  assign N645 = N242 & N243 & (N244 & pe_o_4__0_) & pe_o_4__1_;
  assign N242 = ~pe_o_4__4_;
  assign N243 = ~pe_o_4__3_;
  assign N244 = ~pe_o_4__2_;
  assign N647 = N245 & N246 & (pe_o_4__2_ & N247) & N248;
  assign N245 = ~pe_o_4__4_;
  assign N246 = ~pe_o_4__3_;
  assign N247 = ~pe_o_4__0_;
  assign N248 = ~pe_o_4__1_;
  assign N649 = N249 & N250 & (pe_o_4__2_ & pe_o_4__0_) & N251;
  assign N249 = ~pe_o_4__4_;
  assign N250 = ~pe_o_4__3_;
  assign N251 = ~pe_o_4__1_;
  assign N651 = N252 & N253 & (pe_o_4__2_ & N254) & pe_o_4__1_;
  assign N252 = ~pe_o_4__4_;
  assign N253 = ~pe_o_4__3_;
  assign N254 = ~pe_o_4__0_;
  assign N653 = N255 & N256 & (pe_o_4__2_ & pe_o_4__0_) & pe_o_4__1_;
  assign N255 = ~pe_o_4__4_;
  assign N256 = ~pe_o_4__3_;
  assign N655 = N257 & pe_o_4__3_ & (N258 & N259) & N260;
  assign N257 = ~pe_o_4__4_;
  assign N258 = ~pe_o_4__2_;
  assign N259 = ~pe_o_4__0_;
  assign N260 = ~pe_o_4__1_;
  assign N657 = N261 & pe_o_4__3_ & (N262 & pe_o_4__0_) & N263;
  assign N261 = ~pe_o_4__4_;
  assign N262 = ~pe_o_4__2_;
  assign N263 = ~pe_o_4__1_;
  assign N659 = N264 & pe_o_4__3_ & (N265 & N266) & pe_o_4__1_;
  assign N264 = ~pe_o_4__4_;
  assign N265 = ~pe_o_4__2_;
  assign N266 = ~pe_o_4__0_;
  assign N661 = N267 & pe_o_4__3_ & (N268 & pe_o_4__0_) & pe_o_4__1_;
  assign N267 = ~pe_o_4__4_;
  assign N268 = ~pe_o_4__2_;
  assign N663 = N269 & pe_o_4__3_ & (pe_o_4__2_ & N270) & N271;
  assign N269 = ~pe_o_4__4_;
  assign N270 = ~pe_o_4__0_;
  assign N271 = ~pe_o_4__1_;
  assign N665 = N272 & pe_o_4__3_ & (pe_o_4__2_ & pe_o_4__0_) & N273;
  assign N272 = ~pe_o_4__4_;
  assign N273 = ~pe_o_4__1_;
  assign N667 = N274 & pe_o_4__3_ & (pe_o_4__2_ & N275) & pe_o_4__1_;
  assign N274 = ~pe_o_4__4_;
  assign N275 = ~pe_o_4__0_;
  assign N669 = pe_o_4__3_ & pe_o_4__2_ & (pe_o_4__0_ & pe_o_4__1_);
  assign N642 = pe_o_4__4_ & N276 & (N277 & pe_o_4__0_) & N278;
  assign N276 = ~pe_o_4__3_;
  assign N277 = ~pe_o_4__2_;
  assign N278 = ~pe_o_4__1_;
  assign N644 = pe_o_4__4_ & N279 & (N280 & N281) & pe_o_4__1_;
  assign N279 = ~pe_o_4__3_;
  assign N280 = ~pe_o_4__2_;
  assign N281 = ~pe_o_4__0_;
  assign N646 = pe_o_4__4_ & N282 & (N283 & pe_o_4__0_) & pe_o_4__1_;
  assign N282 = ~pe_o_4__3_;
  assign N283 = ~pe_o_4__2_;
  assign N648 = pe_o_4__4_ & N284 & (pe_o_4__2_ & N285) & N286;
  assign N284 = ~pe_o_4__3_;
  assign N285 = ~pe_o_4__0_;
  assign N286 = ~pe_o_4__1_;
  assign N650 = pe_o_4__4_ & N287 & (pe_o_4__2_ & pe_o_4__0_) & N288;
  assign N287 = ~pe_o_4__3_;
  assign N288 = ~pe_o_4__1_;
  assign N652 = pe_o_4__4_ & N289 & (pe_o_4__2_ & N290) & pe_o_4__1_;
  assign N289 = ~pe_o_4__3_;
  assign N290 = ~pe_o_4__0_;
  assign N654 = pe_o_4__4_ & pe_o_4__2_ & (pe_o_4__0_ & pe_o_4__1_);
  assign N656 = pe_o_4__4_ & pe_o_4__3_ & (N291 & N292) & N293;
  assign N291 = ~pe_o_4__2_;
  assign N292 = ~pe_o_4__0_;
  assign N293 = ~pe_o_4__1_;
  assign N658 = pe_o_4__4_ & pe_o_4__3_ & (N294 & pe_o_4__0_) & N295;
  assign N294 = ~pe_o_4__2_;
  assign N295 = ~pe_o_4__1_;
  assign N660 = pe_o_4__4_ & pe_o_4__3_ & (N296 & N297) & pe_o_4__1_;
  assign N296 = ~pe_o_4__2_;
  assign N297 = ~pe_o_4__0_;
  assign N662 = pe_o_4__4_ & pe_o_4__3_ & (pe_o_4__0_ & pe_o_4__1_);
  assign N664 = pe_o_4__4_ & pe_o_4__3_ & (pe_o_4__2_ & N298) & N299;
  assign N298 = ~pe_o_4__0_;
  assign N299 = ~pe_o_4__1_;
  assign N666 = pe_o_4__4_ & pe_o_4__3_ & (pe_o_4__2_ & pe_o_4__0_);
  assign N668 = pe_o_4__4_ & pe_o_4__3_ & (pe_o_4__2_ & pe_o_4__1_);
  assign way_id_o[3] = (N300)? lru_i[0] : 
                       (N301)? lru_i[1] : 
                       (N302)? lru_i[2] : 
                       (N303)? lru_i[3] : 
                       (N304)? lru_i[4] : 
                       (N305)? lru_i[5] : 
                       (N306)? lru_i[6] : 
                       (N307)? lru_i[7] : 
                       (N308)? lru_i[8] : 
                       (N309)? lru_i[9] : 
                       (N310)? lru_i[10] : 
                       (N311)? lru_i[11] : 
                       (N312)? lru_i[12] : 
                       (N313)? lru_i[13] : 
                       (N314)? lru_i[14] : 
                       (N315)? lru_i[15] : 
                       (N316)? lru_i[16] : 
                       (N317)? lru_i[17] : 
                       (N318)? lru_i[18] : 
                       (N319)? lru_i[19] : 
                       (N320)? lru_i[20] : 
                       (N321)? lru_i[21] : 
                       (N322)? lru_i[22] : 
                       (N323)? lru_i[23] : 
                       (N324)? lru_i[24] : 
                       (N325)? lru_i[25] : 
                       (N326)? lru_i[26] : 
                       (N327)? lru_i[27] : 
                       (N328)? lru_i[28] : 
                       (N329)? lru_i[29] : 
                       (N330)? lru_i[30] : 1'b0;
  assign N300 = N484;
  assign N301 = N486;
  assign N302 = N488;
  assign N303 = N490;
  assign N304 = N492;
  assign N305 = N494;
  assign N306 = N496;
  assign N307 = N498;
  assign N308 = N500;
  assign N309 = N502;
  assign N310 = N504;
  assign N311 = N506;
  assign N312 = N508;
  assign N313 = N510;
  assign N314 = N512;
  assign N315 = N514;
  assign N316 = N485;
  assign N317 = N487;
  assign N318 = N489;
  assign N319 = N491;
  assign N320 = N493;
  assign N321 = N495;
  assign N322 = N497;
  assign N323 = N499;
  assign N324 = N501;
  assign N325 = N503;
  assign N326 = N505;
  assign N327 = N507;
  assign N328 = N509;
  assign N329 = N511;
  assign N330 = N513;
  assign way_id_o[2] = (N331)? lru_i[0] : 
                       (N332)? lru_i[1] : 
                       (N333)? lru_i[2] : 
                       (N334)? lru_i[3] : 
                       (N335)? lru_i[4] : 
                       (N336)? lru_i[5] : 
                       (N337)? lru_i[6] : 
                       (N338)? lru_i[7] : 
                       (N339)? lru_i[8] : 
                       (N340)? lru_i[9] : 
                       (N341)? lru_i[10] : 
                       (N342)? lru_i[11] : 
                       (N343)? lru_i[12] : 
                       (N344)? lru_i[13] : 
                       (N345)? lru_i[14] : 
                       (N346)? lru_i[15] : 
                       (N347)? lru_i[16] : 
                       (N348)? lru_i[17] : 
                       (N349)? lru_i[18] : 
                       (N350)? lru_i[19] : 
                       (N351)? lru_i[20] : 
                       (N352)? lru_i[21] : 
                       (N353)? lru_i[22] : 
                       (N354)? lru_i[23] : 
                       (N355)? lru_i[24] : 
                       (N356)? lru_i[25] : 
                       (N357)? lru_i[26] : 
                       (N358)? lru_i[27] : 
                       (N359)? lru_i[28] : 
                       (N360)? lru_i[29] : 
                       (N361)? lru_i[30] : 1'b0;
  assign N331 = N515;
  assign N332 = N517;
  assign N333 = N519;
  assign N334 = N521;
  assign N335 = N523;
  assign N336 = N525;
  assign N337 = N527;
  assign N338 = N529;
  assign N339 = N531;
  assign N340 = N533;
  assign N341 = N535;
  assign N342 = N537;
  assign N343 = N539;
  assign N344 = N541;
  assign N345 = N543;
  assign N346 = N545;
  assign N347 = N516;
  assign N348 = N518;
  assign N349 = N520;
  assign N350 = N522;
  assign N351 = N524;
  assign N352 = N526;
  assign N353 = N528;
  assign N354 = N530;
  assign N355 = N532;
  assign N356 = N534;
  assign N357 = N536;
  assign N358 = N538;
  assign N359 = N540;
  assign N360 = N542;
  assign N361 = N544;
  assign way_id_o[1] = (N362)? lru_i[0] : 
                       (N363)? lru_i[1] : 
                       (N364)? lru_i[2] : 
                       (N365)? lru_i[3] : 
                       (N366)? lru_i[4] : 
                       (N367)? lru_i[5] : 
                       (N368)? lru_i[6] : 
                       (N369)? lru_i[7] : 
                       (N370)? lru_i[8] : 
                       (N371)? lru_i[9] : 
                       (N372)? lru_i[10] : 
                       (N373)? lru_i[11] : 
                       (N374)? lru_i[12] : 
                       (N375)? lru_i[13] : 
                       (N376)? lru_i[14] : 
                       (N377)? lru_i[15] : 
                       (N378)? lru_i[16] : 
                       (N379)? lru_i[17] : 
                       (N380)? lru_i[18] : 
                       (N381)? lru_i[19] : 
                       (N382)? lru_i[20] : 
                       (N383)? lru_i[21] : 
                       (N384)? lru_i[22] : 
                       (N385)? lru_i[23] : 
                       (N386)? lru_i[24] : 
                       (N387)? lru_i[25] : 
                       (N388)? lru_i[26] : 
                       (N389)? lru_i[27] : 
                       (N390)? lru_i[28] : 
                       (N391)? lru_i[29] : 
                       (N392)? lru_i[30] : 1'b0;
  assign N362 = N577;
  assign N363 = N579;
  assign N364 = N581;
  assign N365 = N583;
  assign N366 = N585;
  assign N367 = N587;
  assign N368 = N589;
  assign N369 = N591;
  assign N370 = N593;
  assign N371 = N595;
  assign N372 = N597;
  assign N373 = N599;
  assign N374 = N601;
  assign N375 = N603;
  assign N376 = N605;
  assign N377 = N607;
  assign N378 = N578;
  assign N379 = N580;
  assign N380 = N582;
  assign N381 = N584;
  assign N382 = N586;
  assign N383 = N588;
  assign N384 = N590;
  assign N385 = N592;
  assign N386 = N594;
  assign N387 = N596;
  assign N388 = N598;
  assign N389 = N600;
  assign N390 = N602;
  assign N391 = N604;
  assign N392 = N606;
  assign way_id_o[0] = (N393)? lru_i[0] : 
                       (N394)? lru_i[1] : 
                       (N395)? lru_i[2] : 
                       (N396)? lru_i[3] : 
                       (N397)? lru_i[4] : 
                       (N398)? lru_i[5] : 
                       (N399)? lru_i[6] : 
                       (N400)? lru_i[7] : 
                       (N401)? lru_i[8] : 
                       (N402)? lru_i[9] : 
                       (N403)? lru_i[10] : 
                       (N404)? lru_i[11] : 
                       (N405)? lru_i[12] : 
                       (N406)? lru_i[13] : 
                       (N407)? lru_i[14] : 
                       (N408)? lru_i[15] : 
                       (N409)? lru_i[16] : 
                       (N410)? lru_i[17] : 
                       (N411)? lru_i[18] : 
                       (N412)? lru_i[19] : 
                       (N413)? lru_i[20] : 
                       (N414)? lru_i[21] : 
                       (N415)? lru_i[22] : 
                       (N416)? lru_i[23] : 
                       (N417)? lru_i[24] : 
                       (N418)? lru_i[25] : 
                       (N419)? lru_i[26] : 
                       (N420)? lru_i[27] : 
                       (N421)? lru_i[28] : 
                       (N422)? lru_i[29] : 
                       (N423)? lru_i[30] : 1'b0;
  assign N393 = N639;
  assign N394 = N641;
  assign N395 = N643;
  assign N396 = N645;
  assign N397 = N647;
  assign N398 = N649;
  assign N399 = N651;
  assign N400 = N653;
  assign N401 = N655;
  assign N402 = N657;
  assign N403 = N659;
  assign N404 = N661;
  assign N405 = N663;
  assign N406 = N665;
  assign N407 = N667;
  assign N408 = N669;
  assign N409 = N640;
  assign N410 = N642;
  assign N411 = N644;
  assign N412 = N646;
  assign N413 = N648;
  assign N414 = N650;
  assign N415 = N652;
  assign N416 = N654;
  assign N417 = N656;
  assign N418 = N658;
  assign N419 = N660;
  assign N420 = N662;
  assign N421 = N664;
  assign N422 = N666;
  assign N423 = N668;
  assign way_id_o[4] = (N453)? lru_i[0] : 
                       (N455)? lru_i[1] : 
                       (N457)? lru_i[2] : 
                       (N459)? lru_i[3] : 
                       (N461)? lru_i[4] : 
                       (N463)? lru_i[5] : 
                       (N465)? lru_i[6] : 
                       (N467)? lru_i[7] : 
                       (N469)? lru_i[8] : 
                       (N471)? lru_i[9] : 
                       (N473)? lru_i[10] : 
                       (N475)? lru_i[11] : 
                       (N477)? lru_i[12] : 
                       (N479)? lru_i[13] : 
                       (N481)? lru_i[14] : 
                       (N483)? lru_i[15] : 
                       (N454)? lru_i[16] : 
                       (N456)? lru_i[17] : 
                       (N458)? lru_i[18] : 
                       (N460)? lru_i[19] : 
                       (N462)? lru_i[20] : 
                       (N464)? lru_i[21] : 
                       (N466)? lru_i[22] : 
                       (N468)? lru_i[23] : 
                       (N470)? lru_i[24] : 
                       (N472)? lru_i[25] : 
                       (N474)? lru_i[26] : 
                       (N476)? lru_i[27] : 
                       (N478)? lru_i[28] : 
                       (N480)? lru_i[29] : 
                       (N482)? lru_i[30] : 1'b0;
  assign mask[1] = 1'b1 & N701;
  assign N701 = ~lru_i[0];
  assign mask[2] = 1'b1 & lru_i[0];
  assign mask[3] = mask[1] & N702;
  assign N702 = ~lru_i[1];
  assign mask[4] = mask[1] & lru_i[1];
  assign mask[5] = mask[2] & N703;
  assign N703 = ~lru_i[2];
  assign mask[6] = mask[2] & lru_i[2];
  assign mask[7] = mask[3] & N704;
  assign N704 = ~lru_i[3];
  assign mask[8] = mask[3] & lru_i[3];
  assign mask[9] = mask[4] & N705;
  assign N705 = ~lru_i[4];
  assign mask[10] = mask[4] & lru_i[4];
  assign mask[11] = mask[5] & N706;
  assign N706 = ~lru_i[5];
  assign mask[12] = mask[5] & lru_i[5];
  assign mask[13] = mask[6] & N707;
  assign N707 = ~lru_i[6];
  assign mask[14] = mask[6] & lru_i[6];
  assign mask[15] = mask[7] & N708;
  assign N708 = ~lru_i[7];
  assign mask[16] = mask[7] & lru_i[7];
  assign mask[17] = mask[8] & N709;
  assign N709 = ~lru_i[8];
  assign mask[18] = mask[8] & lru_i[8];
  assign mask[19] = mask[9] & N710;
  assign N710 = ~lru_i[9];
  assign mask[20] = mask[9] & lru_i[9];
  assign mask[21] = mask[10] & N711;
  assign N711 = ~lru_i[10];
  assign mask[22] = mask[10] & lru_i[10];
  assign mask[23] = mask[11] & N712;
  assign N712 = ~lru_i[11];
  assign mask[24] = mask[11] & lru_i[11];
  assign mask[25] = mask[12] & N713;
  assign N713 = ~lru_i[12];
  assign mask[26] = mask[12] & lru_i[12];
  assign mask[27] = mask[13] & N714;
  assign N714 = ~lru_i[13];
  assign mask[28] = mask[13] & lru_i[13];
  assign mask[29] = mask[14] & N715;
  assign N715 = ~lru_i[14];
  assign mask[30] = mask[14] & lru_i[14];
  assign N424 = N452 & N452;
  assign N425 = N452 & 1'b0;
  assign N426 = 1'b0 & N452;
  assign N427 = 1'b0 & 1'b0;
  assign N428 = N424 & N452;
  assign N429 = N424 & 1'b0;
  assign N430 = N426 & N452;
  assign N431 = N426 & 1'b0;
  assign N432 = N425 & N452;
  assign N433 = N425 & 1'b0;
  assign N434 = N427 & N452;
  assign N435 = N427 & 1'b0;
  assign N436 = N428 & N452;
  assign N437 = N428 & 1'b0;
  assign N438 = N430 & N452;
  assign N439 = N430 & 1'b0;
  assign N440 = N432 & N452;
  assign N441 = N432 & 1'b0;
  assign N442 = N434 & N452;
  assign N443 = N434 & 1'b0;
  assign N444 = N429 & N452;
  assign N445 = N429 & 1'b0;
  assign N446 = N431 & N452;
  assign N447 = N431 & 1'b0;
  assign N448 = N433 & N452;
  assign N449 = N433 & 1'b0;
  assign N450 = N435 & N452;
  assign N451 = N435 & 1'b0;
  assign N452 = ~1'b0;
  assign N453 = N436 & N452;
  assign N454 = N436 & 1'b0;
  assign N455 = N438 & N452;
  assign N456 = N438 & 1'b0;
  assign N457 = N440 & N452;
  assign N458 = N440 & 1'b0;
  assign N459 = N442 & N452;
  assign N460 = N442 & 1'b0;
  assign N461 = N444 & N452;
  assign N462 = N444 & 1'b0;
  assign N463 = N446 & N452;
  assign N464 = N446 & 1'b0;
  assign N465 = N448 & N452;
  assign N466 = N448 & 1'b0;
  assign N467 = N450 & N452;
  assign N468 = N450 & 1'b0;
  assign N469 = N437 & N452;
  assign N470 = N437 & 1'b0;
  assign N471 = N439 & N452;
  assign N472 = N439 & 1'b0;
  assign N473 = N441 & N452;
  assign N474 = N441 & 1'b0;
  assign N475 = N443 & N452;
  assign N476 = N443 & 1'b0;
  assign N477 = N445 & N452;
  assign N478 = N445 & 1'b0;
  assign N479 = N447 & N452;
  assign N480 = N447 & 1'b0;
  assign N481 = N449 & N452;
  assign N482 = N449 & 1'b0;
  assign N483 = N451 & N452;
  assign pe_i_1__30_ = mask[30] ^ 1'b0;
  assign pe_i_1__29_ = mask[29] ^ 1'b0;
  assign pe_i_1__28_ = mask[28] ^ 1'b0;
  assign pe_i_1__27_ = mask[27] ^ 1'b0;
  assign pe_i_1__26_ = mask[26] ^ 1'b0;
  assign pe_i_1__25_ = mask[25] ^ 1'b0;
  assign pe_i_1__24_ = mask[24] ^ 1'b0;
  assign pe_i_1__23_ = mask[23] ^ 1'b0;
  assign pe_i_1__22_ = mask[22] ^ 1'b0;
  assign pe_i_1__21_ = mask[21] ^ 1'b0;
  assign pe_i_1__20_ = mask[20] ^ 1'b0;
  assign pe_i_1__19_ = mask[19] ^ 1'b0;
  assign pe_i_1__18_ = mask[18] ^ 1'b0;
  assign pe_i_1__17_ = mask[17] ^ 1'b0;
  assign pe_i_1__16_ = mask[16] ^ 1'b0;
  assign pe_i_1__15_ = mask[15] ^ 1'b0;
  assign pe_i_1__14_ = mask[14] ^ 1'b0;
  assign pe_i_1__13_ = mask[13] ^ 1'b0;
  assign pe_i_1__12_ = mask[12] ^ 1'b0;
  assign pe_i_1__11_ = mask[11] ^ 1'b0;
  assign pe_i_1__10_ = mask[10] ^ 1'b0;
  assign pe_i_1__9_ = mask[9] ^ 1'b0;
  assign pe_i_1__8_ = mask[8] ^ 1'b0;
  assign pe_i_1__7_ = mask[7] ^ 1'b0;
  assign pe_i_1__6_ = mask[6] ^ 1'b0;
  assign pe_i_1__5_ = mask[5] ^ 1'b0;
  assign pe_i_1__4_ = mask[4] ^ 1'b0;
  assign pe_i_1__3_ = mask[3] ^ 1'b0;
  assign pe_i_1__2_ = mask[2] ^ 1'b0;
  assign pe_i_1__1_ = mask[1] ^ 1'b0;
  assign pe_i_1__0_ = 1'b1 ^ 1'b1;
  assign pe_i_2__30_ = pe_i_1__30_ ^ N576;
  assign pe_i_2__29_ = pe_i_1__29_ ^ N575;
  assign pe_i_2__28_ = pe_i_1__28_ ^ N574;
  assign pe_i_2__27_ = pe_i_1__27_ ^ N573;
  assign pe_i_2__26_ = pe_i_1__26_ ^ N572;
  assign pe_i_2__25_ = pe_i_1__25_ ^ N571;
  assign pe_i_2__24_ = pe_i_1__24_ ^ N570;
  assign pe_i_2__23_ = pe_i_1__23_ ^ N569;
  assign pe_i_2__22_ = pe_i_1__22_ ^ N568;
  assign pe_i_2__21_ = pe_i_1__21_ ^ N567;
  assign pe_i_2__20_ = pe_i_1__20_ ^ N566;
  assign pe_i_2__19_ = pe_i_1__19_ ^ N565;
  assign pe_i_2__18_ = pe_i_1__18_ ^ N564;
  assign pe_i_2__17_ = pe_i_1__17_ ^ N563;
  assign pe_i_2__16_ = pe_i_1__16_ ^ N562;
  assign pe_i_2__15_ = pe_i_1__15_ ^ N561;
  assign pe_i_2__14_ = pe_i_1__14_ ^ N560;
  assign pe_i_2__13_ = pe_i_1__13_ ^ N559;
  assign pe_i_2__12_ = pe_i_1__12_ ^ N558;
  assign pe_i_2__11_ = pe_i_1__11_ ^ N557;
  assign pe_i_2__10_ = pe_i_1__10_ ^ N556;
  assign pe_i_2__9_ = pe_i_1__9_ ^ N555;
  assign pe_i_2__8_ = pe_i_1__8_ ^ N554;
  assign pe_i_2__7_ = pe_i_1__7_ ^ N553;
  assign pe_i_2__6_ = pe_i_1__6_ ^ N552;
  assign pe_i_2__5_ = pe_i_1__5_ ^ N551;
  assign pe_i_2__4_ = pe_i_1__4_ ^ N550;
  assign pe_i_2__3_ = pe_i_1__3_ ^ N549;
  assign pe_i_2__2_ = pe_i_1__2_ ^ N548;
  assign pe_i_2__1_ = pe_i_1__1_ ^ N547;
  assign pe_i_2__0_ = pe_i_1__0_ ^ N546;
  assign pe_i_3__30_ = pe_i_2__30_ ^ N638;
  assign pe_i_3__29_ = pe_i_2__29_ ^ N637;
  assign pe_i_3__28_ = pe_i_2__28_ ^ N636;
  assign pe_i_3__27_ = pe_i_2__27_ ^ N635;
  assign pe_i_3__26_ = pe_i_2__26_ ^ N634;
  assign pe_i_3__25_ = pe_i_2__25_ ^ N633;
  assign pe_i_3__24_ = pe_i_2__24_ ^ N632;
  assign pe_i_3__23_ = pe_i_2__23_ ^ N631;
  assign pe_i_3__22_ = pe_i_2__22_ ^ N630;
  assign pe_i_3__21_ = pe_i_2__21_ ^ N629;
  assign pe_i_3__20_ = pe_i_2__20_ ^ N628;
  assign pe_i_3__19_ = pe_i_2__19_ ^ N627;
  assign pe_i_3__18_ = pe_i_2__18_ ^ N626;
  assign pe_i_3__17_ = pe_i_2__17_ ^ N625;
  assign pe_i_3__16_ = pe_i_2__16_ ^ N624;
  assign pe_i_3__15_ = pe_i_2__15_ ^ N623;
  assign pe_i_3__14_ = pe_i_2__14_ ^ N622;
  assign pe_i_3__13_ = pe_i_2__13_ ^ N621;
  assign pe_i_3__12_ = pe_i_2__12_ ^ N620;
  assign pe_i_3__11_ = pe_i_2__11_ ^ N619;
  assign pe_i_3__10_ = pe_i_2__10_ ^ N618;
  assign pe_i_3__9_ = pe_i_2__9_ ^ N617;
  assign pe_i_3__8_ = pe_i_2__8_ ^ N616;
  assign pe_i_3__7_ = pe_i_2__7_ ^ N615;
  assign pe_i_3__6_ = pe_i_2__6_ ^ N614;
  assign pe_i_3__5_ = pe_i_2__5_ ^ N613;
  assign pe_i_3__4_ = pe_i_2__4_ ^ N612;
  assign pe_i_3__3_ = pe_i_2__3_ ^ N611;
  assign pe_i_3__2_ = pe_i_2__2_ ^ N610;
  assign pe_i_3__1_ = pe_i_2__1_ ^ N609;
  assign pe_i_3__0_ = pe_i_2__0_ ^ N608;
  assign pe_i_4__30_ = pe_i_3__30_ ^ N700;
  assign pe_i_4__29_ = pe_i_3__29_ ^ N699;
  assign pe_i_4__28_ = pe_i_3__28_ ^ N698;
  assign pe_i_4__27_ = pe_i_3__27_ ^ N697;
  assign pe_i_4__26_ = pe_i_3__26_ ^ N696;
  assign pe_i_4__25_ = pe_i_3__25_ ^ N695;
  assign pe_i_4__24_ = pe_i_3__24_ ^ N694;
  assign pe_i_4__23_ = pe_i_3__23_ ^ N693;
  assign pe_i_4__22_ = pe_i_3__22_ ^ N692;
  assign pe_i_4__21_ = pe_i_3__21_ ^ N691;
  assign pe_i_4__20_ = pe_i_3__20_ ^ N690;
  assign pe_i_4__19_ = pe_i_3__19_ ^ N689;
  assign pe_i_4__18_ = pe_i_3__18_ ^ N688;
  assign pe_i_4__17_ = pe_i_3__17_ ^ N687;
  assign pe_i_4__16_ = pe_i_3__16_ ^ N686;
  assign pe_i_4__15_ = pe_i_3__15_ ^ N685;
  assign pe_i_4__14_ = pe_i_3__14_ ^ N684;
  assign pe_i_4__13_ = pe_i_3__13_ ^ N683;
  assign pe_i_4__12_ = pe_i_3__12_ ^ N682;
  assign pe_i_4__11_ = pe_i_3__11_ ^ N681;
  assign pe_i_4__10_ = pe_i_3__10_ ^ N680;
  assign pe_i_4__9_ = pe_i_3__9_ ^ N679;
  assign pe_i_4__8_ = pe_i_3__8_ ^ N678;
  assign pe_i_4__7_ = pe_i_3__7_ ^ N677;
  assign pe_i_4__6_ = pe_i_3__6_ ^ N676;
  assign pe_i_4__5_ = pe_i_3__5_ ^ N675;
  assign pe_i_4__4_ = pe_i_3__4_ ^ N674;
  assign pe_i_4__3_ = pe_i_3__3_ ^ N673;
  assign pe_i_4__2_ = pe_i_3__2_ ^ N672;
  assign pe_i_4__1_ = pe_i_3__1_ ^ N671;
  assign pe_i_4__0_ = pe_i_3__0_ ^ N670;

endmodule

