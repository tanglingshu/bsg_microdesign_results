

module top
(
  clk_i,
  reset_i,
  en_i,
  w_v_i,
  w_set_not_clear_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_data_i,
  r_v_o,
  r_addr_o,
  empty_v_o,
  empty_addr_o
);

  input [8:0] w_addr_i;
  input [15:0] w_data_i;
  input [15:0] r_data_i;
  output [8:0] r_addr_o;
  output [8:0] empty_addr_o;
  input clk_i;
  input reset_i;
  input en_i;
  input w_v_i;
  input w_set_not_clear_i;
  input r_v_i;
  output r_v_o;
  output empty_v_o;

  bsg_cam_1r1w
  wrapper
  (
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_data_i(r_data_i),
    .r_addr_o(r_addr_o),
    .empty_addr_o(empty_addr_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(en_i),
    .w_v_i(w_v_i),
    .w_set_not_clear_i(w_set_not_clear_i),
    .r_v_i(r_v_i),
    .r_v_o(r_v_o),
    .empty_v_o(empty_v_o)
  );


endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_encode_one_hot_width_p8
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_encode_one_hot_width_p16
(
  i,
  addr_o,
  v_o
);

  input [15:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o;
  wire [5:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p8
  aligned_left
  (
    .i(i[7:0]),
    .addr_o(aligned_addrs[2:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p8
  aligned_right
  (
    .i(i[15:8]),
    .addr_o(aligned_addrs[5:3]),
    .v_o(addr_o[3])
  );

  assign v_o = addr_o[3] | aligned_vs[0];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[5];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[4];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[3];

endmodule



module bsg_encode_one_hot_width_p32
(
  i,
  addr_o,
  v_o
);

  input [31:0] i;
  output [4:0] addr_o;
  output v_o;
  wire [4:0] addr_o;
  wire v_o;
  wire [7:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p16
  aligned_left
  (
    .i(i[15:0]),
    .addr_o(aligned_addrs[3:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p16
  aligned_right
  (
    .i(i[31:16]),
    .addr_o(aligned_addrs[7:4]),
    .v_o(addr_o[4])
  );

  assign v_o = addr_o[4] | aligned_vs[0];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[7];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[6];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[5];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[4];

endmodule



module bsg_encode_one_hot_width_p64
(
  i,
  addr_o,
  v_o
);

  input [63:0] i;
  output [5:0] addr_o;
  output v_o;
  wire [5:0] addr_o;
  wire v_o;
  wire [9:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p32
  aligned_left
  (
    .i(i[31:0]),
    .addr_o(aligned_addrs[4:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p32
  aligned_right
  (
    .i(i[63:32]),
    .addr_o(aligned_addrs[9:5]),
    .v_o(addr_o[5])
  );

  assign v_o = addr_o[5] | aligned_vs[0];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[9];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[8];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[7];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[6];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[5];

endmodule



module bsg_encode_one_hot_width_p128
(
  i,
  addr_o,
  v_o
);

  input [127:0] i;
  output [6:0] addr_o;
  output v_o;
  wire [6:0] addr_o;
  wire v_o;
  wire [11:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p64
  aligned_left
  (
    .i(i[63:0]),
    .addr_o(aligned_addrs[5:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p64
  aligned_right
  (
    .i(i[127:64]),
    .addr_o(aligned_addrs[11:6]),
    .v_o(addr_o[6])
  );

  assign v_o = addr_o[6] | aligned_vs[0];
  assign addr_o[5] = aligned_addrs[5] | aligned_addrs[11];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[10];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[9];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[8];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[7];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[6];

endmodule



module bsg_encode_one_hot_width_p256
(
  i,
  addr_o,
  v_o
);

  input [255:0] i;
  output [7:0] addr_o;
  output v_o;
  wire [7:0] addr_o;
  wire v_o;
  wire [13:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p128
  aligned_left
  (
    .i(i[127:0]),
    .addr_o(aligned_addrs[6:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p128
  aligned_right
  (
    .i(i[255:128]),
    .addr_o(aligned_addrs[13:7]),
    .v_o(addr_o[7])
  );

  assign v_o = addr_o[7] | aligned_vs[0];
  assign addr_o[6] = aligned_addrs[6] | aligned_addrs[13];
  assign addr_o[5] = aligned_addrs[5] | aligned_addrs[12];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[11];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[10];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[9];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[8];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[7];

endmodule



module bsg_encode_one_hot_width_p512_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [511:0] i;
  output [8:0] addr_o;
  output v_o;
  wire [8:0] addr_o;
  wire v_o;
  wire [15:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p256
  aligned_left
  (
    .i(i[255:0]),
    .addr_o(aligned_addrs[7:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p256
  aligned_right
  (
    .i(i[511:256]),
    .addr_o(aligned_addrs[15:8]),
    .v_o(addr_o[8])
  );

  assign v_o = addr_o[8] | aligned_vs[0];
  assign addr_o[7] = aligned_addrs[7] | aligned_addrs[15];
  assign addr_o[6] = aligned_addrs[6] | aligned_addrs[14];
  assign addr_o[5] = aligned_addrs[5] | aligned_addrs[13];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[12];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[11];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[10];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[9];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[8];

endmodule



module bsg_scan_width_p512_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [511:0] i;
  output [511:0] o;
  wire [511:0] o;
  wire t_1__511_,t_1__510_,t_1__509_,t_1__508_,t_1__507_,t_1__506_,t_1__505_,t_1__504_,
  t_1__503_,t_1__502_,t_1__501_,t_1__500_,t_1__499_,t_1__498_,t_1__497_,t_1__496_,
  t_1__495_,t_1__494_,t_1__493_,t_1__492_,t_1__491_,t_1__490_,t_1__489_,t_1__488_,
  t_1__487_,t_1__486_,t_1__485_,t_1__484_,t_1__483_,t_1__482_,t_1__481_,t_1__480_,
  t_1__479_,t_1__478_,t_1__477_,t_1__476_,t_1__475_,t_1__474_,t_1__473_,t_1__472_,
  t_1__471_,t_1__470_,t_1__469_,t_1__468_,t_1__467_,t_1__466_,t_1__465_,t_1__464_,
  t_1__463_,t_1__462_,t_1__461_,t_1__460_,t_1__459_,t_1__458_,t_1__457_,t_1__456_,
  t_1__455_,t_1__454_,t_1__453_,t_1__452_,t_1__451_,t_1__450_,t_1__449_,t_1__448_,
  t_1__447_,t_1__446_,t_1__445_,t_1__444_,t_1__443_,t_1__442_,t_1__441_,t_1__440_,
  t_1__439_,t_1__438_,t_1__437_,t_1__436_,t_1__435_,t_1__434_,t_1__433_,t_1__432_,
  t_1__431_,t_1__430_,t_1__429_,t_1__428_,t_1__427_,t_1__426_,t_1__425_,t_1__424_,
  t_1__423_,t_1__422_,t_1__421_,t_1__420_,t_1__419_,t_1__418_,t_1__417_,t_1__416_,
  t_1__415_,t_1__414_,t_1__413_,t_1__412_,t_1__411_,t_1__410_,t_1__409_,t_1__408_,
  t_1__407_,t_1__406_,t_1__405_,t_1__404_,t_1__403_,t_1__402_,t_1__401_,t_1__400_,
  t_1__399_,t_1__398_,t_1__397_,t_1__396_,t_1__395_,t_1__394_,t_1__393_,t_1__392_,
  t_1__391_,t_1__390_,t_1__389_,t_1__388_,t_1__387_,t_1__386_,t_1__385_,t_1__384_,
  t_1__383_,t_1__382_,t_1__381_,t_1__380_,t_1__379_,t_1__378_,t_1__377_,t_1__376_,
  t_1__375_,t_1__374_,t_1__373_,t_1__372_,t_1__371_,t_1__370_,t_1__369_,t_1__368_,
  t_1__367_,t_1__366_,t_1__365_,t_1__364_,t_1__363_,t_1__362_,t_1__361_,t_1__360_,
  t_1__359_,t_1__358_,t_1__357_,t_1__356_,t_1__355_,t_1__354_,t_1__353_,t_1__352_,
  t_1__351_,t_1__350_,t_1__349_,t_1__348_,t_1__347_,t_1__346_,t_1__345_,t_1__344_,
  t_1__343_,t_1__342_,t_1__341_,t_1__340_,t_1__339_,t_1__338_,t_1__337_,t_1__336_,
  t_1__335_,t_1__334_,t_1__333_,t_1__332_,t_1__331_,t_1__330_,t_1__329_,t_1__328_,
  t_1__327_,t_1__326_,t_1__325_,t_1__324_,t_1__323_,t_1__322_,t_1__321_,t_1__320_,
  t_1__319_,t_1__318_,t_1__317_,t_1__316_,t_1__315_,t_1__314_,t_1__313_,t_1__312_,
  t_1__311_,t_1__310_,t_1__309_,t_1__308_,t_1__307_,t_1__306_,t_1__305_,t_1__304_,
  t_1__303_,t_1__302_,t_1__301_,t_1__300_,t_1__299_,t_1__298_,t_1__297_,t_1__296_,
  t_1__295_,t_1__294_,t_1__293_,t_1__292_,t_1__291_,t_1__290_,t_1__289_,t_1__288_,
  t_1__287_,t_1__286_,t_1__285_,t_1__284_,t_1__283_,t_1__282_,t_1__281_,t_1__280_,
  t_1__279_,t_1__278_,t_1__277_,t_1__276_,t_1__275_,t_1__274_,t_1__273_,t_1__272_,
  t_1__271_,t_1__270_,t_1__269_,t_1__268_,t_1__267_,t_1__266_,t_1__265_,t_1__264_,
  t_1__263_,t_1__262_,t_1__261_,t_1__260_,t_1__259_,t_1__258_,t_1__257_,t_1__256_,
  t_1__255_,t_1__254_,t_1__253_,t_1__252_,t_1__251_,t_1__250_,t_1__249_,t_1__248_,
  t_1__247_,t_1__246_,t_1__245_,t_1__244_,t_1__243_,t_1__242_,t_1__241_,t_1__240_,
  t_1__239_,t_1__238_,t_1__237_,t_1__236_,t_1__235_,t_1__234_,t_1__233_,t_1__232_,
  t_1__231_,t_1__230_,t_1__229_,t_1__228_,t_1__227_,t_1__226_,t_1__225_,t_1__224_,
  t_1__223_,t_1__222_,t_1__221_,t_1__220_,t_1__219_,t_1__218_,t_1__217_,t_1__216_,
  t_1__215_,t_1__214_,t_1__213_,t_1__212_,t_1__211_,t_1__210_,t_1__209_,t_1__208_,
  t_1__207_,t_1__206_,t_1__205_,t_1__204_,t_1__203_,t_1__202_,t_1__201_,t_1__200_,
  t_1__199_,t_1__198_,t_1__197_,t_1__196_,t_1__195_,t_1__194_,t_1__193_,t_1__192_,
  t_1__191_,t_1__190_,t_1__189_,t_1__188_,t_1__187_,t_1__186_,t_1__185_,t_1__184_,
  t_1__183_,t_1__182_,t_1__181_,t_1__180_,t_1__179_,t_1__178_,t_1__177_,t_1__176_,
  t_1__175_,t_1__174_,t_1__173_,t_1__172_,t_1__171_,t_1__170_,t_1__169_,t_1__168_,
  t_1__167_,t_1__166_,t_1__165_,t_1__164_,t_1__163_,t_1__162_,t_1__161_,t_1__160_,
  t_1__159_,t_1__158_,t_1__157_,t_1__156_,t_1__155_,t_1__154_,t_1__153_,t_1__152_,
  t_1__151_,t_1__150_,t_1__149_,t_1__148_,t_1__147_,t_1__146_,t_1__145_,t_1__144_,
  t_1__143_,t_1__142_,t_1__141_,t_1__140_,t_1__139_,t_1__138_,t_1__137_,t_1__136_,
  t_1__135_,t_1__134_,t_1__133_,t_1__132_,t_1__131_,t_1__130_,t_1__129_,t_1__128_,
  t_1__127_,t_1__126_,t_1__125_,t_1__124_,t_1__123_,t_1__122_,t_1__121_,t_1__120_,
  t_1__119_,t_1__118_,t_1__117_,t_1__116_,t_1__115_,t_1__114_,t_1__113_,t_1__112_,
  t_1__111_,t_1__110_,t_1__109_,t_1__108_,t_1__107_,t_1__106_,t_1__105_,t_1__104_,
  t_1__103_,t_1__102_,t_1__101_,t_1__100_,t_1__99_,t_1__98_,t_1__97_,t_1__96_,
  t_1__95_,t_1__94_,t_1__93_,t_1__92_,t_1__91_,t_1__90_,t_1__89_,t_1__88_,t_1__87_,
  t_1__86_,t_1__85_,t_1__84_,t_1__83_,t_1__82_,t_1__81_,t_1__80_,t_1__79_,t_1__78_,
  t_1__77_,t_1__76_,t_1__75_,t_1__74_,t_1__73_,t_1__72_,t_1__71_,t_1__70_,t_1__69_,
  t_1__68_,t_1__67_,t_1__66_,t_1__65_,t_1__64_,t_1__63_,t_1__62_,t_1__61_,t_1__60_,
  t_1__59_,t_1__58_,t_1__57_,t_1__56_,t_1__55_,t_1__54_,t_1__53_,t_1__52_,
  t_1__51_,t_1__50_,t_1__49_,t_1__48_,t_1__47_,t_1__46_,t_1__45_,t_1__44_,t_1__43_,
  t_1__42_,t_1__41_,t_1__40_,t_1__39_,t_1__38_,t_1__37_,t_1__36_,t_1__35_,t_1__34_,
  t_1__33_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,t_1__27_,t_1__26_,t_1__25_,
  t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,t_1__18_,t_1__17_,t_1__16_,
  t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,t_1__9_,t_1__8_,t_1__7_,
  t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_,t_2__511_,t_2__510_,t_2__509_,
  t_2__508_,t_2__507_,t_2__506_,t_2__505_,t_2__504_,t_2__503_,t_2__502_,t_2__501_,
  t_2__500_,t_2__499_,t_2__498_,t_2__497_,t_2__496_,t_2__495_,t_2__494_,t_2__493_,
  t_2__492_,t_2__491_,t_2__490_,t_2__489_,t_2__488_,t_2__487_,t_2__486_,t_2__485_,
  t_2__484_,t_2__483_,t_2__482_,t_2__481_,t_2__480_,t_2__479_,t_2__478_,t_2__477_,
  t_2__476_,t_2__475_,t_2__474_,t_2__473_,t_2__472_,t_2__471_,t_2__470_,t_2__469_,
  t_2__468_,t_2__467_,t_2__466_,t_2__465_,t_2__464_,t_2__463_,t_2__462_,t_2__461_,
  t_2__460_,t_2__459_,t_2__458_,t_2__457_,t_2__456_,t_2__455_,t_2__454_,t_2__453_,
  t_2__452_,t_2__451_,t_2__450_,t_2__449_,t_2__448_,t_2__447_,t_2__446_,t_2__445_,
  t_2__444_,t_2__443_,t_2__442_,t_2__441_,t_2__440_,t_2__439_,t_2__438_,t_2__437_,
  t_2__436_,t_2__435_,t_2__434_,t_2__433_,t_2__432_,t_2__431_,t_2__430_,t_2__429_,
  t_2__428_,t_2__427_,t_2__426_,t_2__425_,t_2__424_,t_2__423_,t_2__422_,t_2__421_,
  t_2__420_,t_2__419_,t_2__418_,t_2__417_,t_2__416_,t_2__415_,t_2__414_,t_2__413_,
  t_2__412_,t_2__411_,t_2__410_,t_2__409_,t_2__408_,t_2__407_,t_2__406_,t_2__405_,
  t_2__404_,t_2__403_,t_2__402_,t_2__401_,t_2__400_,t_2__399_,t_2__398_,t_2__397_,
  t_2__396_,t_2__395_,t_2__394_,t_2__393_,t_2__392_,t_2__391_,t_2__390_,t_2__389_,
  t_2__388_,t_2__387_,t_2__386_,t_2__385_,t_2__384_,t_2__383_,t_2__382_,t_2__381_,
  t_2__380_,t_2__379_,t_2__378_,t_2__377_,t_2__376_,t_2__375_,t_2__374_,t_2__373_,
  t_2__372_,t_2__371_,t_2__370_,t_2__369_,t_2__368_,t_2__367_,t_2__366_,t_2__365_,
  t_2__364_,t_2__363_,t_2__362_,t_2__361_,t_2__360_,t_2__359_,t_2__358_,t_2__357_,
  t_2__356_,t_2__355_,t_2__354_,t_2__353_,t_2__352_,t_2__351_,t_2__350_,t_2__349_,
  t_2__348_,t_2__347_,t_2__346_,t_2__345_,t_2__344_,t_2__343_,t_2__342_,t_2__341_,
  t_2__340_,t_2__339_,t_2__338_,t_2__337_,t_2__336_,t_2__335_,t_2__334_,t_2__333_,
  t_2__332_,t_2__331_,t_2__330_,t_2__329_,t_2__328_,t_2__327_,t_2__326_,t_2__325_,
  t_2__324_,t_2__323_,t_2__322_,t_2__321_,t_2__320_,t_2__319_,t_2__318_,t_2__317_,
  t_2__316_,t_2__315_,t_2__314_,t_2__313_,t_2__312_,t_2__311_,t_2__310_,t_2__309_,
  t_2__308_,t_2__307_,t_2__306_,t_2__305_,t_2__304_,t_2__303_,t_2__302_,t_2__301_,
  t_2__300_,t_2__299_,t_2__298_,t_2__297_,t_2__296_,t_2__295_,t_2__294_,t_2__293_,
  t_2__292_,t_2__291_,t_2__290_,t_2__289_,t_2__288_,t_2__287_,t_2__286_,t_2__285_,
  t_2__284_,t_2__283_,t_2__282_,t_2__281_,t_2__280_,t_2__279_,t_2__278_,t_2__277_,
  t_2__276_,t_2__275_,t_2__274_,t_2__273_,t_2__272_,t_2__271_,t_2__270_,t_2__269_,
  t_2__268_,t_2__267_,t_2__266_,t_2__265_,t_2__264_,t_2__263_,t_2__262_,t_2__261_,
  t_2__260_,t_2__259_,t_2__258_,t_2__257_,t_2__256_,t_2__255_,t_2__254_,t_2__253_,
  t_2__252_,t_2__251_,t_2__250_,t_2__249_,t_2__248_,t_2__247_,t_2__246_,t_2__245_,
  t_2__244_,t_2__243_,t_2__242_,t_2__241_,t_2__240_,t_2__239_,t_2__238_,t_2__237_,
  t_2__236_,t_2__235_,t_2__234_,t_2__233_,t_2__232_,t_2__231_,t_2__230_,t_2__229_,
  t_2__228_,t_2__227_,t_2__226_,t_2__225_,t_2__224_,t_2__223_,t_2__222_,t_2__221_,
  t_2__220_,t_2__219_,t_2__218_,t_2__217_,t_2__216_,t_2__215_,t_2__214_,t_2__213_,
  t_2__212_,t_2__211_,t_2__210_,t_2__209_,t_2__208_,t_2__207_,t_2__206_,t_2__205_,
  t_2__204_,t_2__203_,t_2__202_,t_2__201_,t_2__200_,t_2__199_,t_2__198_,t_2__197_,
  t_2__196_,t_2__195_,t_2__194_,t_2__193_,t_2__192_,t_2__191_,t_2__190_,t_2__189_,
  t_2__188_,t_2__187_,t_2__186_,t_2__185_,t_2__184_,t_2__183_,t_2__182_,t_2__181_,
  t_2__180_,t_2__179_,t_2__178_,t_2__177_,t_2__176_,t_2__175_,t_2__174_,t_2__173_,
  t_2__172_,t_2__171_,t_2__170_,t_2__169_,t_2__168_,t_2__167_,t_2__166_,t_2__165_,
  t_2__164_,t_2__163_,t_2__162_,t_2__161_,t_2__160_,t_2__159_,t_2__158_,t_2__157_,
  t_2__156_,t_2__155_,t_2__154_,t_2__153_,t_2__152_,t_2__151_,t_2__150_,t_2__149_,
  t_2__148_,t_2__147_,t_2__146_,t_2__145_,t_2__144_,t_2__143_,t_2__142_,t_2__141_,
  t_2__140_,t_2__139_,t_2__138_,t_2__137_,t_2__136_,t_2__135_,t_2__134_,t_2__133_,
  t_2__132_,t_2__131_,t_2__130_,t_2__129_,t_2__128_,t_2__127_,t_2__126_,t_2__125_,
  t_2__124_,t_2__123_,t_2__122_,t_2__121_,t_2__120_,t_2__119_,t_2__118_,t_2__117_,
  t_2__116_,t_2__115_,t_2__114_,t_2__113_,t_2__112_,t_2__111_,t_2__110_,t_2__109_,
  t_2__108_,t_2__107_,t_2__106_,t_2__105_,t_2__104_,t_2__103_,t_2__102_,t_2__101_,
  t_2__100_,t_2__99_,t_2__98_,t_2__97_,t_2__96_,t_2__95_,t_2__94_,t_2__93_,
  t_2__92_,t_2__91_,t_2__90_,t_2__89_,t_2__88_,t_2__87_,t_2__86_,t_2__85_,t_2__84_,
  t_2__83_,t_2__82_,t_2__81_,t_2__80_,t_2__79_,t_2__78_,t_2__77_,t_2__76_,t_2__75_,
  t_2__74_,t_2__73_,t_2__72_,t_2__71_,t_2__70_,t_2__69_,t_2__68_,t_2__67_,t_2__66_,
  t_2__65_,t_2__64_,t_2__63_,t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,t_2__57_,
  t_2__56_,t_2__55_,t_2__54_,t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,t_2__48_,
  t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,t_2__39_,
  t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,t_2__30_,
  t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,
  t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,
  t_2__2_,t_2__1_,t_2__0_,t_3__511_,t_3__510_,t_3__509_,t_3__508_,t_3__507_,t_3__506_,
  t_3__505_,t_3__504_,t_3__503_,t_3__502_,t_3__501_,t_3__500_,t_3__499_,t_3__498_,
  t_3__497_,t_3__496_,t_3__495_,t_3__494_,t_3__493_,t_3__492_,t_3__491_,t_3__490_,
  t_3__489_,t_3__488_,t_3__487_,t_3__486_,t_3__485_,t_3__484_,t_3__483_,t_3__482_,
  t_3__481_,t_3__480_,t_3__479_,t_3__478_,t_3__477_,t_3__476_,t_3__475_,t_3__474_,
  t_3__473_,t_3__472_,t_3__471_,t_3__470_,t_3__469_,t_3__468_,t_3__467_,t_3__466_,
  t_3__465_,t_3__464_,t_3__463_,t_3__462_,t_3__461_,t_3__460_,t_3__459_,t_3__458_,
  t_3__457_,t_3__456_,t_3__455_,t_3__454_,t_3__453_,t_3__452_,t_3__451_,t_3__450_,
  t_3__449_,t_3__448_,t_3__447_,t_3__446_,t_3__445_,t_3__444_,t_3__443_,t_3__442_,
  t_3__441_,t_3__440_,t_3__439_,t_3__438_,t_3__437_,t_3__436_,t_3__435_,t_3__434_,
  t_3__433_,t_3__432_,t_3__431_,t_3__430_,t_3__429_,t_3__428_,t_3__427_,t_3__426_,
  t_3__425_,t_3__424_,t_3__423_,t_3__422_,t_3__421_,t_3__420_,t_3__419_,t_3__418_,
  t_3__417_,t_3__416_,t_3__415_,t_3__414_,t_3__413_,t_3__412_,t_3__411_,t_3__410_,
  t_3__409_,t_3__408_,t_3__407_,t_3__406_,t_3__405_,t_3__404_,t_3__403_,t_3__402_,
  t_3__401_,t_3__400_,t_3__399_,t_3__398_,t_3__397_,t_3__396_,t_3__395_,t_3__394_,
  t_3__393_,t_3__392_,t_3__391_,t_3__390_,t_3__389_,t_3__388_,t_3__387_,t_3__386_,
  t_3__385_,t_3__384_,t_3__383_,t_3__382_,t_3__381_,t_3__380_,t_3__379_,t_3__378_,
  t_3__377_,t_3__376_,t_3__375_,t_3__374_,t_3__373_,t_3__372_,t_3__371_,t_3__370_,
  t_3__369_,t_3__368_,t_3__367_,t_3__366_,t_3__365_,t_3__364_,t_3__363_,t_3__362_,
  t_3__361_,t_3__360_,t_3__359_,t_3__358_,t_3__357_,t_3__356_,t_3__355_,t_3__354_,
  t_3__353_,t_3__352_,t_3__351_,t_3__350_,t_3__349_,t_3__348_,t_3__347_,t_3__346_,
  t_3__345_,t_3__344_,t_3__343_,t_3__342_,t_3__341_,t_3__340_,t_3__339_,t_3__338_,
  t_3__337_,t_3__336_,t_3__335_,t_3__334_,t_3__333_,t_3__332_,t_3__331_,t_3__330_,
  t_3__329_,t_3__328_,t_3__327_,t_3__326_,t_3__325_,t_3__324_,t_3__323_,t_3__322_,
  t_3__321_,t_3__320_,t_3__319_,t_3__318_,t_3__317_,t_3__316_,t_3__315_,t_3__314_,
  t_3__313_,t_3__312_,t_3__311_,t_3__310_,t_3__309_,t_3__308_,t_3__307_,t_3__306_,
  t_3__305_,t_3__304_,t_3__303_,t_3__302_,t_3__301_,t_3__300_,t_3__299_,t_3__298_,
  t_3__297_,t_3__296_,t_3__295_,t_3__294_,t_3__293_,t_3__292_,t_3__291_,t_3__290_,
  t_3__289_,t_3__288_,t_3__287_,t_3__286_,t_3__285_,t_3__284_,t_3__283_,t_3__282_,
  t_3__281_,t_3__280_,t_3__279_,t_3__278_,t_3__277_,t_3__276_,t_3__275_,t_3__274_,
  t_3__273_,t_3__272_,t_3__271_,t_3__270_,t_3__269_,t_3__268_,t_3__267_,t_3__266_,
  t_3__265_,t_3__264_,t_3__263_,t_3__262_,t_3__261_,t_3__260_,t_3__259_,t_3__258_,
  t_3__257_,t_3__256_,t_3__255_,t_3__254_,t_3__253_,t_3__252_,t_3__251_,t_3__250_,
  t_3__249_,t_3__248_,t_3__247_,t_3__246_,t_3__245_,t_3__244_,t_3__243_,t_3__242_,
  t_3__241_,t_3__240_,t_3__239_,t_3__238_,t_3__237_,t_3__236_,t_3__235_,t_3__234_,
  t_3__233_,t_3__232_,t_3__231_,t_3__230_,t_3__229_,t_3__228_,t_3__227_,t_3__226_,
  t_3__225_,t_3__224_,t_3__223_,t_3__222_,t_3__221_,t_3__220_,t_3__219_,t_3__218_,
  t_3__217_,t_3__216_,t_3__215_,t_3__214_,t_3__213_,t_3__212_,t_3__211_,t_3__210_,
  t_3__209_,t_3__208_,t_3__207_,t_3__206_,t_3__205_,t_3__204_,t_3__203_,t_3__202_,
  t_3__201_,t_3__200_,t_3__199_,t_3__198_,t_3__197_,t_3__196_,t_3__195_,t_3__194_,
  t_3__193_,t_3__192_,t_3__191_,t_3__190_,t_3__189_,t_3__188_,t_3__187_,t_3__186_,
  t_3__185_,t_3__184_,t_3__183_,t_3__182_,t_3__181_,t_3__180_,t_3__179_,t_3__178_,
  t_3__177_,t_3__176_,t_3__175_,t_3__174_,t_3__173_,t_3__172_,t_3__171_,t_3__170_,
  t_3__169_,t_3__168_,t_3__167_,t_3__166_,t_3__165_,t_3__164_,t_3__163_,t_3__162_,
  t_3__161_,t_3__160_,t_3__159_,t_3__158_,t_3__157_,t_3__156_,t_3__155_,t_3__154_,
  t_3__153_,t_3__152_,t_3__151_,t_3__150_,t_3__149_,t_3__148_,t_3__147_,t_3__146_,
  t_3__145_,t_3__144_,t_3__143_,t_3__142_,t_3__141_,t_3__140_,t_3__139_,t_3__138_,
  t_3__137_,t_3__136_,t_3__135_,t_3__134_,t_3__133_,t_3__132_,t_3__131_,t_3__130_,
  t_3__129_,t_3__128_,t_3__127_,t_3__126_,t_3__125_,t_3__124_,t_3__123_,t_3__122_,
  t_3__121_,t_3__120_,t_3__119_,t_3__118_,t_3__117_,t_3__116_,t_3__115_,t_3__114_,
  t_3__113_,t_3__112_,t_3__111_,t_3__110_,t_3__109_,t_3__108_,t_3__107_,t_3__106_,
  t_3__105_,t_3__104_,t_3__103_,t_3__102_,t_3__101_,t_3__100_,t_3__99_,t_3__98_,
  t_3__97_,t_3__96_,t_3__95_,t_3__94_,t_3__93_,t_3__92_,t_3__91_,t_3__90_,t_3__89_,
  t_3__88_,t_3__87_,t_3__86_,t_3__85_,t_3__84_,t_3__83_,t_3__82_,t_3__81_,t_3__80_,
  t_3__79_,t_3__78_,t_3__77_,t_3__76_,t_3__75_,t_3__74_,t_3__73_,t_3__72_,
  t_3__71_,t_3__70_,t_3__69_,t_3__68_,t_3__67_,t_3__66_,t_3__65_,t_3__64_,t_3__63_,
  t_3__62_,t_3__61_,t_3__60_,t_3__59_,t_3__58_,t_3__57_,t_3__56_,t_3__55_,t_3__54_,
  t_3__53_,t_3__52_,t_3__51_,t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,t_3__45_,
  t_3__44_,t_3__43_,t_3__42_,t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,t_3__36_,
  t_3__35_,t_3__34_,t_3__33_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,
  t_3__26_,t_3__25_,t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,
  t_3__17_,t_3__16_,t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,
  t_3__8_,t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_4__511_,
  t_4__510_,t_4__509_,t_4__508_,t_4__507_,t_4__506_,t_4__505_,t_4__504_,t_4__503_,
  t_4__502_,t_4__501_,t_4__500_,t_4__499_,t_4__498_,t_4__497_,t_4__496_,t_4__495_,
  t_4__494_,t_4__493_,t_4__492_,t_4__491_,t_4__490_,t_4__489_,t_4__488_,t_4__487_,
  t_4__486_,t_4__485_,t_4__484_,t_4__483_,t_4__482_,t_4__481_,t_4__480_,t_4__479_,
  t_4__478_,t_4__477_,t_4__476_,t_4__475_,t_4__474_,t_4__473_,t_4__472_,t_4__471_,
  t_4__470_,t_4__469_,t_4__468_,t_4__467_,t_4__466_,t_4__465_,t_4__464_,t_4__463_,
  t_4__462_,t_4__461_,t_4__460_,t_4__459_,t_4__458_,t_4__457_,t_4__456_,t_4__455_,
  t_4__454_,t_4__453_,t_4__452_,t_4__451_,t_4__450_,t_4__449_,t_4__448_,t_4__447_,
  t_4__446_,t_4__445_,t_4__444_,t_4__443_,t_4__442_,t_4__441_,t_4__440_,t_4__439_,
  t_4__438_,t_4__437_,t_4__436_,t_4__435_,t_4__434_,t_4__433_,t_4__432_,t_4__431_,
  t_4__430_,t_4__429_,t_4__428_,t_4__427_,t_4__426_,t_4__425_,t_4__424_,t_4__423_,
  t_4__422_,t_4__421_,t_4__420_,t_4__419_,t_4__418_,t_4__417_,t_4__416_,t_4__415_,
  t_4__414_,t_4__413_,t_4__412_,t_4__411_,t_4__410_,t_4__409_,t_4__408_,t_4__407_,
  t_4__406_,t_4__405_,t_4__404_,t_4__403_,t_4__402_,t_4__401_,t_4__400_,t_4__399_,
  t_4__398_,t_4__397_,t_4__396_,t_4__395_,t_4__394_,t_4__393_,t_4__392_,t_4__391_,
  t_4__390_,t_4__389_,t_4__388_,t_4__387_,t_4__386_,t_4__385_,t_4__384_,t_4__383_,
  t_4__382_,t_4__381_,t_4__380_,t_4__379_,t_4__378_,t_4__377_,t_4__376_,t_4__375_,
  t_4__374_,t_4__373_,t_4__372_,t_4__371_,t_4__370_,t_4__369_,t_4__368_,t_4__367_,
  t_4__366_,t_4__365_,t_4__364_,t_4__363_,t_4__362_,t_4__361_,t_4__360_,t_4__359_,
  t_4__358_,t_4__357_,t_4__356_,t_4__355_,t_4__354_,t_4__353_,t_4__352_,t_4__351_,
  t_4__350_,t_4__349_,t_4__348_,t_4__347_,t_4__346_,t_4__345_,t_4__344_,t_4__343_,
  t_4__342_,t_4__341_,t_4__340_,t_4__339_,t_4__338_,t_4__337_,t_4__336_,t_4__335_,
  t_4__334_,t_4__333_,t_4__332_,t_4__331_,t_4__330_,t_4__329_,t_4__328_,t_4__327_,
  t_4__326_,t_4__325_,t_4__324_,t_4__323_,t_4__322_,t_4__321_,t_4__320_,t_4__319_,
  t_4__318_,t_4__317_,t_4__316_,t_4__315_,t_4__314_,t_4__313_,t_4__312_,t_4__311_,
  t_4__310_,t_4__309_,t_4__308_,t_4__307_,t_4__306_,t_4__305_,t_4__304_,t_4__303_,
  t_4__302_,t_4__301_,t_4__300_,t_4__299_,t_4__298_,t_4__297_,t_4__296_,t_4__295_,
  t_4__294_,t_4__293_,t_4__292_,t_4__291_,t_4__290_,t_4__289_,t_4__288_,t_4__287_,
  t_4__286_,t_4__285_,t_4__284_,t_4__283_,t_4__282_,t_4__281_,t_4__280_,t_4__279_,
  t_4__278_,t_4__277_,t_4__276_,t_4__275_,t_4__274_,t_4__273_,t_4__272_,t_4__271_,
  t_4__270_,t_4__269_,t_4__268_,t_4__267_,t_4__266_,t_4__265_,t_4__264_,t_4__263_,
  t_4__262_,t_4__261_,t_4__260_,t_4__259_,t_4__258_,t_4__257_,t_4__256_,t_4__255_,
  t_4__254_,t_4__253_,t_4__252_,t_4__251_,t_4__250_,t_4__249_,t_4__248_,t_4__247_,
  t_4__246_,t_4__245_,t_4__244_,t_4__243_,t_4__242_,t_4__241_,t_4__240_,t_4__239_,
  t_4__238_,t_4__237_,t_4__236_,t_4__235_,t_4__234_,t_4__233_,t_4__232_,t_4__231_,
  t_4__230_,t_4__229_,t_4__228_,t_4__227_,t_4__226_,t_4__225_,t_4__224_,t_4__223_,
  t_4__222_,t_4__221_,t_4__220_,t_4__219_,t_4__218_,t_4__217_,t_4__216_,t_4__215_,
  t_4__214_,t_4__213_,t_4__212_,t_4__211_,t_4__210_,t_4__209_,t_4__208_,t_4__207_,
  t_4__206_,t_4__205_,t_4__204_,t_4__203_,t_4__202_,t_4__201_,t_4__200_,t_4__199_,
  t_4__198_,t_4__197_,t_4__196_,t_4__195_,t_4__194_,t_4__193_,t_4__192_,t_4__191_,
  t_4__190_,t_4__189_,t_4__188_,t_4__187_,t_4__186_,t_4__185_,t_4__184_,t_4__183_,
  t_4__182_,t_4__181_,t_4__180_,t_4__179_,t_4__178_,t_4__177_,t_4__176_,t_4__175_,
  t_4__174_,t_4__173_,t_4__172_,t_4__171_,t_4__170_,t_4__169_,t_4__168_,t_4__167_,
  t_4__166_,t_4__165_,t_4__164_,t_4__163_,t_4__162_,t_4__161_,t_4__160_,t_4__159_,
  t_4__158_,t_4__157_,t_4__156_,t_4__155_,t_4__154_,t_4__153_,t_4__152_,t_4__151_,
  t_4__150_,t_4__149_,t_4__148_,t_4__147_,t_4__146_,t_4__145_,t_4__144_,t_4__143_,
  t_4__142_,t_4__141_,t_4__140_,t_4__139_,t_4__138_,t_4__137_,t_4__136_,t_4__135_,
  t_4__134_,t_4__133_,t_4__132_,t_4__131_,t_4__130_,t_4__129_,t_4__128_,t_4__127_,
  t_4__126_,t_4__125_,t_4__124_,t_4__123_,t_4__122_,t_4__121_,t_4__120_,t_4__119_,
  t_4__118_,t_4__117_,t_4__116_,t_4__115_,t_4__114_,t_4__113_,t_4__112_,t_4__111_,
  t_4__110_,t_4__109_,t_4__108_,t_4__107_,t_4__106_,t_4__105_,t_4__104_,t_4__103_,
  t_4__102_,t_4__101_,t_4__100_,t_4__99_,t_4__98_,t_4__97_,t_4__96_,t_4__95_,
  t_4__94_,t_4__93_,t_4__92_,t_4__91_,t_4__90_,t_4__89_,t_4__88_,t_4__87_,t_4__86_,
  t_4__85_,t_4__84_,t_4__83_,t_4__82_,t_4__81_,t_4__80_,t_4__79_,t_4__78_,t_4__77_,
  t_4__76_,t_4__75_,t_4__74_,t_4__73_,t_4__72_,t_4__71_,t_4__70_,t_4__69_,t_4__68_,
  t_4__67_,t_4__66_,t_4__65_,t_4__64_,t_4__63_,t_4__62_,t_4__61_,t_4__60_,t_4__59_,
  t_4__58_,t_4__57_,t_4__56_,t_4__55_,t_4__54_,t_4__53_,t_4__52_,t_4__51_,t_4__50_,
  t_4__49_,t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,t_4__43_,t_4__42_,
  t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,t_4__34_,t_4__33_,
  t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,t_4__25_,t_4__24_,
  t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,t_4__16_,t_4__15_,
  t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,t_4__7_,t_4__6_,t_4__5_,
  t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_,t_5__511_,t_5__510_,t_5__509_,t_5__508_,
  t_5__507_,t_5__506_,t_5__505_,t_5__504_,t_5__503_,t_5__502_,t_5__501_,t_5__500_,
  t_5__499_,t_5__498_,t_5__497_,t_5__496_,t_5__495_,t_5__494_,t_5__493_,t_5__492_,
  t_5__491_,t_5__490_,t_5__489_,t_5__488_,t_5__487_,t_5__486_,t_5__485_,t_5__484_,
  t_5__483_,t_5__482_,t_5__481_,t_5__480_,t_5__479_,t_5__478_,t_5__477_,t_5__476_,
  t_5__475_,t_5__474_,t_5__473_,t_5__472_,t_5__471_,t_5__470_,t_5__469_,t_5__468_,
  t_5__467_,t_5__466_,t_5__465_,t_5__464_,t_5__463_,t_5__462_,t_5__461_,t_5__460_,
  t_5__459_,t_5__458_,t_5__457_,t_5__456_,t_5__455_,t_5__454_,t_5__453_,t_5__452_,
  t_5__451_,t_5__450_,t_5__449_,t_5__448_,t_5__447_,t_5__446_,t_5__445_,t_5__444_,
  t_5__443_,t_5__442_,t_5__441_,t_5__440_,t_5__439_,t_5__438_,t_5__437_,t_5__436_,
  t_5__435_,t_5__434_,t_5__433_,t_5__432_,t_5__431_,t_5__430_,t_5__429_,t_5__428_,
  t_5__427_,t_5__426_,t_5__425_,t_5__424_,t_5__423_,t_5__422_,t_5__421_,t_5__420_,
  t_5__419_,t_5__418_,t_5__417_,t_5__416_,t_5__415_,t_5__414_,t_5__413_,t_5__412_,
  t_5__411_,t_5__410_,t_5__409_,t_5__408_,t_5__407_,t_5__406_,t_5__405_,t_5__404_,
  t_5__403_,t_5__402_,t_5__401_,t_5__400_,t_5__399_,t_5__398_,t_5__397_,t_5__396_,
  t_5__395_,t_5__394_,t_5__393_,t_5__392_,t_5__391_,t_5__390_,t_5__389_,t_5__388_,
  t_5__387_,t_5__386_,t_5__385_,t_5__384_,t_5__383_,t_5__382_,t_5__381_,t_5__380_,
  t_5__379_,t_5__378_,t_5__377_,t_5__376_,t_5__375_,t_5__374_,t_5__373_,t_5__372_,
  t_5__371_,t_5__370_,t_5__369_,t_5__368_,t_5__367_,t_5__366_,t_5__365_,t_5__364_,
  t_5__363_,t_5__362_,t_5__361_,t_5__360_,t_5__359_,t_5__358_,t_5__357_,t_5__356_,
  t_5__355_,t_5__354_,t_5__353_,t_5__352_,t_5__351_,t_5__350_,t_5__349_,t_5__348_,
  t_5__347_,t_5__346_,t_5__345_,t_5__344_,t_5__343_,t_5__342_,t_5__341_,t_5__340_,
  t_5__339_,t_5__338_,t_5__337_,t_5__336_,t_5__335_,t_5__334_,t_5__333_,t_5__332_,
  t_5__331_,t_5__330_,t_5__329_,t_5__328_,t_5__327_,t_5__326_,t_5__325_,t_5__324_,
  t_5__323_,t_5__322_,t_5__321_,t_5__320_,t_5__319_,t_5__318_,t_5__317_,t_5__316_,
  t_5__315_,t_5__314_,t_5__313_,t_5__312_,t_5__311_,t_5__310_,t_5__309_,t_5__308_,
  t_5__307_,t_5__306_,t_5__305_,t_5__304_,t_5__303_,t_5__302_,t_5__301_,t_5__300_,
  t_5__299_,t_5__298_,t_5__297_,t_5__296_,t_5__295_,t_5__294_,t_5__293_,t_5__292_,
  t_5__291_,t_5__290_,t_5__289_,t_5__288_,t_5__287_,t_5__286_,t_5__285_,t_5__284_,
  t_5__283_,t_5__282_,t_5__281_,t_5__280_,t_5__279_,t_5__278_,t_5__277_,t_5__276_,
  t_5__275_,t_5__274_,t_5__273_,t_5__272_,t_5__271_,t_5__270_,t_5__269_,t_5__268_,
  t_5__267_,t_5__266_,t_5__265_,t_5__264_,t_5__263_,t_5__262_,t_5__261_,t_5__260_,
  t_5__259_,t_5__258_,t_5__257_,t_5__256_,t_5__255_,t_5__254_,t_5__253_,t_5__252_,
  t_5__251_,t_5__250_,t_5__249_,t_5__248_,t_5__247_,t_5__246_,t_5__245_,t_5__244_,
  t_5__243_,t_5__242_,t_5__241_,t_5__240_,t_5__239_,t_5__238_,t_5__237_,t_5__236_,
  t_5__235_,t_5__234_,t_5__233_,t_5__232_,t_5__231_,t_5__230_,t_5__229_,t_5__228_,
  t_5__227_,t_5__226_,t_5__225_,t_5__224_,t_5__223_,t_5__222_,t_5__221_,t_5__220_,
  t_5__219_,t_5__218_,t_5__217_,t_5__216_,t_5__215_,t_5__214_,t_5__213_,t_5__212_,
  t_5__211_,t_5__210_,t_5__209_,t_5__208_,t_5__207_,t_5__206_,t_5__205_,t_5__204_,
  t_5__203_,t_5__202_,t_5__201_,t_5__200_,t_5__199_,t_5__198_,t_5__197_,t_5__196_,
  t_5__195_,t_5__194_,t_5__193_,t_5__192_,t_5__191_,t_5__190_,t_5__189_,t_5__188_,
  t_5__187_,t_5__186_,t_5__185_,t_5__184_,t_5__183_,t_5__182_,t_5__181_,t_5__180_,
  t_5__179_,t_5__178_,t_5__177_,t_5__176_,t_5__175_,t_5__174_,t_5__173_,t_5__172_,
  t_5__171_,t_5__170_,t_5__169_,t_5__168_,t_5__167_,t_5__166_,t_5__165_,t_5__164_,
  t_5__163_,t_5__162_,t_5__161_,t_5__160_,t_5__159_,t_5__158_,t_5__157_,t_5__156_,
  t_5__155_,t_5__154_,t_5__153_,t_5__152_,t_5__151_,t_5__150_,t_5__149_,t_5__148_,
  t_5__147_,t_5__146_,t_5__145_,t_5__144_,t_5__143_,t_5__142_,t_5__141_,t_5__140_,
  t_5__139_,t_5__138_,t_5__137_,t_5__136_,t_5__135_,t_5__134_,t_5__133_,t_5__132_,
  t_5__131_,t_5__130_,t_5__129_,t_5__128_,t_5__127_,t_5__126_,t_5__125_,t_5__124_,
  t_5__123_,t_5__122_,t_5__121_,t_5__120_,t_5__119_,t_5__118_,t_5__117_,t_5__116_,
  t_5__115_,t_5__114_,t_5__113_,t_5__112_,t_5__111_,t_5__110_,t_5__109_,t_5__108_,
  t_5__107_,t_5__106_,t_5__105_,t_5__104_,t_5__103_,t_5__102_,t_5__101_,t_5__100_,
  t_5__99_,t_5__98_,t_5__97_,t_5__96_,t_5__95_,t_5__94_,t_5__93_,t_5__92_,
  t_5__91_,t_5__90_,t_5__89_,t_5__88_,t_5__87_,t_5__86_,t_5__85_,t_5__84_,t_5__83_,
  t_5__82_,t_5__81_,t_5__80_,t_5__79_,t_5__78_,t_5__77_,t_5__76_,t_5__75_,t_5__74_,
  t_5__73_,t_5__72_,t_5__71_,t_5__70_,t_5__69_,t_5__68_,t_5__67_,t_5__66_,t_5__65_,
  t_5__64_,t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,t_5__58_,t_5__57_,t_5__56_,
  t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,
  t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,
  t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,
  t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,
  t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,
  t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,
  t_5__1_,t_5__0_,t_6__511_,t_6__510_,t_6__509_,t_6__508_,t_6__507_,t_6__506_,t_6__505_,
  t_6__504_,t_6__503_,t_6__502_,t_6__501_,t_6__500_,t_6__499_,t_6__498_,t_6__497_,
  t_6__496_,t_6__495_,t_6__494_,t_6__493_,t_6__492_,t_6__491_,t_6__490_,t_6__489_,
  t_6__488_,t_6__487_,t_6__486_,t_6__485_,t_6__484_,t_6__483_,t_6__482_,t_6__481_,
  t_6__480_,t_6__479_,t_6__478_,t_6__477_,t_6__476_,t_6__475_,t_6__474_,t_6__473_,
  t_6__472_,t_6__471_,t_6__470_,t_6__469_,t_6__468_,t_6__467_,t_6__466_,t_6__465_,
  t_6__464_,t_6__463_,t_6__462_,t_6__461_,t_6__460_,t_6__459_,t_6__458_,t_6__457_,
  t_6__456_,t_6__455_,t_6__454_,t_6__453_,t_6__452_,t_6__451_,t_6__450_,t_6__449_,
  t_6__448_,t_6__447_,t_6__446_,t_6__445_,t_6__444_,t_6__443_,t_6__442_,t_6__441_,
  t_6__440_,t_6__439_,t_6__438_,t_6__437_,t_6__436_,t_6__435_,t_6__434_,t_6__433_,
  t_6__432_,t_6__431_,t_6__430_,t_6__429_,t_6__428_,t_6__427_,t_6__426_,t_6__425_,
  t_6__424_,t_6__423_,t_6__422_,t_6__421_,t_6__420_,t_6__419_,t_6__418_,t_6__417_,
  t_6__416_,t_6__415_,t_6__414_,t_6__413_,t_6__412_,t_6__411_,t_6__410_,t_6__409_,
  t_6__408_,t_6__407_,t_6__406_,t_6__405_,t_6__404_,t_6__403_,t_6__402_,t_6__401_,
  t_6__400_,t_6__399_,t_6__398_,t_6__397_,t_6__396_,t_6__395_,t_6__394_,t_6__393_,
  t_6__392_,t_6__391_,t_6__390_,t_6__389_,t_6__388_,t_6__387_,t_6__386_,t_6__385_,
  t_6__384_,t_6__383_,t_6__382_,t_6__381_,t_6__380_,t_6__379_,t_6__378_,t_6__377_,
  t_6__376_,t_6__375_,t_6__374_,t_6__373_,t_6__372_,t_6__371_,t_6__370_,t_6__369_,
  t_6__368_,t_6__367_,t_6__366_,t_6__365_,t_6__364_,t_6__363_,t_6__362_,t_6__361_,
  t_6__360_,t_6__359_,t_6__358_,t_6__357_,t_6__356_,t_6__355_,t_6__354_,t_6__353_,
  t_6__352_,t_6__351_,t_6__350_,t_6__349_,t_6__348_,t_6__347_,t_6__346_,t_6__345_,
  t_6__344_,t_6__343_,t_6__342_,t_6__341_,t_6__340_,t_6__339_,t_6__338_,t_6__337_,
  t_6__336_,t_6__335_,t_6__334_,t_6__333_,t_6__332_,t_6__331_,t_6__330_,t_6__329_,
  t_6__328_,t_6__327_,t_6__326_,t_6__325_,t_6__324_,t_6__323_,t_6__322_,t_6__321_,
  t_6__320_,t_6__319_,t_6__318_,t_6__317_,t_6__316_,t_6__315_,t_6__314_,t_6__313_,
  t_6__312_,t_6__311_,t_6__310_,t_6__309_,t_6__308_,t_6__307_,t_6__306_,t_6__305_,
  t_6__304_,t_6__303_,t_6__302_,t_6__301_,t_6__300_,t_6__299_,t_6__298_,t_6__297_,
  t_6__296_,t_6__295_,t_6__294_,t_6__293_,t_6__292_,t_6__291_,t_6__290_,t_6__289_,
  t_6__288_,t_6__287_,t_6__286_,t_6__285_,t_6__284_,t_6__283_,t_6__282_,t_6__281_,
  t_6__280_,t_6__279_,t_6__278_,t_6__277_,t_6__276_,t_6__275_,t_6__274_,t_6__273_,
  t_6__272_,t_6__271_,t_6__270_,t_6__269_,t_6__268_,t_6__267_,t_6__266_,t_6__265_,
  t_6__264_,t_6__263_,t_6__262_,t_6__261_,t_6__260_,t_6__259_,t_6__258_,t_6__257_,
  t_6__256_,t_6__255_,t_6__254_,t_6__253_,t_6__252_,t_6__251_,t_6__250_,t_6__249_,
  t_6__248_,t_6__247_,t_6__246_,t_6__245_,t_6__244_,t_6__243_,t_6__242_,t_6__241_,
  t_6__240_,t_6__239_,t_6__238_,t_6__237_,t_6__236_,t_6__235_,t_6__234_,t_6__233_,
  t_6__232_,t_6__231_,t_6__230_,t_6__229_,t_6__228_,t_6__227_,t_6__226_,t_6__225_,
  t_6__224_,t_6__223_,t_6__222_,t_6__221_,t_6__220_,t_6__219_,t_6__218_,t_6__217_,
  t_6__216_,t_6__215_,t_6__214_,t_6__213_,t_6__212_,t_6__211_,t_6__210_,t_6__209_,
  t_6__208_,t_6__207_,t_6__206_,t_6__205_,t_6__204_,t_6__203_,t_6__202_,t_6__201_,
  t_6__200_,t_6__199_,t_6__198_,t_6__197_,t_6__196_,t_6__195_,t_6__194_,t_6__193_,
  t_6__192_,t_6__191_,t_6__190_,t_6__189_,t_6__188_,t_6__187_,t_6__186_,t_6__185_,
  t_6__184_,t_6__183_,t_6__182_,t_6__181_,t_6__180_,t_6__179_,t_6__178_,t_6__177_,
  t_6__176_,t_6__175_,t_6__174_,t_6__173_,t_6__172_,t_6__171_,t_6__170_,t_6__169_,
  t_6__168_,t_6__167_,t_6__166_,t_6__165_,t_6__164_,t_6__163_,t_6__162_,t_6__161_,
  t_6__160_,t_6__159_,t_6__158_,t_6__157_,t_6__156_,t_6__155_,t_6__154_,t_6__153_,
  t_6__152_,t_6__151_,t_6__150_,t_6__149_,t_6__148_,t_6__147_,t_6__146_,t_6__145_,
  t_6__144_,t_6__143_,t_6__142_,t_6__141_,t_6__140_,t_6__139_,t_6__138_,t_6__137_,
  t_6__136_,t_6__135_,t_6__134_,t_6__133_,t_6__132_,t_6__131_,t_6__130_,t_6__129_,
  t_6__128_,t_6__127_,t_6__126_,t_6__125_,t_6__124_,t_6__123_,t_6__122_,t_6__121_,
  t_6__120_,t_6__119_,t_6__118_,t_6__117_,t_6__116_,t_6__115_,t_6__114_,t_6__113_,
  t_6__112_,t_6__111_,t_6__110_,t_6__109_,t_6__108_,t_6__107_,t_6__106_,t_6__105_,
  t_6__104_,t_6__103_,t_6__102_,t_6__101_,t_6__100_,t_6__99_,t_6__98_,t_6__97_,
  t_6__96_,t_6__95_,t_6__94_,t_6__93_,t_6__92_,t_6__91_,t_6__90_,t_6__89_,t_6__88_,
  t_6__87_,t_6__86_,t_6__85_,t_6__84_,t_6__83_,t_6__82_,t_6__81_,t_6__80_,t_6__79_,
  t_6__78_,t_6__77_,t_6__76_,t_6__75_,t_6__74_,t_6__73_,t_6__72_,t_6__71_,t_6__70_,
  t_6__69_,t_6__68_,t_6__67_,t_6__66_,t_6__65_,t_6__64_,t_6__63_,t_6__62_,
  t_6__61_,t_6__60_,t_6__59_,t_6__58_,t_6__57_,t_6__56_,t_6__55_,t_6__54_,t_6__53_,
  t_6__52_,t_6__51_,t_6__50_,t_6__49_,t_6__48_,t_6__47_,t_6__46_,t_6__45_,t_6__44_,
  t_6__43_,t_6__42_,t_6__41_,t_6__40_,t_6__39_,t_6__38_,t_6__37_,t_6__36_,t_6__35_,
  t_6__34_,t_6__33_,t_6__32_,t_6__31_,t_6__30_,t_6__29_,t_6__28_,t_6__27_,t_6__26_,
  t_6__25_,t_6__24_,t_6__23_,t_6__22_,t_6__21_,t_6__20_,t_6__19_,t_6__18_,t_6__17_,
  t_6__16_,t_6__15_,t_6__14_,t_6__13_,t_6__12_,t_6__11_,t_6__10_,t_6__9_,t_6__8_,
  t_6__7_,t_6__6_,t_6__5_,t_6__4_,t_6__3_,t_6__2_,t_6__1_,t_6__0_,t_7__511_,t_7__510_,
  t_7__509_,t_7__508_,t_7__507_,t_7__506_,t_7__505_,t_7__504_,t_7__503_,t_7__502_,
  t_7__501_,t_7__500_,t_7__499_,t_7__498_,t_7__497_,t_7__496_,t_7__495_,t_7__494_,
  t_7__493_,t_7__492_,t_7__491_,t_7__490_,t_7__489_,t_7__488_,t_7__487_,t_7__486_,
  t_7__485_,t_7__484_,t_7__483_,t_7__482_,t_7__481_,t_7__480_,t_7__479_,t_7__478_,
  t_7__477_,t_7__476_,t_7__475_,t_7__474_,t_7__473_,t_7__472_,t_7__471_,t_7__470_,
  t_7__469_,t_7__468_,t_7__467_,t_7__466_,t_7__465_,t_7__464_,t_7__463_,t_7__462_,
  t_7__461_,t_7__460_,t_7__459_,t_7__458_,t_7__457_,t_7__456_,t_7__455_,t_7__454_,
  t_7__453_,t_7__452_,t_7__451_,t_7__450_,t_7__449_,t_7__448_,t_7__447_,t_7__446_,
  t_7__445_,t_7__444_,t_7__443_,t_7__442_,t_7__441_,t_7__440_,t_7__439_,t_7__438_,
  t_7__437_,t_7__436_,t_7__435_,t_7__434_,t_7__433_,t_7__432_,t_7__431_,t_7__430_,
  t_7__429_,t_7__428_,t_7__427_,t_7__426_,t_7__425_,t_7__424_,t_7__423_,t_7__422_,
  t_7__421_,t_7__420_,t_7__419_,t_7__418_,t_7__417_,t_7__416_,t_7__415_,t_7__414_,
  t_7__413_,t_7__412_,t_7__411_,t_7__410_,t_7__409_,t_7__408_,t_7__407_,t_7__406_,
  t_7__405_,t_7__404_,t_7__403_,t_7__402_,t_7__401_,t_7__400_,t_7__399_,t_7__398_,
  t_7__397_,t_7__396_,t_7__395_,t_7__394_,t_7__393_,t_7__392_,t_7__391_,t_7__390_,
  t_7__389_,t_7__388_,t_7__387_,t_7__386_,t_7__385_,t_7__384_,t_7__383_,t_7__382_,
  t_7__381_,t_7__380_,t_7__379_,t_7__378_,t_7__377_,t_7__376_,t_7__375_,t_7__374_,
  t_7__373_,t_7__372_,t_7__371_,t_7__370_,t_7__369_,t_7__368_,t_7__367_,t_7__366_,
  t_7__365_,t_7__364_,t_7__363_,t_7__362_,t_7__361_,t_7__360_,t_7__359_,t_7__358_,
  t_7__357_,t_7__356_,t_7__355_,t_7__354_,t_7__353_,t_7__352_,t_7__351_,t_7__350_,
  t_7__349_,t_7__348_,t_7__347_,t_7__346_,t_7__345_,t_7__344_,t_7__343_,t_7__342_,
  t_7__341_,t_7__340_,t_7__339_,t_7__338_,t_7__337_,t_7__336_,t_7__335_,t_7__334_,
  t_7__333_,t_7__332_,t_7__331_,t_7__330_,t_7__329_,t_7__328_,t_7__327_,t_7__326_,
  t_7__325_,t_7__324_,t_7__323_,t_7__322_,t_7__321_,t_7__320_,t_7__319_,t_7__318_,
  t_7__317_,t_7__316_,t_7__315_,t_7__314_,t_7__313_,t_7__312_,t_7__311_,t_7__310_,
  t_7__309_,t_7__308_,t_7__307_,t_7__306_,t_7__305_,t_7__304_,t_7__303_,t_7__302_,
  t_7__301_,t_7__300_,t_7__299_,t_7__298_,t_7__297_,t_7__296_,t_7__295_,t_7__294_,
  t_7__293_,t_7__292_,t_7__291_,t_7__290_,t_7__289_,t_7__288_,t_7__287_,t_7__286_,
  t_7__285_,t_7__284_,t_7__283_,t_7__282_,t_7__281_,t_7__280_,t_7__279_,t_7__278_,
  t_7__277_,t_7__276_,t_7__275_,t_7__274_,t_7__273_,t_7__272_,t_7__271_,t_7__270_,
  t_7__269_,t_7__268_,t_7__267_,t_7__266_,t_7__265_,t_7__264_,t_7__263_,t_7__262_,
  t_7__261_,t_7__260_,t_7__259_,t_7__258_,t_7__257_,t_7__256_,t_7__255_,t_7__254_,
  t_7__253_,t_7__252_,t_7__251_,t_7__250_,t_7__249_,t_7__248_,t_7__247_,t_7__246_,
  t_7__245_,t_7__244_,t_7__243_,t_7__242_,t_7__241_,t_7__240_,t_7__239_,t_7__238_,
  t_7__237_,t_7__236_,t_7__235_,t_7__234_,t_7__233_,t_7__232_,t_7__231_,t_7__230_,
  t_7__229_,t_7__228_,t_7__227_,t_7__226_,t_7__225_,t_7__224_,t_7__223_,t_7__222_,
  t_7__221_,t_7__220_,t_7__219_,t_7__218_,t_7__217_,t_7__216_,t_7__215_,t_7__214_,
  t_7__213_,t_7__212_,t_7__211_,t_7__210_,t_7__209_,t_7__208_,t_7__207_,t_7__206_,
  t_7__205_,t_7__204_,t_7__203_,t_7__202_,t_7__201_,t_7__200_,t_7__199_,t_7__198_,
  t_7__197_,t_7__196_,t_7__195_,t_7__194_,t_7__193_,t_7__192_,t_7__191_,t_7__190_,
  t_7__189_,t_7__188_,t_7__187_,t_7__186_,t_7__185_,t_7__184_,t_7__183_,t_7__182_,
  t_7__181_,t_7__180_,t_7__179_,t_7__178_,t_7__177_,t_7__176_,t_7__175_,t_7__174_,
  t_7__173_,t_7__172_,t_7__171_,t_7__170_,t_7__169_,t_7__168_,t_7__167_,t_7__166_,
  t_7__165_,t_7__164_,t_7__163_,t_7__162_,t_7__161_,t_7__160_,t_7__159_,t_7__158_,
  t_7__157_,t_7__156_,t_7__155_,t_7__154_,t_7__153_,t_7__152_,t_7__151_,t_7__150_,
  t_7__149_,t_7__148_,t_7__147_,t_7__146_,t_7__145_,t_7__144_,t_7__143_,t_7__142_,
  t_7__141_,t_7__140_,t_7__139_,t_7__138_,t_7__137_,t_7__136_,t_7__135_,t_7__134_,
  t_7__133_,t_7__132_,t_7__131_,t_7__130_,t_7__129_,t_7__128_,t_7__127_,t_7__126_,
  t_7__125_,t_7__124_,t_7__123_,t_7__122_,t_7__121_,t_7__120_,t_7__119_,t_7__118_,
  t_7__117_,t_7__116_,t_7__115_,t_7__114_,t_7__113_,t_7__112_,t_7__111_,t_7__110_,
  t_7__109_,t_7__108_,t_7__107_,t_7__106_,t_7__105_,t_7__104_,t_7__103_,t_7__102_,
  t_7__101_,t_7__100_,t_7__99_,t_7__98_,t_7__97_,t_7__96_,t_7__95_,t_7__94_,
  t_7__93_,t_7__92_,t_7__91_,t_7__90_,t_7__89_,t_7__88_,t_7__87_,t_7__86_,t_7__85_,
  t_7__84_,t_7__83_,t_7__82_,t_7__81_,t_7__80_,t_7__79_,t_7__78_,t_7__77_,t_7__76_,
  t_7__75_,t_7__74_,t_7__73_,t_7__72_,t_7__71_,t_7__70_,t_7__69_,t_7__68_,t_7__67_,
  t_7__66_,t_7__65_,t_7__64_,t_7__63_,t_7__62_,t_7__61_,t_7__60_,t_7__59_,t_7__58_,
  t_7__57_,t_7__56_,t_7__55_,t_7__54_,t_7__53_,t_7__52_,t_7__51_,t_7__50_,t_7__49_,
  t_7__48_,t_7__47_,t_7__46_,t_7__45_,t_7__44_,t_7__43_,t_7__42_,t_7__41_,t_7__40_,
  t_7__39_,t_7__38_,t_7__37_,t_7__36_,t_7__35_,t_7__34_,t_7__33_,t_7__32_,
  t_7__31_,t_7__30_,t_7__29_,t_7__28_,t_7__27_,t_7__26_,t_7__25_,t_7__24_,t_7__23_,
  t_7__22_,t_7__21_,t_7__20_,t_7__19_,t_7__18_,t_7__17_,t_7__16_,t_7__15_,t_7__14_,
  t_7__13_,t_7__12_,t_7__11_,t_7__10_,t_7__9_,t_7__8_,t_7__7_,t_7__6_,t_7__5_,t_7__4_,
  t_7__3_,t_7__2_,t_7__1_,t_7__0_,t_8__511_,t_8__510_,t_8__509_,t_8__508_,t_8__507_,
  t_8__506_,t_8__505_,t_8__504_,t_8__503_,t_8__502_,t_8__501_,t_8__500_,t_8__499_,
  t_8__498_,t_8__497_,t_8__496_,t_8__495_,t_8__494_,t_8__493_,t_8__492_,t_8__491_,
  t_8__490_,t_8__489_,t_8__488_,t_8__487_,t_8__486_,t_8__485_,t_8__484_,t_8__483_,
  t_8__482_,t_8__481_,t_8__480_,t_8__479_,t_8__478_,t_8__477_,t_8__476_,t_8__475_,
  t_8__474_,t_8__473_,t_8__472_,t_8__471_,t_8__470_,t_8__469_,t_8__468_,t_8__467_,
  t_8__466_,t_8__465_,t_8__464_,t_8__463_,t_8__462_,t_8__461_,t_8__460_,t_8__459_,
  t_8__458_,t_8__457_,t_8__456_,t_8__455_,t_8__454_,t_8__453_,t_8__452_,t_8__451_,
  t_8__450_,t_8__449_,t_8__448_,t_8__447_,t_8__446_,t_8__445_,t_8__444_,t_8__443_,
  t_8__442_,t_8__441_,t_8__440_,t_8__439_,t_8__438_,t_8__437_,t_8__436_,t_8__435_,
  t_8__434_,t_8__433_,t_8__432_,t_8__431_,t_8__430_,t_8__429_,t_8__428_,t_8__427_,
  t_8__426_,t_8__425_,t_8__424_,t_8__423_,t_8__422_,t_8__421_,t_8__420_,t_8__419_,
  t_8__418_,t_8__417_,t_8__416_,t_8__415_,t_8__414_,t_8__413_,t_8__412_,t_8__411_,
  t_8__410_,t_8__409_,t_8__408_,t_8__407_,t_8__406_,t_8__405_,t_8__404_,t_8__403_,
  t_8__402_,t_8__401_,t_8__400_,t_8__399_,t_8__398_,t_8__397_,t_8__396_,t_8__395_,
  t_8__394_,t_8__393_,t_8__392_,t_8__391_,t_8__390_,t_8__389_,t_8__388_,t_8__387_,
  t_8__386_,t_8__385_,t_8__384_,t_8__383_,t_8__382_,t_8__381_,t_8__380_,t_8__379_,
  t_8__378_,t_8__377_,t_8__376_,t_8__375_,t_8__374_,t_8__373_,t_8__372_,t_8__371_,
  t_8__370_,t_8__369_,t_8__368_,t_8__367_,t_8__366_,t_8__365_,t_8__364_,t_8__363_,
  t_8__362_,t_8__361_,t_8__360_,t_8__359_,t_8__358_,t_8__357_,t_8__356_,t_8__355_,
  t_8__354_,t_8__353_,t_8__352_,t_8__351_,t_8__350_,t_8__349_,t_8__348_,t_8__347_,
  t_8__346_,t_8__345_,t_8__344_,t_8__343_,t_8__342_,t_8__341_,t_8__340_,t_8__339_,
  t_8__338_,t_8__337_,t_8__336_,t_8__335_,t_8__334_,t_8__333_,t_8__332_,t_8__331_,
  t_8__330_,t_8__329_,t_8__328_,t_8__327_,t_8__326_,t_8__325_,t_8__324_,t_8__323_,
  t_8__322_,t_8__321_,t_8__320_,t_8__319_,t_8__318_,t_8__317_,t_8__316_,t_8__315_,
  t_8__314_,t_8__313_,t_8__312_,t_8__311_,t_8__310_,t_8__309_,t_8__308_,t_8__307_,
  t_8__306_,t_8__305_,t_8__304_,t_8__303_,t_8__302_,t_8__301_,t_8__300_,t_8__299_,
  t_8__298_,t_8__297_,t_8__296_,t_8__295_,t_8__294_,t_8__293_,t_8__292_,t_8__291_,
  t_8__290_,t_8__289_,t_8__288_,t_8__287_,t_8__286_,t_8__285_,t_8__284_,t_8__283_,
  t_8__282_,t_8__281_,t_8__280_,t_8__279_,t_8__278_,t_8__277_,t_8__276_,t_8__275_,
  t_8__274_,t_8__273_,t_8__272_,t_8__271_,t_8__270_,t_8__269_,t_8__268_,t_8__267_,
  t_8__266_,t_8__265_,t_8__264_,t_8__263_,t_8__262_,t_8__261_,t_8__260_,t_8__259_,
  t_8__258_,t_8__257_,t_8__256_,t_8__255_,t_8__254_,t_8__253_,t_8__252_,t_8__251_,
  t_8__250_,t_8__249_,t_8__248_,t_8__247_,t_8__246_,t_8__245_,t_8__244_,t_8__243_,
  t_8__242_,t_8__241_,t_8__240_,t_8__239_,t_8__238_,t_8__237_,t_8__236_,t_8__235_,
  t_8__234_,t_8__233_,t_8__232_,t_8__231_,t_8__230_,t_8__229_,t_8__228_,t_8__227_,
  t_8__226_,t_8__225_,t_8__224_,t_8__223_,t_8__222_,t_8__221_,t_8__220_,t_8__219_,
  t_8__218_,t_8__217_,t_8__216_,t_8__215_,t_8__214_,t_8__213_,t_8__212_,t_8__211_,
  t_8__210_,t_8__209_,t_8__208_,t_8__207_,t_8__206_,t_8__205_,t_8__204_,t_8__203_,
  t_8__202_,t_8__201_,t_8__200_,t_8__199_,t_8__198_,t_8__197_,t_8__196_,t_8__195_,
  t_8__194_,t_8__193_,t_8__192_,t_8__191_,t_8__190_,t_8__189_,t_8__188_,t_8__187_,
  t_8__186_,t_8__185_,t_8__184_,t_8__183_,t_8__182_,t_8__181_,t_8__180_,t_8__179_,
  t_8__178_,t_8__177_,t_8__176_,t_8__175_,t_8__174_,t_8__173_,t_8__172_,t_8__171_,
  t_8__170_,t_8__169_,t_8__168_,t_8__167_,t_8__166_,t_8__165_,t_8__164_,t_8__163_,
  t_8__162_,t_8__161_,t_8__160_,t_8__159_,t_8__158_,t_8__157_,t_8__156_,t_8__155_,
  t_8__154_,t_8__153_,t_8__152_,t_8__151_,t_8__150_,t_8__149_,t_8__148_,t_8__147_,
  t_8__146_,t_8__145_,t_8__144_,t_8__143_,t_8__142_,t_8__141_,t_8__140_,t_8__139_,
  t_8__138_,t_8__137_,t_8__136_,t_8__135_,t_8__134_,t_8__133_,t_8__132_,t_8__131_,
  t_8__130_,t_8__129_,t_8__128_,t_8__127_,t_8__126_,t_8__125_,t_8__124_,t_8__123_,
  t_8__122_,t_8__121_,t_8__120_,t_8__119_,t_8__118_,t_8__117_,t_8__116_,t_8__115_,
  t_8__114_,t_8__113_,t_8__112_,t_8__111_,t_8__110_,t_8__109_,t_8__108_,t_8__107_,
  t_8__106_,t_8__105_,t_8__104_,t_8__103_,t_8__102_,t_8__101_,t_8__100_,t_8__99_,
  t_8__98_,t_8__97_,t_8__96_,t_8__95_,t_8__94_,t_8__93_,t_8__92_,t_8__91_,t_8__90_,
  t_8__89_,t_8__88_,t_8__87_,t_8__86_,t_8__85_,t_8__84_,t_8__83_,t_8__82_,
  t_8__81_,t_8__80_,t_8__79_,t_8__78_,t_8__77_,t_8__76_,t_8__75_,t_8__74_,t_8__73_,
  t_8__72_,t_8__71_,t_8__70_,t_8__69_,t_8__68_,t_8__67_,t_8__66_,t_8__65_,t_8__64_,
  t_8__63_,t_8__62_,t_8__61_,t_8__60_,t_8__59_,t_8__58_,t_8__57_,t_8__56_,t_8__55_,
  t_8__54_,t_8__53_,t_8__52_,t_8__51_,t_8__50_,t_8__49_,t_8__48_,t_8__47_,t_8__46_,
  t_8__45_,t_8__44_,t_8__43_,t_8__42_,t_8__41_,t_8__40_,t_8__39_,t_8__38_,t_8__37_,
  t_8__36_,t_8__35_,t_8__34_,t_8__33_,t_8__32_,t_8__31_,t_8__30_,t_8__29_,t_8__28_,
  t_8__27_,t_8__26_,t_8__25_,t_8__24_,t_8__23_,t_8__22_,t_8__21_,t_8__20_,t_8__19_,
  t_8__18_,t_8__17_,t_8__16_,t_8__15_,t_8__14_,t_8__13_,t_8__12_,t_8__11_,t_8__10_,
  t_8__9_,t_8__8_,t_8__7_,t_8__6_,t_8__5_,t_8__4_,t_8__3_,t_8__2_,t_8__1_,t_8__0_;
  assign t_1__511_ = i[0] | 1'b0;
  assign t_1__510_ = i[1] | i[0];
  assign t_1__509_ = i[2] | i[1];
  assign t_1__508_ = i[3] | i[2];
  assign t_1__507_ = i[4] | i[3];
  assign t_1__506_ = i[5] | i[4];
  assign t_1__505_ = i[6] | i[5];
  assign t_1__504_ = i[7] | i[6];
  assign t_1__503_ = i[8] | i[7];
  assign t_1__502_ = i[9] | i[8];
  assign t_1__501_ = i[10] | i[9];
  assign t_1__500_ = i[11] | i[10];
  assign t_1__499_ = i[12] | i[11];
  assign t_1__498_ = i[13] | i[12];
  assign t_1__497_ = i[14] | i[13];
  assign t_1__496_ = i[15] | i[14];
  assign t_1__495_ = i[16] | i[15];
  assign t_1__494_ = i[17] | i[16];
  assign t_1__493_ = i[18] | i[17];
  assign t_1__492_ = i[19] | i[18];
  assign t_1__491_ = i[20] | i[19];
  assign t_1__490_ = i[21] | i[20];
  assign t_1__489_ = i[22] | i[21];
  assign t_1__488_ = i[23] | i[22];
  assign t_1__487_ = i[24] | i[23];
  assign t_1__486_ = i[25] | i[24];
  assign t_1__485_ = i[26] | i[25];
  assign t_1__484_ = i[27] | i[26];
  assign t_1__483_ = i[28] | i[27];
  assign t_1__482_ = i[29] | i[28];
  assign t_1__481_ = i[30] | i[29];
  assign t_1__480_ = i[31] | i[30];
  assign t_1__479_ = i[32] | i[31];
  assign t_1__478_ = i[33] | i[32];
  assign t_1__477_ = i[34] | i[33];
  assign t_1__476_ = i[35] | i[34];
  assign t_1__475_ = i[36] | i[35];
  assign t_1__474_ = i[37] | i[36];
  assign t_1__473_ = i[38] | i[37];
  assign t_1__472_ = i[39] | i[38];
  assign t_1__471_ = i[40] | i[39];
  assign t_1__470_ = i[41] | i[40];
  assign t_1__469_ = i[42] | i[41];
  assign t_1__468_ = i[43] | i[42];
  assign t_1__467_ = i[44] | i[43];
  assign t_1__466_ = i[45] | i[44];
  assign t_1__465_ = i[46] | i[45];
  assign t_1__464_ = i[47] | i[46];
  assign t_1__463_ = i[48] | i[47];
  assign t_1__462_ = i[49] | i[48];
  assign t_1__461_ = i[50] | i[49];
  assign t_1__460_ = i[51] | i[50];
  assign t_1__459_ = i[52] | i[51];
  assign t_1__458_ = i[53] | i[52];
  assign t_1__457_ = i[54] | i[53];
  assign t_1__456_ = i[55] | i[54];
  assign t_1__455_ = i[56] | i[55];
  assign t_1__454_ = i[57] | i[56];
  assign t_1__453_ = i[58] | i[57];
  assign t_1__452_ = i[59] | i[58];
  assign t_1__451_ = i[60] | i[59];
  assign t_1__450_ = i[61] | i[60];
  assign t_1__449_ = i[62] | i[61];
  assign t_1__448_ = i[63] | i[62];
  assign t_1__447_ = i[64] | i[63];
  assign t_1__446_ = i[65] | i[64];
  assign t_1__445_ = i[66] | i[65];
  assign t_1__444_ = i[67] | i[66];
  assign t_1__443_ = i[68] | i[67];
  assign t_1__442_ = i[69] | i[68];
  assign t_1__441_ = i[70] | i[69];
  assign t_1__440_ = i[71] | i[70];
  assign t_1__439_ = i[72] | i[71];
  assign t_1__438_ = i[73] | i[72];
  assign t_1__437_ = i[74] | i[73];
  assign t_1__436_ = i[75] | i[74];
  assign t_1__435_ = i[76] | i[75];
  assign t_1__434_ = i[77] | i[76];
  assign t_1__433_ = i[78] | i[77];
  assign t_1__432_ = i[79] | i[78];
  assign t_1__431_ = i[80] | i[79];
  assign t_1__430_ = i[81] | i[80];
  assign t_1__429_ = i[82] | i[81];
  assign t_1__428_ = i[83] | i[82];
  assign t_1__427_ = i[84] | i[83];
  assign t_1__426_ = i[85] | i[84];
  assign t_1__425_ = i[86] | i[85];
  assign t_1__424_ = i[87] | i[86];
  assign t_1__423_ = i[88] | i[87];
  assign t_1__422_ = i[89] | i[88];
  assign t_1__421_ = i[90] | i[89];
  assign t_1__420_ = i[91] | i[90];
  assign t_1__419_ = i[92] | i[91];
  assign t_1__418_ = i[93] | i[92];
  assign t_1__417_ = i[94] | i[93];
  assign t_1__416_ = i[95] | i[94];
  assign t_1__415_ = i[96] | i[95];
  assign t_1__414_ = i[97] | i[96];
  assign t_1__413_ = i[98] | i[97];
  assign t_1__412_ = i[99] | i[98];
  assign t_1__411_ = i[100] | i[99];
  assign t_1__410_ = i[101] | i[100];
  assign t_1__409_ = i[102] | i[101];
  assign t_1__408_ = i[103] | i[102];
  assign t_1__407_ = i[104] | i[103];
  assign t_1__406_ = i[105] | i[104];
  assign t_1__405_ = i[106] | i[105];
  assign t_1__404_ = i[107] | i[106];
  assign t_1__403_ = i[108] | i[107];
  assign t_1__402_ = i[109] | i[108];
  assign t_1__401_ = i[110] | i[109];
  assign t_1__400_ = i[111] | i[110];
  assign t_1__399_ = i[112] | i[111];
  assign t_1__398_ = i[113] | i[112];
  assign t_1__397_ = i[114] | i[113];
  assign t_1__396_ = i[115] | i[114];
  assign t_1__395_ = i[116] | i[115];
  assign t_1__394_ = i[117] | i[116];
  assign t_1__393_ = i[118] | i[117];
  assign t_1__392_ = i[119] | i[118];
  assign t_1__391_ = i[120] | i[119];
  assign t_1__390_ = i[121] | i[120];
  assign t_1__389_ = i[122] | i[121];
  assign t_1__388_ = i[123] | i[122];
  assign t_1__387_ = i[124] | i[123];
  assign t_1__386_ = i[125] | i[124];
  assign t_1__385_ = i[126] | i[125];
  assign t_1__384_ = i[127] | i[126];
  assign t_1__383_ = i[128] | i[127];
  assign t_1__382_ = i[129] | i[128];
  assign t_1__381_ = i[130] | i[129];
  assign t_1__380_ = i[131] | i[130];
  assign t_1__379_ = i[132] | i[131];
  assign t_1__378_ = i[133] | i[132];
  assign t_1__377_ = i[134] | i[133];
  assign t_1__376_ = i[135] | i[134];
  assign t_1__375_ = i[136] | i[135];
  assign t_1__374_ = i[137] | i[136];
  assign t_1__373_ = i[138] | i[137];
  assign t_1__372_ = i[139] | i[138];
  assign t_1__371_ = i[140] | i[139];
  assign t_1__370_ = i[141] | i[140];
  assign t_1__369_ = i[142] | i[141];
  assign t_1__368_ = i[143] | i[142];
  assign t_1__367_ = i[144] | i[143];
  assign t_1__366_ = i[145] | i[144];
  assign t_1__365_ = i[146] | i[145];
  assign t_1__364_ = i[147] | i[146];
  assign t_1__363_ = i[148] | i[147];
  assign t_1__362_ = i[149] | i[148];
  assign t_1__361_ = i[150] | i[149];
  assign t_1__360_ = i[151] | i[150];
  assign t_1__359_ = i[152] | i[151];
  assign t_1__358_ = i[153] | i[152];
  assign t_1__357_ = i[154] | i[153];
  assign t_1__356_ = i[155] | i[154];
  assign t_1__355_ = i[156] | i[155];
  assign t_1__354_ = i[157] | i[156];
  assign t_1__353_ = i[158] | i[157];
  assign t_1__352_ = i[159] | i[158];
  assign t_1__351_ = i[160] | i[159];
  assign t_1__350_ = i[161] | i[160];
  assign t_1__349_ = i[162] | i[161];
  assign t_1__348_ = i[163] | i[162];
  assign t_1__347_ = i[164] | i[163];
  assign t_1__346_ = i[165] | i[164];
  assign t_1__345_ = i[166] | i[165];
  assign t_1__344_ = i[167] | i[166];
  assign t_1__343_ = i[168] | i[167];
  assign t_1__342_ = i[169] | i[168];
  assign t_1__341_ = i[170] | i[169];
  assign t_1__340_ = i[171] | i[170];
  assign t_1__339_ = i[172] | i[171];
  assign t_1__338_ = i[173] | i[172];
  assign t_1__337_ = i[174] | i[173];
  assign t_1__336_ = i[175] | i[174];
  assign t_1__335_ = i[176] | i[175];
  assign t_1__334_ = i[177] | i[176];
  assign t_1__333_ = i[178] | i[177];
  assign t_1__332_ = i[179] | i[178];
  assign t_1__331_ = i[180] | i[179];
  assign t_1__330_ = i[181] | i[180];
  assign t_1__329_ = i[182] | i[181];
  assign t_1__328_ = i[183] | i[182];
  assign t_1__327_ = i[184] | i[183];
  assign t_1__326_ = i[185] | i[184];
  assign t_1__325_ = i[186] | i[185];
  assign t_1__324_ = i[187] | i[186];
  assign t_1__323_ = i[188] | i[187];
  assign t_1__322_ = i[189] | i[188];
  assign t_1__321_ = i[190] | i[189];
  assign t_1__320_ = i[191] | i[190];
  assign t_1__319_ = i[192] | i[191];
  assign t_1__318_ = i[193] | i[192];
  assign t_1__317_ = i[194] | i[193];
  assign t_1__316_ = i[195] | i[194];
  assign t_1__315_ = i[196] | i[195];
  assign t_1__314_ = i[197] | i[196];
  assign t_1__313_ = i[198] | i[197];
  assign t_1__312_ = i[199] | i[198];
  assign t_1__311_ = i[200] | i[199];
  assign t_1__310_ = i[201] | i[200];
  assign t_1__309_ = i[202] | i[201];
  assign t_1__308_ = i[203] | i[202];
  assign t_1__307_ = i[204] | i[203];
  assign t_1__306_ = i[205] | i[204];
  assign t_1__305_ = i[206] | i[205];
  assign t_1__304_ = i[207] | i[206];
  assign t_1__303_ = i[208] | i[207];
  assign t_1__302_ = i[209] | i[208];
  assign t_1__301_ = i[210] | i[209];
  assign t_1__300_ = i[211] | i[210];
  assign t_1__299_ = i[212] | i[211];
  assign t_1__298_ = i[213] | i[212];
  assign t_1__297_ = i[214] | i[213];
  assign t_1__296_ = i[215] | i[214];
  assign t_1__295_ = i[216] | i[215];
  assign t_1__294_ = i[217] | i[216];
  assign t_1__293_ = i[218] | i[217];
  assign t_1__292_ = i[219] | i[218];
  assign t_1__291_ = i[220] | i[219];
  assign t_1__290_ = i[221] | i[220];
  assign t_1__289_ = i[222] | i[221];
  assign t_1__288_ = i[223] | i[222];
  assign t_1__287_ = i[224] | i[223];
  assign t_1__286_ = i[225] | i[224];
  assign t_1__285_ = i[226] | i[225];
  assign t_1__284_ = i[227] | i[226];
  assign t_1__283_ = i[228] | i[227];
  assign t_1__282_ = i[229] | i[228];
  assign t_1__281_ = i[230] | i[229];
  assign t_1__280_ = i[231] | i[230];
  assign t_1__279_ = i[232] | i[231];
  assign t_1__278_ = i[233] | i[232];
  assign t_1__277_ = i[234] | i[233];
  assign t_1__276_ = i[235] | i[234];
  assign t_1__275_ = i[236] | i[235];
  assign t_1__274_ = i[237] | i[236];
  assign t_1__273_ = i[238] | i[237];
  assign t_1__272_ = i[239] | i[238];
  assign t_1__271_ = i[240] | i[239];
  assign t_1__270_ = i[241] | i[240];
  assign t_1__269_ = i[242] | i[241];
  assign t_1__268_ = i[243] | i[242];
  assign t_1__267_ = i[244] | i[243];
  assign t_1__266_ = i[245] | i[244];
  assign t_1__265_ = i[246] | i[245];
  assign t_1__264_ = i[247] | i[246];
  assign t_1__263_ = i[248] | i[247];
  assign t_1__262_ = i[249] | i[248];
  assign t_1__261_ = i[250] | i[249];
  assign t_1__260_ = i[251] | i[250];
  assign t_1__259_ = i[252] | i[251];
  assign t_1__258_ = i[253] | i[252];
  assign t_1__257_ = i[254] | i[253];
  assign t_1__256_ = i[255] | i[254];
  assign t_1__255_ = i[256] | i[255];
  assign t_1__254_ = i[257] | i[256];
  assign t_1__253_ = i[258] | i[257];
  assign t_1__252_ = i[259] | i[258];
  assign t_1__251_ = i[260] | i[259];
  assign t_1__250_ = i[261] | i[260];
  assign t_1__249_ = i[262] | i[261];
  assign t_1__248_ = i[263] | i[262];
  assign t_1__247_ = i[264] | i[263];
  assign t_1__246_ = i[265] | i[264];
  assign t_1__245_ = i[266] | i[265];
  assign t_1__244_ = i[267] | i[266];
  assign t_1__243_ = i[268] | i[267];
  assign t_1__242_ = i[269] | i[268];
  assign t_1__241_ = i[270] | i[269];
  assign t_1__240_ = i[271] | i[270];
  assign t_1__239_ = i[272] | i[271];
  assign t_1__238_ = i[273] | i[272];
  assign t_1__237_ = i[274] | i[273];
  assign t_1__236_ = i[275] | i[274];
  assign t_1__235_ = i[276] | i[275];
  assign t_1__234_ = i[277] | i[276];
  assign t_1__233_ = i[278] | i[277];
  assign t_1__232_ = i[279] | i[278];
  assign t_1__231_ = i[280] | i[279];
  assign t_1__230_ = i[281] | i[280];
  assign t_1__229_ = i[282] | i[281];
  assign t_1__228_ = i[283] | i[282];
  assign t_1__227_ = i[284] | i[283];
  assign t_1__226_ = i[285] | i[284];
  assign t_1__225_ = i[286] | i[285];
  assign t_1__224_ = i[287] | i[286];
  assign t_1__223_ = i[288] | i[287];
  assign t_1__222_ = i[289] | i[288];
  assign t_1__221_ = i[290] | i[289];
  assign t_1__220_ = i[291] | i[290];
  assign t_1__219_ = i[292] | i[291];
  assign t_1__218_ = i[293] | i[292];
  assign t_1__217_ = i[294] | i[293];
  assign t_1__216_ = i[295] | i[294];
  assign t_1__215_ = i[296] | i[295];
  assign t_1__214_ = i[297] | i[296];
  assign t_1__213_ = i[298] | i[297];
  assign t_1__212_ = i[299] | i[298];
  assign t_1__211_ = i[300] | i[299];
  assign t_1__210_ = i[301] | i[300];
  assign t_1__209_ = i[302] | i[301];
  assign t_1__208_ = i[303] | i[302];
  assign t_1__207_ = i[304] | i[303];
  assign t_1__206_ = i[305] | i[304];
  assign t_1__205_ = i[306] | i[305];
  assign t_1__204_ = i[307] | i[306];
  assign t_1__203_ = i[308] | i[307];
  assign t_1__202_ = i[309] | i[308];
  assign t_1__201_ = i[310] | i[309];
  assign t_1__200_ = i[311] | i[310];
  assign t_1__199_ = i[312] | i[311];
  assign t_1__198_ = i[313] | i[312];
  assign t_1__197_ = i[314] | i[313];
  assign t_1__196_ = i[315] | i[314];
  assign t_1__195_ = i[316] | i[315];
  assign t_1__194_ = i[317] | i[316];
  assign t_1__193_ = i[318] | i[317];
  assign t_1__192_ = i[319] | i[318];
  assign t_1__191_ = i[320] | i[319];
  assign t_1__190_ = i[321] | i[320];
  assign t_1__189_ = i[322] | i[321];
  assign t_1__188_ = i[323] | i[322];
  assign t_1__187_ = i[324] | i[323];
  assign t_1__186_ = i[325] | i[324];
  assign t_1__185_ = i[326] | i[325];
  assign t_1__184_ = i[327] | i[326];
  assign t_1__183_ = i[328] | i[327];
  assign t_1__182_ = i[329] | i[328];
  assign t_1__181_ = i[330] | i[329];
  assign t_1__180_ = i[331] | i[330];
  assign t_1__179_ = i[332] | i[331];
  assign t_1__178_ = i[333] | i[332];
  assign t_1__177_ = i[334] | i[333];
  assign t_1__176_ = i[335] | i[334];
  assign t_1__175_ = i[336] | i[335];
  assign t_1__174_ = i[337] | i[336];
  assign t_1__173_ = i[338] | i[337];
  assign t_1__172_ = i[339] | i[338];
  assign t_1__171_ = i[340] | i[339];
  assign t_1__170_ = i[341] | i[340];
  assign t_1__169_ = i[342] | i[341];
  assign t_1__168_ = i[343] | i[342];
  assign t_1__167_ = i[344] | i[343];
  assign t_1__166_ = i[345] | i[344];
  assign t_1__165_ = i[346] | i[345];
  assign t_1__164_ = i[347] | i[346];
  assign t_1__163_ = i[348] | i[347];
  assign t_1__162_ = i[349] | i[348];
  assign t_1__161_ = i[350] | i[349];
  assign t_1__160_ = i[351] | i[350];
  assign t_1__159_ = i[352] | i[351];
  assign t_1__158_ = i[353] | i[352];
  assign t_1__157_ = i[354] | i[353];
  assign t_1__156_ = i[355] | i[354];
  assign t_1__155_ = i[356] | i[355];
  assign t_1__154_ = i[357] | i[356];
  assign t_1__153_ = i[358] | i[357];
  assign t_1__152_ = i[359] | i[358];
  assign t_1__151_ = i[360] | i[359];
  assign t_1__150_ = i[361] | i[360];
  assign t_1__149_ = i[362] | i[361];
  assign t_1__148_ = i[363] | i[362];
  assign t_1__147_ = i[364] | i[363];
  assign t_1__146_ = i[365] | i[364];
  assign t_1__145_ = i[366] | i[365];
  assign t_1__144_ = i[367] | i[366];
  assign t_1__143_ = i[368] | i[367];
  assign t_1__142_ = i[369] | i[368];
  assign t_1__141_ = i[370] | i[369];
  assign t_1__140_ = i[371] | i[370];
  assign t_1__139_ = i[372] | i[371];
  assign t_1__138_ = i[373] | i[372];
  assign t_1__137_ = i[374] | i[373];
  assign t_1__136_ = i[375] | i[374];
  assign t_1__135_ = i[376] | i[375];
  assign t_1__134_ = i[377] | i[376];
  assign t_1__133_ = i[378] | i[377];
  assign t_1__132_ = i[379] | i[378];
  assign t_1__131_ = i[380] | i[379];
  assign t_1__130_ = i[381] | i[380];
  assign t_1__129_ = i[382] | i[381];
  assign t_1__128_ = i[383] | i[382];
  assign t_1__127_ = i[384] | i[383];
  assign t_1__126_ = i[385] | i[384];
  assign t_1__125_ = i[386] | i[385];
  assign t_1__124_ = i[387] | i[386];
  assign t_1__123_ = i[388] | i[387];
  assign t_1__122_ = i[389] | i[388];
  assign t_1__121_ = i[390] | i[389];
  assign t_1__120_ = i[391] | i[390];
  assign t_1__119_ = i[392] | i[391];
  assign t_1__118_ = i[393] | i[392];
  assign t_1__117_ = i[394] | i[393];
  assign t_1__116_ = i[395] | i[394];
  assign t_1__115_ = i[396] | i[395];
  assign t_1__114_ = i[397] | i[396];
  assign t_1__113_ = i[398] | i[397];
  assign t_1__112_ = i[399] | i[398];
  assign t_1__111_ = i[400] | i[399];
  assign t_1__110_ = i[401] | i[400];
  assign t_1__109_ = i[402] | i[401];
  assign t_1__108_ = i[403] | i[402];
  assign t_1__107_ = i[404] | i[403];
  assign t_1__106_ = i[405] | i[404];
  assign t_1__105_ = i[406] | i[405];
  assign t_1__104_ = i[407] | i[406];
  assign t_1__103_ = i[408] | i[407];
  assign t_1__102_ = i[409] | i[408];
  assign t_1__101_ = i[410] | i[409];
  assign t_1__100_ = i[411] | i[410];
  assign t_1__99_ = i[412] | i[411];
  assign t_1__98_ = i[413] | i[412];
  assign t_1__97_ = i[414] | i[413];
  assign t_1__96_ = i[415] | i[414];
  assign t_1__95_ = i[416] | i[415];
  assign t_1__94_ = i[417] | i[416];
  assign t_1__93_ = i[418] | i[417];
  assign t_1__92_ = i[419] | i[418];
  assign t_1__91_ = i[420] | i[419];
  assign t_1__90_ = i[421] | i[420];
  assign t_1__89_ = i[422] | i[421];
  assign t_1__88_ = i[423] | i[422];
  assign t_1__87_ = i[424] | i[423];
  assign t_1__86_ = i[425] | i[424];
  assign t_1__85_ = i[426] | i[425];
  assign t_1__84_ = i[427] | i[426];
  assign t_1__83_ = i[428] | i[427];
  assign t_1__82_ = i[429] | i[428];
  assign t_1__81_ = i[430] | i[429];
  assign t_1__80_ = i[431] | i[430];
  assign t_1__79_ = i[432] | i[431];
  assign t_1__78_ = i[433] | i[432];
  assign t_1__77_ = i[434] | i[433];
  assign t_1__76_ = i[435] | i[434];
  assign t_1__75_ = i[436] | i[435];
  assign t_1__74_ = i[437] | i[436];
  assign t_1__73_ = i[438] | i[437];
  assign t_1__72_ = i[439] | i[438];
  assign t_1__71_ = i[440] | i[439];
  assign t_1__70_ = i[441] | i[440];
  assign t_1__69_ = i[442] | i[441];
  assign t_1__68_ = i[443] | i[442];
  assign t_1__67_ = i[444] | i[443];
  assign t_1__66_ = i[445] | i[444];
  assign t_1__65_ = i[446] | i[445];
  assign t_1__64_ = i[447] | i[446];
  assign t_1__63_ = i[448] | i[447];
  assign t_1__62_ = i[449] | i[448];
  assign t_1__61_ = i[450] | i[449];
  assign t_1__60_ = i[451] | i[450];
  assign t_1__59_ = i[452] | i[451];
  assign t_1__58_ = i[453] | i[452];
  assign t_1__57_ = i[454] | i[453];
  assign t_1__56_ = i[455] | i[454];
  assign t_1__55_ = i[456] | i[455];
  assign t_1__54_ = i[457] | i[456];
  assign t_1__53_ = i[458] | i[457];
  assign t_1__52_ = i[459] | i[458];
  assign t_1__51_ = i[460] | i[459];
  assign t_1__50_ = i[461] | i[460];
  assign t_1__49_ = i[462] | i[461];
  assign t_1__48_ = i[463] | i[462];
  assign t_1__47_ = i[464] | i[463];
  assign t_1__46_ = i[465] | i[464];
  assign t_1__45_ = i[466] | i[465];
  assign t_1__44_ = i[467] | i[466];
  assign t_1__43_ = i[468] | i[467];
  assign t_1__42_ = i[469] | i[468];
  assign t_1__41_ = i[470] | i[469];
  assign t_1__40_ = i[471] | i[470];
  assign t_1__39_ = i[472] | i[471];
  assign t_1__38_ = i[473] | i[472];
  assign t_1__37_ = i[474] | i[473];
  assign t_1__36_ = i[475] | i[474];
  assign t_1__35_ = i[476] | i[475];
  assign t_1__34_ = i[477] | i[476];
  assign t_1__33_ = i[478] | i[477];
  assign t_1__32_ = i[479] | i[478];
  assign t_1__31_ = i[480] | i[479];
  assign t_1__30_ = i[481] | i[480];
  assign t_1__29_ = i[482] | i[481];
  assign t_1__28_ = i[483] | i[482];
  assign t_1__27_ = i[484] | i[483];
  assign t_1__26_ = i[485] | i[484];
  assign t_1__25_ = i[486] | i[485];
  assign t_1__24_ = i[487] | i[486];
  assign t_1__23_ = i[488] | i[487];
  assign t_1__22_ = i[489] | i[488];
  assign t_1__21_ = i[490] | i[489];
  assign t_1__20_ = i[491] | i[490];
  assign t_1__19_ = i[492] | i[491];
  assign t_1__18_ = i[493] | i[492];
  assign t_1__17_ = i[494] | i[493];
  assign t_1__16_ = i[495] | i[494];
  assign t_1__15_ = i[496] | i[495];
  assign t_1__14_ = i[497] | i[496];
  assign t_1__13_ = i[498] | i[497];
  assign t_1__12_ = i[499] | i[498];
  assign t_1__11_ = i[500] | i[499];
  assign t_1__10_ = i[501] | i[500];
  assign t_1__9_ = i[502] | i[501];
  assign t_1__8_ = i[503] | i[502];
  assign t_1__7_ = i[504] | i[503];
  assign t_1__6_ = i[505] | i[504];
  assign t_1__5_ = i[506] | i[505];
  assign t_1__4_ = i[507] | i[506];
  assign t_1__3_ = i[508] | i[507];
  assign t_1__2_ = i[509] | i[508];
  assign t_1__1_ = i[510] | i[509];
  assign t_1__0_ = i[511] | i[510];
  assign t_2__511_ = t_1__511_ | 1'b0;
  assign t_2__510_ = t_1__510_ | 1'b0;
  assign t_2__509_ = t_1__509_ | t_1__511_;
  assign t_2__508_ = t_1__508_ | t_1__510_;
  assign t_2__507_ = t_1__507_ | t_1__509_;
  assign t_2__506_ = t_1__506_ | t_1__508_;
  assign t_2__505_ = t_1__505_ | t_1__507_;
  assign t_2__504_ = t_1__504_ | t_1__506_;
  assign t_2__503_ = t_1__503_ | t_1__505_;
  assign t_2__502_ = t_1__502_ | t_1__504_;
  assign t_2__501_ = t_1__501_ | t_1__503_;
  assign t_2__500_ = t_1__500_ | t_1__502_;
  assign t_2__499_ = t_1__499_ | t_1__501_;
  assign t_2__498_ = t_1__498_ | t_1__500_;
  assign t_2__497_ = t_1__497_ | t_1__499_;
  assign t_2__496_ = t_1__496_ | t_1__498_;
  assign t_2__495_ = t_1__495_ | t_1__497_;
  assign t_2__494_ = t_1__494_ | t_1__496_;
  assign t_2__493_ = t_1__493_ | t_1__495_;
  assign t_2__492_ = t_1__492_ | t_1__494_;
  assign t_2__491_ = t_1__491_ | t_1__493_;
  assign t_2__490_ = t_1__490_ | t_1__492_;
  assign t_2__489_ = t_1__489_ | t_1__491_;
  assign t_2__488_ = t_1__488_ | t_1__490_;
  assign t_2__487_ = t_1__487_ | t_1__489_;
  assign t_2__486_ = t_1__486_ | t_1__488_;
  assign t_2__485_ = t_1__485_ | t_1__487_;
  assign t_2__484_ = t_1__484_ | t_1__486_;
  assign t_2__483_ = t_1__483_ | t_1__485_;
  assign t_2__482_ = t_1__482_ | t_1__484_;
  assign t_2__481_ = t_1__481_ | t_1__483_;
  assign t_2__480_ = t_1__480_ | t_1__482_;
  assign t_2__479_ = t_1__479_ | t_1__481_;
  assign t_2__478_ = t_1__478_ | t_1__480_;
  assign t_2__477_ = t_1__477_ | t_1__479_;
  assign t_2__476_ = t_1__476_ | t_1__478_;
  assign t_2__475_ = t_1__475_ | t_1__477_;
  assign t_2__474_ = t_1__474_ | t_1__476_;
  assign t_2__473_ = t_1__473_ | t_1__475_;
  assign t_2__472_ = t_1__472_ | t_1__474_;
  assign t_2__471_ = t_1__471_ | t_1__473_;
  assign t_2__470_ = t_1__470_ | t_1__472_;
  assign t_2__469_ = t_1__469_ | t_1__471_;
  assign t_2__468_ = t_1__468_ | t_1__470_;
  assign t_2__467_ = t_1__467_ | t_1__469_;
  assign t_2__466_ = t_1__466_ | t_1__468_;
  assign t_2__465_ = t_1__465_ | t_1__467_;
  assign t_2__464_ = t_1__464_ | t_1__466_;
  assign t_2__463_ = t_1__463_ | t_1__465_;
  assign t_2__462_ = t_1__462_ | t_1__464_;
  assign t_2__461_ = t_1__461_ | t_1__463_;
  assign t_2__460_ = t_1__460_ | t_1__462_;
  assign t_2__459_ = t_1__459_ | t_1__461_;
  assign t_2__458_ = t_1__458_ | t_1__460_;
  assign t_2__457_ = t_1__457_ | t_1__459_;
  assign t_2__456_ = t_1__456_ | t_1__458_;
  assign t_2__455_ = t_1__455_ | t_1__457_;
  assign t_2__454_ = t_1__454_ | t_1__456_;
  assign t_2__453_ = t_1__453_ | t_1__455_;
  assign t_2__452_ = t_1__452_ | t_1__454_;
  assign t_2__451_ = t_1__451_ | t_1__453_;
  assign t_2__450_ = t_1__450_ | t_1__452_;
  assign t_2__449_ = t_1__449_ | t_1__451_;
  assign t_2__448_ = t_1__448_ | t_1__450_;
  assign t_2__447_ = t_1__447_ | t_1__449_;
  assign t_2__446_ = t_1__446_ | t_1__448_;
  assign t_2__445_ = t_1__445_ | t_1__447_;
  assign t_2__444_ = t_1__444_ | t_1__446_;
  assign t_2__443_ = t_1__443_ | t_1__445_;
  assign t_2__442_ = t_1__442_ | t_1__444_;
  assign t_2__441_ = t_1__441_ | t_1__443_;
  assign t_2__440_ = t_1__440_ | t_1__442_;
  assign t_2__439_ = t_1__439_ | t_1__441_;
  assign t_2__438_ = t_1__438_ | t_1__440_;
  assign t_2__437_ = t_1__437_ | t_1__439_;
  assign t_2__436_ = t_1__436_ | t_1__438_;
  assign t_2__435_ = t_1__435_ | t_1__437_;
  assign t_2__434_ = t_1__434_ | t_1__436_;
  assign t_2__433_ = t_1__433_ | t_1__435_;
  assign t_2__432_ = t_1__432_ | t_1__434_;
  assign t_2__431_ = t_1__431_ | t_1__433_;
  assign t_2__430_ = t_1__430_ | t_1__432_;
  assign t_2__429_ = t_1__429_ | t_1__431_;
  assign t_2__428_ = t_1__428_ | t_1__430_;
  assign t_2__427_ = t_1__427_ | t_1__429_;
  assign t_2__426_ = t_1__426_ | t_1__428_;
  assign t_2__425_ = t_1__425_ | t_1__427_;
  assign t_2__424_ = t_1__424_ | t_1__426_;
  assign t_2__423_ = t_1__423_ | t_1__425_;
  assign t_2__422_ = t_1__422_ | t_1__424_;
  assign t_2__421_ = t_1__421_ | t_1__423_;
  assign t_2__420_ = t_1__420_ | t_1__422_;
  assign t_2__419_ = t_1__419_ | t_1__421_;
  assign t_2__418_ = t_1__418_ | t_1__420_;
  assign t_2__417_ = t_1__417_ | t_1__419_;
  assign t_2__416_ = t_1__416_ | t_1__418_;
  assign t_2__415_ = t_1__415_ | t_1__417_;
  assign t_2__414_ = t_1__414_ | t_1__416_;
  assign t_2__413_ = t_1__413_ | t_1__415_;
  assign t_2__412_ = t_1__412_ | t_1__414_;
  assign t_2__411_ = t_1__411_ | t_1__413_;
  assign t_2__410_ = t_1__410_ | t_1__412_;
  assign t_2__409_ = t_1__409_ | t_1__411_;
  assign t_2__408_ = t_1__408_ | t_1__410_;
  assign t_2__407_ = t_1__407_ | t_1__409_;
  assign t_2__406_ = t_1__406_ | t_1__408_;
  assign t_2__405_ = t_1__405_ | t_1__407_;
  assign t_2__404_ = t_1__404_ | t_1__406_;
  assign t_2__403_ = t_1__403_ | t_1__405_;
  assign t_2__402_ = t_1__402_ | t_1__404_;
  assign t_2__401_ = t_1__401_ | t_1__403_;
  assign t_2__400_ = t_1__400_ | t_1__402_;
  assign t_2__399_ = t_1__399_ | t_1__401_;
  assign t_2__398_ = t_1__398_ | t_1__400_;
  assign t_2__397_ = t_1__397_ | t_1__399_;
  assign t_2__396_ = t_1__396_ | t_1__398_;
  assign t_2__395_ = t_1__395_ | t_1__397_;
  assign t_2__394_ = t_1__394_ | t_1__396_;
  assign t_2__393_ = t_1__393_ | t_1__395_;
  assign t_2__392_ = t_1__392_ | t_1__394_;
  assign t_2__391_ = t_1__391_ | t_1__393_;
  assign t_2__390_ = t_1__390_ | t_1__392_;
  assign t_2__389_ = t_1__389_ | t_1__391_;
  assign t_2__388_ = t_1__388_ | t_1__390_;
  assign t_2__387_ = t_1__387_ | t_1__389_;
  assign t_2__386_ = t_1__386_ | t_1__388_;
  assign t_2__385_ = t_1__385_ | t_1__387_;
  assign t_2__384_ = t_1__384_ | t_1__386_;
  assign t_2__383_ = t_1__383_ | t_1__385_;
  assign t_2__382_ = t_1__382_ | t_1__384_;
  assign t_2__381_ = t_1__381_ | t_1__383_;
  assign t_2__380_ = t_1__380_ | t_1__382_;
  assign t_2__379_ = t_1__379_ | t_1__381_;
  assign t_2__378_ = t_1__378_ | t_1__380_;
  assign t_2__377_ = t_1__377_ | t_1__379_;
  assign t_2__376_ = t_1__376_ | t_1__378_;
  assign t_2__375_ = t_1__375_ | t_1__377_;
  assign t_2__374_ = t_1__374_ | t_1__376_;
  assign t_2__373_ = t_1__373_ | t_1__375_;
  assign t_2__372_ = t_1__372_ | t_1__374_;
  assign t_2__371_ = t_1__371_ | t_1__373_;
  assign t_2__370_ = t_1__370_ | t_1__372_;
  assign t_2__369_ = t_1__369_ | t_1__371_;
  assign t_2__368_ = t_1__368_ | t_1__370_;
  assign t_2__367_ = t_1__367_ | t_1__369_;
  assign t_2__366_ = t_1__366_ | t_1__368_;
  assign t_2__365_ = t_1__365_ | t_1__367_;
  assign t_2__364_ = t_1__364_ | t_1__366_;
  assign t_2__363_ = t_1__363_ | t_1__365_;
  assign t_2__362_ = t_1__362_ | t_1__364_;
  assign t_2__361_ = t_1__361_ | t_1__363_;
  assign t_2__360_ = t_1__360_ | t_1__362_;
  assign t_2__359_ = t_1__359_ | t_1__361_;
  assign t_2__358_ = t_1__358_ | t_1__360_;
  assign t_2__357_ = t_1__357_ | t_1__359_;
  assign t_2__356_ = t_1__356_ | t_1__358_;
  assign t_2__355_ = t_1__355_ | t_1__357_;
  assign t_2__354_ = t_1__354_ | t_1__356_;
  assign t_2__353_ = t_1__353_ | t_1__355_;
  assign t_2__352_ = t_1__352_ | t_1__354_;
  assign t_2__351_ = t_1__351_ | t_1__353_;
  assign t_2__350_ = t_1__350_ | t_1__352_;
  assign t_2__349_ = t_1__349_ | t_1__351_;
  assign t_2__348_ = t_1__348_ | t_1__350_;
  assign t_2__347_ = t_1__347_ | t_1__349_;
  assign t_2__346_ = t_1__346_ | t_1__348_;
  assign t_2__345_ = t_1__345_ | t_1__347_;
  assign t_2__344_ = t_1__344_ | t_1__346_;
  assign t_2__343_ = t_1__343_ | t_1__345_;
  assign t_2__342_ = t_1__342_ | t_1__344_;
  assign t_2__341_ = t_1__341_ | t_1__343_;
  assign t_2__340_ = t_1__340_ | t_1__342_;
  assign t_2__339_ = t_1__339_ | t_1__341_;
  assign t_2__338_ = t_1__338_ | t_1__340_;
  assign t_2__337_ = t_1__337_ | t_1__339_;
  assign t_2__336_ = t_1__336_ | t_1__338_;
  assign t_2__335_ = t_1__335_ | t_1__337_;
  assign t_2__334_ = t_1__334_ | t_1__336_;
  assign t_2__333_ = t_1__333_ | t_1__335_;
  assign t_2__332_ = t_1__332_ | t_1__334_;
  assign t_2__331_ = t_1__331_ | t_1__333_;
  assign t_2__330_ = t_1__330_ | t_1__332_;
  assign t_2__329_ = t_1__329_ | t_1__331_;
  assign t_2__328_ = t_1__328_ | t_1__330_;
  assign t_2__327_ = t_1__327_ | t_1__329_;
  assign t_2__326_ = t_1__326_ | t_1__328_;
  assign t_2__325_ = t_1__325_ | t_1__327_;
  assign t_2__324_ = t_1__324_ | t_1__326_;
  assign t_2__323_ = t_1__323_ | t_1__325_;
  assign t_2__322_ = t_1__322_ | t_1__324_;
  assign t_2__321_ = t_1__321_ | t_1__323_;
  assign t_2__320_ = t_1__320_ | t_1__322_;
  assign t_2__319_ = t_1__319_ | t_1__321_;
  assign t_2__318_ = t_1__318_ | t_1__320_;
  assign t_2__317_ = t_1__317_ | t_1__319_;
  assign t_2__316_ = t_1__316_ | t_1__318_;
  assign t_2__315_ = t_1__315_ | t_1__317_;
  assign t_2__314_ = t_1__314_ | t_1__316_;
  assign t_2__313_ = t_1__313_ | t_1__315_;
  assign t_2__312_ = t_1__312_ | t_1__314_;
  assign t_2__311_ = t_1__311_ | t_1__313_;
  assign t_2__310_ = t_1__310_ | t_1__312_;
  assign t_2__309_ = t_1__309_ | t_1__311_;
  assign t_2__308_ = t_1__308_ | t_1__310_;
  assign t_2__307_ = t_1__307_ | t_1__309_;
  assign t_2__306_ = t_1__306_ | t_1__308_;
  assign t_2__305_ = t_1__305_ | t_1__307_;
  assign t_2__304_ = t_1__304_ | t_1__306_;
  assign t_2__303_ = t_1__303_ | t_1__305_;
  assign t_2__302_ = t_1__302_ | t_1__304_;
  assign t_2__301_ = t_1__301_ | t_1__303_;
  assign t_2__300_ = t_1__300_ | t_1__302_;
  assign t_2__299_ = t_1__299_ | t_1__301_;
  assign t_2__298_ = t_1__298_ | t_1__300_;
  assign t_2__297_ = t_1__297_ | t_1__299_;
  assign t_2__296_ = t_1__296_ | t_1__298_;
  assign t_2__295_ = t_1__295_ | t_1__297_;
  assign t_2__294_ = t_1__294_ | t_1__296_;
  assign t_2__293_ = t_1__293_ | t_1__295_;
  assign t_2__292_ = t_1__292_ | t_1__294_;
  assign t_2__291_ = t_1__291_ | t_1__293_;
  assign t_2__290_ = t_1__290_ | t_1__292_;
  assign t_2__289_ = t_1__289_ | t_1__291_;
  assign t_2__288_ = t_1__288_ | t_1__290_;
  assign t_2__287_ = t_1__287_ | t_1__289_;
  assign t_2__286_ = t_1__286_ | t_1__288_;
  assign t_2__285_ = t_1__285_ | t_1__287_;
  assign t_2__284_ = t_1__284_ | t_1__286_;
  assign t_2__283_ = t_1__283_ | t_1__285_;
  assign t_2__282_ = t_1__282_ | t_1__284_;
  assign t_2__281_ = t_1__281_ | t_1__283_;
  assign t_2__280_ = t_1__280_ | t_1__282_;
  assign t_2__279_ = t_1__279_ | t_1__281_;
  assign t_2__278_ = t_1__278_ | t_1__280_;
  assign t_2__277_ = t_1__277_ | t_1__279_;
  assign t_2__276_ = t_1__276_ | t_1__278_;
  assign t_2__275_ = t_1__275_ | t_1__277_;
  assign t_2__274_ = t_1__274_ | t_1__276_;
  assign t_2__273_ = t_1__273_ | t_1__275_;
  assign t_2__272_ = t_1__272_ | t_1__274_;
  assign t_2__271_ = t_1__271_ | t_1__273_;
  assign t_2__270_ = t_1__270_ | t_1__272_;
  assign t_2__269_ = t_1__269_ | t_1__271_;
  assign t_2__268_ = t_1__268_ | t_1__270_;
  assign t_2__267_ = t_1__267_ | t_1__269_;
  assign t_2__266_ = t_1__266_ | t_1__268_;
  assign t_2__265_ = t_1__265_ | t_1__267_;
  assign t_2__264_ = t_1__264_ | t_1__266_;
  assign t_2__263_ = t_1__263_ | t_1__265_;
  assign t_2__262_ = t_1__262_ | t_1__264_;
  assign t_2__261_ = t_1__261_ | t_1__263_;
  assign t_2__260_ = t_1__260_ | t_1__262_;
  assign t_2__259_ = t_1__259_ | t_1__261_;
  assign t_2__258_ = t_1__258_ | t_1__260_;
  assign t_2__257_ = t_1__257_ | t_1__259_;
  assign t_2__256_ = t_1__256_ | t_1__258_;
  assign t_2__255_ = t_1__255_ | t_1__257_;
  assign t_2__254_ = t_1__254_ | t_1__256_;
  assign t_2__253_ = t_1__253_ | t_1__255_;
  assign t_2__252_ = t_1__252_ | t_1__254_;
  assign t_2__251_ = t_1__251_ | t_1__253_;
  assign t_2__250_ = t_1__250_ | t_1__252_;
  assign t_2__249_ = t_1__249_ | t_1__251_;
  assign t_2__248_ = t_1__248_ | t_1__250_;
  assign t_2__247_ = t_1__247_ | t_1__249_;
  assign t_2__246_ = t_1__246_ | t_1__248_;
  assign t_2__245_ = t_1__245_ | t_1__247_;
  assign t_2__244_ = t_1__244_ | t_1__246_;
  assign t_2__243_ = t_1__243_ | t_1__245_;
  assign t_2__242_ = t_1__242_ | t_1__244_;
  assign t_2__241_ = t_1__241_ | t_1__243_;
  assign t_2__240_ = t_1__240_ | t_1__242_;
  assign t_2__239_ = t_1__239_ | t_1__241_;
  assign t_2__238_ = t_1__238_ | t_1__240_;
  assign t_2__237_ = t_1__237_ | t_1__239_;
  assign t_2__236_ = t_1__236_ | t_1__238_;
  assign t_2__235_ = t_1__235_ | t_1__237_;
  assign t_2__234_ = t_1__234_ | t_1__236_;
  assign t_2__233_ = t_1__233_ | t_1__235_;
  assign t_2__232_ = t_1__232_ | t_1__234_;
  assign t_2__231_ = t_1__231_ | t_1__233_;
  assign t_2__230_ = t_1__230_ | t_1__232_;
  assign t_2__229_ = t_1__229_ | t_1__231_;
  assign t_2__228_ = t_1__228_ | t_1__230_;
  assign t_2__227_ = t_1__227_ | t_1__229_;
  assign t_2__226_ = t_1__226_ | t_1__228_;
  assign t_2__225_ = t_1__225_ | t_1__227_;
  assign t_2__224_ = t_1__224_ | t_1__226_;
  assign t_2__223_ = t_1__223_ | t_1__225_;
  assign t_2__222_ = t_1__222_ | t_1__224_;
  assign t_2__221_ = t_1__221_ | t_1__223_;
  assign t_2__220_ = t_1__220_ | t_1__222_;
  assign t_2__219_ = t_1__219_ | t_1__221_;
  assign t_2__218_ = t_1__218_ | t_1__220_;
  assign t_2__217_ = t_1__217_ | t_1__219_;
  assign t_2__216_ = t_1__216_ | t_1__218_;
  assign t_2__215_ = t_1__215_ | t_1__217_;
  assign t_2__214_ = t_1__214_ | t_1__216_;
  assign t_2__213_ = t_1__213_ | t_1__215_;
  assign t_2__212_ = t_1__212_ | t_1__214_;
  assign t_2__211_ = t_1__211_ | t_1__213_;
  assign t_2__210_ = t_1__210_ | t_1__212_;
  assign t_2__209_ = t_1__209_ | t_1__211_;
  assign t_2__208_ = t_1__208_ | t_1__210_;
  assign t_2__207_ = t_1__207_ | t_1__209_;
  assign t_2__206_ = t_1__206_ | t_1__208_;
  assign t_2__205_ = t_1__205_ | t_1__207_;
  assign t_2__204_ = t_1__204_ | t_1__206_;
  assign t_2__203_ = t_1__203_ | t_1__205_;
  assign t_2__202_ = t_1__202_ | t_1__204_;
  assign t_2__201_ = t_1__201_ | t_1__203_;
  assign t_2__200_ = t_1__200_ | t_1__202_;
  assign t_2__199_ = t_1__199_ | t_1__201_;
  assign t_2__198_ = t_1__198_ | t_1__200_;
  assign t_2__197_ = t_1__197_ | t_1__199_;
  assign t_2__196_ = t_1__196_ | t_1__198_;
  assign t_2__195_ = t_1__195_ | t_1__197_;
  assign t_2__194_ = t_1__194_ | t_1__196_;
  assign t_2__193_ = t_1__193_ | t_1__195_;
  assign t_2__192_ = t_1__192_ | t_1__194_;
  assign t_2__191_ = t_1__191_ | t_1__193_;
  assign t_2__190_ = t_1__190_ | t_1__192_;
  assign t_2__189_ = t_1__189_ | t_1__191_;
  assign t_2__188_ = t_1__188_ | t_1__190_;
  assign t_2__187_ = t_1__187_ | t_1__189_;
  assign t_2__186_ = t_1__186_ | t_1__188_;
  assign t_2__185_ = t_1__185_ | t_1__187_;
  assign t_2__184_ = t_1__184_ | t_1__186_;
  assign t_2__183_ = t_1__183_ | t_1__185_;
  assign t_2__182_ = t_1__182_ | t_1__184_;
  assign t_2__181_ = t_1__181_ | t_1__183_;
  assign t_2__180_ = t_1__180_ | t_1__182_;
  assign t_2__179_ = t_1__179_ | t_1__181_;
  assign t_2__178_ = t_1__178_ | t_1__180_;
  assign t_2__177_ = t_1__177_ | t_1__179_;
  assign t_2__176_ = t_1__176_ | t_1__178_;
  assign t_2__175_ = t_1__175_ | t_1__177_;
  assign t_2__174_ = t_1__174_ | t_1__176_;
  assign t_2__173_ = t_1__173_ | t_1__175_;
  assign t_2__172_ = t_1__172_ | t_1__174_;
  assign t_2__171_ = t_1__171_ | t_1__173_;
  assign t_2__170_ = t_1__170_ | t_1__172_;
  assign t_2__169_ = t_1__169_ | t_1__171_;
  assign t_2__168_ = t_1__168_ | t_1__170_;
  assign t_2__167_ = t_1__167_ | t_1__169_;
  assign t_2__166_ = t_1__166_ | t_1__168_;
  assign t_2__165_ = t_1__165_ | t_1__167_;
  assign t_2__164_ = t_1__164_ | t_1__166_;
  assign t_2__163_ = t_1__163_ | t_1__165_;
  assign t_2__162_ = t_1__162_ | t_1__164_;
  assign t_2__161_ = t_1__161_ | t_1__163_;
  assign t_2__160_ = t_1__160_ | t_1__162_;
  assign t_2__159_ = t_1__159_ | t_1__161_;
  assign t_2__158_ = t_1__158_ | t_1__160_;
  assign t_2__157_ = t_1__157_ | t_1__159_;
  assign t_2__156_ = t_1__156_ | t_1__158_;
  assign t_2__155_ = t_1__155_ | t_1__157_;
  assign t_2__154_ = t_1__154_ | t_1__156_;
  assign t_2__153_ = t_1__153_ | t_1__155_;
  assign t_2__152_ = t_1__152_ | t_1__154_;
  assign t_2__151_ = t_1__151_ | t_1__153_;
  assign t_2__150_ = t_1__150_ | t_1__152_;
  assign t_2__149_ = t_1__149_ | t_1__151_;
  assign t_2__148_ = t_1__148_ | t_1__150_;
  assign t_2__147_ = t_1__147_ | t_1__149_;
  assign t_2__146_ = t_1__146_ | t_1__148_;
  assign t_2__145_ = t_1__145_ | t_1__147_;
  assign t_2__144_ = t_1__144_ | t_1__146_;
  assign t_2__143_ = t_1__143_ | t_1__145_;
  assign t_2__142_ = t_1__142_ | t_1__144_;
  assign t_2__141_ = t_1__141_ | t_1__143_;
  assign t_2__140_ = t_1__140_ | t_1__142_;
  assign t_2__139_ = t_1__139_ | t_1__141_;
  assign t_2__138_ = t_1__138_ | t_1__140_;
  assign t_2__137_ = t_1__137_ | t_1__139_;
  assign t_2__136_ = t_1__136_ | t_1__138_;
  assign t_2__135_ = t_1__135_ | t_1__137_;
  assign t_2__134_ = t_1__134_ | t_1__136_;
  assign t_2__133_ = t_1__133_ | t_1__135_;
  assign t_2__132_ = t_1__132_ | t_1__134_;
  assign t_2__131_ = t_1__131_ | t_1__133_;
  assign t_2__130_ = t_1__130_ | t_1__132_;
  assign t_2__129_ = t_1__129_ | t_1__131_;
  assign t_2__128_ = t_1__128_ | t_1__130_;
  assign t_2__127_ = t_1__127_ | t_1__129_;
  assign t_2__126_ = t_1__126_ | t_1__128_;
  assign t_2__125_ = t_1__125_ | t_1__127_;
  assign t_2__124_ = t_1__124_ | t_1__126_;
  assign t_2__123_ = t_1__123_ | t_1__125_;
  assign t_2__122_ = t_1__122_ | t_1__124_;
  assign t_2__121_ = t_1__121_ | t_1__123_;
  assign t_2__120_ = t_1__120_ | t_1__122_;
  assign t_2__119_ = t_1__119_ | t_1__121_;
  assign t_2__118_ = t_1__118_ | t_1__120_;
  assign t_2__117_ = t_1__117_ | t_1__119_;
  assign t_2__116_ = t_1__116_ | t_1__118_;
  assign t_2__115_ = t_1__115_ | t_1__117_;
  assign t_2__114_ = t_1__114_ | t_1__116_;
  assign t_2__113_ = t_1__113_ | t_1__115_;
  assign t_2__112_ = t_1__112_ | t_1__114_;
  assign t_2__111_ = t_1__111_ | t_1__113_;
  assign t_2__110_ = t_1__110_ | t_1__112_;
  assign t_2__109_ = t_1__109_ | t_1__111_;
  assign t_2__108_ = t_1__108_ | t_1__110_;
  assign t_2__107_ = t_1__107_ | t_1__109_;
  assign t_2__106_ = t_1__106_ | t_1__108_;
  assign t_2__105_ = t_1__105_ | t_1__107_;
  assign t_2__104_ = t_1__104_ | t_1__106_;
  assign t_2__103_ = t_1__103_ | t_1__105_;
  assign t_2__102_ = t_1__102_ | t_1__104_;
  assign t_2__101_ = t_1__101_ | t_1__103_;
  assign t_2__100_ = t_1__100_ | t_1__102_;
  assign t_2__99_ = t_1__99_ | t_1__101_;
  assign t_2__98_ = t_1__98_ | t_1__100_;
  assign t_2__97_ = t_1__97_ | t_1__99_;
  assign t_2__96_ = t_1__96_ | t_1__98_;
  assign t_2__95_ = t_1__95_ | t_1__97_;
  assign t_2__94_ = t_1__94_ | t_1__96_;
  assign t_2__93_ = t_1__93_ | t_1__95_;
  assign t_2__92_ = t_1__92_ | t_1__94_;
  assign t_2__91_ = t_1__91_ | t_1__93_;
  assign t_2__90_ = t_1__90_ | t_1__92_;
  assign t_2__89_ = t_1__89_ | t_1__91_;
  assign t_2__88_ = t_1__88_ | t_1__90_;
  assign t_2__87_ = t_1__87_ | t_1__89_;
  assign t_2__86_ = t_1__86_ | t_1__88_;
  assign t_2__85_ = t_1__85_ | t_1__87_;
  assign t_2__84_ = t_1__84_ | t_1__86_;
  assign t_2__83_ = t_1__83_ | t_1__85_;
  assign t_2__82_ = t_1__82_ | t_1__84_;
  assign t_2__81_ = t_1__81_ | t_1__83_;
  assign t_2__80_ = t_1__80_ | t_1__82_;
  assign t_2__79_ = t_1__79_ | t_1__81_;
  assign t_2__78_ = t_1__78_ | t_1__80_;
  assign t_2__77_ = t_1__77_ | t_1__79_;
  assign t_2__76_ = t_1__76_ | t_1__78_;
  assign t_2__75_ = t_1__75_ | t_1__77_;
  assign t_2__74_ = t_1__74_ | t_1__76_;
  assign t_2__73_ = t_1__73_ | t_1__75_;
  assign t_2__72_ = t_1__72_ | t_1__74_;
  assign t_2__71_ = t_1__71_ | t_1__73_;
  assign t_2__70_ = t_1__70_ | t_1__72_;
  assign t_2__69_ = t_1__69_ | t_1__71_;
  assign t_2__68_ = t_1__68_ | t_1__70_;
  assign t_2__67_ = t_1__67_ | t_1__69_;
  assign t_2__66_ = t_1__66_ | t_1__68_;
  assign t_2__65_ = t_1__65_ | t_1__67_;
  assign t_2__64_ = t_1__64_ | t_1__66_;
  assign t_2__63_ = t_1__63_ | t_1__65_;
  assign t_2__62_ = t_1__62_ | t_1__64_;
  assign t_2__61_ = t_1__61_ | t_1__63_;
  assign t_2__60_ = t_1__60_ | t_1__62_;
  assign t_2__59_ = t_1__59_ | t_1__61_;
  assign t_2__58_ = t_1__58_ | t_1__60_;
  assign t_2__57_ = t_1__57_ | t_1__59_;
  assign t_2__56_ = t_1__56_ | t_1__58_;
  assign t_2__55_ = t_1__55_ | t_1__57_;
  assign t_2__54_ = t_1__54_ | t_1__56_;
  assign t_2__53_ = t_1__53_ | t_1__55_;
  assign t_2__52_ = t_1__52_ | t_1__54_;
  assign t_2__51_ = t_1__51_ | t_1__53_;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__511_ = t_2__511_ | 1'b0;
  assign t_3__510_ = t_2__510_ | 1'b0;
  assign t_3__509_ = t_2__509_ | 1'b0;
  assign t_3__508_ = t_2__508_ | 1'b0;
  assign t_3__507_ = t_2__507_ | t_2__511_;
  assign t_3__506_ = t_2__506_ | t_2__510_;
  assign t_3__505_ = t_2__505_ | t_2__509_;
  assign t_3__504_ = t_2__504_ | t_2__508_;
  assign t_3__503_ = t_2__503_ | t_2__507_;
  assign t_3__502_ = t_2__502_ | t_2__506_;
  assign t_3__501_ = t_2__501_ | t_2__505_;
  assign t_3__500_ = t_2__500_ | t_2__504_;
  assign t_3__499_ = t_2__499_ | t_2__503_;
  assign t_3__498_ = t_2__498_ | t_2__502_;
  assign t_3__497_ = t_2__497_ | t_2__501_;
  assign t_3__496_ = t_2__496_ | t_2__500_;
  assign t_3__495_ = t_2__495_ | t_2__499_;
  assign t_3__494_ = t_2__494_ | t_2__498_;
  assign t_3__493_ = t_2__493_ | t_2__497_;
  assign t_3__492_ = t_2__492_ | t_2__496_;
  assign t_3__491_ = t_2__491_ | t_2__495_;
  assign t_3__490_ = t_2__490_ | t_2__494_;
  assign t_3__489_ = t_2__489_ | t_2__493_;
  assign t_3__488_ = t_2__488_ | t_2__492_;
  assign t_3__487_ = t_2__487_ | t_2__491_;
  assign t_3__486_ = t_2__486_ | t_2__490_;
  assign t_3__485_ = t_2__485_ | t_2__489_;
  assign t_3__484_ = t_2__484_ | t_2__488_;
  assign t_3__483_ = t_2__483_ | t_2__487_;
  assign t_3__482_ = t_2__482_ | t_2__486_;
  assign t_3__481_ = t_2__481_ | t_2__485_;
  assign t_3__480_ = t_2__480_ | t_2__484_;
  assign t_3__479_ = t_2__479_ | t_2__483_;
  assign t_3__478_ = t_2__478_ | t_2__482_;
  assign t_3__477_ = t_2__477_ | t_2__481_;
  assign t_3__476_ = t_2__476_ | t_2__480_;
  assign t_3__475_ = t_2__475_ | t_2__479_;
  assign t_3__474_ = t_2__474_ | t_2__478_;
  assign t_3__473_ = t_2__473_ | t_2__477_;
  assign t_3__472_ = t_2__472_ | t_2__476_;
  assign t_3__471_ = t_2__471_ | t_2__475_;
  assign t_3__470_ = t_2__470_ | t_2__474_;
  assign t_3__469_ = t_2__469_ | t_2__473_;
  assign t_3__468_ = t_2__468_ | t_2__472_;
  assign t_3__467_ = t_2__467_ | t_2__471_;
  assign t_3__466_ = t_2__466_ | t_2__470_;
  assign t_3__465_ = t_2__465_ | t_2__469_;
  assign t_3__464_ = t_2__464_ | t_2__468_;
  assign t_3__463_ = t_2__463_ | t_2__467_;
  assign t_3__462_ = t_2__462_ | t_2__466_;
  assign t_3__461_ = t_2__461_ | t_2__465_;
  assign t_3__460_ = t_2__460_ | t_2__464_;
  assign t_3__459_ = t_2__459_ | t_2__463_;
  assign t_3__458_ = t_2__458_ | t_2__462_;
  assign t_3__457_ = t_2__457_ | t_2__461_;
  assign t_3__456_ = t_2__456_ | t_2__460_;
  assign t_3__455_ = t_2__455_ | t_2__459_;
  assign t_3__454_ = t_2__454_ | t_2__458_;
  assign t_3__453_ = t_2__453_ | t_2__457_;
  assign t_3__452_ = t_2__452_ | t_2__456_;
  assign t_3__451_ = t_2__451_ | t_2__455_;
  assign t_3__450_ = t_2__450_ | t_2__454_;
  assign t_3__449_ = t_2__449_ | t_2__453_;
  assign t_3__448_ = t_2__448_ | t_2__452_;
  assign t_3__447_ = t_2__447_ | t_2__451_;
  assign t_3__446_ = t_2__446_ | t_2__450_;
  assign t_3__445_ = t_2__445_ | t_2__449_;
  assign t_3__444_ = t_2__444_ | t_2__448_;
  assign t_3__443_ = t_2__443_ | t_2__447_;
  assign t_3__442_ = t_2__442_ | t_2__446_;
  assign t_3__441_ = t_2__441_ | t_2__445_;
  assign t_3__440_ = t_2__440_ | t_2__444_;
  assign t_3__439_ = t_2__439_ | t_2__443_;
  assign t_3__438_ = t_2__438_ | t_2__442_;
  assign t_3__437_ = t_2__437_ | t_2__441_;
  assign t_3__436_ = t_2__436_ | t_2__440_;
  assign t_3__435_ = t_2__435_ | t_2__439_;
  assign t_3__434_ = t_2__434_ | t_2__438_;
  assign t_3__433_ = t_2__433_ | t_2__437_;
  assign t_3__432_ = t_2__432_ | t_2__436_;
  assign t_3__431_ = t_2__431_ | t_2__435_;
  assign t_3__430_ = t_2__430_ | t_2__434_;
  assign t_3__429_ = t_2__429_ | t_2__433_;
  assign t_3__428_ = t_2__428_ | t_2__432_;
  assign t_3__427_ = t_2__427_ | t_2__431_;
  assign t_3__426_ = t_2__426_ | t_2__430_;
  assign t_3__425_ = t_2__425_ | t_2__429_;
  assign t_3__424_ = t_2__424_ | t_2__428_;
  assign t_3__423_ = t_2__423_ | t_2__427_;
  assign t_3__422_ = t_2__422_ | t_2__426_;
  assign t_3__421_ = t_2__421_ | t_2__425_;
  assign t_3__420_ = t_2__420_ | t_2__424_;
  assign t_3__419_ = t_2__419_ | t_2__423_;
  assign t_3__418_ = t_2__418_ | t_2__422_;
  assign t_3__417_ = t_2__417_ | t_2__421_;
  assign t_3__416_ = t_2__416_ | t_2__420_;
  assign t_3__415_ = t_2__415_ | t_2__419_;
  assign t_3__414_ = t_2__414_ | t_2__418_;
  assign t_3__413_ = t_2__413_ | t_2__417_;
  assign t_3__412_ = t_2__412_ | t_2__416_;
  assign t_3__411_ = t_2__411_ | t_2__415_;
  assign t_3__410_ = t_2__410_ | t_2__414_;
  assign t_3__409_ = t_2__409_ | t_2__413_;
  assign t_3__408_ = t_2__408_ | t_2__412_;
  assign t_3__407_ = t_2__407_ | t_2__411_;
  assign t_3__406_ = t_2__406_ | t_2__410_;
  assign t_3__405_ = t_2__405_ | t_2__409_;
  assign t_3__404_ = t_2__404_ | t_2__408_;
  assign t_3__403_ = t_2__403_ | t_2__407_;
  assign t_3__402_ = t_2__402_ | t_2__406_;
  assign t_3__401_ = t_2__401_ | t_2__405_;
  assign t_3__400_ = t_2__400_ | t_2__404_;
  assign t_3__399_ = t_2__399_ | t_2__403_;
  assign t_3__398_ = t_2__398_ | t_2__402_;
  assign t_3__397_ = t_2__397_ | t_2__401_;
  assign t_3__396_ = t_2__396_ | t_2__400_;
  assign t_3__395_ = t_2__395_ | t_2__399_;
  assign t_3__394_ = t_2__394_ | t_2__398_;
  assign t_3__393_ = t_2__393_ | t_2__397_;
  assign t_3__392_ = t_2__392_ | t_2__396_;
  assign t_3__391_ = t_2__391_ | t_2__395_;
  assign t_3__390_ = t_2__390_ | t_2__394_;
  assign t_3__389_ = t_2__389_ | t_2__393_;
  assign t_3__388_ = t_2__388_ | t_2__392_;
  assign t_3__387_ = t_2__387_ | t_2__391_;
  assign t_3__386_ = t_2__386_ | t_2__390_;
  assign t_3__385_ = t_2__385_ | t_2__389_;
  assign t_3__384_ = t_2__384_ | t_2__388_;
  assign t_3__383_ = t_2__383_ | t_2__387_;
  assign t_3__382_ = t_2__382_ | t_2__386_;
  assign t_3__381_ = t_2__381_ | t_2__385_;
  assign t_3__380_ = t_2__380_ | t_2__384_;
  assign t_3__379_ = t_2__379_ | t_2__383_;
  assign t_3__378_ = t_2__378_ | t_2__382_;
  assign t_3__377_ = t_2__377_ | t_2__381_;
  assign t_3__376_ = t_2__376_ | t_2__380_;
  assign t_3__375_ = t_2__375_ | t_2__379_;
  assign t_3__374_ = t_2__374_ | t_2__378_;
  assign t_3__373_ = t_2__373_ | t_2__377_;
  assign t_3__372_ = t_2__372_ | t_2__376_;
  assign t_3__371_ = t_2__371_ | t_2__375_;
  assign t_3__370_ = t_2__370_ | t_2__374_;
  assign t_3__369_ = t_2__369_ | t_2__373_;
  assign t_3__368_ = t_2__368_ | t_2__372_;
  assign t_3__367_ = t_2__367_ | t_2__371_;
  assign t_3__366_ = t_2__366_ | t_2__370_;
  assign t_3__365_ = t_2__365_ | t_2__369_;
  assign t_3__364_ = t_2__364_ | t_2__368_;
  assign t_3__363_ = t_2__363_ | t_2__367_;
  assign t_3__362_ = t_2__362_ | t_2__366_;
  assign t_3__361_ = t_2__361_ | t_2__365_;
  assign t_3__360_ = t_2__360_ | t_2__364_;
  assign t_3__359_ = t_2__359_ | t_2__363_;
  assign t_3__358_ = t_2__358_ | t_2__362_;
  assign t_3__357_ = t_2__357_ | t_2__361_;
  assign t_3__356_ = t_2__356_ | t_2__360_;
  assign t_3__355_ = t_2__355_ | t_2__359_;
  assign t_3__354_ = t_2__354_ | t_2__358_;
  assign t_3__353_ = t_2__353_ | t_2__357_;
  assign t_3__352_ = t_2__352_ | t_2__356_;
  assign t_3__351_ = t_2__351_ | t_2__355_;
  assign t_3__350_ = t_2__350_ | t_2__354_;
  assign t_3__349_ = t_2__349_ | t_2__353_;
  assign t_3__348_ = t_2__348_ | t_2__352_;
  assign t_3__347_ = t_2__347_ | t_2__351_;
  assign t_3__346_ = t_2__346_ | t_2__350_;
  assign t_3__345_ = t_2__345_ | t_2__349_;
  assign t_3__344_ = t_2__344_ | t_2__348_;
  assign t_3__343_ = t_2__343_ | t_2__347_;
  assign t_3__342_ = t_2__342_ | t_2__346_;
  assign t_3__341_ = t_2__341_ | t_2__345_;
  assign t_3__340_ = t_2__340_ | t_2__344_;
  assign t_3__339_ = t_2__339_ | t_2__343_;
  assign t_3__338_ = t_2__338_ | t_2__342_;
  assign t_3__337_ = t_2__337_ | t_2__341_;
  assign t_3__336_ = t_2__336_ | t_2__340_;
  assign t_3__335_ = t_2__335_ | t_2__339_;
  assign t_3__334_ = t_2__334_ | t_2__338_;
  assign t_3__333_ = t_2__333_ | t_2__337_;
  assign t_3__332_ = t_2__332_ | t_2__336_;
  assign t_3__331_ = t_2__331_ | t_2__335_;
  assign t_3__330_ = t_2__330_ | t_2__334_;
  assign t_3__329_ = t_2__329_ | t_2__333_;
  assign t_3__328_ = t_2__328_ | t_2__332_;
  assign t_3__327_ = t_2__327_ | t_2__331_;
  assign t_3__326_ = t_2__326_ | t_2__330_;
  assign t_3__325_ = t_2__325_ | t_2__329_;
  assign t_3__324_ = t_2__324_ | t_2__328_;
  assign t_3__323_ = t_2__323_ | t_2__327_;
  assign t_3__322_ = t_2__322_ | t_2__326_;
  assign t_3__321_ = t_2__321_ | t_2__325_;
  assign t_3__320_ = t_2__320_ | t_2__324_;
  assign t_3__319_ = t_2__319_ | t_2__323_;
  assign t_3__318_ = t_2__318_ | t_2__322_;
  assign t_3__317_ = t_2__317_ | t_2__321_;
  assign t_3__316_ = t_2__316_ | t_2__320_;
  assign t_3__315_ = t_2__315_ | t_2__319_;
  assign t_3__314_ = t_2__314_ | t_2__318_;
  assign t_3__313_ = t_2__313_ | t_2__317_;
  assign t_3__312_ = t_2__312_ | t_2__316_;
  assign t_3__311_ = t_2__311_ | t_2__315_;
  assign t_3__310_ = t_2__310_ | t_2__314_;
  assign t_3__309_ = t_2__309_ | t_2__313_;
  assign t_3__308_ = t_2__308_ | t_2__312_;
  assign t_3__307_ = t_2__307_ | t_2__311_;
  assign t_3__306_ = t_2__306_ | t_2__310_;
  assign t_3__305_ = t_2__305_ | t_2__309_;
  assign t_3__304_ = t_2__304_ | t_2__308_;
  assign t_3__303_ = t_2__303_ | t_2__307_;
  assign t_3__302_ = t_2__302_ | t_2__306_;
  assign t_3__301_ = t_2__301_ | t_2__305_;
  assign t_3__300_ = t_2__300_ | t_2__304_;
  assign t_3__299_ = t_2__299_ | t_2__303_;
  assign t_3__298_ = t_2__298_ | t_2__302_;
  assign t_3__297_ = t_2__297_ | t_2__301_;
  assign t_3__296_ = t_2__296_ | t_2__300_;
  assign t_3__295_ = t_2__295_ | t_2__299_;
  assign t_3__294_ = t_2__294_ | t_2__298_;
  assign t_3__293_ = t_2__293_ | t_2__297_;
  assign t_3__292_ = t_2__292_ | t_2__296_;
  assign t_3__291_ = t_2__291_ | t_2__295_;
  assign t_3__290_ = t_2__290_ | t_2__294_;
  assign t_3__289_ = t_2__289_ | t_2__293_;
  assign t_3__288_ = t_2__288_ | t_2__292_;
  assign t_3__287_ = t_2__287_ | t_2__291_;
  assign t_3__286_ = t_2__286_ | t_2__290_;
  assign t_3__285_ = t_2__285_ | t_2__289_;
  assign t_3__284_ = t_2__284_ | t_2__288_;
  assign t_3__283_ = t_2__283_ | t_2__287_;
  assign t_3__282_ = t_2__282_ | t_2__286_;
  assign t_3__281_ = t_2__281_ | t_2__285_;
  assign t_3__280_ = t_2__280_ | t_2__284_;
  assign t_3__279_ = t_2__279_ | t_2__283_;
  assign t_3__278_ = t_2__278_ | t_2__282_;
  assign t_3__277_ = t_2__277_ | t_2__281_;
  assign t_3__276_ = t_2__276_ | t_2__280_;
  assign t_3__275_ = t_2__275_ | t_2__279_;
  assign t_3__274_ = t_2__274_ | t_2__278_;
  assign t_3__273_ = t_2__273_ | t_2__277_;
  assign t_3__272_ = t_2__272_ | t_2__276_;
  assign t_3__271_ = t_2__271_ | t_2__275_;
  assign t_3__270_ = t_2__270_ | t_2__274_;
  assign t_3__269_ = t_2__269_ | t_2__273_;
  assign t_3__268_ = t_2__268_ | t_2__272_;
  assign t_3__267_ = t_2__267_ | t_2__271_;
  assign t_3__266_ = t_2__266_ | t_2__270_;
  assign t_3__265_ = t_2__265_ | t_2__269_;
  assign t_3__264_ = t_2__264_ | t_2__268_;
  assign t_3__263_ = t_2__263_ | t_2__267_;
  assign t_3__262_ = t_2__262_ | t_2__266_;
  assign t_3__261_ = t_2__261_ | t_2__265_;
  assign t_3__260_ = t_2__260_ | t_2__264_;
  assign t_3__259_ = t_2__259_ | t_2__263_;
  assign t_3__258_ = t_2__258_ | t_2__262_;
  assign t_3__257_ = t_2__257_ | t_2__261_;
  assign t_3__256_ = t_2__256_ | t_2__260_;
  assign t_3__255_ = t_2__255_ | t_2__259_;
  assign t_3__254_ = t_2__254_ | t_2__258_;
  assign t_3__253_ = t_2__253_ | t_2__257_;
  assign t_3__252_ = t_2__252_ | t_2__256_;
  assign t_3__251_ = t_2__251_ | t_2__255_;
  assign t_3__250_ = t_2__250_ | t_2__254_;
  assign t_3__249_ = t_2__249_ | t_2__253_;
  assign t_3__248_ = t_2__248_ | t_2__252_;
  assign t_3__247_ = t_2__247_ | t_2__251_;
  assign t_3__246_ = t_2__246_ | t_2__250_;
  assign t_3__245_ = t_2__245_ | t_2__249_;
  assign t_3__244_ = t_2__244_ | t_2__248_;
  assign t_3__243_ = t_2__243_ | t_2__247_;
  assign t_3__242_ = t_2__242_ | t_2__246_;
  assign t_3__241_ = t_2__241_ | t_2__245_;
  assign t_3__240_ = t_2__240_ | t_2__244_;
  assign t_3__239_ = t_2__239_ | t_2__243_;
  assign t_3__238_ = t_2__238_ | t_2__242_;
  assign t_3__237_ = t_2__237_ | t_2__241_;
  assign t_3__236_ = t_2__236_ | t_2__240_;
  assign t_3__235_ = t_2__235_ | t_2__239_;
  assign t_3__234_ = t_2__234_ | t_2__238_;
  assign t_3__233_ = t_2__233_ | t_2__237_;
  assign t_3__232_ = t_2__232_ | t_2__236_;
  assign t_3__231_ = t_2__231_ | t_2__235_;
  assign t_3__230_ = t_2__230_ | t_2__234_;
  assign t_3__229_ = t_2__229_ | t_2__233_;
  assign t_3__228_ = t_2__228_ | t_2__232_;
  assign t_3__227_ = t_2__227_ | t_2__231_;
  assign t_3__226_ = t_2__226_ | t_2__230_;
  assign t_3__225_ = t_2__225_ | t_2__229_;
  assign t_3__224_ = t_2__224_ | t_2__228_;
  assign t_3__223_ = t_2__223_ | t_2__227_;
  assign t_3__222_ = t_2__222_ | t_2__226_;
  assign t_3__221_ = t_2__221_ | t_2__225_;
  assign t_3__220_ = t_2__220_ | t_2__224_;
  assign t_3__219_ = t_2__219_ | t_2__223_;
  assign t_3__218_ = t_2__218_ | t_2__222_;
  assign t_3__217_ = t_2__217_ | t_2__221_;
  assign t_3__216_ = t_2__216_ | t_2__220_;
  assign t_3__215_ = t_2__215_ | t_2__219_;
  assign t_3__214_ = t_2__214_ | t_2__218_;
  assign t_3__213_ = t_2__213_ | t_2__217_;
  assign t_3__212_ = t_2__212_ | t_2__216_;
  assign t_3__211_ = t_2__211_ | t_2__215_;
  assign t_3__210_ = t_2__210_ | t_2__214_;
  assign t_3__209_ = t_2__209_ | t_2__213_;
  assign t_3__208_ = t_2__208_ | t_2__212_;
  assign t_3__207_ = t_2__207_ | t_2__211_;
  assign t_3__206_ = t_2__206_ | t_2__210_;
  assign t_3__205_ = t_2__205_ | t_2__209_;
  assign t_3__204_ = t_2__204_ | t_2__208_;
  assign t_3__203_ = t_2__203_ | t_2__207_;
  assign t_3__202_ = t_2__202_ | t_2__206_;
  assign t_3__201_ = t_2__201_ | t_2__205_;
  assign t_3__200_ = t_2__200_ | t_2__204_;
  assign t_3__199_ = t_2__199_ | t_2__203_;
  assign t_3__198_ = t_2__198_ | t_2__202_;
  assign t_3__197_ = t_2__197_ | t_2__201_;
  assign t_3__196_ = t_2__196_ | t_2__200_;
  assign t_3__195_ = t_2__195_ | t_2__199_;
  assign t_3__194_ = t_2__194_ | t_2__198_;
  assign t_3__193_ = t_2__193_ | t_2__197_;
  assign t_3__192_ = t_2__192_ | t_2__196_;
  assign t_3__191_ = t_2__191_ | t_2__195_;
  assign t_3__190_ = t_2__190_ | t_2__194_;
  assign t_3__189_ = t_2__189_ | t_2__193_;
  assign t_3__188_ = t_2__188_ | t_2__192_;
  assign t_3__187_ = t_2__187_ | t_2__191_;
  assign t_3__186_ = t_2__186_ | t_2__190_;
  assign t_3__185_ = t_2__185_ | t_2__189_;
  assign t_3__184_ = t_2__184_ | t_2__188_;
  assign t_3__183_ = t_2__183_ | t_2__187_;
  assign t_3__182_ = t_2__182_ | t_2__186_;
  assign t_3__181_ = t_2__181_ | t_2__185_;
  assign t_3__180_ = t_2__180_ | t_2__184_;
  assign t_3__179_ = t_2__179_ | t_2__183_;
  assign t_3__178_ = t_2__178_ | t_2__182_;
  assign t_3__177_ = t_2__177_ | t_2__181_;
  assign t_3__176_ = t_2__176_ | t_2__180_;
  assign t_3__175_ = t_2__175_ | t_2__179_;
  assign t_3__174_ = t_2__174_ | t_2__178_;
  assign t_3__173_ = t_2__173_ | t_2__177_;
  assign t_3__172_ = t_2__172_ | t_2__176_;
  assign t_3__171_ = t_2__171_ | t_2__175_;
  assign t_3__170_ = t_2__170_ | t_2__174_;
  assign t_3__169_ = t_2__169_ | t_2__173_;
  assign t_3__168_ = t_2__168_ | t_2__172_;
  assign t_3__167_ = t_2__167_ | t_2__171_;
  assign t_3__166_ = t_2__166_ | t_2__170_;
  assign t_3__165_ = t_2__165_ | t_2__169_;
  assign t_3__164_ = t_2__164_ | t_2__168_;
  assign t_3__163_ = t_2__163_ | t_2__167_;
  assign t_3__162_ = t_2__162_ | t_2__166_;
  assign t_3__161_ = t_2__161_ | t_2__165_;
  assign t_3__160_ = t_2__160_ | t_2__164_;
  assign t_3__159_ = t_2__159_ | t_2__163_;
  assign t_3__158_ = t_2__158_ | t_2__162_;
  assign t_3__157_ = t_2__157_ | t_2__161_;
  assign t_3__156_ = t_2__156_ | t_2__160_;
  assign t_3__155_ = t_2__155_ | t_2__159_;
  assign t_3__154_ = t_2__154_ | t_2__158_;
  assign t_3__153_ = t_2__153_ | t_2__157_;
  assign t_3__152_ = t_2__152_ | t_2__156_;
  assign t_3__151_ = t_2__151_ | t_2__155_;
  assign t_3__150_ = t_2__150_ | t_2__154_;
  assign t_3__149_ = t_2__149_ | t_2__153_;
  assign t_3__148_ = t_2__148_ | t_2__152_;
  assign t_3__147_ = t_2__147_ | t_2__151_;
  assign t_3__146_ = t_2__146_ | t_2__150_;
  assign t_3__145_ = t_2__145_ | t_2__149_;
  assign t_3__144_ = t_2__144_ | t_2__148_;
  assign t_3__143_ = t_2__143_ | t_2__147_;
  assign t_3__142_ = t_2__142_ | t_2__146_;
  assign t_3__141_ = t_2__141_ | t_2__145_;
  assign t_3__140_ = t_2__140_ | t_2__144_;
  assign t_3__139_ = t_2__139_ | t_2__143_;
  assign t_3__138_ = t_2__138_ | t_2__142_;
  assign t_3__137_ = t_2__137_ | t_2__141_;
  assign t_3__136_ = t_2__136_ | t_2__140_;
  assign t_3__135_ = t_2__135_ | t_2__139_;
  assign t_3__134_ = t_2__134_ | t_2__138_;
  assign t_3__133_ = t_2__133_ | t_2__137_;
  assign t_3__132_ = t_2__132_ | t_2__136_;
  assign t_3__131_ = t_2__131_ | t_2__135_;
  assign t_3__130_ = t_2__130_ | t_2__134_;
  assign t_3__129_ = t_2__129_ | t_2__133_;
  assign t_3__128_ = t_2__128_ | t_2__132_;
  assign t_3__127_ = t_2__127_ | t_2__131_;
  assign t_3__126_ = t_2__126_ | t_2__130_;
  assign t_3__125_ = t_2__125_ | t_2__129_;
  assign t_3__124_ = t_2__124_ | t_2__128_;
  assign t_3__123_ = t_2__123_ | t_2__127_;
  assign t_3__122_ = t_2__122_ | t_2__126_;
  assign t_3__121_ = t_2__121_ | t_2__125_;
  assign t_3__120_ = t_2__120_ | t_2__124_;
  assign t_3__119_ = t_2__119_ | t_2__123_;
  assign t_3__118_ = t_2__118_ | t_2__122_;
  assign t_3__117_ = t_2__117_ | t_2__121_;
  assign t_3__116_ = t_2__116_ | t_2__120_;
  assign t_3__115_ = t_2__115_ | t_2__119_;
  assign t_3__114_ = t_2__114_ | t_2__118_;
  assign t_3__113_ = t_2__113_ | t_2__117_;
  assign t_3__112_ = t_2__112_ | t_2__116_;
  assign t_3__111_ = t_2__111_ | t_2__115_;
  assign t_3__110_ = t_2__110_ | t_2__114_;
  assign t_3__109_ = t_2__109_ | t_2__113_;
  assign t_3__108_ = t_2__108_ | t_2__112_;
  assign t_3__107_ = t_2__107_ | t_2__111_;
  assign t_3__106_ = t_2__106_ | t_2__110_;
  assign t_3__105_ = t_2__105_ | t_2__109_;
  assign t_3__104_ = t_2__104_ | t_2__108_;
  assign t_3__103_ = t_2__103_ | t_2__107_;
  assign t_3__102_ = t_2__102_ | t_2__106_;
  assign t_3__101_ = t_2__101_ | t_2__105_;
  assign t_3__100_ = t_2__100_ | t_2__104_;
  assign t_3__99_ = t_2__99_ | t_2__103_;
  assign t_3__98_ = t_2__98_ | t_2__102_;
  assign t_3__97_ = t_2__97_ | t_2__101_;
  assign t_3__96_ = t_2__96_ | t_2__100_;
  assign t_3__95_ = t_2__95_ | t_2__99_;
  assign t_3__94_ = t_2__94_ | t_2__98_;
  assign t_3__93_ = t_2__93_ | t_2__97_;
  assign t_3__92_ = t_2__92_ | t_2__96_;
  assign t_3__91_ = t_2__91_ | t_2__95_;
  assign t_3__90_ = t_2__90_ | t_2__94_;
  assign t_3__89_ = t_2__89_ | t_2__93_;
  assign t_3__88_ = t_2__88_ | t_2__92_;
  assign t_3__87_ = t_2__87_ | t_2__91_;
  assign t_3__86_ = t_2__86_ | t_2__90_;
  assign t_3__85_ = t_2__85_ | t_2__89_;
  assign t_3__84_ = t_2__84_ | t_2__88_;
  assign t_3__83_ = t_2__83_ | t_2__87_;
  assign t_3__82_ = t_2__82_ | t_2__86_;
  assign t_3__81_ = t_2__81_ | t_2__85_;
  assign t_3__80_ = t_2__80_ | t_2__84_;
  assign t_3__79_ = t_2__79_ | t_2__83_;
  assign t_3__78_ = t_2__78_ | t_2__82_;
  assign t_3__77_ = t_2__77_ | t_2__81_;
  assign t_3__76_ = t_2__76_ | t_2__80_;
  assign t_3__75_ = t_2__75_ | t_2__79_;
  assign t_3__74_ = t_2__74_ | t_2__78_;
  assign t_3__73_ = t_2__73_ | t_2__77_;
  assign t_3__72_ = t_2__72_ | t_2__76_;
  assign t_3__71_ = t_2__71_ | t_2__75_;
  assign t_3__70_ = t_2__70_ | t_2__74_;
  assign t_3__69_ = t_2__69_ | t_2__73_;
  assign t_3__68_ = t_2__68_ | t_2__72_;
  assign t_3__67_ = t_2__67_ | t_2__71_;
  assign t_3__66_ = t_2__66_ | t_2__70_;
  assign t_3__65_ = t_2__65_ | t_2__69_;
  assign t_3__64_ = t_2__64_ | t_2__68_;
  assign t_3__63_ = t_2__63_ | t_2__67_;
  assign t_3__62_ = t_2__62_ | t_2__66_;
  assign t_3__61_ = t_2__61_ | t_2__65_;
  assign t_3__60_ = t_2__60_ | t_2__64_;
  assign t_3__59_ = t_2__59_ | t_2__63_;
  assign t_3__58_ = t_2__58_ | t_2__62_;
  assign t_3__57_ = t_2__57_ | t_2__61_;
  assign t_3__56_ = t_2__56_ | t_2__60_;
  assign t_3__55_ = t_2__55_ | t_2__59_;
  assign t_3__54_ = t_2__54_ | t_2__58_;
  assign t_3__53_ = t_2__53_ | t_2__57_;
  assign t_3__52_ = t_2__52_ | t_2__56_;
  assign t_3__51_ = t_2__51_ | t_2__55_;
  assign t_3__50_ = t_2__50_ | t_2__54_;
  assign t_3__49_ = t_2__49_ | t_2__53_;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__511_ = t_3__511_ | 1'b0;
  assign t_4__510_ = t_3__510_ | 1'b0;
  assign t_4__509_ = t_3__509_ | 1'b0;
  assign t_4__508_ = t_3__508_ | 1'b0;
  assign t_4__507_ = t_3__507_ | 1'b0;
  assign t_4__506_ = t_3__506_ | 1'b0;
  assign t_4__505_ = t_3__505_ | 1'b0;
  assign t_4__504_ = t_3__504_ | 1'b0;
  assign t_4__503_ = t_3__503_ | t_3__511_;
  assign t_4__502_ = t_3__502_ | t_3__510_;
  assign t_4__501_ = t_3__501_ | t_3__509_;
  assign t_4__500_ = t_3__500_ | t_3__508_;
  assign t_4__499_ = t_3__499_ | t_3__507_;
  assign t_4__498_ = t_3__498_ | t_3__506_;
  assign t_4__497_ = t_3__497_ | t_3__505_;
  assign t_4__496_ = t_3__496_ | t_3__504_;
  assign t_4__495_ = t_3__495_ | t_3__503_;
  assign t_4__494_ = t_3__494_ | t_3__502_;
  assign t_4__493_ = t_3__493_ | t_3__501_;
  assign t_4__492_ = t_3__492_ | t_3__500_;
  assign t_4__491_ = t_3__491_ | t_3__499_;
  assign t_4__490_ = t_3__490_ | t_3__498_;
  assign t_4__489_ = t_3__489_ | t_3__497_;
  assign t_4__488_ = t_3__488_ | t_3__496_;
  assign t_4__487_ = t_3__487_ | t_3__495_;
  assign t_4__486_ = t_3__486_ | t_3__494_;
  assign t_4__485_ = t_3__485_ | t_3__493_;
  assign t_4__484_ = t_3__484_ | t_3__492_;
  assign t_4__483_ = t_3__483_ | t_3__491_;
  assign t_4__482_ = t_3__482_ | t_3__490_;
  assign t_4__481_ = t_3__481_ | t_3__489_;
  assign t_4__480_ = t_3__480_ | t_3__488_;
  assign t_4__479_ = t_3__479_ | t_3__487_;
  assign t_4__478_ = t_3__478_ | t_3__486_;
  assign t_4__477_ = t_3__477_ | t_3__485_;
  assign t_4__476_ = t_3__476_ | t_3__484_;
  assign t_4__475_ = t_3__475_ | t_3__483_;
  assign t_4__474_ = t_3__474_ | t_3__482_;
  assign t_4__473_ = t_3__473_ | t_3__481_;
  assign t_4__472_ = t_3__472_ | t_3__480_;
  assign t_4__471_ = t_3__471_ | t_3__479_;
  assign t_4__470_ = t_3__470_ | t_3__478_;
  assign t_4__469_ = t_3__469_ | t_3__477_;
  assign t_4__468_ = t_3__468_ | t_3__476_;
  assign t_4__467_ = t_3__467_ | t_3__475_;
  assign t_4__466_ = t_3__466_ | t_3__474_;
  assign t_4__465_ = t_3__465_ | t_3__473_;
  assign t_4__464_ = t_3__464_ | t_3__472_;
  assign t_4__463_ = t_3__463_ | t_3__471_;
  assign t_4__462_ = t_3__462_ | t_3__470_;
  assign t_4__461_ = t_3__461_ | t_3__469_;
  assign t_4__460_ = t_3__460_ | t_3__468_;
  assign t_4__459_ = t_3__459_ | t_3__467_;
  assign t_4__458_ = t_3__458_ | t_3__466_;
  assign t_4__457_ = t_3__457_ | t_3__465_;
  assign t_4__456_ = t_3__456_ | t_3__464_;
  assign t_4__455_ = t_3__455_ | t_3__463_;
  assign t_4__454_ = t_3__454_ | t_3__462_;
  assign t_4__453_ = t_3__453_ | t_3__461_;
  assign t_4__452_ = t_3__452_ | t_3__460_;
  assign t_4__451_ = t_3__451_ | t_3__459_;
  assign t_4__450_ = t_3__450_ | t_3__458_;
  assign t_4__449_ = t_3__449_ | t_3__457_;
  assign t_4__448_ = t_3__448_ | t_3__456_;
  assign t_4__447_ = t_3__447_ | t_3__455_;
  assign t_4__446_ = t_3__446_ | t_3__454_;
  assign t_4__445_ = t_3__445_ | t_3__453_;
  assign t_4__444_ = t_3__444_ | t_3__452_;
  assign t_4__443_ = t_3__443_ | t_3__451_;
  assign t_4__442_ = t_3__442_ | t_3__450_;
  assign t_4__441_ = t_3__441_ | t_3__449_;
  assign t_4__440_ = t_3__440_ | t_3__448_;
  assign t_4__439_ = t_3__439_ | t_3__447_;
  assign t_4__438_ = t_3__438_ | t_3__446_;
  assign t_4__437_ = t_3__437_ | t_3__445_;
  assign t_4__436_ = t_3__436_ | t_3__444_;
  assign t_4__435_ = t_3__435_ | t_3__443_;
  assign t_4__434_ = t_3__434_ | t_3__442_;
  assign t_4__433_ = t_3__433_ | t_3__441_;
  assign t_4__432_ = t_3__432_ | t_3__440_;
  assign t_4__431_ = t_3__431_ | t_3__439_;
  assign t_4__430_ = t_3__430_ | t_3__438_;
  assign t_4__429_ = t_3__429_ | t_3__437_;
  assign t_4__428_ = t_3__428_ | t_3__436_;
  assign t_4__427_ = t_3__427_ | t_3__435_;
  assign t_4__426_ = t_3__426_ | t_3__434_;
  assign t_4__425_ = t_3__425_ | t_3__433_;
  assign t_4__424_ = t_3__424_ | t_3__432_;
  assign t_4__423_ = t_3__423_ | t_3__431_;
  assign t_4__422_ = t_3__422_ | t_3__430_;
  assign t_4__421_ = t_3__421_ | t_3__429_;
  assign t_4__420_ = t_3__420_ | t_3__428_;
  assign t_4__419_ = t_3__419_ | t_3__427_;
  assign t_4__418_ = t_3__418_ | t_3__426_;
  assign t_4__417_ = t_3__417_ | t_3__425_;
  assign t_4__416_ = t_3__416_ | t_3__424_;
  assign t_4__415_ = t_3__415_ | t_3__423_;
  assign t_4__414_ = t_3__414_ | t_3__422_;
  assign t_4__413_ = t_3__413_ | t_3__421_;
  assign t_4__412_ = t_3__412_ | t_3__420_;
  assign t_4__411_ = t_3__411_ | t_3__419_;
  assign t_4__410_ = t_3__410_ | t_3__418_;
  assign t_4__409_ = t_3__409_ | t_3__417_;
  assign t_4__408_ = t_3__408_ | t_3__416_;
  assign t_4__407_ = t_3__407_ | t_3__415_;
  assign t_4__406_ = t_3__406_ | t_3__414_;
  assign t_4__405_ = t_3__405_ | t_3__413_;
  assign t_4__404_ = t_3__404_ | t_3__412_;
  assign t_4__403_ = t_3__403_ | t_3__411_;
  assign t_4__402_ = t_3__402_ | t_3__410_;
  assign t_4__401_ = t_3__401_ | t_3__409_;
  assign t_4__400_ = t_3__400_ | t_3__408_;
  assign t_4__399_ = t_3__399_ | t_3__407_;
  assign t_4__398_ = t_3__398_ | t_3__406_;
  assign t_4__397_ = t_3__397_ | t_3__405_;
  assign t_4__396_ = t_3__396_ | t_3__404_;
  assign t_4__395_ = t_3__395_ | t_3__403_;
  assign t_4__394_ = t_3__394_ | t_3__402_;
  assign t_4__393_ = t_3__393_ | t_3__401_;
  assign t_4__392_ = t_3__392_ | t_3__400_;
  assign t_4__391_ = t_3__391_ | t_3__399_;
  assign t_4__390_ = t_3__390_ | t_3__398_;
  assign t_4__389_ = t_3__389_ | t_3__397_;
  assign t_4__388_ = t_3__388_ | t_3__396_;
  assign t_4__387_ = t_3__387_ | t_3__395_;
  assign t_4__386_ = t_3__386_ | t_3__394_;
  assign t_4__385_ = t_3__385_ | t_3__393_;
  assign t_4__384_ = t_3__384_ | t_3__392_;
  assign t_4__383_ = t_3__383_ | t_3__391_;
  assign t_4__382_ = t_3__382_ | t_3__390_;
  assign t_4__381_ = t_3__381_ | t_3__389_;
  assign t_4__380_ = t_3__380_ | t_3__388_;
  assign t_4__379_ = t_3__379_ | t_3__387_;
  assign t_4__378_ = t_3__378_ | t_3__386_;
  assign t_4__377_ = t_3__377_ | t_3__385_;
  assign t_4__376_ = t_3__376_ | t_3__384_;
  assign t_4__375_ = t_3__375_ | t_3__383_;
  assign t_4__374_ = t_3__374_ | t_3__382_;
  assign t_4__373_ = t_3__373_ | t_3__381_;
  assign t_4__372_ = t_3__372_ | t_3__380_;
  assign t_4__371_ = t_3__371_ | t_3__379_;
  assign t_4__370_ = t_3__370_ | t_3__378_;
  assign t_4__369_ = t_3__369_ | t_3__377_;
  assign t_4__368_ = t_3__368_ | t_3__376_;
  assign t_4__367_ = t_3__367_ | t_3__375_;
  assign t_4__366_ = t_3__366_ | t_3__374_;
  assign t_4__365_ = t_3__365_ | t_3__373_;
  assign t_4__364_ = t_3__364_ | t_3__372_;
  assign t_4__363_ = t_3__363_ | t_3__371_;
  assign t_4__362_ = t_3__362_ | t_3__370_;
  assign t_4__361_ = t_3__361_ | t_3__369_;
  assign t_4__360_ = t_3__360_ | t_3__368_;
  assign t_4__359_ = t_3__359_ | t_3__367_;
  assign t_4__358_ = t_3__358_ | t_3__366_;
  assign t_4__357_ = t_3__357_ | t_3__365_;
  assign t_4__356_ = t_3__356_ | t_3__364_;
  assign t_4__355_ = t_3__355_ | t_3__363_;
  assign t_4__354_ = t_3__354_ | t_3__362_;
  assign t_4__353_ = t_3__353_ | t_3__361_;
  assign t_4__352_ = t_3__352_ | t_3__360_;
  assign t_4__351_ = t_3__351_ | t_3__359_;
  assign t_4__350_ = t_3__350_ | t_3__358_;
  assign t_4__349_ = t_3__349_ | t_3__357_;
  assign t_4__348_ = t_3__348_ | t_3__356_;
  assign t_4__347_ = t_3__347_ | t_3__355_;
  assign t_4__346_ = t_3__346_ | t_3__354_;
  assign t_4__345_ = t_3__345_ | t_3__353_;
  assign t_4__344_ = t_3__344_ | t_3__352_;
  assign t_4__343_ = t_3__343_ | t_3__351_;
  assign t_4__342_ = t_3__342_ | t_3__350_;
  assign t_4__341_ = t_3__341_ | t_3__349_;
  assign t_4__340_ = t_3__340_ | t_3__348_;
  assign t_4__339_ = t_3__339_ | t_3__347_;
  assign t_4__338_ = t_3__338_ | t_3__346_;
  assign t_4__337_ = t_3__337_ | t_3__345_;
  assign t_4__336_ = t_3__336_ | t_3__344_;
  assign t_4__335_ = t_3__335_ | t_3__343_;
  assign t_4__334_ = t_3__334_ | t_3__342_;
  assign t_4__333_ = t_3__333_ | t_3__341_;
  assign t_4__332_ = t_3__332_ | t_3__340_;
  assign t_4__331_ = t_3__331_ | t_3__339_;
  assign t_4__330_ = t_3__330_ | t_3__338_;
  assign t_4__329_ = t_3__329_ | t_3__337_;
  assign t_4__328_ = t_3__328_ | t_3__336_;
  assign t_4__327_ = t_3__327_ | t_3__335_;
  assign t_4__326_ = t_3__326_ | t_3__334_;
  assign t_4__325_ = t_3__325_ | t_3__333_;
  assign t_4__324_ = t_3__324_ | t_3__332_;
  assign t_4__323_ = t_3__323_ | t_3__331_;
  assign t_4__322_ = t_3__322_ | t_3__330_;
  assign t_4__321_ = t_3__321_ | t_3__329_;
  assign t_4__320_ = t_3__320_ | t_3__328_;
  assign t_4__319_ = t_3__319_ | t_3__327_;
  assign t_4__318_ = t_3__318_ | t_3__326_;
  assign t_4__317_ = t_3__317_ | t_3__325_;
  assign t_4__316_ = t_3__316_ | t_3__324_;
  assign t_4__315_ = t_3__315_ | t_3__323_;
  assign t_4__314_ = t_3__314_ | t_3__322_;
  assign t_4__313_ = t_3__313_ | t_3__321_;
  assign t_4__312_ = t_3__312_ | t_3__320_;
  assign t_4__311_ = t_3__311_ | t_3__319_;
  assign t_4__310_ = t_3__310_ | t_3__318_;
  assign t_4__309_ = t_3__309_ | t_3__317_;
  assign t_4__308_ = t_3__308_ | t_3__316_;
  assign t_4__307_ = t_3__307_ | t_3__315_;
  assign t_4__306_ = t_3__306_ | t_3__314_;
  assign t_4__305_ = t_3__305_ | t_3__313_;
  assign t_4__304_ = t_3__304_ | t_3__312_;
  assign t_4__303_ = t_3__303_ | t_3__311_;
  assign t_4__302_ = t_3__302_ | t_3__310_;
  assign t_4__301_ = t_3__301_ | t_3__309_;
  assign t_4__300_ = t_3__300_ | t_3__308_;
  assign t_4__299_ = t_3__299_ | t_3__307_;
  assign t_4__298_ = t_3__298_ | t_3__306_;
  assign t_4__297_ = t_3__297_ | t_3__305_;
  assign t_4__296_ = t_3__296_ | t_3__304_;
  assign t_4__295_ = t_3__295_ | t_3__303_;
  assign t_4__294_ = t_3__294_ | t_3__302_;
  assign t_4__293_ = t_3__293_ | t_3__301_;
  assign t_4__292_ = t_3__292_ | t_3__300_;
  assign t_4__291_ = t_3__291_ | t_3__299_;
  assign t_4__290_ = t_3__290_ | t_3__298_;
  assign t_4__289_ = t_3__289_ | t_3__297_;
  assign t_4__288_ = t_3__288_ | t_3__296_;
  assign t_4__287_ = t_3__287_ | t_3__295_;
  assign t_4__286_ = t_3__286_ | t_3__294_;
  assign t_4__285_ = t_3__285_ | t_3__293_;
  assign t_4__284_ = t_3__284_ | t_3__292_;
  assign t_4__283_ = t_3__283_ | t_3__291_;
  assign t_4__282_ = t_3__282_ | t_3__290_;
  assign t_4__281_ = t_3__281_ | t_3__289_;
  assign t_4__280_ = t_3__280_ | t_3__288_;
  assign t_4__279_ = t_3__279_ | t_3__287_;
  assign t_4__278_ = t_3__278_ | t_3__286_;
  assign t_4__277_ = t_3__277_ | t_3__285_;
  assign t_4__276_ = t_3__276_ | t_3__284_;
  assign t_4__275_ = t_3__275_ | t_3__283_;
  assign t_4__274_ = t_3__274_ | t_3__282_;
  assign t_4__273_ = t_3__273_ | t_3__281_;
  assign t_4__272_ = t_3__272_ | t_3__280_;
  assign t_4__271_ = t_3__271_ | t_3__279_;
  assign t_4__270_ = t_3__270_ | t_3__278_;
  assign t_4__269_ = t_3__269_ | t_3__277_;
  assign t_4__268_ = t_3__268_ | t_3__276_;
  assign t_4__267_ = t_3__267_ | t_3__275_;
  assign t_4__266_ = t_3__266_ | t_3__274_;
  assign t_4__265_ = t_3__265_ | t_3__273_;
  assign t_4__264_ = t_3__264_ | t_3__272_;
  assign t_4__263_ = t_3__263_ | t_3__271_;
  assign t_4__262_ = t_3__262_ | t_3__270_;
  assign t_4__261_ = t_3__261_ | t_3__269_;
  assign t_4__260_ = t_3__260_ | t_3__268_;
  assign t_4__259_ = t_3__259_ | t_3__267_;
  assign t_4__258_ = t_3__258_ | t_3__266_;
  assign t_4__257_ = t_3__257_ | t_3__265_;
  assign t_4__256_ = t_3__256_ | t_3__264_;
  assign t_4__255_ = t_3__255_ | t_3__263_;
  assign t_4__254_ = t_3__254_ | t_3__262_;
  assign t_4__253_ = t_3__253_ | t_3__261_;
  assign t_4__252_ = t_3__252_ | t_3__260_;
  assign t_4__251_ = t_3__251_ | t_3__259_;
  assign t_4__250_ = t_3__250_ | t_3__258_;
  assign t_4__249_ = t_3__249_ | t_3__257_;
  assign t_4__248_ = t_3__248_ | t_3__256_;
  assign t_4__247_ = t_3__247_ | t_3__255_;
  assign t_4__246_ = t_3__246_ | t_3__254_;
  assign t_4__245_ = t_3__245_ | t_3__253_;
  assign t_4__244_ = t_3__244_ | t_3__252_;
  assign t_4__243_ = t_3__243_ | t_3__251_;
  assign t_4__242_ = t_3__242_ | t_3__250_;
  assign t_4__241_ = t_3__241_ | t_3__249_;
  assign t_4__240_ = t_3__240_ | t_3__248_;
  assign t_4__239_ = t_3__239_ | t_3__247_;
  assign t_4__238_ = t_3__238_ | t_3__246_;
  assign t_4__237_ = t_3__237_ | t_3__245_;
  assign t_4__236_ = t_3__236_ | t_3__244_;
  assign t_4__235_ = t_3__235_ | t_3__243_;
  assign t_4__234_ = t_3__234_ | t_3__242_;
  assign t_4__233_ = t_3__233_ | t_3__241_;
  assign t_4__232_ = t_3__232_ | t_3__240_;
  assign t_4__231_ = t_3__231_ | t_3__239_;
  assign t_4__230_ = t_3__230_ | t_3__238_;
  assign t_4__229_ = t_3__229_ | t_3__237_;
  assign t_4__228_ = t_3__228_ | t_3__236_;
  assign t_4__227_ = t_3__227_ | t_3__235_;
  assign t_4__226_ = t_3__226_ | t_3__234_;
  assign t_4__225_ = t_3__225_ | t_3__233_;
  assign t_4__224_ = t_3__224_ | t_3__232_;
  assign t_4__223_ = t_3__223_ | t_3__231_;
  assign t_4__222_ = t_3__222_ | t_3__230_;
  assign t_4__221_ = t_3__221_ | t_3__229_;
  assign t_4__220_ = t_3__220_ | t_3__228_;
  assign t_4__219_ = t_3__219_ | t_3__227_;
  assign t_4__218_ = t_3__218_ | t_3__226_;
  assign t_4__217_ = t_3__217_ | t_3__225_;
  assign t_4__216_ = t_3__216_ | t_3__224_;
  assign t_4__215_ = t_3__215_ | t_3__223_;
  assign t_4__214_ = t_3__214_ | t_3__222_;
  assign t_4__213_ = t_3__213_ | t_3__221_;
  assign t_4__212_ = t_3__212_ | t_3__220_;
  assign t_4__211_ = t_3__211_ | t_3__219_;
  assign t_4__210_ = t_3__210_ | t_3__218_;
  assign t_4__209_ = t_3__209_ | t_3__217_;
  assign t_4__208_ = t_3__208_ | t_3__216_;
  assign t_4__207_ = t_3__207_ | t_3__215_;
  assign t_4__206_ = t_3__206_ | t_3__214_;
  assign t_4__205_ = t_3__205_ | t_3__213_;
  assign t_4__204_ = t_3__204_ | t_3__212_;
  assign t_4__203_ = t_3__203_ | t_3__211_;
  assign t_4__202_ = t_3__202_ | t_3__210_;
  assign t_4__201_ = t_3__201_ | t_3__209_;
  assign t_4__200_ = t_3__200_ | t_3__208_;
  assign t_4__199_ = t_3__199_ | t_3__207_;
  assign t_4__198_ = t_3__198_ | t_3__206_;
  assign t_4__197_ = t_3__197_ | t_3__205_;
  assign t_4__196_ = t_3__196_ | t_3__204_;
  assign t_4__195_ = t_3__195_ | t_3__203_;
  assign t_4__194_ = t_3__194_ | t_3__202_;
  assign t_4__193_ = t_3__193_ | t_3__201_;
  assign t_4__192_ = t_3__192_ | t_3__200_;
  assign t_4__191_ = t_3__191_ | t_3__199_;
  assign t_4__190_ = t_3__190_ | t_3__198_;
  assign t_4__189_ = t_3__189_ | t_3__197_;
  assign t_4__188_ = t_3__188_ | t_3__196_;
  assign t_4__187_ = t_3__187_ | t_3__195_;
  assign t_4__186_ = t_3__186_ | t_3__194_;
  assign t_4__185_ = t_3__185_ | t_3__193_;
  assign t_4__184_ = t_3__184_ | t_3__192_;
  assign t_4__183_ = t_3__183_ | t_3__191_;
  assign t_4__182_ = t_3__182_ | t_3__190_;
  assign t_4__181_ = t_3__181_ | t_3__189_;
  assign t_4__180_ = t_3__180_ | t_3__188_;
  assign t_4__179_ = t_3__179_ | t_3__187_;
  assign t_4__178_ = t_3__178_ | t_3__186_;
  assign t_4__177_ = t_3__177_ | t_3__185_;
  assign t_4__176_ = t_3__176_ | t_3__184_;
  assign t_4__175_ = t_3__175_ | t_3__183_;
  assign t_4__174_ = t_3__174_ | t_3__182_;
  assign t_4__173_ = t_3__173_ | t_3__181_;
  assign t_4__172_ = t_3__172_ | t_3__180_;
  assign t_4__171_ = t_3__171_ | t_3__179_;
  assign t_4__170_ = t_3__170_ | t_3__178_;
  assign t_4__169_ = t_3__169_ | t_3__177_;
  assign t_4__168_ = t_3__168_ | t_3__176_;
  assign t_4__167_ = t_3__167_ | t_3__175_;
  assign t_4__166_ = t_3__166_ | t_3__174_;
  assign t_4__165_ = t_3__165_ | t_3__173_;
  assign t_4__164_ = t_3__164_ | t_3__172_;
  assign t_4__163_ = t_3__163_ | t_3__171_;
  assign t_4__162_ = t_3__162_ | t_3__170_;
  assign t_4__161_ = t_3__161_ | t_3__169_;
  assign t_4__160_ = t_3__160_ | t_3__168_;
  assign t_4__159_ = t_3__159_ | t_3__167_;
  assign t_4__158_ = t_3__158_ | t_3__166_;
  assign t_4__157_ = t_3__157_ | t_3__165_;
  assign t_4__156_ = t_3__156_ | t_3__164_;
  assign t_4__155_ = t_3__155_ | t_3__163_;
  assign t_4__154_ = t_3__154_ | t_3__162_;
  assign t_4__153_ = t_3__153_ | t_3__161_;
  assign t_4__152_ = t_3__152_ | t_3__160_;
  assign t_4__151_ = t_3__151_ | t_3__159_;
  assign t_4__150_ = t_3__150_ | t_3__158_;
  assign t_4__149_ = t_3__149_ | t_3__157_;
  assign t_4__148_ = t_3__148_ | t_3__156_;
  assign t_4__147_ = t_3__147_ | t_3__155_;
  assign t_4__146_ = t_3__146_ | t_3__154_;
  assign t_4__145_ = t_3__145_ | t_3__153_;
  assign t_4__144_ = t_3__144_ | t_3__152_;
  assign t_4__143_ = t_3__143_ | t_3__151_;
  assign t_4__142_ = t_3__142_ | t_3__150_;
  assign t_4__141_ = t_3__141_ | t_3__149_;
  assign t_4__140_ = t_3__140_ | t_3__148_;
  assign t_4__139_ = t_3__139_ | t_3__147_;
  assign t_4__138_ = t_3__138_ | t_3__146_;
  assign t_4__137_ = t_3__137_ | t_3__145_;
  assign t_4__136_ = t_3__136_ | t_3__144_;
  assign t_4__135_ = t_3__135_ | t_3__143_;
  assign t_4__134_ = t_3__134_ | t_3__142_;
  assign t_4__133_ = t_3__133_ | t_3__141_;
  assign t_4__132_ = t_3__132_ | t_3__140_;
  assign t_4__131_ = t_3__131_ | t_3__139_;
  assign t_4__130_ = t_3__130_ | t_3__138_;
  assign t_4__129_ = t_3__129_ | t_3__137_;
  assign t_4__128_ = t_3__128_ | t_3__136_;
  assign t_4__127_ = t_3__127_ | t_3__135_;
  assign t_4__126_ = t_3__126_ | t_3__134_;
  assign t_4__125_ = t_3__125_ | t_3__133_;
  assign t_4__124_ = t_3__124_ | t_3__132_;
  assign t_4__123_ = t_3__123_ | t_3__131_;
  assign t_4__122_ = t_3__122_ | t_3__130_;
  assign t_4__121_ = t_3__121_ | t_3__129_;
  assign t_4__120_ = t_3__120_ | t_3__128_;
  assign t_4__119_ = t_3__119_ | t_3__127_;
  assign t_4__118_ = t_3__118_ | t_3__126_;
  assign t_4__117_ = t_3__117_ | t_3__125_;
  assign t_4__116_ = t_3__116_ | t_3__124_;
  assign t_4__115_ = t_3__115_ | t_3__123_;
  assign t_4__114_ = t_3__114_ | t_3__122_;
  assign t_4__113_ = t_3__113_ | t_3__121_;
  assign t_4__112_ = t_3__112_ | t_3__120_;
  assign t_4__111_ = t_3__111_ | t_3__119_;
  assign t_4__110_ = t_3__110_ | t_3__118_;
  assign t_4__109_ = t_3__109_ | t_3__117_;
  assign t_4__108_ = t_3__108_ | t_3__116_;
  assign t_4__107_ = t_3__107_ | t_3__115_;
  assign t_4__106_ = t_3__106_ | t_3__114_;
  assign t_4__105_ = t_3__105_ | t_3__113_;
  assign t_4__104_ = t_3__104_ | t_3__112_;
  assign t_4__103_ = t_3__103_ | t_3__111_;
  assign t_4__102_ = t_3__102_ | t_3__110_;
  assign t_4__101_ = t_3__101_ | t_3__109_;
  assign t_4__100_ = t_3__100_ | t_3__108_;
  assign t_4__99_ = t_3__99_ | t_3__107_;
  assign t_4__98_ = t_3__98_ | t_3__106_;
  assign t_4__97_ = t_3__97_ | t_3__105_;
  assign t_4__96_ = t_3__96_ | t_3__104_;
  assign t_4__95_ = t_3__95_ | t_3__103_;
  assign t_4__94_ = t_3__94_ | t_3__102_;
  assign t_4__93_ = t_3__93_ | t_3__101_;
  assign t_4__92_ = t_3__92_ | t_3__100_;
  assign t_4__91_ = t_3__91_ | t_3__99_;
  assign t_4__90_ = t_3__90_ | t_3__98_;
  assign t_4__89_ = t_3__89_ | t_3__97_;
  assign t_4__88_ = t_3__88_ | t_3__96_;
  assign t_4__87_ = t_3__87_ | t_3__95_;
  assign t_4__86_ = t_3__86_ | t_3__94_;
  assign t_4__85_ = t_3__85_ | t_3__93_;
  assign t_4__84_ = t_3__84_ | t_3__92_;
  assign t_4__83_ = t_3__83_ | t_3__91_;
  assign t_4__82_ = t_3__82_ | t_3__90_;
  assign t_4__81_ = t_3__81_ | t_3__89_;
  assign t_4__80_ = t_3__80_ | t_3__88_;
  assign t_4__79_ = t_3__79_ | t_3__87_;
  assign t_4__78_ = t_3__78_ | t_3__86_;
  assign t_4__77_ = t_3__77_ | t_3__85_;
  assign t_4__76_ = t_3__76_ | t_3__84_;
  assign t_4__75_ = t_3__75_ | t_3__83_;
  assign t_4__74_ = t_3__74_ | t_3__82_;
  assign t_4__73_ = t_3__73_ | t_3__81_;
  assign t_4__72_ = t_3__72_ | t_3__80_;
  assign t_4__71_ = t_3__71_ | t_3__79_;
  assign t_4__70_ = t_3__70_ | t_3__78_;
  assign t_4__69_ = t_3__69_ | t_3__77_;
  assign t_4__68_ = t_3__68_ | t_3__76_;
  assign t_4__67_ = t_3__67_ | t_3__75_;
  assign t_4__66_ = t_3__66_ | t_3__74_;
  assign t_4__65_ = t_3__65_ | t_3__73_;
  assign t_4__64_ = t_3__64_ | t_3__72_;
  assign t_4__63_ = t_3__63_ | t_3__71_;
  assign t_4__62_ = t_3__62_ | t_3__70_;
  assign t_4__61_ = t_3__61_ | t_3__69_;
  assign t_4__60_ = t_3__60_ | t_3__68_;
  assign t_4__59_ = t_3__59_ | t_3__67_;
  assign t_4__58_ = t_3__58_ | t_3__66_;
  assign t_4__57_ = t_3__57_ | t_3__65_;
  assign t_4__56_ = t_3__56_ | t_3__64_;
  assign t_4__55_ = t_3__55_ | t_3__63_;
  assign t_4__54_ = t_3__54_ | t_3__62_;
  assign t_4__53_ = t_3__53_ | t_3__61_;
  assign t_4__52_ = t_3__52_ | t_3__60_;
  assign t_4__51_ = t_3__51_ | t_3__59_;
  assign t_4__50_ = t_3__50_ | t_3__58_;
  assign t_4__49_ = t_3__49_ | t_3__57_;
  assign t_4__48_ = t_3__48_ | t_3__56_;
  assign t_4__47_ = t_3__47_ | t_3__55_;
  assign t_4__46_ = t_3__46_ | t_3__54_;
  assign t_4__45_ = t_3__45_ | t_3__53_;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__511_ = t_4__511_ | 1'b0;
  assign t_5__510_ = t_4__510_ | 1'b0;
  assign t_5__509_ = t_4__509_ | 1'b0;
  assign t_5__508_ = t_4__508_ | 1'b0;
  assign t_5__507_ = t_4__507_ | 1'b0;
  assign t_5__506_ = t_4__506_ | 1'b0;
  assign t_5__505_ = t_4__505_ | 1'b0;
  assign t_5__504_ = t_4__504_ | 1'b0;
  assign t_5__503_ = t_4__503_ | 1'b0;
  assign t_5__502_ = t_4__502_ | 1'b0;
  assign t_5__501_ = t_4__501_ | 1'b0;
  assign t_5__500_ = t_4__500_ | 1'b0;
  assign t_5__499_ = t_4__499_ | 1'b0;
  assign t_5__498_ = t_4__498_ | 1'b0;
  assign t_5__497_ = t_4__497_ | 1'b0;
  assign t_5__496_ = t_4__496_ | 1'b0;
  assign t_5__495_ = t_4__495_ | t_4__511_;
  assign t_5__494_ = t_4__494_ | t_4__510_;
  assign t_5__493_ = t_4__493_ | t_4__509_;
  assign t_5__492_ = t_4__492_ | t_4__508_;
  assign t_5__491_ = t_4__491_ | t_4__507_;
  assign t_5__490_ = t_4__490_ | t_4__506_;
  assign t_5__489_ = t_4__489_ | t_4__505_;
  assign t_5__488_ = t_4__488_ | t_4__504_;
  assign t_5__487_ = t_4__487_ | t_4__503_;
  assign t_5__486_ = t_4__486_ | t_4__502_;
  assign t_5__485_ = t_4__485_ | t_4__501_;
  assign t_5__484_ = t_4__484_ | t_4__500_;
  assign t_5__483_ = t_4__483_ | t_4__499_;
  assign t_5__482_ = t_4__482_ | t_4__498_;
  assign t_5__481_ = t_4__481_ | t_4__497_;
  assign t_5__480_ = t_4__480_ | t_4__496_;
  assign t_5__479_ = t_4__479_ | t_4__495_;
  assign t_5__478_ = t_4__478_ | t_4__494_;
  assign t_5__477_ = t_4__477_ | t_4__493_;
  assign t_5__476_ = t_4__476_ | t_4__492_;
  assign t_5__475_ = t_4__475_ | t_4__491_;
  assign t_5__474_ = t_4__474_ | t_4__490_;
  assign t_5__473_ = t_4__473_ | t_4__489_;
  assign t_5__472_ = t_4__472_ | t_4__488_;
  assign t_5__471_ = t_4__471_ | t_4__487_;
  assign t_5__470_ = t_4__470_ | t_4__486_;
  assign t_5__469_ = t_4__469_ | t_4__485_;
  assign t_5__468_ = t_4__468_ | t_4__484_;
  assign t_5__467_ = t_4__467_ | t_4__483_;
  assign t_5__466_ = t_4__466_ | t_4__482_;
  assign t_5__465_ = t_4__465_ | t_4__481_;
  assign t_5__464_ = t_4__464_ | t_4__480_;
  assign t_5__463_ = t_4__463_ | t_4__479_;
  assign t_5__462_ = t_4__462_ | t_4__478_;
  assign t_5__461_ = t_4__461_ | t_4__477_;
  assign t_5__460_ = t_4__460_ | t_4__476_;
  assign t_5__459_ = t_4__459_ | t_4__475_;
  assign t_5__458_ = t_4__458_ | t_4__474_;
  assign t_5__457_ = t_4__457_ | t_4__473_;
  assign t_5__456_ = t_4__456_ | t_4__472_;
  assign t_5__455_ = t_4__455_ | t_4__471_;
  assign t_5__454_ = t_4__454_ | t_4__470_;
  assign t_5__453_ = t_4__453_ | t_4__469_;
  assign t_5__452_ = t_4__452_ | t_4__468_;
  assign t_5__451_ = t_4__451_ | t_4__467_;
  assign t_5__450_ = t_4__450_ | t_4__466_;
  assign t_5__449_ = t_4__449_ | t_4__465_;
  assign t_5__448_ = t_4__448_ | t_4__464_;
  assign t_5__447_ = t_4__447_ | t_4__463_;
  assign t_5__446_ = t_4__446_ | t_4__462_;
  assign t_5__445_ = t_4__445_ | t_4__461_;
  assign t_5__444_ = t_4__444_ | t_4__460_;
  assign t_5__443_ = t_4__443_ | t_4__459_;
  assign t_5__442_ = t_4__442_ | t_4__458_;
  assign t_5__441_ = t_4__441_ | t_4__457_;
  assign t_5__440_ = t_4__440_ | t_4__456_;
  assign t_5__439_ = t_4__439_ | t_4__455_;
  assign t_5__438_ = t_4__438_ | t_4__454_;
  assign t_5__437_ = t_4__437_ | t_4__453_;
  assign t_5__436_ = t_4__436_ | t_4__452_;
  assign t_5__435_ = t_4__435_ | t_4__451_;
  assign t_5__434_ = t_4__434_ | t_4__450_;
  assign t_5__433_ = t_4__433_ | t_4__449_;
  assign t_5__432_ = t_4__432_ | t_4__448_;
  assign t_5__431_ = t_4__431_ | t_4__447_;
  assign t_5__430_ = t_4__430_ | t_4__446_;
  assign t_5__429_ = t_4__429_ | t_4__445_;
  assign t_5__428_ = t_4__428_ | t_4__444_;
  assign t_5__427_ = t_4__427_ | t_4__443_;
  assign t_5__426_ = t_4__426_ | t_4__442_;
  assign t_5__425_ = t_4__425_ | t_4__441_;
  assign t_5__424_ = t_4__424_ | t_4__440_;
  assign t_5__423_ = t_4__423_ | t_4__439_;
  assign t_5__422_ = t_4__422_ | t_4__438_;
  assign t_5__421_ = t_4__421_ | t_4__437_;
  assign t_5__420_ = t_4__420_ | t_4__436_;
  assign t_5__419_ = t_4__419_ | t_4__435_;
  assign t_5__418_ = t_4__418_ | t_4__434_;
  assign t_5__417_ = t_4__417_ | t_4__433_;
  assign t_5__416_ = t_4__416_ | t_4__432_;
  assign t_5__415_ = t_4__415_ | t_4__431_;
  assign t_5__414_ = t_4__414_ | t_4__430_;
  assign t_5__413_ = t_4__413_ | t_4__429_;
  assign t_5__412_ = t_4__412_ | t_4__428_;
  assign t_5__411_ = t_4__411_ | t_4__427_;
  assign t_5__410_ = t_4__410_ | t_4__426_;
  assign t_5__409_ = t_4__409_ | t_4__425_;
  assign t_5__408_ = t_4__408_ | t_4__424_;
  assign t_5__407_ = t_4__407_ | t_4__423_;
  assign t_5__406_ = t_4__406_ | t_4__422_;
  assign t_5__405_ = t_4__405_ | t_4__421_;
  assign t_5__404_ = t_4__404_ | t_4__420_;
  assign t_5__403_ = t_4__403_ | t_4__419_;
  assign t_5__402_ = t_4__402_ | t_4__418_;
  assign t_5__401_ = t_4__401_ | t_4__417_;
  assign t_5__400_ = t_4__400_ | t_4__416_;
  assign t_5__399_ = t_4__399_ | t_4__415_;
  assign t_5__398_ = t_4__398_ | t_4__414_;
  assign t_5__397_ = t_4__397_ | t_4__413_;
  assign t_5__396_ = t_4__396_ | t_4__412_;
  assign t_5__395_ = t_4__395_ | t_4__411_;
  assign t_5__394_ = t_4__394_ | t_4__410_;
  assign t_5__393_ = t_4__393_ | t_4__409_;
  assign t_5__392_ = t_4__392_ | t_4__408_;
  assign t_5__391_ = t_4__391_ | t_4__407_;
  assign t_5__390_ = t_4__390_ | t_4__406_;
  assign t_5__389_ = t_4__389_ | t_4__405_;
  assign t_5__388_ = t_4__388_ | t_4__404_;
  assign t_5__387_ = t_4__387_ | t_4__403_;
  assign t_5__386_ = t_4__386_ | t_4__402_;
  assign t_5__385_ = t_4__385_ | t_4__401_;
  assign t_5__384_ = t_4__384_ | t_4__400_;
  assign t_5__383_ = t_4__383_ | t_4__399_;
  assign t_5__382_ = t_4__382_ | t_4__398_;
  assign t_5__381_ = t_4__381_ | t_4__397_;
  assign t_5__380_ = t_4__380_ | t_4__396_;
  assign t_5__379_ = t_4__379_ | t_4__395_;
  assign t_5__378_ = t_4__378_ | t_4__394_;
  assign t_5__377_ = t_4__377_ | t_4__393_;
  assign t_5__376_ = t_4__376_ | t_4__392_;
  assign t_5__375_ = t_4__375_ | t_4__391_;
  assign t_5__374_ = t_4__374_ | t_4__390_;
  assign t_5__373_ = t_4__373_ | t_4__389_;
  assign t_5__372_ = t_4__372_ | t_4__388_;
  assign t_5__371_ = t_4__371_ | t_4__387_;
  assign t_5__370_ = t_4__370_ | t_4__386_;
  assign t_5__369_ = t_4__369_ | t_4__385_;
  assign t_5__368_ = t_4__368_ | t_4__384_;
  assign t_5__367_ = t_4__367_ | t_4__383_;
  assign t_5__366_ = t_4__366_ | t_4__382_;
  assign t_5__365_ = t_4__365_ | t_4__381_;
  assign t_5__364_ = t_4__364_ | t_4__380_;
  assign t_5__363_ = t_4__363_ | t_4__379_;
  assign t_5__362_ = t_4__362_ | t_4__378_;
  assign t_5__361_ = t_4__361_ | t_4__377_;
  assign t_5__360_ = t_4__360_ | t_4__376_;
  assign t_5__359_ = t_4__359_ | t_4__375_;
  assign t_5__358_ = t_4__358_ | t_4__374_;
  assign t_5__357_ = t_4__357_ | t_4__373_;
  assign t_5__356_ = t_4__356_ | t_4__372_;
  assign t_5__355_ = t_4__355_ | t_4__371_;
  assign t_5__354_ = t_4__354_ | t_4__370_;
  assign t_5__353_ = t_4__353_ | t_4__369_;
  assign t_5__352_ = t_4__352_ | t_4__368_;
  assign t_5__351_ = t_4__351_ | t_4__367_;
  assign t_5__350_ = t_4__350_ | t_4__366_;
  assign t_5__349_ = t_4__349_ | t_4__365_;
  assign t_5__348_ = t_4__348_ | t_4__364_;
  assign t_5__347_ = t_4__347_ | t_4__363_;
  assign t_5__346_ = t_4__346_ | t_4__362_;
  assign t_5__345_ = t_4__345_ | t_4__361_;
  assign t_5__344_ = t_4__344_ | t_4__360_;
  assign t_5__343_ = t_4__343_ | t_4__359_;
  assign t_5__342_ = t_4__342_ | t_4__358_;
  assign t_5__341_ = t_4__341_ | t_4__357_;
  assign t_5__340_ = t_4__340_ | t_4__356_;
  assign t_5__339_ = t_4__339_ | t_4__355_;
  assign t_5__338_ = t_4__338_ | t_4__354_;
  assign t_5__337_ = t_4__337_ | t_4__353_;
  assign t_5__336_ = t_4__336_ | t_4__352_;
  assign t_5__335_ = t_4__335_ | t_4__351_;
  assign t_5__334_ = t_4__334_ | t_4__350_;
  assign t_5__333_ = t_4__333_ | t_4__349_;
  assign t_5__332_ = t_4__332_ | t_4__348_;
  assign t_5__331_ = t_4__331_ | t_4__347_;
  assign t_5__330_ = t_4__330_ | t_4__346_;
  assign t_5__329_ = t_4__329_ | t_4__345_;
  assign t_5__328_ = t_4__328_ | t_4__344_;
  assign t_5__327_ = t_4__327_ | t_4__343_;
  assign t_5__326_ = t_4__326_ | t_4__342_;
  assign t_5__325_ = t_4__325_ | t_4__341_;
  assign t_5__324_ = t_4__324_ | t_4__340_;
  assign t_5__323_ = t_4__323_ | t_4__339_;
  assign t_5__322_ = t_4__322_ | t_4__338_;
  assign t_5__321_ = t_4__321_ | t_4__337_;
  assign t_5__320_ = t_4__320_ | t_4__336_;
  assign t_5__319_ = t_4__319_ | t_4__335_;
  assign t_5__318_ = t_4__318_ | t_4__334_;
  assign t_5__317_ = t_4__317_ | t_4__333_;
  assign t_5__316_ = t_4__316_ | t_4__332_;
  assign t_5__315_ = t_4__315_ | t_4__331_;
  assign t_5__314_ = t_4__314_ | t_4__330_;
  assign t_5__313_ = t_4__313_ | t_4__329_;
  assign t_5__312_ = t_4__312_ | t_4__328_;
  assign t_5__311_ = t_4__311_ | t_4__327_;
  assign t_5__310_ = t_4__310_ | t_4__326_;
  assign t_5__309_ = t_4__309_ | t_4__325_;
  assign t_5__308_ = t_4__308_ | t_4__324_;
  assign t_5__307_ = t_4__307_ | t_4__323_;
  assign t_5__306_ = t_4__306_ | t_4__322_;
  assign t_5__305_ = t_4__305_ | t_4__321_;
  assign t_5__304_ = t_4__304_ | t_4__320_;
  assign t_5__303_ = t_4__303_ | t_4__319_;
  assign t_5__302_ = t_4__302_ | t_4__318_;
  assign t_5__301_ = t_4__301_ | t_4__317_;
  assign t_5__300_ = t_4__300_ | t_4__316_;
  assign t_5__299_ = t_4__299_ | t_4__315_;
  assign t_5__298_ = t_4__298_ | t_4__314_;
  assign t_5__297_ = t_4__297_ | t_4__313_;
  assign t_5__296_ = t_4__296_ | t_4__312_;
  assign t_5__295_ = t_4__295_ | t_4__311_;
  assign t_5__294_ = t_4__294_ | t_4__310_;
  assign t_5__293_ = t_4__293_ | t_4__309_;
  assign t_5__292_ = t_4__292_ | t_4__308_;
  assign t_5__291_ = t_4__291_ | t_4__307_;
  assign t_5__290_ = t_4__290_ | t_4__306_;
  assign t_5__289_ = t_4__289_ | t_4__305_;
  assign t_5__288_ = t_4__288_ | t_4__304_;
  assign t_5__287_ = t_4__287_ | t_4__303_;
  assign t_5__286_ = t_4__286_ | t_4__302_;
  assign t_5__285_ = t_4__285_ | t_4__301_;
  assign t_5__284_ = t_4__284_ | t_4__300_;
  assign t_5__283_ = t_4__283_ | t_4__299_;
  assign t_5__282_ = t_4__282_ | t_4__298_;
  assign t_5__281_ = t_4__281_ | t_4__297_;
  assign t_5__280_ = t_4__280_ | t_4__296_;
  assign t_5__279_ = t_4__279_ | t_4__295_;
  assign t_5__278_ = t_4__278_ | t_4__294_;
  assign t_5__277_ = t_4__277_ | t_4__293_;
  assign t_5__276_ = t_4__276_ | t_4__292_;
  assign t_5__275_ = t_4__275_ | t_4__291_;
  assign t_5__274_ = t_4__274_ | t_4__290_;
  assign t_5__273_ = t_4__273_ | t_4__289_;
  assign t_5__272_ = t_4__272_ | t_4__288_;
  assign t_5__271_ = t_4__271_ | t_4__287_;
  assign t_5__270_ = t_4__270_ | t_4__286_;
  assign t_5__269_ = t_4__269_ | t_4__285_;
  assign t_5__268_ = t_4__268_ | t_4__284_;
  assign t_5__267_ = t_4__267_ | t_4__283_;
  assign t_5__266_ = t_4__266_ | t_4__282_;
  assign t_5__265_ = t_4__265_ | t_4__281_;
  assign t_5__264_ = t_4__264_ | t_4__280_;
  assign t_5__263_ = t_4__263_ | t_4__279_;
  assign t_5__262_ = t_4__262_ | t_4__278_;
  assign t_5__261_ = t_4__261_ | t_4__277_;
  assign t_5__260_ = t_4__260_ | t_4__276_;
  assign t_5__259_ = t_4__259_ | t_4__275_;
  assign t_5__258_ = t_4__258_ | t_4__274_;
  assign t_5__257_ = t_4__257_ | t_4__273_;
  assign t_5__256_ = t_4__256_ | t_4__272_;
  assign t_5__255_ = t_4__255_ | t_4__271_;
  assign t_5__254_ = t_4__254_ | t_4__270_;
  assign t_5__253_ = t_4__253_ | t_4__269_;
  assign t_5__252_ = t_4__252_ | t_4__268_;
  assign t_5__251_ = t_4__251_ | t_4__267_;
  assign t_5__250_ = t_4__250_ | t_4__266_;
  assign t_5__249_ = t_4__249_ | t_4__265_;
  assign t_5__248_ = t_4__248_ | t_4__264_;
  assign t_5__247_ = t_4__247_ | t_4__263_;
  assign t_5__246_ = t_4__246_ | t_4__262_;
  assign t_5__245_ = t_4__245_ | t_4__261_;
  assign t_5__244_ = t_4__244_ | t_4__260_;
  assign t_5__243_ = t_4__243_ | t_4__259_;
  assign t_5__242_ = t_4__242_ | t_4__258_;
  assign t_5__241_ = t_4__241_ | t_4__257_;
  assign t_5__240_ = t_4__240_ | t_4__256_;
  assign t_5__239_ = t_4__239_ | t_4__255_;
  assign t_5__238_ = t_4__238_ | t_4__254_;
  assign t_5__237_ = t_4__237_ | t_4__253_;
  assign t_5__236_ = t_4__236_ | t_4__252_;
  assign t_5__235_ = t_4__235_ | t_4__251_;
  assign t_5__234_ = t_4__234_ | t_4__250_;
  assign t_5__233_ = t_4__233_ | t_4__249_;
  assign t_5__232_ = t_4__232_ | t_4__248_;
  assign t_5__231_ = t_4__231_ | t_4__247_;
  assign t_5__230_ = t_4__230_ | t_4__246_;
  assign t_5__229_ = t_4__229_ | t_4__245_;
  assign t_5__228_ = t_4__228_ | t_4__244_;
  assign t_5__227_ = t_4__227_ | t_4__243_;
  assign t_5__226_ = t_4__226_ | t_4__242_;
  assign t_5__225_ = t_4__225_ | t_4__241_;
  assign t_5__224_ = t_4__224_ | t_4__240_;
  assign t_5__223_ = t_4__223_ | t_4__239_;
  assign t_5__222_ = t_4__222_ | t_4__238_;
  assign t_5__221_ = t_4__221_ | t_4__237_;
  assign t_5__220_ = t_4__220_ | t_4__236_;
  assign t_5__219_ = t_4__219_ | t_4__235_;
  assign t_5__218_ = t_4__218_ | t_4__234_;
  assign t_5__217_ = t_4__217_ | t_4__233_;
  assign t_5__216_ = t_4__216_ | t_4__232_;
  assign t_5__215_ = t_4__215_ | t_4__231_;
  assign t_5__214_ = t_4__214_ | t_4__230_;
  assign t_5__213_ = t_4__213_ | t_4__229_;
  assign t_5__212_ = t_4__212_ | t_4__228_;
  assign t_5__211_ = t_4__211_ | t_4__227_;
  assign t_5__210_ = t_4__210_ | t_4__226_;
  assign t_5__209_ = t_4__209_ | t_4__225_;
  assign t_5__208_ = t_4__208_ | t_4__224_;
  assign t_5__207_ = t_4__207_ | t_4__223_;
  assign t_5__206_ = t_4__206_ | t_4__222_;
  assign t_5__205_ = t_4__205_ | t_4__221_;
  assign t_5__204_ = t_4__204_ | t_4__220_;
  assign t_5__203_ = t_4__203_ | t_4__219_;
  assign t_5__202_ = t_4__202_ | t_4__218_;
  assign t_5__201_ = t_4__201_ | t_4__217_;
  assign t_5__200_ = t_4__200_ | t_4__216_;
  assign t_5__199_ = t_4__199_ | t_4__215_;
  assign t_5__198_ = t_4__198_ | t_4__214_;
  assign t_5__197_ = t_4__197_ | t_4__213_;
  assign t_5__196_ = t_4__196_ | t_4__212_;
  assign t_5__195_ = t_4__195_ | t_4__211_;
  assign t_5__194_ = t_4__194_ | t_4__210_;
  assign t_5__193_ = t_4__193_ | t_4__209_;
  assign t_5__192_ = t_4__192_ | t_4__208_;
  assign t_5__191_ = t_4__191_ | t_4__207_;
  assign t_5__190_ = t_4__190_ | t_4__206_;
  assign t_5__189_ = t_4__189_ | t_4__205_;
  assign t_5__188_ = t_4__188_ | t_4__204_;
  assign t_5__187_ = t_4__187_ | t_4__203_;
  assign t_5__186_ = t_4__186_ | t_4__202_;
  assign t_5__185_ = t_4__185_ | t_4__201_;
  assign t_5__184_ = t_4__184_ | t_4__200_;
  assign t_5__183_ = t_4__183_ | t_4__199_;
  assign t_5__182_ = t_4__182_ | t_4__198_;
  assign t_5__181_ = t_4__181_ | t_4__197_;
  assign t_5__180_ = t_4__180_ | t_4__196_;
  assign t_5__179_ = t_4__179_ | t_4__195_;
  assign t_5__178_ = t_4__178_ | t_4__194_;
  assign t_5__177_ = t_4__177_ | t_4__193_;
  assign t_5__176_ = t_4__176_ | t_4__192_;
  assign t_5__175_ = t_4__175_ | t_4__191_;
  assign t_5__174_ = t_4__174_ | t_4__190_;
  assign t_5__173_ = t_4__173_ | t_4__189_;
  assign t_5__172_ = t_4__172_ | t_4__188_;
  assign t_5__171_ = t_4__171_ | t_4__187_;
  assign t_5__170_ = t_4__170_ | t_4__186_;
  assign t_5__169_ = t_4__169_ | t_4__185_;
  assign t_5__168_ = t_4__168_ | t_4__184_;
  assign t_5__167_ = t_4__167_ | t_4__183_;
  assign t_5__166_ = t_4__166_ | t_4__182_;
  assign t_5__165_ = t_4__165_ | t_4__181_;
  assign t_5__164_ = t_4__164_ | t_4__180_;
  assign t_5__163_ = t_4__163_ | t_4__179_;
  assign t_5__162_ = t_4__162_ | t_4__178_;
  assign t_5__161_ = t_4__161_ | t_4__177_;
  assign t_5__160_ = t_4__160_ | t_4__176_;
  assign t_5__159_ = t_4__159_ | t_4__175_;
  assign t_5__158_ = t_4__158_ | t_4__174_;
  assign t_5__157_ = t_4__157_ | t_4__173_;
  assign t_5__156_ = t_4__156_ | t_4__172_;
  assign t_5__155_ = t_4__155_ | t_4__171_;
  assign t_5__154_ = t_4__154_ | t_4__170_;
  assign t_5__153_ = t_4__153_ | t_4__169_;
  assign t_5__152_ = t_4__152_ | t_4__168_;
  assign t_5__151_ = t_4__151_ | t_4__167_;
  assign t_5__150_ = t_4__150_ | t_4__166_;
  assign t_5__149_ = t_4__149_ | t_4__165_;
  assign t_5__148_ = t_4__148_ | t_4__164_;
  assign t_5__147_ = t_4__147_ | t_4__163_;
  assign t_5__146_ = t_4__146_ | t_4__162_;
  assign t_5__145_ = t_4__145_ | t_4__161_;
  assign t_5__144_ = t_4__144_ | t_4__160_;
  assign t_5__143_ = t_4__143_ | t_4__159_;
  assign t_5__142_ = t_4__142_ | t_4__158_;
  assign t_5__141_ = t_4__141_ | t_4__157_;
  assign t_5__140_ = t_4__140_ | t_4__156_;
  assign t_5__139_ = t_4__139_ | t_4__155_;
  assign t_5__138_ = t_4__138_ | t_4__154_;
  assign t_5__137_ = t_4__137_ | t_4__153_;
  assign t_5__136_ = t_4__136_ | t_4__152_;
  assign t_5__135_ = t_4__135_ | t_4__151_;
  assign t_5__134_ = t_4__134_ | t_4__150_;
  assign t_5__133_ = t_4__133_ | t_4__149_;
  assign t_5__132_ = t_4__132_ | t_4__148_;
  assign t_5__131_ = t_4__131_ | t_4__147_;
  assign t_5__130_ = t_4__130_ | t_4__146_;
  assign t_5__129_ = t_4__129_ | t_4__145_;
  assign t_5__128_ = t_4__128_ | t_4__144_;
  assign t_5__127_ = t_4__127_ | t_4__143_;
  assign t_5__126_ = t_4__126_ | t_4__142_;
  assign t_5__125_ = t_4__125_ | t_4__141_;
  assign t_5__124_ = t_4__124_ | t_4__140_;
  assign t_5__123_ = t_4__123_ | t_4__139_;
  assign t_5__122_ = t_4__122_ | t_4__138_;
  assign t_5__121_ = t_4__121_ | t_4__137_;
  assign t_5__120_ = t_4__120_ | t_4__136_;
  assign t_5__119_ = t_4__119_ | t_4__135_;
  assign t_5__118_ = t_4__118_ | t_4__134_;
  assign t_5__117_ = t_4__117_ | t_4__133_;
  assign t_5__116_ = t_4__116_ | t_4__132_;
  assign t_5__115_ = t_4__115_ | t_4__131_;
  assign t_5__114_ = t_4__114_ | t_4__130_;
  assign t_5__113_ = t_4__113_ | t_4__129_;
  assign t_5__112_ = t_4__112_ | t_4__128_;
  assign t_5__111_ = t_4__111_ | t_4__127_;
  assign t_5__110_ = t_4__110_ | t_4__126_;
  assign t_5__109_ = t_4__109_ | t_4__125_;
  assign t_5__108_ = t_4__108_ | t_4__124_;
  assign t_5__107_ = t_4__107_ | t_4__123_;
  assign t_5__106_ = t_4__106_ | t_4__122_;
  assign t_5__105_ = t_4__105_ | t_4__121_;
  assign t_5__104_ = t_4__104_ | t_4__120_;
  assign t_5__103_ = t_4__103_ | t_4__119_;
  assign t_5__102_ = t_4__102_ | t_4__118_;
  assign t_5__101_ = t_4__101_ | t_4__117_;
  assign t_5__100_ = t_4__100_ | t_4__116_;
  assign t_5__99_ = t_4__99_ | t_4__115_;
  assign t_5__98_ = t_4__98_ | t_4__114_;
  assign t_5__97_ = t_4__97_ | t_4__113_;
  assign t_5__96_ = t_4__96_ | t_4__112_;
  assign t_5__95_ = t_4__95_ | t_4__111_;
  assign t_5__94_ = t_4__94_ | t_4__110_;
  assign t_5__93_ = t_4__93_ | t_4__109_;
  assign t_5__92_ = t_4__92_ | t_4__108_;
  assign t_5__91_ = t_4__91_ | t_4__107_;
  assign t_5__90_ = t_4__90_ | t_4__106_;
  assign t_5__89_ = t_4__89_ | t_4__105_;
  assign t_5__88_ = t_4__88_ | t_4__104_;
  assign t_5__87_ = t_4__87_ | t_4__103_;
  assign t_5__86_ = t_4__86_ | t_4__102_;
  assign t_5__85_ = t_4__85_ | t_4__101_;
  assign t_5__84_ = t_4__84_ | t_4__100_;
  assign t_5__83_ = t_4__83_ | t_4__99_;
  assign t_5__82_ = t_4__82_ | t_4__98_;
  assign t_5__81_ = t_4__81_ | t_4__97_;
  assign t_5__80_ = t_4__80_ | t_4__96_;
  assign t_5__79_ = t_4__79_ | t_4__95_;
  assign t_5__78_ = t_4__78_ | t_4__94_;
  assign t_5__77_ = t_4__77_ | t_4__93_;
  assign t_5__76_ = t_4__76_ | t_4__92_;
  assign t_5__75_ = t_4__75_ | t_4__91_;
  assign t_5__74_ = t_4__74_ | t_4__90_;
  assign t_5__73_ = t_4__73_ | t_4__89_;
  assign t_5__72_ = t_4__72_ | t_4__88_;
  assign t_5__71_ = t_4__71_ | t_4__87_;
  assign t_5__70_ = t_4__70_ | t_4__86_;
  assign t_5__69_ = t_4__69_ | t_4__85_;
  assign t_5__68_ = t_4__68_ | t_4__84_;
  assign t_5__67_ = t_4__67_ | t_4__83_;
  assign t_5__66_ = t_4__66_ | t_4__82_;
  assign t_5__65_ = t_4__65_ | t_4__81_;
  assign t_5__64_ = t_4__64_ | t_4__80_;
  assign t_5__63_ = t_4__63_ | t_4__79_;
  assign t_5__62_ = t_4__62_ | t_4__78_;
  assign t_5__61_ = t_4__61_ | t_4__77_;
  assign t_5__60_ = t_4__60_ | t_4__76_;
  assign t_5__59_ = t_4__59_ | t_4__75_;
  assign t_5__58_ = t_4__58_ | t_4__74_;
  assign t_5__57_ = t_4__57_ | t_4__73_;
  assign t_5__56_ = t_4__56_ | t_4__72_;
  assign t_5__55_ = t_4__55_ | t_4__71_;
  assign t_5__54_ = t_4__54_ | t_4__70_;
  assign t_5__53_ = t_4__53_ | t_4__69_;
  assign t_5__52_ = t_4__52_ | t_4__68_;
  assign t_5__51_ = t_4__51_ | t_4__67_;
  assign t_5__50_ = t_4__50_ | t_4__66_;
  assign t_5__49_ = t_4__49_ | t_4__65_;
  assign t_5__48_ = t_4__48_ | t_4__64_;
  assign t_5__47_ = t_4__47_ | t_4__63_;
  assign t_5__46_ = t_4__46_ | t_4__62_;
  assign t_5__45_ = t_4__45_ | t_4__61_;
  assign t_5__44_ = t_4__44_ | t_4__60_;
  assign t_5__43_ = t_4__43_ | t_4__59_;
  assign t_5__42_ = t_4__42_ | t_4__58_;
  assign t_5__41_ = t_4__41_ | t_4__57_;
  assign t_5__40_ = t_4__40_ | t_4__56_;
  assign t_5__39_ = t_4__39_ | t_4__55_;
  assign t_5__38_ = t_4__38_ | t_4__54_;
  assign t_5__37_ = t_4__37_ | t_4__53_;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign t_6__511_ = t_5__511_ | 1'b0;
  assign t_6__510_ = t_5__510_ | 1'b0;
  assign t_6__509_ = t_5__509_ | 1'b0;
  assign t_6__508_ = t_5__508_ | 1'b0;
  assign t_6__507_ = t_5__507_ | 1'b0;
  assign t_6__506_ = t_5__506_ | 1'b0;
  assign t_6__505_ = t_5__505_ | 1'b0;
  assign t_6__504_ = t_5__504_ | 1'b0;
  assign t_6__503_ = t_5__503_ | 1'b0;
  assign t_6__502_ = t_5__502_ | 1'b0;
  assign t_6__501_ = t_5__501_ | 1'b0;
  assign t_6__500_ = t_5__500_ | 1'b0;
  assign t_6__499_ = t_5__499_ | 1'b0;
  assign t_6__498_ = t_5__498_ | 1'b0;
  assign t_6__497_ = t_5__497_ | 1'b0;
  assign t_6__496_ = t_5__496_ | 1'b0;
  assign t_6__495_ = t_5__495_ | 1'b0;
  assign t_6__494_ = t_5__494_ | 1'b0;
  assign t_6__493_ = t_5__493_ | 1'b0;
  assign t_6__492_ = t_5__492_ | 1'b0;
  assign t_6__491_ = t_5__491_ | 1'b0;
  assign t_6__490_ = t_5__490_ | 1'b0;
  assign t_6__489_ = t_5__489_ | 1'b0;
  assign t_6__488_ = t_5__488_ | 1'b0;
  assign t_6__487_ = t_5__487_ | 1'b0;
  assign t_6__486_ = t_5__486_ | 1'b0;
  assign t_6__485_ = t_5__485_ | 1'b0;
  assign t_6__484_ = t_5__484_ | 1'b0;
  assign t_6__483_ = t_5__483_ | 1'b0;
  assign t_6__482_ = t_5__482_ | 1'b0;
  assign t_6__481_ = t_5__481_ | 1'b0;
  assign t_6__480_ = t_5__480_ | 1'b0;
  assign t_6__479_ = t_5__479_ | t_5__511_;
  assign t_6__478_ = t_5__478_ | t_5__510_;
  assign t_6__477_ = t_5__477_ | t_5__509_;
  assign t_6__476_ = t_5__476_ | t_5__508_;
  assign t_6__475_ = t_5__475_ | t_5__507_;
  assign t_6__474_ = t_5__474_ | t_5__506_;
  assign t_6__473_ = t_5__473_ | t_5__505_;
  assign t_6__472_ = t_5__472_ | t_5__504_;
  assign t_6__471_ = t_5__471_ | t_5__503_;
  assign t_6__470_ = t_5__470_ | t_5__502_;
  assign t_6__469_ = t_5__469_ | t_5__501_;
  assign t_6__468_ = t_5__468_ | t_5__500_;
  assign t_6__467_ = t_5__467_ | t_5__499_;
  assign t_6__466_ = t_5__466_ | t_5__498_;
  assign t_6__465_ = t_5__465_ | t_5__497_;
  assign t_6__464_ = t_5__464_ | t_5__496_;
  assign t_6__463_ = t_5__463_ | t_5__495_;
  assign t_6__462_ = t_5__462_ | t_5__494_;
  assign t_6__461_ = t_5__461_ | t_5__493_;
  assign t_6__460_ = t_5__460_ | t_5__492_;
  assign t_6__459_ = t_5__459_ | t_5__491_;
  assign t_6__458_ = t_5__458_ | t_5__490_;
  assign t_6__457_ = t_5__457_ | t_5__489_;
  assign t_6__456_ = t_5__456_ | t_5__488_;
  assign t_6__455_ = t_5__455_ | t_5__487_;
  assign t_6__454_ = t_5__454_ | t_5__486_;
  assign t_6__453_ = t_5__453_ | t_5__485_;
  assign t_6__452_ = t_5__452_ | t_5__484_;
  assign t_6__451_ = t_5__451_ | t_5__483_;
  assign t_6__450_ = t_5__450_ | t_5__482_;
  assign t_6__449_ = t_5__449_ | t_5__481_;
  assign t_6__448_ = t_5__448_ | t_5__480_;
  assign t_6__447_ = t_5__447_ | t_5__479_;
  assign t_6__446_ = t_5__446_ | t_5__478_;
  assign t_6__445_ = t_5__445_ | t_5__477_;
  assign t_6__444_ = t_5__444_ | t_5__476_;
  assign t_6__443_ = t_5__443_ | t_5__475_;
  assign t_6__442_ = t_5__442_ | t_5__474_;
  assign t_6__441_ = t_5__441_ | t_5__473_;
  assign t_6__440_ = t_5__440_ | t_5__472_;
  assign t_6__439_ = t_5__439_ | t_5__471_;
  assign t_6__438_ = t_5__438_ | t_5__470_;
  assign t_6__437_ = t_5__437_ | t_5__469_;
  assign t_6__436_ = t_5__436_ | t_5__468_;
  assign t_6__435_ = t_5__435_ | t_5__467_;
  assign t_6__434_ = t_5__434_ | t_5__466_;
  assign t_6__433_ = t_5__433_ | t_5__465_;
  assign t_6__432_ = t_5__432_ | t_5__464_;
  assign t_6__431_ = t_5__431_ | t_5__463_;
  assign t_6__430_ = t_5__430_ | t_5__462_;
  assign t_6__429_ = t_5__429_ | t_5__461_;
  assign t_6__428_ = t_5__428_ | t_5__460_;
  assign t_6__427_ = t_5__427_ | t_5__459_;
  assign t_6__426_ = t_5__426_ | t_5__458_;
  assign t_6__425_ = t_5__425_ | t_5__457_;
  assign t_6__424_ = t_5__424_ | t_5__456_;
  assign t_6__423_ = t_5__423_ | t_5__455_;
  assign t_6__422_ = t_5__422_ | t_5__454_;
  assign t_6__421_ = t_5__421_ | t_5__453_;
  assign t_6__420_ = t_5__420_ | t_5__452_;
  assign t_6__419_ = t_5__419_ | t_5__451_;
  assign t_6__418_ = t_5__418_ | t_5__450_;
  assign t_6__417_ = t_5__417_ | t_5__449_;
  assign t_6__416_ = t_5__416_ | t_5__448_;
  assign t_6__415_ = t_5__415_ | t_5__447_;
  assign t_6__414_ = t_5__414_ | t_5__446_;
  assign t_6__413_ = t_5__413_ | t_5__445_;
  assign t_6__412_ = t_5__412_ | t_5__444_;
  assign t_6__411_ = t_5__411_ | t_5__443_;
  assign t_6__410_ = t_5__410_ | t_5__442_;
  assign t_6__409_ = t_5__409_ | t_5__441_;
  assign t_6__408_ = t_5__408_ | t_5__440_;
  assign t_6__407_ = t_5__407_ | t_5__439_;
  assign t_6__406_ = t_5__406_ | t_5__438_;
  assign t_6__405_ = t_5__405_ | t_5__437_;
  assign t_6__404_ = t_5__404_ | t_5__436_;
  assign t_6__403_ = t_5__403_ | t_5__435_;
  assign t_6__402_ = t_5__402_ | t_5__434_;
  assign t_6__401_ = t_5__401_ | t_5__433_;
  assign t_6__400_ = t_5__400_ | t_5__432_;
  assign t_6__399_ = t_5__399_ | t_5__431_;
  assign t_6__398_ = t_5__398_ | t_5__430_;
  assign t_6__397_ = t_5__397_ | t_5__429_;
  assign t_6__396_ = t_5__396_ | t_5__428_;
  assign t_6__395_ = t_5__395_ | t_5__427_;
  assign t_6__394_ = t_5__394_ | t_5__426_;
  assign t_6__393_ = t_5__393_ | t_5__425_;
  assign t_6__392_ = t_5__392_ | t_5__424_;
  assign t_6__391_ = t_5__391_ | t_5__423_;
  assign t_6__390_ = t_5__390_ | t_5__422_;
  assign t_6__389_ = t_5__389_ | t_5__421_;
  assign t_6__388_ = t_5__388_ | t_5__420_;
  assign t_6__387_ = t_5__387_ | t_5__419_;
  assign t_6__386_ = t_5__386_ | t_5__418_;
  assign t_6__385_ = t_5__385_ | t_5__417_;
  assign t_6__384_ = t_5__384_ | t_5__416_;
  assign t_6__383_ = t_5__383_ | t_5__415_;
  assign t_6__382_ = t_5__382_ | t_5__414_;
  assign t_6__381_ = t_5__381_ | t_5__413_;
  assign t_6__380_ = t_5__380_ | t_5__412_;
  assign t_6__379_ = t_5__379_ | t_5__411_;
  assign t_6__378_ = t_5__378_ | t_5__410_;
  assign t_6__377_ = t_5__377_ | t_5__409_;
  assign t_6__376_ = t_5__376_ | t_5__408_;
  assign t_6__375_ = t_5__375_ | t_5__407_;
  assign t_6__374_ = t_5__374_ | t_5__406_;
  assign t_6__373_ = t_5__373_ | t_5__405_;
  assign t_6__372_ = t_5__372_ | t_5__404_;
  assign t_6__371_ = t_5__371_ | t_5__403_;
  assign t_6__370_ = t_5__370_ | t_5__402_;
  assign t_6__369_ = t_5__369_ | t_5__401_;
  assign t_6__368_ = t_5__368_ | t_5__400_;
  assign t_6__367_ = t_5__367_ | t_5__399_;
  assign t_6__366_ = t_5__366_ | t_5__398_;
  assign t_6__365_ = t_5__365_ | t_5__397_;
  assign t_6__364_ = t_5__364_ | t_5__396_;
  assign t_6__363_ = t_5__363_ | t_5__395_;
  assign t_6__362_ = t_5__362_ | t_5__394_;
  assign t_6__361_ = t_5__361_ | t_5__393_;
  assign t_6__360_ = t_5__360_ | t_5__392_;
  assign t_6__359_ = t_5__359_ | t_5__391_;
  assign t_6__358_ = t_5__358_ | t_5__390_;
  assign t_6__357_ = t_5__357_ | t_5__389_;
  assign t_6__356_ = t_5__356_ | t_5__388_;
  assign t_6__355_ = t_5__355_ | t_5__387_;
  assign t_6__354_ = t_5__354_ | t_5__386_;
  assign t_6__353_ = t_5__353_ | t_5__385_;
  assign t_6__352_ = t_5__352_ | t_5__384_;
  assign t_6__351_ = t_5__351_ | t_5__383_;
  assign t_6__350_ = t_5__350_ | t_5__382_;
  assign t_6__349_ = t_5__349_ | t_5__381_;
  assign t_6__348_ = t_5__348_ | t_5__380_;
  assign t_6__347_ = t_5__347_ | t_5__379_;
  assign t_6__346_ = t_5__346_ | t_5__378_;
  assign t_6__345_ = t_5__345_ | t_5__377_;
  assign t_6__344_ = t_5__344_ | t_5__376_;
  assign t_6__343_ = t_5__343_ | t_5__375_;
  assign t_6__342_ = t_5__342_ | t_5__374_;
  assign t_6__341_ = t_5__341_ | t_5__373_;
  assign t_6__340_ = t_5__340_ | t_5__372_;
  assign t_6__339_ = t_5__339_ | t_5__371_;
  assign t_6__338_ = t_5__338_ | t_5__370_;
  assign t_6__337_ = t_5__337_ | t_5__369_;
  assign t_6__336_ = t_5__336_ | t_5__368_;
  assign t_6__335_ = t_5__335_ | t_5__367_;
  assign t_6__334_ = t_5__334_ | t_5__366_;
  assign t_6__333_ = t_5__333_ | t_5__365_;
  assign t_6__332_ = t_5__332_ | t_5__364_;
  assign t_6__331_ = t_5__331_ | t_5__363_;
  assign t_6__330_ = t_5__330_ | t_5__362_;
  assign t_6__329_ = t_5__329_ | t_5__361_;
  assign t_6__328_ = t_5__328_ | t_5__360_;
  assign t_6__327_ = t_5__327_ | t_5__359_;
  assign t_6__326_ = t_5__326_ | t_5__358_;
  assign t_6__325_ = t_5__325_ | t_5__357_;
  assign t_6__324_ = t_5__324_ | t_5__356_;
  assign t_6__323_ = t_5__323_ | t_5__355_;
  assign t_6__322_ = t_5__322_ | t_5__354_;
  assign t_6__321_ = t_5__321_ | t_5__353_;
  assign t_6__320_ = t_5__320_ | t_5__352_;
  assign t_6__319_ = t_5__319_ | t_5__351_;
  assign t_6__318_ = t_5__318_ | t_5__350_;
  assign t_6__317_ = t_5__317_ | t_5__349_;
  assign t_6__316_ = t_5__316_ | t_5__348_;
  assign t_6__315_ = t_5__315_ | t_5__347_;
  assign t_6__314_ = t_5__314_ | t_5__346_;
  assign t_6__313_ = t_5__313_ | t_5__345_;
  assign t_6__312_ = t_5__312_ | t_5__344_;
  assign t_6__311_ = t_5__311_ | t_5__343_;
  assign t_6__310_ = t_5__310_ | t_5__342_;
  assign t_6__309_ = t_5__309_ | t_5__341_;
  assign t_6__308_ = t_5__308_ | t_5__340_;
  assign t_6__307_ = t_5__307_ | t_5__339_;
  assign t_6__306_ = t_5__306_ | t_5__338_;
  assign t_6__305_ = t_5__305_ | t_5__337_;
  assign t_6__304_ = t_5__304_ | t_5__336_;
  assign t_6__303_ = t_5__303_ | t_5__335_;
  assign t_6__302_ = t_5__302_ | t_5__334_;
  assign t_6__301_ = t_5__301_ | t_5__333_;
  assign t_6__300_ = t_5__300_ | t_5__332_;
  assign t_6__299_ = t_5__299_ | t_5__331_;
  assign t_6__298_ = t_5__298_ | t_5__330_;
  assign t_6__297_ = t_5__297_ | t_5__329_;
  assign t_6__296_ = t_5__296_ | t_5__328_;
  assign t_6__295_ = t_5__295_ | t_5__327_;
  assign t_6__294_ = t_5__294_ | t_5__326_;
  assign t_6__293_ = t_5__293_ | t_5__325_;
  assign t_6__292_ = t_5__292_ | t_5__324_;
  assign t_6__291_ = t_5__291_ | t_5__323_;
  assign t_6__290_ = t_5__290_ | t_5__322_;
  assign t_6__289_ = t_5__289_ | t_5__321_;
  assign t_6__288_ = t_5__288_ | t_5__320_;
  assign t_6__287_ = t_5__287_ | t_5__319_;
  assign t_6__286_ = t_5__286_ | t_5__318_;
  assign t_6__285_ = t_5__285_ | t_5__317_;
  assign t_6__284_ = t_5__284_ | t_5__316_;
  assign t_6__283_ = t_5__283_ | t_5__315_;
  assign t_6__282_ = t_5__282_ | t_5__314_;
  assign t_6__281_ = t_5__281_ | t_5__313_;
  assign t_6__280_ = t_5__280_ | t_5__312_;
  assign t_6__279_ = t_5__279_ | t_5__311_;
  assign t_6__278_ = t_5__278_ | t_5__310_;
  assign t_6__277_ = t_5__277_ | t_5__309_;
  assign t_6__276_ = t_5__276_ | t_5__308_;
  assign t_6__275_ = t_5__275_ | t_5__307_;
  assign t_6__274_ = t_5__274_ | t_5__306_;
  assign t_6__273_ = t_5__273_ | t_5__305_;
  assign t_6__272_ = t_5__272_ | t_5__304_;
  assign t_6__271_ = t_5__271_ | t_5__303_;
  assign t_6__270_ = t_5__270_ | t_5__302_;
  assign t_6__269_ = t_5__269_ | t_5__301_;
  assign t_6__268_ = t_5__268_ | t_5__300_;
  assign t_6__267_ = t_5__267_ | t_5__299_;
  assign t_6__266_ = t_5__266_ | t_5__298_;
  assign t_6__265_ = t_5__265_ | t_5__297_;
  assign t_6__264_ = t_5__264_ | t_5__296_;
  assign t_6__263_ = t_5__263_ | t_5__295_;
  assign t_6__262_ = t_5__262_ | t_5__294_;
  assign t_6__261_ = t_5__261_ | t_5__293_;
  assign t_6__260_ = t_5__260_ | t_5__292_;
  assign t_6__259_ = t_5__259_ | t_5__291_;
  assign t_6__258_ = t_5__258_ | t_5__290_;
  assign t_6__257_ = t_5__257_ | t_5__289_;
  assign t_6__256_ = t_5__256_ | t_5__288_;
  assign t_6__255_ = t_5__255_ | t_5__287_;
  assign t_6__254_ = t_5__254_ | t_5__286_;
  assign t_6__253_ = t_5__253_ | t_5__285_;
  assign t_6__252_ = t_5__252_ | t_5__284_;
  assign t_6__251_ = t_5__251_ | t_5__283_;
  assign t_6__250_ = t_5__250_ | t_5__282_;
  assign t_6__249_ = t_5__249_ | t_5__281_;
  assign t_6__248_ = t_5__248_ | t_5__280_;
  assign t_6__247_ = t_5__247_ | t_5__279_;
  assign t_6__246_ = t_5__246_ | t_5__278_;
  assign t_6__245_ = t_5__245_ | t_5__277_;
  assign t_6__244_ = t_5__244_ | t_5__276_;
  assign t_6__243_ = t_5__243_ | t_5__275_;
  assign t_6__242_ = t_5__242_ | t_5__274_;
  assign t_6__241_ = t_5__241_ | t_5__273_;
  assign t_6__240_ = t_5__240_ | t_5__272_;
  assign t_6__239_ = t_5__239_ | t_5__271_;
  assign t_6__238_ = t_5__238_ | t_5__270_;
  assign t_6__237_ = t_5__237_ | t_5__269_;
  assign t_6__236_ = t_5__236_ | t_5__268_;
  assign t_6__235_ = t_5__235_ | t_5__267_;
  assign t_6__234_ = t_5__234_ | t_5__266_;
  assign t_6__233_ = t_5__233_ | t_5__265_;
  assign t_6__232_ = t_5__232_ | t_5__264_;
  assign t_6__231_ = t_5__231_ | t_5__263_;
  assign t_6__230_ = t_5__230_ | t_5__262_;
  assign t_6__229_ = t_5__229_ | t_5__261_;
  assign t_6__228_ = t_5__228_ | t_5__260_;
  assign t_6__227_ = t_5__227_ | t_5__259_;
  assign t_6__226_ = t_5__226_ | t_5__258_;
  assign t_6__225_ = t_5__225_ | t_5__257_;
  assign t_6__224_ = t_5__224_ | t_5__256_;
  assign t_6__223_ = t_5__223_ | t_5__255_;
  assign t_6__222_ = t_5__222_ | t_5__254_;
  assign t_6__221_ = t_5__221_ | t_5__253_;
  assign t_6__220_ = t_5__220_ | t_5__252_;
  assign t_6__219_ = t_5__219_ | t_5__251_;
  assign t_6__218_ = t_5__218_ | t_5__250_;
  assign t_6__217_ = t_5__217_ | t_5__249_;
  assign t_6__216_ = t_5__216_ | t_5__248_;
  assign t_6__215_ = t_5__215_ | t_5__247_;
  assign t_6__214_ = t_5__214_ | t_5__246_;
  assign t_6__213_ = t_5__213_ | t_5__245_;
  assign t_6__212_ = t_5__212_ | t_5__244_;
  assign t_6__211_ = t_5__211_ | t_5__243_;
  assign t_6__210_ = t_5__210_ | t_5__242_;
  assign t_6__209_ = t_5__209_ | t_5__241_;
  assign t_6__208_ = t_5__208_ | t_5__240_;
  assign t_6__207_ = t_5__207_ | t_5__239_;
  assign t_6__206_ = t_5__206_ | t_5__238_;
  assign t_6__205_ = t_5__205_ | t_5__237_;
  assign t_6__204_ = t_5__204_ | t_5__236_;
  assign t_6__203_ = t_5__203_ | t_5__235_;
  assign t_6__202_ = t_5__202_ | t_5__234_;
  assign t_6__201_ = t_5__201_ | t_5__233_;
  assign t_6__200_ = t_5__200_ | t_5__232_;
  assign t_6__199_ = t_5__199_ | t_5__231_;
  assign t_6__198_ = t_5__198_ | t_5__230_;
  assign t_6__197_ = t_5__197_ | t_5__229_;
  assign t_6__196_ = t_5__196_ | t_5__228_;
  assign t_6__195_ = t_5__195_ | t_5__227_;
  assign t_6__194_ = t_5__194_ | t_5__226_;
  assign t_6__193_ = t_5__193_ | t_5__225_;
  assign t_6__192_ = t_5__192_ | t_5__224_;
  assign t_6__191_ = t_5__191_ | t_5__223_;
  assign t_6__190_ = t_5__190_ | t_5__222_;
  assign t_6__189_ = t_5__189_ | t_5__221_;
  assign t_6__188_ = t_5__188_ | t_5__220_;
  assign t_6__187_ = t_5__187_ | t_5__219_;
  assign t_6__186_ = t_5__186_ | t_5__218_;
  assign t_6__185_ = t_5__185_ | t_5__217_;
  assign t_6__184_ = t_5__184_ | t_5__216_;
  assign t_6__183_ = t_5__183_ | t_5__215_;
  assign t_6__182_ = t_5__182_ | t_5__214_;
  assign t_6__181_ = t_5__181_ | t_5__213_;
  assign t_6__180_ = t_5__180_ | t_5__212_;
  assign t_6__179_ = t_5__179_ | t_5__211_;
  assign t_6__178_ = t_5__178_ | t_5__210_;
  assign t_6__177_ = t_5__177_ | t_5__209_;
  assign t_6__176_ = t_5__176_ | t_5__208_;
  assign t_6__175_ = t_5__175_ | t_5__207_;
  assign t_6__174_ = t_5__174_ | t_5__206_;
  assign t_6__173_ = t_5__173_ | t_5__205_;
  assign t_6__172_ = t_5__172_ | t_5__204_;
  assign t_6__171_ = t_5__171_ | t_5__203_;
  assign t_6__170_ = t_5__170_ | t_5__202_;
  assign t_6__169_ = t_5__169_ | t_5__201_;
  assign t_6__168_ = t_5__168_ | t_5__200_;
  assign t_6__167_ = t_5__167_ | t_5__199_;
  assign t_6__166_ = t_5__166_ | t_5__198_;
  assign t_6__165_ = t_5__165_ | t_5__197_;
  assign t_6__164_ = t_5__164_ | t_5__196_;
  assign t_6__163_ = t_5__163_ | t_5__195_;
  assign t_6__162_ = t_5__162_ | t_5__194_;
  assign t_6__161_ = t_5__161_ | t_5__193_;
  assign t_6__160_ = t_5__160_ | t_5__192_;
  assign t_6__159_ = t_5__159_ | t_5__191_;
  assign t_6__158_ = t_5__158_ | t_5__190_;
  assign t_6__157_ = t_5__157_ | t_5__189_;
  assign t_6__156_ = t_5__156_ | t_5__188_;
  assign t_6__155_ = t_5__155_ | t_5__187_;
  assign t_6__154_ = t_5__154_ | t_5__186_;
  assign t_6__153_ = t_5__153_ | t_5__185_;
  assign t_6__152_ = t_5__152_ | t_5__184_;
  assign t_6__151_ = t_5__151_ | t_5__183_;
  assign t_6__150_ = t_5__150_ | t_5__182_;
  assign t_6__149_ = t_5__149_ | t_5__181_;
  assign t_6__148_ = t_5__148_ | t_5__180_;
  assign t_6__147_ = t_5__147_ | t_5__179_;
  assign t_6__146_ = t_5__146_ | t_5__178_;
  assign t_6__145_ = t_5__145_ | t_5__177_;
  assign t_6__144_ = t_5__144_ | t_5__176_;
  assign t_6__143_ = t_5__143_ | t_5__175_;
  assign t_6__142_ = t_5__142_ | t_5__174_;
  assign t_6__141_ = t_5__141_ | t_5__173_;
  assign t_6__140_ = t_5__140_ | t_5__172_;
  assign t_6__139_ = t_5__139_ | t_5__171_;
  assign t_6__138_ = t_5__138_ | t_5__170_;
  assign t_6__137_ = t_5__137_ | t_5__169_;
  assign t_6__136_ = t_5__136_ | t_5__168_;
  assign t_6__135_ = t_5__135_ | t_5__167_;
  assign t_6__134_ = t_5__134_ | t_5__166_;
  assign t_6__133_ = t_5__133_ | t_5__165_;
  assign t_6__132_ = t_5__132_ | t_5__164_;
  assign t_6__131_ = t_5__131_ | t_5__163_;
  assign t_6__130_ = t_5__130_ | t_5__162_;
  assign t_6__129_ = t_5__129_ | t_5__161_;
  assign t_6__128_ = t_5__128_ | t_5__160_;
  assign t_6__127_ = t_5__127_ | t_5__159_;
  assign t_6__126_ = t_5__126_ | t_5__158_;
  assign t_6__125_ = t_5__125_ | t_5__157_;
  assign t_6__124_ = t_5__124_ | t_5__156_;
  assign t_6__123_ = t_5__123_ | t_5__155_;
  assign t_6__122_ = t_5__122_ | t_5__154_;
  assign t_6__121_ = t_5__121_ | t_5__153_;
  assign t_6__120_ = t_5__120_ | t_5__152_;
  assign t_6__119_ = t_5__119_ | t_5__151_;
  assign t_6__118_ = t_5__118_ | t_5__150_;
  assign t_6__117_ = t_5__117_ | t_5__149_;
  assign t_6__116_ = t_5__116_ | t_5__148_;
  assign t_6__115_ = t_5__115_ | t_5__147_;
  assign t_6__114_ = t_5__114_ | t_5__146_;
  assign t_6__113_ = t_5__113_ | t_5__145_;
  assign t_6__112_ = t_5__112_ | t_5__144_;
  assign t_6__111_ = t_5__111_ | t_5__143_;
  assign t_6__110_ = t_5__110_ | t_5__142_;
  assign t_6__109_ = t_5__109_ | t_5__141_;
  assign t_6__108_ = t_5__108_ | t_5__140_;
  assign t_6__107_ = t_5__107_ | t_5__139_;
  assign t_6__106_ = t_5__106_ | t_5__138_;
  assign t_6__105_ = t_5__105_ | t_5__137_;
  assign t_6__104_ = t_5__104_ | t_5__136_;
  assign t_6__103_ = t_5__103_ | t_5__135_;
  assign t_6__102_ = t_5__102_ | t_5__134_;
  assign t_6__101_ = t_5__101_ | t_5__133_;
  assign t_6__100_ = t_5__100_ | t_5__132_;
  assign t_6__99_ = t_5__99_ | t_5__131_;
  assign t_6__98_ = t_5__98_ | t_5__130_;
  assign t_6__97_ = t_5__97_ | t_5__129_;
  assign t_6__96_ = t_5__96_ | t_5__128_;
  assign t_6__95_ = t_5__95_ | t_5__127_;
  assign t_6__94_ = t_5__94_ | t_5__126_;
  assign t_6__93_ = t_5__93_ | t_5__125_;
  assign t_6__92_ = t_5__92_ | t_5__124_;
  assign t_6__91_ = t_5__91_ | t_5__123_;
  assign t_6__90_ = t_5__90_ | t_5__122_;
  assign t_6__89_ = t_5__89_ | t_5__121_;
  assign t_6__88_ = t_5__88_ | t_5__120_;
  assign t_6__87_ = t_5__87_ | t_5__119_;
  assign t_6__86_ = t_5__86_ | t_5__118_;
  assign t_6__85_ = t_5__85_ | t_5__117_;
  assign t_6__84_ = t_5__84_ | t_5__116_;
  assign t_6__83_ = t_5__83_ | t_5__115_;
  assign t_6__82_ = t_5__82_ | t_5__114_;
  assign t_6__81_ = t_5__81_ | t_5__113_;
  assign t_6__80_ = t_5__80_ | t_5__112_;
  assign t_6__79_ = t_5__79_ | t_5__111_;
  assign t_6__78_ = t_5__78_ | t_5__110_;
  assign t_6__77_ = t_5__77_ | t_5__109_;
  assign t_6__76_ = t_5__76_ | t_5__108_;
  assign t_6__75_ = t_5__75_ | t_5__107_;
  assign t_6__74_ = t_5__74_ | t_5__106_;
  assign t_6__73_ = t_5__73_ | t_5__105_;
  assign t_6__72_ = t_5__72_ | t_5__104_;
  assign t_6__71_ = t_5__71_ | t_5__103_;
  assign t_6__70_ = t_5__70_ | t_5__102_;
  assign t_6__69_ = t_5__69_ | t_5__101_;
  assign t_6__68_ = t_5__68_ | t_5__100_;
  assign t_6__67_ = t_5__67_ | t_5__99_;
  assign t_6__66_ = t_5__66_ | t_5__98_;
  assign t_6__65_ = t_5__65_ | t_5__97_;
  assign t_6__64_ = t_5__64_ | t_5__96_;
  assign t_6__63_ = t_5__63_ | t_5__95_;
  assign t_6__62_ = t_5__62_ | t_5__94_;
  assign t_6__61_ = t_5__61_ | t_5__93_;
  assign t_6__60_ = t_5__60_ | t_5__92_;
  assign t_6__59_ = t_5__59_ | t_5__91_;
  assign t_6__58_ = t_5__58_ | t_5__90_;
  assign t_6__57_ = t_5__57_ | t_5__89_;
  assign t_6__56_ = t_5__56_ | t_5__88_;
  assign t_6__55_ = t_5__55_ | t_5__87_;
  assign t_6__54_ = t_5__54_ | t_5__86_;
  assign t_6__53_ = t_5__53_ | t_5__85_;
  assign t_6__52_ = t_5__52_ | t_5__84_;
  assign t_6__51_ = t_5__51_ | t_5__83_;
  assign t_6__50_ = t_5__50_ | t_5__82_;
  assign t_6__49_ = t_5__49_ | t_5__81_;
  assign t_6__48_ = t_5__48_ | t_5__80_;
  assign t_6__47_ = t_5__47_ | t_5__79_;
  assign t_6__46_ = t_5__46_ | t_5__78_;
  assign t_6__45_ = t_5__45_ | t_5__77_;
  assign t_6__44_ = t_5__44_ | t_5__76_;
  assign t_6__43_ = t_5__43_ | t_5__75_;
  assign t_6__42_ = t_5__42_ | t_5__74_;
  assign t_6__41_ = t_5__41_ | t_5__73_;
  assign t_6__40_ = t_5__40_ | t_5__72_;
  assign t_6__39_ = t_5__39_ | t_5__71_;
  assign t_6__38_ = t_5__38_ | t_5__70_;
  assign t_6__37_ = t_5__37_ | t_5__69_;
  assign t_6__36_ = t_5__36_ | t_5__68_;
  assign t_6__35_ = t_5__35_ | t_5__67_;
  assign t_6__34_ = t_5__34_ | t_5__66_;
  assign t_6__33_ = t_5__33_ | t_5__65_;
  assign t_6__32_ = t_5__32_ | t_5__64_;
  assign t_6__31_ = t_5__31_ | t_5__63_;
  assign t_6__30_ = t_5__30_ | t_5__62_;
  assign t_6__29_ = t_5__29_ | t_5__61_;
  assign t_6__28_ = t_5__28_ | t_5__60_;
  assign t_6__27_ = t_5__27_ | t_5__59_;
  assign t_6__26_ = t_5__26_ | t_5__58_;
  assign t_6__25_ = t_5__25_ | t_5__57_;
  assign t_6__24_ = t_5__24_ | t_5__56_;
  assign t_6__23_ = t_5__23_ | t_5__55_;
  assign t_6__22_ = t_5__22_ | t_5__54_;
  assign t_6__21_ = t_5__21_ | t_5__53_;
  assign t_6__20_ = t_5__20_ | t_5__52_;
  assign t_6__19_ = t_5__19_ | t_5__51_;
  assign t_6__18_ = t_5__18_ | t_5__50_;
  assign t_6__17_ = t_5__17_ | t_5__49_;
  assign t_6__16_ = t_5__16_ | t_5__48_;
  assign t_6__15_ = t_5__15_ | t_5__47_;
  assign t_6__14_ = t_5__14_ | t_5__46_;
  assign t_6__13_ = t_5__13_ | t_5__45_;
  assign t_6__12_ = t_5__12_ | t_5__44_;
  assign t_6__11_ = t_5__11_ | t_5__43_;
  assign t_6__10_ = t_5__10_ | t_5__42_;
  assign t_6__9_ = t_5__9_ | t_5__41_;
  assign t_6__8_ = t_5__8_ | t_5__40_;
  assign t_6__7_ = t_5__7_ | t_5__39_;
  assign t_6__6_ = t_5__6_ | t_5__38_;
  assign t_6__5_ = t_5__5_ | t_5__37_;
  assign t_6__4_ = t_5__4_ | t_5__36_;
  assign t_6__3_ = t_5__3_ | t_5__35_;
  assign t_6__2_ = t_5__2_ | t_5__34_;
  assign t_6__1_ = t_5__1_ | t_5__33_;
  assign t_6__0_ = t_5__0_ | t_5__32_;
  assign t_7__511_ = t_6__511_ | 1'b0;
  assign t_7__510_ = t_6__510_ | 1'b0;
  assign t_7__509_ = t_6__509_ | 1'b0;
  assign t_7__508_ = t_6__508_ | 1'b0;
  assign t_7__507_ = t_6__507_ | 1'b0;
  assign t_7__506_ = t_6__506_ | 1'b0;
  assign t_7__505_ = t_6__505_ | 1'b0;
  assign t_7__504_ = t_6__504_ | 1'b0;
  assign t_7__503_ = t_6__503_ | 1'b0;
  assign t_7__502_ = t_6__502_ | 1'b0;
  assign t_7__501_ = t_6__501_ | 1'b0;
  assign t_7__500_ = t_6__500_ | 1'b0;
  assign t_7__499_ = t_6__499_ | 1'b0;
  assign t_7__498_ = t_6__498_ | 1'b0;
  assign t_7__497_ = t_6__497_ | 1'b0;
  assign t_7__496_ = t_6__496_ | 1'b0;
  assign t_7__495_ = t_6__495_ | 1'b0;
  assign t_7__494_ = t_6__494_ | 1'b0;
  assign t_7__493_ = t_6__493_ | 1'b0;
  assign t_7__492_ = t_6__492_ | 1'b0;
  assign t_7__491_ = t_6__491_ | 1'b0;
  assign t_7__490_ = t_6__490_ | 1'b0;
  assign t_7__489_ = t_6__489_ | 1'b0;
  assign t_7__488_ = t_6__488_ | 1'b0;
  assign t_7__487_ = t_6__487_ | 1'b0;
  assign t_7__486_ = t_6__486_ | 1'b0;
  assign t_7__485_ = t_6__485_ | 1'b0;
  assign t_7__484_ = t_6__484_ | 1'b0;
  assign t_7__483_ = t_6__483_ | 1'b0;
  assign t_7__482_ = t_6__482_ | 1'b0;
  assign t_7__481_ = t_6__481_ | 1'b0;
  assign t_7__480_ = t_6__480_ | 1'b0;
  assign t_7__479_ = t_6__479_ | 1'b0;
  assign t_7__478_ = t_6__478_ | 1'b0;
  assign t_7__477_ = t_6__477_ | 1'b0;
  assign t_7__476_ = t_6__476_ | 1'b0;
  assign t_7__475_ = t_6__475_ | 1'b0;
  assign t_7__474_ = t_6__474_ | 1'b0;
  assign t_7__473_ = t_6__473_ | 1'b0;
  assign t_7__472_ = t_6__472_ | 1'b0;
  assign t_7__471_ = t_6__471_ | 1'b0;
  assign t_7__470_ = t_6__470_ | 1'b0;
  assign t_7__469_ = t_6__469_ | 1'b0;
  assign t_7__468_ = t_6__468_ | 1'b0;
  assign t_7__467_ = t_6__467_ | 1'b0;
  assign t_7__466_ = t_6__466_ | 1'b0;
  assign t_7__465_ = t_6__465_ | 1'b0;
  assign t_7__464_ = t_6__464_ | 1'b0;
  assign t_7__463_ = t_6__463_ | 1'b0;
  assign t_7__462_ = t_6__462_ | 1'b0;
  assign t_7__461_ = t_6__461_ | 1'b0;
  assign t_7__460_ = t_6__460_ | 1'b0;
  assign t_7__459_ = t_6__459_ | 1'b0;
  assign t_7__458_ = t_6__458_ | 1'b0;
  assign t_7__457_ = t_6__457_ | 1'b0;
  assign t_7__456_ = t_6__456_ | 1'b0;
  assign t_7__455_ = t_6__455_ | 1'b0;
  assign t_7__454_ = t_6__454_ | 1'b0;
  assign t_7__453_ = t_6__453_ | 1'b0;
  assign t_7__452_ = t_6__452_ | 1'b0;
  assign t_7__451_ = t_6__451_ | 1'b0;
  assign t_7__450_ = t_6__450_ | 1'b0;
  assign t_7__449_ = t_6__449_ | 1'b0;
  assign t_7__448_ = t_6__448_ | 1'b0;
  assign t_7__447_ = t_6__447_ | t_6__511_;
  assign t_7__446_ = t_6__446_ | t_6__510_;
  assign t_7__445_ = t_6__445_ | t_6__509_;
  assign t_7__444_ = t_6__444_ | t_6__508_;
  assign t_7__443_ = t_6__443_ | t_6__507_;
  assign t_7__442_ = t_6__442_ | t_6__506_;
  assign t_7__441_ = t_6__441_ | t_6__505_;
  assign t_7__440_ = t_6__440_ | t_6__504_;
  assign t_7__439_ = t_6__439_ | t_6__503_;
  assign t_7__438_ = t_6__438_ | t_6__502_;
  assign t_7__437_ = t_6__437_ | t_6__501_;
  assign t_7__436_ = t_6__436_ | t_6__500_;
  assign t_7__435_ = t_6__435_ | t_6__499_;
  assign t_7__434_ = t_6__434_ | t_6__498_;
  assign t_7__433_ = t_6__433_ | t_6__497_;
  assign t_7__432_ = t_6__432_ | t_6__496_;
  assign t_7__431_ = t_6__431_ | t_6__495_;
  assign t_7__430_ = t_6__430_ | t_6__494_;
  assign t_7__429_ = t_6__429_ | t_6__493_;
  assign t_7__428_ = t_6__428_ | t_6__492_;
  assign t_7__427_ = t_6__427_ | t_6__491_;
  assign t_7__426_ = t_6__426_ | t_6__490_;
  assign t_7__425_ = t_6__425_ | t_6__489_;
  assign t_7__424_ = t_6__424_ | t_6__488_;
  assign t_7__423_ = t_6__423_ | t_6__487_;
  assign t_7__422_ = t_6__422_ | t_6__486_;
  assign t_7__421_ = t_6__421_ | t_6__485_;
  assign t_7__420_ = t_6__420_ | t_6__484_;
  assign t_7__419_ = t_6__419_ | t_6__483_;
  assign t_7__418_ = t_6__418_ | t_6__482_;
  assign t_7__417_ = t_6__417_ | t_6__481_;
  assign t_7__416_ = t_6__416_ | t_6__480_;
  assign t_7__415_ = t_6__415_ | t_6__479_;
  assign t_7__414_ = t_6__414_ | t_6__478_;
  assign t_7__413_ = t_6__413_ | t_6__477_;
  assign t_7__412_ = t_6__412_ | t_6__476_;
  assign t_7__411_ = t_6__411_ | t_6__475_;
  assign t_7__410_ = t_6__410_ | t_6__474_;
  assign t_7__409_ = t_6__409_ | t_6__473_;
  assign t_7__408_ = t_6__408_ | t_6__472_;
  assign t_7__407_ = t_6__407_ | t_6__471_;
  assign t_7__406_ = t_6__406_ | t_6__470_;
  assign t_7__405_ = t_6__405_ | t_6__469_;
  assign t_7__404_ = t_6__404_ | t_6__468_;
  assign t_7__403_ = t_6__403_ | t_6__467_;
  assign t_7__402_ = t_6__402_ | t_6__466_;
  assign t_7__401_ = t_6__401_ | t_6__465_;
  assign t_7__400_ = t_6__400_ | t_6__464_;
  assign t_7__399_ = t_6__399_ | t_6__463_;
  assign t_7__398_ = t_6__398_ | t_6__462_;
  assign t_7__397_ = t_6__397_ | t_6__461_;
  assign t_7__396_ = t_6__396_ | t_6__460_;
  assign t_7__395_ = t_6__395_ | t_6__459_;
  assign t_7__394_ = t_6__394_ | t_6__458_;
  assign t_7__393_ = t_6__393_ | t_6__457_;
  assign t_7__392_ = t_6__392_ | t_6__456_;
  assign t_7__391_ = t_6__391_ | t_6__455_;
  assign t_7__390_ = t_6__390_ | t_6__454_;
  assign t_7__389_ = t_6__389_ | t_6__453_;
  assign t_7__388_ = t_6__388_ | t_6__452_;
  assign t_7__387_ = t_6__387_ | t_6__451_;
  assign t_7__386_ = t_6__386_ | t_6__450_;
  assign t_7__385_ = t_6__385_ | t_6__449_;
  assign t_7__384_ = t_6__384_ | t_6__448_;
  assign t_7__383_ = t_6__383_ | t_6__447_;
  assign t_7__382_ = t_6__382_ | t_6__446_;
  assign t_7__381_ = t_6__381_ | t_6__445_;
  assign t_7__380_ = t_6__380_ | t_6__444_;
  assign t_7__379_ = t_6__379_ | t_6__443_;
  assign t_7__378_ = t_6__378_ | t_6__442_;
  assign t_7__377_ = t_6__377_ | t_6__441_;
  assign t_7__376_ = t_6__376_ | t_6__440_;
  assign t_7__375_ = t_6__375_ | t_6__439_;
  assign t_7__374_ = t_6__374_ | t_6__438_;
  assign t_7__373_ = t_6__373_ | t_6__437_;
  assign t_7__372_ = t_6__372_ | t_6__436_;
  assign t_7__371_ = t_6__371_ | t_6__435_;
  assign t_7__370_ = t_6__370_ | t_6__434_;
  assign t_7__369_ = t_6__369_ | t_6__433_;
  assign t_7__368_ = t_6__368_ | t_6__432_;
  assign t_7__367_ = t_6__367_ | t_6__431_;
  assign t_7__366_ = t_6__366_ | t_6__430_;
  assign t_7__365_ = t_6__365_ | t_6__429_;
  assign t_7__364_ = t_6__364_ | t_6__428_;
  assign t_7__363_ = t_6__363_ | t_6__427_;
  assign t_7__362_ = t_6__362_ | t_6__426_;
  assign t_7__361_ = t_6__361_ | t_6__425_;
  assign t_7__360_ = t_6__360_ | t_6__424_;
  assign t_7__359_ = t_6__359_ | t_6__423_;
  assign t_7__358_ = t_6__358_ | t_6__422_;
  assign t_7__357_ = t_6__357_ | t_6__421_;
  assign t_7__356_ = t_6__356_ | t_6__420_;
  assign t_7__355_ = t_6__355_ | t_6__419_;
  assign t_7__354_ = t_6__354_ | t_6__418_;
  assign t_7__353_ = t_6__353_ | t_6__417_;
  assign t_7__352_ = t_6__352_ | t_6__416_;
  assign t_7__351_ = t_6__351_ | t_6__415_;
  assign t_7__350_ = t_6__350_ | t_6__414_;
  assign t_7__349_ = t_6__349_ | t_6__413_;
  assign t_7__348_ = t_6__348_ | t_6__412_;
  assign t_7__347_ = t_6__347_ | t_6__411_;
  assign t_7__346_ = t_6__346_ | t_6__410_;
  assign t_7__345_ = t_6__345_ | t_6__409_;
  assign t_7__344_ = t_6__344_ | t_6__408_;
  assign t_7__343_ = t_6__343_ | t_6__407_;
  assign t_7__342_ = t_6__342_ | t_6__406_;
  assign t_7__341_ = t_6__341_ | t_6__405_;
  assign t_7__340_ = t_6__340_ | t_6__404_;
  assign t_7__339_ = t_6__339_ | t_6__403_;
  assign t_7__338_ = t_6__338_ | t_6__402_;
  assign t_7__337_ = t_6__337_ | t_6__401_;
  assign t_7__336_ = t_6__336_ | t_6__400_;
  assign t_7__335_ = t_6__335_ | t_6__399_;
  assign t_7__334_ = t_6__334_ | t_6__398_;
  assign t_7__333_ = t_6__333_ | t_6__397_;
  assign t_7__332_ = t_6__332_ | t_6__396_;
  assign t_7__331_ = t_6__331_ | t_6__395_;
  assign t_7__330_ = t_6__330_ | t_6__394_;
  assign t_7__329_ = t_6__329_ | t_6__393_;
  assign t_7__328_ = t_6__328_ | t_6__392_;
  assign t_7__327_ = t_6__327_ | t_6__391_;
  assign t_7__326_ = t_6__326_ | t_6__390_;
  assign t_7__325_ = t_6__325_ | t_6__389_;
  assign t_7__324_ = t_6__324_ | t_6__388_;
  assign t_7__323_ = t_6__323_ | t_6__387_;
  assign t_7__322_ = t_6__322_ | t_6__386_;
  assign t_7__321_ = t_6__321_ | t_6__385_;
  assign t_7__320_ = t_6__320_ | t_6__384_;
  assign t_7__319_ = t_6__319_ | t_6__383_;
  assign t_7__318_ = t_6__318_ | t_6__382_;
  assign t_7__317_ = t_6__317_ | t_6__381_;
  assign t_7__316_ = t_6__316_ | t_6__380_;
  assign t_7__315_ = t_6__315_ | t_6__379_;
  assign t_7__314_ = t_6__314_ | t_6__378_;
  assign t_7__313_ = t_6__313_ | t_6__377_;
  assign t_7__312_ = t_6__312_ | t_6__376_;
  assign t_7__311_ = t_6__311_ | t_6__375_;
  assign t_7__310_ = t_6__310_ | t_6__374_;
  assign t_7__309_ = t_6__309_ | t_6__373_;
  assign t_7__308_ = t_6__308_ | t_6__372_;
  assign t_7__307_ = t_6__307_ | t_6__371_;
  assign t_7__306_ = t_6__306_ | t_6__370_;
  assign t_7__305_ = t_6__305_ | t_6__369_;
  assign t_7__304_ = t_6__304_ | t_6__368_;
  assign t_7__303_ = t_6__303_ | t_6__367_;
  assign t_7__302_ = t_6__302_ | t_6__366_;
  assign t_7__301_ = t_6__301_ | t_6__365_;
  assign t_7__300_ = t_6__300_ | t_6__364_;
  assign t_7__299_ = t_6__299_ | t_6__363_;
  assign t_7__298_ = t_6__298_ | t_6__362_;
  assign t_7__297_ = t_6__297_ | t_6__361_;
  assign t_7__296_ = t_6__296_ | t_6__360_;
  assign t_7__295_ = t_6__295_ | t_6__359_;
  assign t_7__294_ = t_6__294_ | t_6__358_;
  assign t_7__293_ = t_6__293_ | t_6__357_;
  assign t_7__292_ = t_6__292_ | t_6__356_;
  assign t_7__291_ = t_6__291_ | t_6__355_;
  assign t_7__290_ = t_6__290_ | t_6__354_;
  assign t_7__289_ = t_6__289_ | t_6__353_;
  assign t_7__288_ = t_6__288_ | t_6__352_;
  assign t_7__287_ = t_6__287_ | t_6__351_;
  assign t_7__286_ = t_6__286_ | t_6__350_;
  assign t_7__285_ = t_6__285_ | t_6__349_;
  assign t_7__284_ = t_6__284_ | t_6__348_;
  assign t_7__283_ = t_6__283_ | t_6__347_;
  assign t_7__282_ = t_6__282_ | t_6__346_;
  assign t_7__281_ = t_6__281_ | t_6__345_;
  assign t_7__280_ = t_6__280_ | t_6__344_;
  assign t_7__279_ = t_6__279_ | t_6__343_;
  assign t_7__278_ = t_6__278_ | t_6__342_;
  assign t_7__277_ = t_6__277_ | t_6__341_;
  assign t_7__276_ = t_6__276_ | t_6__340_;
  assign t_7__275_ = t_6__275_ | t_6__339_;
  assign t_7__274_ = t_6__274_ | t_6__338_;
  assign t_7__273_ = t_6__273_ | t_6__337_;
  assign t_7__272_ = t_6__272_ | t_6__336_;
  assign t_7__271_ = t_6__271_ | t_6__335_;
  assign t_7__270_ = t_6__270_ | t_6__334_;
  assign t_7__269_ = t_6__269_ | t_6__333_;
  assign t_7__268_ = t_6__268_ | t_6__332_;
  assign t_7__267_ = t_6__267_ | t_6__331_;
  assign t_7__266_ = t_6__266_ | t_6__330_;
  assign t_7__265_ = t_6__265_ | t_6__329_;
  assign t_7__264_ = t_6__264_ | t_6__328_;
  assign t_7__263_ = t_6__263_ | t_6__327_;
  assign t_7__262_ = t_6__262_ | t_6__326_;
  assign t_7__261_ = t_6__261_ | t_6__325_;
  assign t_7__260_ = t_6__260_ | t_6__324_;
  assign t_7__259_ = t_6__259_ | t_6__323_;
  assign t_7__258_ = t_6__258_ | t_6__322_;
  assign t_7__257_ = t_6__257_ | t_6__321_;
  assign t_7__256_ = t_6__256_ | t_6__320_;
  assign t_7__255_ = t_6__255_ | t_6__319_;
  assign t_7__254_ = t_6__254_ | t_6__318_;
  assign t_7__253_ = t_6__253_ | t_6__317_;
  assign t_7__252_ = t_6__252_ | t_6__316_;
  assign t_7__251_ = t_6__251_ | t_6__315_;
  assign t_7__250_ = t_6__250_ | t_6__314_;
  assign t_7__249_ = t_6__249_ | t_6__313_;
  assign t_7__248_ = t_6__248_ | t_6__312_;
  assign t_7__247_ = t_6__247_ | t_6__311_;
  assign t_7__246_ = t_6__246_ | t_6__310_;
  assign t_7__245_ = t_6__245_ | t_6__309_;
  assign t_7__244_ = t_6__244_ | t_6__308_;
  assign t_7__243_ = t_6__243_ | t_6__307_;
  assign t_7__242_ = t_6__242_ | t_6__306_;
  assign t_7__241_ = t_6__241_ | t_6__305_;
  assign t_7__240_ = t_6__240_ | t_6__304_;
  assign t_7__239_ = t_6__239_ | t_6__303_;
  assign t_7__238_ = t_6__238_ | t_6__302_;
  assign t_7__237_ = t_6__237_ | t_6__301_;
  assign t_7__236_ = t_6__236_ | t_6__300_;
  assign t_7__235_ = t_6__235_ | t_6__299_;
  assign t_7__234_ = t_6__234_ | t_6__298_;
  assign t_7__233_ = t_6__233_ | t_6__297_;
  assign t_7__232_ = t_6__232_ | t_6__296_;
  assign t_7__231_ = t_6__231_ | t_6__295_;
  assign t_7__230_ = t_6__230_ | t_6__294_;
  assign t_7__229_ = t_6__229_ | t_6__293_;
  assign t_7__228_ = t_6__228_ | t_6__292_;
  assign t_7__227_ = t_6__227_ | t_6__291_;
  assign t_7__226_ = t_6__226_ | t_6__290_;
  assign t_7__225_ = t_6__225_ | t_6__289_;
  assign t_7__224_ = t_6__224_ | t_6__288_;
  assign t_7__223_ = t_6__223_ | t_6__287_;
  assign t_7__222_ = t_6__222_ | t_6__286_;
  assign t_7__221_ = t_6__221_ | t_6__285_;
  assign t_7__220_ = t_6__220_ | t_6__284_;
  assign t_7__219_ = t_6__219_ | t_6__283_;
  assign t_7__218_ = t_6__218_ | t_6__282_;
  assign t_7__217_ = t_6__217_ | t_6__281_;
  assign t_7__216_ = t_6__216_ | t_6__280_;
  assign t_7__215_ = t_6__215_ | t_6__279_;
  assign t_7__214_ = t_6__214_ | t_6__278_;
  assign t_7__213_ = t_6__213_ | t_6__277_;
  assign t_7__212_ = t_6__212_ | t_6__276_;
  assign t_7__211_ = t_6__211_ | t_6__275_;
  assign t_7__210_ = t_6__210_ | t_6__274_;
  assign t_7__209_ = t_6__209_ | t_6__273_;
  assign t_7__208_ = t_6__208_ | t_6__272_;
  assign t_7__207_ = t_6__207_ | t_6__271_;
  assign t_7__206_ = t_6__206_ | t_6__270_;
  assign t_7__205_ = t_6__205_ | t_6__269_;
  assign t_7__204_ = t_6__204_ | t_6__268_;
  assign t_7__203_ = t_6__203_ | t_6__267_;
  assign t_7__202_ = t_6__202_ | t_6__266_;
  assign t_7__201_ = t_6__201_ | t_6__265_;
  assign t_7__200_ = t_6__200_ | t_6__264_;
  assign t_7__199_ = t_6__199_ | t_6__263_;
  assign t_7__198_ = t_6__198_ | t_6__262_;
  assign t_7__197_ = t_6__197_ | t_6__261_;
  assign t_7__196_ = t_6__196_ | t_6__260_;
  assign t_7__195_ = t_6__195_ | t_6__259_;
  assign t_7__194_ = t_6__194_ | t_6__258_;
  assign t_7__193_ = t_6__193_ | t_6__257_;
  assign t_7__192_ = t_6__192_ | t_6__256_;
  assign t_7__191_ = t_6__191_ | t_6__255_;
  assign t_7__190_ = t_6__190_ | t_6__254_;
  assign t_7__189_ = t_6__189_ | t_6__253_;
  assign t_7__188_ = t_6__188_ | t_6__252_;
  assign t_7__187_ = t_6__187_ | t_6__251_;
  assign t_7__186_ = t_6__186_ | t_6__250_;
  assign t_7__185_ = t_6__185_ | t_6__249_;
  assign t_7__184_ = t_6__184_ | t_6__248_;
  assign t_7__183_ = t_6__183_ | t_6__247_;
  assign t_7__182_ = t_6__182_ | t_6__246_;
  assign t_7__181_ = t_6__181_ | t_6__245_;
  assign t_7__180_ = t_6__180_ | t_6__244_;
  assign t_7__179_ = t_6__179_ | t_6__243_;
  assign t_7__178_ = t_6__178_ | t_6__242_;
  assign t_7__177_ = t_6__177_ | t_6__241_;
  assign t_7__176_ = t_6__176_ | t_6__240_;
  assign t_7__175_ = t_6__175_ | t_6__239_;
  assign t_7__174_ = t_6__174_ | t_6__238_;
  assign t_7__173_ = t_6__173_ | t_6__237_;
  assign t_7__172_ = t_6__172_ | t_6__236_;
  assign t_7__171_ = t_6__171_ | t_6__235_;
  assign t_7__170_ = t_6__170_ | t_6__234_;
  assign t_7__169_ = t_6__169_ | t_6__233_;
  assign t_7__168_ = t_6__168_ | t_6__232_;
  assign t_7__167_ = t_6__167_ | t_6__231_;
  assign t_7__166_ = t_6__166_ | t_6__230_;
  assign t_7__165_ = t_6__165_ | t_6__229_;
  assign t_7__164_ = t_6__164_ | t_6__228_;
  assign t_7__163_ = t_6__163_ | t_6__227_;
  assign t_7__162_ = t_6__162_ | t_6__226_;
  assign t_7__161_ = t_6__161_ | t_6__225_;
  assign t_7__160_ = t_6__160_ | t_6__224_;
  assign t_7__159_ = t_6__159_ | t_6__223_;
  assign t_7__158_ = t_6__158_ | t_6__222_;
  assign t_7__157_ = t_6__157_ | t_6__221_;
  assign t_7__156_ = t_6__156_ | t_6__220_;
  assign t_7__155_ = t_6__155_ | t_6__219_;
  assign t_7__154_ = t_6__154_ | t_6__218_;
  assign t_7__153_ = t_6__153_ | t_6__217_;
  assign t_7__152_ = t_6__152_ | t_6__216_;
  assign t_7__151_ = t_6__151_ | t_6__215_;
  assign t_7__150_ = t_6__150_ | t_6__214_;
  assign t_7__149_ = t_6__149_ | t_6__213_;
  assign t_7__148_ = t_6__148_ | t_6__212_;
  assign t_7__147_ = t_6__147_ | t_6__211_;
  assign t_7__146_ = t_6__146_ | t_6__210_;
  assign t_7__145_ = t_6__145_ | t_6__209_;
  assign t_7__144_ = t_6__144_ | t_6__208_;
  assign t_7__143_ = t_6__143_ | t_6__207_;
  assign t_7__142_ = t_6__142_ | t_6__206_;
  assign t_7__141_ = t_6__141_ | t_6__205_;
  assign t_7__140_ = t_6__140_ | t_6__204_;
  assign t_7__139_ = t_6__139_ | t_6__203_;
  assign t_7__138_ = t_6__138_ | t_6__202_;
  assign t_7__137_ = t_6__137_ | t_6__201_;
  assign t_7__136_ = t_6__136_ | t_6__200_;
  assign t_7__135_ = t_6__135_ | t_6__199_;
  assign t_7__134_ = t_6__134_ | t_6__198_;
  assign t_7__133_ = t_6__133_ | t_6__197_;
  assign t_7__132_ = t_6__132_ | t_6__196_;
  assign t_7__131_ = t_6__131_ | t_6__195_;
  assign t_7__130_ = t_6__130_ | t_6__194_;
  assign t_7__129_ = t_6__129_ | t_6__193_;
  assign t_7__128_ = t_6__128_ | t_6__192_;
  assign t_7__127_ = t_6__127_ | t_6__191_;
  assign t_7__126_ = t_6__126_ | t_6__190_;
  assign t_7__125_ = t_6__125_ | t_6__189_;
  assign t_7__124_ = t_6__124_ | t_6__188_;
  assign t_7__123_ = t_6__123_ | t_6__187_;
  assign t_7__122_ = t_6__122_ | t_6__186_;
  assign t_7__121_ = t_6__121_ | t_6__185_;
  assign t_7__120_ = t_6__120_ | t_6__184_;
  assign t_7__119_ = t_6__119_ | t_6__183_;
  assign t_7__118_ = t_6__118_ | t_6__182_;
  assign t_7__117_ = t_6__117_ | t_6__181_;
  assign t_7__116_ = t_6__116_ | t_6__180_;
  assign t_7__115_ = t_6__115_ | t_6__179_;
  assign t_7__114_ = t_6__114_ | t_6__178_;
  assign t_7__113_ = t_6__113_ | t_6__177_;
  assign t_7__112_ = t_6__112_ | t_6__176_;
  assign t_7__111_ = t_6__111_ | t_6__175_;
  assign t_7__110_ = t_6__110_ | t_6__174_;
  assign t_7__109_ = t_6__109_ | t_6__173_;
  assign t_7__108_ = t_6__108_ | t_6__172_;
  assign t_7__107_ = t_6__107_ | t_6__171_;
  assign t_7__106_ = t_6__106_ | t_6__170_;
  assign t_7__105_ = t_6__105_ | t_6__169_;
  assign t_7__104_ = t_6__104_ | t_6__168_;
  assign t_7__103_ = t_6__103_ | t_6__167_;
  assign t_7__102_ = t_6__102_ | t_6__166_;
  assign t_7__101_ = t_6__101_ | t_6__165_;
  assign t_7__100_ = t_6__100_ | t_6__164_;
  assign t_7__99_ = t_6__99_ | t_6__163_;
  assign t_7__98_ = t_6__98_ | t_6__162_;
  assign t_7__97_ = t_6__97_ | t_6__161_;
  assign t_7__96_ = t_6__96_ | t_6__160_;
  assign t_7__95_ = t_6__95_ | t_6__159_;
  assign t_7__94_ = t_6__94_ | t_6__158_;
  assign t_7__93_ = t_6__93_ | t_6__157_;
  assign t_7__92_ = t_6__92_ | t_6__156_;
  assign t_7__91_ = t_6__91_ | t_6__155_;
  assign t_7__90_ = t_6__90_ | t_6__154_;
  assign t_7__89_ = t_6__89_ | t_6__153_;
  assign t_7__88_ = t_6__88_ | t_6__152_;
  assign t_7__87_ = t_6__87_ | t_6__151_;
  assign t_7__86_ = t_6__86_ | t_6__150_;
  assign t_7__85_ = t_6__85_ | t_6__149_;
  assign t_7__84_ = t_6__84_ | t_6__148_;
  assign t_7__83_ = t_6__83_ | t_6__147_;
  assign t_7__82_ = t_6__82_ | t_6__146_;
  assign t_7__81_ = t_6__81_ | t_6__145_;
  assign t_7__80_ = t_6__80_ | t_6__144_;
  assign t_7__79_ = t_6__79_ | t_6__143_;
  assign t_7__78_ = t_6__78_ | t_6__142_;
  assign t_7__77_ = t_6__77_ | t_6__141_;
  assign t_7__76_ = t_6__76_ | t_6__140_;
  assign t_7__75_ = t_6__75_ | t_6__139_;
  assign t_7__74_ = t_6__74_ | t_6__138_;
  assign t_7__73_ = t_6__73_ | t_6__137_;
  assign t_7__72_ = t_6__72_ | t_6__136_;
  assign t_7__71_ = t_6__71_ | t_6__135_;
  assign t_7__70_ = t_6__70_ | t_6__134_;
  assign t_7__69_ = t_6__69_ | t_6__133_;
  assign t_7__68_ = t_6__68_ | t_6__132_;
  assign t_7__67_ = t_6__67_ | t_6__131_;
  assign t_7__66_ = t_6__66_ | t_6__130_;
  assign t_7__65_ = t_6__65_ | t_6__129_;
  assign t_7__64_ = t_6__64_ | t_6__128_;
  assign t_7__63_ = t_6__63_ | t_6__127_;
  assign t_7__62_ = t_6__62_ | t_6__126_;
  assign t_7__61_ = t_6__61_ | t_6__125_;
  assign t_7__60_ = t_6__60_ | t_6__124_;
  assign t_7__59_ = t_6__59_ | t_6__123_;
  assign t_7__58_ = t_6__58_ | t_6__122_;
  assign t_7__57_ = t_6__57_ | t_6__121_;
  assign t_7__56_ = t_6__56_ | t_6__120_;
  assign t_7__55_ = t_6__55_ | t_6__119_;
  assign t_7__54_ = t_6__54_ | t_6__118_;
  assign t_7__53_ = t_6__53_ | t_6__117_;
  assign t_7__52_ = t_6__52_ | t_6__116_;
  assign t_7__51_ = t_6__51_ | t_6__115_;
  assign t_7__50_ = t_6__50_ | t_6__114_;
  assign t_7__49_ = t_6__49_ | t_6__113_;
  assign t_7__48_ = t_6__48_ | t_6__112_;
  assign t_7__47_ = t_6__47_ | t_6__111_;
  assign t_7__46_ = t_6__46_ | t_6__110_;
  assign t_7__45_ = t_6__45_ | t_6__109_;
  assign t_7__44_ = t_6__44_ | t_6__108_;
  assign t_7__43_ = t_6__43_ | t_6__107_;
  assign t_7__42_ = t_6__42_ | t_6__106_;
  assign t_7__41_ = t_6__41_ | t_6__105_;
  assign t_7__40_ = t_6__40_ | t_6__104_;
  assign t_7__39_ = t_6__39_ | t_6__103_;
  assign t_7__38_ = t_6__38_ | t_6__102_;
  assign t_7__37_ = t_6__37_ | t_6__101_;
  assign t_7__36_ = t_6__36_ | t_6__100_;
  assign t_7__35_ = t_6__35_ | t_6__99_;
  assign t_7__34_ = t_6__34_ | t_6__98_;
  assign t_7__33_ = t_6__33_ | t_6__97_;
  assign t_7__32_ = t_6__32_ | t_6__96_;
  assign t_7__31_ = t_6__31_ | t_6__95_;
  assign t_7__30_ = t_6__30_ | t_6__94_;
  assign t_7__29_ = t_6__29_ | t_6__93_;
  assign t_7__28_ = t_6__28_ | t_6__92_;
  assign t_7__27_ = t_6__27_ | t_6__91_;
  assign t_7__26_ = t_6__26_ | t_6__90_;
  assign t_7__25_ = t_6__25_ | t_6__89_;
  assign t_7__24_ = t_6__24_ | t_6__88_;
  assign t_7__23_ = t_6__23_ | t_6__87_;
  assign t_7__22_ = t_6__22_ | t_6__86_;
  assign t_7__21_ = t_6__21_ | t_6__85_;
  assign t_7__20_ = t_6__20_ | t_6__84_;
  assign t_7__19_ = t_6__19_ | t_6__83_;
  assign t_7__18_ = t_6__18_ | t_6__82_;
  assign t_7__17_ = t_6__17_ | t_6__81_;
  assign t_7__16_ = t_6__16_ | t_6__80_;
  assign t_7__15_ = t_6__15_ | t_6__79_;
  assign t_7__14_ = t_6__14_ | t_6__78_;
  assign t_7__13_ = t_6__13_ | t_6__77_;
  assign t_7__12_ = t_6__12_ | t_6__76_;
  assign t_7__11_ = t_6__11_ | t_6__75_;
  assign t_7__10_ = t_6__10_ | t_6__74_;
  assign t_7__9_ = t_6__9_ | t_6__73_;
  assign t_7__8_ = t_6__8_ | t_6__72_;
  assign t_7__7_ = t_6__7_ | t_6__71_;
  assign t_7__6_ = t_6__6_ | t_6__70_;
  assign t_7__5_ = t_6__5_ | t_6__69_;
  assign t_7__4_ = t_6__4_ | t_6__68_;
  assign t_7__3_ = t_6__3_ | t_6__67_;
  assign t_7__2_ = t_6__2_ | t_6__66_;
  assign t_7__1_ = t_6__1_ | t_6__65_;
  assign t_7__0_ = t_6__0_ | t_6__64_;
  assign t_8__511_ = t_7__511_ | 1'b0;
  assign t_8__510_ = t_7__510_ | 1'b0;
  assign t_8__509_ = t_7__509_ | 1'b0;
  assign t_8__508_ = t_7__508_ | 1'b0;
  assign t_8__507_ = t_7__507_ | 1'b0;
  assign t_8__506_ = t_7__506_ | 1'b0;
  assign t_8__505_ = t_7__505_ | 1'b0;
  assign t_8__504_ = t_7__504_ | 1'b0;
  assign t_8__503_ = t_7__503_ | 1'b0;
  assign t_8__502_ = t_7__502_ | 1'b0;
  assign t_8__501_ = t_7__501_ | 1'b0;
  assign t_8__500_ = t_7__500_ | 1'b0;
  assign t_8__499_ = t_7__499_ | 1'b0;
  assign t_8__498_ = t_7__498_ | 1'b0;
  assign t_8__497_ = t_7__497_ | 1'b0;
  assign t_8__496_ = t_7__496_ | 1'b0;
  assign t_8__495_ = t_7__495_ | 1'b0;
  assign t_8__494_ = t_7__494_ | 1'b0;
  assign t_8__493_ = t_7__493_ | 1'b0;
  assign t_8__492_ = t_7__492_ | 1'b0;
  assign t_8__491_ = t_7__491_ | 1'b0;
  assign t_8__490_ = t_7__490_ | 1'b0;
  assign t_8__489_ = t_7__489_ | 1'b0;
  assign t_8__488_ = t_7__488_ | 1'b0;
  assign t_8__487_ = t_7__487_ | 1'b0;
  assign t_8__486_ = t_7__486_ | 1'b0;
  assign t_8__485_ = t_7__485_ | 1'b0;
  assign t_8__484_ = t_7__484_ | 1'b0;
  assign t_8__483_ = t_7__483_ | 1'b0;
  assign t_8__482_ = t_7__482_ | 1'b0;
  assign t_8__481_ = t_7__481_ | 1'b0;
  assign t_8__480_ = t_7__480_ | 1'b0;
  assign t_8__479_ = t_7__479_ | 1'b0;
  assign t_8__478_ = t_7__478_ | 1'b0;
  assign t_8__477_ = t_7__477_ | 1'b0;
  assign t_8__476_ = t_7__476_ | 1'b0;
  assign t_8__475_ = t_7__475_ | 1'b0;
  assign t_8__474_ = t_7__474_ | 1'b0;
  assign t_8__473_ = t_7__473_ | 1'b0;
  assign t_8__472_ = t_7__472_ | 1'b0;
  assign t_8__471_ = t_7__471_ | 1'b0;
  assign t_8__470_ = t_7__470_ | 1'b0;
  assign t_8__469_ = t_7__469_ | 1'b0;
  assign t_8__468_ = t_7__468_ | 1'b0;
  assign t_8__467_ = t_7__467_ | 1'b0;
  assign t_8__466_ = t_7__466_ | 1'b0;
  assign t_8__465_ = t_7__465_ | 1'b0;
  assign t_8__464_ = t_7__464_ | 1'b0;
  assign t_8__463_ = t_7__463_ | 1'b0;
  assign t_8__462_ = t_7__462_ | 1'b0;
  assign t_8__461_ = t_7__461_ | 1'b0;
  assign t_8__460_ = t_7__460_ | 1'b0;
  assign t_8__459_ = t_7__459_ | 1'b0;
  assign t_8__458_ = t_7__458_ | 1'b0;
  assign t_8__457_ = t_7__457_ | 1'b0;
  assign t_8__456_ = t_7__456_ | 1'b0;
  assign t_8__455_ = t_7__455_ | 1'b0;
  assign t_8__454_ = t_7__454_ | 1'b0;
  assign t_8__453_ = t_7__453_ | 1'b0;
  assign t_8__452_ = t_7__452_ | 1'b0;
  assign t_8__451_ = t_7__451_ | 1'b0;
  assign t_8__450_ = t_7__450_ | 1'b0;
  assign t_8__449_ = t_7__449_ | 1'b0;
  assign t_8__448_ = t_7__448_ | 1'b0;
  assign t_8__447_ = t_7__447_ | 1'b0;
  assign t_8__446_ = t_7__446_ | 1'b0;
  assign t_8__445_ = t_7__445_ | 1'b0;
  assign t_8__444_ = t_7__444_ | 1'b0;
  assign t_8__443_ = t_7__443_ | 1'b0;
  assign t_8__442_ = t_7__442_ | 1'b0;
  assign t_8__441_ = t_7__441_ | 1'b0;
  assign t_8__440_ = t_7__440_ | 1'b0;
  assign t_8__439_ = t_7__439_ | 1'b0;
  assign t_8__438_ = t_7__438_ | 1'b0;
  assign t_8__437_ = t_7__437_ | 1'b0;
  assign t_8__436_ = t_7__436_ | 1'b0;
  assign t_8__435_ = t_7__435_ | 1'b0;
  assign t_8__434_ = t_7__434_ | 1'b0;
  assign t_8__433_ = t_7__433_ | 1'b0;
  assign t_8__432_ = t_7__432_ | 1'b0;
  assign t_8__431_ = t_7__431_ | 1'b0;
  assign t_8__430_ = t_7__430_ | 1'b0;
  assign t_8__429_ = t_7__429_ | 1'b0;
  assign t_8__428_ = t_7__428_ | 1'b0;
  assign t_8__427_ = t_7__427_ | 1'b0;
  assign t_8__426_ = t_7__426_ | 1'b0;
  assign t_8__425_ = t_7__425_ | 1'b0;
  assign t_8__424_ = t_7__424_ | 1'b0;
  assign t_8__423_ = t_7__423_ | 1'b0;
  assign t_8__422_ = t_7__422_ | 1'b0;
  assign t_8__421_ = t_7__421_ | 1'b0;
  assign t_8__420_ = t_7__420_ | 1'b0;
  assign t_8__419_ = t_7__419_ | 1'b0;
  assign t_8__418_ = t_7__418_ | 1'b0;
  assign t_8__417_ = t_7__417_ | 1'b0;
  assign t_8__416_ = t_7__416_ | 1'b0;
  assign t_8__415_ = t_7__415_ | 1'b0;
  assign t_8__414_ = t_7__414_ | 1'b0;
  assign t_8__413_ = t_7__413_ | 1'b0;
  assign t_8__412_ = t_7__412_ | 1'b0;
  assign t_8__411_ = t_7__411_ | 1'b0;
  assign t_8__410_ = t_7__410_ | 1'b0;
  assign t_8__409_ = t_7__409_ | 1'b0;
  assign t_8__408_ = t_7__408_ | 1'b0;
  assign t_8__407_ = t_7__407_ | 1'b0;
  assign t_8__406_ = t_7__406_ | 1'b0;
  assign t_8__405_ = t_7__405_ | 1'b0;
  assign t_8__404_ = t_7__404_ | 1'b0;
  assign t_8__403_ = t_7__403_ | 1'b0;
  assign t_8__402_ = t_7__402_ | 1'b0;
  assign t_8__401_ = t_7__401_ | 1'b0;
  assign t_8__400_ = t_7__400_ | 1'b0;
  assign t_8__399_ = t_7__399_ | 1'b0;
  assign t_8__398_ = t_7__398_ | 1'b0;
  assign t_8__397_ = t_7__397_ | 1'b0;
  assign t_8__396_ = t_7__396_ | 1'b0;
  assign t_8__395_ = t_7__395_ | 1'b0;
  assign t_8__394_ = t_7__394_ | 1'b0;
  assign t_8__393_ = t_7__393_ | 1'b0;
  assign t_8__392_ = t_7__392_ | 1'b0;
  assign t_8__391_ = t_7__391_ | 1'b0;
  assign t_8__390_ = t_7__390_ | 1'b0;
  assign t_8__389_ = t_7__389_ | 1'b0;
  assign t_8__388_ = t_7__388_ | 1'b0;
  assign t_8__387_ = t_7__387_ | 1'b0;
  assign t_8__386_ = t_7__386_ | 1'b0;
  assign t_8__385_ = t_7__385_ | 1'b0;
  assign t_8__384_ = t_7__384_ | 1'b0;
  assign t_8__383_ = t_7__383_ | t_7__511_;
  assign t_8__382_ = t_7__382_ | t_7__510_;
  assign t_8__381_ = t_7__381_ | t_7__509_;
  assign t_8__380_ = t_7__380_ | t_7__508_;
  assign t_8__379_ = t_7__379_ | t_7__507_;
  assign t_8__378_ = t_7__378_ | t_7__506_;
  assign t_8__377_ = t_7__377_ | t_7__505_;
  assign t_8__376_ = t_7__376_ | t_7__504_;
  assign t_8__375_ = t_7__375_ | t_7__503_;
  assign t_8__374_ = t_7__374_ | t_7__502_;
  assign t_8__373_ = t_7__373_ | t_7__501_;
  assign t_8__372_ = t_7__372_ | t_7__500_;
  assign t_8__371_ = t_7__371_ | t_7__499_;
  assign t_8__370_ = t_7__370_ | t_7__498_;
  assign t_8__369_ = t_7__369_ | t_7__497_;
  assign t_8__368_ = t_7__368_ | t_7__496_;
  assign t_8__367_ = t_7__367_ | t_7__495_;
  assign t_8__366_ = t_7__366_ | t_7__494_;
  assign t_8__365_ = t_7__365_ | t_7__493_;
  assign t_8__364_ = t_7__364_ | t_7__492_;
  assign t_8__363_ = t_7__363_ | t_7__491_;
  assign t_8__362_ = t_7__362_ | t_7__490_;
  assign t_8__361_ = t_7__361_ | t_7__489_;
  assign t_8__360_ = t_7__360_ | t_7__488_;
  assign t_8__359_ = t_7__359_ | t_7__487_;
  assign t_8__358_ = t_7__358_ | t_7__486_;
  assign t_8__357_ = t_7__357_ | t_7__485_;
  assign t_8__356_ = t_7__356_ | t_7__484_;
  assign t_8__355_ = t_7__355_ | t_7__483_;
  assign t_8__354_ = t_7__354_ | t_7__482_;
  assign t_8__353_ = t_7__353_ | t_7__481_;
  assign t_8__352_ = t_7__352_ | t_7__480_;
  assign t_8__351_ = t_7__351_ | t_7__479_;
  assign t_8__350_ = t_7__350_ | t_7__478_;
  assign t_8__349_ = t_7__349_ | t_7__477_;
  assign t_8__348_ = t_7__348_ | t_7__476_;
  assign t_8__347_ = t_7__347_ | t_7__475_;
  assign t_8__346_ = t_7__346_ | t_7__474_;
  assign t_8__345_ = t_7__345_ | t_7__473_;
  assign t_8__344_ = t_7__344_ | t_7__472_;
  assign t_8__343_ = t_7__343_ | t_7__471_;
  assign t_8__342_ = t_7__342_ | t_7__470_;
  assign t_8__341_ = t_7__341_ | t_7__469_;
  assign t_8__340_ = t_7__340_ | t_7__468_;
  assign t_8__339_ = t_7__339_ | t_7__467_;
  assign t_8__338_ = t_7__338_ | t_7__466_;
  assign t_8__337_ = t_7__337_ | t_7__465_;
  assign t_8__336_ = t_7__336_ | t_7__464_;
  assign t_8__335_ = t_7__335_ | t_7__463_;
  assign t_8__334_ = t_7__334_ | t_7__462_;
  assign t_8__333_ = t_7__333_ | t_7__461_;
  assign t_8__332_ = t_7__332_ | t_7__460_;
  assign t_8__331_ = t_7__331_ | t_7__459_;
  assign t_8__330_ = t_7__330_ | t_7__458_;
  assign t_8__329_ = t_7__329_ | t_7__457_;
  assign t_8__328_ = t_7__328_ | t_7__456_;
  assign t_8__327_ = t_7__327_ | t_7__455_;
  assign t_8__326_ = t_7__326_ | t_7__454_;
  assign t_8__325_ = t_7__325_ | t_7__453_;
  assign t_8__324_ = t_7__324_ | t_7__452_;
  assign t_8__323_ = t_7__323_ | t_7__451_;
  assign t_8__322_ = t_7__322_ | t_7__450_;
  assign t_8__321_ = t_7__321_ | t_7__449_;
  assign t_8__320_ = t_7__320_ | t_7__448_;
  assign t_8__319_ = t_7__319_ | t_7__447_;
  assign t_8__318_ = t_7__318_ | t_7__446_;
  assign t_8__317_ = t_7__317_ | t_7__445_;
  assign t_8__316_ = t_7__316_ | t_7__444_;
  assign t_8__315_ = t_7__315_ | t_7__443_;
  assign t_8__314_ = t_7__314_ | t_7__442_;
  assign t_8__313_ = t_7__313_ | t_7__441_;
  assign t_8__312_ = t_7__312_ | t_7__440_;
  assign t_8__311_ = t_7__311_ | t_7__439_;
  assign t_8__310_ = t_7__310_ | t_7__438_;
  assign t_8__309_ = t_7__309_ | t_7__437_;
  assign t_8__308_ = t_7__308_ | t_7__436_;
  assign t_8__307_ = t_7__307_ | t_7__435_;
  assign t_8__306_ = t_7__306_ | t_7__434_;
  assign t_8__305_ = t_7__305_ | t_7__433_;
  assign t_8__304_ = t_7__304_ | t_7__432_;
  assign t_8__303_ = t_7__303_ | t_7__431_;
  assign t_8__302_ = t_7__302_ | t_7__430_;
  assign t_8__301_ = t_7__301_ | t_7__429_;
  assign t_8__300_ = t_7__300_ | t_7__428_;
  assign t_8__299_ = t_7__299_ | t_7__427_;
  assign t_8__298_ = t_7__298_ | t_7__426_;
  assign t_8__297_ = t_7__297_ | t_7__425_;
  assign t_8__296_ = t_7__296_ | t_7__424_;
  assign t_8__295_ = t_7__295_ | t_7__423_;
  assign t_8__294_ = t_7__294_ | t_7__422_;
  assign t_8__293_ = t_7__293_ | t_7__421_;
  assign t_8__292_ = t_7__292_ | t_7__420_;
  assign t_8__291_ = t_7__291_ | t_7__419_;
  assign t_8__290_ = t_7__290_ | t_7__418_;
  assign t_8__289_ = t_7__289_ | t_7__417_;
  assign t_8__288_ = t_7__288_ | t_7__416_;
  assign t_8__287_ = t_7__287_ | t_7__415_;
  assign t_8__286_ = t_7__286_ | t_7__414_;
  assign t_8__285_ = t_7__285_ | t_7__413_;
  assign t_8__284_ = t_7__284_ | t_7__412_;
  assign t_8__283_ = t_7__283_ | t_7__411_;
  assign t_8__282_ = t_7__282_ | t_7__410_;
  assign t_8__281_ = t_7__281_ | t_7__409_;
  assign t_8__280_ = t_7__280_ | t_7__408_;
  assign t_8__279_ = t_7__279_ | t_7__407_;
  assign t_8__278_ = t_7__278_ | t_7__406_;
  assign t_8__277_ = t_7__277_ | t_7__405_;
  assign t_8__276_ = t_7__276_ | t_7__404_;
  assign t_8__275_ = t_7__275_ | t_7__403_;
  assign t_8__274_ = t_7__274_ | t_7__402_;
  assign t_8__273_ = t_7__273_ | t_7__401_;
  assign t_8__272_ = t_7__272_ | t_7__400_;
  assign t_8__271_ = t_7__271_ | t_7__399_;
  assign t_8__270_ = t_7__270_ | t_7__398_;
  assign t_8__269_ = t_7__269_ | t_7__397_;
  assign t_8__268_ = t_7__268_ | t_7__396_;
  assign t_8__267_ = t_7__267_ | t_7__395_;
  assign t_8__266_ = t_7__266_ | t_7__394_;
  assign t_8__265_ = t_7__265_ | t_7__393_;
  assign t_8__264_ = t_7__264_ | t_7__392_;
  assign t_8__263_ = t_7__263_ | t_7__391_;
  assign t_8__262_ = t_7__262_ | t_7__390_;
  assign t_8__261_ = t_7__261_ | t_7__389_;
  assign t_8__260_ = t_7__260_ | t_7__388_;
  assign t_8__259_ = t_7__259_ | t_7__387_;
  assign t_8__258_ = t_7__258_ | t_7__386_;
  assign t_8__257_ = t_7__257_ | t_7__385_;
  assign t_8__256_ = t_7__256_ | t_7__384_;
  assign t_8__255_ = t_7__255_ | t_7__383_;
  assign t_8__254_ = t_7__254_ | t_7__382_;
  assign t_8__253_ = t_7__253_ | t_7__381_;
  assign t_8__252_ = t_7__252_ | t_7__380_;
  assign t_8__251_ = t_7__251_ | t_7__379_;
  assign t_8__250_ = t_7__250_ | t_7__378_;
  assign t_8__249_ = t_7__249_ | t_7__377_;
  assign t_8__248_ = t_7__248_ | t_7__376_;
  assign t_8__247_ = t_7__247_ | t_7__375_;
  assign t_8__246_ = t_7__246_ | t_7__374_;
  assign t_8__245_ = t_7__245_ | t_7__373_;
  assign t_8__244_ = t_7__244_ | t_7__372_;
  assign t_8__243_ = t_7__243_ | t_7__371_;
  assign t_8__242_ = t_7__242_ | t_7__370_;
  assign t_8__241_ = t_7__241_ | t_7__369_;
  assign t_8__240_ = t_7__240_ | t_7__368_;
  assign t_8__239_ = t_7__239_ | t_7__367_;
  assign t_8__238_ = t_7__238_ | t_7__366_;
  assign t_8__237_ = t_7__237_ | t_7__365_;
  assign t_8__236_ = t_7__236_ | t_7__364_;
  assign t_8__235_ = t_7__235_ | t_7__363_;
  assign t_8__234_ = t_7__234_ | t_7__362_;
  assign t_8__233_ = t_7__233_ | t_7__361_;
  assign t_8__232_ = t_7__232_ | t_7__360_;
  assign t_8__231_ = t_7__231_ | t_7__359_;
  assign t_8__230_ = t_7__230_ | t_7__358_;
  assign t_8__229_ = t_7__229_ | t_7__357_;
  assign t_8__228_ = t_7__228_ | t_7__356_;
  assign t_8__227_ = t_7__227_ | t_7__355_;
  assign t_8__226_ = t_7__226_ | t_7__354_;
  assign t_8__225_ = t_7__225_ | t_7__353_;
  assign t_8__224_ = t_7__224_ | t_7__352_;
  assign t_8__223_ = t_7__223_ | t_7__351_;
  assign t_8__222_ = t_7__222_ | t_7__350_;
  assign t_8__221_ = t_7__221_ | t_7__349_;
  assign t_8__220_ = t_7__220_ | t_7__348_;
  assign t_8__219_ = t_7__219_ | t_7__347_;
  assign t_8__218_ = t_7__218_ | t_7__346_;
  assign t_8__217_ = t_7__217_ | t_7__345_;
  assign t_8__216_ = t_7__216_ | t_7__344_;
  assign t_8__215_ = t_7__215_ | t_7__343_;
  assign t_8__214_ = t_7__214_ | t_7__342_;
  assign t_8__213_ = t_7__213_ | t_7__341_;
  assign t_8__212_ = t_7__212_ | t_7__340_;
  assign t_8__211_ = t_7__211_ | t_7__339_;
  assign t_8__210_ = t_7__210_ | t_7__338_;
  assign t_8__209_ = t_7__209_ | t_7__337_;
  assign t_8__208_ = t_7__208_ | t_7__336_;
  assign t_8__207_ = t_7__207_ | t_7__335_;
  assign t_8__206_ = t_7__206_ | t_7__334_;
  assign t_8__205_ = t_7__205_ | t_7__333_;
  assign t_8__204_ = t_7__204_ | t_7__332_;
  assign t_8__203_ = t_7__203_ | t_7__331_;
  assign t_8__202_ = t_7__202_ | t_7__330_;
  assign t_8__201_ = t_7__201_ | t_7__329_;
  assign t_8__200_ = t_7__200_ | t_7__328_;
  assign t_8__199_ = t_7__199_ | t_7__327_;
  assign t_8__198_ = t_7__198_ | t_7__326_;
  assign t_8__197_ = t_7__197_ | t_7__325_;
  assign t_8__196_ = t_7__196_ | t_7__324_;
  assign t_8__195_ = t_7__195_ | t_7__323_;
  assign t_8__194_ = t_7__194_ | t_7__322_;
  assign t_8__193_ = t_7__193_ | t_7__321_;
  assign t_8__192_ = t_7__192_ | t_7__320_;
  assign t_8__191_ = t_7__191_ | t_7__319_;
  assign t_8__190_ = t_7__190_ | t_7__318_;
  assign t_8__189_ = t_7__189_ | t_7__317_;
  assign t_8__188_ = t_7__188_ | t_7__316_;
  assign t_8__187_ = t_7__187_ | t_7__315_;
  assign t_8__186_ = t_7__186_ | t_7__314_;
  assign t_8__185_ = t_7__185_ | t_7__313_;
  assign t_8__184_ = t_7__184_ | t_7__312_;
  assign t_8__183_ = t_7__183_ | t_7__311_;
  assign t_8__182_ = t_7__182_ | t_7__310_;
  assign t_8__181_ = t_7__181_ | t_7__309_;
  assign t_8__180_ = t_7__180_ | t_7__308_;
  assign t_8__179_ = t_7__179_ | t_7__307_;
  assign t_8__178_ = t_7__178_ | t_7__306_;
  assign t_8__177_ = t_7__177_ | t_7__305_;
  assign t_8__176_ = t_7__176_ | t_7__304_;
  assign t_8__175_ = t_7__175_ | t_7__303_;
  assign t_8__174_ = t_7__174_ | t_7__302_;
  assign t_8__173_ = t_7__173_ | t_7__301_;
  assign t_8__172_ = t_7__172_ | t_7__300_;
  assign t_8__171_ = t_7__171_ | t_7__299_;
  assign t_8__170_ = t_7__170_ | t_7__298_;
  assign t_8__169_ = t_7__169_ | t_7__297_;
  assign t_8__168_ = t_7__168_ | t_7__296_;
  assign t_8__167_ = t_7__167_ | t_7__295_;
  assign t_8__166_ = t_7__166_ | t_7__294_;
  assign t_8__165_ = t_7__165_ | t_7__293_;
  assign t_8__164_ = t_7__164_ | t_7__292_;
  assign t_8__163_ = t_7__163_ | t_7__291_;
  assign t_8__162_ = t_7__162_ | t_7__290_;
  assign t_8__161_ = t_7__161_ | t_7__289_;
  assign t_8__160_ = t_7__160_ | t_7__288_;
  assign t_8__159_ = t_7__159_ | t_7__287_;
  assign t_8__158_ = t_7__158_ | t_7__286_;
  assign t_8__157_ = t_7__157_ | t_7__285_;
  assign t_8__156_ = t_7__156_ | t_7__284_;
  assign t_8__155_ = t_7__155_ | t_7__283_;
  assign t_8__154_ = t_7__154_ | t_7__282_;
  assign t_8__153_ = t_7__153_ | t_7__281_;
  assign t_8__152_ = t_7__152_ | t_7__280_;
  assign t_8__151_ = t_7__151_ | t_7__279_;
  assign t_8__150_ = t_7__150_ | t_7__278_;
  assign t_8__149_ = t_7__149_ | t_7__277_;
  assign t_8__148_ = t_7__148_ | t_7__276_;
  assign t_8__147_ = t_7__147_ | t_7__275_;
  assign t_8__146_ = t_7__146_ | t_7__274_;
  assign t_8__145_ = t_7__145_ | t_7__273_;
  assign t_8__144_ = t_7__144_ | t_7__272_;
  assign t_8__143_ = t_7__143_ | t_7__271_;
  assign t_8__142_ = t_7__142_ | t_7__270_;
  assign t_8__141_ = t_7__141_ | t_7__269_;
  assign t_8__140_ = t_7__140_ | t_7__268_;
  assign t_8__139_ = t_7__139_ | t_7__267_;
  assign t_8__138_ = t_7__138_ | t_7__266_;
  assign t_8__137_ = t_7__137_ | t_7__265_;
  assign t_8__136_ = t_7__136_ | t_7__264_;
  assign t_8__135_ = t_7__135_ | t_7__263_;
  assign t_8__134_ = t_7__134_ | t_7__262_;
  assign t_8__133_ = t_7__133_ | t_7__261_;
  assign t_8__132_ = t_7__132_ | t_7__260_;
  assign t_8__131_ = t_7__131_ | t_7__259_;
  assign t_8__130_ = t_7__130_ | t_7__258_;
  assign t_8__129_ = t_7__129_ | t_7__257_;
  assign t_8__128_ = t_7__128_ | t_7__256_;
  assign t_8__127_ = t_7__127_ | t_7__255_;
  assign t_8__126_ = t_7__126_ | t_7__254_;
  assign t_8__125_ = t_7__125_ | t_7__253_;
  assign t_8__124_ = t_7__124_ | t_7__252_;
  assign t_8__123_ = t_7__123_ | t_7__251_;
  assign t_8__122_ = t_7__122_ | t_7__250_;
  assign t_8__121_ = t_7__121_ | t_7__249_;
  assign t_8__120_ = t_7__120_ | t_7__248_;
  assign t_8__119_ = t_7__119_ | t_7__247_;
  assign t_8__118_ = t_7__118_ | t_7__246_;
  assign t_8__117_ = t_7__117_ | t_7__245_;
  assign t_8__116_ = t_7__116_ | t_7__244_;
  assign t_8__115_ = t_7__115_ | t_7__243_;
  assign t_8__114_ = t_7__114_ | t_7__242_;
  assign t_8__113_ = t_7__113_ | t_7__241_;
  assign t_8__112_ = t_7__112_ | t_7__240_;
  assign t_8__111_ = t_7__111_ | t_7__239_;
  assign t_8__110_ = t_7__110_ | t_7__238_;
  assign t_8__109_ = t_7__109_ | t_7__237_;
  assign t_8__108_ = t_7__108_ | t_7__236_;
  assign t_8__107_ = t_7__107_ | t_7__235_;
  assign t_8__106_ = t_7__106_ | t_7__234_;
  assign t_8__105_ = t_7__105_ | t_7__233_;
  assign t_8__104_ = t_7__104_ | t_7__232_;
  assign t_8__103_ = t_7__103_ | t_7__231_;
  assign t_8__102_ = t_7__102_ | t_7__230_;
  assign t_8__101_ = t_7__101_ | t_7__229_;
  assign t_8__100_ = t_7__100_ | t_7__228_;
  assign t_8__99_ = t_7__99_ | t_7__227_;
  assign t_8__98_ = t_7__98_ | t_7__226_;
  assign t_8__97_ = t_7__97_ | t_7__225_;
  assign t_8__96_ = t_7__96_ | t_7__224_;
  assign t_8__95_ = t_7__95_ | t_7__223_;
  assign t_8__94_ = t_7__94_ | t_7__222_;
  assign t_8__93_ = t_7__93_ | t_7__221_;
  assign t_8__92_ = t_7__92_ | t_7__220_;
  assign t_8__91_ = t_7__91_ | t_7__219_;
  assign t_8__90_ = t_7__90_ | t_7__218_;
  assign t_8__89_ = t_7__89_ | t_7__217_;
  assign t_8__88_ = t_7__88_ | t_7__216_;
  assign t_8__87_ = t_7__87_ | t_7__215_;
  assign t_8__86_ = t_7__86_ | t_7__214_;
  assign t_8__85_ = t_7__85_ | t_7__213_;
  assign t_8__84_ = t_7__84_ | t_7__212_;
  assign t_8__83_ = t_7__83_ | t_7__211_;
  assign t_8__82_ = t_7__82_ | t_7__210_;
  assign t_8__81_ = t_7__81_ | t_7__209_;
  assign t_8__80_ = t_7__80_ | t_7__208_;
  assign t_8__79_ = t_7__79_ | t_7__207_;
  assign t_8__78_ = t_7__78_ | t_7__206_;
  assign t_8__77_ = t_7__77_ | t_7__205_;
  assign t_8__76_ = t_7__76_ | t_7__204_;
  assign t_8__75_ = t_7__75_ | t_7__203_;
  assign t_8__74_ = t_7__74_ | t_7__202_;
  assign t_8__73_ = t_7__73_ | t_7__201_;
  assign t_8__72_ = t_7__72_ | t_7__200_;
  assign t_8__71_ = t_7__71_ | t_7__199_;
  assign t_8__70_ = t_7__70_ | t_7__198_;
  assign t_8__69_ = t_7__69_ | t_7__197_;
  assign t_8__68_ = t_7__68_ | t_7__196_;
  assign t_8__67_ = t_7__67_ | t_7__195_;
  assign t_8__66_ = t_7__66_ | t_7__194_;
  assign t_8__65_ = t_7__65_ | t_7__193_;
  assign t_8__64_ = t_7__64_ | t_7__192_;
  assign t_8__63_ = t_7__63_ | t_7__191_;
  assign t_8__62_ = t_7__62_ | t_7__190_;
  assign t_8__61_ = t_7__61_ | t_7__189_;
  assign t_8__60_ = t_7__60_ | t_7__188_;
  assign t_8__59_ = t_7__59_ | t_7__187_;
  assign t_8__58_ = t_7__58_ | t_7__186_;
  assign t_8__57_ = t_7__57_ | t_7__185_;
  assign t_8__56_ = t_7__56_ | t_7__184_;
  assign t_8__55_ = t_7__55_ | t_7__183_;
  assign t_8__54_ = t_7__54_ | t_7__182_;
  assign t_8__53_ = t_7__53_ | t_7__181_;
  assign t_8__52_ = t_7__52_ | t_7__180_;
  assign t_8__51_ = t_7__51_ | t_7__179_;
  assign t_8__50_ = t_7__50_ | t_7__178_;
  assign t_8__49_ = t_7__49_ | t_7__177_;
  assign t_8__48_ = t_7__48_ | t_7__176_;
  assign t_8__47_ = t_7__47_ | t_7__175_;
  assign t_8__46_ = t_7__46_ | t_7__174_;
  assign t_8__45_ = t_7__45_ | t_7__173_;
  assign t_8__44_ = t_7__44_ | t_7__172_;
  assign t_8__43_ = t_7__43_ | t_7__171_;
  assign t_8__42_ = t_7__42_ | t_7__170_;
  assign t_8__41_ = t_7__41_ | t_7__169_;
  assign t_8__40_ = t_7__40_ | t_7__168_;
  assign t_8__39_ = t_7__39_ | t_7__167_;
  assign t_8__38_ = t_7__38_ | t_7__166_;
  assign t_8__37_ = t_7__37_ | t_7__165_;
  assign t_8__36_ = t_7__36_ | t_7__164_;
  assign t_8__35_ = t_7__35_ | t_7__163_;
  assign t_8__34_ = t_7__34_ | t_7__162_;
  assign t_8__33_ = t_7__33_ | t_7__161_;
  assign t_8__32_ = t_7__32_ | t_7__160_;
  assign t_8__31_ = t_7__31_ | t_7__159_;
  assign t_8__30_ = t_7__30_ | t_7__158_;
  assign t_8__29_ = t_7__29_ | t_7__157_;
  assign t_8__28_ = t_7__28_ | t_7__156_;
  assign t_8__27_ = t_7__27_ | t_7__155_;
  assign t_8__26_ = t_7__26_ | t_7__154_;
  assign t_8__25_ = t_7__25_ | t_7__153_;
  assign t_8__24_ = t_7__24_ | t_7__152_;
  assign t_8__23_ = t_7__23_ | t_7__151_;
  assign t_8__22_ = t_7__22_ | t_7__150_;
  assign t_8__21_ = t_7__21_ | t_7__149_;
  assign t_8__20_ = t_7__20_ | t_7__148_;
  assign t_8__19_ = t_7__19_ | t_7__147_;
  assign t_8__18_ = t_7__18_ | t_7__146_;
  assign t_8__17_ = t_7__17_ | t_7__145_;
  assign t_8__16_ = t_7__16_ | t_7__144_;
  assign t_8__15_ = t_7__15_ | t_7__143_;
  assign t_8__14_ = t_7__14_ | t_7__142_;
  assign t_8__13_ = t_7__13_ | t_7__141_;
  assign t_8__12_ = t_7__12_ | t_7__140_;
  assign t_8__11_ = t_7__11_ | t_7__139_;
  assign t_8__10_ = t_7__10_ | t_7__138_;
  assign t_8__9_ = t_7__9_ | t_7__137_;
  assign t_8__8_ = t_7__8_ | t_7__136_;
  assign t_8__7_ = t_7__7_ | t_7__135_;
  assign t_8__6_ = t_7__6_ | t_7__134_;
  assign t_8__5_ = t_7__5_ | t_7__133_;
  assign t_8__4_ = t_7__4_ | t_7__132_;
  assign t_8__3_ = t_7__3_ | t_7__131_;
  assign t_8__2_ = t_7__2_ | t_7__130_;
  assign t_8__1_ = t_7__1_ | t_7__129_;
  assign t_8__0_ = t_7__0_ | t_7__128_;
  assign o[0] = t_8__511_ | 1'b0;
  assign o[1] = t_8__510_ | 1'b0;
  assign o[2] = t_8__509_ | 1'b0;
  assign o[3] = t_8__508_ | 1'b0;
  assign o[4] = t_8__507_ | 1'b0;
  assign o[5] = t_8__506_ | 1'b0;
  assign o[6] = t_8__505_ | 1'b0;
  assign o[7] = t_8__504_ | 1'b0;
  assign o[8] = t_8__503_ | 1'b0;
  assign o[9] = t_8__502_ | 1'b0;
  assign o[10] = t_8__501_ | 1'b0;
  assign o[11] = t_8__500_ | 1'b0;
  assign o[12] = t_8__499_ | 1'b0;
  assign o[13] = t_8__498_ | 1'b0;
  assign o[14] = t_8__497_ | 1'b0;
  assign o[15] = t_8__496_ | 1'b0;
  assign o[16] = t_8__495_ | 1'b0;
  assign o[17] = t_8__494_ | 1'b0;
  assign o[18] = t_8__493_ | 1'b0;
  assign o[19] = t_8__492_ | 1'b0;
  assign o[20] = t_8__491_ | 1'b0;
  assign o[21] = t_8__490_ | 1'b0;
  assign o[22] = t_8__489_ | 1'b0;
  assign o[23] = t_8__488_ | 1'b0;
  assign o[24] = t_8__487_ | 1'b0;
  assign o[25] = t_8__486_ | 1'b0;
  assign o[26] = t_8__485_ | 1'b0;
  assign o[27] = t_8__484_ | 1'b0;
  assign o[28] = t_8__483_ | 1'b0;
  assign o[29] = t_8__482_ | 1'b0;
  assign o[30] = t_8__481_ | 1'b0;
  assign o[31] = t_8__480_ | 1'b0;
  assign o[32] = t_8__479_ | 1'b0;
  assign o[33] = t_8__478_ | 1'b0;
  assign o[34] = t_8__477_ | 1'b0;
  assign o[35] = t_8__476_ | 1'b0;
  assign o[36] = t_8__475_ | 1'b0;
  assign o[37] = t_8__474_ | 1'b0;
  assign o[38] = t_8__473_ | 1'b0;
  assign o[39] = t_8__472_ | 1'b0;
  assign o[40] = t_8__471_ | 1'b0;
  assign o[41] = t_8__470_ | 1'b0;
  assign o[42] = t_8__469_ | 1'b0;
  assign o[43] = t_8__468_ | 1'b0;
  assign o[44] = t_8__467_ | 1'b0;
  assign o[45] = t_8__466_ | 1'b0;
  assign o[46] = t_8__465_ | 1'b0;
  assign o[47] = t_8__464_ | 1'b0;
  assign o[48] = t_8__463_ | 1'b0;
  assign o[49] = t_8__462_ | 1'b0;
  assign o[50] = t_8__461_ | 1'b0;
  assign o[51] = t_8__460_ | 1'b0;
  assign o[52] = t_8__459_ | 1'b0;
  assign o[53] = t_8__458_ | 1'b0;
  assign o[54] = t_8__457_ | 1'b0;
  assign o[55] = t_8__456_ | 1'b0;
  assign o[56] = t_8__455_ | 1'b0;
  assign o[57] = t_8__454_ | 1'b0;
  assign o[58] = t_8__453_ | 1'b0;
  assign o[59] = t_8__452_ | 1'b0;
  assign o[60] = t_8__451_ | 1'b0;
  assign o[61] = t_8__450_ | 1'b0;
  assign o[62] = t_8__449_ | 1'b0;
  assign o[63] = t_8__448_ | 1'b0;
  assign o[64] = t_8__447_ | 1'b0;
  assign o[65] = t_8__446_ | 1'b0;
  assign o[66] = t_8__445_ | 1'b0;
  assign o[67] = t_8__444_ | 1'b0;
  assign o[68] = t_8__443_ | 1'b0;
  assign o[69] = t_8__442_ | 1'b0;
  assign o[70] = t_8__441_ | 1'b0;
  assign o[71] = t_8__440_ | 1'b0;
  assign o[72] = t_8__439_ | 1'b0;
  assign o[73] = t_8__438_ | 1'b0;
  assign o[74] = t_8__437_ | 1'b0;
  assign o[75] = t_8__436_ | 1'b0;
  assign o[76] = t_8__435_ | 1'b0;
  assign o[77] = t_8__434_ | 1'b0;
  assign o[78] = t_8__433_ | 1'b0;
  assign o[79] = t_8__432_ | 1'b0;
  assign o[80] = t_8__431_ | 1'b0;
  assign o[81] = t_8__430_ | 1'b0;
  assign o[82] = t_8__429_ | 1'b0;
  assign o[83] = t_8__428_ | 1'b0;
  assign o[84] = t_8__427_ | 1'b0;
  assign o[85] = t_8__426_ | 1'b0;
  assign o[86] = t_8__425_ | 1'b0;
  assign o[87] = t_8__424_ | 1'b0;
  assign o[88] = t_8__423_ | 1'b0;
  assign o[89] = t_8__422_ | 1'b0;
  assign o[90] = t_8__421_ | 1'b0;
  assign o[91] = t_8__420_ | 1'b0;
  assign o[92] = t_8__419_ | 1'b0;
  assign o[93] = t_8__418_ | 1'b0;
  assign o[94] = t_8__417_ | 1'b0;
  assign o[95] = t_8__416_ | 1'b0;
  assign o[96] = t_8__415_ | 1'b0;
  assign o[97] = t_8__414_ | 1'b0;
  assign o[98] = t_8__413_ | 1'b0;
  assign o[99] = t_8__412_ | 1'b0;
  assign o[100] = t_8__411_ | 1'b0;
  assign o[101] = t_8__410_ | 1'b0;
  assign o[102] = t_8__409_ | 1'b0;
  assign o[103] = t_8__408_ | 1'b0;
  assign o[104] = t_8__407_ | 1'b0;
  assign o[105] = t_8__406_ | 1'b0;
  assign o[106] = t_8__405_ | 1'b0;
  assign o[107] = t_8__404_ | 1'b0;
  assign o[108] = t_8__403_ | 1'b0;
  assign o[109] = t_8__402_ | 1'b0;
  assign o[110] = t_8__401_ | 1'b0;
  assign o[111] = t_8__400_ | 1'b0;
  assign o[112] = t_8__399_ | 1'b0;
  assign o[113] = t_8__398_ | 1'b0;
  assign o[114] = t_8__397_ | 1'b0;
  assign o[115] = t_8__396_ | 1'b0;
  assign o[116] = t_8__395_ | 1'b0;
  assign o[117] = t_8__394_ | 1'b0;
  assign o[118] = t_8__393_ | 1'b0;
  assign o[119] = t_8__392_ | 1'b0;
  assign o[120] = t_8__391_ | 1'b0;
  assign o[121] = t_8__390_ | 1'b0;
  assign o[122] = t_8__389_ | 1'b0;
  assign o[123] = t_8__388_ | 1'b0;
  assign o[124] = t_8__387_ | 1'b0;
  assign o[125] = t_8__386_ | 1'b0;
  assign o[126] = t_8__385_ | 1'b0;
  assign o[127] = t_8__384_ | 1'b0;
  assign o[128] = t_8__383_ | 1'b0;
  assign o[129] = t_8__382_ | 1'b0;
  assign o[130] = t_8__381_ | 1'b0;
  assign o[131] = t_8__380_ | 1'b0;
  assign o[132] = t_8__379_ | 1'b0;
  assign o[133] = t_8__378_ | 1'b0;
  assign o[134] = t_8__377_ | 1'b0;
  assign o[135] = t_8__376_ | 1'b0;
  assign o[136] = t_8__375_ | 1'b0;
  assign o[137] = t_8__374_ | 1'b0;
  assign o[138] = t_8__373_ | 1'b0;
  assign o[139] = t_8__372_ | 1'b0;
  assign o[140] = t_8__371_ | 1'b0;
  assign o[141] = t_8__370_ | 1'b0;
  assign o[142] = t_8__369_ | 1'b0;
  assign o[143] = t_8__368_ | 1'b0;
  assign o[144] = t_8__367_ | 1'b0;
  assign o[145] = t_8__366_ | 1'b0;
  assign o[146] = t_8__365_ | 1'b0;
  assign o[147] = t_8__364_ | 1'b0;
  assign o[148] = t_8__363_ | 1'b0;
  assign o[149] = t_8__362_ | 1'b0;
  assign o[150] = t_8__361_ | 1'b0;
  assign o[151] = t_8__360_ | 1'b0;
  assign o[152] = t_8__359_ | 1'b0;
  assign o[153] = t_8__358_ | 1'b0;
  assign o[154] = t_8__357_ | 1'b0;
  assign o[155] = t_8__356_ | 1'b0;
  assign o[156] = t_8__355_ | 1'b0;
  assign o[157] = t_8__354_ | 1'b0;
  assign o[158] = t_8__353_ | 1'b0;
  assign o[159] = t_8__352_ | 1'b0;
  assign o[160] = t_8__351_ | 1'b0;
  assign o[161] = t_8__350_ | 1'b0;
  assign o[162] = t_8__349_ | 1'b0;
  assign o[163] = t_8__348_ | 1'b0;
  assign o[164] = t_8__347_ | 1'b0;
  assign o[165] = t_8__346_ | 1'b0;
  assign o[166] = t_8__345_ | 1'b0;
  assign o[167] = t_8__344_ | 1'b0;
  assign o[168] = t_8__343_ | 1'b0;
  assign o[169] = t_8__342_ | 1'b0;
  assign o[170] = t_8__341_ | 1'b0;
  assign o[171] = t_8__340_ | 1'b0;
  assign o[172] = t_8__339_ | 1'b0;
  assign o[173] = t_8__338_ | 1'b0;
  assign o[174] = t_8__337_ | 1'b0;
  assign o[175] = t_8__336_ | 1'b0;
  assign o[176] = t_8__335_ | 1'b0;
  assign o[177] = t_8__334_ | 1'b0;
  assign o[178] = t_8__333_ | 1'b0;
  assign o[179] = t_8__332_ | 1'b0;
  assign o[180] = t_8__331_ | 1'b0;
  assign o[181] = t_8__330_ | 1'b0;
  assign o[182] = t_8__329_ | 1'b0;
  assign o[183] = t_8__328_ | 1'b0;
  assign o[184] = t_8__327_ | 1'b0;
  assign o[185] = t_8__326_ | 1'b0;
  assign o[186] = t_8__325_ | 1'b0;
  assign o[187] = t_8__324_ | 1'b0;
  assign o[188] = t_8__323_ | 1'b0;
  assign o[189] = t_8__322_ | 1'b0;
  assign o[190] = t_8__321_ | 1'b0;
  assign o[191] = t_8__320_ | 1'b0;
  assign o[192] = t_8__319_ | 1'b0;
  assign o[193] = t_8__318_ | 1'b0;
  assign o[194] = t_8__317_ | 1'b0;
  assign o[195] = t_8__316_ | 1'b0;
  assign o[196] = t_8__315_ | 1'b0;
  assign o[197] = t_8__314_ | 1'b0;
  assign o[198] = t_8__313_ | 1'b0;
  assign o[199] = t_8__312_ | 1'b0;
  assign o[200] = t_8__311_ | 1'b0;
  assign o[201] = t_8__310_ | 1'b0;
  assign o[202] = t_8__309_ | 1'b0;
  assign o[203] = t_8__308_ | 1'b0;
  assign o[204] = t_8__307_ | 1'b0;
  assign o[205] = t_8__306_ | 1'b0;
  assign o[206] = t_8__305_ | 1'b0;
  assign o[207] = t_8__304_ | 1'b0;
  assign o[208] = t_8__303_ | 1'b0;
  assign o[209] = t_8__302_ | 1'b0;
  assign o[210] = t_8__301_ | 1'b0;
  assign o[211] = t_8__300_ | 1'b0;
  assign o[212] = t_8__299_ | 1'b0;
  assign o[213] = t_8__298_ | 1'b0;
  assign o[214] = t_8__297_ | 1'b0;
  assign o[215] = t_8__296_ | 1'b0;
  assign o[216] = t_8__295_ | 1'b0;
  assign o[217] = t_8__294_ | 1'b0;
  assign o[218] = t_8__293_ | 1'b0;
  assign o[219] = t_8__292_ | 1'b0;
  assign o[220] = t_8__291_ | 1'b0;
  assign o[221] = t_8__290_ | 1'b0;
  assign o[222] = t_8__289_ | 1'b0;
  assign o[223] = t_8__288_ | 1'b0;
  assign o[224] = t_8__287_ | 1'b0;
  assign o[225] = t_8__286_ | 1'b0;
  assign o[226] = t_8__285_ | 1'b0;
  assign o[227] = t_8__284_ | 1'b0;
  assign o[228] = t_8__283_ | 1'b0;
  assign o[229] = t_8__282_ | 1'b0;
  assign o[230] = t_8__281_ | 1'b0;
  assign o[231] = t_8__280_ | 1'b0;
  assign o[232] = t_8__279_ | 1'b0;
  assign o[233] = t_8__278_ | 1'b0;
  assign o[234] = t_8__277_ | 1'b0;
  assign o[235] = t_8__276_ | 1'b0;
  assign o[236] = t_8__275_ | 1'b0;
  assign o[237] = t_8__274_ | 1'b0;
  assign o[238] = t_8__273_ | 1'b0;
  assign o[239] = t_8__272_ | 1'b0;
  assign o[240] = t_8__271_ | 1'b0;
  assign o[241] = t_8__270_ | 1'b0;
  assign o[242] = t_8__269_ | 1'b0;
  assign o[243] = t_8__268_ | 1'b0;
  assign o[244] = t_8__267_ | 1'b0;
  assign o[245] = t_8__266_ | 1'b0;
  assign o[246] = t_8__265_ | 1'b0;
  assign o[247] = t_8__264_ | 1'b0;
  assign o[248] = t_8__263_ | 1'b0;
  assign o[249] = t_8__262_ | 1'b0;
  assign o[250] = t_8__261_ | 1'b0;
  assign o[251] = t_8__260_ | 1'b0;
  assign o[252] = t_8__259_ | 1'b0;
  assign o[253] = t_8__258_ | 1'b0;
  assign o[254] = t_8__257_ | 1'b0;
  assign o[255] = t_8__256_ | 1'b0;
  assign o[256] = t_8__255_ | t_8__511_;
  assign o[257] = t_8__254_ | t_8__510_;
  assign o[258] = t_8__253_ | t_8__509_;
  assign o[259] = t_8__252_ | t_8__508_;
  assign o[260] = t_8__251_ | t_8__507_;
  assign o[261] = t_8__250_ | t_8__506_;
  assign o[262] = t_8__249_ | t_8__505_;
  assign o[263] = t_8__248_ | t_8__504_;
  assign o[264] = t_8__247_ | t_8__503_;
  assign o[265] = t_8__246_ | t_8__502_;
  assign o[266] = t_8__245_ | t_8__501_;
  assign o[267] = t_8__244_ | t_8__500_;
  assign o[268] = t_8__243_ | t_8__499_;
  assign o[269] = t_8__242_ | t_8__498_;
  assign o[270] = t_8__241_ | t_8__497_;
  assign o[271] = t_8__240_ | t_8__496_;
  assign o[272] = t_8__239_ | t_8__495_;
  assign o[273] = t_8__238_ | t_8__494_;
  assign o[274] = t_8__237_ | t_8__493_;
  assign o[275] = t_8__236_ | t_8__492_;
  assign o[276] = t_8__235_ | t_8__491_;
  assign o[277] = t_8__234_ | t_8__490_;
  assign o[278] = t_8__233_ | t_8__489_;
  assign o[279] = t_8__232_ | t_8__488_;
  assign o[280] = t_8__231_ | t_8__487_;
  assign o[281] = t_8__230_ | t_8__486_;
  assign o[282] = t_8__229_ | t_8__485_;
  assign o[283] = t_8__228_ | t_8__484_;
  assign o[284] = t_8__227_ | t_8__483_;
  assign o[285] = t_8__226_ | t_8__482_;
  assign o[286] = t_8__225_ | t_8__481_;
  assign o[287] = t_8__224_ | t_8__480_;
  assign o[288] = t_8__223_ | t_8__479_;
  assign o[289] = t_8__222_ | t_8__478_;
  assign o[290] = t_8__221_ | t_8__477_;
  assign o[291] = t_8__220_ | t_8__476_;
  assign o[292] = t_8__219_ | t_8__475_;
  assign o[293] = t_8__218_ | t_8__474_;
  assign o[294] = t_8__217_ | t_8__473_;
  assign o[295] = t_8__216_ | t_8__472_;
  assign o[296] = t_8__215_ | t_8__471_;
  assign o[297] = t_8__214_ | t_8__470_;
  assign o[298] = t_8__213_ | t_8__469_;
  assign o[299] = t_8__212_ | t_8__468_;
  assign o[300] = t_8__211_ | t_8__467_;
  assign o[301] = t_8__210_ | t_8__466_;
  assign o[302] = t_8__209_ | t_8__465_;
  assign o[303] = t_8__208_ | t_8__464_;
  assign o[304] = t_8__207_ | t_8__463_;
  assign o[305] = t_8__206_ | t_8__462_;
  assign o[306] = t_8__205_ | t_8__461_;
  assign o[307] = t_8__204_ | t_8__460_;
  assign o[308] = t_8__203_ | t_8__459_;
  assign o[309] = t_8__202_ | t_8__458_;
  assign o[310] = t_8__201_ | t_8__457_;
  assign o[311] = t_8__200_ | t_8__456_;
  assign o[312] = t_8__199_ | t_8__455_;
  assign o[313] = t_8__198_ | t_8__454_;
  assign o[314] = t_8__197_ | t_8__453_;
  assign o[315] = t_8__196_ | t_8__452_;
  assign o[316] = t_8__195_ | t_8__451_;
  assign o[317] = t_8__194_ | t_8__450_;
  assign o[318] = t_8__193_ | t_8__449_;
  assign o[319] = t_8__192_ | t_8__448_;
  assign o[320] = t_8__191_ | t_8__447_;
  assign o[321] = t_8__190_ | t_8__446_;
  assign o[322] = t_8__189_ | t_8__445_;
  assign o[323] = t_8__188_ | t_8__444_;
  assign o[324] = t_8__187_ | t_8__443_;
  assign o[325] = t_8__186_ | t_8__442_;
  assign o[326] = t_8__185_ | t_8__441_;
  assign o[327] = t_8__184_ | t_8__440_;
  assign o[328] = t_8__183_ | t_8__439_;
  assign o[329] = t_8__182_ | t_8__438_;
  assign o[330] = t_8__181_ | t_8__437_;
  assign o[331] = t_8__180_ | t_8__436_;
  assign o[332] = t_8__179_ | t_8__435_;
  assign o[333] = t_8__178_ | t_8__434_;
  assign o[334] = t_8__177_ | t_8__433_;
  assign o[335] = t_8__176_ | t_8__432_;
  assign o[336] = t_8__175_ | t_8__431_;
  assign o[337] = t_8__174_ | t_8__430_;
  assign o[338] = t_8__173_ | t_8__429_;
  assign o[339] = t_8__172_ | t_8__428_;
  assign o[340] = t_8__171_ | t_8__427_;
  assign o[341] = t_8__170_ | t_8__426_;
  assign o[342] = t_8__169_ | t_8__425_;
  assign o[343] = t_8__168_ | t_8__424_;
  assign o[344] = t_8__167_ | t_8__423_;
  assign o[345] = t_8__166_ | t_8__422_;
  assign o[346] = t_8__165_ | t_8__421_;
  assign o[347] = t_8__164_ | t_8__420_;
  assign o[348] = t_8__163_ | t_8__419_;
  assign o[349] = t_8__162_ | t_8__418_;
  assign o[350] = t_8__161_ | t_8__417_;
  assign o[351] = t_8__160_ | t_8__416_;
  assign o[352] = t_8__159_ | t_8__415_;
  assign o[353] = t_8__158_ | t_8__414_;
  assign o[354] = t_8__157_ | t_8__413_;
  assign o[355] = t_8__156_ | t_8__412_;
  assign o[356] = t_8__155_ | t_8__411_;
  assign o[357] = t_8__154_ | t_8__410_;
  assign o[358] = t_8__153_ | t_8__409_;
  assign o[359] = t_8__152_ | t_8__408_;
  assign o[360] = t_8__151_ | t_8__407_;
  assign o[361] = t_8__150_ | t_8__406_;
  assign o[362] = t_8__149_ | t_8__405_;
  assign o[363] = t_8__148_ | t_8__404_;
  assign o[364] = t_8__147_ | t_8__403_;
  assign o[365] = t_8__146_ | t_8__402_;
  assign o[366] = t_8__145_ | t_8__401_;
  assign o[367] = t_8__144_ | t_8__400_;
  assign o[368] = t_8__143_ | t_8__399_;
  assign o[369] = t_8__142_ | t_8__398_;
  assign o[370] = t_8__141_ | t_8__397_;
  assign o[371] = t_8__140_ | t_8__396_;
  assign o[372] = t_8__139_ | t_8__395_;
  assign o[373] = t_8__138_ | t_8__394_;
  assign o[374] = t_8__137_ | t_8__393_;
  assign o[375] = t_8__136_ | t_8__392_;
  assign o[376] = t_8__135_ | t_8__391_;
  assign o[377] = t_8__134_ | t_8__390_;
  assign o[378] = t_8__133_ | t_8__389_;
  assign o[379] = t_8__132_ | t_8__388_;
  assign o[380] = t_8__131_ | t_8__387_;
  assign o[381] = t_8__130_ | t_8__386_;
  assign o[382] = t_8__129_ | t_8__385_;
  assign o[383] = t_8__128_ | t_8__384_;
  assign o[384] = t_8__127_ | t_8__383_;
  assign o[385] = t_8__126_ | t_8__382_;
  assign o[386] = t_8__125_ | t_8__381_;
  assign o[387] = t_8__124_ | t_8__380_;
  assign o[388] = t_8__123_ | t_8__379_;
  assign o[389] = t_8__122_ | t_8__378_;
  assign o[390] = t_8__121_ | t_8__377_;
  assign o[391] = t_8__120_ | t_8__376_;
  assign o[392] = t_8__119_ | t_8__375_;
  assign o[393] = t_8__118_ | t_8__374_;
  assign o[394] = t_8__117_ | t_8__373_;
  assign o[395] = t_8__116_ | t_8__372_;
  assign o[396] = t_8__115_ | t_8__371_;
  assign o[397] = t_8__114_ | t_8__370_;
  assign o[398] = t_8__113_ | t_8__369_;
  assign o[399] = t_8__112_ | t_8__368_;
  assign o[400] = t_8__111_ | t_8__367_;
  assign o[401] = t_8__110_ | t_8__366_;
  assign o[402] = t_8__109_ | t_8__365_;
  assign o[403] = t_8__108_ | t_8__364_;
  assign o[404] = t_8__107_ | t_8__363_;
  assign o[405] = t_8__106_ | t_8__362_;
  assign o[406] = t_8__105_ | t_8__361_;
  assign o[407] = t_8__104_ | t_8__360_;
  assign o[408] = t_8__103_ | t_8__359_;
  assign o[409] = t_8__102_ | t_8__358_;
  assign o[410] = t_8__101_ | t_8__357_;
  assign o[411] = t_8__100_ | t_8__356_;
  assign o[412] = t_8__99_ | t_8__355_;
  assign o[413] = t_8__98_ | t_8__354_;
  assign o[414] = t_8__97_ | t_8__353_;
  assign o[415] = t_8__96_ | t_8__352_;
  assign o[416] = t_8__95_ | t_8__351_;
  assign o[417] = t_8__94_ | t_8__350_;
  assign o[418] = t_8__93_ | t_8__349_;
  assign o[419] = t_8__92_ | t_8__348_;
  assign o[420] = t_8__91_ | t_8__347_;
  assign o[421] = t_8__90_ | t_8__346_;
  assign o[422] = t_8__89_ | t_8__345_;
  assign o[423] = t_8__88_ | t_8__344_;
  assign o[424] = t_8__87_ | t_8__343_;
  assign o[425] = t_8__86_ | t_8__342_;
  assign o[426] = t_8__85_ | t_8__341_;
  assign o[427] = t_8__84_ | t_8__340_;
  assign o[428] = t_8__83_ | t_8__339_;
  assign o[429] = t_8__82_ | t_8__338_;
  assign o[430] = t_8__81_ | t_8__337_;
  assign o[431] = t_8__80_ | t_8__336_;
  assign o[432] = t_8__79_ | t_8__335_;
  assign o[433] = t_8__78_ | t_8__334_;
  assign o[434] = t_8__77_ | t_8__333_;
  assign o[435] = t_8__76_ | t_8__332_;
  assign o[436] = t_8__75_ | t_8__331_;
  assign o[437] = t_8__74_ | t_8__330_;
  assign o[438] = t_8__73_ | t_8__329_;
  assign o[439] = t_8__72_ | t_8__328_;
  assign o[440] = t_8__71_ | t_8__327_;
  assign o[441] = t_8__70_ | t_8__326_;
  assign o[442] = t_8__69_ | t_8__325_;
  assign o[443] = t_8__68_ | t_8__324_;
  assign o[444] = t_8__67_ | t_8__323_;
  assign o[445] = t_8__66_ | t_8__322_;
  assign o[446] = t_8__65_ | t_8__321_;
  assign o[447] = t_8__64_ | t_8__320_;
  assign o[448] = t_8__63_ | t_8__319_;
  assign o[449] = t_8__62_ | t_8__318_;
  assign o[450] = t_8__61_ | t_8__317_;
  assign o[451] = t_8__60_ | t_8__316_;
  assign o[452] = t_8__59_ | t_8__315_;
  assign o[453] = t_8__58_ | t_8__314_;
  assign o[454] = t_8__57_ | t_8__313_;
  assign o[455] = t_8__56_ | t_8__312_;
  assign o[456] = t_8__55_ | t_8__311_;
  assign o[457] = t_8__54_ | t_8__310_;
  assign o[458] = t_8__53_ | t_8__309_;
  assign o[459] = t_8__52_ | t_8__308_;
  assign o[460] = t_8__51_ | t_8__307_;
  assign o[461] = t_8__50_ | t_8__306_;
  assign o[462] = t_8__49_ | t_8__305_;
  assign o[463] = t_8__48_ | t_8__304_;
  assign o[464] = t_8__47_ | t_8__303_;
  assign o[465] = t_8__46_ | t_8__302_;
  assign o[466] = t_8__45_ | t_8__301_;
  assign o[467] = t_8__44_ | t_8__300_;
  assign o[468] = t_8__43_ | t_8__299_;
  assign o[469] = t_8__42_ | t_8__298_;
  assign o[470] = t_8__41_ | t_8__297_;
  assign o[471] = t_8__40_ | t_8__296_;
  assign o[472] = t_8__39_ | t_8__295_;
  assign o[473] = t_8__38_ | t_8__294_;
  assign o[474] = t_8__37_ | t_8__293_;
  assign o[475] = t_8__36_ | t_8__292_;
  assign o[476] = t_8__35_ | t_8__291_;
  assign o[477] = t_8__34_ | t_8__290_;
  assign o[478] = t_8__33_ | t_8__289_;
  assign o[479] = t_8__32_ | t_8__288_;
  assign o[480] = t_8__31_ | t_8__287_;
  assign o[481] = t_8__30_ | t_8__286_;
  assign o[482] = t_8__29_ | t_8__285_;
  assign o[483] = t_8__28_ | t_8__284_;
  assign o[484] = t_8__27_ | t_8__283_;
  assign o[485] = t_8__26_ | t_8__282_;
  assign o[486] = t_8__25_ | t_8__281_;
  assign o[487] = t_8__24_ | t_8__280_;
  assign o[488] = t_8__23_ | t_8__279_;
  assign o[489] = t_8__22_ | t_8__278_;
  assign o[490] = t_8__21_ | t_8__277_;
  assign o[491] = t_8__20_ | t_8__276_;
  assign o[492] = t_8__19_ | t_8__275_;
  assign o[493] = t_8__18_ | t_8__274_;
  assign o[494] = t_8__17_ | t_8__273_;
  assign o[495] = t_8__16_ | t_8__272_;
  assign o[496] = t_8__15_ | t_8__271_;
  assign o[497] = t_8__14_ | t_8__270_;
  assign o[498] = t_8__13_ | t_8__269_;
  assign o[499] = t_8__12_ | t_8__268_;
  assign o[500] = t_8__11_ | t_8__267_;
  assign o[501] = t_8__10_ | t_8__266_;
  assign o[502] = t_8__9_ | t_8__265_;
  assign o[503] = t_8__8_ | t_8__264_;
  assign o[504] = t_8__7_ | t_8__263_;
  assign o[505] = t_8__6_ | t_8__262_;
  assign o[506] = t_8__5_ | t_8__261_;
  assign o[507] = t_8__4_ | t_8__260_;
  assign o[508] = t_8__3_ | t_8__259_;
  assign o[509] = t_8__2_ | t_8__258_;
  assign o[510] = t_8__1_ | t_8__257_;
  assign o[511] = t_8__0_ | t_8__256_;

endmodule



module bsg_priority_encode_one_hot_out_width_p512_lo_to_hi_p1
(
  i,
  o
);

  input [511:0] i;
  output [511:0] o;
  wire [511:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510;
  wire [511:1] scan_lo;

  bsg_scan_width_p512_or_p1_lo_to_hi_p1
  genblk1_scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[511] = scan_lo[511] & N0;
  assign N0 = ~scan_lo[510];
  assign o[510] = scan_lo[510] & N1;
  assign N1 = ~scan_lo[509];
  assign o[509] = scan_lo[509] & N2;
  assign N2 = ~scan_lo[508];
  assign o[508] = scan_lo[508] & N3;
  assign N3 = ~scan_lo[507];
  assign o[507] = scan_lo[507] & N4;
  assign N4 = ~scan_lo[506];
  assign o[506] = scan_lo[506] & N5;
  assign N5 = ~scan_lo[505];
  assign o[505] = scan_lo[505] & N6;
  assign N6 = ~scan_lo[504];
  assign o[504] = scan_lo[504] & N7;
  assign N7 = ~scan_lo[503];
  assign o[503] = scan_lo[503] & N8;
  assign N8 = ~scan_lo[502];
  assign o[502] = scan_lo[502] & N9;
  assign N9 = ~scan_lo[501];
  assign o[501] = scan_lo[501] & N10;
  assign N10 = ~scan_lo[500];
  assign o[500] = scan_lo[500] & N11;
  assign N11 = ~scan_lo[499];
  assign o[499] = scan_lo[499] & N12;
  assign N12 = ~scan_lo[498];
  assign o[498] = scan_lo[498] & N13;
  assign N13 = ~scan_lo[497];
  assign o[497] = scan_lo[497] & N14;
  assign N14 = ~scan_lo[496];
  assign o[496] = scan_lo[496] & N15;
  assign N15 = ~scan_lo[495];
  assign o[495] = scan_lo[495] & N16;
  assign N16 = ~scan_lo[494];
  assign o[494] = scan_lo[494] & N17;
  assign N17 = ~scan_lo[493];
  assign o[493] = scan_lo[493] & N18;
  assign N18 = ~scan_lo[492];
  assign o[492] = scan_lo[492] & N19;
  assign N19 = ~scan_lo[491];
  assign o[491] = scan_lo[491] & N20;
  assign N20 = ~scan_lo[490];
  assign o[490] = scan_lo[490] & N21;
  assign N21 = ~scan_lo[489];
  assign o[489] = scan_lo[489] & N22;
  assign N22 = ~scan_lo[488];
  assign o[488] = scan_lo[488] & N23;
  assign N23 = ~scan_lo[487];
  assign o[487] = scan_lo[487] & N24;
  assign N24 = ~scan_lo[486];
  assign o[486] = scan_lo[486] & N25;
  assign N25 = ~scan_lo[485];
  assign o[485] = scan_lo[485] & N26;
  assign N26 = ~scan_lo[484];
  assign o[484] = scan_lo[484] & N27;
  assign N27 = ~scan_lo[483];
  assign o[483] = scan_lo[483] & N28;
  assign N28 = ~scan_lo[482];
  assign o[482] = scan_lo[482] & N29;
  assign N29 = ~scan_lo[481];
  assign o[481] = scan_lo[481] & N30;
  assign N30 = ~scan_lo[480];
  assign o[480] = scan_lo[480] & N31;
  assign N31 = ~scan_lo[479];
  assign o[479] = scan_lo[479] & N32;
  assign N32 = ~scan_lo[478];
  assign o[478] = scan_lo[478] & N33;
  assign N33 = ~scan_lo[477];
  assign o[477] = scan_lo[477] & N34;
  assign N34 = ~scan_lo[476];
  assign o[476] = scan_lo[476] & N35;
  assign N35 = ~scan_lo[475];
  assign o[475] = scan_lo[475] & N36;
  assign N36 = ~scan_lo[474];
  assign o[474] = scan_lo[474] & N37;
  assign N37 = ~scan_lo[473];
  assign o[473] = scan_lo[473] & N38;
  assign N38 = ~scan_lo[472];
  assign o[472] = scan_lo[472] & N39;
  assign N39 = ~scan_lo[471];
  assign o[471] = scan_lo[471] & N40;
  assign N40 = ~scan_lo[470];
  assign o[470] = scan_lo[470] & N41;
  assign N41 = ~scan_lo[469];
  assign o[469] = scan_lo[469] & N42;
  assign N42 = ~scan_lo[468];
  assign o[468] = scan_lo[468] & N43;
  assign N43 = ~scan_lo[467];
  assign o[467] = scan_lo[467] & N44;
  assign N44 = ~scan_lo[466];
  assign o[466] = scan_lo[466] & N45;
  assign N45 = ~scan_lo[465];
  assign o[465] = scan_lo[465] & N46;
  assign N46 = ~scan_lo[464];
  assign o[464] = scan_lo[464] & N47;
  assign N47 = ~scan_lo[463];
  assign o[463] = scan_lo[463] & N48;
  assign N48 = ~scan_lo[462];
  assign o[462] = scan_lo[462] & N49;
  assign N49 = ~scan_lo[461];
  assign o[461] = scan_lo[461] & N50;
  assign N50 = ~scan_lo[460];
  assign o[460] = scan_lo[460] & N51;
  assign N51 = ~scan_lo[459];
  assign o[459] = scan_lo[459] & N52;
  assign N52 = ~scan_lo[458];
  assign o[458] = scan_lo[458] & N53;
  assign N53 = ~scan_lo[457];
  assign o[457] = scan_lo[457] & N54;
  assign N54 = ~scan_lo[456];
  assign o[456] = scan_lo[456] & N55;
  assign N55 = ~scan_lo[455];
  assign o[455] = scan_lo[455] & N56;
  assign N56 = ~scan_lo[454];
  assign o[454] = scan_lo[454] & N57;
  assign N57 = ~scan_lo[453];
  assign o[453] = scan_lo[453] & N58;
  assign N58 = ~scan_lo[452];
  assign o[452] = scan_lo[452] & N59;
  assign N59 = ~scan_lo[451];
  assign o[451] = scan_lo[451] & N60;
  assign N60 = ~scan_lo[450];
  assign o[450] = scan_lo[450] & N61;
  assign N61 = ~scan_lo[449];
  assign o[449] = scan_lo[449] & N62;
  assign N62 = ~scan_lo[448];
  assign o[448] = scan_lo[448] & N63;
  assign N63 = ~scan_lo[447];
  assign o[447] = scan_lo[447] & N64;
  assign N64 = ~scan_lo[446];
  assign o[446] = scan_lo[446] & N65;
  assign N65 = ~scan_lo[445];
  assign o[445] = scan_lo[445] & N66;
  assign N66 = ~scan_lo[444];
  assign o[444] = scan_lo[444] & N67;
  assign N67 = ~scan_lo[443];
  assign o[443] = scan_lo[443] & N68;
  assign N68 = ~scan_lo[442];
  assign o[442] = scan_lo[442] & N69;
  assign N69 = ~scan_lo[441];
  assign o[441] = scan_lo[441] & N70;
  assign N70 = ~scan_lo[440];
  assign o[440] = scan_lo[440] & N71;
  assign N71 = ~scan_lo[439];
  assign o[439] = scan_lo[439] & N72;
  assign N72 = ~scan_lo[438];
  assign o[438] = scan_lo[438] & N73;
  assign N73 = ~scan_lo[437];
  assign o[437] = scan_lo[437] & N74;
  assign N74 = ~scan_lo[436];
  assign o[436] = scan_lo[436] & N75;
  assign N75 = ~scan_lo[435];
  assign o[435] = scan_lo[435] & N76;
  assign N76 = ~scan_lo[434];
  assign o[434] = scan_lo[434] & N77;
  assign N77 = ~scan_lo[433];
  assign o[433] = scan_lo[433] & N78;
  assign N78 = ~scan_lo[432];
  assign o[432] = scan_lo[432] & N79;
  assign N79 = ~scan_lo[431];
  assign o[431] = scan_lo[431] & N80;
  assign N80 = ~scan_lo[430];
  assign o[430] = scan_lo[430] & N81;
  assign N81 = ~scan_lo[429];
  assign o[429] = scan_lo[429] & N82;
  assign N82 = ~scan_lo[428];
  assign o[428] = scan_lo[428] & N83;
  assign N83 = ~scan_lo[427];
  assign o[427] = scan_lo[427] & N84;
  assign N84 = ~scan_lo[426];
  assign o[426] = scan_lo[426] & N85;
  assign N85 = ~scan_lo[425];
  assign o[425] = scan_lo[425] & N86;
  assign N86 = ~scan_lo[424];
  assign o[424] = scan_lo[424] & N87;
  assign N87 = ~scan_lo[423];
  assign o[423] = scan_lo[423] & N88;
  assign N88 = ~scan_lo[422];
  assign o[422] = scan_lo[422] & N89;
  assign N89 = ~scan_lo[421];
  assign o[421] = scan_lo[421] & N90;
  assign N90 = ~scan_lo[420];
  assign o[420] = scan_lo[420] & N91;
  assign N91 = ~scan_lo[419];
  assign o[419] = scan_lo[419] & N92;
  assign N92 = ~scan_lo[418];
  assign o[418] = scan_lo[418] & N93;
  assign N93 = ~scan_lo[417];
  assign o[417] = scan_lo[417] & N94;
  assign N94 = ~scan_lo[416];
  assign o[416] = scan_lo[416] & N95;
  assign N95 = ~scan_lo[415];
  assign o[415] = scan_lo[415] & N96;
  assign N96 = ~scan_lo[414];
  assign o[414] = scan_lo[414] & N97;
  assign N97 = ~scan_lo[413];
  assign o[413] = scan_lo[413] & N98;
  assign N98 = ~scan_lo[412];
  assign o[412] = scan_lo[412] & N99;
  assign N99 = ~scan_lo[411];
  assign o[411] = scan_lo[411] & N100;
  assign N100 = ~scan_lo[410];
  assign o[410] = scan_lo[410] & N101;
  assign N101 = ~scan_lo[409];
  assign o[409] = scan_lo[409] & N102;
  assign N102 = ~scan_lo[408];
  assign o[408] = scan_lo[408] & N103;
  assign N103 = ~scan_lo[407];
  assign o[407] = scan_lo[407] & N104;
  assign N104 = ~scan_lo[406];
  assign o[406] = scan_lo[406] & N105;
  assign N105 = ~scan_lo[405];
  assign o[405] = scan_lo[405] & N106;
  assign N106 = ~scan_lo[404];
  assign o[404] = scan_lo[404] & N107;
  assign N107 = ~scan_lo[403];
  assign o[403] = scan_lo[403] & N108;
  assign N108 = ~scan_lo[402];
  assign o[402] = scan_lo[402] & N109;
  assign N109 = ~scan_lo[401];
  assign o[401] = scan_lo[401] & N110;
  assign N110 = ~scan_lo[400];
  assign o[400] = scan_lo[400] & N111;
  assign N111 = ~scan_lo[399];
  assign o[399] = scan_lo[399] & N112;
  assign N112 = ~scan_lo[398];
  assign o[398] = scan_lo[398] & N113;
  assign N113 = ~scan_lo[397];
  assign o[397] = scan_lo[397] & N114;
  assign N114 = ~scan_lo[396];
  assign o[396] = scan_lo[396] & N115;
  assign N115 = ~scan_lo[395];
  assign o[395] = scan_lo[395] & N116;
  assign N116 = ~scan_lo[394];
  assign o[394] = scan_lo[394] & N117;
  assign N117 = ~scan_lo[393];
  assign o[393] = scan_lo[393] & N118;
  assign N118 = ~scan_lo[392];
  assign o[392] = scan_lo[392] & N119;
  assign N119 = ~scan_lo[391];
  assign o[391] = scan_lo[391] & N120;
  assign N120 = ~scan_lo[390];
  assign o[390] = scan_lo[390] & N121;
  assign N121 = ~scan_lo[389];
  assign o[389] = scan_lo[389] & N122;
  assign N122 = ~scan_lo[388];
  assign o[388] = scan_lo[388] & N123;
  assign N123 = ~scan_lo[387];
  assign o[387] = scan_lo[387] & N124;
  assign N124 = ~scan_lo[386];
  assign o[386] = scan_lo[386] & N125;
  assign N125 = ~scan_lo[385];
  assign o[385] = scan_lo[385] & N126;
  assign N126 = ~scan_lo[384];
  assign o[384] = scan_lo[384] & N127;
  assign N127 = ~scan_lo[383];
  assign o[383] = scan_lo[383] & N128;
  assign N128 = ~scan_lo[382];
  assign o[382] = scan_lo[382] & N129;
  assign N129 = ~scan_lo[381];
  assign o[381] = scan_lo[381] & N130;
  assign N130 = ~scan_lo[380];
  assign o[380] = scan_lo[380] & N131;
  assign N131 = ~scan_lo[379];
  assign o[379] = scan_lo[379] & N132;
  assign N132 = ~scan_lo[378];
  assign o[378] = scan_lo[378] & N133;
  assign N133 = ~scan_lo[377];
  assign o[377] = scan_lo[377] & N134;
  assign N134 = ~scan_lo[376];
  assign o[376] = scan_lo[376] & N135;
  assign N135 = ~scan_lo[375];
  assign o[375] = scan_lo[375] & N136;
  assign N136 = ~scan_lo[374];
  assign o[374] = scan_lo[374] & N137;
  assign N137 = ~scan_lo[373];
  assign o[373] = scan_lo[373] & N138;
  assign N138 = ~scan_lo[372];
  assign o[372] = scan_lo[372] & N139;
  assign N139 = ~scan_lo[371];
  assign o[371] = scan_lo[371] & N140;
  assign N140 = ~scan_lo[370];
  assign o[370] = scan_lo[370] & N141;
  assign N141 = ~scan_lo[369];
  assign o[369] = scan_lo[369] & N142;
  assign N142 = ~scan_lo[368];
  assign o[368] = scan_lo[368] & N143;
  assign N143 = ~scan_lo[367];
  assign o[367] = scan_lo[367] & N144;
  assign N144 = ~scan_lo[366];
  assign o[366] = scan_lo[366] & N145;
  assign N145 = ~scan_lo[365];
  assign o[365] = scan_lo[365] & N146;
  assign N146 = ~scan_lo[364];
  assign o[364] = scan_lo[364] & N147;
  assign N147 = ~scan_lo[363];
  assign o[363] = scan_lo[363] & N148;
  assign N148 = ~scan_lo[362];
  assign o[362] = scan_lo[362] & N149;
  assign N149 = ~scan_lo[361];
  assign o[361] = scan_lo[361] & N150;
  assign N150 = ~scan_lo[360];
  assign o[360] = scan_lo[360] & N151;
  assign N151 = ~scan_lo[359];
  assign o[359] = scan_lo[359] & N152;
  assign N152 = ~scan_lo[358];
  assign o[358] = scan_lo[358] & N153;
  assign N153 = ~scan_lo[357];
  assign o[357] = scan_lo[357] & N154;
  assign N154 = ~scan_lo[356];
  assign o[356] = scan_lo[356] & N155;
  assign N155 = ~scan_lo[355];
  assign o[355] = scan_lo[355] & N156;
  assign N156 = ~scan_lo[354];
  assign o[354] = scan_lo[354] & N157;
  assign N157 = ~scan_lo[353];
  assign o[353] = scan_lo[353] & N158;
  assign N158 = ~scan_lo[352];
  assign o[352] = scan_lo[352] & N159;
  assign N159 = ~scan_lo[351];
  assign o[351] = scan_lo[351] & N160;
  assign N160 = ~scan_lo[350];
  assign o[350] = scan_lo[350] & N161;
  assign N161 = ~scan_lo[349];
  assign o[349] = scan_lo[349] & N162;
  assign N162 = ~scan_lo[348];
  assign o[348] = scan_lo[348] & N163;
  assign N163 = ~scan_lo[347];
  assign o[347] = scan_lo[347] & N164;
  assign N164 = ~scan_lo[346];
  assign o[346] = scan_lo[346] & N165;
  assign N165 = ~scan_lo[345];
  assign o[345] = scan_lo[345] & N166;
  assign N166 = ~scan_lo[344];
  assign o[344] = scan_lo[344] & N167;
  assign N167 = ~scan_lo[343];
  assign o[343] = scan_lo[343] & N168;
  assign N168 = ~scan_lo[342];
  assign o[342] = scan_lo[342] & N169;
  assign N169 = ~scan_lo[341];
  assign o[341] = scan_lo[341] & N170;
  assign N170 = ~scan_lo[340];
  assign o[340] = scan_lo[340] & N171;
  assign N171 = ~scan_lo[339];
  assign o[339] = scan_lo[339] & N172;
  assign N172 = ~scan_lo[338];
  assign o[338] = scan_lo[338] & N173;
  assign N173 = ~scan_lo[337];
  assign o[337] = scan_lo[337] & N174;
  assign N174 = ~scan_lo[336];
  assign o[336] = scan_lo[336] & N175;
  assign N175 = ~scan_lo[335];
  assign o[335] = scan_lo[335] & N176;
  assign N176 = ~scan_lo[334];
  assign o[334] = scan_lo[334] & N177;
  assign N177 = ~scan_lo[333];
  assign o[333] = scan_lo[333] & N178;
  assign N178 = ~scan_lo[332];
  assign o[332] = scan_lo[332] & N179;
  assign N179 = ~scan_lo[331];
  assign o[331] = scan_lo[331] & N180;
  assign N180 = ~scan_lo[330];
  assign o[330] = scan_lo[330] & N181;
  assign N181 = ~scan_lo[329];
  assign o[329] = scan_lo[329] & N182;
  assign N182 = ~scan_lo[328];
  assign o[328] = scan_lo[328] & N183;
  assign N183 = ~scan_lo[327];
  assign o[327] = scan_lo[327] & N184;
  assign N184 = ~scan_lo[326];
  assign o[326] = scan_lo[326] & N185;
  assign N185 = ~scan_lo[325];
  assign o[325] = scan_lo[325] & N186;
  assign N186 = ~scan_lo[324];
  assign o[324] = scan_lo[324] & N187;
  assign N187 = ~scan_lo[323];
  assign o[323] = scan_lo[323] & N188;
  assign N188 = ~scan_lo[322];
  assign o[322] = scan_lo[322] & N189;
  assign N189 = ~scan_lo[321];
  assign o[321] = scan_lo[321] & N190;
  assign N190 = ~scan_lo[320];
  assign o[320] = scan_lo[320] & N191;
  assign N191 = ~scan_lo[319];
  assign o[319] = scan_lo[319] & N192;
  assign N192 = ~scan_lo[318];
  assign o[318] = scan_lo[318] & N193;
  assign N193 = ~scan_lo[317];
  assign o[317] = scan_lo[317] & N194;
  assign N194 = ~scan_lo[316];
  assign o[316] = scan_lo[316] & N195;
  assign N195 = ~scan_lo[315];
  assign o[315] = scan_lo[315] & N196;
  assign N196 = ~scan_lo[314];
  assign o[314] = scan_lo[314] & N197;
  assign N197 = ~scan_lo[313];
  assign o[313] = scan_lo[313] & N198;
  assign N198 = ~scan_lo[312];
  assign o[312] = scan_lo[312] & N199;
  assign N199 = ~scan_lo[311];
  assign o[311] = scan_lo[311] & N200;
  assign N200 = ~scan_lo[310];
  assign o[310] = scan_lo[310] & N201;
  assign N201 = ~scan_lo[309];
  assign o[309] = scan_lo[309] & N202;
  assign N202 = ~scan_lo[308];
  assign o[308] = scan_lo[308] & N203;
  assign N203 = ~scan_lo[307];
  assign o[307] = scan_lo[307] & N204;
  assign N204 = ~scan_lo[306];
  assign o[306] = scan_lo[306] & N205;
  assign N205 = ~scan_lo[305];
  assign o[305] = scan_lo[305] & N206;
  assign N206 = ~scan_lo[304];
  assign o[304] = scan_lo[304] & N207;
  assign N207 = ~scan_lo[303];
  assign o[303] = scan_lo[303] & N208;
  assign N208 = ~scan_lo[302];
  assign o[302] = scan_lo[302] & N209;
  assign N209 = ~scan_lo[301];
  assign o[301] = scan_lo[301] & N210;
  assign N210 = ~scan_lo[300];
  assign o[300] = scan_lo[300] & N211;
  assign N211 = ~scan_lo[299];
  assign o[299] = scan_lo[299] & N212;
  assign N212 = ~scan_lo[298];
  assign o[298] = scan_lo[298] & N213;
  assign N213 = ~scan_lo[297];
  assign o[297] = scan_lo[297] & N214;
  assign N214 = ~scan_lo[296];
  assign o[296] = scan_lo[296] & N215;
  assign N215 = ~scan_lo[295];
  assign o[295] = scan_lo[295] & N216;
  assign N216 = ~scan_lo[294];
  assign o[294] = scan_lo[294] & N217;
  assign N217 = ~scan_lo[293];
  assign o[293] = scan_lo[293] & N218;
  assign N218 = ~scan_lo[292];
  assign o[292] = scan_lo[292] & N219;
  assign N219 = ~scan_lo[291];
  assign o[291] = scan_lo[291] & N220;
  assign N220 = ~scan_lo[290];
  assign o[290] = scan_lo[290] & N221;
  assign N221 = ~scan_lo[289];
  assign o[289] = scan_lo[289] & N222;
  assign N222 = ~scan_lo[288];
  assign o[288] = scan_lo[288] & N223;
  assign N223 = ~scan_lo[287];
  assign o[287] = scan_lo[287] & N224;
  assign N224 = ~scan_lo[286];
  assign o[286] = scan_lo[286] & N225;
  assign N225 = ~scan_lo[285];
  assign o[285] = scan_lo[285] & N226;
  assign N226 = ~scan_lo[284];
  assign o[284] = scan_lo[284] & N227;
  assign N227 = ~scan_lo[283];
  assign o[283] = scan_lo[283] & N228;
  assign N228 = ~scan_lo[282];
  assign o[282] = scan_lo[282] & N229;
  assign N229 = ~scan_lo[281];
  assign o[281] = scan_lo[281] & N230;
  assign N230 = ~scan_lo[280];
  assign o[280] = scan_lo[280] & N231;
  assign N231 = ~scan_lo[279];
  assign o[279] = scan_lo[279] & N232;
  assign N232 = ~scan_lo[278];
  assign o[278] = scan_lo[278] & N233;
  assign N233 = ~scan_lo[277];
  assign o[277] = scan_lo[277] & N234;
  assign N234 = ~scan_lo[276];
  assign o[276] = scan_lo[276] & N235;
  assign N235 = ~scan_lo[275];
  assign o[275] = scan_lo[275] & N236;
  assign N236 = ~scan_lo[274];
  assign o[274] = scan_lo[274] & N237;
  assign N237 = ~scan_lo[273];
  assign o[273] = scan_lo[273] & N238;
  assign N238 = ~scan_lo[272];
  assign o[272] = scan_lo[272] & N239;
  assign N239 = ~scan_lo[271];
  assign o[271] = scan_lo[271] & N240;
  assign N240 = ~scan_lo[270];
  assign o[270] = scan_lo[270] & N241;
  assign N241 = ~scan_lo[269];
  assign o[269] = scan_lo[269] & N242;
  assign N242 = ~scan_lo[268];
  assign o[268] = scan_lo[268] & N243;
  assign N243 = ~scan_lo[267];
  assign o[267] = scan_lo[267] & N244;
  assign N244 = ~scan_lo[266];
  assign o[266] = scan_lo[266] & N245;
  assign N245 = ~scan_lo[265];
  assign o[265] = scan_lo[265] & N246;
  assign N246 = ~scan_lo[264];
  assign o[264] = scan_lo[264] & N247;
  assign N247 = ~scan_lo[263];
  assign o[263] = scan_lo[263] & N248;
  assign N248 = ~scan_lo[262];
  assign o[262] = scan_lo[262] & N249;
  assign N249 = ~scan_lo[261];
  assign o[261] = scan_lo[261] & N250;
  assign N250 = ~scan_lo[260];
  assign o[260] = scan_lo[260] & N251;
  assign N251 = ~scan_lo[259];
  assign o[259] = scan_lo[259] & N252;
  assign N252 = ~scan_lo[258];
  assign o[258] = scan_lo[258] & N253;
  assign N253 = ~scan_lo[257];
  assign o[257] = scan_lo[257] & N254;
  assign N254 = ~scan_lo[256];
  assign o[256] = scan_lo[256] & N255;
  assign N255 = ~scan_lo[255];
  assign o[255] = scan_lo[255] & N256;
  assign N256 = ~scan_lo[254];
  assign o[254] = scan_lo[254] & N257;
  assign N257 = ~scan_lo[253];
  assign o[253] = scan_lo[253] & N258;
  assign N258 = ~scan_lo[252];
  assign o[252] = scan_lo[252] & N259;
  assign N259 = ~scan_lo[251];
  assign o[251] = scan_lo[251] & N260;
  assign N260 = ~scan_lo[250];
  assign o[250] = scan_lo[250] & N261;
  assign N261 = ~scan_lo[249];
  assign o[249] = scan_lo[249] & N262;
  assign N262 = ~scan_lo[248];
  assign o[248] = scan_lo[248] & N263;
  assign N263 = ~scan_lo[247];
  assign o[247] = scan_lo[247] & N264;
  assign N264 = ~scan_lo[246];
  assign o[246] = scan_lo[246] & N265;
  assign N265 = ~scan_lo[245];
  assign o[245] = scan_lo[245] & N266;
  assign N266 = ~scan_lo[244];
  assign o[244] = scan_lo[244] & N267;
  assign N267 = ~scan_lo[243];
  assign o[243] = scan_lo[243] & N268;
  assign N268 = ~scan_lo[242];
  assign o[242] = scan_lo[242] & N269;
  assign N269 = ~scan_lo[241];
  assign o[241] = scan_lo[241] & N270;
  assign N270 = ~scan_lo[240];
  assign o[240] = scan_lo[240] & N271;
  assign N271 = ~scan_lo[239];
  assign o[239] = scan_lo[239] & N272;
  assign N272 = ~scan_lo[238];
  assign o[238] = scan_lo[238] & N273;
  assign N273 = ~scan_lo[237];
  assign o[237] = scan_lo[237] & N274;
  assign N274 = ~scan_lo[236];
  assign o[236] = scan_lo[236] & N275;
  assign N275 = ~scan_lo[235];
  assign o[235] = scan_lo[235] & N276;
  assign N276 = ~scan_lo[234];
  assign o[234] = scan_lo[234] & N277;
  assign N277 = ~scan_lo[233];
  assign o[233] = scan_lo[233] & N278;
  assign N278 = ~scan_lo[232];
  assign o[232] = scan_lo[232] & N279;
  assign N279 = ~scan_lo[231];
  assign o[231] = scan_lo[231] & N280;
  assign N280 = ~scan_lo[230];
  assign o[230] = scan_lo[230] & N281;
  assign N281 = ~scan_lo[229];
  assign o[229] = scan_lo[229] & N282;
  assign N282 = ~scan_lo[228];
  assign o[228] = scan_lo[228] & N283;
  assign N283 = ~scan_lo[227];
  assign o[227] = scan_lo[227] & N284;
  assign N284 = ~scan_lo[226];
  assign o[226] = scan_lo[226] & N285;
  assign N285 = ~scan_lo[225];
  assign o[225] = scan_lo[225] & N286;
  assign N286 = ~scan_lo[224];
  assign o[224] = scan_lo[224] & N287;
  assign N287 = ~scan_lo[223];
  assign o[223] = scan_lo[223] & N288;
  assign N288 = ~scan_lo[222];
  assign o[222] = scan_lo[222] & N289;
  assign N289 = ~scan_lo[221];
  assign o[221] = scan_lo[221] & N290;
  assign N290 = ~scan_lo[220];
  assign o[220] = scan_lo[220] & N291;
  assign N291 = ~scan_lo[219];
  assign o[219] = scan_lo[219] & N292;
  assign N292 = ~scan_lo[218];
  assign o[218] = scan_lo[218] & N293;
  assign N293 = ~scan_lo[217];
  assign o[217] = scan_lo[217] & N294;
  assign N294 = ~scan_lo[216];
  assign o[216] = scan_lo[216] & N295;
  assign N295 = ~scan_lo[215];
  assign o[215] = scan_lo[215] & N296;
  assign N296 = ~scan_lo[214];
  assign o[214] = scan_lo[214] & N297;
  assign N297 = ~scan_lo[213];
  assign o[213] = scan_lo[213] & N298;
  assign N298 = ~scan_lo[212];
  assign o[212] = scan_lo[212] & N299;
  assign N299 = ~scan_lo[211];
  assign o[211] = scan_lo[211] & N300;
  assign N300 = ~scan_lo[210];
  assign o[210] = scan_lo[210] & N301;
  assign N301 = ~scan_lo[209];
  assign o[209] = scan_lo[209] & N302;
  assign N302 = ~scan_lo[208];
  assign o[208] = scan_lo[208] & N303;
  assign N303 = ~scan_lo[207];
  assign o[207] = scan_lo[207] & N304;
  assign N304 = ~scan_lo[206];
  assign o[206] = scan_lo[206] & N305;
  assign N305 = ~scan_lo[205];
  assign o[205] = scan_lo[205] & N306;
  assign N306 = ~scan_lo[204];
  assign o[204] = scan_lo[204] & N307;
  assign N307 = ~scan_lo[203];
  assign o[203] = scan_lo[203] & N308;
  assign N308 = ~scan_lo[202];
  assign o[202] = scan_lo[202] & N309;
  assign N309 = ~scan_lo[201];
  assign o[201] = scan_lo[201] & N310;
  assign N310 = ~scan_lo[200];
  assign o[200] = scan_lo[200] & N311;
  assign N311 = ~scan_lo[199];
  assign o[199] = scan_lo[199] & N312;
  assign N312 = ~scan_lo[198];
  assign o[198] = scan_lo[198] & N313;
  assign N313 = ~scan_lo[197];
  assign o[197] = scan_lo[197] & N314;
  assign N314 = ~scan_lo[196];
  assign o[196] = scan_lo[196] & N315;
  assign N315 = ~scan_lo[195];
  assign o[195] = scan_lo[195] & N316;
  assign N316 = ~scan_lo[194];
  assign o[194] = scan_lo[194] & N317;
  assign N317 = ~scan_lo[193];
  assign o[193] = scan_lo[193] & N318;
  assign N318 = ~scan_lo[192];
  assign o[192] = scan_lo[192] & N319;
  assign N319 = ~scan_lo[191];
  assign o[191] = scan_lo[191] & N320;
  assign N320 = ~scan_lo[190];
  assign o[190] = scan_lo[190] & N321;
  assign N321 = ~scan_lo[189];
  assign o[189] = scan_lo[189] & N322;
  assign N322 = ~scan_lo[188];
  assign o[188] = scan_lo[188] & N323;
  assign N323 = ~scan_lo[187];
  assign o[187] = scan_lo[187] & N324;
  assign N324 = ~scan_lo[186];
  assign o[186] = scan_lo[186] & N325;
  assign N325 = ~scan_lo[185];
  assign o[185] = scan_lo[185] & N326;
  assign N326 = ~scan_lo[184];
  assign o[184] = scan_lo[184] & N327;
  assign N327 = ~scan_lo[183];
  assign o[183] = scan_lo[183] & N328;
  assign N328 = ~scan_lo[182];
  assign o[182] = scan_lo[182] & N329;
  assign N329 = ~scan_lo[181];
  assign o[181] = scan_lo[181] & N330;
  assign N330 = ~scan_lo[180];
  assign o[180] = scan_lo[180] & N331;
  assign N331 = ~scan_lo[179];
  assign o[179] = scan_lo[179] & N332;
  assign N332 = ~scan_lo[178];
  assign o[178] = scan_lo[178] & N333;
  assign N333 = ~scan_lo[177];
  assign o[177] = scan_lo[177] & N334;
  assign N334 = ~scan_lo[176];
  assign o[176] = scan_lo[176] & N335;
  assign N335 = ~scan_lo[175];
  assign o[175] = scan_lo[175] & N336;
  assign N336 = ~scan_lo[174];
  assign o[174] = scan_lo[174] & N337;
  assign N337 = ~scan_lo[173];
  assign o[173] = scan_lo[173] & N338;
  assign N338 = ~scan_lo[172];
  assign o[172] = scan_lo[172] & N339;
  assign N339 = ~scan_lo[171];
  assign o[171] = scan_lo[171] & N340;
  assign N340 = ~scan_lo[170];
  assign o[170] = scan_lo[170] & N341;
  assign N341 = ~scan_lo[169];
  assign o[169] = scan_lo[169] & N342;
  assign N342 = ~scan_lo[168];
  assign o[168] = scan_lo[168] & N343;
  assign N343 = ~scan_lo[167];
  assign o[167] = scan_lo[167] & N344;
  assign N344 = ~scan_lo[166];
  assign o[166] = scan_lo[166] & N345;
  assign N345 = ~scan_lo[165];
  assign o[165] = scan_lo[165] & N346;
  assign N346 = ~scan_lo[164];
  assign o[164] = scan_lo[164] & N347;
  assign N347 = ~scan_lo[163];
  assign o[163] = scan_lo[163] & N348;
  assign N348 = ~scan_lo[162];
  assign o[162] = scan_lo[162] & N349;
  assign N349 = ~scan_lo[161];
  assign o[161] = scan_lo[161] & N350;
  assign N350 = ~scan_lo[160];
  assign o[160] = scan_lo[160] & N351;
  assign N351 = ~scan_lo[159];
  assign o[159] = scan_lo[159] & N352;
  assign N352 = ~scan_lo[158];
  assign o[158] = scan_lo[158] & N353;
  assign N353 = ~scan_lo[157];
  assign o[157] = scan_lo[157] & N354;
  assign N354 = ~scan_lo[156];
  assign o[156] = scan_lo[156] & N355;
  assign N355 = ~scan_lo[155];
  assign o[155] = scan_lo[155] & N356;
  assign N356 = ~scan_lo[154];
  assign o[154] = scan_lo[154] & N357;
  assign N357 = ~scan_lo[153];
  assign o[153] = scan_lo[153] & N358;
  assign N358 = ~scan_lo[152];
  assign o[152] = scan_lo[152] & N359;
  assign N359 = ~scan_lo[151];
  assign o[151] = scan_lo[151] & N360;
  assign N360 = ~scan_lo[150];
  assign o[150] = scan_lo[150] & N361;
  assign N361 = ~scan_lo[149];
  assign o[149] = scan_lo[149] & N362;
  assign N362 = ~scan_lo[148];
  assign o[148] = scan_lo[148] & N363;
  assign N363 = ~scan_lo[147];
  assign o[147] = scan_lo[147] & N364;
  assign N364 = ~scan_lo[146];
  assign o[146] = scan_lo[146] & N365;
  assign N365 = ~scan_lo[145];
  assign o[145] = scan_lo[145] & N366;
  assign N366 = ~scan_lo[144];
  assign o[144] = scan_lo[144] & N367;
  assign N367 = ~scan_lo[143];
  assign o[143] = scan_lo[143] & N368;
  assign N368 = ~scan_lo[142];
  assign o[142] = scan_lo[142] & N369;
  assign N369 = ~scan_lo[141];
  assign o[141] = scan_lo[141] & N370;
  assign N370 = ~scan_lo[140];
  assign o[140] = scan_lo[140] & N371;
  assign N371 = ~scan_lo[139];
  assign o[139] = scan_lo[139] & N372;
  assign N372 = ~scan_lo[138];
  assign o[138] = scan_lo[138] & N373;
  assign N373 = ~scan_lo[137];
  assign o[137] = scan_lo[137] & N374;
  assign N374 = ~scan_lo[136];
  assign o[136] = scan_lo[136] & N375;
  assign N375 = ~scan_lo[135];
  assign o[135] = scan_lo[135] & N376;
  assign N376 = ~scan_lo[134];
  assign o[134] = scan_lo[134] & N377;
  assign N377 = ~scan_lo[133];
  assign o[133] = scan_lo[133] & N378;
  assign N378 = ~scan_lo[132];
  assign o[132] = scan_lo[132] & N379;
  assign N379 = ~scan_lo[131];
  assign o[131] = scan_lo[131] & N380;
  assign N380 = ~scan_lo[130];
  assign o[130] = scan_lo[130] & N381;
  assign N381 = ~scan_lo[129];
  assign o[129] = scan_lo[129] & N382;
  assign N382 = ~scan_lo[128];
  assign o[128] = scan_lo[128] & N383;
  assign N383 = ~scan_lo[127];
  assign o[127] = scan_lo[127] & N384;
  assign N384 = ~scan_lo[126];
  assign o[126] = scan_lo[126] & N385;
  assign N385 = ~scan_lo[125];
  assign o[125] = scan_lo[125] & N386;
  assign N386 = ~scan_lo[124];
  assign o[124] = scan_lo[124] & N387;
  assign N387 = ~scan_lo[123];
  assign o[123] = scan_lo[123] & N388;
  assign N388 = ~scan_lo[122];
  assign o[122] = scan_lo[122] & N389;
  assign N389 = ~scan_lo[121];
  assign o[121] = scan_lo[121] & N390;
  assign N390 = ~scan_lo[120];
  assign o[120] = scan_lo[120] & N391;
  assign N391 = ~scan_lo[119];
  assign o[119] = scan_lo[119] & N392;
  assign N392 = ~scan_lo[118];
  assign o[118] = scan_lo[118] & N393;
  assign N393 = ~scan_lo[117];
  assign o[117] = scan_lo[117] & N394;
  assign N394 = ~scan_lo[116];
  assign o[116] = scan_lo[116] & N395;
  assign N395 = ~scan_lo[115];
  assign o[115] = scan_lo[115] & N396;
  assign N396 = ~scan_lo[114];
  assign o[114] = scan_lo[114] & N397;
  assign N397 = ~scan_lo[113];
  assign o[113] = scan_lo[113] & N398;
  assign N398 = ~scan_lo[112];
  assign o[112] = scan_lo[112] & N399;
  assign N399 = ~scan_lo[111];
  assign o[111] = scan_lo[111] & N400;
  assign N400 = ~scan_lo[110];
  assign o[110] = scan_lo[110] & N401;
  assign N401 = ~scan_lo[109];
  assign o[109] = scan_lo[109] & N402;
  assign N402 = ~scan_lo[108];
  assign o[108] = scan_lo[108] & N403;
  assign N403 = ~scan_lo[107];
  assign o[107] = scan_lo[107] & N404;
  assign N404 = ~scan_lo[106];
  assign o[106] = scan_lo[106] & N405;
  assign N405 = ~scan_lo[105];
  assign o[105] = scan_lo[105] & N406;
  assign N406 = ~scan_lo[104];
  assign o[104] = scan_lo[104] & N407;
  assign N407 = ~scan_lo[103];
  assign o[103] = scan_lo[103] & N408;
  assign N408 = ~scan_lo[102];
  assign o[102] = scan_lo[102] & N409;
  assign N409 = ~scan_lo[101];
  assign o[101] = scan_lo[101] & N410;
  assign N410 = ~scan_lo[100];
  assign o[100] = scan_lo[100] & N411;
  assign N411 = ~scan_lo[99];
  assign o[99] = scan_lo[99] & N412;
  assign N412 = ~scan_lo[98];
  assign o[98] = scan_lo[98] & N413;
  assign N413 = ~scan_lo[97];
  assign o[97] = scan_lo[97] & N414;
  assign N414 = ~scan_lo[96];
  assign o[96] = scan_lo[96] & N415;
  assign N415 = ~scan_lo[95];
  assign o[95] = scan_lo[95] & N416;
  assign N416 = ~scan_lo[94];
  assign o[94] = scan_lo[94] & N417;
  assign N417 = ~scan_lo[93];
  assign o[93] = scan_lo[93] & N418;
  assign N418 = ~scan_lo[92];
  assign o[92] = scan_lo[92] & N419;
  assign N419 = ~scan_lo[91];
  assign o[91] = scan_lo[91] & N420;
  assign N420 = ~scan_lo[90];
  assign o[90] = scan_lo[90] & N421;
  assign N421 = ~scan_lo[89];
  assign o[89] = scan_lo[89] & N422;
  assign N422 = ~scan_lo[88];
  assign o[88] = scan_lo[88] & N423;
  assign N423 = ~scan_lo[87];
  assign o[87] = scan_lo[87] & N424;
  assign N424 = ~scan_lo[86];
  assign o[86] = scan_lo[86] & N425;
  assign N425 = ~scan_lo[85];
  assign o[85] = scan_lo[85] & N426;
  assign N426 = ~scan_lo[84];
  assign o[84] = scan_lo[84] & N427;
  assign N427 = ~scan_lo[83];
  assign o[83] = scan_lo[83] & N428;
  assign N428 = ~scan_lo[82];
  assign o[82] = scan_lo[82] & N429;
  assign N429 = ~scan_lo[81];
  assign o[81] = scan_lo[81] & N430;
  assign N430 = ~scan_lo[80];
  assign o[80] = scan_lo[80] & N431;
  assign N431 = ~scan_lo[79];
  assign o[79] = scan_lo[79] & N432;
  assign N432 = ~scan_lo[78];
  assign o[78] = scan_lo[78] & N433;
  assign N433 = ~scan_lo[77];
  assign o[77] = scan_lo[77] & N434;
  assign N434 = ~scan_lo[76];
  assign o[76] = scan_lo[76] & N435;
  assign N435 = ~scan_lo[75];
  assign o[75] = scan_lo[75] & N436;
  assign N436 = ~scan_lo[74];
  assign o[74] = scan_lo[74] & N437;
  assign N437 = ~scan_lo[73];
  assign o[73] = scan_lo[73] & N438;
  assign N438 = ~scan_lo[72];
  assign o[72] = scan_lo[72] & N439;
  assign N439 = ~scan_lo[71];
  assign o[71] = scan_lo[71] & N440;
  assign N440 = ~scan_lo[70];
  assign o[70] = scan_lo[70] & N441;
  assign N441 = ~scan_lo[69];
  assign o[69] = scan_lo[69] & N442;
  assign N442 = ~scan_lo[68];
  assign o[68] = scan_lo[68] & N443;
  assign N443 = ~scan_lo[67];
  assign o[67] = scan_lo[67] & N444;
  assign N444 = ~scan_lo[66];
  assign o[66] = scan_lo[66] & N445;
  assign N445 = ~scan_lo[65];
  assign o[65] = scan_lo[65] & N446;
  assign N446 = ~scan_lo[64];
  assign o[64] = scan_lo[64] & N447;
  assign N447 = ~scan_lo[63];
  assign o[63] = scan_lo[63] & N448;
  assign N448 = ~scan_lo[62];
  assign o[62] = scan_lo[62] & N449;
  assign N449 = ~scan_lo[61];
  assign o[61] = scan_lo[61] & N450;
  assign N450 = ~scan_lo[60];
  assign o[60] = scan_lo[60] & N451;
  assign N451 = ~scan_lo[59];
  assign o[59] = scan_lo[59] & N452;
  assign N452 = ~scan_lo[58];
  assign o[58] = scan_lo[58] & N453;
  assign N453 = ~scan_lo[57];
  assign o[57] = scan_lo[57] & N454;
  assign N454 = ~scan_lo[56];
  assign o[56] = scan_lo[56] & N455;
  assign N455 = ~scan_lo[55];
  assign o[55] = scan_lo[55] & N456;
  assign N456 = ~scan_lo[54];
  assign o[54] = scan_lo[54] & N457;
  assign N457 = ~scan_lo[53];
  assign o[53] = scan_lo[53] & N458;
  assign N458 = ~scan_lo[52];
  assign o[52] = scan_lo[52] & N459;
  assign N459 = ~scan_lo[51];
  assign o[51] = scan_lo[51] & N460;
  assign N460 = ~scan_lo[50];
  assign o[50] = scan_lo[50] & N461;
  assign N461 = ~scan_lo[49];
  assign o[49] = scan_lo[49] & N462;
  assign N462 = ~scan_lo[48];
  assign o[48] = scan_lo[48] & N463;
  assign N463 = ~scan_lo[47];
  assign o[47] = scan_lo[47] & N464;
  assign N464 = ~scan_lo[46];
  assign o[46] = scan_lo[46] & N465;
  assign N465 = ~scan_lo[45];
  assign o[45] = scan_lo[45] & N466;
  assign N466 = ~scan_lo[44];
  assign o[44] = scan_lo[44] & N467;
  assign N467 = ~scan_lo[43];
  assign o[43] = scan_lo[43] & N468;
  assign N468 = ~scan_lo[42];
  assign o[42] = scan_lo[42] & N469;
  assign N469 = ~scan_lo[41];
  assign o[41] = scan_lo[41] & N470;
  assign N470 = ~scan_lo[40];
  assign o[40] = scan_lo[40] & N471;
  assign N471 = ~scan_lo[39];
  assign o[39] = scan_lo[39] & N472;
  assign N472 = ~scan_lo[38];
  assign o[38] = scan_lo[38] & N473;
  assign N473 = ~scan_lo[37];
  assign o[37] = scan_lo[37] & N474;
  assign N474 = ~scan_lo[36];
  assign o[36] = scan_lo[36] & N475;
  assign N475 = ~scan_lo[35];
  assign o[35] = scan_lo[35] & N476;
  assign N476 = ~scan_lo[34];
  assign o[34] = scan_lo[34] & N477;
  assign N477 = ~scan_lo[33];
  assign o[33] = scan_lo[33] & N478;
  assign N478 = ~scan_lo[32];
  assign o[32] = scan_lo[32] & N479;
  assign N479 = ~scan_lo[31];
  assign o[31] = scan_lo[31] & N480;
  assign N480 = ~scan_lo[30];
  assign o[30] = scan_lo[30] & N481;
  assign N481 = ~scan_lo[29];
  assign o[29] = scan_lo[29] & N482;
  assign N482 = ~scan_lo[28];
  assign o[28] = scan_lo[28] & N483;
  assign N483 = ~scan_lo[27];
  assign o[27] = scan_lo[27] & N484;
  assign N484 = ~scan_lo[26];
  assign o[26] = scan_lo[26] & N485;
  assign N485 = ~scan_lo[25];
  assign o[25] = scan_lo[25] & N486;
  assign N486 = ~scan_lo[24];
  assign o[24] = scan_lo[24] & N487;
  assign N487 = ~scan_lo[23];
  assign o[23] = scan_lo[23] & N488;
  assign N488 = ~scan_lo[22];
  assign o[22] = scan_lo[22] & N489;
  assign N489 = ~scan_lo[21];
  assign o[21] = scan_lo[21] & N490;
  assign N490 = ~scan_lo[20];
  assign o[20] = scan_lo[20] & N491;
  assign N491 = ~scan_lo[19];
  assign o[19] = scan_lo[19] & N492;
  assign N492 = ~scan_lo[18];
  assign o[18] = scan_lo[18] & N493;
  assign N493 = ~scan_lo[17];
  assign o[17] = scan_lo[17] & N494;
  assign N494 = ~scan_lo[16];
  assign o[16] = scan_lo[16] & N495;
  assign N495 = ~scan_lo[15];
  assign o[15] = scan_lo[15] & N496;
  assign N496 = ~scan_lo[14];
  assign o[14] = scan_lo[14] & N497;
  assign N497 = ~scan_lo[13];
  assign o[13] = scan_lo[13] & N498;
  assign N498 = ~scan_lo[12];
  assign o[12] = scan_lo[12] & N499;
  assign N499 = ~scan_lo[11];
  assign o[11] = scan_lo[11] & N500;
  assign N500 = ~scan_lo[10];
  assign o[10] = scan_lo[10] & N501;
  assign N501 = ~scan_lo[9];
  assign o[9] = scan_lo[9] & N502;
  assign N502 = ~scan_lo[8];
  assign o[8] = scan_lo[8] & N503;
  assign N503 = ~scan_lo[7];
  assign o[7] = scan_lo[7] & N504;
  assign N504 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N505;
  assign N505 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N506;
  assign N506 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N507;
  assign N507 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N508;
  assign N508 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N509;
  assign N509 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N510;
  assign N510 = ~o[0];

endmodule



module bsg_priority_encode_width_p512_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [511:0] i;
  output [8:0] addr_o;
  output v_o;
  wire [8:0] addr_o;
  wire v_o;
  wire [511:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p512_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_width_p512_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_cam_1r1w
(
  clk_i,
  reset_i,
  en_i,
  w_v_i,
  w_set_not_clear_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_data_i,
  r_v_o,
  r_addr_o,
  empty_v_o,
  empty_addr_o
);

  input [8:0] w_addr_i;
  input [15:0] w_data_i;
  input [15:0] r_data_i;
  output [8:0] r_addr_o;
  output [8:0] empty_addr_o;
  input clk_i;
  input reset_i;
  input en_i;
  input w_v_i;
  input w_set_not_clear_i;
  input r_v_i;
  output r_v_o;
  output empty_v_o;
  wire [8:0] r_addr_o,empty_addr_o;
  wire r_v_o,empty_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  matched,empty_found,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,
  N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,
  N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,
  N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,
  N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
  N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,
  N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,
  N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,
  N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,
  N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,
  N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,
  N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,
  N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,
  N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,
  N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,
  N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,
  N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,
  N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,
  N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,
  N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
  N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,
  N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,
  N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,
  N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
  N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,
  N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,
  N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,
  N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,
  N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,
  N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,
  N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,
  N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,
  N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,
  N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
  N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,
  N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,
  N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,
  N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,
  N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,
  N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,
  N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,
  N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,
  N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,
  N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,
  N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,
  N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,
  N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,
  N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,
  N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,
  N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,
  N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,
  N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,
  N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,
  N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,
  N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,
  N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
  N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,
  N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,
  N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
  N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,
  N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,
  N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,
  N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,
  N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,
  N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,
  N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,
  N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,
  N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
  N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,
  N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,
  N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,
  N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,
  N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,
  N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,
  N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,
  N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,
  N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,
  N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,
  N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,
  N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,
  N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,
  N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,
  N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
  N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,
  N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,
  N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,
  N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,
  N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,
  N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,
  N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,
  N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,
  N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
  N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,
  N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,
  N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,
  N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,
  N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,
  N1765,N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,
  N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,
  N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,
  N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,
  N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,
  N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,
  N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,
  N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,
  N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,
  N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,
  N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,
  N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,
  N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,
  N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,
  N1952,N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,
  N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,
  N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,
  N1992,N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,
  N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,
  N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,
  N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,
  N2045,N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,
  N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,
  N2072,N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,
  N2085,N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,
  N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,
  N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,
  N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,
  N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,
  N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,
  N2165,N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,
  N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,
  N2192,N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,
  N2205,N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,
  N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,
  N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,
  N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,
  N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,
  N2272,N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,
  N2285,N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,
  N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,
  N2312,N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,
  N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
  N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,
  N2352,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,
  N2365,N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,
  N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,
  N2392,N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,
  N2405,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,
  N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,
  N2432,N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,
  N2445,N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,
  N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,
  N2472,N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,
  N2485,N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,
  N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,
  N2512,N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,
  N2525,N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,
  N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,
  N2552,N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,
  N2565,N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,
  N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,
  N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,
  N2605,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,
  N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,
  N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,
  N2645,N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,
  N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,
  N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,
  N2685,N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,
  N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,
  N2712,N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,
  N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
  N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,
  N2752,N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,
  N2765,N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,
  N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,
  N2792,N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,
  N2805,N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,
  N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,
  N2832,N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,
  N2845,N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,
  N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,
  N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,
  N2885,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,
  N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,
  N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,
  N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,
  N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,
  N2952,N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,
  N2965,N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,
  N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,
  N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,
  N3005,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,
  N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,
  N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,
  N3045,N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,
  N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,
  N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,
  N3085,N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,
  N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,
  N3112,N3113,N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,
  N3125,N3126,N3127,N3128,N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,
  N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,
  N3152,N3153,N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,
  N3165,N3166,N3167,N3168,N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,
  N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,
  N3192,N3193,N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,
  N3205,N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,
  N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,
  N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,
  N3245,N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,
  N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,
  N3272,N3273,N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,
  N3285,N3286,N3287,N3288,N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,
  N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,
  N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,
  N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,
  N3339,N3340,N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,
  N3352,N3353,N3354,N3355,N3356,N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,
  N3365,N3366,N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,
  N3379,N3380,N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,
  N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,
  N3405,N3406,N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,
  N3419,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,
  N3432,N3433,N3434,N3435,N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,
  N3445,N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,
  N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,
  N3472,N3473,N3474,N3475,N3476,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,
  N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,
  N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,
  N3512,N3513,N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,
  N3525,N3526,N3527,N3528,N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,
  N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,
  N3552,N3553,N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,
  N3565,N3566,N3567,N3568,N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,
  N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,
  N3592,N3593,N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,
  N3605,N3606,N3607,N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,
  N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,
  N3632,N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,
  N3645,N3646,N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,
  N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,
  N3672,N3673,N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,
  N3685,N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,
  N3699,N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,
  N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,
  N3725,N3726,N3727,N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,
  N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,
  N3752,N3753,N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,
  N3765,N3766,N3767,N3768,N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,
  N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,
  N3792,N3793,N3794,N3795,N3796,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,
  N3805,N3806,N3807,N3808,N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,
  N3819,N3820,N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,
  N3832,N3833,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,
  N3845,N3846,N3847,N3848,N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,
  N3859,N3860,N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,
  N3872,N3873,N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,
  N3885,N3886,N3887,N3888,N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,
  N3899,N3900,N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,
  N3912,N3913,N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,
  N3925,N3926,N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,
  N3939,N3940,N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,
  N3952,N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,
  N3965,N3966,N3967,N3968,N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,
  N3979,N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,
  N3992,N3993,N3994,N3995,N3996,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,
  N4005,N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,
  N4019,N4020,N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,
  N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,
  N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,
  N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,
  N4072,N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,
  N4085,N4086,N4087,N4088,N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,
  N4099,N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,
  N4112,N4113,N4114,N4115,N4116,N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,
  N4125,N4126,N4127,N4128,N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,
  N4139,N4140,N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,
  N4152,N4153,N4154,N4155,N4156,N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,
  N4165,N4166,N4167,N4168,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,
  N4179,N4180,N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,
  N4192,N4193,N4194,N4195,N4196,N4197,N4198;
  wire [511:0] match_array,empty_array;
  reg [8191:0] mem;
  reg [511:0] valid;
  assign N1564 = mem[8191:8176] == r_data_i;
  assign N1565 = mem[8175:8160] == r_data_i;
  assign N1566 = mem[8159:8144] == r_data_i;
  assign N1567 = mem[8143:8128] == r_data_i;
  assign N1568 = mem[8127:8112] == r_data_i;
  assign N1569 = mem[8111:8096] == r_data_i;
  assign N1570 = mem[8095:8080] == r_data_i;
  assign N1571 = mem[8079:8064] == r_data_i;
  assign N1572 = mem[8063:8048] == r_data_i;
  assign N1573 = mem[8047:8032] == r_data_i;
  assign N1574 = mem[8031:8016] == r_data_i;
  assign N1575 = mem[8015:8000] == r_data_i;
  assign N1576 = mem[7999:7984] == r_data_i;
  assign N1577 = mem[7983:7968] == r_data_i;
  assign N1578 = mem[7967:7952] == r_data_i;
  assign N1579 = mem[7951:7936] == r_data_i;
  assign N1580 = mem[7935:7920] == r_data_i;
  assign N1581 = mem[7919:7904] == r_data_i;
  assign N1582 = mem[7903:7888] == r_data_i;
  assign N1583 = mem[7887:7872] == r_data_i;
  assign N1584 = mem[7871:7856] == r_data_i;
  assign N1585 = mem[7855:7840] == r_data_i;
  assign N1586 = mem[7839:7824] == r_data_i;
  assign N1587 = mem[7823:7808] == r_data_i;
  assign N1588 = mem[7807:7792] == r_data_i;
  assign N1589 = mem[7791:7776] == r_data_i;
  assign N1590 = mem[7775:7760] == r_data_i;
  assign N1591 = mem[7759:7744] == r_data_i;
  assign N1592 = mem[7743:7728] == r_data_i;
  assign N1593 = mem[7727:7712] == r_data_i;
  assign N1594 = mem[7711:7696] == r_data_i;
  assign N1595 = mem[7695:7680] == r_data_i;
  assign N1596 = mem[7679:7664] == r_data_i;
  assign N1597 = mem[7663:7648] == r_data_i;
  assign N1598 = mem[7647:7632] == r_data_i;
  assign N1599 = mem[7631:7616] == r_data_i;
  assign N1600 = mem[7615:7600] == r_data_i;
  assign N1601 = mem[7599:7584] == r_data_i;
  assign N1602 = mem[7583:7568] == r_data_i;
  assign N1603 = mem[7567:7552] == r_data_i;
  assign N1604 = mem[7551:7536] == r_data_i;
  assign N1605 = mem[7535:7520] == r_data_i;
  assign N1606 = mem[7519:7504] == r_data_i;
  assign N1607 = mem[7503:7488] == r_data_i;
  assign N1608 = mem[7487:7472] == r_data_i;
  assign N1609 = mem[7471:7456] == r_data_i;
  assign N1610 = mem[7455:7440] == r_data_i;
  assign N1611 = mem[7439:7424] == r_data_i;
  assign N1612 = mem[7423:7408] == r_data_i;
  assign N1613 = mem[7407:7392] == r_data_i;
  assign N1614 = mem[7391:7376] == r_data_i;
  assign N1615 = mem[7375:7360] == r_data_i;
  assign N1616 = mem[7359:7344] == r_data_i;
  assign N1617 = mem[7343:7328] == r_data_i;
  assign N1618 = mem[7327:7312] == r_data_i;
  assign N1619 = mem[7311:7296] == r_data_i;
  assign N1620 = mem[7295:7280] == r_data_i;
  assign N1621 = mem[7279:7264] == r_data_i;
  assign N1622 = mem[7263:7248] == r_data_i;
  assign N1623 = mem[7247:7232] == r_data_i;
  assign N1624 = mem[7231:7216] == r_data_i;
  assign N1625 = mem[7215:7200] == r_data_i;
  assign N1626 = mem[7199:7184] == r_data_i;
  assign N1627 = mem[7183:7168] == r_data_i;
  assign N1628 = mem[7167:7152] == r_data_i;
  assign N1629 = mem[7151:7136] == r_data_i;
  assign N1630 = mem[7135:7120] == r_data_i;
  assign N1631 = mem[7119:7104] == r_data_i;
  assign N1632 = mem[7103:7088] == r_data_i;
  assign N1633 = mem[7087:7072] == r_data_i;
  assign N1634 = mem[7071:7056] == r_data_i;
  assign N1635 = mem[7055:7040] == r_data_i;
  assign N1636 = mem[7039:7024] == r_data_i;
  assign N1637 = mem[7023:7008] == r_data_i;
  assign N1638 = mem[7007:6992] == r_data_i;
  assign N1639 = mem[6991:6976] == r_data_i;
  assign N1640 = mem[6975:6960] == r_data_i;
  assign N1641 = mem[6959:6944] == r_data_i;
  assign N1642 = mem[6943:6928] == r_data_i;
  assign N1643 = mem[6927:6912] == r_data_i;
  assign N1644 = mem[6911:6896] == r_data_i;
  assign N1645 = mem[6895:6880] == r_data_i;
  assign N1646 = mem[6879:6864] == r_data_i;
  assign N1647 = mem[6863:6848] == r_data_i;
  assign N1648 = mem[6847:6832] == r_data_i;
  assign N1649 = mem[6831:6816] == r_data_i;
  assign N1650 = mem[6815:6800] == r_data_i;
  assign N1651 = mem[6799:6784] == r_data_i;
  assign N1652 = mem[6783:6768] == r_data_i;
  assign N1653 = mem[6767:6752] == r_data_i;
  assign N1654 = mem[6751:6736] == r_data_i;
  assign N1655 = mem[6735:6720] == r_data_i;
  assign N1656 = mem[6719:6704] == r_data_i;
  assign N1657 = mem[6703:6688] == r_data_i;
  assign N1658 = mem[6687:6672] == r_data_i;
  assign N1659 = mem[6671:6656] == r_data_i;
  assign N1660 = mem[6655:6640] == r_data_i;
  assign N1661 = mem[6639:6624] == r_data_i;
  assign N1662 = mem[6623:6608] == r_data_i;
  assign N1663 = mem[6607:6592] == r_data_i;
  assign N1664 = mem[6591:6576] == r_data_i;
  assign N1665 = mem[6575:6560] == r_data_i;
  assign N1666 = mem[6559:6544] == r_data_i;
  assign N1667 = mem[6543:6528] == r_data_i;
  assign N1668 = mem[6527:6512] == r_data_i;
  assign N1669 = mem[6511:6496] == r_data_i;
  assign N1670 = mem[6495:6480] == r_data_i;
  assign N1671 = mem[6479:6464] == r_data_i;
  assign N1672 = mem[6463:6448] == r_data_i;
  assign N1673 = mem[6447:6432] == r_data_i;
  assign N1674 = mem[6431:6416] == r_data_i;
  assign N1675 = mem[6415:6400] == r_data_i;
  assign N1676 = mem[6399:6384] == r_data_i;
  assign N1677 = mem[6383:6368] == r_data_i;
  assign N1678 = mem[6367:6352] == r_data_i;
  assign N1679 = mem[6351:6336] == r_data_i;
  assign N1680 = mem[6335:6320] == r_data_i;
  assign N1681 = mem[6319:6304] == r_data_i;
  assign N1682 = mem[6303:6288] == r_data_i;
  assign N1683 = mem[6287:6272] == r_data_i;
  assign N1684 = mem[6271:6256] == r_data_i;
  assign N1685 = mem[6255:6240] == r_data_i;
  assign N1686 = mem[6239:6224] == r_data_i;
  assign N1687 = mem[6223:6208] == r_data_i;
  assign N1688 = mem[6207:6192] == r_data_i;
  assign N1689 = mem[6191:6176] == r_data_i;
  assign N1690 = mem[6175:6160] == r_data_i;
  assign N1691 = mem[6159:6144] == r_data_i;
  assign N1692 = mem[6143:6128] == r_data_i;
  assign N1693 = mem[6127:6112] == r_data_i;
  assign N1694 = mem[6111:6096] == r_data_i;
  assign N1695 = mem[6095:6080] == r_data_i;
  assign N1696 = mem[6079:6064] == r_data_i;
  assign N1697 = mem[6063:6048] == r_data_i;
  assign N1698 = mem[6047:6032] == r_data_i;
  assign N1699 = mem[6031:6016] == r_data_i;
  assign N1700 = mem[6015:6000] == r_data_i;
  assign N1701 = mem[5999:5984] == r_data_i;
  assign N1702 = mem[5983:5968] == r_data_i;
  assign N1703 = mem[5967:5952] == r_data_i;
  assign N1704 = mem[5951:5936] == r_data_i;
  assign N1705 = mem[5935:5920] == r_data_i;
  assign N1706 = mem[5919:5904] == r_data_i;
  assign N1707 = mem[5903:5888] == r_data_i;
  assign N1708 = mem[5887:5872] == r_data_i;
  assign N1709 = mem[5871:5856] == r_data_i;
  assign N1710 = mem[5855:5840] == r_data_i;
  assign N1711 = mem[5839:5824] == r_data_i;
  assign N1712 = mem[5823:5808] == r_data_i;
  assign N1713 = mem[5807:5792] == r_data_i;
  assign N1714 = mem[5791:5776] == r_data_i;
  assign N1715 = mem[5775:5760] == r_data_i;
  assign N1716 = mem[5759:5744] == r_data_i;
  assign N1717 = mem[5743:5728] == r_data_i;
  assign N1718 = mem[5727:5712] == r_data_i;
  assign N1719 = mem[5711:5696] == r_data_i;
  assign N1720 = mem[5695:5680] == r_data_i;
  assign N1721 = mem[5679:5664] == r_data_i;
  assign N1722 = mem[5663:5648] == r_data_i;
  assign N1723 = mem[5647:5632] == r_data_i;
  assign N1724 = mem[5631:5616] == r_data_i;
  assign N1725 = mem[5615:5600] == r_data_i;
  assign N1726 = mem[5599:5584] == r_data_i;
  assign N1727 = mem[5583:5568] == r_data_i;
  assign N1728 = mem[5567:5552] == r_data_i;
  assign N1729 = mem[5551:5536] == r_data_i;
  assign N1730 = mem[5535:5520] == r_data_i;
  assign N1731 = mem[5519:5504] == r_data_i;
  assign N1732 = mem[5503:5488] == r_data_i;
  assign N1733 = mem[5487:5472] == r_data_i;
  assign N1734 = mem[5471:5456] == r_data_i;
  assign N1735 = mem[5455:5440] == r_data_i;
  assign N1736 = mem[5439:5424] == r_data_i;
  assign N1737 = mem[5423:5408] == r_data_i;
  assign N1738 = mem[5407:5392] == r_data_i;
  assign N1739 = mem[5391:5376] == r_data_i;
  assign N1740 = mem[5375:5360] == r_data_i;
  assign N1741 = mem[5359:5344] == r_data_i;
  assign N1742 = mem[5343:5328] == r_data_i;
  assign N1743 = mem[5327:5312] == r_data_i;
  assign N1744 = mem[5311:5296] == r_data_i;
  assign N1745 = mem[5295:5280] == r_data_i;
  assign N1746 = mem[5279:5264] == r_data_i;
  assign N1747 = mem[5263:5248] == r_data_i;
  assign N1748 = mem[5247:5232] == r_data_i;
  assign N1749 = mem[5231:5216] == r_data_i;
  assign N1750 = mem[5215:5200] == r_data_i;
  assign N1751 = mem[5199:5184] == r_data_i;
  assign N1752 = mem[5183:5168] == r_data_i;
  assign N1753 = mem[5167:5152] == r_data_i;
  assign N1754 = mem[5151:5136] == r_data_i;
  assign N1755 = mem[5135:5120] == r_data_i;
  assign N1756 = mem[5119:5104] == r_data_i;
  assign N1757 = mem[5103:5088] == r_data_i;
  assign N1758 = mem[5087:5072] == r_data_i;
  assign N1759 = mem[5071:5056] == r_data_i;
  assign N1760 = mem[5055:5040] == r_data_i;
  assign N1761 = mem[5039:5024] == r_data_i;
  assign N1762 = mem[5023:5008] == r_data_i;
  assign N1763 = mem[5007:4992] == r_data_i;
  assign N1764 = mem[4991:4976] == r_data_i;
  assign N1765 = mem[4975:4960] == r_data_i;
  assign N1766 = mem[4959:4944] == r_data_i;
  assign N1767 = mem[4943:4928] == r_data_i;
  assign N1768 = mem[4927:4912] == r_data_i;
  assign N1769 = mem[4911:4896] == r_data_i;
  assign N1770 = mem[4895:4880] == r_data_i;
  assign N1771 = mem[4879:4864] == r_data_i;
  assign N1772 = mem[4863:4848] == r_data_i;
  assign N1773 = mem[4847:4832] == r_data_i;
  assign N1774 = mem[4831:4816] == r_data_i;
  assign N1775 = mem[4815:4800] == r_data_i;
  assign N1776 = mem[4799:4784] == r_data_i;
  assign N1777 = mem[4783:4768] == r_data_i;
  assign N1778 = mem[4767:4752] == r_data_i;
  assign N1779 = mem[4751:4736] == r_data_i;
  assign N1780 = mem[4735:4720] == r_data_i;
  assign N1781 = mem[4719:4704] == r_data_i;
  assign N1782 = mem[4703:4688] == r_data_i;
  assign N1783 = mem[4687:4672] == r_data_i;
  assign N1784 = mem[4671:4656] == r_data_i;
  assign N1785 = mem[4655:4640] == r_data_i;
  assign N1786 = mem[4639:4624] == r_data_i;
  assign N1787 = mem[4623:4608] == r_data_i;
  assign N1788 = mem[4607:4592] == r_data_i;
  assign N1789 = mem[4591:4576] == r_data_i;
  assign N1790 = mem[4575:4560] == r_data_i;
  assign N1791 = mem[4559:4544] == r_data_i;
  assign N1792 = mem[4543:4528] == r_data_i;
  assign N1793 = mem[4527:4512] == r_data_i;
  assign N1794 = mem[4511:4496] == r_data_i;
  assign N1795 = mem[4495:4480] == r_data_i;
  assign N1796 = mem[4479:4464] == r_data_i;
  assign N1797 = mem[4463:4448] == r_data_i;
  assign N1798 = mem[4447:4432] == r_data_i;
  assign N1799 = mem[4431:4416] == r_data_i;
  assign N1800 = mem[4415:4400] == r_data_i;
  assign N1801 = mem[4399:4384] == r_data_i;
  assign N1802 = mem[4383:4368] == r_data_i;
  assign N1803 = mem[4367:4352] == r_data_i;
  assign N1804 = mem[4351:4336] == r_data_i;
  assign N1805 = mem[4335:4320] == r_data_i;
  assign N1806 = mem[4319:4304] == r_data_i;
  assign N1807 = mem[4303:4288] == r_data_i;
  assign N1808 = mem[4287:4272] == r_data_i;
  assign N1809 = mem[4271:4256] == r_data_i;
  assign N1810 = mem[4255:4240] == r_data_i;
  assign N1811 = mem[4239:4224] == r_data_i;
  assign N1812 = mem[4223:4208] == r_data_i;
  assign N1813 = mem[4207:4192] == r_data_i;
  assign N1814 = mem[4191:4176] == r_data_i;
  assign N1815 = mem[4175:4160] == r_data_i;
  assign N1816 = mem[4159:4144] == r_data_i;
  assign N1817 = mem[4143:4128] == r_data_i;
  assign N1818 = mem[4127:4112] == r_data_i;
  assign N1819 = mem[4111:4096] == r_data_i;
  assign N1820 = mem[4095:4080] == r_data_i;
  assign N1821 = mem[4079:4064] == r_data_i;
  assign N1822 = mem[4063:4048] == r_data_i;
  assign N1823 = mem[4047:4032] == r_data_i;
  assign N1824 = mem[4031:4016] == r_data_i;
  assign N1825 = mem[4015:4000] == r_data_i;
  assign N1826 = mem[3999:3984] == r_data_i;
  assign N1827 = mem[3983:3968] == r_data_i;
  assign N1828 = mem[3967:3952] == r_data_i;
  assign N1829 = mem[3951:3936] == r_data_i;
  assign N1830 = mem[3935:3920] == r_data_i;
  assign N1831 = mem[3919:3904] == r_data_i;
  assign N1832 = mem[3903:3888] == r_data_i;
  assign N1833 = mem[3887:3872] == r_data_i;
  assign N1834 = mem[3871:3856] == r_data_i;
  assign N1835 = mem[3855:3840] == r_data_i;
  assign N1836 = mem[3839:3824] == r_data_i;
  assign N1837 = mem[3823:3808] == r_data_i;
  assign N1838 = mem[3807:3792] == r_data_i;
  assign N1839 = mem[3791:3776] == r_data_i;
  assign N1840 = mem[3775:3760] == r_data_i;
  assign N1841 = mem[3759:3744] == r_data_i;
  assign N1842 = mem[3743:3728] == r_data_i;
  assign N1843 = mem[3727:3712] == r_data_i;
  assign N1844 = mem[3711:3696] == r_data_i;
  assign N1845 = mem[3695:3680] == r_data_i;
  assign N1846 = mem[3679:3664] == r_data_i;
  assign N1847 = mem[3663:3648] == r_data_i;
  assign N1848 = mem[3647:3632] == r_data_i;
  assign N1849 = mem[3631:3616] == r_data_i;
  assign N1850 = mem[3615:3600] == r_data_i;
  assign N1851 = mem[3599:3584] == r_data_i;
  assign N1852 = mem[3583:3568] == r_data_i;
  assign N1853 = mem[3567:3552] == r_data_i;
  assign N1854 = mem[3551:3536] == r_data_i;
  assign N1855 = mem[3535:3520] == r_data_i;
  assign N1856 = mem[3519:3504] == r_data_i;
  assign N1857 = mem[3503:3488] == r_data_i;
  assign N1858 = mem[3487:3472] == r_data_i;
  assign N1859 = mem[3471:3456] == r_data_i;
  assign N1860 = mem[3455:3440] == r_data_i;
  assign N1861 = mem[3439:3424] == r_data_i;
  assign N1862 = mem[3423:3408] == r_data_i;
  assign N1863 = mem[3407:3392] == r_data_i;
  assign N1864 = mem[3391:3376] == r_data_i;
  assign N1865 = mem[3375:3360] == r_data_i;
  assign N1866 = mem[3359:3344] == r_data_i;
  assign N1867 = mem[3343:3328] == r_data_i;
  assign N1868 = mem[3327:3312] == r_data_i;
  assign N1869 = mem[3311:3296] == r_data_i;
  assign N1870 = mem[3295:3280] == r_data_i;
  assign N1871 = mem[3279:3264] == r_data_i;
  assign N1872 = mem[3263:3248] == r_data_i;
  assign N1873 = mem[3247:3232] == r_data_i;
  assign N1874 = mem[3231:3216] == r_data_i;
  assign N1875 = mem[3215:3200] == r_data_i;
  assign N1876 = mem[3199:3184] == r_data_i;
  assign N1877 = mem[3183:3168] == r_data_i;
  assign N1878 = mem[3167:3152] == r_data_i;
  assign N1879 = mem[3151:3136] == r_data_i;
  assign N1880 = mem[3135:3120] == r_data_i;
  assign N1881 = mem[3119:3104] == r_data_i;
  assign N1882 = mem[3103:3088] == r_data_i;
  assign N1883 = mem[3087:3072] == r_data_i;
  assign N1884 = mem[3071:3056] == r_data_i;
  assign N1885 = mem[3055:3040] == r_data_i;
  assign N1886 = mem[3039:3024] == r_data_i;
  assign N1887 = mem[3023:3008] == r_data_i;
  assign N1888 = mem[3007:2992] == r_data_i;
  assign N1889 = mem[2991:2976] == r_data_i;
  assign N1890 = mem[2975:2960] == r_data_i;
  assign N1891 = mem[2959:2944] == r_data_i;
  assign N1892 = mem[2943:2928] == r_data_i;
  assign N1893 = mem[2927:2912] == r_data_i;
  assign N1894 = mem[2911:2896] == r_data_i;
  assign N1895 = mem[2895:2880] == r_data_i;
  assign N1896 = mem[2879:2864] == r_data_i;
  assign N1897 = mem[2863:2848] == r_data_i;
  assign N1898 = mem[2847:2832] == r_data_i;
  assign N1899 = mem[2831:2816] == r_data_i;
  assign N1900 = mem[2815:2800] == r_data_i;
  assign N1901 = mem[2799:2784] == r_data_i;
  assign N1902 = mem[2783:2768] == r_data_i;
  assign N1903 = mem[2767:2752] == r_data_i;
  assign N1904 = mem[2751:2736] == r_data_i;
  assign N1905 = mem[2735:2720] == r_data_i;
  assign N1906 = mem[2719:2704] == r_data_i;
  assign N1907 = mem[2703:2688] == r_data_i;
  assign N1908 = mem[2687:2672] == r_data_i;
  assign N1909 = mem[2671:2656] == r_data_i;
  assign N1910 = mem[2655:2640] == r_data_i;
  assign N1911 = mem[2639:2624] == r_data_i;
  assign N1912 = mem[2623:2608] == r_data_i;
  assign N1913 = mem[2607:2592] == r_data_i;
  assign N1914 = mem[2591:2576] == r_data_i;
  assign N1915 = mem[2575:2560] == r_data_i;
  assign N1916 = mem[2559:2544] == r_data_i;
  assign N1917 = mem[2543:2528] == r_data_i;
  assign N1918 = mem[2527:2512] == r_data_i;
  assign N1919 = mem[2511:2496] == r_data_i;
  assign N1920 = mem[2495:2480] == r_data_i;
  assign N1921 = mem[2479:2464] == r_data_i;
  assign N1922 = mem[2463:2448] == r_data_i;
  assign N1923 = mem[2447:2432] == r_data_i;
  assign N1924 = mem[2431:2416] == r_data_i;
  assign N1925 = mem[2415:2400] == r_data_i;
  assign N1926 = mem[2399:2384] == r_data_i;
  assign N1927 = mem[2383:2368] == r_data_i;
  assign N1928 = mem[2367:2352] == r_data_i;
  assign N1929 = mem[2351:2336] == r_data_i;
  assign N1930 = mem[2335:2320] == r_data_i;
  assign N1931 = mem[2319:2304] == r_data_i;
  assign N1932 = mem[2303:2288] == r_data_i;
  assign N1933 = mem[2287:2272] == r_data_i;
  assign N1934 = mem[2271:2256] == r_data_i;
  assign N1935 = mem[2255:2240] == r_data_i;
  assign N1936 = mem[2239:2224] == r_data_i;
  assign N1937 = mem[2223:2208] == r_data_i;
  assign N1938 = mem[2207:2192] == r_data_i;
  assign N1939 = mem[2191:2176] == r_data_i;
  assign N1940 = mem[2175:2160] == r_data_i;
  assign N1941 = mem[2159:2144] == r_data_i;
  assign N1942 = mem[2143:2128] == r_data_i;
  assign N1943 = mem[2127:2112] == r_data_i;
  assign N1944 = mem[2111:2096] == r_data_i;
  assign N1945 = mem[2095:2080] == r_data_i;
  assign N1946 = mem[2079:2064] == r_data_i;
  assign N1947 = mem[2063:2048] == r_data_i;
  assign N1948 = mem[2047:2032] == r_data_i;
  assign N1949 = mem[2031:2016] == r_data_i;
  assign N1950 = mem[2015:2000] == r_data_i;
  assign N1951 = mem[1999:1984] == r_data_i;
  assign N1952 = mem[1983:1968] == r_data_i;
  assign N1953 = mem[1967:1952] == r_data_i;
  assign N1954 = mem[1951:1936] == r_data_i;
  assign N1955 = mem[1935:1920] == r_data_i;
  assign N1956 = mem[1919:1904] == r_data_i;
  assign N1957 = mem[1903:1888] == r_data_i;
  assign N1958 = mem[1887:1872] == r_data_i;
  assign N1959 = mem[1871:1856] == r_data_i;
  assign N1960 = mem[1855:1840] == r_data_i;
  assign N1961 = mem[1839:1824] == r_data_i;
  assign N1962 = mem[1823:1808] == r_data_i;
  assign N1963 = mem[1807:1792] == r_data_i;
  assign N1964 = mem[1791:1776] == r_data_i;
  assign N1965 = mem[1775:1760] == r_data_i;
  assign N1966 = mem[1759:1744] == r_data_i;
  assign N1967 = mem[1743:1728] == r_data_i;
  assign N1968 = mem[1727:1712] == r_data_i;
  assign N1969 = mem[1711:1696] == r_data_i;
  assign N1970 = mem[1695:1680] == r_data_i;
  assign N1971 = mem[1679:1664] == r_data_i;
  assign N1972 = mem[1663:1648] == r_data_i;
  assign N1973 = mem[1647:1632] == r_data_i;
  assign N1974 = mem[1631:1616] == r_data_i;
  assign N1975 = mem[1615:1600] == r_data_i;
  assign N1976 = mem[1599:1584] == r_data_i;
  assign N1977 = mem[1583:1568] == r_data_i;
  assign N1978 = mem[1567:1552] == r_data_i;
  assign N1979 = mem[1551:1536] == r_data_i;
  assign N1980 = mem[1535:1520] == r_data_i;
  assign N1981 = mem[1519:1504] == r_data_i;
  assign N1982 = mem[1503:1488] == r_data_i;
  assign N1983 = mem[1487:1472] == r_data_i;
  assign N1984 = mem[1471:1456] == r_data_i;
  assign N1985 = mem[1455:1440] == r_data_i;
  assign N1986 = mem[1439:1424] == r_data_i;
  assign N1987 = mem[1423:1408] == r_data_i;
  assign N1988 = mem[1407:1392] == r_data_i;
  assign N1989 = mem[1391:1376] == r_data_i;
  assign N1990 = mem[1375:1360] == r_data_i;
  assign N1991 = mem[1359:1344] == r_data_i;
  assign N1992 = mem[1343:1328] == r_data_i;
  assign N1993 = mem[1327:1312] == r_data_i;
  assign N1994 = mem[1311:1296] == r_data_i;
  assign N1995 = mem[1295:1280] == r_data_i;
  assign N1996 = mem[1279:1264] == r_data_i;
  assign N1997 = mem[1263:1248] == r_data_i;
  assign N1998 = mem[1247:1232] == r_data_i;
  assign N1999 = mem[1231:1216] == r_data_i;
  assign N2000 = mem[1215:1200] == r_data_i;
  assign N2001 = mem[1199:1184] == r_data_i;
  assign N2002 = mem[1183:1168] == r_data_i;
  assign N2003 = mem[1167:1152] == r_data_i;
  assign N2004 = mem[1151:1136] == r_data_i;
  assign N2005 = mem[1135:1120] == r_data_i;
  assign N2006 = mem[1119:1104] == r_data_i;
  assign N2007 = mem[1103:1088] == r_data_i;
  assign N2008 = mem[1087:1072] == r_data_i;
  assign N2009 = mem[1071:1056] == r_data_i;
  assign N2010 = mem[1055:1040] == r_data_i;
  assign N2011 = mem[1039:1024] == r_data_i;
  assign N2012 = mem[1023:1008] == r_data_i;
  assign N2013 = mem[1007:992] == r_data_i;
  assign N2014 = mem[991:976] == r_data_i;
  assign N2015 = mem[975:960] == r_data_i;
  assign N2016 = mem[959:944] == r_data_i;
  assign N2017 = mem[943:928] == r_data_i;
  assign N2018 = mem[927:912] == r_data_i;
  assign N2019 = mem[911:896] == r_data_i;
  assign N2020 = mem[895:880] == r_data_i;
  assign N2021 = mem[879:864] == r_data_i;
  assign N2022 = mem[863:848] == r_data_i;
  assign N2023 = mem[847:832] == r_data_i;
  assign N2024 = mem[831:816] == r_data_i;
  assign N2025 = mem[815:800] == r_data_i;
  assign N2026 = mem[799:784] == r_data_i;
  assign N2027 = mem[783:768] == r_data_i;
  assign N2028 = mem[767:752] == r_data_i;
  assign N2029 = mem[751:736] == r_data_i;
  assign N2030 = mem[735:720] == r_data_i;
  assign N2031 = mem[719:704] == r_data_i;
  assign N2032 = mem[703:688] == r_data_i;
  assign N2033 = mem[687:672] == r_data_i;
  assign N2034 = mem[671:656] == r_data_i;
  assign N2035 = mem[655:640] == r_data_i;
  assign N2036 = mem[639:624] == r_data_i;
  assign N2037 = mem[623:608] == r_data_i;
  assign N2038 = mem[607:592] == r_data_i;
  assign N2039 = mem[591:576] == r_data_i;
  assign N2040 = mem[575:560] == r_data_i;
  assign N2041 = mem[559:544] == r_data_i;
  assign N2042 = mem[543:528] == r_data_i;
  assign N2043 = mem[527:512] == r_data_i;
  assign N2044 = mem[511:496] == r_data_i;
  assign N2045 = mem[495:480] == r_data_i;
  assign N2046 = mem[479:464] == r_data_i;
  assign N2047 = mem[463:448] == r_data_i;
  assign N2048 = mem[447:432] == r_data_i;
  assign N2049 = mem[431:416] == r_data_i;
  assign N2050 = mem[415:400] == r_data_i;
  assign N2051 = mem[399:384] == r_data_i;
  assign N2052 = mem[383:368] == r_data_i;
  assign N2053 = mem[367:352] == r_data_i;
  assign N2054 = mem[351:336] == r_data_i;
  assign N2055 = mem[335:320] == r_data_i;
  assign N2056 = mem[319:304] == r_data_i;
  assign N2057 = mem[303:288] == r_data_i;
  assign N2058 = mem[287:272] == r_data_i;
  assign N2059 = mem[271:256] == r_data_i;
  assign N2060 = mem[255:240] == r_data_i;
  assign N2061 = mem[239:224] == r_data_i;
  assign N2062 = mem[223:208] == r_data_i;
  assign N2063 = mem[207:192] == r_data_i;
  assign N2064 = mem[191:176] == r_data_i;
  assign N2065 = mem[175:160] == r_data_i;
  assign N2066 = mem[159:144] == r_data_i;
  assign N2067 = mem[143:128] == r_data_i;
  assign N2068 = mem[127:112] == r_data_i;
  assign N2069 = mem[111:96] == r_data_i;
  assign N2070 = mem[95:80] == r_data_i;
  assign N2071 = mem[79:64] == r_data_i;
  assign N2072 = mem[63:48] == r_data_i;
  assign N2073 = mem[47:32] == r_data_i;
  assign N2074 = mem[31:16] == r_data_i;
  assign N2075 = mem[15:0] == r_data_i;

  bsg_encode_one_hot_width_p512_lo_to_hi_p1
  fi4_ohe
  (
    .i(match_array),
    .addr_o(r_addr_o),
    .v_o(matched)
  );


  bsg_priority_encode_width_p512_lo_to_hi_p1
  fi5_epe
  (
    .i(empty_array),
    .addr_o(empty_addr_o),
    .v_o(empty_found)
  );

  assign N2076 = w_addr_i[7] & w_addr_i[8];
  assign N2077 = N0 & w_addr_i[8];
  assign N0 = ~w_addr_i[7];
  assign N2078 = w_addr_i[7] & N1;
  assign N1 = ~w_addr_i[8];
  assign N2079 = N2 & N3;
  assign N2 = ~w_addr_i[7];
  assign N3 = ~w_addr_i[8];
  assign N2080 = w_addr_i[5] & w_addr_i[6];
  assign N2081 = N4 & w_addr_i[6];
  assign N4 = ~w_addr_i[5];
  assign N2082 = w_addr_i[5] & N5;
  assign N5 = ~w_addr_i[6];
  assign N2083 = N6 & N7;
  assign N6 = ~w_addr_i[5];
  assign N7 = ~w_addr_i[6];
  assign N2084 = N2076 & N2080;
  assign N2085 = N2076 & N2081;
  assign N2086 = N2076 & N2082;
  assign N2087 = N2076 & N2083;
  assign N2088 = N2077 & N2080;
  assign N2089 = N2077 & N2081;
  assign N2090 = N2077 & N2082;
  assign N2091 = N2077 & N2083;
  assign N2092 = N2078 & N2080;
  assign N2093 = N2078 & N2081;
  assign N2094 = N2078 & N2082;
  assign N2095 = N2078 & N2083;
  assign N2096 = N2079 & N2080;
  assign N2097 = N2079 & N2081;
  assign N2098 = N2079 & N2082;
  assign N2099 = N2079 & N2083;
  assign N2100 = w_addr_i[3] & w_addr_i[4];
  assign N2101 = N8 & w_addr_i[4];
  assign N8 = ~w_addr_i[3];
  assign N2102 = w_addr_i[3] & N9;
  assign N9 = ~w_addr_i[4];
  assign N2103 = N10 & N11;
  assign N10 = ~w_addr_i[3];
  assign N11 = ~w_addr_i[4];
  assign N2104 = ~w_addr_i[2];
  assign N2105 = w_addr_i[0] & w_addr_i[1];
  assign N2106 = N12 & w_addr_i[1];
  assign N12 = ~w_addr_i[0];
  assign N2107 = w_addr_i[0] & N13;
  assign N13 = ~w_addr_i[1];
  assign N2108 = N14 & N15;
  assign N14 = ~w_addr_i[0];
  assign N15 = ~w_addr_i[1];
  assign N2109 = w_addr_i[2] & N2105;
  assign N2110 = w_addr_i[2] & N2106;
  assign N2111 = w_addr_i[2] & N2107;
  assign N2112 = w_addr_i[2] & N2108;
  assign N2113 = N2104 & N2105;
  assign N2114 = N2104 & N2106;
  assign N2115 = N2104 & N2107;
  assign N2116 = N2104 & N2108;
  assign N2117 = N2100 & N2109;
  assign N2118 = N2100 & N2110;
  assign N2119 = N2100 & N2111;
  assign N2120 = N2100 & N2112;
  assign N2121 = N2100 & N2113;
  assign N2122 = N2100 & N2114;
  assign N2123 = N2100 & N2115;
  assign N2124 = N2100 & N2116;
  assign N2125 = N2101 & N2109;
  assign N2126 = N2101 & N2110;
  assign N2127 = N2101 & N2111;
  assign N2128 = N2101 & N2112;
  assign N2129 = N2101 & N2113;
  assign N2130 = N2101 & N2114;
  assign N2131 = N2101 & N2115;
  assign N2132 = N2101 & N2116;
  assign N2133 = N2102 & N2109;
  assign N2134 = N2102 & N2110;
  assign N2135 = N2102 & N2111;
  assign N2136 = N2102 & N2112;
  assign N2137 = N2102 & N2113;
  assign N2138 = N2102 & N2114;
  assign N2139 = N2102 & N2115;
  assign N2140 = N2102 & N2116;
  assign N2141 = N2103 & N2109;
  assign N2142 = N2103 & N2110;
  assign N2143 = N2103 & N2111;
  assign N2144 = N2103 & N2112;
  assign N2145 = N2103 & N2113;
  assign N2146 = N2103 & N2114;
  assign N2147 = N2103 & N2115;
  assign N2148 = N2103 & N2116;
  assign N531 = N2084 & N2117;
  assign N530 = N2084 & N2118;
  assign N529 = N2084 & N2119;
  assign N528 = N2084 & N2120;
  assign N527 = N2084 & N2121;
  assign N526 = N2084 & N2122;
  assign N525 = N2084 & N2123;
  assign N524 = N2084 & N2124;
  assign N523 = N2084 & N2125;
  assign N522 = N2084 & N2126;
  assign N521 = N2084 & N2127;
  assign N520 = N2084 & N2128;
  assign N519 = N2084 & N2129;
  assign N518 = N2084 & N2130;
  assign N517 = N2084 & N2131;
  assign N516 = N2084 & N2132;
  assign N515 = N2084 & N2133;
  assign N514 = N2084 & N2134;
  assign N513 = N2084 & N2135;
  assign N512 = N2084 & N2136;
  assign N511 = N2084 & N2137;
  assign N510 = N2084 & N2138;
  assign N509 = N2084 & N2139;
  assign N508 = N2084 & N2140;
  assign N507 = N2084 & N2141;
  assign N506 = N2084 & N2142;
  assign N505 = N2084 & N2143;
  assign N504 = N2084 & N2144;
  assign N503 = N2084 & N2145;
  assign N502 = N2084 & N2146;
  assign N501 = N2084 & N2147;
  assign N500 = N2084 & N2148;
  assign N499 = N2085 & N2117;
  assign N498 = N2085 & N2118;
  assign N497 = N2085 & N2119;
  assign N496 = N2085 & N2120;
  assign N495 = N2085 & N2121;
  assign N494 = N2085 & N2122;
  assign N493 = N2085 & N2123;
  assign N492 = N2085 & N2124;
  assign N491 = N2085 & N2125;
  assign N490 = N2085 & N2126;
  assign N489 = N2085 & N2127;
  assign N488 = N2085 & N2128;
  assign N487 = N2085 & N2129;
  assign N486 = N2085 & N2130;
  assign N485 = N2085 & N2131;
  assign N484 = N2085 & N2132;
  assign N483 = N2085 & N2133;
  assign N482 = N2085 & N2134;
  assign N481 = N2085 & N2135;
  assign N480 = N2085 & N2136;
  assign N479 = N2085 & N2137;
  assign N478 = N2085 & N2138;
  assign N477 = N2085 & N2139;
  assign N476 = N2085 & N2140;
  assign N475 = N2085 & N2141;
  assign N474 = N2085 & N2142;
  assign N473 = N2085 & N2143;
  assign N472 = N2085 & N2144;
  assign N471 = N2085 & N2145;
  assign N470 = N2085 & N2146;
  assign N469 = N2085 & N2147;
  assign N468 = N2085 & N2148;
  assign N467 = N2086 & N2117;
  assign N466 = N2086 & N2118;
  assign N465 = N2086 & N2119;
  assign N464 = N2086 & N2120;
  assign N463 = N2086 & N2121;
  assign N462 = N2086 & N2122;
  assign N461 = N2086 & N2123;
  assign N460 = N2086 & N2124;
  assign N459 = N2086 & N2125;
  assign N458 = N2086 & N2126;
  assign N457 = N2086 & N2127;
  assign N456 = N2086 & N2128;
  assign N455 = N2086 & N2129;
  assign N454 = N2086 & N2130;
  assign N453 = N2086 & N2131;
  assign N452 = N2086 & N2132;
  assign N451 = N2086 & N2133;
  assign N450 = N2086 & N2134;
  assign N449 = N2086 & N2135;
  assign N448 = N2086 & N2136;
  assign N447 = N2086 & N2137;
  assign N446 = N2086 & N2138;
  assign N445 = N2086 & N2139;
  assign N444 = N2086 & N2140;
  assign N443 = N2086 & N2141;
  assign N442 = N2086 & N2142;
  assign N441 = N2086 & N2143;
  assign N440 = N2086 & N2144;
  assign N439 = N2086 & N2145;
  assign N438 = N2086 & N2146;
  assign N437 = N2086 & N2147;
  assign N436 = N2086 & N2148;
  assign N435 = N2087 & N2117;
  assign N434 = N2087 & N2118;
  assign N433 = N2087 & N2119;
  assign N432 = N2087 & N2120;
  assign N431 = N2087 & N2121;
  assign N430 = N2087 & N2122;
  assign N429 = N2087 & N2123;
  assign N428 = N2087 & N2124;
  assign N427 = N2087 & N2125;
  assign N426 = N2087 & N2126;
  assign N425 = N2087 & N2127;
  assign N424 = N2087 & N2128;
  assign N423 = N2087 & N2129;
  assign N422 = N2087 & N2130;
  assign N421 = N2087 & N2131;
  assign N420 = N2087 & N2132;
  assign N419 = N2087 & N2133;
  assign N418 = N2087 & N2134;
  assign N417 = N2087 & N2135;
  assign N416 = N2087 & N2136;
  assign N415 = N2087 & N2137;
  assign N414 = N2087 & N2138;
  assign N413 = N2087 & N2139;
  assign N412 = N2087 & N2140;
  assign N411 = N2087 & N2141;
  assign N410 = N2087 & N2142;
  assign N409 = N2087 & N2143;
  assign N408 = N2087 & N2144;
  assign N407 = N2087 & N2145;
  assign N406 = N2087 & N2146;
  assign N405 = N2087 & N2147;
  assign N404 = N2087 & N2148;
  assign N403 = N2088 & N2117;
  assign N402 = N2088 & N2118;
  assign N401 = N2088 & N2119;
  assign N400 = N2088 & N2120;
  assign N399 = N2088 & N2121;
  assign N398 = N2088 & N2122;
  assign N397 = N2088 & N2123;
  assign N396 = N2088 & N2124;
  assign N395 = N2088 & N2125;
  assign N394 = N2088 & N2126;
  assign N393 = N2088 & N2127;
  assign N392 = N2088 & N2128;
  assign N391 = N2088 & N2129;
  assign N390 = N2088 & N2130;
  assign N389 = N2088 & N2131;
  assign N388 = N2088 & N2132;
  assign N387 = N2088 & N2133;
  assign N386 = N2088 & N2134;
  assign N385 = N2088 & N2135;
  assign N384 = N2088 & N2136;
  assign N383 = N2088 & N2137;
  assign N382 = N2088 & N2138;
  assign N381 = N2088 & N2139;
  assign N380 = N2088 & N2140;
  assign N379 = N2088 & N2141;
  assign N378 = N2088 & N2142;
  assign N377 = N2088 & N2143;
  assign N376 = N2088 & N2144;
  assign N375 = N2088 & N2145;
  assign N374 = N2088 & N2146;
  assign N373 = N2088 & N2147;
  assign N372 = N2088 & N2148;
  assign N371 = N2089 & N2117;
  assign N370 = N2089 & N2118;
  assign N369 = N2089 & N2119;
  assign N368 = N2089 & N2120;
  assign N367 = N2089 & N2121;
  assign N366 = N2089 & N2122;
  assign N365 = N2089 & N2123;
  assign N364 = N2089 & N2124;
  assign N363 = N2089 & N2125;
  assign N362 = N2089 & N2126;
  assign N361 = N2089 & N2127;
  assign N360 = N2089 & N2128;
  assign N359 = N2089 & N2129;
  assign N358 = N2089 & N2130;
  assign N357 = N2089 & N2131;
  assign N356 = N2089 & N2132;
  assign N355 = N2089 & N2133;
  assign N354 = N2089 & N2134;
  assign N353 = N2089 & N2135;
  assign N352 = N2089 & N2136;
  assign N351 = N2089 & N2137;
  assign N350 = N2089 & N2138;
  assign N349 = N2089 & N2139;
  assign N348 = N2089 & N2140;
  assign N347 = N2089 & N2141;
  assign N346 = N2089 & N2142;
  assign N345 = N2089 & N2143;
  assign N344 = N2089 & N2144;
  assign N343 = N2089 & N2145;
  assign N342 = N2089 & N2146;
  assign N341 = N2089 & N2147;
  assign N340 = N2089 & N2148;
  assign N339 = N2090 & N2117;
  assign N338 = N2090 & N2118;
  assign N337 = N2090 & N2119;
  assign N336 = N2090 & N2120;
  assign N335 = N2090 & N2121;
  assign N334 = N2090 & N2122;
  assign N333 = N2090 & N2123;
  assign N332 = N2090 & N2124;
  assign N331 = N2090 & N2125;
  assign N330 = N2090 & N2126;
  assign N329 = N2090 & N2127;
  assign N328 = N2090 & N2128;
  assign N327 = N2090 & N2129;
  assign N326 = N2090 & N2130;
  assign N325 = N2090 & N2131;
  assign N324 = N2090 & N2132;
  assign N323 = N2090 & N2133;
  assign N322 = N2090 & N2134;
  assign N321 = N2090 & N2135;
  assign N320 = N2090 & N2136;
  assign N319 = N2090 & N2137;
  assign N318 = N2090 & N2138;
  assign N317 = N2090 & N2139;
  assign N316 = N2090 & N2140;
  assign N315 = N2090 & N2141;
  assign N314 = N2090 & N2142;
  assign N313 = N2090 & N2143;
  assign N312 = N2090 & N2144;
  assign N311 = N2090 & N2145;
  assign N310 = N2090 & N2146;
  assign N309 = N2090 & N2147;
  assign N308 = N2090 & N2148;
  assign N307 = N2091 & N2117;
  assign N306 = N2091 & N2118;
  assign N305 = N2091 & N2119;
  assign N304 = N2091 & N2120;
  assign N303 = N2091 & N2121;
  assign N302 = N2091 & N2122;
  assign N301 = N2091 & N2123;
  assign N300 = N2091 & N2124;
  assign N299 = N2091 & N2125;
  assign N298 = N2091 & N2126;
  assign N297 = N2091 & N2127;
  assign N296 = N2091 & N2128;
  assign N295 = N2091 & N2129;
  assign N294 = N2091 & N2130;
  assign N293 = N2091 & N2131;
  assign N292 = N2091 & N2132;
  assign N291 = N2091 & N2133;
  assign N290 = N2091 & N2134;
  assign N289 = N2091 & N2135;
  assign N288 = N2091 & N2136;
  assign N287 = N2091 & N2137;
  assign N286 = N2091 & N2138;
  assign N285 = N2091 & N2139;
  assign N284 = N2091 & N2140;
  assign N283 = N2091 & N2141;
  assign N282 = N2091 & N2142;
  assign N281 = N2091 & N2143;
  assign N280 = N2091 & N2144;
  assign N279 = N2091 & N2145;
  assign N278 = N2091 & N2146;
  assign N277 = N2091 & N2147;
  assign N276 = N2091 & N2148;
  assign N275 = N2092 & N2117;
  assign N274 = N2092 & N2118;
  assign N273 = N2092 & N2119;
  assign N272 = N2092 & N2120;
  assign N271 = N2092 & N2121;
  assign N270 = N2092 & N2122;
  assign N269 = N2092 & N2123;
  assign N268 = N2092 & N2124;
  assign N267 = N2092 & N2125;
  assign N266 = N2092 & N2126;
  assign N265 = N2092 & N2127;
  assign N264 = N2092 & N2128;
  assign N263 = N2092 & N2129;
  assign N262 = N2092 & N2130;
  assign N261 = N2092 & N2131;
  assign N260 = N2092 & N2132;
  assign N259 = N2092 & N2133;
  assign N258 = N2092 & N2134;
  assign N257 = N2092 & N2135;
  assign N256 = N2092 & N2136;
  assign N255 = N2092 & N2137;
  assign N254 = N2092 & N2138;
  assign N253 = N2092 & N2139;
  assign N252 = N2092 & N2140;
  assign N251 = N2092 & N2141;
  assign N250 = N2092 & N2142;
  assign N249 = N2092 & N2143;
  assign N248 = N2092 & N2144;
  assign N247 = N2092 & N2145;
  assign N246 = N2092 & N2146;
  assign N245 = N2092 & N2147;
  assign N244 = N2092 & N2148;
  assign N243 = N2093 & N2117;
  assign N242 = N2093 & N2118;
  assign N241 = N2093 & N2119;
  assign N240 = N2093 & N2120;
  assign N239 = N2093 & N2121;
  assign N238 = N2093 & N2122;
  assign N237 = N2093 & N2123;
  assign N236 = N2093 & N2124;
  assign N235 = N2093 & N2125;
  assign N234 = N2093 & N2126;
  assign N233 = N2093 & N2127;
  assign N232 = N2093 & N2128;
  assign N231 = N2093 & N2129;
  assign N230 = N2093 & N2130;
  assign N229 = N2093 & N2131;
  assign N228 = N2093 & N2132;
  assign N227 = N2093 & N2133;
  assign N226 = N2093 & N2134;
  assign N225 = N2093 & N2135;
  assign N224 = N2093 & N2136;
  assign N223 = N2093 & N2137;
  assign N222 = N2093 & N2138;
  assign N221 = N2093 & N2139;
  assign N220 = N2093 & N2140;
  assign N219 = N2093 & N2141;
  assign N218 = N2093 & N2142;
  assign N217 = N2093 & N2143;
  assign N216 = N2093 & N2144;
  assign N215 = N2093 & N2145;
  assign N214 = N2093 & N2146;
  assign N213 = N2093 & N2147;
  assign N212 = N2093 & N2148;
  assign N211 = N2094 & N2117;
  assign N210 = N2094 & N2118;
  assign N209 = N2094 & N2119;
  assign N208 = N2094 & N2120;
  assign N207 = N2094 & N2121;
  assign N206 = N2094 & N2122;
  assign N205 = N2094 & N2123;
  assign N204 = N2094 & N2124;
  assign N203 = N2094 & N2125;
  assign N202 = N2094 & N2126;
  assign N201 = N2094 & N2127;
  assign N200 = N2094 & N2128;
  assign N199 = N2094 & N2129;
  assign N198 = N2094 & N2130;
  assign N197 = N2094 & N2131;
  assign N196 = N2094 & N2132;
  assign N195 = N2094 & N2133;
  assign N194 = N2094 & N2134;
  assign N193 = N2094 & N2135;
  assign N192 = N2094 & N2136;
  assign N191 = N2094 & N2137;
  assign N190 = N2094 & N2138;
  assign N189 = N2094 & N2139;
  assign N188 = N2094 & N2140;
  assign N187 = N2094 & N2141;
  assign N186 = N2094 & N2142;
  assign N185 = N2094 & N2143;
  assign N184 = N2094 & N2144;
  assign N183 = N2094 & N2145;
  assign N182 = N2094 & N2146;
  assign N181 = N2094 & N2147;
  assign N180 = N2094 & N2148;
  assign N179 = N2095 & N2117;
  assign N178 = N2095 & N2118;
  assign N177 = N2095 & N2119;
  assign N176 = N2095 & N2120;
  assign N175 = N2095 & N2121;
  assign N174 = N2095 & N2122;
  assign N173 = N2095 & N2123;
  assign N172 = N2095 & N2124;
  assign N171 = N2095 & N2125;
  assign N170 = N2095 & N2126;
  assign N169 = N2095 & N2127;
  assign N168 = N2095 & N2128;
  assign N167 = N2095 & N2129;
  assign N166 = N2095 & N2130;
  assign N165 = N2095 & N2131;
  assign N164 = N2095 & N2132;
  assign N163 = N2095 & N2133;
  assign N162 = N2095 & N2134;
  assign N161 = N2095 & N2135;
  assign N160 = N2095 & N2136;
  assign N159 = N2095 & N2137;
  assign N158 = N2095 & N2138;
  assign N157 = N2095 & N2139;
  assign N156 = N2095 & N2140;
  assign N155 = N2095 & N2141;
  assign N154 = N2095 & N2142;
  assign N153 = N2095 & N2143;
  assign N152 = N2095 & N2144;
  assign N151 = N2095 & N2145;
  assign N150 = N2095 & N2146;
  assign N149 = N2095 & N2147;
  assign N148 = N2095 & N2148;
  assign N147 = N2096 & N2117;
  assign N146 = N2096 & N2118;
  assign N145 = N2096 & N2119;
  assign N144 = N2096 & N2120;
  assign N143 = N2096 & N2121;
  assign N142 = N2096 & N2122;
  assign N141 = N2096 & N2123;
  assign N140 = N2096 & N2124;
  assign N139 = N2096 & N2125;
  assign N138 = N2096 & N2126;
  assign N137 = N2096 & N2127;
  assign N136 = N2096 & N2128;
  assign N135 = N2096 & N2129;
  assign N134 = N2096 & N2130;
  assign N133 = N2096 & N2131;
  assign N132 = N2096 & N2132;
  assign N131 = N2096 & N2133;
  assign N130 = N2096 & N2134;
  assign N129 = N2096 & N2135;
  assign N128 = N2096 & N2136;
  assign N127 = N2096 & N2137;
  assign N126 = N2096 & N2138;
  assign N125 = N2096 & N2139;
  assign N124 = N2096 & N2140;
  assign N123 = N2096 & N2141;
  assign N122 = N2096 & N2142;
  assign N121 = N2096 & N2143;
  assign N120 = N2096 & N2144;
  assign N119 = N2096 & N2145;
  assign N118 = N2096 & N2146;
  assign N117 = N2096 & N2147;
  assign N116 = N2096 & N2148;
  assign N115 = N2097 & N2117;
  assign N114 = N2097 & N2118;
  assign N113 = N2097 & N2119;
  assign N112 = N2097 & N2120;
  assign N111 = N2097 & N2121;
  assign N110 = N2097 & N2122;
  assign N109 = N2097 & N2123;
  assign N108 = N2097 & N2124;
  assign N107 = N2097 & N2125;
  assign N106 = N2097 & N2126;
  assign N105 = N2097 & N2127;
  assign N104 = N2097 & N2128;
  assign N103 = N2097 & N2129;
  assign N102 = N2097 & N2130;
  assign N101 = N2097 & N2131;
  assign N100 = N2097 & N2132;
  assign N99 = N2097 & N2133;
  assign N98 = N2097 & N2134;
  assign N97 = N2097 & N2135;
  assign N96 = N2097 & N2136;
  assign N95 = N2097 & N2137;
  assign N94 = N2097 & N2138;
  assign N93 = N2097 & N2139;
  assign N92 = N2097 & N2140;
  assign N91 = N2097 & N2141;
  assign N90 = N2097 & N2142;
  assign N89 = N2097 & N2143;
  assign N88 = N2097 & N2144;
  assign N87 = N2097 & N2145;
  assign N86 = N2097 & N2146;
  assign N85 = N2097 & N2147;
  assign N84 = N2097 & N2148;
  assign N83 = N2098 & N2117;
  assign N82 = N2098 & N2118;
  assign N81 = N2098 & N2119;
  assign N80 = N2098 & N2120;
  assign N79 = N2098 & N2121;
  assign N78 = N2098 & N2122;
  assign N77 = N2098 & N2123;
  assign N76 = N2098 & N2124;
  assign N75 = N2098 & N2125;
  assign N74 = N2098 & N2126;
  assign N73 = N2098 & N2127;
  assign N72 = N2098 & N2128;
  assign N71 = N2098 & N2129;
  assign N70 = N2098 & N2130;
  assign N69 = N2098 & N2131;
  assign N68 = N2098 & N2132;
  assign N67 = N2098 & N2133;
  assign N66 = N2098 & N2134;
  assign N65 = N2098 & N2135;
  assign N64 = N2098 & N2136;
  assign N63 = N2098 & N2137;
  assign N62 = N2098 & N2138;
  assign N61 = N2098 & N2139;
  assign N60 = N2098 & N2140;
  assign N59 = N2098 & N2141;
  assign N58 = N2098 & N2142;
  assign N57 = N2098 & N2143;
  assign N56 = N2098 & N2144;
  assign N55 = N2098 & N2145;
  assign N54 = N2098 & N2146;
  assign N53 = N2098 & N2147;
  assign N52 = N2098 & N2148;
  assign N51 = N2099 & N2117;
  assign N50 = N2099 & N2118;
  assign N49 = N2099 & N2119;
  assign N48 = N2099 & N2120;
  assign N47 = N2099 & N2121;
  assign N46 = N2099 & N2122;
  assign N45 = N2099 & N2123;
  assign N44 = N2099 & N2124;
  assign N43 = N2099 & N2125;
  assign N42 = N2099 & N2126;
  assign N41 = N2099 & N2127;
  assign N40 = N2099 & N2128;
  assign N39 = N2099 & N2129;
  assign N38 = N2099 & N2130;
  assign N37 = N2099 & N2131;
  assign N36 = N2099 & N2132;
  assign N35 = N2099 & N2133;
  assign N34 = N2099 & N2134;
  assign N33 = N2099 & N2135;
  assign N32 = N2099 & N2136;
  assign N31 = N2099 & N2137;
  assign N30 = N2099 & N2138;
  assign N29 = N2099 & N2139;
  assign N28 = N2099 & N2140;
  assign N27 = N2099 & N2141;
  assign N26 = N2099 & N2142;
  assign N25 = N2099 & N2143;
  assign N24 = N2099 & N2144;
  assign N23 = N2099 & N2145;
  assign N22 = N2099 & N2146;
  assign N21 = N2099 & N2147;
  assign N20 = N2099 & N2148;
  assign { N1049, N1048, N1047, N1046, N1045, N1044, N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N542, N540, N538, N536, N534, N532 } = (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N1563)? { N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = reset_i;
  assign { N543, N541, N539, N537, N535, N533 } = (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                  (N1563)? { w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i } : 1'b0;
  assign { N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064, N1063, N1062, N1061, N1060, N1059, N1058, N1057, N1056, N1055, N1054, N1053, N1052, N1051, N1050 } = (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N1563)? { N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign r_v_o = N2149 & matched;
  assign N2149 = en_i & r_v_i;
  assign empty_v_o = en_i & empty_found;
  assign N17 = en_i & w_v_i;
  assign N18 = N17 | reset_i;
  assign N19 = ~N18;
  assign N1562 = ~reset_i;
  assign N1563 = N17 & N1562;
  assign match_array[0] = N2152 & valid[0];
  assign N2152 = N2151 & N1564;
  assign N2151 = N2150 & en_i;
  assign N2150 = ~reset_i;
  assign empty_array[0] = N2153 & N2154;
  assign N2153 = N2150 & en_i;
  assign N2154 = ~valid[0];
  assign match_array[1] = N2156 & valid[1];
  assign N2156 = N2155 & N1565;
  assign N2155 = N2150 & en_i;
  assign empty_array[1] = N2157 & N2158;
  assign N2157 = N2150 & en_i;
  assign N2158 = ~valid[1];
  assign match_array[2] = N2160 & valid[2];
  assign N2160 = N2159 & N1566;
  assign N2159 = N2150 & en_i;
  assign empty_array[2] = N2161 & N2162;
  assign N2161 = N2150 & en_i;
  assign N2162 = ~valid[2];
  assign match_array[3] = N2164 & valid[3];
  assign N2164 = N2163 & N1567;
  assign N2163 = N2150 & en_i;
  assign empty_array[3] = N2165 & N2166;
  assign N2165 = N2150 & en_i;
  assign N2166 = ~valid[3];
  assign match_array[4] = N2168 & valid[4];
  assign N2168 = N2167 & N1568;
  assign N2167 = N2150 & en_i;
  assign empty_array[4] = N2169 & N2170;
  assign N2169 = N2150 & en_i;
  assign N2170 = ~valid[4];
  assign match_array[5] = N2172 & valid[5];
  assign N2172 = N2171 & N1569;
  assign N2171 = N2150 & en_i;
  assign empty_array[5] = N2173 & N2174;
  assign N2173 = N2150 & en_i;
  assign N2174 = ~valid[5];
  assign match_array[6] = N2176 & valid[6];
  assign N2176 = N2175 & N1570;
  assign N2175 = N2150 & en_i;
  assign empty_array[6] = N2177 & N2178;
  assign N2177 = N2150 & en_i;
  assign N2178 = ~valid[6];
  assign match_array[7] = N2180 & valid[7];
  assign N2180 = N2179 & N1571;
  assign N2179 = N2150 & en_i;
  assign empty_array[7] = N2181 & N2182;
  assign N2181 = N2150 & en_i;
  assign N2182 = ~valid[7];
  assign match_array[8] = N2184 & valid[8];
  assign N2184 = N2183 & N1572;
  assign N2183 = N2150 & en_i;
  assign empty_array[8] = N2185 & N2186;
  assign N2185 = N2150 & en_i;
  assign N2186 = ~valid[8];
  assign match_array[9] = N2188 & valid[9];
  assign N2188 = N2187 & N1573;
  assign N2187 = N2150 & en_i;
  assign empty_array[9] = N2189 & N2190;
  assign N2189 = N2150 & en_i;
  assign N2190 = ~valid[9];
  assign match_array[10] = N2192 & valid[10];
  assign N2192 = N2191 & N1574;
  assign N2191 = N2150 & en_i;
  assign empty_array[10] = N2193 & N2194;
  assign N2193 = N2150 & en_i;
  assign N2194 = ~valid[10];
  assign match_array[11] = N2196 & valid[11];
  assign N2196 = N2195 & N1575;
  assign N2195 = N2150 & en_i;
  assign empty_array[11] = N2197 & N2198;
  assign N2197 = N2150 & en_i;
  assign N2198 = ~valid[11];
  assign match_array[12] = N2200 & valid[12];
  assign N2200 = N2199 & N1576;
  assign N2199 = N2150 & en_i;
  assign empty_array[12] = N2201 & N2202;
  assign N2201 = N2150 & en_i;
  assign N2202 = ~valid[12];
  assign match_array[13] = N2204 & valid[13];
  assign N2204 = N2203 & N1577;
  assign N2203 = N2150 & en_i;
  assign empty_array[13] = N2205 & N2206;
  assign N2205 = N2150 & en_i;
  assign N2206 = ~valid[13];
  assign match_array[14] = N2208 & valid[14];
  assign N2208 = N2207 & N1578;
  assign N2207 = N2150 & en_i;
  assign empty_array[14] = N2209 & N2210;
  assign N2209 = N2150 & en_i;
  assign N2210 = ~valid[14];
  assign match_array[15] = N2212 & valid[15];
  assign N2212 = N2211 & N1579;
  assign N2211 = N2150 & en_i;
  assign empty_array[15] = N2213 & N2214;
  assign N2213 = N2150 & en_i;
  assign N2214 = ~valid[15];
  assign match_array[16] = N2216 & valid[16];
  assign N2216 = N2215 & N1580;
  assign N2215 = N2150 & en_i;
  assign empty_array[16] = N2217 & N2218;
  assign N2217 = N2150 & en_i;
  assign N2218 = ~valid[16];
  assign match_array[17] = N2220 & valid[17];
  assign N2220 = N2219 & N1581;
  assign N2219 = N2150 & en_i;
  assign empty_array[17] = N2221 & N2222;
  assign N2221 = N2150 & en_i;
  assign N2222 = ~valid[17];
  assign match_array[18] = N2224 & valid[18];
  assign N2224 = N2223 & N1582;
  assign N2223 = N2150 & en_i;
  assign empty_array[18] = N2225 & N2226;
  assign N2225 = N2150 & en_i;
  assign N2226 = ~valid[18];
  assign match_array[19] = N2228 & valid[19];
  assign N2228 = N2227 & N1583;
  assign N2227 = N2150 & en_i;
  assign empty_array[19] = N2229 & N2230;
  assign N2229 = N2150 & en_i;
  assign N2230 = ~valid[19];
  assign match_array[20] = N2232 & valid[20];
  assign N2232 = N2231 & N1584;
  assign N2231 = N2150 & en_i;
  assign empty_array[20] = N2233 & N2234;
  assign N2233 = N2150 & en_i;
  assign N2234 = ~valid[20];
  assign match_array[21] = N2236 & valid[21];
  assign N2236 = N2235 & N1585;
  assign N2235 = N2150 & en_i;
  assign empty_array[21] = N2237 & N2238;
  assign N2237 = N2150 & en_i;
  assign N2238 = ~valid[21];
  assign match_array[22] = N2240 & valid[22];
  assign N2240 = N2239 & N1586;
  assign N2239 = N2150 & en_i;
  assign empty_array[22] = N2241 & N2242;
  assign N2241 = N2150 & en_i;
  assign N2242 = ~valid[22];
  assign match_array[23] = N2244 & valid[23];
  assign N2244 = N2243 & N1587;
  assign N2243 = N2150 & en_i;
  assign empty_array[23] = N2245 & N2246;
  assign N2245 = N2150 & en_i;
  assign N2246 = ~valid[23];
  assign match_array[24] = N2248 & valid[24];
  assign N2248 = N2247 & N1588;
  assign N2247 = N2150 & en_i;
  assign empty_array[24] = N2249 & N2250;
  assign N2249 = N2150 & en_i;
  assign N2250 = ~valid[24];
  assign match_array[25] = N2252 & valid[25];
  assign N2252 = N2251 & N1589;
  assign N2251 = N2150 & en_i;
  assign empty_array[25] = N2253 & N2254;
  assign N2253 = N2150 & en_i;
  assign N2254 = ~valid[25];
  assign match_array[26] = N2256 & valid[26];
  assign N2256 = N2255 & N1590;
  assign N2255 = N2150 & en_i;
  assign empty_array[26] = N2257 & N2258;
  assign N2257 = N2150 & en_i;
  assign N2258 = ~valid[26];
  assign match_array[27] = N2260 & valid[27];
  assign N2260 = N2259 & N1591;
  assign N2259 = N2150 & en_i;
  assign empty_array[27] = N2261 & N2262;
  assign N2261 = N2150 & en_i;
  assign N2262 = ~valid[27];
  assign match_array[28] = N2264 & valid[28];
  assign N2264 = N2263 & N1592;
  assign N2263 = N2150 & en_i;
  assign empty_array[28] = N2265 & N2266;
  assign N2265 = N2150 & en_i;
  assign N2266 = ~valid[28];
  assign match_array[29] = N2268 & valid[29];
  assign N2268 = N2267 & N1593;
  assign N2267 = N2150 & en_i;
  assign empty_array[29] = N2269 & N2270;
  assign N2269 = N2150 & en_i;
  assign N2270 = ~valid[29];
  assign match_array[30] = N2272 & valid[30];
  assign N2272 = N2271 & N1594;
  assign N2271 = N2150 & en_i;
  assign empty_array[30] = N2273 & N2274;
  assign N2273 = N2150 & en_i;
  assign N2274 = ~valid[30];
  assign match_array[31] = N2276 & valid[31];
  assign N2276 = N2275 & N1595;
  assign N2275 = N2150 & en_i;
  assign empty_array[31] = N2277 & N2278;
  assign N2277 = N2150 & en_i;
  assign N2278 = ~valid[31];
  assign match_array[32] = N2280 & valid[32];
  assign N2280 = N2279 & N1596;
  assign N2279 = N2150 & en_i;
  assign empty_array[32] = N2281 & N2282;
  assign N2281 = N2150 & en_i;
  assign N2282 = ~valid[32];
  assign match_array[33] = N2284 & valid[33];
  assign N2284 = N2283 & N1597;
  assign N2283 = N2150 & en_i;
  assign empty_array[33] = N2285 & N2286;
  assign N2285 = N2150 & en_i;
  assign N2286 = ~valid[33];
  assign match_array[34] = N2288 & valid[34];
  assign N2288 = N2287 & N1598;
  assign N2287 = N2150 & en_i;
  assign empty_array[34] = N2289 & N2290;
  assign N2289 = N2150 & en_i;
  assign N2290 = ~valid[34];
  assign match_array[35] = N2292 & valid[35];
  assign N2292 = N2291 & N1599;
  assign N2291 = N2150 & en_i;
  assign empty_array[35] = N2293 & N2294;
  assign N2293 = N2150 & en_i;
  assign N2294 = ~valid[35];
  assign match_array[36] = N2296 & valid[36];
  assign N2296 = N2295 & N1600;
  assign N2295 = N2150 & en_i;
  assign empty_array[36] = N2297 & N2298;
  assign N2297 = N2150 & en_i;
  assign N2298 = ~valid[36];
  assign match_array[37] = N2300 & valid[37];
  assign N2300 = N2299 & N1601;
  assign N2299 = N2150 & en_i;
  assign empty_array[37] = N2301 & N2302;
  assign N2301 = N2150 & en_i;
  assign N2302 = ~valid[37];
  assign match_array[38] = N2304 & valid[38];
  assign N2304 = N2303 & N1602;
  assign N2303 = N2150 & en_i;
  assign empty_array[38] = N2305 & N2306;
  assign N2305 = N2150 & en_i;
  assign N2306 = ~valid[38];
  assign match_array[39] = N2308 & valid[39];
  assign N2308 = N2307 & N1603;
  assign N2307 = N2150 & en_i;
  assign empty_array[39] = N2309 & N2310;
  assign N2309 = N2150 & en_i;
  assign N2310 = ~valid[39];
  assign match_array[40] = N2312 & valid[40];
  assign N2312 = N2311 & N1604;
  assign N2311 = N2150 & en_i;
  assign empty_array[40] = N2313 & N2314;
  assign N2313 = N2150 & en_i;
  assign N2314 = ~valid[40];
  assign match_array[41] = N2316 & valid[41];
  assign N2316 = N2315 & N1605;
  assign N2315 = N2150 & en_i;
  assign empty_array[41] = N2317 & N2318;
  assign N2317 = N2150 & en_i;
  assign N2318 = ~valid[41];
  assign match_array[42] = N2320 & valid[42];
  assign N2320 = N2319 & N1606;
  assign N2319 = N2150 & en_i;
  assign empty_array[42] = N2321 & N2322;
  assign N2321 = N2150 & en_i;
  assign N2322 = ~valid[42];
  assign match_array[43] = N2324 & valid[43];
  assign N2324 = N2323 & N1607;
  assign N2323 = N2150 & en_i;
  assign empty_array[43] = N2325 & N2326;
  assign N2325 = N2150 & en_i;
  assign N2326 = ~valid[43];
  assign match_array[44] = N2328 & valid[44];
  assign N2328 = N2327 & N1608;
  assign N2327 = N2150 & en_i;
  assign empty_array[44] = N2329 & N2330;
  assign N2329 = N2150 & en_i;
  assign N2330 = ~valid[44];
  assign match_array[45] = N2332 & valid[45];
  assign N2332 = N2331 & N1609;
  assign N2331 = N2150 & en_i;
  assign empty_array[45] = N2333 & N2334;
  assign N2333 = N2150 & en_i;
  assign N2334 = ~valid[45];
  assign match_array[46] = N2336 & valid[46];
  assign N2336 = N2335 & N1610;
  assign N2335 = N2150 & en_i;
  assign empty_array[46] = N2337 & N2338;
  assign N2337 = N2150 & en_i;
  assign N2338 = ~valid[46];
  assign match_array[47] = N2340 & valid[47];
  assign N2340 = N2339 & N1611;
  assign N2339 = N2150 & en_i;
  assign empty_array[47] = N2341 & N2342;
  assign N2341 = N2150 & en_i;
  assign N2342 = ~valid[47];
  assign match_array[48] = N2344 & valid[48];
  assign N2344 = N2343 & N1612;
  assign N2343 = N2150 & en_i;
  assign empty_array[48] = N2345 & N2346;
  assign N2345 = N2150 & en_i;
  assign N2346 = ~valid[48];
  assign match_array[49] = N2348 & valid[49];
  assign N2348 = N2347 & N1613;
  assign N2347 = N2150 & en_i;
  assign empty_array[49] = N2349 & N2350;
  assign N2349 = N2150 & en_i;
  assign N2350 = ~valid[49];
  assign match_array[50] = N2352 & valid[50];
  assign N2352 = N2351 & N1614;
  assign N2351 = N2150 & en_i;
  assign empty_array[50] = N2353 & N2354;
  assign N2353 = N2150 & en_i;
  assign N2354 = ~valid[50];
  assign match_array[51] = N2356 & valid[51];
  assign N2356 = N2355 & N1615;
  assign N2355 = N2150 & en_i;
  assign empty_array[51] = N2357 & N2358;
  assign N2357 = N2150 & en_i;
  assign N2358 = ~valid[51];
  assign match_array[52] = N2360 & valid[52];
  assign N2360 = N2359 & N1616;
  assign N2359 = N2150 & en_i;
  assign empty_array[52] = N2361 & N2362;
  assign N2361 = N2150 & en_i;
  assign N2362 = ~valid[52];
  assign match_array[53] = N2364 & valid[53];
  assign N2364 = N2363 & N1617;
  assign N2363 = N2150 & en_i;
  assign empty_array[53] = N2365 & N2366;
  assign N2365 = N2150 & en_i;
  assign N2366 = ~valid[53];
  assign match_array[54] = N2368 & valid[54];
  assign N2368 = N2367 & N1618;
  assign N2367 = N2150 & en_i;
  assign empty_array[54] = N2369 & N2370;
  assign N2369 = N2150 & en_i;
  assign N2370 = ~valid[54];
  assign match_array[55] = N2372 & valid[55];
  assign N2372 = N2371 & N1619;
  assign N2371 = N2150 & en_i;
  assign empty_array[55] = N2373 & N2374;
  assign N2373 = N2150 & en_i;
  assign N2374 = ~valid[55];
  assign match_array[56] = N2376 & valid[56];
  assign N2376 = N2375 & N1620;
  assign N2375 = N2150 & en_i;
  assign empty_array[56] = N2377 & N2378;
  assign N2377 = N2150 & en_i;
  assign N2378 = ~valid[56];
  assign match_array[57] = N2380 & valid[57];
  assign N2380 = N2379 & N1621;
  assign N2379 = N2150 & en_i;
  assign empty_array[57] = N2381 & N2382;
  assign N2381 = N2150 & en_i;
  assign N2382 = ~valid[57];
  assign match_array[58] = N2384 & valid[58];
  assign N2384 = N2383 & N1622;
  assign N2383 = N2150 & en_i;
  assign empty_array[58] = N2385 & N2386;
  assign N2385 = N2150 & en_i;
  assign N2386 = ~valid[58];
  assign match_array[59] = N2388 & valid[59];
  assign N2388 = N2387 & N1623;
  assign N2387 = N2150 & en_i;
  assign empty_array[59] = N2389 & N2390;
  assign N2389 = N2150 & en_i;
  assign N2390 = ~valid[59];
  assign match_array[60] = N2392 & valid[60];
  assign N2392 = N2391 & N1624;
  assign N2391 = N2150 & en_i;
  assign empty_array[60] = N2393 & N2394;
  assign N2393 = N2150 & en_i;
  assign N2394 = ~valid[60];
  assign match_array[61] = N2396 & valid[61];
  assign N2396 = N2395 & N1625;
  assign N2395 = N2150 & en_i;
  assign empty_array[61] = N2397 & N2398;
  assign N2397 = N2150 & en_i;
  assign N2398 = ~valid[61];
  assign match_array[62] = N2400 & valid[62];
  assign N2400 = N2399 & N1626;
  assign N2399 = N2150 & en_i;
  assign empty_array[62] = N2401 & N2402;
  assign N2401 = N2150 & en_i;
  assign N2402 = ~valid[62];
  assign match_array[63] = N2404 & valid[63];
  assign N2404 = N2403 & N1627;
  assign N2403 = N2150 & en_i;
  assign empty_array[63] = N2405 & N2406;
  assign N2405 = N2150 & en_i;
  assign N2406 = ~valid[63];
  assign match_array[64] = N2408 & valid[64];
  assign N2408 = N2407 & N1628;
  assign N2407 = N2150 & en_i;
  assign empty_array[64] = N2409 & N2410;
  assign N2409 = N2150 & en_i;
  assign N2410 = ~valid[64];
  assign match_array[65] = N2412 & valid[65];
  assign N2412 = N2411 & N1629;
  assign N2411 = N2150 & en_i;
  assign empty_array[65] = N2413 & N2414;
  assign N2413 = N2150 & en_i;
  assign N2414 = ~valid[65];
  assign match_array[66] = N2416 & valid[66];
  assign N2416 = N2415 & N1630;
  assign N2415 = N2150 & en_i;
  assign empty_array[66] = N2417 & N2418;
  assign N2417 = N2150 & en_i;
  assign N2418 = ~valid[66];
  assign match_array[67] = N2420 & valid[67];
  assign N2420 = N2419 & N1631;
  assign N2419 = N2150 & en_i;
  assign empty_array[67] = N2421 & N2422;
  assign N2421 = N2150 & en_i;
  assign N2422 = ~valid[67];
  assign match_array[68] = N2424 & valid[68];
  assign N2424 = N2423 & N1632;
  assign N2423 = N2150 & en_i;
  assign empty_array[68] = N2425 & N2426;
  assign N2425 = N2150 & en_i;
  assign N2426 = ~valid[68];
  assign match_array[69] = N2428 & valid[69];
  assign N2428 = N2427 & N1633;
  assign N2427 = N2150 & en_i;
  assign empty_array[69] = N2429 & N2430;
  assign N2429 = N2150 & en_i;
  assign N2430 = ~valid[69];
  assign match_array[70] = N2432 & valid[70];
  assign N2432 = N2431 & N1634;
  assign N2431 = N2150 & en_i;
  assign empty_array[70] = N2433 & N2434;
  assign N2433 = N2150 & en_i;
  assign N2434 = ~valid[70];
  assign match_array[71] = N2436 & valid[71];
  assign N2436 = N2435 & N1635;
  assign N2435 = N2150 & en_i;
  assign empty_array[71] = N2437 & N2438;
  assign N2437 = N2150 & en_i;
  assign N2438 = ~valid[71];
  assign match_array[72] = N2440 & valid[72];
  assign N2440 = N2439 & N1636;
  assign N2439 = N2150 & en_i;
  assign empty_array[72] = N2441 & N2442;
  assign N2441 = N2150 & en_i;
  assign N2442 = ~valid[72];
  assign match_array[73] = N2444 & valid[73];
  assign N2444 = N2443 & N1637;
  assign N2443 = N2150 & en_i;
  assign empty_array[73] = N2445 & N2446;
  assign N2445 = N2150 & en_i;
  assign N2446 = ~valid[73];
  assign match_array[74] = N2448 & valid[74];
  assign N2448 = N2447 & N1638;
  assign N2447 = N2150 & en_i;
  assign empty_array[74] = N2449 & N2450;
  assign N2449 = N2150 & en_i;
  assign N2450 = ~valid[74];
  assign match_array[75] = N2452 & valid[75];
  assign N2452 = N2451 & N1639;
  assign N2451 = N2150 & en_i;
  assign empty_array[75] = N2453 & N2454;
  assign N2453 = N2150 & en_i;
  assign N2454 = ~valid[75];
  assign match_array[76] = N2456 & valid[76];
  assign N2456 = N2455 & N1640;
  assign N2455 = N2150 & en_i;
  assign empty_array[76] = N2457 & N2458;
  assign N2457 = N2150 & en_i;
  assign N2458 = ~valid[76];
  assign match_array[77] = N2460 & valid[77];
  assign N2460 = N2459 & N1641;
  assign N2459 = N2150 & en_i;
  assign empty_array[77] = N2461 & N2462;
  assign N2461 = N2150 & en_i;
  assign N2462 = ~valid[77];
  assign match_array[78] = N2464 & valid[78];
  assign N2464 = N2463 & N1642;
  assign N2463 = N2150 & en_i;
  assign empty_array[78] = N2465 & N2466;
  assign N2465 = N2150 & en_i;
  assign N2466 = ~valid[78];
  assign match_array[79] = N2468 & valid[79];
  assign N2468 = N2467 & N1643;
  assign N2467 = N2150 & en_i;
  assign empty_array[79] = N2469 & N2470;
  assign N2469 = N2150 & en_i;
  assign N2470 = ~valid[79];
  assign match_array[80] = N2472 & valid[80];
  assign N2472 = N2471 & N1644;
  assign N2471 = N2150 & en_i;
  assign empty_array[80] = N2473 & N2474;
  assign N2473 = N2150 & en_i;
  assign N2474 = ~valid[80];
  assign match_array[81] = N2476 & valid[81];
  assign N2476 = N2475 & N1645;
  assign N2475 = N2150 & en_i;
  assign empty_array[81] = N2477 & N2478;
  assign N2477 = N2150 & en_i;
  assign N2478 = ~valid[81];
  assign match_array[82] = N2480 & valid[82];
  assign N2480 = N2479 & N1646;
  assign N2479 = N2150 & en_i;
  assign empty_array[82] = N2481 & N2482;
  assign N2481 = N2150 & en_i;
  assign N2482 = ~valid[82];
  assign match_array[83] = N2484 & valid[83];
  assign N2484 = N2483 & N1647;
  assign N2483 = N2150 & en_i;
  assign empty_array[83] = N2485 & N2486;
  assign N2485 = N2150 & en_i;
  assign N2486 = ~valid[83];
  assign match_array[84] = N2488 & valid[84];
  assign N2488 = N2487 & N1648;
  assign N2487 = N2150 & en_i;
  assign empty_array[84] = N2489 & N2490;
  assign N2489 = N2150 & en_i;
  assign N2490 = ~valid[84];
  assign match_array[85] = N2492 & valid[85];
  assign N2492 = N2491 & N1649;
  assign N2491 = N2150 & en_i;
  assign empty_array[85] = N2493 & N2494;
  assign N2493 = N2150 & en_i;
  assign N2494 = ~valid[85];
  assign match_array[86] = N2496 & valid[86];
  assign N2496 = N2495 & N1650;
  assign N2495 = N2150 & en_i;
  assign empty_array[86] = N2497 & N2498;
  assign N2497 = N2150 & en_i;
  assign N2498 = ~valid[86];
  assign match_array[87] = N2500 & valid[87];
  assign N2500 = N2499 & N1651;
  assign N2499 = N2150 & en_i;
  assign empty_array[87] = N2501 & N2502;
  assign N2501 = N2150 & en_i;
  assign N2502 = ~valid[87];
  assign match_array[88] = N2504 & valid[88];
  assign N2504 = N2503 & N1652;
  assign N2503 = N2150 & en_i;
  assign empty_array[88] = N2505 & N2506;
  assign N2505 = N2150 & en_i;
  assign N2506 = ~valid[88];
  assign match_array[89] = N2508 & valid[89];
  assign N2508 = N2507 & N1653;
  assign N2507 = N2150 & en_i;
  assign empty_array[89] = N2509 & N2510;
  assign N2509 = N2150 & en_i;
  assign N2510 = ~valid[89];
  assign match_array[90] = N2512 & valid[90];
  assign N2512 = N2511 & N1654;
  assign N2511 = N2150 & en_i;
  assign empty_array[90] = N2513 & N2514;
  assign N2513 = N2150 & en_i;
  assign N2514 = ~valid[90];
  assign match_array[91] = N2516 & valid[91];
  assign N2516 = N2515 & N1655;
  assign N2515 = N2150 & en_i;
  assign empty_array[91] = N2517 & N2518;
  assign N2517 = N2150 & en_i;
  assign N2518 = ~valid[91];
  assign match_array[92] = N2520 & valid[92];
  assign N2520 = N2519 & N1656;
  assign N2519 = N2150 & en_i;
  assign empty_array[92] = N2521 & N2522;
  assign N2521 = N2150 & en_i;
  assign N2522 = ~valid[92];
  assign match_array[93] = N2524 & valid[93];
  assign N2524 = N2523 & N1657;
  assign N2523 = N2150 & en_i;
  assign empty_array[93] = N2525 & N2526;
  assign N2525 = N2150 & en_i;
  assign N2526 = ~valid[93];
  assign match_array[94] = N2528 & valid[94];
  assign N2528 = N2527 & N1658;
  assign N2527 = N2150 & en_i;
  assign empty_array[94] = N2529 & N2530;
  assign N2529 = N2150 & en_i;
  assign N2530 = ~valid[94];
  assign match_array[95] = N2532 & valid[95];
  assign N2532 = N2531 & N1659;
  assign N2531 = N2150 & en_i;
  assign empty_array[95] = N2533 & N2534;
  assign N2533 = N2150 & en_i;
  assign N2534 = ~valid[95];
  assign match_array[96] = N2536 & valid[96];
  assign N2536 = N2535 & N1660;
  assign N2535 = N2150 & en_i;
  assign empty_array[96] = N2537 & N2538;
  assign N2537 = N2150 & en_i;
  assign N2538 = ~valid[96];
  assign match_array[97] = N2540 & valid[97];
  assign N2540 = N2539 & N1661;
  assign N2539 = N2150 & en_i;
  assign empty_array[97] = N2541 & N2542;
  assign N2541 = N2150 & en_i;
  assign N2542 = ~valid[97];
  assign match_array[98] = N2544 & valid[98];
  assign N2544 = N2543 & N1662;
  assign N2543 = N2150 & en_i;
  assign empty_array[98] = N2545 & N2546;
  assign N2545 = N2150 & en_i;
  assign N2546 = ~valid[98];
  assign match_array[99] = N2548 & valid[99];
  assign N2548 = N2547 & N1663;
  assign N2547 = N2150 & en_i;
  assign empty_array[99] = N2549 & N2550;
  assign N2549 = N2150 & en_i;
  assign N2550 = ~valid[99];
  assign match_array[100] = N2552 & valid[100];
  assign N2552 = N2551 & N1664;
  assign N2551 = N2150 & en_i;
  assign empty_array[100] = N2553 & N2554;
  assign N2553 = N2150 & en_i;
  assign N2554 = ~valid[100];
  assign match_array[101] = N2556 & valid[101];
  assign N2556 = N2555 & N1665;
  assign N2555 = N2150 & en_i;
  assign empty_array[101] = N2557 & N2558;
  assign N2557 = N2150 & en_i;
  assign N2558 = ~valid[101];
  assign match_array[102] = N2560 & valid[102];
  assign N2560 = N2559 & N1666;
  assign N2559 = N2150 & en_i;
  assign empty_array[102] = N2561 & N2562;
  assign N2561 = N2150 & en_i;
  assign N2562 = ~valid[102];
  assign match_array[103] = N2564 & valid[103];
  assign N2564 = N2563 & N1667;
  assign N2563 = N2150 & en_i;
  assign empty_array[103] = N2565 & N2566;
  assign N2565 = N2150 & en_i;
  assign N2566 = ~valid[103];
  assign match_array[104] = N2568 & valid[104];
  assign N2568 = N2567 & N1668;
  assign N2567 = N2150 & en_i;
  assign empty_array[104] = N2569 & N2570;
  assign N2569 = N2150 & en_i;
  assign N2570 = ~valid[104];
  assign match_array[105] = N2572 & valid[105];
  assign N2572 = N2571 & N1669;
  assign N2571 = N2150 & en_i;
  assign empty_array[105] = N2573 & N2574;
  assign N2573 = N2150 & en_i;
  assign N2574 = ~valid[105];
  assign match_array[106] = N2576 & valid[106];
  assign N2576 = N2575 & N1670;
  assign N2575 = N2150 & en_i;
  assign empty_array[106] = N2577 & N2578;
  assign N2577 = N2150 & en_i;
  assign N2578 = ~valid[106];
  assign match_array[107] = N2580 & valid[107];
  assign N2580 = N2579 & N1671;
  assign N2579 = N2150 & en_i;
  assign empty_array[107] = N2581 & N2582;
  assign N2581 = N2150 & en_i;
  assign N2582 = ~valid[107];
  assign match_array[108] = N2584 & valid[108];
  assign N2584 = N2583 & N1672;
  assign N2583 = N2150 & en_i;
  assign empty_array[108] = N2585 & N2586;
  assign N2585 = N2150 & en_i;
  assign N2586 = ~valid[108];
  assign match_array[109] = N2588 & valid[109];
  assign N2588 = N2587 & N1673;
  assign N2587 = N2150 & en_i;
  assign empty_array[109] = N2589 & N2590;
  assign N2589 = N2150 & en_i;
  assign N2590 = ~valid[109];
  assign match_array[110] = N2592 & valid[110];
  assign N2592 = N2591 & N1674;
  assign N2591 = N2150 & en_i;
  assign empty_array[110] = N2593 & N2594;
  assign N2593 = N2150 & en_i;
  assign N2594 = ~valid[110];
  assign match_array[111] = N2596 & valid[111];
  assign N2596 = N2595 & N1675;
  assign N2595 = N2150 & en_i;
  assign empty_array[111] = N2597 & N2598;
  assign N2597 = N2150 & en_i;
  assign N2598 = ~valid[111];
  assign match_array[112] = N2600 & valid[112];
  assign N2600 = N2599 & N1676;
  assign N2599 = N2150 & en_i;
  assign empty_array[112] = N2601 & N2602;
  assign N2601 = N2150 & en_i;
  assign N2602 = ~valid[112];
  assign match_array[113] = N2604 & valid[113];
  assign N2604 = N2603 & N1677;
  assign N2603 = N2150 & en_i;
  assign empty_array[113] = N2605 & N2606;
  assign N2605 = N2150 & en_i;
  assign N2606 = ~valid[113];
  assign match_array[114] = N2608 & valid[114];
  assign N2608 = N2607 & N1678;
  assign N2607 = N2150 & en_i;
  assign empty_array[114] = N2609 & N2610;
  assign N2609 = N2150 & en_i;
  assign N2610 = ~valid[114];
  assign match_array[115] = N2612 & valid[115];
  assign N2612 = N2611 & N1679;
  assign N2611 = N2150 & en_i;
  assign empty_array[115] = N2613 & N2614;
  assign N2613 = N2150 & en_i;
  assign N2614 = ~valid[115];
  assign match_array[116] = N2616 & valid[116];
  assign N2616 = N2615 & N1680;
  assign N2615 = N2150 & en_i;
  assign empty_array[116] = N2617 & N2618;
  assign N2617 = N2150 & en_i;
  assign N2618 = ~valid[116];
  assign match_array[117] = N2620 & valid[117];
  assign N2620 = N2619 & N1681;
  assign N2619 = N2150 & en_i;
  assign empty_array[117] = N2621 & N2622;
  assign N2621 = N2150 & en_i;
  assign N2622 = ~valid[117];
  assign match_array[118] = N2624 & valid[118];
  assign N2624 = N2623 & N1682;
  assign N2623 = N2150 & en_i;
  assign empty_array[118] = N2625 & N2626;
  assign N2625 = N2150 & en_i;
  assign N2626 = ~valid[118];
  assign match_array[119] = N2628 & valid[119];
  assign N2628 = N2627 & N1683;
  assign N2627 = N2150 & en_i;
  assign empty_array[119] = N2629 & N2630;
  assign N2629 = N2150 & en_i;
  assign N2630 = ~valid[119];
  assign match_array[120] = N2632 & valid[120];
  assign N2632 = N2631 & N1684;
  assign N2631 = N2150 & en_i;
  assign empty_array[120] = N2633 & N2634;
  assign N2633 = N2150 & en_i;
  assign N2634 = ~valid[120];
  assign match_array[121] = N2636 & valid[121];
  assign N2636 = N2635 & N1685;
  assign N2635 = N2150 & en_i;
  assign empty_array[121] = N2637 & N2638;
  assign N2637 = N2150 & en_i;
  assign N2638 = ~valid[121];
  assign match_array[122] = N2640 & valid[122];
  assign N2640 = N2639 & N1686;
  assign N2639 = N2150 & en_i;
  assign empty_array[122] = N2641 & N2642;
  assign N2641 = N2150 & en_i;
  assign N2642 = ~valid[122];
  assign match_array[123] = N2644 & valid[123];
  assign N2644 = N2643 & N1687;
  assign N2643 = N2150 & en_i;
  assign empty_array[123] = N2645 & N2646;
  assign N2645 = N2150 & en_i;
  assign N2646 = ~valid[123];
  assign match_array[124] = N2648 & valid[124];
  assign N2648 = N2647 & N1688;
  assign N2647 = N2150 & en_i;
  assign empty_array[124] = N2649 & N2650;
  assign N2649 = N2150 & en_i;
  assign N2650 = ~valid[124];
  assign match_array[125] = N2652 & valid[125];
  assign N2652 = N2651 & N1689;
  assign N2651 = N2150 & en_i;
  assign empty_array[125] = N2653 & N2654;
  assign N2653 = N2150 & en_i;
  assign N2654 = ~valid[125];
  assign match_array[126] = N2656 & valid[126];
  assign N2656 = N2655 & N1690;
  assign N2655 = N2150 & en_i;
  assign empty_array[126] = N2657 & N2658;
  assign N2657 = N2150 & en_i;
  assign N2658 = ~valid[126];
  assign match_array[127] = N2660 & valid[127];
  assign N2660 = N2659 & N1691;
  assign N2659 = N2150 & en_i;
  assign empty_array[127] = N2661 & N2662;
  assign N2661 = N2150 & en_i;
  assign N2662 = ~valid[127];
  assign match_array[128] = N2664 & valid[128];
  assign N2664 = N2663 & N1692;
  assign N2663 = N2150 & en_i;
  assign empty_array[128] = N2665 & N2666;
  assign N2665 = N2150 & en_i;
  assign N2666 = ~valid[128];
  assign match_array[129] = N2668 & valid[129];
  assign N2668 = N2667 & N1693;
  assign N2667 = N2150 & en_i;
  assign empty_array[129] = N2669 & N2670;
  assign N2669 = N2150 & en_i;
  assign N2670 = ~valid[129];
  assign match_array[130] = N2672 & valid[130];
  assign N2672 = N2671 & N1694;
  assign N2671 = N2150 & en_i;
  assign empty_array[130] = N2673 & N2674;
  assign N2673 = N2150 & en_i;
  assign N2674 = ~valid[130];
  assign match_array[131] = N2676 & valid[131];
  assign N2676 = N2675 & N1695;
  assign N2675 = N2150 & en_i;
  assign empty_array[131] = N2677 & N2678;
  assign N2677 = N2150 & en_i;
  assign N2678 = ~valid[131];
  assign match_array[132] = N2680 & valid[132];
  assign N2680 = N2679 & N1696;
  assign N2679 = N2150 & en_i;
  assign empty_array[132] = N2681 & N2682;
  assign N2681 = N2150 & en_i;
  assign N2682 = ~valid[132];
  assign match_array[133] = N2684 & valid[133];
  assign N2684 = N2683 & N1697;
  assign N2683 = N2150 & en_i;
  assign empty_array[133] = N2685 & N2686;
  assign N2685 = N2150 & en_i;
  assign N2686 = ~valid[133];
  assign match_array[134] = N2688 & valid[134];
  assign N2688 = N2687 & N1698;
  assign N2687 = N2150 & en_i;
  assign empty_array[134] = N2689 & N2690;
  assign N2689 = N2150 & en_i;
  assign N2690 = ~valid[134];
  assign match_array[135] = N2692 & valid[135];
  assign N2692 = N2691 & N1699;
  assign N2691 = N2150 & en_i;
  assign empty_array[135] = N2693 & N2694;
  assign N2693 = N2150 & en_i;
  assign N2694 = ~valid[135];
  assign match_array[136] = N2696 & valid[136];
  assign N2696 = N2695 & N1700;
  assign N2695 = N2150 & en_i;
  assign empty_array[136] = N2697 & N2698;
  assign N2697 = N2150 & en_i;
  assign N2698 = ~valid[136];
  assign match_array[137] = N2700 & valid[137];
  assign N2700 = N2699 & N1701;
  assign N2699 = N2150 & en_i;
  assign empty_array[137] = N2701 & N2702;
  assign N2701 = N2150 & en_i;
  assign N2702 = ~valid[137];
  assign match_array[138] = N2704 & valid[138];
  assign N2704 = N2703 & N1702;
  assign N2703 = N2150 & en_i;
  assign empty_array[138] = N2705 & N2706;
  assign N2705 = N2150 & en_i;
  assign N2706 = ~valid[138];
  assign match_array[139] = N2708 & valid[139];
  assign N2708 = N2707 & N1703;
  assign N2707 = N2150 & en_i;
  assign empty_array[139] = N2709 & N2710;
  assign N2709 = N2150 & en_i;
  assign N2710 = ~valid[139];
  assign match_array[140] = N2712 & valid[140];
  assign N2712 = N2711 & N1704;
  assign N2711 = N2150 & en_i;
  assign empty_array[140] = N2713 & N2714;
  assign N2713 = N2150 & en_i;
  assign N2714 = ~valid[140];
  assign match_array[141] = N2716 & valid[141];
  assign N2716 = N2715 & N1705;
  assign N2715 = N2150 & en_i;
  assign empty_array[141] = N2717 & N2718;
  assign N2717 = N2150 & en_i;
  assign N2718 = ~valid[141];
  assign match_array[142] = N2720 & valid[142];
  assign N2720 = N2719 & N1706;
  assign N2719 = N2150 & en_i;
  assign empty_array[142] = N2721 & N2722;
  assign N2721 = N2150 & en_i;
  assign N2722 = ~valid[142];
  assign match_array[143] = N2724 & valid[143];
  assign N2724 = N2723 & N1707;
  assign N2723 = N2150 & en_i;
  assign empty_array[143] = N2725 & N2726;
  assign N2725 = N2150 & en_i;
  assign N2726 = ~valid[143];
  assign match_array[144] = N2728 & valid[144];
  assign N2728 = N2727 & N1708;
  assign N2727 = N2150 & en_i;
  assign empty_array[144] = N2729 & N2730;
  assign N2729 = N2150 & en_i;
  assign N2730 = ~valid[144];
  assign match_array[145] = N2732 & valid[145];
  assign N2732 = N2731 & N1709;
  assign N2731 = N2150 & en_i;
  assign empty_array[145] = N2733 & N2734;
  assign N2733 = N2150 & en_i;
  assign N2734 = ~valid[145];
  assign match_array[146] = N2736 & valid[146];
  assign N2736 = N2735 & N1710;
  assign N2735 = N2150 & en_i;
  assign empty_array[146] = N2737 & N2738;
  assign N2737 = N2150 & en_i;
  assign N2738 = ~valid[146];
  assign match_array[147] = N2740 & valid[147];
  assign N2740 = N2739 & N1711;
  assign N2739 = N2150 & en_i;
  assign empty_array[147] = N2741 & N2742;
  assign N2741 = N2150 & en_i;
  assign N2742 = ~valid[147];
  assign match_array[148] = N2744 & valid[148];
  assign N2744 = N2743 & N1712;
  assign N2743 = N2150 & en_i;
  assign empty_array[148] = N2745 & N2746;
  assign N2745 = N2150 & en_i;
  assign N2746 = ~valid[148];
  assign match_array[149] = N2748 & valid[149];
  assign N2748 = N2747 & N1713;
  assign N2747 = N2150 & en_i;
  assign empty_array[149] = N2749 & N2750;
  assign N2749 = N2150 & en_i;
  assign N2750 = ~valid[149];
  assign match_array[150] = N2752 & valid[150];
  assign N2752 = N2751 & N1714;
  assign N2751 = N2150 & en_i;
  assign empty_array[150] = N2753 & N2754;
  assign N2753 = N2150 & en_i;
  assign N2754 = ~valid[150];
  assign match_array[151] = N2756 & valid[151];
  assign N2756 = N2755 & N1715;
  assign N2755 = N2150 & en_i;
  assign empty_array[151] = N2757 & N2758;
  assign N2757 = N2150 & en_i;
  assign N2758 = ~valid[151];
  assign match_array[152] = N2760 & valid[152];
  assign N2760 = N2759 & N1716;
  assign N2759 = N2150 & en_i;
  assign empty_array[152] = N2761 & N2762;
  assign N2761 = N2150 & en_i;
  assign N2762 = ~valid[152];
  assign match_array[153] = N2764 & valid[153];
  assign N2764 = N2763 & N1717;
  assign N2763 = N2150 & en_i;
  assign empty_array[153] = N2765 & N2766;
  assign N2765 = N2150 & en_i;
  assign N2766 = ~valid[153];
  assign match_array[154] = N2768 & valid[154];
  assign N2768 = N2767 & N1718;
  assign N2767 = N2150 & en_i;
  assign empty_array[154] = N2769 & N2770;
  assign N2769 = N2150 & en_i;
  assign N2770 = ~valid[154];
  assign match_array[155] = N2772 & valid[155];
  assign N2772 = N2771 & N1719;
  assign N2771 = N2150 & en_i;
  assign empty_array[155] = N2773 & N2774;
  assign N2773 = N2150 & en_i;
  assign N2774 = ~valid[155];
  assign match_array[156] = N2776 & valid[156];
  assign N2776 = N2775 & N1720;
  assign N2775 = N2150 & en_i;
  assign empty_array[156] = N2777 & N2778;
  assign N2777 = N2150 & en_i;
  assign N2778 = ~valid[156];
  assign match_array[157] = N2780 & valid[157];
  assign N2780 = N2779 & N1721;
  assign N2779 = N2150 & en_i;
  assign empty_array[157] = N2781 & N2782;
  assign N2781 = N2150 & en_i;
  assign N2782 = ~valid[157];
  assign match_array[158] = N2784 & valid[158];
  assign N2784 = N2783 & N1722;
  assign N2783 = N2150 & en_i;
  assign empty_array[158] = N2785 & N2786;
  assign N2785 = N2150 & en_i;
  assign N2786 = ~valid[158];
  assign match_array[159] = N2788 & valid[159];
  assign N2788 = N2787 & N1723;
  assign N2787 = N2150 & en_i;
  assign empty_array[159] = N2789 & N2790;
  assign N2789 = N2150 & en_i;
  assign N2790 = ~valid[159];
  assign match_array[160] = N2792 & valid[160];
  assign N2792 = N2791 & N1724;
  assign N2791 = N2150 & en_i;
  assign empty_array[160] = N2793 & N2794;
  assign N2793 = N2150 & en_i;
  assign N2794 = ~valid[160];
  assign match_array[161] = N2796 & valid[161];
  assign N2796 = N2795 & N1725;
  assign N2795 = N2150 & en_i;
  assign empty_array[161] = N2797 & N2798;
  assign N2797 = N2150 & en_i;
  assign N2798 = ~valid[161];
  assign match_array[162] = N2800 & valid[162];
  assign N2800 = N2799 & N1726;
  assign N2799 = N2150 & en_i;
  assign empty_array[162] = N2801 & N2802;
  assign N2801 = N2150 & en_i;
  assign N2802 = ~valid[162];
  assign match_array[163] = N2804 & valid[163];
  assign N2804 = N2803 & N1727;
  assign N2803 = N2150 & en_i;
  assign empty_array[163] = N2805 & N2806;
  assign N2805 = N2150 & en_i;
  assign N2806 = ~valid[163];
  assign match_array[164] = N2808 & valid[164];
  assign N2808 = N2807 & N1728;
  assign N2807 = N2150 & en_i;
  assign empty_array[164] = N2809 & N2810;
  assign N2809 = N2150 & en_i;
  assign N2810 = ~valid[164];
  assign match_array[165] = N2812 & valid[165];
  assign N2812 = N2811 & N1729;
  assign N2811 = N2150 & en_i;
  assign empty_array[165] = N2813 & N2814;
  assign N2813 = N2150 & en_i;
  assign N2814 = ~valid[165];
  assign match_array[166] = N2816 & valid[166];
  assign N2816 = N2815 & N1730;
  assign N2815 = N2150 & en_i;
  assign empty_array[166] = N2817 & N2818;
  assign N2817 = N2150 & en_i;
  assign N2818 = ~valid[166];
  assign match_array[167] = N2820 & valid[167];
  assign N2820 = N2819 & N1731;
  assign N2819 = N2150 & en_i;
  assign empty_array[167] = N2821 & N2822;
  assign N2821 = N2150 & en_i;
  assign N2822 = ~valid[167];
  assign match_array[168] = N2824 & valid[168];
  assign N2824 = N2823 & N1732;
  assign N2823 = N2150 & en_i;
  assign empty_array[168] = N2825 & N2826;
  assign N2825 = N2150 & en_i;
  assign N2826 = ~valid[168];
  assign match_array[169] = N2828 & valid[169];
  assign N2828 = N2827 & N1733;
  assign N2827 = N2150 & en_i;
  assign empty_array[169] = N2829 & N2830;
  assign N2829 = N2150 & en_i;
  assign N2830 = ~valid[169];
  assign match_array[170] = N2832 & valid[170];
  assign N2832 = N2831 & N1734;
  assign N2831 = N2150 & en_i;
  assign empty_array[170] = N2833 & N2834;
  assign N2833 = N2150 & en_i;
  assign N2834 = ~valid[170];
  assign match_array[171] = N2836 & valid[171];
  assign N2836 = N2835 & N1735;
  assign N2835 = N2150 & en_i;
  assign empty_array[171] = N2837 & N2838;
  assign N2837 = N2150 & en_i;
  assign N2838 = ~valid[171];
  assign match_array[172] = N2840 & valid[172];
  assign N2840 = N2839 & N1736;
  assign N2839 = N2150 & en_i;
  assign empty_array[172] = N2841 & N2842;
  assign N2841 = N2150 & en_i;
  assign N2842 = ~valid[172];
  assign match_array[173] = N2844 & valid[173];
  assign N2844 = N2843 & N1737;
  assign N2843 = N2150 & en_i;
  assign empty_array[173] = N2845 & N2846;
  assign N2845 = N2150 & en_i;
  assign N2846 = ~valid[173];
  assign match_array[174] = N2848 & valid[174];
  assign N2848 = N2847 & N1738;
  assign N2847 = N2150 & en_i;
  assign empty_array[174] = N2849 & N2850;
  assign N2849 = N2150 & en_i;
  assign N2850 = ~valid[174];
  assign match_array[175] = N2852 & valid[175];
  assign N2852 = N2851 & N1739;
  assign N2851 = N2150 & en_i;
  assign empty_array[175] = N2853 & N2854;
  assign N2853 = N2150 & en_i;
  assign N2854 = ~valid[175];
  assign match_array[176] = N2856 & valid[176];
  assign N2856 = N2855 & N1740;
  assign N2855 = N2150 & en_i;
  assign empty_array[176] = N2857 & N2858;
  assign N2857 = N2150 & en_i;
  assign N2858 = ~valid[176];
  assign match_array[177] = N2860 & valid[177];
  assign N2860 = N2859 & N1741;
  assign N2859 = N2150 & en_i;
  assign empty_array[177] = N2861 & N2862;
  assign N2861 = N2150 & en_i;
  assign N2862 = ~valid[177];
  assign match_array[178] = N2864 & valid[178];
  assign N2864 = N2863 & N1742;
  assign N2863 = N2150 & en_i;
  assign empty_array[178] = N2865 & N2866;
  assign N2865 = N2150 & en_i;
  assign N2866 = ~valid[178];
  assign match_array[179] = N2868 & valid[179];
  assign N2868 = N2867 & N1743;
  assign N2867 = N2150 & en_i;
  assign empty_array[179] = N2869 & N2870;
  assign N2869 = N2150 & en_i;
  assign N2870 = ~valid[179];
  assign match_array[180] = N2872 & valid[180];
  assign N2872 = N2871 & N1744;
  assign N2871 = N2150 & en_i;
  assign empty_array[180] = N2873 & N2874;
  assign N2873 = N2150 & en_i;
  assign N2874 = ~valid[180];
  assign match_array[181] = N2876 & valid[181];
  assign N2876 = N2875 & N1745;
  assign N2875 = N2150 & en_i;
  assign empty_array[181] = N2877 & N2878;
  assign N2877 = N2150 & en_i;
  assign N2878 = ~valid[181];
  assign match_array[182] = N2880 & valid[182];
  assign N2880 = N2879 & N1746;
  assign N2879 = N2150 & en_i;
  assign empty_array[182] = N2881 & N2882;
  assign N2881 = N2150 & en_i;
  assign N2882 = ~valid[182];
  assign match_array[183] = N2884 & valid[183];
  assign N2884 = N2883 & N1747;
  assign N2883 = N2150 & en_i;
  assign empty_array[183] = N2885 & N2886;
  assign N2885 = N2150 & en_i;
  assign N2886 = ~valid[183];
  assign match_array[184] = N2888 & valid[184];
  assign N2888 = N2887 & N1748;
  assign N2887 = N2150 & en_i;
  assign empty_array[184] = N2889 & N2890;
  assign N2889 = N2150 & en_i;
  assign N2890 = ~valid[184];
  assign match_array[185] = N2892 & valid[185];
  assign N2892 = N2891 & N1749;
  assign N2891 = N2150 & en_i;
  assign empty_array[185] = N2893 & N2894;
  assign N2893 = N2150 & en_i;
  assign N2894 = ~valid[185];
  assign match_array[186] = N2896 & valid[186];
  assign N2896 = N2895 & N1750;
  assign N2895 = N2150 & en_i;
  assign empty_array[186] = N2897 & N2898;
  assign N2897 = N2150 & en_i;
  assign N2898 = ~valid[186];
  assign match_array[187] = N2900 & valid[187];
  assign N2900 = N2899 & N1751;
  assign N2899 = N2150 & en_i;
  assign empty_array[187] = N2901 & N2902;
  assign N2901 = N2150 & en_i;
  assign N2902 = ~valid[187];
  assign match_array[188] = N2904 & valid[188];
  assign N2904 = N2903 & N1752;
  assign N2903 = N2150 & en_i;
  assign empty_array[188] = N2905 & N2906;
  assign N2905 = N2150 & en_i;
  assign N2906 = ~valid[188];
  assign match_array[189] = N2908 & valid[189];
  assign N2908 = N2907 & N1753;
  assign N2907 = N2150 & en_i;
  assign empty_array[189] = N2909 & N2910;
  assign N2909 = N2150 & en_i;
  assign N2910 = ~valid[189];
  assign match_array[190] = N2912 & valid[190];
  assign N2912 = N2911 & N1754;
  assign N2911 = N2150 & en_i;
  assign empty_array[190] = N2913 & N2914;
  assign N2913 = N2150 & en_i;
  assign N2914 = ~valid[190];
  assign match_array[191] = N2916 & valid[191];
  assign N2916 = N2915 & N1755;
  assign N2915 = N2150 & en_i;
  assign empty_array[191] = N2917 & N2918;
  assign N2917 = N2150 & en_i;
  assign N2918 = ~valid[191];
  assign match_array[192] = N2920 & valid[192];
  assign N2920 = N2919 & N1756;
  assign N2919 = N2150 & en_i;
  assign empty_array[192] = N2921 & N2922;
  assign N2921 = N2150 & en_i;
  assign N2922 = ~valid[192];
  assign match_array[193] = N2924 & valid[193];
  assign N2924 = N2923 & N1757;
  assign N2923 = N2150 & en_i;
  assign empty_array[193] = N2925 & N2926;
  assign N2925 = N2150 & en_i;
  assign N2926 = ~valid[193];
  assign match_array[194] = N2928 & valid[194];
  assign N2928 = N2927 & N1758;
  assign N2927 = N2150 & en_i;
  assign empty_array[194] = N2929 & N2930;
  assign N2929 = N2150 & en_i;
  assign N2930 = ~valid[194];
  assign match_array[195] = N2932 & valid[195];
  assign N2932 = N2931 & N1759;
  assign N2931 = N2150 & en_i;
  assign empty_array[195] = N2933 & N2934;
  assign N2933 = N2150 & en_i;
  assign N2934 = ~valid[195];
  assign match_array[196] = N2936 & valid[196];
  assign N2936 = N2935 & N1760;
  assign N2935 = N2150 & en_i;
  assign empty_array[196] = N2937 & N2938;
  assign N2937 = N2150 & en_i;
  assign N2938 = ~valid[196];
  assign match_array[197] = N2940 & valid[197];
  assign N2940 = N2939 & N1761;
  assign N2939 = N2150 & en_i;
  assign empty_array[197] = N2941 & N2942;
  assign N2941 = N2150 & en_i;
  assign N2942 = ~valid[197];
  assign match_array[198] = N2944 & valid[198];
  assign N2944 = N2943 & N1762;
  assign N2943 = N2150 & en_i;
  assign empty_array[198] = N2945 & N2946;
  assign N2945 = N2150 & en_i;
  assign N2946 = ~valid[198];
  assign match_array[199] = N2948 & valid[199];
  assign N2948 = N2947 & N1763;
  assign N2947 = N2150 & en_i;
  assign empty_array[199] = N2949 & N2950;
  assign N2949 = N2150 & en_i;
  assign N2950 = ~valid[199];
  assign match_array[200] = N2952 & valid[200];
  assign N2952 = N2951 & N1764;
  assign N2951 = N2150 & en_i;
  assign empty_array[200] = N2953 & N2954;
  assign N2953 = N2150 & en_i;
  assign N2954 = ~valid[200];
  assign match_array[201] = N2956 & valid[201];
  assign N2956 = N2955 & N1765;
  assign N2955 = N2150 & en_i;
  assign empty_array[201] = N2957 & N2958;
  assign N2957 = N2150 & en_i;
  assign N2958 = ~valid[201];
  assign match_array[202] = N2960 & valid[202];
  assign N2960 = N2959 & N1766;
  assign N2959 = N2150 & en_i;
  assign empty_array[202] = N2961 & N2962;
  assign N2961 = N2150 & en_i;
  assign N2962 = ~valid[202];
  assign match_array[203] = N2964 & valid[203];
  assign N2964 = N2963 & N1767;
  assign N2963 = N2150 & en_i;
  assign empty_array[203] = N2965 & N2966;
  assign N2965 = N2150 & en_i;
  assign N2966 = ~valid[203];
  assign match_array[204] = N2968 & valid[204];
  assign N2968 = N2967 & N1768;
  assign N2967 = N2150 & en_i;
  assign empty_array[204] = N2969 & N2970;
  assign N2969 = N2150 & en_i;
  assign N2970 = ~valid[204];
  assign match_array[205] = N2972 & valid[205];
  assign N2972 = N2971 & N1769;
  assign N2971 = N2150 & en_i;
  assign empty_array[205] = N2973 & N2974;
  assign N2973 = N2150 & en_i;
  assign N2974 = ~valid[205];
  assign match_array[206] = N2976 & valid[206];
  assign N2976 = N2975 & N1770;
  assign N2975 = N2150 & en_i;
  assign empty_array[206] = N2977 & N2978;
  assign N2977 = N2150 & en_i;
  assign N2978 = ~valid[206];
  assign match_array[207] = N2980 & valid[207];
  assign N2980 = N2979 & N1771;
  assign N2979 = N2150 & en_i;
  assign empty_array[207] = N2981 & N2982;
  assign N2981 = N2150 & en_i;
  assign N2982 = ~valid[207];
  assign match_array[208] = N2984 & valid[208];
  assign N2984 = N2983 & N1772;
  assign N2983 = N2150 & en_i;
  assign empty_array[208] = N2985 & N2986;
  assign N2985 = N2150 & en_i;
  assign N2986 = ~valid[208];
  assign match_array[209] = N2988 & valid[209];
  assign N2988 = N2987 & N1773;
  assign N2987 = N2150 & en_i;
  assign empty_array[209] = N2989 & N2990;
  assign N2989 = N2150 & en_i;
  assign N2990 = ~valid[209];
  assign match_array[210] = N2992 & valid[210];
  assign N2992 = N2991 & N1774;
  assign N2991 = N2150 & en_i;
  assign empty_array[210] = N2993 & N2994;
  assign N2993 = N2150 & en_i;
  assign N2994 = ~valid[210];
  assign match_array[211] = N2996 & valid[211];
  assign N2996 = N2995 & N1775;
  assign N2995 = N2150 & en_i;
  assign empty_array[211] = N2997 & N2998;
  assign N2997 = N2150 & en_i;
  assign N2998 = ~valid[211];
  assign match_array[212] = N3000 & valid[212];
  assign N3000 = N2999 & N1776;
  assign N2999 = N2150 & en_i;
  assign empty_array[212] = N3001 & N3002;
  assign N3001 = N2150 & en_i;
  assign N3002 = ~valid[212];
  assign match_array[213] = N3004 & valid[213];
  assign N3004 = N3003 & N1777;
  assign N3003 = N2150 & en_i;
  assign empty_array[213] = N3005 & N3006;
  assign N3005 = N2150 & en_i;
  assign N3006 = ~valid[213];
  assign match_array[214] = N3008 & valid[214];
  assign N3008 = N3007 & N1778;
  assign N3007 = N2150 & en_i;
  assign empty_array[214] = N3009 & N3010;
  assign N3009 = N2150 & en_i;
  assign N3010 = ~valid[214];
  assign match_array[215] = N3012 & valid[215];
  assign N3012 = N3011 & N1779;
  assign N3011 = N2150 & en_i;
  assign empty_array[215] = N3013 & N3014;
  assign N3013 = N2150 & en_i;
  assign N3014 = ~valid[215];
  assign match_array[216] = N3016 & valid[216];
  assign N3016 = N3015 & N1780;
  assign N3015 = N2150 & en_i;
  assign empty_array[216] = N3017 & N3018;
  assign N3017 = N2150 & en_i;
  assign N3018 = ~valid[216];
  assign match_array[217] = N3020 & valid[217];
  assign N3020 = N3019 & N1781;
  assign N3019 = N2150 & en_i;
  assign empty_array[217] = N3021 & N3022;
  assign N3021 = N2150 & en_i;
  assign N3022 = ~valid[217];
  assign match_array[218] = N3024 & valid[218];
  assign N3024 = N3023 & N1782;
  assign N3023 = N2150 & en_i;
  assign empty_array[218] = N3025 & N3026;
  assign N3025 = N2150 & en_i;
  assign N3026 = ~valid[218];
  assign match_array[219] = N3028 & valid[219];
  assign N3028 = N3027 & N1783;
  assign N3027 = N2150 & en_i;
  assign empty_array[219] = N3029 & N3030;
  assign N3029 = N2150 & en_i;
  assign N3030 = ~valid[219];
  assign match_array[220] = N3032 & valid[220];
  assign N3032 = N3031 & N1784;
  assign N3031 = N2150 & en_i;
  assign empty_array[220] = N3033 & N3034;
  assign N3033 = N2150 & en_i;
  assign N3034 = ~valid[220];
  assign match_array[221] = N3036 & valid[221];
  assign N3036 = N3035 & N1785;
  assign N3035 = N2150 & en_i;
  assign empty_array[221] = N3037 & N3038;
  assign N3037 = N2150 & en_i;
  assign N3038 = ~valid[221];
  assign match_array[222] = N3040 & valid[222];
  assign N3040 = N3039 & N1786;
  assign N3039 = N2150 & en_i;
  assign empty_array[222] = N3041 & N3042;
  assign N3041 = N2150 & en_i;
  assign N3042 = ~valid[222];
  assign match_array[223] = N3044 & valid[223];
  assign N3044 = N3043 & N1787;
  assign N3043 = N2150 & en_i;
  assign empty_array[223] = N3045 & N3046;
  assign N3045 = N2150 & en_i;
  assign N3046 = ~valid[223];
  assign match_array[224] = N3048 & valid[224];
  assign N3048 = N3047 & N1788;
  assign N3047 = N2150 & en_i;
  assign empty_array[224] = N3049 & N3050;
  assign N3049 = N2150 & en_i;
  assign N3050 = ~valid[224];
  assign match_array[225] = N3052 & valid[225];
  assign N3052 = N3051 & N1789;
  assign N3051 = N2150 & en_i;
  assign empty_array[225] = N3053 & N3054;
  assign N3053 = N2150 & en_i;
  assign N3054 = ~valid[225];
  assign match_array[226] = N3056 & valid[226];
  assign N3056 = N3055 & N1790;
  assign N3055 = N2150 & en_i;
  assign empty_array[226] = N3057 & N3058;
  assign N3057 = N2150 & en_i;
  assign N3058 = ~valid[226];
  assign match_array[227] = N3060 & valid[227];
  assign N3060 = N3059 & N1791;
  assign N3059 = N2150 & en_i;
  assign empty_array[227] = N3061 & N3062;
  assign N3061 = N2150 & en_i;
  assign N3062 = ~valid[227];
  assign match_array[228] = N3064 & valid[228];
  assign N3064 = N3063 & N1792;
  assign N3063 = N2150 & en_i;
  assign empty_array[228] = N3065 & N3066;
  assign N3065 = N2150 & en_i;
  assign N3066 = ~valid[228];
  assign match_array[229] = N3068 & valid[229];
  assign N3068 = N3067 & N1793;
  assign N3067 = N2150 & en_i;
  assign empty_array[229] = N3069 & N3070;
  assign N3069 = N2150 & en_i;
  assign N3070 = ~valid[229];
  assign match_array[230] = N3072 & valid[230];
  assign N3072 = N3071 & N1794;
  assign N3071 = N2150 & en_i;
  assign empty_array[230] = N3073 & N3074;
  assign N3073 = N2150 & en_i;
  assign N3074 = ~valid[230];
  assign match_array[231] = N3076 & valid[231];
  assign N3076 = N3075 & N1795;
  assign N3075 = N2150 & en_i;
  assign empty_array[231] = N3077 & N3078;
  assign N3077 = N2150 & en_i;
  assign N3078 = ~valid[231];
  assign match_array[232] = N3080 & valid[232];
  assign N3080 = N3079 & N1796;
  assign N3079 = N2150 & en_i;
  assign empty_array[232] = N3081 & N3082;
  assign N3081 = N2150 & en_i;
  assign N3082 = ~valid[232];
  assign match_array[233] = N3084 & valid[233];
  assign N3084 = N3083 & N1797;
  assign N3083 = N2150 & en_i;
  assign empty_array[233] = N3085 & N3086;
  assign N3085 = N2150 & en_i;
  assign N3086 = ~valid[233];
  assign match_array[234] = N3088 & valid[234];
  assign N3088 = N3087 & N1798;
  assign N3087 = N2150 & en_i;
  assign empty_array[234] = N3089 & N3090;
  assign N3089 = N2150 & en_i;
  assign N3090 = ~valid[234];
  assign match_array[235] = N3092 & valid[235];
  assign N3092 = N3091 & N1799;
  assign N3091 = N2150 & en_i;
  assign empty_array[235] = N3093 & N3094;
  assign N3093 = N2150 & en_i;
  assign N3094 = ~valid[235];
  assign match_array[236] = N3096 & valid[236];
  assign N3096 = N3095 & N1800;
  assign N3095 = N2150 & en_i;
  assign empty_array[236] = N3097 & N3098;
  assign N3097 = N2150 & en_i;
  assign N3098 = ~valid[236];
  assign match_array[237] = N3100 & valid[237];
  assign N3100 = N3099 & N1801;
  assign N3099 = N2150 & en_i;
  assign empty_array[237] = N3101 & N3102;
  assign N3101 = N2150 & en_i;
  assign N3102 = ~valid[237];
  assign match_array[238] = N3104 & valid[238];
  assign N3104 = N3103 & N1802;
  assign N3103 = N2150 & en_i;
  assign empty_array[238] = N3105 & N3106;
  assign N3105 = N2150 & en_i;
  assign N3106 = ~valid[238];
  assign match_array[239] = N3108 & valid[239];
  assign N3108 = N3107 & N1803;
  assign N3107 = N2150 & en_i;
  assign empty_array[239] = N3109 & N3110;
  assign N3109 = N2150 & en_i;
  assign N3110 = ~valid[239];
  assign match_array[240] = N3112 & valid[240];
  assign N3112 = N3111 & N1804;
  assign N3111 = N2150 & en_i;
  assign empty_array[240] = N3113 & N3114;
  assign N3113 = N2150 & en_i;
  assign N3114 = ~valid[240];
  assign match_array[241] = N3116 & valid[241];
  assign N3116 = N3115 & N1805;
  assign N3115 = N2150 & en_i;
  assign empty_array[241] = N3117 & N3118;
  assign N3117 = N2150 & en_i;
  assign N3118 = ~valid[241];
  assign match_array[242] = N3120 & valid[242];
  assign N3120 = N3119 & N1806;
  assign N3119 = N2150 & en_i;
  assign empty_array[242] = N3121 & N3122;
  assign N3121 = N2150 & en_i;
  assign N3122 = ~valid[242];
  assign match_array[243] = N3124 & valid[243];
  assign N3124 = N3123 & N1807;
  assign N3123 = N2150 & en_i;
  assign empty_array[243] = N3125 & N3126;
  assign N3125 = N2150 & en_i;
  assign N3126 = ~valid[243];
  assign match_array[244] = N3128 & valid[244];
  assign N3128 = N3127 & N1808;
  assign N3127 = N2150 & en_i;
  assign empty_array[244] = N3129 & N3130;
  assign N3129 = N2150 & en_i;
  assign N3130 = ~valid[244];
  assign match_array[245] = N3132 & valid[245];
  assign N3132 = N3131 & N1809;
  assign N3131 = N2150 & en_i;
  assign empty_array[245] = N3133 & N3134;
  assign N3133 = N2150 & en_i;
  assign N3134 = ~valid[245];
  assign match_array[246] = N3136 & valid[246];
  assign N3136 = N3135 & N1810;
  assign N3135 = N2150 & en_i;
  assign empty_array[246] = N3137 & N3138;
  assign N3137 = N2150 & en_i;
  assign N3138 = ~valid[246];
  assign match_array[247] = N3140 & valid[247];
  assign N3140 = N3139 & N1811;
  assign N3139 = N2150 & en_i;
  assign empty_array[247] = N3141 & N3142;
  assign N3141 = N2150 & en_i;
  assign N3142 = ~valid[247];
  assign match_array[248] = N3144 & valid[248];
  assign N3144 = N3143 & N1812;
  assign N3143 = N2150 & en_i;
  assign empty_array[248] = N3145 & N3146;
  assign N3145 = N2150 & en_i;
  assign N3146 = ~valid[248];
  assign match_array[249] = N3148 & valid[249];
  assign N3148 = N3147 & N1813;
  assign N3147 = N2150 & en_i;
  assign empty_array[249] = N3149 & N3150;
  assign N3149 = N2150 & en_i;
  assign N3150 = ~valid[249];
  assign match_array[250] = N3152 & valid[250];
  assign N3152 = N3151 & N1814;
  assign N3151 = N2150 & en_i;
  assign empty_array[250] = N3153 & N3154;
  assign N3153 = N2150 & en_i;
  assign N3154 = ~valid[250];
  assign match_array[251] = N3156 & valid[251];
  assign N3156 = N3155 & N1815;
  assign N3155 = N2150 & en_i;
  assign empty_array[251] = N3157 & N3158;
  assign N3157 = N2150 & en_i;
  assign N3158 = ~valid[251];
  assign match_array[252] = N3160 & valid[252];
  assign N3160 = N3159 & N1816;
  assign N3159 = N2150 & en_i;
  assign empty_array[252] = N3161 & N3162;
  assign N3161 = N2150 & en_i;
  assign N3162 = ~valid[252];
  assign match_array[253] = N3164 & valid[253];
  assign N3164 = N3163 & N1817;
  assign N3163 = N2150 & en_i;
  assign empty_array[253] = N3165 & N3166;
  assign N3165 = N2150 & en_i;
  assign N3166 = ~valid[253];
  assign match_array[254] = N3168 & valid[254];
  assign N3168 = N3167 & N1818;
  assign N3167 = N2150 & en_i;
  assign empty_array[254] = N3169 & N3170;
  assign N3169 = N2150 & en_i;
  assign N3170 = ~valid[254];
  assign match_array[255] = N3172 & valid[255];
  assign N3172 = N3171 & N1819;
  assign N3171 = N2150 & en_i;
  assign empty_array[255] = N3173 & N3174;
  assign N3173 = N2150 & en_i;
  assign N3174 = ~valid[255];
  assign match_array[256] = N3176 & valid[256];
  assign N3176 = N3175 & N1820;
  assign N3175 = N2150 & en_i;
  assign empty_array[256] = N3177 & N3178;
  assign N3177 = N2150 & en_i;
  assign N3178 = ~valid[256];
  assign match_array[257] = N3180 & valid[257];
  assign N3180 = N3179 & N1821;
  assign N3179 = N2150 & en_i;
  assign empty_array[257] = N3181 & N3182;
  assign N3181 = N2150 & en_i;
  assign N3182 = ~valid[257];
  assign match_array[258] = N3184 & valid[258];
  assign N3184 = N3183 & N1822;
  assign N3183 = N2150 & en_i;
  assign empty_array[258] = N3185 & N3186;
  assign N3185 = N2150 & en_i;
  assign N3186 = ~valid[258];
  assign match_array[259] = N3188 & valid[259];
  assign N3188 = N3187 & N1823;
  assign N3187 = N2150 & en_i;
  assign empty_array[259] = N3189 & N3190;
  assign N3189 = N2150 & en_i;
  assign N3190 = ~valid[259];
  assign match_array[260] = N3192 & valid[260];
  assign N3192 = N3191 & N1824;
  assign N3191 = N2150 & en_i;
  assign empty_array[260] = N3193 & N3194;
  assign N3193 = N2150 & en_i;
  assign N3194 = ~valid[260];
  assign match_array[261] = N3196 & valid[261];
  assign N3196 = N3195 & N1825;
  assign N3195 = N2150 & en_i;
  assign empty_array[261] = N3197 & N3198;
  assign N3197 = N2150 & en_i;
  assign N3198 = ~valid[261];
  assign match_array[262] = N3200 & valid[262];
  assign N3200 = N3199 & N1826;
  assign N3199 = N2150 & en_i;
  assign empty_array[262] = N3201 & N3202;
  assign N3201 = N2150 & en_i;
  assign N3202 = ~valid[262];
  assign match_array[263] = N3204 & valid[263];
  assign N3204 = N3203 & N1827;
  assign N3203 = N2150 & en_i;
  assign empty_array[263] = N3205 & N3206;
  assign N3205 = N2150 & en_i;
  assign N3206 = ~valid[263];
  assign match_array[264] = N3208 & valid[264];
  assign N3208 = N3207 & N1828;
  assign N3207 = N2150 & en_i;
  assign empty_array[264] = N3209 & N3210;
  assign N3209 = N2150 & en_i;
  assign N3210 = ~valid[264];
  assign match_array[265] = N3212 & valid[265];
  assign N3212 = N3211 & N1829;
  assign N3211 = N2150 & en_i;
  assign empty_array[265] = N3213 & N3214;
  assign N3213 = N2150 & en_i;
  assign N3214 = ~valid[265];
  assign match_array[266] = N3216 & valid[266];
  assign N3216 = N3215 & N1830;
  assign N3215 = N2150 & en_i;
  assign empty_array[266] = N3217 & N3218;
  assign N3217 = N2150 & en_i;
  assign N3218 = ~valid[266];
  assign match_array[267] = N3220 & valid[267];
  assign N3220 = N3219 & N1831;
  assign N3219 = N2150 & en_i;
  assign empty_array[267] = N3221 & N3222;
  assign N3221 = N2150 & en_i;
  assign N3222 = ~valid[267];
  assign match_array[268] = N3224 & valid[268];
  assign N3224 = N3223 & N1832;
  assign N3223 = N2150 & en_i;
  assign empty_array[268] = N3225 & N3226;
  assign N3225 = N2150 & en_i;
  assign N3226 = ~valid[268];
  assign match_array[269] = N3228 & valid[269];
  assign N3228 = N3227 & N1833;
  assign N3227 = N2150 & en_i;
  assign empty_array[269] = N3229 & N3230;
  assign N3229 = N2150 & en_i;
  assign N3230 = ~valid[269];
  assign match_array[270] = N3232 & valid[270];
  assign N3232 = N3231 & N1834;
  assign N3231 = N2150 & en_i;
  assign empty_array[270] = N3233 & N3234;
  assign N3233 = N2150 & en_i;
  assign N3234 = ~valid[270];
  assign match_array[271] = N3236 & valid[271];
  assign N3236 = N3235 & N1835;
  assign N3235 = N2150 & en_i;
  assign empty_array[271] = N3237 & N3238;
  assign N3237 = N2150 & en_i;
  assign N3238 = ~valid[271];
  assign match_array[272] = N3240 & valid[272];
  assign N3240 = N3239 & N1836;
  assign N3239 = N2150 & en_i;
  assign empty_array[272] = N3241 & N3242;
  assign N3241 = N2150 & en_i;
  assign N3242 = ~valid[272];
  assign match_array[273] = N3244 & valid[273];
  assign N3244 = N3243 & N1837;
  assign N3243 = N2150 & en_i;
  assign empty_array[273] = N3245 & N3246;
  assign N3245 = N2150 & en_i;
  assign N3246 = ~valid[273];
  assign match_array[274] = N3248 & valid[274];
  assign N3248 = N3247 & N1838;
  assign N3247 = N2150 & en_i;
  assign empty_array[274] = N3249 & N3250;
  assign N3249 = N2150 & en_i;
  assign N3250 = ~valid[274];
  assign match_array[275] = N3252 & valid[275];
  assign N3252 = N3251 & N1839;
  assign N3251 = N2150 & en_i;
  assign empty_array[275] = N3253 & N3254;
  assign N3253 = N2150 & en_i;
  assign N3254 = ~valid[275];
  assign match_array[276] = N3256 & valid[276];
  assign N3256 = N3255 & N1840;
  assign N3255 = N2150 & en_i;
  assign empty_array[276] = N3257 & N3258;
  assign N3257 = N2150 & en_i;
  assign N3258 = ~valid[276];
  assign match_array[277] = N3260 & valid[277];
  assign N3260 = N3259 & N1841;
  assign N3259 = N2150 & en_i;
  assign empty_array[277] = N3261 & N3262;
  assign N3261 = N2150 & en_i;
  assign N3262 = ~valid[277];
  assign match_array[278] = N3264 & valid[278];
  assign N3264 = N3263 & N1842;
  assign N3263 = N2150 & en_i;
  assign empty_array[278] = N3265 & N3266;
  assign N3265 = N2150 & en_i;
  assign N3266 = ~valid[278];
  assign match_array[279] = N3268 & valid[279];
  assign N3268 = N3267 & N1843;
  assign N3267 = N2150 & en_i;
  assign empty_array[279] = N3269 & N3270;
  assign N3269 = N2150 & en_i;
  assign N3270 = ~valid[279];
  assign match_array[280] = N3272 & valid[280];
  assign N3272 = N3271 & N1844;
  assign N3271 = N2150 & en_i;
  assign empty_array[280] = N3273 & N3274;
  assign N3273 = N2150 & en_i;
  assign N3274 = ~valid[280];
  assign match_array[281] = N3276 & valid[281];
  assign N3276 = N3275 & N1845;
  assign N3275 = N2150 & en_i;
  assign empty_array[281] = N3277 & N3278;
  assign N3277 = N2150 & en_i;
  assign N3278 = ~valid[281];
  assign match_array[282] = N3280 & valid[282];
  assign N3280 = N3279 & N1846;
  assign N3279 = N2150 & en_i;
  assign empty_array[282] = N3281 & N3282;
  assign N3281 = N2150 & en_i;
  assign N3282 = ~valid[282];
  assign match_array[283] = N3284 & valid[283];
  assign N3284 = N3283 & N1847;
  assign N3283 = N2150 & en_i;
  assign empty_array[283] = N3285 & N3286;
  assign N3285 = N2150 & en_i;
  assign N3286 = ~valid[283];
  assign match_array[284] = N3288 & valid[284];
  assign N3288 = N3287 & N1848;
  assign N3287 = N2150 & en_i;
  assign empty_array[284] = N3289 & N3290;
  assign N3289 = N2150 & en_i;
  assign N3290 = ~valid[284];
  assign match_array[285] = N3292 & valid[285];
  assign N3292 = N3291 & N1849;
  assign N3291 = N2150 & en_i;
  assign empty_array[285] = N3293 & N3294;
  assign N3293 = N2150 & en_i;
  assign N3294 = ~valid[285];
  assign match_array[286] = N3296 & valid[286];
  assign N3296 = N3295 & N1850;
  assign N3295 = N2150 & en_i;
  assign empty_array[286] = N3297 & N3298;
  assign N3297 = N2150 & en_i;
  assign N3298 = ~valid[286];
  assign match_array[287] = N3300 & valid[287];
  assign N3300 = N3299 & N1851;
  assign N3299 = N2150 & en_i;
  assign empty_array[287] = N3301 & N3302;
  assign N3301 = N2150 & en_i;
  assign N3302 = ~valid[287];
  assign match_array[288] = N3304 & valid[288];
  assign N3304 = N3303 & N1852;
  assign N3303 = N2150 & en_i;
  assign empty_array[288] = N3305 & N3306;
  assign N3305 = N2150 & en_i;
  assign N3306 = ~valid[288];
  assign match_array[289] = N3308 & valid[289];
  assign N3308 = N3307 & N1853;
  assign N3307 = N2150 & en_i;
  assign empty_array[289] = N3309 & N3310;
  assign N3309 = N2150 & en_i;
  assign N3310 = ~valid[289];
  assign match_array[290] = N3312 & valid[290];
  assign N3312 = N3311 & N1854;
  assign N3311 = N2150 & en_i;
  assign empty_array[290] = N3313 & N3314;
  assign N3313 = N2150 & en_i;
  assign N3314 = ~valid[290];
  assign match_array[291] = N3316 & valid[291];
  assign N3316 = N3315 & N1855;
  assign N3315 = N2150 & en_i;
  assign empty_array[291] = N3317 & N3318;
  assign N3317 = N2150 & en_i;
  assign N3318 = ~valid[291];
  assign match_array[292] = N3320 & valid[292];
  assign N3320 = N3319 & N1856;
  assign N3319 = N2150 & en_i;
  assign empty_array[292] = N3321 & N3322;
  assign N3321 = N2150 & en_i;
  assign N3322 = ~valid[292];
  assign match_array[293] = N3324 & valid[293];
  assign N3324 = N3323 & N1857;
  assign N3323 = N2150 & en_i;
  assign empty_array[293] = N3325 & N3326;
  assign N3325 = N2150 & en_i;
  assign N3326 = ~valid[293];
  assign match_array[294] = N3328 & valid[294];
  assign N3328 = N3327 & N1858;
  assign N3327 = N2150 & en_i;
  assign empty_array[294] = N3329 & N3330;
  assign N3329 = N2150 & en_i;
  assign N3330 = ~valid[294];
  assign match_array[295] = N3332 & valid[295];
  assign N3332 = N3331 & N1859;
  assign N3331 = N2150 & en_i;
  assign empty_array[295] = N3333 & N3334;
  assign N3333 = N2150 & en_i;
  assign N3334 = ~valid[295];
  assign match_array[296] = N3336 & valid[296];
  assign N3336 = N3335 & N1860;
  assign N3335 = N2150 & en_i;
  assign empty_array[296] = N3337 & N3338;
  assign N3337 = N2150 & en_i;
  assign N3338 = ~valid[296];
  assign match_array[297] = N3340 & valid[297];
  assign N3340 = N3339 & N1861;
  assign N3339 = N2150 & en_i;
  assign empty_array[297] = N3341 & N3342;
  assign N3341 = N2150 & en_i;
  assign N3342 = ~valid[297];
  assign match_array[298] = N3344 & valid[298];
  assign N3344 = N3343 & N1862;
  assign N3343 = N2150 & en_i;
  assign empty_array[298] = N3345 & N3346;
  assign N3345 = N2150 & en_i;
  assign N3346 = ~valid[298];
  assign match_array[299] = N3348 & valid[299];
  assign N3348 = N3347 & N1863;
  assign N3347 = N2150 & en_i;
  assign empty_array[299] = N3349 & N3350;
  assign N3349 = N2150 & en_i;
  assign N3350 = ~valid[299];
  assign match_array[300] = N3352 & valid[300];
  assign N3352 = N3351 & N1864;
  assign N3351 = N2150 & en_i;
  assign empty_array[300] = N3353 & N3354;
  assign N3353 = N2150 & en_i;
  assign N3354 = ~valid[300];
  assign match_array[301] = N3356 & valid[301];
  assign N3356 = N3355 & N1865;
  assign N3355 = N2150 & en_i;
  assign empty_array[301] = N3357 & N3358;
  assign N3357 = N2150 & en_i;
  assign N3358 = ~valid[301];
  assign match_array[302] = N3360 & valid[302];
  assign N3360 = N3359 & N1866;
  assign N3359 = N2150 & en_i;
  assign empty_array[302] = N3361 & N3362;
  assign N3361 = N2150 & en_i;
  assign N3362 = ~valid[302];
  assign match_array[303] = N3364 & valid[303];
  assign N3364 = N3363 & N1867;
  assign N3363 = N2150 & en_i;
  assign empty_array[303] = N3365 & N3366;
  assign N3365 = N2150 & en_i;
  assign N3366 = ~valid[303];
  assign match_array[304] = N3368 & valid[304];
  assign N3368 = N3367 & N1868;
  assign N3367 = N2150 & en_i;
  assign empty_array[304] = N3369 & N3370;
  assign N3369 = N2150 & en_i;
  assign N3370 = ~valid[304];
  assign match_array[305] = N3372 & valid[305];
  assign N3372 = N3371 & N1869;
  assign N3371 = N2150 & en_i;
  assign empty_array[305] = N3373 & N3374;
  assign N3373 = N2150 & en_i;
  assign N3374 = ~valid[305];
  assign match_array[306] = N3376 & valid[306];
  assign N3376 = N3375 & N1870;
  assign N3375 = N2150 & en_i;
  assign empty_array[306] = N3377 & N3378;
  assign N3377 = N2150 & en_i;
  assign N3378 = ~valid[306];
  assign match_array[307] = N3380 & valid[307];
  assign N3380 = N3379 & N1871;
  assign N3379 = N2150 & en_i;
  assign empty_array[307] = N3381 & N3382;
  assign N3381 = N2150 & en_i;
  assign N3382 = ~valid[307];
  assign match_array[308] = N3384 & valid[308];
  assign N3384 = N3383 & N1872;
  assign N3383 = N2150 & en_i;
  assign empty_array[308] = N3385 & N3386;
  assign N3385 = N2150 & en_i;
  assign N3386 = ~valid[308];
  assign match_array[309] = N3388 & valid[309];
  assign N3388 = N3387 & N1873;
  assign N3387 = N2150 & en_i;
  assign empty_array[309] = N3389 & N3390;
  assign N3389 = N2150 & en_i;
  assign N3390 = ~valid[309];
  assign match_array[310] = N3392 & valid[310];
  assign N3392 = N3391 & N1874;
  assign N3391 = N2150 & en_i;
  assign empty_array[310] = N3393 & N3394;
  assign N3393 = N2150 & en_i;
  assign N3394 = ~valid[310];
  assign match_array[311] = N3396 & valid[311];
  assign N3396 = N3395 & N1875;
  assign N3395 = N2150 & en_i;
  assign empty_array[311] = N3397 & N3398;
  assign N3397 = N2150 & en_i;
  assign N3398 = ~valid[311];
  assign match_array[312] = N3400 & valid[312];
  assign N3400 = N3399 & N1876;
  assign N3399 = N2150 & en_i;
  assign empty_array[312] = N3401 & N3402;
  assign N3401 = N2150 & en_i;
  assign N3402 = ~valid[312];
  assign match_array[313] = N3404 & valid[313];
  assign N3404 = N3403 & N1877;
  assign N3403 = N2150 & en_i;
  assign empty_array[313] = N3405 & N3406;
  assign N3405 = N2150 & en_i;
  assign N3406 = ~valid[313];
  assign match_array[314] = N3408 & valid[314];
  assign N3408 = N3407 & N1878;
  assign N3407 = N2150 & en_i;
  assign empty_array[314] = N3409 & N3410;
  assign N3409 = N2150 & en_i;
  assign N3410 = ~valid[314];
  assign match_array[315] = N3412 & valid[315];
  assign N3412 = N3411 & N1879;
  assign N3411 = N2150 & en_i;
  assign empty_array[315] = N3413 & N3414;
  assign N3413 = N2150 & en_i;
  assign N3414 = ~valid[315];
  assign match_array[316] = N3416 & valid[316];
  assign N3416 = N3415 & N1880;
  assign N3415 = N2150 & en_i;
  assign empty_array[316] = N3417 & N3418;
  assign N3417 = N2150 & en_i;
  assign N3418 = ~valid[316];
  assign match_array[317] = N3420 & valid[317];
  assign N3420 = N3419 & N1881;
  assign N3419 = N2150 & en_i;
  assign empty_array[317] = N3421 & N3422;
  assign N3421 = N2150 & en_i;
  assign N3422 = ~valid[317];
  assign match_array[318] = N3424 & valid[318];
  assign N3424 = N3423 & N1882;
  assign N3423 = N2150 & en_i;
  assign empty_array[318] = N3425 & N3426;
  assign N3425 = N2150 & en_i;
  assign N3426 = ~valid[318];
  assign match_array[319] = N3428 & valid[319];
  assign N3428 = N3427 & N1883;
  assign N3427 = N2150 & en_i;
  assign empty_array[319] = N3429 & N3430;
  assign N3429 = N2150 & en_i;
  assign N3430 = ~valid[319];
  assign match_array[320] = N3432 & valid[320];
  assign N3432 = N3431 & N1884;
  assign N3431 = N2150 & en_i;
  assign empty_array[320] = N3433 & N3434;
  assign N3433 = N2150 & en_i;
  assign N3434 = ~valid[320];
  assign match_array[321] = N3436 & valid[321];
  assign N3436 = N3435 & N1885;
  assign N3435 = N2150 & en_i;
  assign empty_array[321] = N3437 & N3438;
  assign N3437 = N2150 & en_i;
  assign N3438 = ~valid[321];
  assign match_array[322] = N3440 & valid[322];
  assign N3440 = N3439 & N1886;
  assign N3439 = N2150 & en_i;
  assign empty_array[322] = N3441 & N3442;
  assign N3441 = N2150 & en_i;
  assign N3442 = ~valid[322];
  assign match_array[323] = N3444 & valid[323];
  assign N3444 = N3443 & N1887;
  assign N3443 = N2150 & en_i;
  assign empty_array[323] = N3445 & N3446;
  assign N3445 = N2150 & en_i;
  assign N3446 = ~valid[323];
  assign match_array[324] = N3448 & valid[324];
  assign N3448 = N3447 & N1888;
  assign N3447 = N2150 & en_i;
  assign empty_array[324] = N3449 & N3450;
  assign N3449 = N2150 & en_i;
  assign N3450 = ~valid[324];
  assign match_array[325] = N3452 & valid[325];
  assign N3452 = N3451 & N1889;
  assign N3451 = N2150 & en_i;
  assign empty_array[325] = N3453 & N3454;
  assign N3453 = N2150 & en_i;
  assign N3454 = ~valid[325];
  assign match_array[326] = N3456 & valid[326];
  assign N3456 = N3455 & N1890;
  assign N3455 = N2150 & en_i;
  assign empty_array[326] = N3457 & N3458;
  assign N3457 = N2150 & en_i;
  assign N3458 = ~valid[326];
  assign match_array[327] = N3460 & valid[327];
  assign N3460 = N3459 & N1891;
  assign N3459 = N2150 & en_i;
  assign empty_array[327] = N3461 & N3462;
  assign N3461 = N2150 & en_i;
  assign N3462 = ~valid[327];
  assign match_array[328] = N3464 & valid[328];
  assign N3464 = N3463 & N1892;
  assign N3463 = N2150 & en_i;
  assign empty_array[328] = N3465 & N3466;
  assign N3465 = N2150 & en_i;
  assign N3466 = ~valid[328];
  assign match_array[329] = N3468 & valid[329];
  assign N3468 = N3467 & N1893;
  assign N3467 = N2150 & en_i;
  assign empty_array[329] = N3469 & N3470;
  assign N3469 = N2150 & en_i;
  assign N3470 = ~valid[329];
  assign match_array[330] = N3472 & valid[330];
  assign N3472 = N3471 & N1894;
  assign N3471 = N2150 & en_i;
  assign empty_array[330] = N3473 & N3474;
  assign N3473 = N2150 & en_i;
  assign N3474 = ~valid[330];
  assign match_array[331] = N3476 & valid[331];
  assign N3476 = N3475 & N1895;
  assign N3475 = N2150 & en_i;
  assign empty_array[331] = N3477 & N3478;
  assign N3477 = N2150 & en_i;
  assign N3478 = ~valid[331];
  assign match_array[332] = N3480 & valid[332];
  assign N3480 = N3479 & N1896;
  assign N3479 = N2150 & en_i;
  assign empty_array[332] = N3481 & N3482;
  assign N3481 = N2150 & en_i;
  assign N3482 = ~valid[332];
  assign match_array[333] = N3484 & valid[333];
  assign N3484 = N3483 & N1897;
  assign N3483 = N2150 & en_i;
  assign empty_array[333] = N3485 & N3486;
  assign N3485 = N2150 & en_i;
  assign N3486 = ~valid[333];
  assign match_array[334] = N3488 & valid[334];
  assign N3488 = N3487 & N1898;
  assign N3487 = N2150 & en_i;
  assign empty_array[334] = N3489 & N3490;
  assign N3489 = N2150 & en_i;
  assign N3490 = ~valid[334];
  assign match_array[335] = N3492 & valid[335];
  assign N3492 = N3491 & N1899;
  assign N3491 = N2150 & en_i;
  assign empty_array[335] = N3493 & N3494;
  assign N3493 = N2150 & en_i;
  assign N3494 = ~valid[335];
  assign match_array[336] = N3496 & valid[336];
  assign N3496 = N3495 & N1900;
  assign N3495 = N2150 & en_i;
  assign empty_array[336] = N3497 & N3498;
  assign N3497 = N2150 & en_i;
  assign N3498 = ~valid[336];
  assign match_array[337] = N3500 & valid[337];
  assign N3500 = N3499 & N1901;
  assign N3499 = N2150 & en_i;
  assign empty_array[337] = N3501 & N3502;
  assign N3501 = N2150 & en_i;
  assign N3502 = ~valid[337];
  assign match_array[338] = N3504 & valid[338];
  assign N3504 = N3503 & N1902;
  assign N3503 = N2150 & en_i;
  assign empty_array[338] = N3505 & N3506;
  assign N3505 = N2150 & en_i;
  assign N3506 = ~valid[338];
  assign match_array[339] = N3508 & valid[339];
  assign N3508 = N3507 & N1903;
  assign N3507 = N2150 & en_i;
  assign empty_array[339] = N3509 & N3510;
  assign N3509 = N2150 & en_i;
  assign N3510 = ~valid[339];
  assign match_array[340] = N3512 & valid[340];
  assign N3512 = N3511 & N1904;
  assign N3511 = N2150 & en_i;
  assign empty_array[340] = N3513 & N3514;
  assign N3513 = N2150 & en_i;
  assign N3514 = ~valid[340];
  assign match_array[341] = N3516 & valid[341];
  assign N3516 = N3515 & N1905;
  assign N3515 = N2150 & en_i;
  assign empty_array[341] = N3517 & N3518;
  assign N3517 = N2150 & en_i;
  assign N3518 = ~valid[341];
  assign match_array[342] = N3520 & valid[342];
  assign N3520 = N3519 & N1906;
  assign N3519 = N2150 & en_i;
  assign empty_array[342] = N3521 & N3522;
  assign N3521 = N2150 & en_i;
  assign N3522 = ~valid[342];
  assign match_array[343] = N3524 & valid[343];
  assign N3524 = N3523 & N1907;
  assign N3523 = N2150 & en_i;
  assign empty_array[343] = N3525 & N3526;
  assign N3525 = N2150 & en_i;
  assign N3526 = ~valid[343];
  assign match_array[344] = N3528 & valid[344];
  assign N3528 = N3527 & N1908;
  assign N3527 = N2150 & en_i;
  assign empty_array[344] = N3529 & N3530;
  assign N3529 = N2150 & en_i;
  assign N3530 = ~valid[344];
  assign match_array[345] = N3532 & valid[345];
  assign N3532 = N3531 & N1909;
  assign N3531 = N2150 & en_i;
  assign empty_array[345] = N3533 & N3534;
  assign N3533 = N2150 & en_i;
  assign N3534 = ~valid[345];
  assign match_array[346] = N3536 & valid[346];
  assign N3536 = N3535 & N1910;
  assign N3535 = N2150 & en_i;
  assign empty_array[346] = N3537 & N3538;
  assign N3537 = N2150 & en_i;
  assign N3538 = ~valid[346];
  assign match_array[347] = N3540 & valid[347];
  assign N3540 = N3539 & N1911;
  assign N3539 = N2150 & en_i;
  assign empty_array[347] = N3541 & N3542;
  assign N3541 = N2150 & en_i;
  assign N3542 = ~valid[347];
  assign match_array[348] = N3544 & valid[348];
  assign N3544 = N3543 & N1912;
  assign N3543 = N2150 & en_i;
  assign empty_array[348] = N3545 & N3546;
  assign N3545 = N2150 & en_i;
  assign N3546 = ~valid[348];
  assign match_array[349] = N3548 & valid[349];
  assign N3548 = N3547 & N1913;
  assign N3547 = N2150 & en_i;
  assign empty_array[349] = N3549 & N3550;
  assign N3549 = N2150 & en_i;
  assign N3550 = ~valid[349];
  assign match_array[350] = N3552 & valid[350];
  assign N3552 = N3551 & N1914;
  assign N3551 = N2150 & en_i;
  assign empty_array[350] = N3553 & N3554;
  assign N3553 = N2150 & en_i;
  assign N3554 = ~valid[350];
  assign match_array[351] = N3556 & valid[351];
  assign N3556 = N3555 & N1915;
  assign N3555 = N2150 & en_i;
  assign empty_array[351] = N3557 & N3558;
  assign N3557 = N2150 & en_i;
  assign N3558 = ~valid[351];
  assign match_array[352] = N3560 & valid[352];
  assign N3560 = N3559 & N1916;
  assign N3559 = N2150 & en_i;
  assign empty_array[352] = N3561 & N3562;
  assign N3561 = N2150 & en_i;
  assign N3562 = ~valid[352];
  assign match_array[353] = N3564 & valid[353];
  assign N3564 = N3563 & N1917;
  assign N3563 = N2150 & en_i;
  assign empty_array[353] = N3565 & N3566;
  assign N3565 = N2150 & en_i;
  assign N3566 = ~valid[353];
  assign match_array[354] = N3568 & valid[354];
  assign N3568 = N3567 & N1918;
  assign N3567 = N2150 & en_i;
  assign empty_array[354] = N3569 & N3570;
  assign N3569 = N2150 & en_i;
  assign N3570 = ~valid[354];
  assign match_array[355] = N3572 & valid[355];
  assign N3572 = N3571 & N1919;
  assign N3571 = N2150 & en_i;
  assign empty_array[355] = N3573 & N3574;
  assign N3573 = N2150 & en_i;
  assign N3574 = ~valid[355];
  assign match_array[356] = N3576 & valid[356];
  assign N3576 = N3575 & N1920;
  assign N3575 = N2150 & en_i;
  assign empty_array[356] = N3577 & N3578;
  assign N3577 = N2150 & en_i;
  assign N3578 = ~valid[356];
  assign match_array[357] = N3580 & valid[357];
  assign N3580 = N3579 & N1921;
  assign N3579 = N2150 & en_i;
  assign empty_array[357] = N3581 & N3582;
  assign N3581 = N2150 & en_i;
  assign N3582 = ~valid[357];
  assign match_array[358] = N3584 & valid[358];
  assign N3584 = N3583 & N1922;
  assign N3583 = N2150 & en_i;
  assign empty_array[358] = N3585 & N3586;
  assign N3585 = N2150 & en_i;
  assign N3586 = ~valid[358];
  assign match_array[359] = N3588 & valid[359];
  assign N3588 = N3587 & N1923;
  assign N3587 = N2150 & en_i;
  assign empty_array[359] = N3589 & N3590;
  assign N3589 = N2150 & en_i;
  assign N3590 = ~valid[359];
  assign match_array[360] = N3592 & valid[360];
  assign N3592 = N3591 & N1924;
  assign N3591 = N2150 & en_i;
  assign empty_array[360] = N3593 & N3594;
  assign N3593 = N2150 & en_i;
  assign N3594 = ~valid[360];
  assign match_array[361] = N3596 & valid[361];
  assign N3596 = N3595 & N1925;
  assign N3595 = N2150 & en_i;
  assign empty_array[361] = N3597 & N3598;
  assign N3597 = N2150 & en_i;
  assign N3598 = ~valid[361];
  assign match_array[362] = N3600 & valid[362];
  assign N3600 = N3599 & N1926;
  assign N3599 = N2150 & en_i;
  assign empty_array[362] = N3601 & N3602;
  assign N3601 = N2150 & en_i;
  assign N3602 = ~valid[362];
  assign match_array[363] = N3604 & valid[363];
  assign N3604 = N3603 & N1927;
  assign N3603 = N2150 & en_i;
  assign empty_array[363] = N3605 & N3606;
  assign N3605 = N2150 & en_i;
  assign N3606 = ~valid[363];
  assign match_array[364] = N3608 & valid[364];
  assign N3608 = N3607 & N1928;
  assign N3607 = N2150 & en_i;
  assign empty_array[364] = N3609 & N3610;
  assign N3609 = N2150 & en_i;
  assign N3610 = ~valid[364];
  assign match_array[365] = N3612 & valid[365];
  assign N3612 = N3611 & N1929;
  assign N3611 = N2150 & en_i;
  assign empty_array[365] = N3613 & N3614;
  assign N3613 = N2150 & en_i;
  assign N3614 = ~valid[365];
  assign match_array[366] = N3616 & valid[366];
  assign N3616 = N3615 & N1930;
  assign N3615 = N2150 & en_i;
  assign empty_array[366] = N3617 & N3618;
  assign N3617 = N2150 & en_i;
  assign N3618 = ~valid[366];
  assign match_array[367] = N3620 & valid[367];
  assign N3620 = N3619 & N1931;
  assign N3619 = N2150 & en_i;
  assign empty_array[367] = N3621 & N3622;
  assign N3621 = N2150 & en_i;
  assign N3622 = ~valid[367];
  assign match_array[368] = N3624 & valid[368];
  assign N3624 = N3623 & N1932;
  assign N3623 = N2150 & en_i;
  assign empty_array[368] = N3625 & N3626;
  assign N3625 = N2150 & en_i;
  assign N3626 = ~valid[368];
  assign match_array[369] = N3628 & valid[369];
  assign N3628 = N3627 & N1933;
  assign N3627 = N2150 & en_i;
  assign empty_array[369] = N3629 & N3630;
  assign N3629 = N2150 & en_i;
  assign N3630 = ~valid[369];
  assign match_array[370] = N3632 & valid[370];
  assign N3632 = N3631 & N1934;
  assign N3631 = N2150 & en_i;
  assign empty_array[370] = N3633 & N3634;
  assign N3633 = N2150 & en_i;
  assign N3634 = ~valid[370];
  assign match_array[371] = N3636 & valid[371];
  assign N3636 = N3635 & N1935;
  assign N3635 = N2150 & en_i;
  assign empty_array[371] = N3637 & N3638;
  assign N3637 = N2150 & en_i;
  assign N3638 = ~valid[371];
  assign match_array[372] = N3640 & valid[372];
  assign N3640 = N3639 & N1936;
  assign N3639 = N2150 & en_i;
  assign empty_array[372] = N3641 & N3642;
  assign N3641 = N2150 & en_i;
  assign N3642 = ~valid[372];
  assign match_array[373] = N3644 & valid[373];
  assign N3644 = N3643 & N1937;
  assign N3643 = N2150 & en_i;
  assign empty_array[373] = N3645 & N3646;
  assign N3645 = N2150 & en_i;
  assign N3646 = ~valid[373];
  assign match_array[374] = N3648 & valid[374];
  assign N3648 = N3647 & N1938;
  assign N3647 = N2150 & en_i;
  assign empty_array[374] = N3649 & N3650;
  assign N3649 = N2150 & en_i;
  assign N3650 = ~valid[374];
  assign match_array[375] = N3652 & valid[375];
  assign N3652 = N3651 & N1939;
  assign N3651 = N2150 & en_i;
  assign empty_array[375] = N3653 & N3654;
  assign N3653 = N2150 & en_i;
  assign N3654 = ~valid[375];
  assign match_array[376] = N3656 & valid[376];
  assign N3656 = N3655 & N1940;
  assign N3655 = N2150 & en_i;
  assign empty_array[376] = N3657 & N3658;
  assign N3657 = N2150 & en_i;
  assign N3658 = ~valid[376];
  assign match_array[377] = N3660 & valid[377];
  assign N3660 = N3659 & N1941;
  assign N3659 = N2150 & en_i;
  assign empty_array[377] = N3661 & N3662;
  assign N3661 = N2150 & en_i;
  assign N3662 = ~valid[377];
  assign match_array[378] = N3664 & valid[378];
  assign N3664 = N3663 & N1942;
  assign N3663 = N2150 & en_i;
  assign empty_array[378] = N3665 & N3666;
  assign N3665 = N2150 & en_i;
  assign N3666 = ~valid[378];
  assign match_array[379] = N3668 & valid[379];
  assign N3668 = N3667 & N1943;
  assign N3667 = N2150 & en_i;
  assign empty_array[379] = N3669 & N3670;
  assign N3669 = N2150 & en_i;
  assign N3670 = ~valid[379];
  assign match_array[380] = N3672 & valid[380];
  assign N3672 = N3671 & N1944;
  assign N3671 = N2150 & en_i;
  assign empty_array[380] = N3673 & N3674;
  assign N3673 = N2150 & en_i;
  assign N3674 = ~valid[380];
  assign match_array[381] = N3676 & valid[381];
  assign N3676 = N3675 & N1945;
  assign N3675 = N2150 & en_i;
  assign empty_array[381] = N3677 & N3678;
  assign N3677 = N2150 & en_i;
  assign N3678 = ~valid[381];
  assign match_array[382] = N3680 & valid[382];
  assign N3680 = N3679 & N1946;
  assign N3679 = N2150 & en_i;
  assign empty_array[382] = N3681 & N3682;
  assign N3681 = N2150 & en_i;
  assign N3682 = ~valid[382];
  assign match_array[383] = N3684 & valid[383];
  assign N3684 = N3683 & N1947;
  assign N3683 = N2150 & en_i;
  assign empty_array[383] = N3685 & N3686;
  assign N3685 = N2150 & en_i;
  assign N3686 = ~valid[383];
  assign match_array[384] = N3688 & valid[384];
  assign N3688 = N3687 & N1948;
  assign N3687 = N2150 & en_i;
  assign empty_array[384] = N3689 & N3690;
  assign N3689 = N2150 & en_i;
  assign N3690 = ~valid[384];
  assign match_array[385] = N3692 & valid[385];
  assign N3692 = N3691 & N1949;
  assign N3691 = N2150 & en_i;
  assign empty_array[385] = N3693 & N3694;
  assign N3693 = N2150 & en_i;
  assign N3694 = ~valid[385];
  assign match_array[386] = N3696 & valid[386];
  assign N3696 = N3695 & N1950;
  assign N3695 = N2150 & en_i;
  assign empty_array[386] = N3697 & N3698;
  assign N3697 = N2150 & en_i;
  assign N3698 = ~valid[386];
  assign match_array[387] = N3700 & valid[387];
  assign N3700 = N3699 & N1951;
  assign N3699 = N2150 & en_i;
  assign empty_array[387] = N3701 & N3702;
  assign N3701 = N2150 & en_i;
  assign N3702 = ~valid[387];
  assign match_array[388] = N3704 & valid[388];
  assign N3704 = N3703 & N1952;
  assign N3703 = N2150 & en_i;
  assign empty_array[388] = N3705 & N3706;
  assign N3705 = N2150 & en_i;
  assign N3706 = ~valid[388];
  assign match_array[389] = N3708 & valid[389];
  assign N3708 = N3707 & N1953;
  assign N3707 = N2150 & en_i;
  assign empty_array[389] = N3709 & N3710;
  assign N3709 = N2150 & en_i;
  assign N3710 = ~valid[389];
  assign match_array[390] = N3712 & valid[390];
  assign N3712 = N3711 & N1954;
  assign N3711 = N2150 & en_i;
  assign empty_array[390] = N3713 & N3714;
  assign N3713 = N2150 & en_i;
  assign N3714 = ~valid[390];
  assign match_array[391] = N3716 & valid[391];
  assign N3716 = N3715 & N1955;
  assign N3715 = N2150 & en_i;
  assign empty_array[391] = N3717 & N3718;
  assign N3717 = N2150 & en_i;
  assign N3718 = ~valid[391];
  assign match_array[392] = N3720 & valid[392];
  assign N3720 = N3719 & N1956;
  assign N3719 = N2150 & en_i;
  assign empty_array[392] = N3721 & N3722;
  assign N3721 = N2150 & en_i;
  assign N3722 = ~valid[392];
  assign match_array[393] = N3724 & valid[393];
  assign N3724 = N3723 & N1957;
  assign N3723 = N2150 & en_i;
  assign empty_array[393] = N3725 & N3726;
  assign N3725 = N2150 & en_i;
  assign N3726 = ~valid[393];
  assign match_array[394] = N3728 & valid[394];
  assign N3728 = N3727 & N1958;
  assign N3727 = N2150 & en_i;
  assign empty_array[394] = N3729 & N3730;
  assign N3729 = N2150 & en_i;
  assign N3730 = ~valid[394];
  assign match_array[395] = N3732 & valid[395];
  assign N3732 = N3731 & N1959;
  assign N3731 = N2150 & en_i;
  assign empty_array[395] = N3733 & N3734;
  assign N3733 = N2150 & en_i;
  assign N3734 = ~valid[395];
  assign match_array[396] = N3736 & valid[396];
  assign N3736 = N3735 & N1960;
  assign N3735 = N2150 & en_i;
  assign empty_array[396] = N3737 & N3738;
  assign N3737 = N2150 & en_i;
  assign N3738 = ~valid[396];
  assign match_array[397] = N3740 & valid[397];
  assign N3740 = N3739 & N1961;
  assign N3739 = N2150 & en_i;
  assign empty_array[397] = N3741 & N3742;
  assign N3741 = N2150 & en_i;
  assign N3742 = ~valid[397];
  assign match_array[398] = N3744 & valid[398];
  assign N3744 = N3743 & N1962;
  assign N3743 = N2150 & en_i;
  assign empty_array[398] = N3745 & N3746;
  assign N3745 = N2150 & en_i;
  assign N3746 = ~valid[398];
  assign match_array[399] = N3748 & valid[399];
  assign N3748 = N3747 & N1963;
  assign N3747 = N2150 & en_i;
  assign empty_array[399] = N3749 & N3750;
  assign N3749 = N2150 & en_i;
  assign N3750 = ~valid[399];
  assign match_array[400] = N3752 & valid[400];
  assign N3752 = N3751 & N1964;
  assign N3751 = N2150 & en_i;
  assign empty_array[400] = N3753 & N3754;
  assign N3753 = N2150 & en_i;
  assign N3754 = ~valid[400];
  assign match_array[401] = N3756 & valid[401];
  assign N3756 = N3755 & N1965;
  assign N3755 = N2150 & en_i;
  assign empty_array[401] = N3757 & N3758;
  assign N3757 = N2150 & en_i;
  assign N3758 = ~valid[401];
  assign match_array[402] = N3760 & valid[402];
  assign N3760 = N3759 & N1966;
  assign N3759 = N2150 & en_i;
  assign empty_array[402] = N3761 & N3762;
  assign N3761 = N2150 & en_i;
  assign N3762 = ~valid[402];
  assign match_array[403] = N3764 & valid[403];
  assign N3764 = N3763 & N1967;
  assign N3763 = N2150 & en_i;
  assign empty_array[403] = N3765 & N3766;
  assign N3765 = N2150 & en_i;
  assign N3766 = ~valid[403];
  assign match_array[404] = N3768 & valid[404];
  assign N3768 = N3767 & N1968;
  assign N3767 = N2150 & en_i;
  assign empty_array[404] = N3769 & N3770;
  assign N3769 = N2150 & en_i;
  assign N3770 = ~valid[404];
  assign match_array[405] = N3772 & valid[405];
  assign N3772 = N3771 & N1969;
  assign N3771 = N2150 & en_i;
  assign empty_array[405] = N3773 & N3774;
  assign N3773 = N2150 & en_i;
  assign N3774 = ~valid[405];
  assign match_array[406] = N3776 & valid[406];
  assign N3776 = N3775 & N1970;
  assign N3775 = N2150 & en_i;
  assign empty_array[406] = N3777 & N3778;
  assign N3777 = N2150 & en_i;
  assign N3778 = ~valid[406];
  assign match_array[407] = N3780 & valid[407];
  assign N3780 = N3779 & N1971;
  assign N3779 = N2150 & en_i;
  assign empty_array[407] = N3781 & N3782;
  assign N3781 = N2150 & en_i;
  assign N3782 = ~valid[407];
  assign match_array[408] = N3784 & valid[408];
  assign N3784 = N3783 & N1972;
  assign N3783 = N2150 & en_i;
  assign empty_array[408] = N3785 & N3786;
  assign N3785 = N2150 & en_i;
  assign N3786 = ~valid[408];
  assign match_array[409] = N3788 & valid[409];
  assign N3788 = N3787 & N1973;
  assign N3787 = N2150 & en_i;
  assign empty_array[409] = N3789 & N3790;
  assign N3789 = N2150 & en_i;
  assign N3790 = ~valid[409];
  assign match_array[410] = N3792 & valid[410];
  assign N3792 = N3791 & N1974;
  assign N3791 = N2150 & en_i;
  assign empty_array[410] = N3793 & N3794;
  assign N3793 = N2150 & en_i;
  assign N3794 = ~valid[410];
  assign match_array[411] = N3796 & valid[411];
  assign N3796 = N3795 & N1975;
  assign N3795 = N2150 & en_i;
  assign empty_array[411] = N3797 & N3798;
  assign N3797 = N2150 & en_i;
  assign N3798 = ~valid[411];
  assign match_array[412] = N3800 & valid[412];
  assign N3800 = N3799 & N1976;
  assign N3799 = N2150 & en_i;
  assign empty_array[412] = N3801 & N3802;
  assign N3801 = N2150 & en_i;
  assign N3802 = ~valid[412];
  assign match_array[413] = N3804 & valid[413];
  assign N3804 = N3803 & N1977;
  assign N3803 = N2150 & en_i;
  assign empty_array[413] = N3805 & N3806;
  assign N3805 = N2150 & en_i;
  assign N3806 = ~valid[413];
  assign match_array[414] = N3808 & valid[414];
  assign N3808 = N3807 & N1978;
  assign N3807 = N2150 & en_i;
  assign empty_array[414] = N3809 & N3810;
  assign N3809 = N2150 & en_i;
  assign N3810 = ~valid[414];
  assign match_array[415] = N3812 & valid[415];
  assign N3812 = N3811 & N1979;
  assign N3811 = N2150 & en_i;
  assign empty_array[415] = N3813 & N3814;
  assign N3813 = N2150 & en_i;
  assign N3814 = ~valid[415];
  assign match_array[416] = N3816 & valid[416];
  assign N3816 = N3815 & N1980;
  assign N3815 = N2150 & en_i;
  assign empty_array[416] = N3817 & N3818;
  assign N3817 = N2150 & en_i;
  assign N3818 = ~valid[416];
  assign match_array[417] = N3820 & valid[417];
  assign N3820 = N3819 & N1981;
  assign N3819 = N2150 & en_i;
  assign empty_array[417] = N3821 & N3822;
  assign N3821 = N2150 & en_i;
  assign N3822 = ~valid[417];
  assign match_array[418] = N3824 & valid[418];
  assign N3824 = N3823 & N1982;
  assign N3823 = N2150 & en_i;
  assign empty_array[418] = N3825 & N3826;
  assign N3825 = N2150 & en_i;
  assign N3826 = ~valid[418];
  assign match_array[419] = N3828 & valid[419];
  assign N3828 = N3827 & N1983;
  assign N3827 = N2150 & en_i;
  assign empty_array[419] = N3829 & N3830;
  assign N3829 = N2150 & en_i;
  assign N3830 = ~valid[419];
  assign match_array[420] = N3832 & valid[420];
  assign N3832 = N3831 & N1984;
  assign N3831 = N2150 & en_i;
  assign empty_array[420] = N3833 & N3834;
  assign N3833 = N2150 & en_i;
  assign N3834 = ~valid[420];
  assign match_array[421] = N3836 & valid[421];
  assign N3836 = N3835 & N1985;
  assign N3835 = N2150 & en_i;
  assign empty_array[421] = N3837 & N3838;
  assign N3837 = N2150 & en_i;
  assign N3838 = ~valid[421];
  assign match_array[422] = N3840 & valid[422];
  assign N3840 = N3839 & N1986;
  assign N3839 = N2150 & en_i;
  assign empty_array[422] = N3841 & N3842;
  assign N3841 = N2150 & en_i;
  assign N3842 = ~valid[422];
  assign match_array[423] = N3844 & valid[423];
  assign N3844 = N3843 & N1987;
  assign N3843 = N2150 & en_i;
  assign empty_array[423] = N3845 & N3846;
  assign N3845 = N2150 & en_i;
  assign N3846 = ~valid[423];
  assign match_array[424] = N3848 & valid[424];
  assign N3848 = N3847 & N1988;
  assign N3847 = N2150 & en_i;
  assign empty_array[424] = N3849 & N3850;
  assign N3849 = N2150 & en_i;
  assign N3850 = ~valid[424];
  assign match_array[425] = N3852 & valid[425];
  assign N3852 = N3851 & N1989;
  assign N3851 = N2150 & en_i;
  assign empty_array[425] = N3853 & N3854;
  assign N3853 = N2150 & en_i;
  assign N3854 = ~valid[425];
  assign match_array[426] = N3856 & valid[426];
  assign N3856 = N3855 & N1990;
  assign N3855 = N2150 & en_i;
  assign empty_array[426] = N3857 & N3858;
  assign N3857 = N2150 & en_i;
  assign N3858 = ~valid[426];
  assign match_array[427] = N3860 & valid[427];
  assign N3860 = N3859 & N1991;
  assign N3859 = N2150 & en_i;
  assign empty_array[427] = N3861 & N3862;
  assign N3861 = N2150 & en_i;
  assign N3862 = ~valid[427];
  assign match_array[428] = N3864 & valid[428];
  assign N3864 = N3863 & N1992;
  assign N3863 = N2150 & en_i;
  assign empty_array[428] = N3865 & N3866;
  assign N3865 = N2150 & en_i;
  assign N3866 = ~valid[428];
  assign match_array[429] = N3868 & valid[429];
  assign N3868 = N3867 & N1993;
  assign N3867 = N2150 & en_i;
  assign empty_array[429] = N3869 & N3870;
  assign N3869 = N2150 & en_i;
  assign N3870 = ~valid[429];
  assign match_array[430] = N3872 & valid[430];
  assign N3872 = N3871 & N1994;
  assign N3871 = N2150 & en_i;
  assign empty_array[430] = N3873 & N3874;
  assign N3873 = N2150 & en_i;
  assign N3874 = ~valid[430];
  assign match_array[431] = N3876 & valid[431];
  assign N3876 = N3875 & N1995;
  assign N3875 = N2150 & en_i;
  assign empty_array[431] = N3877 & N3878;
  assign N3877 = N2150 & en_i;
  assign N3878 = ~valid[431];
  assign match_array[432] = N3880 & valid[432];
  assign N3880 = N3879 & N1996;
  assign N3879 = N2150 & en_i;
  assign empty_array[432] = N3881 & N3882;
  assign N3881 = N2150 & en_i;
  assign N3882 = ~valid[432];
  assign match_array[433] = N3884 & valid[433];
  assign N3884 = N3883 & N1997;
  assign N3883 = N2150 & en_i;
  assign empty_array[433] = N3885 & N3886;
  assign N3885 = N2150 & en_i;
  assign N3886 = ~valid[433];
  assign match_array[434] = N3888 & valid[434];
  assign N3888 = N3887 & N1998;
  assign N3887 = N2150 & en_i;
  assign empty_array[434] = N3889 & N3890;
  assign N3889 = N2150 & en_i;
  assign N3890 = ~valid[434];
  assign match_array[435] = N3892 & valid[435];
  assign N3892 = N3891 & N1999;
  assign N3891 = N2150 & en_i;
  assign empty_array[435] = N3893 & N3894;
  assign N3893 = N2150 & en_i;
  assign N3894 = ~valid[435];
  assign match_array[436] = N3896 & valid[436];
  assign N3896 = N3895 & N2000;
  assign N3895 = N2150 & en_i;
  assign empty_array[436] = N3897 & N3898;
  assign N3897 = N2150 & en_i;
  assign N3898 = ~valid[436];
  assign match_array[437] = N3900 & valid[437];
  assign N3900 = N3899 & N2001;
  assign N3899 = N2150 & en_i;
  assign empty_array[437] = N3901 & N3902;
  assign N3901 = N2150 & en_i;
  assign N3902 = ~valid[437];
  assign match_array[438] = N3904 & valid[438];
  assign N3904 = N3903 & N2002;
  assign N3903 = N2150 & en_i;
  assign empty_array[438] = N3905 & N3906;
  assign N3905 = N2150 & en_i;
  assign N3906 = ~valid[438];
  assign match_array[439] = N3908 & valid[439];
  assign N3908 = N3907 & N2003;
  assign N3907 = N2150 & en_i;
  assign empty_array[439] = N3909 & N3910;
  assign N3909 = N2150 & en_i;
  assign N3910 = ~valid[439];
  assign match_array[440] = N3912 & valid[440];
  assign N3912 = N3911 & N2004;
  assign N3911 = N2150 & en_i;
  assign empty_array[440] = N3913 & N3914;
  assign N3913 = N2150 & en_i;
  assign N3914 = ~valid[440];
  assign match_array[441] = N3916 & valid[441];
  assign N3916 = N3915 & N2005;
  assign N3915 = N2150 & en_i;
  assign empty_array[441] = N3917 & N3918;
  assign N3917 = N2150 & en_i;
  assign N3918 = ~valid[441];
  assign match_array[442] = N3920 & valid[442];
  assign N3920 = N3919 & N2006;
  assign N3919 = N2150 & en_i;
  assign empty_array[442] = N3921 & N3922;
  assign N3921 = N2150 & en_i;
  assign N3922 = ~valid[442];
  assign match_array[443] = N3924 & valid[443];
  assign N3924 = N3923 & N2007;
  assign N3923 = N2150 & en_i;
  assign empty_array[443] = N3925 & N3926;
  assign N3925 = N2150 & en_i;
  assign N3926 = ~valid[443];
  assign match_array[444] = N3928 & valid[444];
  assign N3928 = N3927 & N2008;
  assign N3927 = N2150 & en_i;
  assign empty_array[444] = N3929 & N3930;
  assign N3929 = N2150 & en_i;
  assign N3930 = ~valid[444];
  assign match_array[445] = N3932 & valid[445];
  assign N3932 = N3931 & N2009;
  assign N3931 = N2150 & en_i;
  assign empty_array[445] = N3933 & N3934;
  assign N3933 = N2150 & en_i;
  assign N3934 = ~valid[445];
  assign match_array[446] = N3936 & valid[446];
  assign N3936 = N3935 & N2010;
  assign N3935 = N2150 & en_i;
  assign empty_array[446] = N3937 & N3938;
  assign N3937 = N2150 & en_i;
  assign N3938 = ~valid[446];
  assign match_array[447] = N3940 & valid[447];
  assign N3940 = N3939 & N2011;
  assign N3939 = N2150 & en_i;
  assign empty_array[447] = N3941 & N3942;
  assign N3941 = N2150 & en_i;
  assign N3942 = ~valid[447];
  assign match_array[448] = N3944 & valid[448];
  assign N3944 = N3943 & N2012;
  assign N3943 = N2150 & en_i;
  assign empty_array[448] = N3945 & N3946;
  assign N3945 = N2150 & en_i;
  assign N3946 = ~valid[448];
  assign match_array[449] = N3948 & valid[449];
  assign N3948 = N3947 & N2013;
  assign N3947 = N2150 & en_i;
  assign empty_array[449] = N3949 & N3950;
  assign N3949 = N2150 & en_i;
  assign N3950 = ~valid[449];
  assign match_array[450] = N3952 & valid[450];
  assign N3952 = N3951 & N2014;
  assign N3951 = N2150 & en_i;
  assign empty_array[450] = N3953 & N3954;
  assign N3953 = N2150 & en_i;
  assign N3954 = ~valid[450];
  assign match_array[451] = N3956 & valid[451];
  assign N3956 = N3955 & N2015;
  assign N3955 = N2150 & en_i;
  assign empty_array[451] = N3957 & N3958;
  assign N3957 = N2150 & en_i;
  assign N3958 = ~valid[451];
  assign match_array[452] = N3960 & valid[452];
  assign N3960 = N3959 & N2016;
  assign N3959 = N2150 & en_i;
  assign empty_array[452] = N3961 & N3962;
  assign N3961 = N2150 & en_i;
  assign N3962 = ~valid[452];
  assign match_array[453] = N3964 & valid[453];
  assign N3964 = N3963 & N2017;
  assign N3963 = N2150 & en_i;
  assign empty_array[453] = N3965 & N3966;
  assign N3965 = N2150 & en_i;
  assign N3966 = ~valid[453];
  assign match_array[454] = N3968 & valid[454];
  assign N3968 = N3967 & N2018;
  assign N3967 = N2150 & en_i;
  assign empty_array[454] = N3969 & N3970;
  assign N3969 = N2150 & en_i;
  assign N3970 = ~valid[454];
  assign match_array[455] = N3972 & valid[455];
  assign N3972 = N3971 & N2019;
  assign N3971 = N2150 & en_i;
  assign empty_array[455] = N3973 & N3974;
  assign N3973 = N2150 & en_i;
  assign N3974 = ~valid[455];
  assign match_array[456] = N3976 & valid[456];
  assign N3976 = N3975 & N2020;
  assign N3975 = N2150 & en_i;
  assign empty_array[456] = N3977 & N3978;
  assign N3977 = N2150 & en_i;
  assign N3978 = ~valid[456];
  assign match_array[457] = N3980 & valid[457];
  assign N3980 = N3979 & N2021;
  assign N3979 = N2150 & en_i;
  assign empty_array[457] = N3981 & N3982;
  assign N3981 = N2150 & en_i;
  assign N3982 = ~valid[457];
  assign match_array[458] = N3984 & valid[458];
  assign N3984 = N3983 & N2022;
  assign N3983 = N2150 & en_i;
  assign empty_array[458] = N3985 & N3986;
  assign N3985 = N2150 & en_i;
  assign N3986 = ~valid[458];
  assign match_array[459] = N3988 & valid[459];
  assign N3988 = N3987 & N2023;
  assign N3987 = N2150 & en_i;
  assign empty_array[459] = N3989 & N3990;
  assign N3989 = N2150 & en_i;
  assign N3990 = ~valid[459];
  assign match_array[460] = N3992 & valid[460];
  assign N3992 = N3991 & N2024;
  assign N3991 = N2150 & en_i;
  assign empty_array[460] = N3993 & N3994;
  assign N3993 = N2150 & en_i;
  assign N3994 = ~valid[460];
  assign match_array[461] = N3996 & valid[461];
  assign N3996 = N3995 & N2025;
  assign N3995 = N2150 & en_i;
  assign empty_array[461] = N3997 & N3998;
  assign N3997 = N2150 & en_i;
  assign N3998 = ~valid[461];
  assign match_array[462] = N4000 & valid[462];
  assign N4000 = N3999 & N2026;
  assign N3999 = N2150 & en_i;
  assign empty_array[462] = N4001 & N4002;
  assign N4001 = N2150 & en_i;
  assign N4002 = ~valid[462];
  assign match_array[463] = N4004 & valid[463];
  assign N4004 = N4003 & N2027;
  assign N4003 = N2150 & en_i;
  assign empty_array[463] = N4005 & N4006;
  assign N4005 = N2150 & en_i;
  assign N4006 = ~valid[463];
  assign match_array[464] = N4008 & valid[464];
  assign N4008 = N4007 & N2028;
  assign N4007 = N2150 & en_i;
  assign empty_array[464] = N4009 & N4010;
  assign N4009 = N2150 & en_i;
  assign N4010 = ~valid[464];
  assign match_array[465] = N4012 & valid[465];
  assign N4012 = N4011 & N2029;
  assign N4011 = N2150 & en_i;
  assign empty_array[465] = N4013 & N4014;
  assign N4013 = N2150 & en_i;
  assign N4014 = ~valid[465];
  assign match_array[466] = N4016 & valid[466];
  assign N4016 = N4015 & N2030;
  assign N4015 = N2150 & en_i;
  assign empty_array[466] = N4017 & N4018;
  assign N4017 = N2150 & en_i;
  assign N4018 = ~valid[466];
  assign match_array[467] = N4020 & valid[467];
  assign N4020 = N4019 & N2031;
  assign N4019 = N2150 & en_i;
  assign empty_array[467] = N4021 & N4022;
  assign N4021 = N2150 & en_i;
  assign N4022 = ~valid[467];
  assign match_array[468] = N4024 & valid[468];
  assign N4024 = N4023 & N2032;
  assign N4023 = N2150 & en_i;
  assign empty_array[468] = N4025 & N4026;
  assign N4025 = N2150 & en_i;
  assign N4026 = ~valid[468];
  assign match_array[469] = N4028 & valid[469];
  assign N4028 = N4027 & N2033;
  assign N4027 = N2150 & en_i;
  assign empty_array[469] = N4029 & N4030;
  assign N4029 = N2150 & en_i;
  assign N4030 = ~valid[469];
  assign match_array[470] = N4032 & valid[470];
  assign N4032 = N4031 & N2034;
  assign N4031 = N2150 & en_i;
  assign empty_array[470] = N4033 & N4034;
  assign N4033 = N2150 & en_i;
  assign N4034 = ~valid[470];
  assign match_array[471] = N4036 & valid[471];
  assign N4036 = N4035 & N2035;
  assign N4035 = N2150 & en_i;
  assign empty_array[471] = N4037 & N4038;
  assign N4037 = N2150 & en_i;
  assign N4038 = ~valid[471];
  assign match_array[472] = N4040 & valid[472];
  assign N4040 = N4039 & N2036;
  assign N4039 = N2150 & en_i;
  assign empty_array[472] = N4041 & N4042;
  assign N4041 = N2150 & en_i;
  assign N4042 = ~valid[472];
  assign match_array[473] = N4044 & valid[473];
  assign N4044 = N4043 & N2037;
  assign N4043 = N2150 & en_i;
  assign empty_array[473] = N4045 & N4046;
  assign N4045 = N2150 & en_i;
  assign N4046 = ~valid[473];
  assign match_array[474] = N4048 & valid[474];
  assign N4048 = N4047 & N2038;
  assign N4047 = N2150 & en_i;
  assign empty_array[474] = N4049 & N4050;
  assign N4049 = N2150 & en_i;
  assign N4050 = ~valid[474];
  assign match_array[475] = N4052 & valid[475];
  assign N4052 = N4051 & N2039;
  assign N4051 = N2150 & en_i;
  assign empty_array[475] = N4053 & N4054;
  assign N4053 = N2150 & en_i;
  assign N4054 = ~valid[475];
  assign match_array[476] = N4056 & valid[476];
  assign N4056 = N4055 & N2040;
  assign N4055 = N2150 & en_i;
  assign empty_array[476] = N4057 & N4058;
  assign N4057 = N2150 & en_i;
  assign N4058 = ~valid[476];
  assign match_array[477] = N4060 & valid[477];
  assign N4060 = N4059 & N2041;
  assign N4059 = N2150 & en_i;
  assign empty_array[477] = N4061 & N4062;
  assign N4061 = N2150 & en_i;
  assign N4062 = ~valid[477];
  assign match_array[478] = N4064 & valid[478];
  assign N4064 = N4063 & N2042;
  assign N4063 = N2150 & en_i;
  assign empty_array[478] = N4065 & N4066;
  assign N4065 = N2150 & en_i;
  assign N4066 = ~valid[478];
  assign match_array[479] = N4068 & valid[479];
  assign N4068 = N4067 & N2043;
  assign N4067 = N2150 & en_i;
  assign empty_array[479] = N4069 & N4070;
  assign N4069 = N2150 & en_i;
  assign N4070 = ~valid[479];
  assign match_array[480] = N4072 & valid[480];
  assign N4072 = N4071 & N2044;
  assign N4071 = N2150 & en_i;
  assign empty_array[480] = N4073 & N4074;
  assign N4073 = N2150 & en_i;
  assign N4074 = ~valid[480];
  assign match_array[481] = N4076 & valid[481];
  assign N4076 = N4075 & N2045;
  assign N4075 = N2150 & en_i;
  assign empty_array[481] = N4077 & N4078;
  assign N4077 = N2150 & en_i;
  assign N4078 = ~valid[481];
  assign match_array[482] = N4080 & valid[482];
  assign N4080 = N4079 & N2046;
  assign N4079 = N2150 & en_i;
  assign empty_array[482] = N4081 & N4082;
  assign N4081 = N2150 & en_i;
  assign N4082 = ~valid[482];
  assign match_array[483] = N4084 & valid[483];
  assign N4084 = N4083 & N2047;
  assign N4083 = N2150 & en_i;
  assign empty_array[483] = N4085 & N4086;
  assign N4085 = N2150 & en_i;
  assign N4086 = ~valid[483];
  assign match_array[484] = N4088 & valid[484];
  assign N4088 = N4087 & N2048;
  assign N4087 = N2150 & en_i;
  assign empty_array[484] = N4089 & N4090;
  assign N4089 = N2150 & en_i;
  assign N4090 = ~valid[484];
  assign match_array[485] = N4092 & valid[485];
  assign N4092 = N4091 & N2049;
  assign N4091 = N2150 & en_i;
  assign empty_array[485] = N4093 & N4094;
  assign N4093 = N2150 & en_i;
  assign N4094 = ~valid[485];
  assign match_array[486] = N4096 & valid[486];
  assign N4096 = N4095 & N2050;
  assign N4095 = N2150 & en_i;
  assign empty_array[486] = N4097 & N4098;
  assign N4097 = N2150 & en_i;
  assign N4098 = ~valid[486];
  assign match_array[487] = N4100 & valid[487];
  assign N4100 = N4099 & N2051;
  assign N4099 = N2150 & en_i;
  assign empty_array[487] = N4101 & N4102;
  assign N4101 = N2150 & en_i;
  assign N4102 = ~valid[487];
  assign match_array[488] = N4104 & valid[488];
  assign N4104 = N4103 & N2052;
  assign N4103 = N2150 & en_i;
  assign empty_array[488] = N4105 & N4106;
  assign N4105 = N2150 & en_i;
  assign N4106 = ~valid[488];
  assign match_array[489] = N4108 & valid[489];
  assign N4108 = N4107 & N2053;
  assign N4107 = N2150 & en_i;
  assign empty_array[489] = N4109 & N4110;
  assign N4109 = N2150 & en_i;
  assign N4110 = ~valid[489];
  assign match_array[490] = N4112 & valid[490];
  assign N4112 = N4111 & N2054;
  assign N4111 = N2150 & en_i;
  assign empty_array[490] = N4113 & N4114;
  assign N4113 = N2150 & en_i;
  assign N4114 = ~valid[490];
  assign match_array[491] = N4116 & valid[491];
  assign N4116 = N4115 & N2055;
  assign N4115 = N2150 & en_i;
  assign empty_array[491] = N4117 & N4118;
  assign N4117 = N2150 & en_i;
  assign N4118 = ~valid[491];
  assign match_array[492] = N4120 & valid[492];
  assign N4120 = N4119 & N2056;
  assign N4119 = N2150 & en_i;
  assign empty_array[492] = N4121 & N4122;
  assign N4121 = N2150 & en_i;
  assign N4122 = ~valid[492];
  assign match_array[493] = N4124 & valid[493];
  assign N4124 = N4123 & N2057;
  assign N4123 = N2150 & en_i;
  assign empty_array[493] = N4125 & N4126;
  assign N4125 = N2150 & en_i;
  assign N4126 = ~valid[493];
  assign match_array[494] = N4128 & valid[494];
  assign N4128 = N4127 & N2058;
  assign N4127 = N2150 & en_i;
  assign empty_array[494] = N4129 & N4130;
  assign N4129 = N2150 & en_i;
  assign N4130 = ~valid[494];
  assign match_array[495] = N4132 & valid[495];
  assign N4132 = N4131 & N2059;
  assign N4131 = N2150 & en_i;
  assign empty_array[495] = N4133 & N4134;
  assign N4133 = N2150 & en_i;
  assign N4134 = ~valid[495];
  assign match_array[496] = N4136 & valid[496];
  assign N4136 = N4135 & N2060;
  assign N4135 = N2150 & en_i;
  assign empty_array[496] = N4137 & N4138;
  assign N4137 = N2150 & en_i;
  assign N4138 = ~valid[496];
  assign match_array[497] = N4140 & valid[497];
  assign N4140 = N4139 & N2061;
  assign N4139 = N2150 & en_i;
  assign empty_array[497] = N4141 & N4142;
  assign N4141 = N2150 & en_i;
  assign N4142 = ~valid[497];
  assign match_array[498] = N4144 & valid[498];
  assign N4144 = N4143 & N2062;
  assign N4143 = N2150 & en_i;
  assign empty_array[498] = N4145 & N4146;
  assign N4145 = N2150 & en_i;
  assign N4146 = ~valid[498];
  assign match_array[499] = N4148 & valid[499];
  assign N4148 = N4147 & N2063;
  assign N4147 = N2150 & en_i;
  assign empty_array[499] = N4149 & N4150;
  assign N4149 = N2150 & en_i;
  assign N4150 = ~valid[499];
  assign match_array[500] = N4152 & valid[500];
  assign N4152 = N4151 & N2064;
  assign N4151 = N2150 & en_i;
  assign empty_array[500] = N4153 & N4154;
  assign N4153 = N2150 & en_i;
  assign N4154 = ~valid[500];
  assign match_array[501] = N4156 & valid[501];
  assign N4156 = N4155 & N2065;
  assign N4155 = N2150 & en_i;
  assign empty_array[501] = N4157 & N4158;
  assign N4157 = N2150 & en_i;
  assign N4158 = ~valid[501];
  assign match_array[502] = N4160 & valid[502];
  assign N4160 = N4159 & N2066;
  assign N4159 = N2150 & en_i;
  assign empty_array[502] = N4161 & N4162;
  assign N4161 = N2150 & en_i;
  assign N4162 = ~valid[502];
  assign match_array[503] = N4164 & valid[503];
  assign N4164 = N4163 & N2067;
  assign N4163 = N2150 & en_i;
  assign empty_array[503] = N4165 & N4166;
  assign N4165 = N2150 & en_i;
  assign N4166 = ~valid[503];
  assign match_array[504] = N4168 & valid[504];
  assign N4168 = N4167 & N2068;
  assign N4167 = N2150 & en_i;
  assign empty_array[504] = N4169 & N4170;
  assign N4169 = N2150 & en_i;
  assign N4170 = ~valid[504];
  assign match_array[505] = N4172 & valid[505];
  assign N4172 = N4171 & N2069;
  assign N4171 = N2150 & en_i;
  assign empty_array[505] = N4173 & N4174;
  assign N4173 = N2150 & en_i;
  assign N4174 = ~valid[505];
  assign match_array[506] = N4176 & valid[506];
  assign N4176 = N4175 & N2070;
  assign N4175 = N2150 & en_i;
  assign empty_array[506] = N4177 & N4178;
  assign N4177 = N2150 & en_i;
  assign N4178 = ~valid[506];
  assign match_array[507] = N4180 & valid[507];
  assign N4180 = N4179 & N2071;
  assign N4179 = N2150 & en_i;
  assign empty_array[507] = N4181 & N4182;
  assign N4181 = N2150 & en_i;
  assign N4182 = ~valid[507];
  assign match_array[508] = N4184 & valid[508];
  assign N4184 = N4183 & N2072;
  assign N4183 = N2150 & en_i;
  assign empty_array[508] = N4185 & N4186;
  assign N4185 = N2150 & en_i;
  assign N4186 = ~valid[508];
  assign match_array[509] = N4188 & valid[509];
  assign N4188 = N4187 & N2073;
  assign N4187 = N2150 & en_i;
  assign empty_array[509] = N4189 & N4190;
  assign N4189 = N2150 & en_i;
  assign N4190 = ~valid[509];
  assign match_array[510] = N4192 & valid[510];
  assign N4192 = N4191 & N2074;
  assign N4191 = N2150 & en_i;
  assign empty_array[510] = N4193 & N4194;
  assign N4193 = N2150 & en_i;
  assign N4194 = ~valid[510];
  assign match_array[511] = N4196 & valid[511];
  assign N4196 = N4195 & N2075;
  assign N4195 = N2150 & en_i;
  assign empty_array[511] = N4197 & N4198;
  assign N4197 = N2150 & en_i;
  assign N4198 = ~valid[511];

  always @(posedge clk_i) begin
    if(N1561) begin
      { mem[8191:8176] } <= { w_data_i[15:0] };
    end 
    if(N1560) begin
      { mem[8175:8160] } <= { w_data_i[15:0] };
    end 
    if(N1559) begin
      { mem[8159:8144] } <= { w_data_i[15:0] };
    end 
    if(N1558) begin
      { mem[8143:8128] } <= { w_data_i[15:0] };
    end 
    if(N1557) begin
      { mem[8127:8112] } <= { w_data_i[15:0] };
    end 
    if(N1556) begin
      { mem[8111:8096] } <= { w_data_i[15:0] };
    end 
    if(N1555) begin
      { mem[8095:8080] } <= { w_data_i[15:0] };
    end 
    if(N1554) begin
      { mem[8079:8064] } <= { w_data_i[15:0] };
    end 
    if(N1553) begin
      { mem[8063:8048] } <= { w_data_i[15:0] };
    end 
    if(N1552) begin
      { mem[8047:8032] } <= { w_data_i[15:0] };
    end 
    if(N1551) begin
      { mem[8031:8016] } <= { w_data_i[15:0] };
    end 
    if(N1550) begin
      { mem[8015:8000] } <= { w_data_i[15:0] };
    end 
    if(N1549) begin
      { mem[7999:7984] } <= { w_data_i[15:0] };
    end 
    if(N1548) begin
      { mem[7983:7968] } <= { w_data_i[15:0] };
    end 
    if(N1547) begin
      { mem[7967:7952] } <= { w_data_i[15:0] };
    end 
    if(N1546) begin
      { mem[7951:7936] } <= { w_data_i[15:0] };
    end 
    if(N1545) begin
      { mem[7935:7920] } <= { w_data_i[15:0] };
    end 
    if(N1544) begin
      { mem[7919:7904] } <= { w_data_i[15:0] };
    end 
    if(N1543) begin
      { mem[7903:7888] } <= { w_data_i[15:0] };
    end 
    if(N1542) begin
      { mem[7887:7872] } <= { w_data_i[15:0] };
    end 
    if(N1541) begin
      { mem[7871:7856] } <= { w_data_i[15:0] };
    end 
    if(N1540) begin
      { mem[7855:7840] } <= { w_data_i[15:0] };
    end 
    if(N1539) begin
      { mem[7839:7824] } <= { w_data_i[15:0] };
    end 
    if(N1538) begin
      { mem[7823:7808] } <= { w_data_i[15:0] };
    end 
    if(N1537) begin
      { mem[7807:7792] } <= { w_data_i[15:0] };
    end 
    if(N1536) begin
      { mem[7791:7776] } <= { w_data_i[15:0] };
    end 
    if(N1535) begin
      { mem[7775:7760] } <= { w_data_i[15:0] };
    end 
    if(N1534) begin
      { mem[7759:7744] } <= { w_data_i[15:0] };
    end 
    if(N1533) begin
      { mem[7743:7728] } <= { w_data_i[15:0] };
    end 
    if(N1532) begin
      { mem[7727:7712] } <= { w_data_i[15:0] };
    end 
    if(N1531) begin
      { mem[7711:7696] } <= { w_data_i[15:0] };
    end 
    if(N1530) begin
      { mem[7695:7680] } <= { w_data_i[15:0] };
    end 
    if(N1529) begin
      { mem[7679:7664] } <= { w_data_i[15:0] };
    end 
    if(N1528) begin
      { mem[7663:7648] } <= { w_data_i[15:0] };
    end 
    if(N1527) begin
      { mem[7647:7632] } <= { w_data_i[15:0] };
    end 
    if(N1526) begin
      { mem[7631:7616] } <= { w_data_i[15:0] };
    end 
    if(N1525) begin
      { mem[7615:7600] } <= { w_data_i[15:0] };
    end 
    if(N1524) begin
      { mem[7599:7584] } <= { w_data_i[15:0] };
    end 
    if(N1523) begin
      { mem[7583:7568] } <= { w_data_i[15:0] };
    end 
    if(N1522) begin
      { mem[7567:7552] } <= { w_data_i[15:0] };
    end 
    if(N1521) begin
      { mem[7551:7536] } <= { w_data_i[15:0] };
    end 
    if(N1520) begin
      { mem[7535:7520] } <= { w_data_i[15:0] };
    end 
    if(N1519) begin
      { mem[7519:7504] } <= { w_data_i[15:0] };
    end 
    if(N1518) begin
      { mem[7503:7488] } <= { w_data_i[15:0] };
    end 
    if(N1517) begin
      { mem[7487:7472] } <= { w_data_i[15:0] };
    end 
    if(N1516) begin
      { mem[7471:7456] } <= { w_data_i[15:0] };
    end 
    if(N1515) begin
      { mem[7455:7440] } <= { w_data_i[15:0] };
    end 
    if(N1514) begin
      { mem[7439:7424] } <= { w_data_i[15:0] };
    end 
    if(N1513) begin
      { mem[7423:7408] } <= { w_data_i[15:0] };
    end 
    if(N1512) begin
      { mem[7407:7392] } <= { w_data_i[15:0] };
    end 
    if(N1511) begin
      { mem[7391:7376] } <= { w_data_i[15:0] };
    end 
    if(N1510) begin
      { mem[7375:7360] } <= { w_data_i[15:0] };
    end 
    if(N1509) begin
      { mem[7359:7344] } <= { w_data_i[15:0] };
    end 
    if(N1508) begin
      { mem[7343:7328] } <= { w_data_i[15:0] };
    end 
    if(N1507) begin
      { mem[7327:7312] } <= { w_data_i[15:0] };
    end 
    if(N1506) begin
      { mem[7311:7296] } <= { w_data_i[15:0] };
    end 
    if(N1505) begin
      { mem[7295:7280] } <= { w_data_i[15:0] };
    end 
    if(N1504) begin
      { mem[7279:7264] } <= { w_data_i[15:0] };
    end 
    if(N1503) begin
      { mem[7263:7248] } <= { w_data_i[15:0] };
    end 
    if(N1502) begin
      { mem[7247:7232] } <= { w_data_i[15:0] };
    end 
    if(N1501) begin
      { mem[7231:7216] } <= { w_data_i[15:0] };
    end 
    if(N1500) begin
      { mem[7215:7200] } <= { w_data_i[15:0] };
    end 
    if(N1499) begin
      { mem[7199:7184] } <= { w_data_i[15:0] };
    end 
    if(N1498) begin
      { mem[7183:7168] } <= { w_data_i[15:0] };
    end 
    if(N1497) begin
      { mem[7167:7152] } <= { w_data_i[15:0] };
    end 
    if(N1496) begin
      { mem[7151:7136] } <= { w_data_i[15:0] };
    end 
    if(N1495) begin
      { mem[7135:7120] } <= { w_data_i[15:0] };
    end 
    if(N1494) begin
      { mem[7119:7104] } <= { w_data_i[15:0] };
    end 
    if(N1493) begin
      { mem[7103:7088] } <= { w_data_i[15:0] };
    end 
    if(N1492) begin
      { mem[7087:7072] } <= { w_data_i[15:0] };
    end 
    if(N1491) begin
      { mem[7071:7056] } <= { w_data_i[15:0] };
    end 
    if(N1490) begin
      { mem[7055:7040] } <= { w_data_i[15:0] };
    end 
    if(N1489) begin
      { mem[7039:7024] } <= { w_data_i[15:0] };
    end 
    if(N1488) begin
      { mem[7023:7008] } <= { w_data_i[15:0] };
    end 
    if(N1487) begin
      { mem[7007:6992] } <= { w_data_i[15:0] };
    end 
    if(N1486) begin
      { mem[6991:6976] } <= { w_data_i[15:0] };
    end 
    if(N1485) begin
      { mem[6975:6960] } <= { w_data_i[15:0] };
    end 
    if(N1484) begin
      { mem[6959:6944] } <= { w_data_i[15:0] };
    end 
    if(N1483) begin
      { mem[6943:6928] } <= { w_data_i[15:0] };
    end 
    if(N1482) begin
      { mem[6927:6912] } <= { w_data_i[15:0] };
    end 
    if(N1481) begin
      { mem[6911:6896] } <= { w_data_i[15:0] };
    end 
    if(N1480) begin
      { mem[6895:6880] } <= { w_data_i[15:0] };
    end 
    if(N1479) begin
      { mem[6879:6864] } <= { w_data_i[15:0] };
    end 
    if(N1478) begin
      { mem[6863:6848] } <= { w_data_i[15:0] };
    end 
    if(N1477) begin
      { mem[6847:6832] } <= { w_data_i[15:0] };
    end 
    if(N1476) begin
      { mem[6831:6816] } <= { w_data_i[15:0] };
    end 
    if(N1475) begin
      { mem[6815:6800] } <= { w_data_i[15:0] };
    end 
    if(N1474) begin
      { mem[6799:6784] } <= { w_data_i[15:0] };
    end 
    if(N1473) begin
      { mem[6783:6768] } <= { w_data_i[15:0] };
    end 
    if(N1472) begin
      { mem[6767:6752] } <= { w_data_i[15:0] };
    end 
    if(N1471) begin
      { mem[6751:6736] } <= { w_data_i[15:0] };
    end 
    if(N1470) begin
      { mem[6735:6720] } <= { w_data_i[15:0] };
    end 
    if(N1469) begin
      { mem[6719:6704] } <= { w_data_i[15:0] };
    end 
    if(N1468) begin
      { mem[6703:6688] } <= { w_data_i[15:0] };
    end 
    if(N1467) begin
      { mem[6687:6672] } <= { w_data_i[15:0] };
    end 
    if(N1466) begin
      { mem[6671:6656] } <= { w_data_i[15:0] };
    end 
    if(N1465) begin
      { mem[6655:6640] } <= { w_data_i[15:0] };
    end 
    if(N1464) begin
      { mem[6639:6624] } <= { w_data_i[15:0] };
    end 
    if(N1463) begin
      { mem[6623:6608] } <= { w_data_i[15:0] };
    end 
    if(N1462) begin
      { mem[6607:6592] } <= { w_data_i[15:0] };
    end 
    if(N1461) begin
      { mem[6591:6576] } <= { w_data_i[15:0] };
    end 
    if(N1460) begin
      { mem[6575:6560] } <= { w_data_i[15:0] };
    end 
    if(N1459) begin
      { mem[6559:6544] } <= { w_data_i[15:0] };
    end 
    if(N1458) begin
      { mem[6543:6528] } <= { w_data_i[15:0] };
    end 
    if(N1457) begin
      { mem[6527:6512] } <= { w_data_i[15:0] };
    end 
    if(N1456) begin
      { mem[6511:6496] } <= { w_data_i[15:0] };
    end 
    if(N1455) begin
      { mem[6495:6480] } <= { w_data_i[15:0] };
    end 
    if(N1454) begin
      { mem[6479:6464] } <= { w_data_i[15:0] };
    end 
    if(N1453) begin
      { mem[6463:6448] } <= { w_data_i[15:0] };
    end 
    if(N1452) begin
      { mem[6447:6432] } <= { w_data_i[15:0] };
    end 
    if(N1451) begin
      { mem[6431:6416] } <= { w_data_i[15:0] };
    end 
    if(N1450) begin
      { mem[6415:6400] } <= { w_data_i[15:0] };
    end 
    if(N1449) begin
      { mem[6399:6384] } <= { w_data_i[15:0] };
    end 
    if(N1448) begin
      { mem[6383:6368] } <= { w_data_i[15:0] };
    end 
    if(N1447) begin
      { mem[6367:6352] } <= { w_data_i[15:0] };
    end 
    if(N1446) begin
      { mem[6351:6336] } <= { w_data_i[15:0] };
    end 
    if(N1445) begin
      { mem[6335:6320] } <= { w_data_i[15:0] };
    end 
    if(N1444) begin
      { mem[6319:6304] } <= { w_data_i[15:0] };
    end 
    if(N1443) begin
      { mem[6303:6288] } <= { w_data_i[15:0] };
    end 
    if(N1442) begin
      { mem[6287:6272] } <= { w_data_i[15:0] };
    end 
    if(N1441) begin
      { mem[6271:6256] } <= { w_data_i[15:0] };
    end 
    if(N1440) begin
      { mem[6255:6240] } <= { w_data_i[15:0] };
    end 
    if(N1439) begin
      { mem[6239:6224] } <= { w_data_i[15:0] };
    end 
    if(N1438) begin
      { mem[6223:6208] } <= { w_data_i[15:0] };
    end 
    if(N1437) begin
      { mem[6207:6192] } <= { w_data_i[15:0] };
    end 
    if(N1436) begin
      { mem[6191:6176] } <= { w_data_i[15:0] };
    end 
    if(N1435) begin
      { mem[6175:6160] } <= { w_data_i[15:0] };
    end 
    if(N1434) begin
      { mem[6159:6144] } <= { w_data_i[15:0] };
    end 
    if(N1433) begin
      { mem[6143:6128] } <= { w_data_i[15:0] };
    end 
    if(N1432) begin
      { mem[6127:6112] } <= { w_data_i[15:0] };
    end 
    if(N1431) begin
      { mem[6111:6096] } <= { w_data_i[15:0] };
    end 
    if(N1430) begin
      { mem[6095:6080] } <= { w_data_i[15:0] };
    end 
    if(N1429) begin
      { mem[6079:6064] } <= { w_data_i[15:0] };
    end 
    if(N1428) begin
      { mem[6063:6048] } <= { w_data_i[15:0] };
    end 
    if(N1427) begin
      { mem[6047:6032] } <= { w_data_i[15:0] };
    end 
    if(N1426) begin
      { mem[6031:6016] } <= { w_data_i[15:0] };
    end 
    if(N1425) begin
      { mem[6015:6000] } <= { w_data_i[15:0] };
    end 
    if(N1424) begin
      { mem[5999:5984] } <= { w_data_i[15:0] };
    end 
    if(N1423) begin
      { mem[5983:5968] } <= { w_data_i[15:0] };
    end 
    if(N1422) begin
      { mem[5967:5952] } <= { w_data_i[15:0] };
    end 
    if(N1421) begin
      { mem[5951:5936] } <= { w_data_i[15:0] };
    end 
    if(N1420) begin
      { mem[5935:5920] } <= { w_data_i[15:0] };
    end 
    if(N1419) begin
      { mem[5919:5904] } <= { w_data_i[15:0] };
    end 
    if(N1418) begin
      { mem[5903:5888] } <= { w_data_i[15:0] };
    end 
    if(N1417) begin
      { mem[5887:5872] } <= { w_data_i[15:0] };
    end 
    if(N1416) begin
      { mem[5871:5856] } <= { w_data_i[15:0] };
    end 
    if(N1415) begin
      { mem[5855:5840] } <= { w_data_i[15:0] };
    end 
    if(N1414) begin
      { mem[5839:5824] } <= { w_data_i[15:0] };
    end 
    if(N1413) begin
      { mem[5823:5808] } <= { w_data_i[15:0] };
    end 
    if(N1412) begin
      { mem[5807:5792] } <= { w_data_i[15:0] };
    end 
    if(N1411) begin
      { mem[5791:5776] } <= { w_data_i[15:0] };
    end 
    if(N1410) begin
      { mem[5775:5760] } <= { w_data_i[15:0] };
    end 
    if(N1409) begin
      { mem[5759:5744] } <= { w_data_i[15:0] };
    end 
    if(N1408) begin
      { mem[5743:5728] } <= { w_data_i[15:0] };
    end 
    if(N1407) begin
      { mem[5727:5712] } <= { w_data_i[15:0] };
    end 
    if(N1406) begin
      { mem[5711:5696] } <= { w_data_i[15:0] };
    end 
    if(N1405) begin
      { mem[5695:5680] } <= { w_data_i[15:0] };
    end 
    if(N1404) begin
      { mem[5679:5664] } <= { w_data_i[15:0] };
    end 
    if(N1403) begin
      { mem[5663:5648] } <= { w_data_i[15:0] };
    end 
    if(N1402) begin
      { mem[5647:5632] } <= { w_data_i[15:0] };
    end 
    if(N1401) begin
      { mem[5631:5616] } <= { w_data_i[15:0] };
    end 
    if(N1400) begin
      { mem[5615:5600] } <= { w_data_i[15:0] };
    end 
    if(N1399) begin
      { mem[5599:5584] } <= { w_data_i[15:0] };
    end 
    if(N1398) begin
      { mem[5583:5568] } <= { w_data_i[15:0] };
    end 
    if(N1397) begin
      { mem[5567:5552] } <= { w_data_i[15:0] };
    end 
    if(N1396) begin
      { mem[5551:5536] } <= { w_data_i[15:0] };
    end 
    if(N1395) begin
      { mem[5535:5520] } <= { w_data_i[15:0] };
    end 
    if(N1394) begin
      { mem[5519:5504] } <= { w_data_i[15:0] };
    end 
    if(N1393) begin
      { mem[5503:5488] } <= { w_data_i[15:0] };
    end 
    if(N1392) begin
      { mem[5487:5472] } <= { w_data_i[15:0] };
    end 
    if(N1391) begin
      { mem[5471:5456] } <= { w_data_i[15:0] };
    end 
    if(N1390) begin
      { mem[5455:5440] } <= { w_data_i[15:0] };
    end 
    if(N1389) begin
      { mem[5439:5424] } <= { w_data_i[15:0] };
    end 
    if(N1388) begin
      { mem[5423:5408] } <= { w_data_i[15:0] };
    end 
    if(N1387) begin
      { mem[5407:5392] } <= { w_data_i[15:0] };
    end 
    if(N1386) begin
      { mem[5391:5376] } <= { w_data_i[15:0] };
    end 
    if(N1385) begin
      { mem[5375:5360] } <= { w_data_i[15:0] };
    end 
    if(N1384) begin
      { mem[5359:5344] } <= { w_data_i[15:0] };
    end 
    if(N1383) begin
      { mem[5343:5328] } <= { w_data_i[15:0] };
    end 
    if(N1382) begin
      { mem[5327:5312] } <= { w_data_i[15:0] };
    end 
    if(N1381) begin
      { mem[5311:5296] } <= { w_data_i[15:0] };
    end 
    if(N1380) begin
      { mem[5295:5280] } <= { w_data_i[15:0] };
    end 
    if(N1379) begin
      { mem[5279:5264] } <= { w_data_i[15:0] };
    end 
    if(N1378) begin
      { mem[5263:5248] } <= { w_data_i[15:0] };
    end 
    if(N1377) begin
      { mem[5247:5232] } <= { w_data_i[15:0] };
    end 
    if(N1376) begin
      { mem[5231:5216] } <= { w_data_i[15:0] };
    end 
    if(N1375) begin
      { mem[5215:5200] } <= { w_data_i[15:0] };
    end 
    if(N1374) begin
      { mem[5199:5184] } <= { w_data_i[15:0] };
    end 
    if(N1373) begin
      { mem[5183:5168] } <= { w_data_i[15:0] };
    end 
    if(N1372) begin
      { mem[5167:5152] } <= { w_data_i[15:0] };
    end 
    if(N1371) begin
      { mem[5151:5136] } <= { w_data_i[15:0] };
    end 
    if(N1370) begin
      { mem[5135:5120] } <= { w_data_i[15:0] };
    end 
    if(N1369) begin
      { mem[5119:5104] } <= { w_data_i[15:0] };
    end 
    if(N1368) begin
      { mem[5103:5088] } <= { w_data_i[15:0] };
    end 
    if(N1367) begin
      { mem[5087:5072] } <= { w_data_i[15:0] };
    end 
    if(N1366) begin
      { mem[5071:5056] } <= { w_data_i[15:0] };
    end 
    if(N1365) begin
      { mem[5055:5040] } <= { w_data_i[15:0] };
    end 
    if(N1364) begin
      { mem[5039:5024] } <= { w_data_i[15:0] };
    end 
    if(N1363) begin
      { mem[5023:5008] } <= { w_data_i[15:0] };
    end 
    if(N1362) begin
      { mem[5007:4992] } <= { w_data_i[15:0] };
    end 
    if(N1361) begin
      { mem[4991:4976] } <= { w_data_i[15:0] };
    end 
    if(N1360) begin
      { mem[4975:4960] } <= { w_data_i[15:0] };
    end 
    if(N1359) begin
      { mem[4959:4944] } <= { w_data_i[15:0] };
    end 
    if(N1358) begin
      { mem[4943:4928] } <= { w_data_i[15:0] };
    end 
    if(N1357) begin
      { mem[4927:4912] } <= { w_data_i[15:0] };
    end 
    if(N1356) begin
      { mem[4911:4896] } <= { w_data_i[15:0] };
    end 
    if(N1355) begin
      { mem[4895:4880] } <= { w_data_i[15:0] };
    end 
    if(N1354) begin
      { mem[4879:4864] } <= { w_data_i[15:0] };
    end 
    if(N1353) begin
      { mem[4863:4848] } <= { w_data_i[15:0] };
    end 
    if(N1352) begin
      { mem[4847:4832] } <= { w_data_i[15:0] };
    end 
    if(N1351) begin
      { mem[4831:4816] } <= { w_data_i[15:0] };
    end 
    if(N1350) begin
      { mem[4815:4800] } <= { w_data_i[15:0] };
    end 
    if(N1349) begin
      { mem[4799:4784] } <= { w_data_i[15:0] };
    end 
    if(N1348) begin
      { mem[4783:4768] } <= { w_data_i[15:0] };
    end 
    if(N1347) begin
      { mem[4767:4752] } <= { w_data_i[15:0] };
    end 
    if(N1346) begin
      { mem[4751:4736] } <= { w_data_i[15:0] };
    end 
    if(N1345) begin
      { mem[4735:4720] } <= { w_data_i[15:0] };
    end 
    if(N1344) begin
      { mem[4719:4704] } <= { w_data_i[15:0] };
    end 
    if(N1343) begin
      { mem[4703:4688] } <= { w_data_i[15:0] };
    end 
    if(N1342) begin
      { mem[4687:4672] } <= { w_data_i[15:0] };
    end 
    if(N1341) begin
      { mem[4671:4656] } <= { w_data_i[15:0] };
    end 
    if(N1340) begin
      { mem[4655:4640] } <= { w_data_i[15:0] };
    end 
    if(N1339) begin
      { mem[4639:4624] } <= { w_data_i[15:0] };
    end 
    if(N1338) begin
      { mem[4623:4608] } <= { w_data_i[15:0] };
    end 
    if(N1337) begin
      { mem[4607:4592] } <= { w_data_i[15:0] };
    end 
    if(N1336) begin
      { mem[4591:4576] } <= { w_data_i[15:0] };
    end 
    if(N1335) begin
      { mem[4575:4560] } <= { w_data_i[15:0] };
    end 
    if(N1334) begin
      { mem[4559:4544] } <= { w_data_i[15:0] };
    end 
    if(N1333) begin
      { mem[4543:4528] } <= { w_data_i[15:0] };
    end 
    if(N1332) begin
      { mem[4527:4512] } <= { w_data_i[15:0] };
    end 
    if(N1331) begin
      { mem[4511:4496] } <= { w_data_i[15:0] };
    end 
    if(N1330) begin
      { mem[4495:4480] } <= { w_data_i[15:0] };
    end 
    if(N1329) begin
      { mem[4479:4464] } <= { w_data_i[15:0] };
    end 
    if(N1328) begin
      { mem[4463:4448] } <= { w_data_i[15:0] };
    end 
    if(N1327) begin
      { mem[4447:4432] } <= { w_data_i[15:0] };
    end 
    if(N1326) begin
      { mem[4431:4416] } <= { w_data_i[15:0] };
    end 
    if(N1325) begin
      { mem[4415:4400] } <= { w_data_i[15:0] };
    end 
    if(N1324) begin
      { mem[4399:4384] } <= { w_data_i[15:0] };
    end 
    if(N1323) begin
      { mem[4383:4368] } <= { w_data_i[15:0] };
    end 
    if(N1322) begin
      { mem[4367:4352] } <= { w_data_i[15:0] };
    end 
    if(N1321) begin
      { mem[4351:4336] } <= { w_data_i[15:0] };
    end 
    if(N1320) begin
      { mem[4335:4320] } <= { w_data_i[15:0] };
    end 
    if(N1319) begin
      { mem[4319:4304] } <= { w_data_i[15:0] };
    end 
    if(N1318) begin
      { mem[4303:4288] } <= { w_data_i[15:0] };
    end 
    if(N1317) begin
      { mem[4287:4272] } <= { w_data_i[15:0] };
    end 
    if(N1316) begin
      { mem[4271:4256] } <= { w_data_i[15:0] };
    end 
    if(N1315) begin
      { mem[4255:4240] } <= { w_data_i[15:0] };
    end 
    if(N1314) begin
      { mem[4239:4224] } <= { w_data_i[15:0] };
    end 
    if(N1313) begin
      { mem[4223:4208] } <= { w_data_i[15:0] };
    end 
    if(N1312) begin
      { mem[4207:4192] } <= { w_data_i[15:0] };
    end 
    if(N1311) begin
      { mem[4191:4176] } <= { w_data_i[15:0] };
    end 
    if(N1310) begin
      { mem[4175:4160] } <= { w_data_i[15:0] };
    end 
    if(N1309) begin
      { mem[4159:4144] } <= { w_data_i[15:0] };
    end 
    if(N1308) begin
      { mem[4143:4128] } <= { w_data_i[15:0] };
    end 
    if(N1307) begin
      { mem[4127:4112] } <= { w_data_i[15:0] };
    end 
    if(N1306) begin
      { mem[4111:4096] } <= { w_data_i[15:0] };
    end 
    if(N1305) begin
      { mem[4095:4080] } <= { w_data_i[15:0] };
    end 
    if(N1304) begin
      { mem[4079:4064] } <= { w_data_i[15:0] };
    end 
    if(N1303) begin
      { mem[4063:4048] } <= { w_data_i[15:0] };
    end 
    if(N1302) begin
      { mem[4047:4032] } <= { w_data_i[15:0] };
    end 
    if(N1301) begin
      { mem[4031:4016] } <= { w_data_i[15:0] };
    end 
    if(N1300) begin
      { mem[4015:4000] } <= { w_data_i[15:0] };
    end 
    if(N1299) begin
      { mem[3999:3984] } <= { w_data_i[15:0] };
    end 
    if(N1298) begin
      { mem[3983:3968] } <= { w_data_i[15:0] };
    end 
    if(N1297) begin
      { mem[3967:3952] } <= { w_data_i[15:0] };
    end 
    if(N1296) begin
      { mem[3951:3936] } <= { w_data_i[15:0] };
    end 
    if(N1295) begin
      { mem[3935:3920] } <= { w_data_i[15:0] };
    end 
    if(N1294) begin
      { mem[3919:3904] } <= { w_data_i[15:0] };
    end 
    if(N1293) begin
      { mem[3903:3888] } <= { w_data_i[15:0] };
    end 
    if(N1292) begin
      { mem[3887:3872] } <= { w_data_i[15:0] };
    end 
    if(N1291) begin
      { mem[3871:3856] } <= { w_data_i[15:0] };
    end 
    if(N1290) begin
      { mem[3855:3840] } <= { w_data_i[15:0] };
    end 
    if(N1289) begin
      { mem[3839:3824] } <= { w_data_i[15:0] };
    end 
    if(N1288) begin
      { mem[3823:3808] } <= { w_data_i[15:0] };
    end 
    if(N1287) begin
      { mem[3807:3792] } <= { w_data_i[15:0] };
    end 
    if(N1286) begin
      { mem[3791:3776] } <= { w_data_i[15:0] };
    end 
    if(N1285) begin
      { mem[3775:3760] } <= { w_data_i[15:0] };
    end 
    if(N1284) begin
      { mem[3759:3744] } <= { w_data_i[15:0] };
    end 
    if(N1283) begin
      { mem[3743:3728] } <= { w_data_i[15:0] };
    end 
    if(N1282) begin
      { mem[3727:3712] } <= { w_data_i[15:0] };
    end 
    if(N1281) begin
      { mem[3711:3696] } <= { w_data_i[15:0] };
    end 
    if(N1280) begin
      { mem[3695:3680] } <= { w_data_i[15:0] };
    end 
    if(N1279) begin
      { mem[3679:3664] } <= { w_data_i[15:0] };
    end 
    if(N1278) begin
      { mem[3663:3648] } <= { w_data_i[15:0] };
    end 
    if(N1277) begin
      { mem[3647:3632] } <= { w_data_i[15:0] };
    end 
    if(N1276) begin
      { mem[3631:3616] } <= { w_data_i[15:0] };
    end 
    if(N1275) begin
      { mem[3615:3600] } <= { w_data_i[15:0] };
    end 
    if(N1274) begin
      { mem[3599:3584] } <= { w_data_i[15:0] };
    end 
    if(N1273) begin
      { mem[3583:3568] } <= { w_data_i[15:0] };
    end 
    if(N1272) begin
      { mem[3567:3552] } <= { w_data_i[15:0] };
    end 
    if(N1271) begin
      { mem[3551:3536] } <= { w_data_i[15:0] };
    end 
    if(N1270) begin
      { mem[3535:3520] } <= { w_data_i[15:0] };
    end 
    if(N1269) begin
      { mem[3519:3504] } <= { w_data_i[15:0] };
    end 
    if(N1268) begin
      { mem[3503:3488] } <= { w_data_i[15:0] };
    end 
    if(N1267) begin
      { mem[3487:3472] } <= { w_data_i[15:0] };
    end 
    if(N1266) begin
      { mem[3471:3456] } <= { w_data_i[15:0] };
    end 
    if(N1265) begin
      { mem[3455:3440] } <= { w_data_i[15:0] };
    end 
    if(N1264) begin
      { mem[3439:3424] } <= { w_data_i[15:0] };
    end 
    if(N1263) begin
      { mem[3423:3408] } <= { w_data_i[15:0] };
    end 
    if(N1262) begin
      { mem[3407:3392] } <= { w_data_i[15:0] };
    end 
    if(N1261) begin
      { mem[3391:3376] } <= { w_data_i[15:0] };
    end 
    if(N1260) begin
      { mem[3375:3360] } <= { w_data_i[15:0] };
    end 
    if(N1259) begin
      { mem[3359:3344] } <= { w_data_i[15:0] };
    end 
    if(N1258) begin
      { mem[3343:3328] } <= { w_data_i[15:0] };
    end 
    if(N1257) begin
      { mem[3327:3312] } <= { w_data_i[15:0] };
    end 
    if(N1256) begin
      { mem[3311:3296] } <= { w_data_i[15:0] };
    end 
    if(N1255) begin
      { mem[3295:3280] } <= { w_data_i[15:0] };
    end 
    if(N1254) begin
      { mem[3279:3264] } <= { w_data_i[15:0] };
    end 
    if(N1253) begin
      { mem[3263:3248] } <= { w_data_i[15:0] };
    end 
    if(N1252) begin
      { mem[3247:3232] } <= { w_data_i[15:0] };
    end 
    if(N1251) begin
      { mem[3231:3216] } <= { w_data_i[15:0] };
    end 
    if(N1250) begin
      { mem[3215:3200] } <= { w_data_i[15:0] };
    end 
    if(N1249) begin
      { mem[3199:3184] } <= { w_data_i[15:0] };
    end 
    if(N1248) begin
      { mem[3183:3168] } <= { w_data_i[15:0] };
    end 
    if(N1247) begin
      { mem[3167:3152] } <= { w_data_i[15:0] };
    end 
    if(N1246) begin
      { mem[3151:3136] } <= { w_data_i[15:0] };
    end 
    if(N1245) begin
      { mem[3135:3120] } <= { w_data_i[15:0] };
    end 
    if(N1244) begin
      { mem[3119:3104] } <= { w_data_i[15:0] };
    end 
    if(N1243) begin
      { mem[3103:3088] } <= { w_data_i[15:0] };
    end 
    if(N1242) begin
      { mem[3087:3072] } <= { w_data_i[15:0] };
    end 
    if(N1241) begin
      { mem[3071:3056] } <= { w_data_i[15:0] };
    end 
    if(N1240) begin
      { mem[3055:3040] } <= { w_data_i[15:0] };
    end 
    if(N1239) begin
      { mem[3039:3024] } <= { w_data_i[15:0] };
    end 
    if(N1238) begin
      { mem[3023:3008] } <= { w_data_i[15:0] };
    end 
    if(N1237) begin
      { mem[3007:2992] } <= { w_data_i[15:0] };
    end 
    if(N1236) begin
      { mem[2991:2976] } <= { w_data_i[15:0] };
    end 
    if(N1235) begin
      { mem[2975:2960] } <= { w_data_i[15:0] };
    end 
    if(N1234) begin
      { mem[2959:2944] } <= { w_data_i[15:0] };
    end 
    if(N1233) begin
      { mem[2943:2928] } <= { w_data_i[15:0] };
    end 
    if(N1232) begin
      { mem[2927:2912] } <= { w_data_i[15:0] };
    end 
    if(N1231) begin
      { mem[2911:2896] } <= { w_data_i[15:0] };
    end 
    if(N1230) begin
      { mem[2895:2880] } <= { w_data_i[15:0] };
    end 
    if(N1229) begin
      { mem[2879:2864] } <= { w_data_i[15:0] };
    end 
    if(N1228) begin
      { mem[2863:2848] } <= { w_data_i[15:0] };
    end 
    if(N1227) begin
      { mem[2847:2832] } <= { w_data_i[15:0] };
    end 
    if(N1226) begin
      { mem[2831:2816] } <= { w_data_i[15:0] };
    end 
    if(N1225) begin
      { mem[2815:2800] } <= { w_data_i[15:0] };
    end 
    if(N1224) begin
      { mem[2799:2784] } <= { w_data_i[15:0] };
    end 
    if(N1223) begin
      { mem[2783:2768] } <= { w_data_i[15:0] };
    end 
    if(N1222) begin
      { mem[2767:2752] } <= { w_data_i[15:0] };
    end 
    if(N1221) begin
      { mem[2751:2736] } <= { w_data_i[15:0] };
    end 
    if(N1220) begin
      { mem[2735:2720] } <= { w_data_i[15:0] };
    end 
    if(N1219) begin
      { mem[2719:2704] } <= { w_data_i[15:0] };
    end 
    if(N1218) begin
      { mem[2703:2688] } <= { w_data_i[15:0] };
    end 
    if(N1217) begin
      { mem[2687:2672] } <= { w_data_i[15:0] };
    end 
    if(N1216) begin
      { mem[2671:2656] } <= { w_data_i[15:0] };
    end 
    if(N1215) begin
      { mem[2655:2640] } <= { w_data_i[15:0] };
    end 
    if(N1214) begin
      { mem[2639:2624] } <= { w_data_i[15:0] };
    end 
    if(N1213) begin
      { mem[2623:2608] } <= { w_data_i[15:0] };
    end 
    if(N1212) begin
      { mem[2607:2592] } <= { w_data_i[15:0] };
    end 
    if(N1211) begin
      { mem[2591:2576] } <= { w_data_i[15:0] };
    end 
    if(N1210) begin
      { mem[2575:2560] } <= { w_data_i[15:0] };
    end 
    if(N1209) begin
      { mem[2559:2544] } <= { w_data_i[15:0] };
    end 
    if(N1208) begin
      { mem[2543:2528] } <= { w_data_i[15:0] };
    end 
    if(N1207) begin
      { mem[2527:2512] } <= { w_data_i[15:0] };
    end 
    if(N1206) begin
      { mem[2511:2496] } <= { w_data_i[15:0] };
    end 
    if(N1205) begin
      { mem[2495:2480] } <= { w_data_i[15:0] };
    end 
    if(N1204) begin
      { mem[2479:2464] } <= { w_data_i[15:0] };
    end 
    if(N1203) begin
      { mem[2463:2448] } <= { w_data_i[15:0] };
    end 
    if(N1202) begin
      { mem[2447:2432] } <= { w_data_i[15:0] };
    end 
    if(N1201) begin
      { mem[2431:2416] } <= { w_data_i[15:0] };
    end 
    if(N1200) begin
      { mem[2415:2400] } <= { w_data_i[15:0] };
    end 
    if(N1199) begin
      { mem[2399:2384] } <= { w_data_i[15:0] };
    end 
    if(N1198) begin
      { mem[2383:2368] } <= { w_data_i[15:0] };
    end 
    if(N1197) begin
      { mem[2367:2352] } <= { w_data_i[15:0] };
    end 
    if(N1196) begin
      { mem[2351:2336] } <= { w_data_i[15:0] };
    end 
    if(N1195) begin
      { mem[2335:2320] } <= { w_data_i[15:0] };
    end 
    if(N1194) begin
      { mem[2319:2304] } <= { w_data_i[15:0] };
    end 
    if(N1193) begin
      { mem[2303:2288] } <= { w_data_i[15:0] };
    end 
    if(N1192) begin
      { mem[2287:2272] } <= { w_data_i[15:0] };
    end 
    if(N1191) begin
      { mem[2271:2256] } <= { w_data_i[15:0] };
    end 
    if(N1190) begin
      { mem[2255:2240] } <= { w_data_i[15:0] };
    end 
    if(N1189) begin
      { mem[2239:2224] } <= { w_data_i[15:0] };
    end 
    if(N1188) begin
      { mem[2223:2208] } <= { w_data_i[15:0] };
    end 
    if(N1187) begin
      { mem[2207:2192] } <= { w_data_i[15:0] };
    end 
    if(N1186) begin
      { mem[2191:2176] } <= { w_data_i[15:0] };
    end 
    if(N1185) begin
      { mem[2175:2160] } <= { w_data_i[15:0] };
    end 
    if(N1184) begin
      { mem[2159:2144] } <= { w_data_i[15:0] };
    end 
    if(N1183) begin
      { mem[2143:2128] } <= { w_data_i[15:0] };
    end 
    if(N1182) begin
      { mem[2127:2112] } <= { w_data_i[15:0] };
    end 
    if(N1181) begin
      { mem[2111:2096] } <= { w_data_i[15:0] };
    end 
    if(N1180) begin
      { mem[2095:2080] } <= { w_data_i[15:0] };
    end 
    if(N1179) begin
      { mem[2079:2064] } <= { w_data_i[15:0] };
    end 
    if(N1178) begin
      { mem[2063:2048] } <= { w_data_i[15:0] };
    end 
    if(N1177) begin
      { mem[2047:2032] } <= { w_data_i[15:0] };
    end 
    if(N1176) begin
      { mem[2031:2016] } <= { w_data_i[15:0] };
    end 
    if(N1175) begin
      { mem[2015:2000] } <= { w_data_i[15:0] };
    end 
    if(N1174) begin
      { mem[1999:1984] } <= { w_data_i[15:0] };
    end 
    if(N1173) begin
      { mem[1983:1968] } <= { w_data_i[15:0] };
    end 
    if(N1172) begin
      { mem[1967:1952] } <= { w_data_i[15:0] };
    end 
    if(N1171) begin
      { mem[1951:1936] } <= { w_data_i[15:0] };
    end 
    if(N1170) begin
      { mem[1935:1920] } <= { w_data_i[15:0] };
    end 
    if(N1169) begin
      { mem[1919:1904] } <= { w_data_i[15:0] };
    end 
    if(N1168) begin
      { mem[1903:1888] } <= { w_data_i[15:0] };
    end 
    if(N1167) begin
      { mem[1887:1872] } <= { w_data_i[15:0] };
    end 
    if(N1166) begin
      { mem[1871:1856] } <= { w_data_i[15:0] };
    end 
    if(N1165) begin
      { mem[1855:1840] } <= { w_data_i[15:0] };
    end 
    if(N1164) begin
      { mem[1839:1824] } <= { w_data_i[15:0] };
    end 
    if(N1163) begin
      { mem[1823:1808] } <= { w_data_i[15:0] };
    end 
    if(N1162) begin
      { mem[1807:1792] } <= { w_data_i[15:0] };
    end 
    if(N1161) begin
      { mem[1791:1776] } <= { w_data_i[15:0] };
    end 
    if(N1160) begin
      { mem[1775:1760] } <= { w_data_i[15:0] };
    end 
    if(N1159) begin
      { mem[1759:1744] } <= { w_data_i[15:0] };
    end 
    if(N1158) begin
      { mem[1743:1728] } <= { w_data_i[15:0] };
    end 
    if(N1157) begin
      { mem[1727:1712] } <= { w_data_i[15:0] };
    end 
    if(N1156) begin
      { mem[1711:1696] } <= { w_data_i[15:0] };
    end 
    if(N1155) begin
      { mem[1695:1680] } <= { w_data_i[15:0] };
    end 
    if(N1154) begin
      { mem[1679:1664] } <= { w_data_i[15:0] };
    end 
    if(N1153) begin
      { mem[1663:1648] } <= { w_data_i[15:0] };
    end 
    if(N1152) begin
      { mem[1647:1632] } <= { w_data_i[15:0] };
    end 
    if(N1151) begin
      { mem[1631:1616] } <= { w_data_i[15:0] };
    end 
    if(N1150) begin
      { mem[1615:1600] } <= { w_data_i[15:0] };
    end 
    if(N1149) begin
      { mem[1599:1584] } <= { w_data_i[15:0] };
    end 
    if(N1148) begin
      { mem[1583:1568] } <= { w_data_i[15:0] };
    end 
    if(N1147) begin
      { mem[1567:1552] } <= { w_data_i[15:0] };
    end 
    if(N1146) begin
      { mem[1551:1536] } <= { w_data_i[15:0] };
    end 
    if(N1145) begin
      { mem[1535:1520] } <= { w_data_i[15:0] };
    end 
    if(N1144) begin
      { mem[1519:1504] } <= { w_data_i[15:0] };
    end 
    if(N1143) begin
      { mem[1503:1488] } <= { w_data_i[15:0] };
    end 
    if(N1142) begin
      { mem[1487:1472] } <= { w_data_i[15:0] };
    end 
    if(N1141) begin
      { mem[1471:1456] } <= { w_data_i[15:0] };
    end 
    if(N1140) begin
      { mem[1455:1440] } <= { w_data_i[15:0] };
    end 
    if(N1139) begin
      { mem[1439:1424] } <= { w_data_i[15:0] };
    end 
    if(N1138) begin
      { mem[1423:1408] } <= { w_data_i[15:0] };
    end 
    if(N1137) begin
      { mem[1407:1392] } <= { w_data_i[15:0] };
    end 
    if(N1136) begin
      { mem[1391:1376] } <= { w_data_i[15:0] };
    end 
    if(N1135) begin
      { mem[1375:1360] } <= { w_data_i[15:0] };
    end 
    if(N1134) begin
      { mem[1359:1344] } <= { w_data_i[15:0] };
    end 
    if(N1133) begin
      { mem[1343:1328] } <= { w_data_i[15:0] };
    end 
    if(N1132) begin
      { mem[1327:1312] } <= { w_data_i[15:0] };
    end 
    if(N1131) begin
      { mem[1311:1296] } <= { w_data_i[15:0] };
    end 
    if(N1130) begin
      { mem[1295:1280] } <= { w_data_i[15:0] };
    end 
    if(N1129) begin
      { mem[1279:1264] } <= { w_data_i[15:0] };
    end 
    if(N1128) begin
      { mem[1263:1248] } <= { w_data_i[15:0] };
    end 
    if(N1127) begin
      { mem[1247:1232] } <= { w_data_i[15:0] };
    end 
    if(N1126) begin
      { mem[1231:1216] } <= { w_data_i[15:0] };
    end 
    if(N1125) begin
      { mem[1215:1200] } <= { w_data_i[15:0] };
    end 
    if(N1124) begin
      { mem[1199:1184] } <= { w_data_i[15:0] };
    end 
    if(N1123) begin
      { mem[1183:1168] } <= { w_data_i[15:0] };
    end 
    if(N1122) begin
      { mem[1167:1152] } <= { w_data_i[15:0] };
    end 
    if(N1121) begin
      { mem[1151:1136] } <= { w_data_i[15:0] };
    end 
    if(N1120) begin
      { mem[1135:1120] } <= { w_data_i[15:0] };
    end 
    if(N1119) begin
      { mem[1119:1104] } <= { w_data_i[15:0] };
    end 
    if(N1118) begin
      { mem[1103:1088] } <= { w_data_i[15:0] };
    end 
    if(N1117) begin
      { mem[1087:1072] } <= { w_data_i[15:0] };
    end 
    if(N1116) begin
      { mem[1071:1056] } <= { w_data_i[15:0] };
    end 
    if(N1115) begin
      { mem[1055:1040] } <= { w_data_i[15:0] };
    end 
    if(N1114) begin
      { mem[1039:1024] } <= { w_data_i[15:0] };
    end 
    if(N1113) begin
      { mem[1023:1008] } <= { w_data_i[15:0] };
    end 
    if(N1112) begin
      { mem[1007:992] } <= { w_data_i[15:0] };
    end 
    if(N1111) begin
      { mem[991:976] } <= { w_data_i[15:0] };
    end 
    if(N1110) begin
      { mem[975:960] } <= { w_data_i[15:0] };
    end 
    if(N1109) begin
      { mem[959:944] } <= { w_data_i[15:0] };
    end 
    if(N1108) begin
      { mem[943:928] } <= { w_data_i[15:0] };
    end 
    if(N1107) begin
      { mem[927:912] } <= { w_data_i[15:0] };
    end 
    if(N1106) begin
      { mem[911:896] } <= { w_data_i[15:0] };
    end 
    if(N1105) begin
      { mem[895:880] } <= { w_data_i[15:0] };
    end 
    if(N1104) begin
      { mem[879:864] } <= { w_data_i[15:0] };
    end 
    if(N1103) begin
      { mem[863:848] } <= { w_data_i[15:0] };
    end 
    if(N1102) begin
      { mem[847:832] } <= { w_data_i[15:0] };
    end 
    if(N1101) begin
      { mem[831:816] } <= { w_data_i[15:0] };
    end 
    if(N1100) begin
      { mem[815:800] } <= { w_data_i[15:0] };
    end 
    if(N1099) begin
      { mem[799:784] } <= { w_data_i[15:0] };
    end 
    if(N1098) begin
      { mem[783:768] } <= { w_data_i[15:0] };
    end 
    if(N1097) begin
      { mem[767:752] } <= { w_data_i[15:0] };
    end 
    if(N1096) begin
      { mem[751:736] } <= { w_data_i[15:0] };
    end 
    if(N1095) begin
      { mem[735:720] } <= { w_data_i[15:0] };
    end 
    if(N1094) begin
      { mem[719:704] } <= { w_data_i[15:0] };
    end 
    if(N1093) begin
      { mem[703:688] } <= { w_data_i[15:0] };
    end 
    if(N1092) begin
      { mem[687:672] } <= { w_data_i[15:0] };
    end 
    if(N1091) begin
      { mem[671:656] } <= { w_data_i[15:0] };
    end 
    if(N1090) begin
      { mem[655:640] } <= { w_data_i[15:0] };
    end 
    if(N1089) begin
      { mem[639:624] } <= { w_data_i[15:0] };
    end 
    if(N1088) begin
      { mem[623:608] } <= { w_data_i[15:0] };
    end 
    if(N1087) begin
      { mem[607:592] } <= { w_data_i[15:0] };
    end 
    if(N1086) begin
      { mem[591:576] } <= { w_data_i[15:0] };
    end 
    if(N1085) begin
      { mem[575:560] } <= { w_data_i[15:0] };
    end 
    if(N1084) begin
      { mem[559:544] } <= { w_data_i[15:0] };
    end 
    if(N1083) begin
      { mem[543:528] } <= { w_data_i[15:0] };
    end 
    if(N1082) begin
      { mem[527:512] } <= { w_data_i[15:0] };
    end 
    if(N1081) begin
      { mem[511:496] } <= { w_data_i[15:0] };
    end 
    if(N1080) begin
      { mem[495:480] } <= { w_data_i[15:0] };
    end 
    if(N1079) begin
      { mem[479:464] } <= { w_data_i[15:0] };
    end 
    if(N1078) begin
      { mem[463:448] } <= { w_data_i[15:0] };
    end 
    if(N1077) begin
      { mem[447:432] } <= { w_data_i[15:0] };
    end 
    if(N1076) begin
      { mem[431:416] } <= { w_data_i[15:0] };
    end 
    if(N1075) begin
      { mem[415:400] } <= { w_data_i[15:0] };
    end 
    if(N1074) begin
      { mem[399:384] } <= { w_data_i[15:0] };
    end 
    if(N1073) begin
      { mem[383:368] } <= { w_data_i[15:0] };
    end 
    if(N1072) begin
      { mem[367:352] } <= { w_data_i[15:0] };
    end 
    if(N1071) begin
      { mem[351:336] } <= { w_data_i[15:0] };
    end 
    if(N1070) begin
      { mem[335:320] } <= { w_data_i[15:0] };
    end 
    if(N1069) begin
      { mem[319:304] } <= { w_data_i[15:0] };
    end 
    if(N1068) begin
      { mem[303:288] } <= { w_data_i[15:0] };
    end 
    if(N1067) begin
      { mem[287:272] } <= { w_data_i[15:0] };
    end 
    if(N1066) begin
      { mem[271:256] } <= { w_data_i[15:0] };
    end 
    if(N1065) begin
      { mem[255:240] } <= { w_data_i[15:0] };
    end 
    if(N1064) begin
      { mem[239:224] } <= { w_data_i[15:0] };
    end 
    if(N1063) begin
      { mem[223:208] } <= { w_data_i[15:0] };
    end 
    if(N1062) begin
      { mem[207:192] } <= { w_data_i[15:0] };
    end 
    if(N1061) begin
      { mem[191:176] } <= { w_data_i[15:0] };
    end 
    if(N1060) begin
      { mem[175:160] } <= { w_data_i[15:0] };
    end 
    if(N1059) begin
      { mem[159:144] } <= { w_data_i[15:0] };
    end 
    if(N1058) begin
      { mem[143:128] } <= { w_data_i[15:0] };
    end 
    if(N1057) begin
      { mem[127:112] } <= { w_data_i[15:0] };
    end 
    if(N1056) begin
      { mem[111:96] } <= { w_data_i[15:0] };
    end 
    if(N1055) begin
      { mem[95:80] } <= { w_data_i[15:0] };
    end 
    if(N1054) begin
      { mem[79:64] } <= { w_data_i[15:0] };
    end 
    if(N1053) begin
      { mem[63:48] } <= { w_data_i[15:0] };
    end 
    if(N1052) begin
      { mem[47:32] } <= { w_data_i[15:0] };
    end 
    if(N1051) begin
      { mem[31:16] } <= { w_data_i[15:0] };
    end 
    if(N1050) begin
      { mem[15:0] } <= { w_data_i[15:0] };
    end 
    if(N1049) begin
      { valid[511:511] } <= { N533 };
    end 
    if(N1048) begin
      { valid[510:510] } <= { N533 };
    end 
    if(N1047) begin
      { valid[509:509] } <= { N533 };
    end 
    if(N1046) begin
      { valid[508:508] } <= { N533 };
    end 
    if(N1045) begin
      { valid[507:507] } <= { N533 };
    end 
    if(N1044) begin
      { valid[506:506] } <= { N533 };
    end 
    if(N1043) begin
      { valid[505:505] } <= { N533 };
    end 
    if(N1042) begin
      { valid[504:504] } <= { N533 };
    end 
    if(N1041) begin
      { valid[503:503] } <= { N533 };
    end 
    if(N1040) begin
      { valid[502:502] } <= { N533 };
    end 
    if(N1039) begin
      { valid[501:501] } <= { N533 };
    end 
    if(N1038) begin
      { valid[500:500] } <= { N533 };
    end 
    if(N1037) begin
      { valid[499:499] } <= { N533 };
    end 
    if(N1036) begin
      { valid[498:498] } <= { N533 };
    end 
    if(N1035) begin
      { valid[497:497] } <= { N533 };
    end 
    if(N1034) begin
      { valid[496:496] } <= { N533 };
    end 
    if(N1033) begin
      { valid[495:495] } <= { N533 };
    end 
    if(N1032) begin
      { valid[494:494] } <= { N533 };
    end 
    if(N1031) begin
      { valid[493:493] } <= { N533 };
    end 
    if(N1030) begin
      { valid[492:492] } <= { N533 };
    end 
    if(N1029) begin
      { valid[491:491] } <= { N533 };
    end 
    if(N1028) begin
      { valid[490:490] } <= { N533 };
    end 
    if(N1027) begin
      { valid[489:489] } <= { N533 };
    end 
    if(N1026) begin
      { valid[488:488] } <= { N533 };
    end 
    if(N1025) begin
      { valid[487:487] } <= { N533 };
    end 
    if(N1024) begin
      { valid[486:486] } <= { N533 };
    end 
    if(N1023) begin
      { valid[485:485] } <= { N533 };
    end 
    if(N1022) begin
      { valid[484:484] } <= { N533 };
    end 
    if(N1021) begin
      { valid[483:483] } <= { N533 };
    end 
    if(N1020) begin
      { valid[482:482] } <= { N533 };
    end 
    if(N1019) begin
      { valid[481:481] } <= { N533 };
    end 
    if(N1018) begin
      { valid[480:480] } <= { N533 };
    end 
    if(N1017) begin
      { valid[479:479] } <= { N533 };
    end 
    if(N1016) begin
      { valid[478:478] } <= { N533 };
    end 
    if(N1015) begin
      { valid[477:477] } <= { N533 };
    end 
    if(N1014) begin
      { valid[476:476] } <= { N533 };
    end 
    if(N1013) begin
      { valid[475:475] } <= { N533 };
    end 
    if(N1012) begin
      { valid[474:474] } <= { N533 };
    end 
    if(N1011) begin
      { valid[473:473] } <= { N533 };
    end 
    if(N1010) begin
      { valid[472:472] } <= { N533 };
    end 
    if(N1009) begin
      { valid[471:471] } <= { N533 };
    end 
    if(N1008) begin
      { valid[470:470] } <= { N533 };
    end 
    if(N1007) begin
      { valid[469:469] } <= { N533 };
    end 
    if(N1006) begin
      { valid[468:468] } <= { N533 };
    end 
    if(N1005) begin
      { valid[467:467] } <= { N533 };
    end 
    if(N1004) begin
      { valid[466:466] } <= { N533 };
    end 
    if(N1003) begin
      { valid[465:465] } <= { N533 };
    end 
    if(N1002) begin
      { valid[464:464] } <= { N533 };
    end 
    if(N1001) begin
      { valid[463:463] } <= { N533 };
    end 
    if(N1000) begin
      { valid[462:462] } <= { N533 };
    end 
    if(N999) begin
      { valid[461:461] } <= { N533 };
    end 
    if(N998) begin
      { valid[460:460] } <= { N533 };
    end 
    if(N997) begin
      { valid[459:459] } <= { N533 };
    end 
    if(N996) begin
      { valid[458:458] } <= { N533 };
    end 
    if(N995) begin
      { valid[457:457] } <= { N533 };
    end 
    if(N994) begin
      { valid[456:456] } <= { N533 };
    end 
    if(N993) begin
      { valid[455:455] } <= { N533 };
    end 
    if(N992) begin
      { valid[454:454] } <= { N533 };
    end 
    if(N991) begin
      { valid[453:453] } <= { N533 };
    end 
    if(N990) begin
      { valid[452:452] } <= { N533 };
    end 
    if(N989) begin
      { valid[451:451] } <= { N533 };
    end 
    if(N988) begin
      { valid[450:450] } <= { N533 };
    end 
    if(N987) begin
      { valid[449:449] } <= { N533 };
    end 
    if(N986) begin
      { valid[448:448] } <= { N533 };
    end 
    if(N985) begin
      { valid[447:447] } <= { N533 };
    end 
    if(N984) begin
      { valid[446:446] } <= { N533 };
    end 
    if(N983) begin
      { valid[445:445] } <= { N533 };
    end 
    if(N982) begin
      { valid[444:444] } <= { N533 };
    end 
    if(N981) begin
      { valid[443:443] } <= { N533 };
    end 
    if(N980) begin
      { valid[442:442] } <= { N533 };
    end 
    if(N979) begin
      { valid[441:441] } <= { N533 };
    end 
    if(N978) begin
      { valid[440:440] } <= { N533 };
    end 
    if(N977) begin
      { valid[439:439] } <= { N533 };
    end 
    if(N976) begin
      { valid[438:438] } <= { N533 };
    end 
    if(N975) begin
      { valid[437:437] } <= { N533 };
    end 
    if(N974) begin
      { valid[436:436] } <= { N533 };
    end 
    if(N973) begin
      { valid[435:435] } <= { N533 };
    end 
    if(N972) begin
      { valid[434:434] } <= { N533 };
    end 
    if(N971) begin
      { valid[433:433] } <= { N533 };
    end 
    if(N970) begin
      { valid[432:432] } <= { N533 };
    end 
    if(N969) begin
      { valid[431:431] } <= { N533 };
    end 
    if(N968) begin
      { valid[430:430] } <= { N533 };
    end 
    if(N967) begin
      { valid[429:429] } <= { N533 };
    end 
    if(N966) begin
      { valid[428:428] } <= { N533 };
    end 
    if(N965) begin
      { valid[427:427] } <= { N533 };
    end 
    if(N964) begin
      { valid[426:426] } <= { N533 };
    end 
    if(N963) begin
      { valid[425:425] } <= { N533 };
    end 
    if(N962) begin
      { valid[424:424] } <= { N533 };
    end 
    if(N961) begin
      { valid[423:423] } <= { N533 };
    end 
    if(N960) begin
      { valid[422:422] } <= { N533 };
    end 
    if(N959) begin
      { valid[421:421] } <= { N533 };
    end 
    if(N958) begin
      { valid[420:420] } <= { N533 };
    end 
    if(N957) begin
      { valid[419:419] } <= { N533 };
    end 
    if(N956) begin
      { valid[418:418] } <= { N533 };
    end 
    if(N955) begin
      { valid[417:417] } <= { N533 };
    end 
    if(N954) begin
      { valid[416:416] } <= { N533 };
    end 
    if(N953) begin
      { valid[415:415] } <= { N533 };
    end 
    if(N952) begin
      { valid[414:414] } <= { N533 };
    end 
    if(N951) begin
      { valid[413:413] } <= { N533 };
    end 
    if(N950) begin
      { valid[412:412] } <= { N535 };
    end 
    if(N949) begin
      { valid[411:411] } <= { N535 };
    end 
    if(N948) begin
      { valid[410:410] } <= { N535 };
    end 
    if(N947) begin
      { valid[409:409] } <= { N535 };
    end 
    if(N946) begin
      { valid[408:408] } <= { N535 };
    end 
    if(N945) begin
      { valid[407:407] } <= { N535 };
    end 
    if(N944) begin
      { valid[406:406] } <= { N535 };
    end 
    if(N943) begin
      { valid[405:405] } <= { N535 };
    end 
    if(N942) begin
      { valid[404:404] } <= { N535 };
    end 
    if(N941) begin
      { valid[403:403] } <= { N535 };
    end 
    if(N940) begin
      { valid[402:402] } <= { N535 };
    end 
    if(N939) begin
      { valid[401:401] } <= { N535 };
    end 
    if(N938) begin
      { valid[400:400] } <= { N535 };
    end 
    if(N937) begin
      { valid[399:399] } <= { N535 };
    end 
    if(N936) begin
      { valid[398:398] } <= { N535 };
    end 
    if(N935) begin
      { valid[397:397] } <= { N535 };
    end 
    if(N934) begin
      { valid[396:396] } <= { N535 };
    end 
    if(N933) begin
      { valid[395:395] } <= { N535 };
    end 
    if(N932) begin
      { valid[394:394] } <= { N535 };
    end 
    if(N931) begin
      { valid[393:393] } <= { N535 };
    end 
    if(N930) begin
      { valid[392:392] } <= { N535 };
    end 
    if(N929) begin
      { valid[391:391] } <= { N535 };
    end 
    if(N928) begin
      { valid[390:390] } <= { N535 };
    end 
    if(N927) begin
      { valid[389:389] } <= { N535 };
    end 
    if(N926) begin
      { valid[388:388] } <= { N535 };
    end 
    if(N925) begin
      { valid[387:387] } <= { N535 };
    end 
    if(N924) begin
      { valid[386:386] } <= { N535 };
    end 
    if(N923) begin
      { valid[385:385] } <= { N535 };
    end 
    if(N922) begin
      { valid[384:384] } <= { N535 };
    end 
    if(N921) begin
      { valid[383:383] } <= { N535 };
    end 
    if(N920) begin
      { valid[382:382] } <= { N535 };
    end 
    if(N919) begin
      { valid[381:381] } <= { N535 };
    end 
    if(N918) begin
      { valid[380:380] } <= { N535 };
    end 
    if(N917) begin
      { valid[379:379] } <= { N535 };
    end 
    if(N916) begin
      { valid[378:378] } <= { N535 };
    end 
    if(N915) begin
      { valid[377:377] } <= { N535 };
    end 
    if(N914) begin
      { valid[376:376] } <= { N535 };
    end 
    if(N913) begin
      { valid[375:375] } <= { N535 };
    end 
    if(N912) begin
      { valid[374:374] } <= { N535 };
    end 
    if(N911) begin
      { valid[373:373] } <= { N535 };
    end 
    if(N910) begin
      { valid[372:372] } <= { N535 };
    end 
    if(N909) begin
      { valid[371:371] } <= { N535 };
    end 
    if(N908) begin
      { valid[370:370] } <= { N535 };
    end 
    if(N907) begin
      { valid[369:369] } <= { N535 };
    end 
    if(N906) begin
      { valid[368:368] } <= { N535 };
    end 
    if(N905) begin
      { valid[367:367] } <= { N535 };
    end 
    if(N904) begin
      { valid[366:366] } <= { N535 };
    end 
    if(N903) begin
      { valid[365:365] } <= { N535 };
    end 
    if(N902) begin
      { valid[364:364] } <= { N535 };
    end 
    if(N901) begin
      { valid[363:363] } <= { N535 };
    end 
    if(N900) begin
      { valid[362:362] } <= { N535 };
    end 
    if(N899) begin
      { valid[361:361] } <= { N535 };
    end 
    if(N898) begin
      { valid[360:360] } <= { N535 };
    end 
    if(N897) begin
      { valid[359:359] } <= { N535 };
    end 
    if(N896) begin
      { valid[358:358] } <= { N535 };
    end 
    if(N895) begin
      { valid[357:357] } <= { N535 };
    end 
    if(N894) begin
      { valid[356:356] } <= { N535 };
    end 
    if(N893) begin
      { valid[355:355] } <= { N535 };
    end 
    if(N892) begin
      { valid[354:354] } <= { N535 };
    end 
    if(N891) begin
      { valid[353:353] } <= { N535 };
    end 
    if(N890) begin
      { valid[352:352] } <= { N535 };
    end 
    if(N889) begin
      { valid[351:351] } <= { N535 };
    end 
    if(N888) begin
      { valid[350:350] } <= { N535 };
    end 
    if(N887) begin
      { valid[349:349] } <= { N535 };
    end 
    if(N886) begin
      { valid[348:348] } <= { N535 };
    end 
    if(N885) begin
      { valid[347:347] } <= { N535 };
    end 
    if(N884) begin
      { valid[346:346] } <= { N535 };
    end 
    if(N883) begin
      { valid[345:345] } <= { N535 };
    end 
    if(N882) begin
      { valid[344:344] } <= { N535 };
    end 
    if(N881) begin
      { valid[343:343] } <= { N535 };
    end 
    if(N880) begin
      { valid[342:342] } <= { N535 };
    end 
    if(N879) begin
      { valid[341:341] } <= { N535 };
    end 
    if(N878) begin
      { valid[340:340] } <= { N535 };
    end 
    if(N877) begin
      { valid[339:339] } <= { N535 };
    end 
    if(N876) begin
      { valid[338:338] } <= { N535 };
    end 
    if(N875) begin
      { valid[337:337] } <= { N535 };
    end 
    if(N874) begin
      { valid[336:336] } <= { N535 };
    end 
    if(N873) begin
      { valid[335:335] } <= { N535 };
    end 
    if(N872) begin
      { valid[334:334] } <= { N535 };
    end 
    if(N871) begin
      { valid[333:333] } <= { N535 };
    end 
    if(N870) begin
      { valid[332:332] } <= { N535 };
    end 
    if(N869) begin
      { valid[331:331] } <= { N535 };
    end 
    if(N868) begin
      { valid[330:330] } <= { N535 };
    end 
    if(N867) begin
      { valid[329:329] } <= { N535 };
    end 
    if(N866) begin
      { valid[328:328] } <= { N535 };
    end 
    if(N865) begin
      { valid[327:327] } <= { N535 };
    end 
    if(N864) begin
      { valid[326:326] } <= { N535 };
    end 
    if(N863) begin
      { valid[325:325] } <= { N535 };
    end 
    if(N862) begin
      { valid[324:324] } <= { N535 };
    end 
    if(N861) begin
      { valid[323:323] } <= { N535 };
    end 
    if(N860) begin
      { valid[322:322] } <= { N535 };
    end 
    if(N859) begin
      { valid[321:321] } <= { N535 };
    end 
    if(N858) begin
      { valid[320:320] } <= { N535 };
    end 
    if(N857) begin
      { valid[319:319] } <= { N535 };
    end 
    if(N856) begin
      { valid[318:318] } <= { N535 };
    end 
    if(N855) begin
      { valid[317:317] } <= { N535 };
    end 
    if(N854) begin
      { valid[316:316] } <= { N535 };
    end 
    if(N853) begin
      { valid[315:315] } <= { N535 };
    end 
    if(N852) begin
      { valid[314:314] } <= { N535 };
    end 
    if(N851) begin
      { valid[313:313] } <= { N537 };
    end 
    if(N850) begin
      { valid[312:312] } <= { N537 };
    end 
    if(N849) begin
      { valid[311:311] } <= { N537 };
    end 
    if(N848) begin
      { valid[310:310] } <= { N537 };
    end 
    if(N847) begin
      { valid[309:309] } <= { N537 };
    end 
    if(N846) begin
      { valid[308:308] } <= { N537 };
    end 
    if(N845) begin
      { valid[307:307] } <= { N537 };
    end 
    if(N844) begin
      { valid[306:306] } <= { N537 };
    end 
    if(N843) begin
      { valid[305:305] } <= { N537 };
    end 
    if(N842) begin
      { valid[304:304] } <= { N537 };
    end 
    if(N841) begin
      { valid[303:303] } <= { N537 };
    end 
    if(N840) begin
      { valid[302:302] } <= { N537 };
    end 
    if(N839) begin
      { valid[301:301] } <= { N537 };
    end 
    if(N838) begin
      { valid[300:300] } <= { N537 };
    end 
    if(N837) begin
      { valid[299:299] } <= { N537 };
    end 
    if(N836) begin
      { valid[298:298] } <= { N537 };
    end 
    if(N835) begin
      { valid[297:297] } <= { N537 };
    end 
    if(N834) begin
      { valid[296:296] } <= { N537 };
    end 
    if(N833) begin
      { valid[295:295] } <= { N537 };
    end 
    if(N832) begin
      { valid[294:294] } <= { N537 };
    end 
    if(N831) begin
      { valid[293:293] } <= { N537 };
    end 
    if(N830) begin
      { valid[292:292] } <= { N537 };
    end 
    if(N829) begin
      { valid[291:291] } <= { N537 };
    end 
    if(N828) begin
      { valid[290:290] } <= { N537 };
    end 
    if(N827) begin
      { valid[289:289] } <= { N537 };
    end 
    if(N826) begin
      { valid[288:288] } <= { N537 };
    end 
    if(N825) begin
      { valid[287:287] } <= { N537 };
    end 
    if(N824) begin
      { valid[286:286] } <= { N537 };
    end 
    if(N823) begin
      { valid[285:285] } <= { N537 };
    end 
    if(N822) begin
      { valid[284:284] } <= { N537 };
    end 
    if(N821) begin
      { valid[283:283] } <= { N537 };
    end 
    if(N820) begin
      { valid[282:282] } <= { N537 };
    end 
    if(N819) begin
      { valid[281:281] } <= { N537 };
    end 
    if(N818) begin
      { valid[280:280] } <= { N537 };
    end 
    if(N817) begin
      { valid[279:279] } <= { N537 };
    end 
    if(N816) begin
      { valid[278:278] } <= { N537 };
    end 
    if(N815) begin
      { valid[277:277] } <= { N537 };
    end 
    if(N814) begin
      { valid[276:276] } <= { N537 };
    end 
    if(N813) begin
      { valid[275:275] } <= { N537 };
    end 
    if(N812) begin
      { valid[274:274] } <= { N537 };
    end 
    if(N811) begin
      { valid[273:273] } <= { N537 };
    end 
    if(N810) begin
      { valid[272:272] } <= { N537 };
    end 
    if(N809) begin
      { valid[271:271] } <= { N537 };
    end 
    if(N808) begin
      { valid[270:270] } <= { N537 };
    end 
    if(N807) begin
      { valid[269:269] } <= { N537 };
    end 
    if(N806) begin
      { valid[268:268] } <= { N537 };
    end 
    if(N805) begin
      { valid[267:267] } <= { N537 };
    end 
    if(N804) begin
      { valid[266:266] } <= { N537 };
    end 
    if(N803) begin
      { valid[265:265] } <= { N537 };
    end 
    if(N802) begin
      { valid[264:264] } <= { N537 };
    end 
    if(N801) begin
      { valid[263:263] } <= { N537 };
    end 
    if(N800) begin
      { valid[262:262] } <= { N537 };
    end 
    if(N799) begin
      { valid[261:261] } <= { N537 };
    end 
    if(N798) begin
      { valid[260:260] } <= { N537 };
    end 
    if(N797) begin
      { valid[259:259] } <= { N537 };
    end 
    if(N796) begin
      { valid[258:258] } <= { N537 };
    end 
    if(N795) begin
      { valid[257:257] } <= { N537 };
    end 
    if(N794) begin
      { valid[256:256] } <= { N537 };
    end 
    if(N793) begin
      { valid[255:255] } <= { N537 };
    end 
    if(N792) begin
      { valid[254:254] } <= { N537 };
    end 
    if(N791) begin
      { valid[253:253] } <= { N537 };
    end 
    if(N790) begin
      { valid[252:252] } <= { N537 };
    end 
    if(N789) begin
      { valid[251:251] } <= { N537 };
    end 
    if(N788) begin
      { valid[250:250] } <= { N537 };
    end 
    if(N787) begin
      { valid[249:249] } <= { N537 };
    end 
    if(N786) begin
      { valid[248:248] } <= { N537 };
    end 
    if(N785) begin
      { valid[247:247] } <= { N537 };
    end 
    if(N784) begin
      { valid[246:246] } <= { N537 };
    end 
    if(N783) begin
      { valid[245:245] } <= { N537 };
    end 
    if(N782) begin
      { valid[244:244] } <= { N537 };
    end 
    if(N781) begin
      { valid[243:243] } <= { N537 };
    end 
    if(N780) begin
      { valid[242:242] } <= { N537 };
    end 
    if(N779) begin
      { valid[241:241] } <= { N537 };
    end 
    if(N778) begin
      { valid[240:240] } <= { N537 };
    end 
    if(N777) begin
      { valid[239:239] } <= { N537 };
    end 
    if(N776) begin
      { valid[238:238] } <= { N537 };
    end 
    if(N775) begin
      { valid[237:237] } <= { N537 };
    end 
    if(N774) begin
      { valid[236:236] } <= { N537 };
    end 
    if(N773) begin
      { valid[235:235] } <= { N537 };
    end 
    if(N772) begin
      { valid[234:234] } <= { N537 };
    end 
    if(N771) begin
      { valid[233:233] } <= { N537 };
    end 
    if(N770) begin
      { valid[232:232] } <= { N537 };
    end 
    if(N769) begin
      { valid[231:231] } <= { N537 };
    end 
    if(N768) begin
      { valid[230:230] } <= { N537 };
    end 
    if(N767) begin
      { valid[229:229] } <= { N537 };
    end 
    if(N766) begin
      { valid[228:228] } <= { N537 };
    end 
    if(N765) begin
      { valid[227:227] } <= { N537 };
    end 
    if(N764) begin
      { valid[226:226] } <= { N537 };
    end 
    if(N763) begin
      { valid[225:225] } <= { N537 };
    end 
    if(N762) begin
      { valid[224:224] } <= { N537 };
    end 
    if(N761) begin
      { valid[223:223] } <= { N537 };
    end 
    if(N760) begin
      { valid[222:222] } <= { N537 };
    end 
    if(N759) begin
      { valid[221:221] } <= { N537 };
    end 
    if(N758) begin
      { valid[220:220] } <= { N537 };
    end 
    if(N757) begin
      { valid[219:219] } <= { N537 };
    end 
    if(N756) begin
      { valid[218:218] } <= { N537 };
    end 
    if(N755) begin
      { valid[217:217] } <= { N537 };
    end 
    if(N754) begin
      { valid[216:216] } <= { N537 };
    end 
    if(N753) begin
      { valid[215:215] } <= { N537 };
    end 
    if(N752) begin
      { valid[214:214] } <= { N539 };
    end 
    if(N751) begin
      { valid[213:213] } <= { N539 };
    end 
    if(N750) begin
      { valid[212:212] } <= { N539 };
    end 
    if(N749) begin
      { valid[211:211] } <= { N539 };
    end 
    if(N748) begin
      { valid[210:210] } <= { N539 };
    end 
    if(N747) begin
      { valid[209:209] } <= { N539 };
    end 
    if(N746) begin
      { valid[208:208] } <= { N539 };
    end 
    if(N745) begin
      { valid[207:207] } <= { N539 };
    end 
    if(N744) begin
      { valid[206:206] } <= { N539 };
    end 
    if(N743) begin
      { valid[205:205] } <= { N539 };
    end 
    if(N742) begin
      { valid[204:204] } <= { N539 };
    end 
    if(N741) begin
      { valid[203:203] } <= { N539 };
    end 
    if(N740) begin
      { valid[202:202] } <= { N539 };
    end 
    if(N739) begin
      { valid[201:201] } <= { N539 };
    end 
    if(N738) begin
      { valid[200:200] } <= { N539 };
    end 
    if(N737) begin
      { valid[199:199] } <= { N539 };
    end 
    if(N736) begin
      { valid[198:198] } <= { N539 };
    end 
    if(N735) begin
      { valid[197:197] } <= { N539 };
    end 
    if(N734) begin
      { valid[196:196] } <= { N539 };
    end 
    if(N733) begin
      { valid[195:195] } <= { N539 };
    end 
    if(N732) begin
      { valid[194:194] } <= { N539 };
    end 
    if(N731) begin
      { valid[193:193] } <= { N539 };
    end 
    if(N730) begin
      { valid[192:192] } <= { N539 };
    end 
    if(N729) begin
      { valid[191:191] } <= { N539 };
    end 
    if(N728) begin
      { valid[190:190] } <= { N539 };
    end 
    if(N727) begin
      { valid[189:189] } <= { N539 };
    end 
    if(N726) begin
      { valid[188:188] } <= { N539 };
    end 
    if(N725) begin
      { valid[187:187] } <= { N539 };
    end 
    if(N724) begin
      { valid[186:186] } <= { N539 };
    end 
    if(N723) begin
      { valid[185:185] } <= { N539 };
    end 
    if(N722) begin
      { valid[184:184] } <= { N539 };
    end 
    if(N721) begin
      { valid[183:183] } <= { N539 };
    end 
    if(N720) begin
      { valid[182:182] } <= { N539 };
    end 
    if(N719) begin
      { valid[181:181] } <= { N539 };
    end 
    if(N718) begin
      { valid[180:180] } <= { N539 };
    end 
    if(N717) begin
      { valid[179:179] } <= { N539 };
    end 
    if(N716) begin
      { valid[178:178] } <= { N539 };
    end 
    if(N715) begin
      { valid[177:177] } <= { N539 };
    end 
    if(N714) begin
      { valid[176:176] } <= { N539 };
    end 
    if(N713) begin
      { valid[175:175] } <= { N539 };
    end 
    if(N712) begin
      { valid[174:174] } <= { N539 };
    end 
    if(N711) begin
      { valid[173:173] } <= { N539 };
    end 
    if(N710) begin
      { valid[172:172] } <= { N539 };
    end 
    if(N709) begin
      { valid[171:171] } <= { N539 };
    end 
    if(N708) begin
      { valid[170:170] } <= { N539 };
    end 
    if(N707) begin
      { valid[169:169] } <= { N539 };
    end 
    if(N706) begin
      { valid[168:168] } <= { N539 };
    end 
    if(N705) begin
      { valid[167:167] } <= { N539 };
    end 
    if(N704) begin
      { valid[166:166] } <= { N539 };
    end 
    if(N703) begin
      { valid[165:165] } <= { N539 };
    end 
    if(N702) begin
      { valid[164:164] } <= { N539 };
    end 
    if(N701) begin
      { valid[163:163] } <= { N539 };
    end 
    if(N700) begin
      { valid[162:162] } <= { N539 };
    end 
    if(N699) begin
      { valid[161:161] } <= { N539 };
    end 
    if(N698) begin
      { valid[160:160] } <= { N539 };
    end 
    if(N697) begin
      { valid[159:159] } <= { N539 };
    end 
    if(N696) begin
      { valid[158:158] } <= { N539 };
    end 
    if(N695) begin
      { valid[157:157] } <= { N539 };
    end 
    if(N694) begin
      { valid[156:156] } <= { N539 };
    end 
    if(N693) begin
      { valid[155:155] } <= { N539 };
    end 
    if(N692) begin
      { valid[154:154] } <= { N539 };
    end 
    if(N691) begin
      { valid[153:153] } <= { N539 };
    end 
    if(N690) begin
      { valid[152:152] } <= { N539 };
    end 
    if(N689) begin
      { valid[151:151] } <= { N539 };
    end 
    if(N688) begin
      { valid[150:150] } <= { N539 };
    end 
    if(N687) begin
      { valid[149:149] } <= { N539 };
    end 
    if(N686) begin
      { valid[148:148] } <= { N539 };
    end 
    if(N685) begin
      { valid[147:147] } <= { N539 };
    end 
    if(N684) begin
      { valid[146:146] } <= { N539 };
    end 
    if(N683) begin
      { valid[145:145] } <= { N539 };
    end 
    if(N682) begin
      { valid[144:144] } <= { N539 };
    end 
    if(N681) begin
      { valid[143:143] } <= { N539 };
    end 
    if(N680) begin
      { valid[142:142] } <= { N539 };
    end 
    if(N679) begin
      { valid[141:141] } <= { N539 };
    end 
    if(N678) begin
      { valid[140:140] } <= { N539 };
    end 
    if(N677) begin
      { valid[139:139] } <= { N539 };
    end 
    if(N676) begin
      { valid[138:138] } <= { N539 };
    end 
    if(N675) begin
      { valid[137:137] } <= { N539 };
    end 
    if(N674) begin
      { valid[136:136] } <= { N539 };
    end 
    if(N673) begin
      { valid[135:135] } <= { N539 };
    end 
    if(N672) begin
      { valid[134:134] } <= { N539 };
    end 
    if(N671) begin
      { valid[133:133] } <= { N539 };
    end 
    if(N670) begin
      { valid[132:132] } <= { N539 };
    end 
    if(N669) begin
      { valid[131:131] } <= { N539 };
    end 
    if(N668) begin
      { valid[130:130] } <= { N539 };
    end 
    if(N667) begin
      { valid[129:129] } <= { N539 };
    end 
    if(N666) begin
      { valid[128:128] } <= { N539 };
    end 
    if(N665) begin
      { valid[127:127] } <= { N539 };
    end 
    if(N664) begin
      { valid[126:126] } <= { N539 };
    end 
    if(N663) begin
      { valid[125:125] } <= { N539 };
    end 
    if(N662) begin
      { valid[124:124] } <= { N539 };
    end 
    if(N661) begin
      { valid[123:123] } <= { N539 };
    end 
    if(N660) begin
      { valid[122:122] } <= { N539 };
    end 
    if(N659) begin
      { valid[121:121] } <= { N539 };
    end 
    if(N658) begin
      { valid[120:120] } <= { N539 };
    end 
    if(N657) begin
      { valid[119:119] } <= { N539 };
    end 
    if(N656) begin
      { valid[118:118] } <= { N539 };
    end 
    if(N655) begin
      { valid[117:117] } <= { N539 };
    end 
    if(N654) begin
      { valid[116:116] } <= { N539 };
    end 
    if(N653) begin
      { valid[115:115] } <= { N541 };
    end 
    if(N652) begin
      { valid[114:114] } <= { N541 };
    end 
    if(N651) begin
      { valid[113:113] } <= { N541 };
    end 
    if(N650) begin
      { valid[112:112] } <= { N541 };
    end 
    if(N649) begin
      { valid[111:111] } <= { N541 };
    end 
    if(N648) begin
      { valid[110:110] } <= { N541 };
    end 
    if(N647) begin
      { valid[109:109] } <= { N541 };
    end 
    if(N646) begin
      { valid[108:108] } <= { N541 };
    end 
    if(N645) begin
      { valid[107:107] } <= { N541 };
    end 
    if(N644) begin
      { valid[106:106] } <= { N541 };
    end 
    if(N643) begin
      { valid[105:105] } <= { N541 };
    end 
    if(N642) begin
      { valid[104:104] } <= { N541 };
    end 
    if(N641) begin
      { valid[103:103] } <= { N541 };
    end 
    if(N640) begin
      { valid[102:102] } <= { N541 };
    end 
    if(N639) begin
      { valid[101:101] } <= { N541 };
    end 
    if(N638) begin
      { valid[100:100] } <= { N541 };
    end 
    if(N637) begin
      { valid[99:99] } <= { N541 };
    end 
    if(N636) begin
      { valid[98:98] } <= { N541 };
    end 
    if(N635) begin
      { valid[97:97] } <= { N541 };
    end 
    if(N634) begin
      { valid[96:96] } <= { N541 };
    end 
    if(N633) begin
      { valid[95:95] } <= { N541 };
    end 
    if(N632) begin
      { valid[94:94] } <= { N541 };
    end 
    if(N631) begin
      { valid[93:93] } <= { N541 };
    end 
    if(N630) begin
      { valid[92:92] } <= { N541 };
    end 
    if(N629) begin
      { valid[91:91] } <= { N541 };
    end 
    if(N628) begin
      { valid[90:90] } <= { N541 };
    end 
    if(N627) begin
      { valid[89:89] } <= { N541 };
    end 
    if(N626) begin
      { valid[88:88] } <= { N541 };
    end 
    if(N625) begin
      { valid[87:87] } <= { N541 };
    end 
    if(N624) begin
      { valid[86:86] } <= { N541 };
    end 
    if(N623) begin
      { valid[85:85] } <= { N541 };
    end 
    if(N622) begin
      { valid[84:84] } <= { N541 };
    end 
    if(N621) begin
      { valid[83:83] } <= { N541 };
    end 
    if(N620) begin
      { valid[82:82] } <= { N541 };
    end 
    if(N619) begin
      { valid[81:81] } <= { N541 };
    end 
    if(N618) begin
      { valid[80:80] } <= { N541 };
    end 
    if(N617) begin
      { valid[79:79] } <= { N541 };
    end 
    if(N616) begin
      { valid[78:78] } <= { N541 };
    end 
    if(N615) begin
      { valid[77:77] } <= { N541 };
    end 
    if(N614) begin
      { valid[76:76] } <= { N541 };
    end 
    if(N613) begin
      { valid[75:75] } <= { N541 };
    end 
    if(N612) begin
      { valid[74:74] } <= { N541 };
    end 
    if(N611) begin
      { valid[73:73] } <= { N541 };
    end 
    if(N610) begin
      { valid[72:72] } <= { N541 };
    end 
    if(N609) begin
      { valid[71:71] } <= { N541 };
    end 
    if(N608) begin
      { valid[70:70] } <= { N541 };
    end 
    if(N607) begin
      { valid[69:69] } <= { N541 };
    end 
    if(N606) begin
      { valid[68:68] } <= { N541 };
    end 
    if(N605) begin
      { valid[67:67] } <= { N541 };
    end 
    if(N604) begin
      { valid[66:66] } <= { N541 };
    end 
    if(N603) begin
      { valid[65:65] } <= { N541 };
    end 
    if(N602) begin
      { valid[64:64] } <= { N541 };
    end 
    if(N601) begin
      { valid[63:63] } <= { N541 };
    end 
    if(N600) begin
      { valid[62:62] } <= { N541 };
    end 
    if(N599) begin
      { valid[61:61] } <= { N541 };
    end 
    if(N598) begin
      { valid[60:60] } <= { N541 };
    end 
    if(N597) begin
      { valid[59:59] } <= { N541 };
    end 
    if(N596) begin
      { valid[58:58] } <= { N541 };
    end 
    if(N595) begin
      { valid[57:57] } <= { N541 };
    end 
    if(N594) begin
      { valid[56:56] } <= { N541 };
    end 
    if(N593) begin
      { valid[55:55] } <= { N541 };
    end 
    if(N592) begin
      { valid[54:54] } <= { N541 };
    end 
    if(N591) begin
      { valid[53:53] } <= { N541 };
    end 
    if(N590) begin
      { valid[52:52] } <= { N541 };
    end 
    if(N589) begin
      { valid[51:51] } <= { N541 };
    end 
    if(N588) begin
      { valid[50:50] } <= { N541 };
    end 
    if(N587) begin
      { valid[49:49] } <= { N541 };
    end 
    if(N586) begin
      { valid[48:48] } <= { N541 };
    end 
    if(N585) begin
      { valid[47:47] } <= { N541 };
    end 
    if(N584) begin
      { valid[46:46] } <= { N541 };
    end 
    if(N583) begin
      { valid[45:45] } <= { N541 };
    end 
    if(N582) begin
      { valid[44:44] } <= { N541 };
    end 
    if(N581) begin
      { valid[43:43] } <= { N541 };
    end 
    if(N580) begin
      { valid[42:42] } <= { N541 };
    end 
    if(N579) begin
      { valid[41:41] } <= { N541 };
    end 
    if(N578) begin
      { valid[40:40] } <= { N541 };
    end 
    if(N577) begin
      { valid[39:39] } <= { N541 };
    end 
    if(N576) begin
      { valid[38:38] } <= { N541 };
    end 
    if(N575) begin
      { valid[37:37] } <= { N541 };
    end 
    if(N574) begin
      { valid[36:36] } <= { N541 };
    end 
    if(N573) begin
      { valid[35:35] } <= { N541 };
    end 
    if(N572) begin
      { valid[34:34] } <= { N541 };
    end 
    if(N571) begin
      { valid[33:33] } <= { N541 };
    end 
    if(N570) begin
      { valid[32:32] } <= { N541 };
    end 
    if(N569) begin
      { valid[31:31] } <= { N541 };
    end 
    if(N568) begin
      { valid[30:30] } <= { N541 };
    end 
    if(N567) begin
      { valid[29:29] } <= { N541 };
    end 
    if(N566) begin
      { valid[28:28] } <= { N541 };
    end 
    if(N565) begin
      { valid[27:27] } <= { N541 };
    end 
    if(N564) begin
      { valid[26:26] } <= { N541 };
    end 
    if(N563) begin
      { valid[25:25] } <= { N541 };
    end 
    if(N562) begin
      { valid[24:24] } <= { N541 };
    end 
    if(N561) begin
      { valid[23:23] } <= { N541 };
    end 
    if(N560) begin
      { valid[22:22] } <= { N541 };
    end 
    if(N559) begin
      { valid[21:21] } <= { N541 };
    end 
    if(N558) begin
      { valid[20:20] } <= { N541 };
    end 
    if(N557) begin
      { valid[19:19] } <= { N541 };
    end 
    if(N556) begin
      { valid[18:18] } <= { N541 };
    end 
    if(N555) begin
      { valid[17:17] } <= { N541 };
    end 
    if(N554) begin
      { valid[16:16] } <= { N543 };
    end 
    if(N553) begin
      { valid[15:15] } <= { N543 };
    end 
    if(N552) begin
      { valid[14:14] } <= { N543 };
    end 
    if(N551) begin
      { valid[13:13] } <= { N543 };
    end 
    if(N550) begin
      { valid[12:12] } <= { N543 };
    end 
    if(N549) begin
      { valid[11:11] } <= { N543 };
    end 
    if(N548) begin
      { valid[10:10] } <= { N543 };
    end 
    if(N547) begin
      { valid[9:9] } <= { N543 };
    end 
    if(N546) begin
      { valid[8:8] } <= { N543 };
    end 
    if(N545) begin
      { valid[7:7] } <= { N543 };
    end 
    if(N544) begin
      { valid[6:6] } <= { N543 };
    end 
    if(N542) begin
      { valid[5:5] } <= { N543 };
    end 
    if(N540) begin
      { valid[4:4] } <= { N541 };
    end 
    if(N538) begin
      { valid[3:3] } <= { N539 };
    end 
    if(N536) begin
      { valid[2:2] } <= { N537 };
    end 
    if(N534) begin
      { valid[1:1] } <= { N535 };
    end 
    if(N532) begin
      { valid[0:0] } <= { N533 };
    end 
  end


endmodule

