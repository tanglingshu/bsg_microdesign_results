

module top
(
  clk_i,
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [511:0] sel_i;
  output [31:0] data_o;
  input clk_i;

  bsg_fifo_shift_datapath
  wrapper
  (
    .data_i(data_i),
    .sel_i(sel_i),
    .data_o(data_o),
    .clk_i(clk_i)
  );


endmodule



module bsg_fifo_shift_datapath
(
  clk_i,
  data_i,
  sel_i,
  data_o
);

  input [31:0] data_i;
  input [511:0] sel_i;
  output [31:0] data_o;
  input clk_i;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,
  r_n_0__31_,r_n_0__30_,r_n_0__29_,r_n_0__28_,r_n_0__27_,r_n_0__26_,r_n_0__25_,
  r_n_0__24_,r_n_0__23_,r_n_0__22_,r_n_0__21_,r_n_0__20_,r_n_0__19_,r_n_0__18_,r_n_0__17_,
  r_n_0__16_,r_n_0__15_,r_n_0__14_,r_n_0__13_,r_n_0__12_,r_n_0__11_,r_n_0__10_,
  r_n_0__9_,r_n_0__8_,r_n_0__7_,r_n_0__6_,r_n_0__5_,r_n_0__4_,r_n_0__3_,r_n_0__2_,
  r_n_0__1_,r_n_0__0_,r_n_16__31_,r_n_16__30_,r_n_16__29_,r_n_16__28_,r_n_16__27_,
  r_n_16__26_,r_n_16__25_,r_n_16__24_,r_n_16__23_,r_n_16__22_,r_n_16__21_,
  r_n_16__20_,r_n_16__19_,r_n_16__18_,r_n_16__17_,r_n_16__16_,r_n_16__15_,r_n_16__14_,
  r_n_16__13_,r_n_16__12_,r_n_16__11_,r_n_16__10_,r_n_16__9_,r_n_16__8_,r_n_16__7_,
  r_n_16__6_,r_n_16__5_,r_n_16__4_,r_n_16__3_,r_n_16__2_,r_n_16__1_,r_n_16__0_,
  r_n_15__31_,r_n_15__30_,r_n_15__29_,r_n_15__28_,r_n_15__27_,r_n_15__26_,r_n_15__25_,
  r_n_15__24_,r_n_15__23_,r_n_15__22_,r_n_15__21_,r_n_15__20_,r_n_15__19_,r_n_15__18_,
  r_n_15__17_,r_n_15__16_,r_n_15__15_,r_n_15__14_,r_n_15__13_,r_n_15__12_,
  r_n_15__11_,r_n_15__10_,r_n_15__9_,r_n_15__8_,r_n_15__7_,r_n_15__6_,r_n_15__5_,
  r_n_15__4_,r_n_15__3_,r_n_15__2_,r_n_15__1_,r_n_15__0_,r_n_14__31_,r_n_14__30_,
  r_n_14__29_,r_n_14__28_,r_n_14__27_,r_n_14__26_,r_n_14__25_,r_n_14__24_,r_n_14__23_,
  r_n_14__22_,r_n_14__21_,r_n_14__20_,r_n_14__19_,r_n_14__18_,r_n_14__17_,r_n_14__16_,
  r_n_14__15_,r_n_14__14_,r_n_14__13_,r_n_14__12_,r_n_14__11_,r_n_14__10_,r_n_14__9_,
  r_n_14__8_,r_n_14__7_,r_n_14__6_,r_n_14__5_,r_n_14__4_,r_n_14__3_,r_n_14__2_,
  r_n_14__1_,r_n_14__0_,r_n_13__31_,r_n_13__30_,r_n_13__29_,r_n_13__28_,r_n_13__27_,
  r_n_13__26_,r_n_13__25_,r_n_13__24_,r_n_13__23_,r_n_13__22_,r_n_13__21_,
  r_n_13__20_,r_n_13__19_,r_n_13__18_,r_n_13__17_,r_n_13__16_,r_n_13__15_,r_n_13__14_,
  r_n_13__13_,r_n_13__12_,r_n_13__11_,r_n_13__10_,r_n_13__9_,r_n_13__8_,r_n_13__7_,
  r_n_13__6_,r_n_13__5_,r_n_13__4_,r_n_13__3_,r_n_13__2_,r_n_13__1_,r_n_13__0_,
  r_n_12__31_,r_n_12__30_,r_n_12__29_,r_n_12__28_,r_n_12__27_,r_n_12__26_,r_n_12__25_,
  r_n_12__24_,r_n_12__23_,r_n_12__22_,r_n_12__21_,r_n_12__20_,r_n_12__19_,
  r_n_12__18_,r_n_12__17_,r_n_12__16_,r_n_12__15_,r_n_12__14_,r_n_12__13_,r_n_12__12_,
  r_n_12__11_,r_n_12__10_,r_n_12__9_,r_n_12__8_,r_n_12__7_,r_n_12__6_,r_n_12__5_,
  r_n_12__4_,r_n_12__3_,r_n_12__2_,r_n_12__1_,r_n_12__0_,r_n_11__31_,r_n_11__30_,
  r_n_11__29_,r_n_11__28_,r_n_11__27_,r_n_11__26_,r_n_11__25_,r_n_11__24_,r_n_11__23_,
  r_n_11__22_,r_n_11__21_,r_n_11__20_,r_n_11__19_,r_n_11__18_,r_n_11__17_,r_n_11__16_,
  r_n_11__15_,r_n_11__14_,r_n_11__13_,r_n_11__12_,r_n_11__11_,r_n_11__10_,
  r_n_11__9_,r_n_11__8_,r_n_11__7_,r_n_11__6_,r_n_11__5_,r_n_11__4_,r_n_11__3_,r_n_11__2_,
  r_n_11__1_,r_n_11__0_,r_n_10__31_,r_n_10__30_,r_n_10__29_,r_n_10__28_,
  r_n_10__27_,r_n_10__26_,r_n_10__25_,r_n_10__24_,r_n_10__23_,r_n_10__22_,r_n_10__21_,
  r_n_10__20_,r_n_10__19_,r_n_10__18_,r_n_10__17_,r_n_10__16_,r_n_10__15_,r_n_10__14_,
  r_n_10__13_,r_n_10__12_,r_n_10__11_,r_n_10__10_,r_n_10__9_,r_n_10__8_,r_n_10__7_,
  r_n_10__6_,r_n_10__5_,r_n_10__4_,r_n_10__3_,r_n_10__2_,r_n_10__1_,r_n_10__0_,
  r_n_9__31_,r_n_9__30_,r_n_9__29_,r_n_9__28_,r_n_9__27_,r_n_9__26_,r_n_9__25_,
  r_n_9__24_,r_n_9__23_,r_n_9__22_,r_n_9__21_,r_n_9__20_,r_n_9__19_,r_n_9__18_,r_n_9__17_,
  r_n_9__16_,r_n_9__15_,r_n_9__14_,r_n_9__13_,r_n_9__12_,r_n_9__11_,r_n_9__10_,
  r_n_9__9_,r_n_9__8_,r_n_9__7_,r_n_9__6_,r_n_9__5_,r_n_9__4_,r_n_9__3_,r_n_9__2_,
  r_n_9__1_,r_n_9__0_,r_n_8__31_,r_n_8__30_,r_n_8__29_,r_n_8__28_,r_n_8__27_,
  r_n_8__26_,r_n_8__25_,r_n_8__24_,r_n_8__23_,r_n_8__22_,r_n_8__21_,r_n_8__20_,r_n_8__19_,
  r_n_8__18_,r_n_8__17_,r_n_8__16_,r_n_8__15_,r_n_8__14_,r_n_8__13_,r_n_8__12_,
  r_n_8__11_,r_n_8__10_,r_n_8__9_,r_n_8__8_,r_n_8__7_,r_n_8__6_,r_n_8__5_,r_n_8__4_,
  r_n_8__3_,r_n_8__2_,r_n_8__1_,r_n_8__0_,r_n_7__31_,r_n_7__30_,r_n_7__29_,
  r_n_7__28_,r_n_7__27_,r_n_7__26_,r_n_7__25_,r_n_7__24_,r_n_7__23_,r_n_7__22_,r_n_7__21_,
  r_n_7__20_,r_n_7__19_,r_n_7__18_,r_n_7__17_,r_n_7__16_,r_n_7__15_,r_n_7__14_,
  r_n_7__13_,r_n_7__12_,r_n_7__11_,r_n_7__10_,r_n_7__9_,r_n_7__8_,r_n_7__7_,
  r_n_7__6_,r_n_7__5_,r_n_7__4_,r_n_7__3_,r_n_7__2_,r_n_7__1_,r_n_7__0_,r_n_6__31_,
  r_n_6__30_,r_n_6__29_,r_n_6__28_,r_n_6__27_,r_n_6__26_,r_n_6__25_,r_n_6__24_,r_n_6__23_,
  r_n_6__22_,r_n_6__21_,r_n_6__20_,r_n_6__19_,r_n_6__18_,r_n_6__17_,r_n_6__16_,
  r_n_6__15_,r_n_6__14_,r_n_6__13_,r_n_6__12_,r_n_6__11_,r_n_6__10_,r_n_6__9_,
  r_n_6__8_,r_n_6__7_,r_n_6__6_,r_n_6__5_,r_n_6__4_,r_n_6__3_,r_n_6__2_,r_n_6__1_,
  r_n_6__0_,r_n_5__31_,r_n_5__30_,r_n_5__29_,r_n_5__28_,r_n_5__27_,r_n_5__26_,r_n_5__25_,
  r_n_5__24_,r_n_5__23_,r_n_5__22_,r_n_5__21_,r_n_5__20_,r_n_5__19_,r_n_5__18_,
  r_n_5__17_,r_n_5__16_,r_n_5__15_,r_n_5__14_,r_n_5__13_,r_n_5__12_,r_n_5__11_,
  r_n_5__10_,r_n_5__9_,r_n_5__8_,r_n_5__7_,r_n_5__6_,r_n_5__5_,r_n_5__4_,r_n_5__3_,
  r_n_5__2_,r_n_5__1_,r_n_5__0_,r_n_4__31_,r_n_4__30_,r_n_4__29_,r_n_4__28_,r_n_4__27_,
  r_n_4__26_,r_n_4__25_,r_n_4__24_,r_n_4__23_,r_n_4__22_,r_n_4__21_,r_n_4__20_,
  r_n_4__19_,r_n_4__18_,r_n_4__17_,r_n_4__16_,r_n_4__15_,r_n_4__14_,r_n_4__13_,
  r_n_4__12_,r_n_4__11_,r_n_4__10_,r_n_4__9_,r_n_4__8_,r_n_4__7_,r_n_4__6_,r_n_4__5_,
  r_n_4__4_,r_n_4__3_,r_n_4__2_,r_n_4__1_,r_n_4__0_,r_n_3__31_,r_n_3__30_,r_n_3__29_,
  r_n_3__28_,r_n_3__27_,r_n_3__26_,r_n_3__25_,r_n_3__24_,r_n_3__23_,r_n_3__22_,
  r_n_3__21_,r_n_3__20_,r_n_3__19_,r_n_3__18_,r_n_3__17_,r_n_3__16_,r_n_3__15_,
  r_n_3__14_,r_n_3__13_,r_n_3__12_,r_n_3__11_,r_n_3__10_,r_n_3__9_,r_n_3__8_,r_n_3__7_,
  r_n_3__6_,r_n_3__5_,r_n_3__4_,r_n_3__3_,r_n_3__2_,r_n_3__1_,r_n_3__0_,r_n_2__31_,
  r_n_2__30_,r_n_2__29_,r_n_2__28_,r_n_2__27_,r_n_2__26_,r_n_2__25_,r_n_2__24_,
  r_n_2__23_,r_n_2__22_,r_n_2__21_,r_n_2__20_,r_n_2__19_,r_n_2__18_,r_n_2__17_,
  r_n_2__16_,r_n_2__15_,r_n_2__14_,r_n_2__13_,r_n_2__12_,r_n_2__11_,r_n_2__10_,
  r_n_2__9_,r_n_2__8_,r_n_2__7_,r_n_2__6_,r_n_2__5_,r_n_2__4_,r_n_2__3_,r_n_2__2_,
  r_n_2__1_,r_n_2__0_,r_n_1__31_,r_n_1__30_,r_n_1__29_,r_n_1__28_,r_n_1__27_,r_n_1__26_,
  r_n_1__25_,r_n_1__24_,r_n_1__23_,r_n_1__22_,r_n_1__21_,r_n_1__20_,r_n_1__19_,
  r_n_1__18_,r_n_1__17_,r_n_1__16_,r_n_1__15_,r_n_1__14_,r_n_1__13_,r_n_1__12_,
  r_n_1__11_,r_n_1__10_,r_n_1__9_,r_n_1__8_,r_n_1__7_,r_n_1__6_,r_n_1__5_,r_n_1__4_,
  r_n_1__3_,r_n_1__2_,r_n_1__1_,r_n_1__0_,r_n_32__31_,r_n_32__30_,r_n_32__29_,
  r_n_32__28_,r_n_32__27_,r_n_32__26_,r_n_32__25_,r_n_32__24_,r_n_32__23_,r_n_32__22_,
  r_n_32__21_,r_n_32__20_,r_n_32__19_,r_n_32__18_,r_n_32__17_,r_n_32__16_,r_n_32__15_,
  r_n_32__14_,r_n_32__13_,r_n_32__12_,r_n_32__11_,r_n_32__10_,r_n_32__9_,r_n_32__8_,
  r_n_32__7_,r_n_32__6_,r_n_32__5_,r_n_32__4_,r_n_32__3_,r_n_32__2_,r_n_32__1_,
  r_n_32__0_,r_n_31__31_,r_n_31__30_,r_n_31__29_,r_n_31__28_,r_n_31__27_,r_n_31__26_,
  r_n_31__25_,r_n_31__24_,r_n_31__23_,r_n_31__22_,r_n_31__21_,r_n_31__20_,
  r_n_31__19_,r_n_31__18_,r_n_31__17_,r_n_31__16_,r_n_31__15_,r_n_31__14_,r_n_31__13_,
  r_n_31__12_,r_n_31__11_,r_n_31__10_,r_n_31__9_,r_n_31__8_,r_n_31__7_,r_n_31__6_,
  r_n_31__5_,r_n_31__4_,r_n_31__3_,r_n_31__2_,r_n_31__1_,r_n_31__0_,r_n_30__31_,
  r_n_30__30_,r_n_30__29_,r_n_30__28_,r_n_30__27_,r_n_30__26_,r_n_30__25_,r_n_30__24_,
  r_n_30__23_,r_n_30__22_,r_n_30__21_,r_n_30__20_,r_n_30__19_,r_n_30__18_,
  r_n_30__17_,r_n_30__16_,r_n_30__15_,r_n_30__14_,r_n_30__13_,r_n_30__12_,r_n_30__11_,
  r_n_30__10_,r_n_30__9_,r_n_30__8_,r_n_30__7_,r_n_30__6_,r_n_30__5_,r_n_30__4_,
  r_n_30__3_,r_n_30__2_,r_n_30__1_,r_n_30__0_,r_n_29__31_,r_n_29__30_,r_n_29__29_,
  r_n_29__28_,r_n_29__27_,r_n_29__26_,r_n_29__25_,r_n_29__24_,r_n_29__23_,r_n_29__22_,
  r_n_29__21_,r_n_29__20_,r_n_29__19_,r_n_29__18_,r_n_29__17_,r_n_29__16_,r_n_29__15_,
  r_n_29__14_,r_n_29__13_,r_n_29__12_,r_n_29__11_,r_n_29__10_,r_n_29__9_,
  r_n_29__8_,r_n_29__7_,r_n_29__6_,r_n_29__5_,r_n_29__4_,r_n_29__3_,r_n_29__2_,r_n_29__1_,
  r_n_29__0_,r_n_28__31_,r_n_28__30_,r_n_28__29_,r_n_28__28_,r_n_28__27_,
  r_n_28__26_,r_n_28__25_,r_n_28__24_,r_n_28__23_,r_n_28__22_,r_n_28__21_,r_n_28__20_,
  r_n_28__19_,r_n_28__18_,r_n_28__17_,r_n_28__16_,r_n_28__15_,r_n_28__14_,r_n_28__13_,
  r_n_28__12_,r_n_28__11_,r_n_28__10_,r_n_28__9_,r_n_28__8_,r_n_28__7_,r_n_28__6_,
  r_n_28__5_,r_n_28__4_,r_n_28__3_,r_n_28__2_,r_n_28__1_,r_n_28__0_,r_n_27__31_,
  r_n_27__30_,r_n_27__29_,r_n_27__28_,r_n_27__27_,r_n_27__26_,r_n_27__25_,r_n_27__24_,
  r_n_27__23_,r_n_27__22_,r_n_27__21_,r_n_27__20_,r_n_27__19_,r_n_27__18_,
  r_n_27__17_,r_n_27__16_,r_n_27__15_,r_n_27__14_,r_n_27__13_,r_n_27__12_,r_n_27__11_,
  r_n_27__10_,r_n_27__9_,r_n_27__8_,r_n_27__7_,r_n_27__6_,r_n_27__5_,r_n_27__4_,
  r_n_27__3_,r_n_27__2_,r_n_27__1_,r_n_27__0_,r_n_26__31_,r_n_26__30_,r_n_26__29_,
  r_n_26__28_,r_n_26__27_,r_n_26__26_,r_n_26__25_,r_n_26__24_,r_n_26__23_,r_n_26__22_,
  r_n_26__21_,r_n_26__20_,r_n_26__19_,r_n_26__18_,r_n_26__17_,r_n_26__16_,
  r_n_26__15_,r_n_26__14_,r_n_26__13_,r_n_26__12_,r_n_26__11_,r_n_26__10_,r_n_26__9_,
  r_n_26__8_,r_n_26__7_,r_n_26__6_,r_n_26__5_,r_n_26__4_,r_n_26__3_,r_n_26__2_,r_n_26__1_,
  r_n_26__0_,r_n_25__31_,r_n_25__30_,r_n_25__29_,r_n_25__28_,r_n_25__27_,
  r_n_25__26_,r_n_25__25_,r_n_25__24_,r_n_25__23_,r_n_25__22_,r_n_25__21_,r_n_25__20_,
  r_n_25__19_,r_n_25__18_,r_n_25__17_,r_n_25__16_,r_n_25__15_,r_n_25__14_,r_n_25__13_,
  r_n_25__12_,r_n_25__11_,r_n_25__10_,r_n_25__9_,r_n_25__8_,r_n_25__7_,r_n_25__6_,
  r_n_25__5_,r_n_25__4_,r_n_25__3_,r_n_25__2_,r_n_25__1_,r_n_25__0_,r_n_24__31_,
  r_n_24__30_,r_n_24__29_,r_n_24__28_,r_n_24__27_,r_n_24__26_,r_n_24__25_,
  r_n_24__24_,r_n_24__23_,r_n_24__22_,r_n_24__21_,r_n_24__20_,r_n_24__19_,r_n_24__18_,
  r_n_24__17_,r_n_24__16_,r_n_24__15_,r_n_24__14_,r_n_24__13_,r_n_24__12_,r_n_24__11_,
  r_n_24__10_,r_n_24__9_,r_n_24__8_,r_n_24__7_,r_n_24__6_,r_n_24__5_,r_n_24__4_,
  r_n_24__3_,r_n_24__2_,r_n_24__1_,r_n_24__0_,r_n_23__31_,r_n_23__30_,r_n_23__29_,
  r_n_23__28_,r_n_23__27_,r_n_23__26_,r_n_23__25_,r_n_23__24_,r_n_23__23_,r_n_23__22_,
  r_n_23__21_,r_n_23__20_,r_n_23__19_,r_n_23__18_,r_n_23__17_,r_n_23__16_,
  r_n_23__15_,r_n_23__14_,r_n_23__13_,r_n_23__12_,r_n_23__11_,r_n_23__10_,r_n_23__9_,
  r_n_23__8_,r_n_23__7_,r_n_23__6_,r_n_23__5_,r_n_23__4_,r_n_23__3_,r_n_23__2_,
  r_n_23__1_,r_n_23__0_,r_n_22__31_,r_n_22__30_,r_n_22__29_,r_n_22__28_,r_n_22__27_,
  r_n_22__26_,r_n_22__25_,r_n_22__24_,r_n_22__23_,r_n_22__22_,r_n_22__21_,r_n_22__20_,
  r_n_22__19_,r_n_22__18_,r_n_22__17_,r_n_22__16_,r_n_22__15_,r_n_22__14_,
  r_n_22__13_,r_n_22__12_,r_n_22__11_,r_n_22__10_,r_n_22__9_,r_n_22__8_,r_n_22__7_,
  r_n_22__6_,r_n_22__5_,r_n_22__4_,r_n_22__3_,r_n_22__2_,r_n_22__1_,r_n_22__0_,r_n_21__31_,
  r_n_21__30_,r_n_21__29_,r_n_21__28_,r_n_21__27_,r_n_21__26_,r_n_21__25_,
  r_n_21__24_,r_n_21__23_,r_n_21__22_,r_n_21__21_,r_n_21__20_,r_n_21__19_,r_n_21__18_,
  r_n_21__17_,r_n_21__16_,r_n_21__15_,r_n_21__14_,r_n_21__13_,r_n_21__12_,r_n_21__11_,
  r_n_21__10_,r_n_21__9_,r_n_21__8_,r_n_21__7_,r_n_21__6_,r_n_21__5_,r_n_21__4_,
  r_n_21__3_,r_n_21__2_,r_n_21__1_,r_n_21__0_,r_n_20__31_,r_n_20__30_,r_n_20__29_,
  r_n_20__28_,r_n_20__27_,r_n_20__26_,r_n_20__25_,r_n_20__24_,r_n_20__23_,
  r_n_20__22_,r_n_20__21_,r_n_20__20_,r_n_20__19_,r_n_20__18_,r_n_20__17_,r_n_20__16_,
  r_n_20__15_,r_n_20__14_,r_n_20__13_,r_n_20__12_,r_n_20__11_,r_n_20__10_,r_n_20__9_,
  r_n_20__8_,r_n_20__7_,r_n_20__6_,r_n_20__5_,r_n_20__4_,r_n_20__3_,r_n_20__2_,
  r_n_20__1_,r_n_20__0_,r_n_19__31_,r_n_19__30_,r_n_19__29_,r_n_19__28_,r_n_19__27_,
  r_n_19__26_,r_n_19__25_,r_n_19__24_,r_n_19__23_,r_n_19__22_,r_n_19__21_,r_n_19__20_,
  r_n_19__19_,r_n_19__18_,r_n_19__17_,r_n_19__16_,r_n_19__15_,r_n_19__14_,
  r_n_19__13_,r_n_19__12_,r_n_19__11_,r_n_19__10_,r_n_19__9_,r_n_19__8_,r_n_19__7_,
  r_n_19__6_,r_n_19__5_,r_n_19__4_,r_n_19__3_,r_n_19__2_,r_n_19__1_,r_n_19__0_,
  r_n_18__31_,r_n_18__30_,r_n_18__29_,r_n_18__28_,r_n_18__27_,r_n_18__26_,r_n_18__25_,
  r_n_18__24_,r_n_18__23_,r_n_18__22_,r_n_18__21_,r_n_18__20_,r_n_18__19_,r_n_18__18_,
  r_n_18__17_,r_n_18__16_,r_n_18__15_,r_n_18__14_,r_n_18__13_,r_n_18__12_,
  r_n_18__11_,r_n_18__10_,r_n_18__9_,r_n_18__8_,r_n_18__7_,r_n_18__6_,r_n_18__5_,r_n_18__4_,
  r_n_18__3_,r_n_18__2_,r_n_18__1_,r_n_18__0_,r_n_17__31_,r_n_17__30_,r_n_17__29_,
  r_n_17__28_,r_n_17__27_,r_n_17__26_,r_n_17__25_,r_n_17__24_,r_n_17__23_,
  r_n_17__22_,r_n_17__21_,r_n_17__20_,r_n_17__19_,r_n_17__18_,r_n_17__17_,r_n_17__16_,
  r_n_17__15_,r_n_17__14_,r_n_17__13_,r_n_17__12_,r_n_17__11_,r_n_17__10_,r_n_17__9_,
  r_n_17__8_,r_n_17__7_,r_n_17__6_,r_n_17__5_,r_n_17__4_,r_n_17__3_,r_n_17__2_,
  r_n_17__1_,r_n_17__0_,r_n_48__31_,r_n_48__30_,r_n_48__29_,r_n_48__28_,r_n_48__27_,
  r_n_48__26_,r_n_48__25_,r_n_48__24_,r_n_48__23_,r_n_48__22_,r_n_48__21_,
  r_n_48__20_,r_n_48__19_,r_n_48__18_,r_n_48__17_,r_n_48__16_,r_n_48__15_,r_n_48__14_,
  r_n_48__13_,r_n_48__12_,r_n_48__11_,r_n_48__10_,r_n_48__9_,r_n_48__8_,r_n_48__7_,
  r_n_48__6_,r_n_48__5_,r_n_48__4_,r_n_48__3_,r_n_48__2_,r_n_48__1_,r_n_48__0_,
  r_n_47__31_,r_n_47__30_,r_n_47__29_,r_n_47__28_,r_n_47__27_,r_n_47__26_,r_n_47__25_,
  r_n_47__24_,r_n_47__23_,r_n_47__22_,r_n_47__21_,r_n_47__20_,r_n_47__19_,r_n_47__18_,
  r_n_47__17_,r_n_47__16_,r_n_47__15_,r_n_47__14_,r_n_47__13_,r_n_47__12_,
  r_n_47__11_,r_n_47__10_,r_n_47__9_,r_n_47__8_,r_n_47__7_,r_n_47__6_,r_n_47__5_,
  r_n_47__4_,r_n_47__3_,r_n_47__2_,r_n_47__1_,r_n_47__0_,r_n_46__31_,r_n_46__30_,
  r_n_46__29_,r_n_46__28_,r_n_46__27_,r_n_46__26_,r_n_46__25_,r_n_46__24_,r_n_46__23_,
  r_n_46__22_,r_n_46__21_,r_n_46__20_,r_n_46__19_,r_n_46__18_,r_n_46__17_,r_n_46__16_,
  r_n_46__15_,r_n_46__14_,r_n_46__13_,r_n_46__12_,r_n_46__11_,r_n_46__10_,r_n_46__9_,
  r_n_46__8_,r_n_46__7_,r_n_46__6_,r_n_46__5_,r_n_46__4_,r_n_46__3_,r_n_46__2_,
  r_n_46__1_,r_n_46__0_,r_n_45__31_,r_n_45__30_,r_n_45__29_,r_n_45__28_,r_n_45__27_,
  r_n_45__26_,r_n_45__25_,r_n_45__24_,r_n_45__23_,r_n_45__22_,r_n_45__21_,
  r_n_45__20_,r_n_45__19_,r_n_45__18_,r_n_45__17_,r_n_45__16_,r_n_45__15_,r_n_45__14_,
  r_n_45__13_,r_n_45__12_,r_n_45__11_,r_n_45__10_,r_n_45__9_,r_n_45__8_,r_n_45__7_,
  r_n_45__6_,r_n_45__5_,r_n_45__4_,r_n_45__3_,r_n_45__2_,r_n_45__1_,r_n_45__0_,
  r_n_44__31_,r_n_44__30_,r_n_44__29_,r_n_44__28_,r_n_44__27_,r_n_44__26_,r_n_44__25_,
  r_n_44__24_,r_n_44__23_,r_n_44__22_,r_n_44__21_,r_n_44__20_,r_n_44__19_,
  r_n_44__18_,r_n_44__17_,r_n_44__16_,r_n_44__15_,r_n_44__14_,r_n_44__13_,r_n_44__12_,
  r_n_44__11_,r_n_44__10_,r_n_44__9_,r_n_44__8_,r_n_44__7_,r_n_44__6_,r_n_44__5_,
  r_n_44__4_,r_n_44__3_,r_n_44__2_,r_n_44__1_,r_n_44__0_,r_n_43__31_,r_n_43__30_,
  r_n_43__29_,r_n_43__28_,r_n_43__27_,r_n_43__26_,r_n_43__25_,r_n_43__24_,r_n_43__23_,
  r_n_43__22_,r_n_43__21_,r_n_43__20_,r_n_43__19_,r_n_43__18_,r_n_43__17_,r_n_43__16_,
  r_n_43__15_,r_n_43__14_,r_n_43__13_,r_n_43__12_,r_n_43__11_,r_n_43__10_,
  r_n_43__9_,r_n_43__8_,r_n_43__7_,r_n_43__6_,r_n_43__5_,r_n_43__4_,r_n_43__3_,r_n_43__2_,
  r_n_43__1_,r_n_43__0_,r_n_42__31_,r_n_42__30_,r_n_42__29_,r_n_42__28_,
  r_n_42__27_,r_n_42__26_,r_n_42__25_,r_n_42__24_,r_n_42__23_,r_n_42__22_,r_n_42__21_,
  r_n_42__20_,r_n_42__19_,r_n_42__18_,r_n_42__17_,r_n_42__16_,r_n_42__15_,r_n_42__14_,
  r_n_42__13_,r_n_42__12_,r_n_42__11_,r_n_42__10_,r_n_42__9_,r_n_42__8_,r_n_42__7_,
  r_n_42__6_,r_n_42__5_,r_n_42__4_,r_n_42__3_,r_n_42__2_,r_n_42__1_,r_n_42__0_,
  r_n_41__31_,r_n_41__30_,r_n_41__29_,r_n_41__28_,r_n_41__27_,r_n_41__26_,r_n_41__25_,
  r_n_41__24_,r_n_41__23_,r_n_41__22_,r_n_41__21_,r_n_41__20_,r_n_41__19_,
  r_n_41__18_,r_n_41__17_,r_n_41__16_,r_n_41__15_,r_n_41__14_,r_n_41__13_,r_n_41__12_,
  r_n_41__11_,r_n_41__10_,r_n_41__9_,r_n_41__8_,r_n_41__7_,r_n_41__6_,r_n_41__5_,
  r_n_41__4_,r_n_41__3_,r_n_41__2_,r_n_41__1_,r_n_41__0_,r_n_40__31_,r_n_40__30_,
  r_n_40__29_,r_n_40__28_,r_n_40__27_,r_n_40__26_,r_n_40__25_,r_n_40__24_,r_n_40__23_,
  r_n_40__22_,r_n_40__21_,r_n_40__20_,r_n_40__19_,r_n_40__18_,r_n_40__17_,
  r_n_40__16_,r_n_40__15_,r_n_40__14_,r_n_40__13_,r_n_40__12_,r_n_40__11_,r_n_40__10_,
  r_n_40__9_,r_n_40__8_,r_n_40__7_,r_n_40__6_,r_n_40__5_,r_n_40__4_,r_n_40__3_,
  r_n_40__2_,r_n_40__1_,r_n_40__0_,r_n_39__31_,r_n_39__30_,r_n_39__29_,r_n_39__28_,
  r_n_39__27_,r_n_39__26_,r_n_39__25_,r_n_39__24_,r_n_39__23_,r_n_39__22_,r_n_39__21_,
  r_n_39__20_,r_n_39__19_,r_n_39__18_,r_n_39__17_,r_n_39__16_,r_n_39__15_,r_n_39__14_,
  r_n_39__13_,r_n_39__12_,r_n_39__11_,r_n_39__10_,r_n_39__9_,r_n_39__8_,r_n_39__7_,
  r_n_39__6_,r_n_39__5_,r_n_39__4_,r_n_39__3_,r_n_39__2_,r_n_39__1_,r_n_39__0_,
  r_n_38__31_,r_n_38__30_,r_n_38__29_,r_n_38__28_,r_n_38__27_,r_n_38__26_,
  r_n_38__25_,r_n_38__24_,r_n_38__23_,r_n_38__22_,r_n_38__21_,r_n_38__20_,r_n_38__19_,
  r_n_38__18_,r_n_38__17_,r_n_38__16_,r_n_38__15_,r_n_38__14_,r_n_38__13_,r_n_38__12_,
  r_n_38__11_,r_n_38__10_,r_n_38__9_,r_n_38__8_,r_n_38__7_,r_n_38__6_,r_n_38__5_,
  r_n_38__4_,r_n_38__3_,r_n_38__2_,r_n_38__1_,r_n_38__0_,r_n_37__31_,r_n_37__30_,
  r_n_37__29_,r_n_37__28_,r_n_37__27_,r_n_37__26_,r_n_37__25_,r_n_37__24_,r_n_37__23_,
  r_n_37__22_,r_n_37__21_,r_n_37__20_,r_n_37__19_,r_n_37__18_,r_n_37__17_,
  r_n_37__16_,r_n_37__15_,r_n_37__14_,r_n_37__13_,r_n_37__12_,r_n_37__11_,r_n_37__10_,
  r_n_37__9_,r_n_37__8_,r_n_37__7_,r_n_37__6_,r_n_37__5_,r_n_37__4_,r_n_37__3_,
  r_n_37__2_,r_n_37__1_,r_n_37__0_,r_n_36__31_,r_n_36__30_,r_n_36__29_,r_n_36__28_,
  r_n_36__27_,r_n_36__26_,r_n_36__25_,r_n_36__24_,r_n_36__23_,r_n_36__22_,r_n_36__21_,
  r_n_36__20_,r_n_36__19_,r_n_36__18_,r_n_36__17_,r_n_36__16_,r_n_36__15_,
  r_n_36__14_,r_n_36__13_,r_n_36__12_,r_n_36__11_,r_n_36__10_,r_n_36__9_,r_n_36__8_,
  r_n_36__7_,r_n_36__6_,r_n_36__5_,r_n_36__4_,r_n_36__3_,r_n_36__2_,r_n_36__1_,r_n_36__0_,
  r_n_35__31_,r_n_35__30_,r_n_35__29_,r_n_35__28_,r_n_35__27_,r_n_35__26_,
  r_n_35__25_,r_n_35__24_,r_n_35__23_,r_n_35__22_,r_n_35__21_,r_n_35__20_,r_n_35__19_,
  r_n_35__18_,r_n_35__17_,r_n_35__16_,r_n_35__15_,r_n_35__14_,r_n_35__13_,r_n_35__12_,
  r_n_35__11_,r_n_35__10_,r_n_35__9_,r_n_35__8_,r_n_35__7_,r_n_35__6_,r_n_35__5_,
  r_n_35__4_,r_n_35__3_,r_n_35__2_,r_n_35__1_,r_n_35__0_,r_n_34__31_,r_n_34__30_,
  r_n_34__29_,r_n_34__28_,r_n_34__27_,r_n_34__26_,r_n_34__25_,r_n_34__24_,
  r_n_34__23_,r_n_34__22_,r_n_34__21_,r_n_34__20_,r_n_34__19_,r_n_34__18_,r_n_34__17_,
  r_n_34__16_,r_n_34__15_,r_n_34__14_,r_n_34__13_,r_n_34__12_,r_n_34__11_,r_n_34__10_,
  r_n_34__9_,r_n_34__8_,r_n_34__7_,r_n_34__6_,r_n_34__5_,r_n_34__4_,r_n_34__3_,
  r_n_34__2_,r_n_34__1_,r_n_34__0_,r_n_33__31_,r_n_33__30_,r_n_33__29_,r_n_33__28_,
  r_n_33__27_,r_n_33__26_,r_n_33__25_,r_n_33__24_,r_n_33__23_,r_n_33__22_,r_n_33__21_,
  r_n_33__20_,r_n_33__19_,r_n_33__18_,r_n_33__17_,r_n_33__16_,r_n_33__15_,
  r_n_33__14_,r_n_33__13_,r_n_33__12_,r_n_33__11_,r_n_33__10_,r_n_33__9_,r_n_33__8_,
  r_n_33__7_,r_n_33__6_,r_n_33__5_,r_n_33__4_,r_n_33__3_,r_n_33__2_,r_n_33__1_,
  r_n_33__0_,r_n_64__31_,r_n_64__30_,r_n_64__29_,r_n_64__28_,r_n_64__27_,r_n_64__26_,
  r_n_64__25_,r_n_64__24_,r_n_64__23_,r_n_64__22_,r_n_64__21_,r_n_64__20_,r_n_64__19_,
  r_n_64__18_,r_n_64__17_,r_n_64__16_,r_n_64__15_,r_n_64__14_,r_n_64__13_,
  r_n_64__12_,r_n_64__11_,r_n_64__10_,r_n_64__9_,r_n_64__8_,r_n_64__7_,r_n_64__6_,r_n_64__5_,
  r_n_64__4_,r_n_64__3_,r_n_64__2_,r_n_64__1_,r_n_64__0_,r_n_63__31_,r_n_63__30_,
  r_n_63__29_,r_n_63__28_,r_n_63__27_,r_n_63__26_,r_n_63__25_,r_n_63__24_,
  r_n_63__23_,r_n_63__22_,r_n_63__21_,r_n_63__20_,r_n_63__19_,r_n_63__18_,r_n_63__17_,
  r_n_63__16_,r_n_63__15_,r_n_63__14_,r_n_63__13_,r_n_63__12_,r_n_63__11_,r_n_63__10_,
  r_n_63__9_,r_n_63__8_,r_n_63__7_,r_n_63__6_,r_n_63__5_,r_n_63__4_,r_n_63__3_,
  r_n_63__2_,r_n_63__1_,r_n_63__0_,r_n_62__31_,r_n_62__30_,r_n_62__29_,r_n_62__28_,
  r_n_62__27_,r_n_62__26_,r_n_62__25_,r_n_62__24_,r_n_62__23_,r_n_62__22_,
  r_n_62__21_,r_n_62__20_,r_n_62__19_,r_n_62__18_,r_n_62__17_,r_n_62__16_,r_n_62__15_,
  r_n_62__14_,r_n_62__13_,r_n_62__12_,r_n_62__11_,r_n_62__10_,r_n_62__9_,r_n_62__8_,
  r_n_62__7_,r_n_62__6_,r_n_62__5_,r_n_62__4_,r_n_62__3_,r_n_62__2_,r_n_62__1_,
  r_n_62__0_,r_n_61__31_,r_n_61__30_,r_n_61__29_,r_n_61__28_,r_n_61__27_,r_n_61__26_,
  r_n_61__25_,r_n_61__24_,r_n_61__23_,r_n_61__22_,r_n_61__21_,r_n_61__20_,r_n_61__19_,
  r_n_61__18_,r_n_61__17_,r_n_61__16_,r_n_61__15_,r_n_61__14_,r_n_61__13_,
  r_n_61__12_,r_n_61__11_,r_n_61__10_,r_n_61__9_,r_n_61__8_,r_n_61__7_,r_n_61__6_,
  r_n_61__5_,r_n_61__4_,r_n_61__3_,r_n_61__2_,r_n_61__1_,r_n_61__0_,r_n_60__31_,
  r_n_60__30_,r_n_60__29_,r_n_60__28_,r_n_60__27_,r_n_60__26_,r_n_60__25_,r_n_60__24_,
  r_n_60__23_,r_n_60__22_,r_n_60__21_,r_n_60__20_,r_n_60__19_,r_n_60__18_,r_n_60__17_,
  r_n_60__16_,r_n_60__15_,r_n_60__14_,r_n_60__13_,r_n_60__12_,r_n_60__11_,
  r_n_60__10_,r_n_60__9_,r_n_60__8_,r_n_60__7_,r_n_60__6_,r_n_60__5_,r_n_60__4_,r_n_60__3_,
  r_n_60__2_,r_n_60__1_,r_n_60__0_,r_n_59__31_,r_n_59__30_,r_n_59__29_,r_n_59__28_,
  r_n_59__27_,r_n_59__26_,r_n_59__25_,r_n_59__24_,r_n_59__23_,r_n_59__22_,
  r_n_59__21_,r_n_59__20_,r_n_59__19_,r_n_59__18_,r_n_59__17_,r_n_59__16_,r_n_59__15_,
  r_n_59__14_,r_n_59__13_,r_n_59__12_,r_n_59__11_,r_n_59__10_,r_n_59__9_,r_n_59__8_,
  r_n_59__7_,r_n_59__6_,r_n_59__5_,r_n_59__4_,r_n_59__3_,r_n_59__2_,r_n_59__1_,
  r_n_59__0_,r_n_58__31_,r_n_58__30_,r_n_58__29_,r_n_58__28_,r_n_58__27_,r_n_58__26_,
  r_n_58__25_,r_n_58__24_,r_n_58__23_,r_n_58__22_,r_n_58__21_,r_n_58__20_,
  r_n_58__19_,r_n_58__18_,r_n_58__17_,r_n_58__16_,r_n_58__15_,r_n_58__14_,r_n_58__13_,
  r_n_58__12_,r_n_58__11_,r_n_58__10_,r_n_58__9_,r_n_58__8_,r_n_58__7_,r_n_58__6_,
  r_n_58__5_,r_n_58__4_,r_n_58__3_,r_n_58__2_,r_n_58__1_,r_n_58__0_,r_n_57__31_,
  r_n_57__30_,r_n_57__29_,r_n_57__28_,r_n_57__27_,r_n_57__26_,r_n_57__25_,r_n_57__24_,
  r_n_57__23_,r_n_57__22_,r_n_57__21_,r_n_57__20_,r_n_57__19_,r_n_57__18_,r_n_57__17_,
  r_n_57__16_,r_n_57__15_,r_n_57__14_,r_n_57__13_,r_n_57__12_,r_n_57__11_,
  r_n_57__10_,r_n_57__9_,r_n_57__8_,r_n_57__7_,r_n_57__6_,r_n_57__5_,r_n_57__4_,r_n_57__3_,
  r_n_57__2_,r_n_57__1_,r_n_57__0_,r_n_56__31_,r_n_56__30_,r_n_56__29_,
  r_n_56__28_,r_n_56__27_,r_n_56__26_,r_n_56__25_,r_n_56__24_,r_n_56__23_,r_n_56__22_,
  r_n_56__21_,r_n_56__20_,r_n_56__19_,r_n_56__18_,r_n_56__17_,r_n_56__16_,r_n_56__15_,
  r_n_56__14_,r_n_56__13_,r_n_56__12_,r_n_56__11_,r_n_56__10_,r_n_56__9_,r_n_56__8_,
  r_n_56__7_,r_n_56__6_,r_n_56__5_,r_n_56__4_,r_n_56__3_,r_n_56__2_,r_n_56__1_,
  r_n_56__0_,r_n_55__31_,r_n_55__30_,r_n_55__29_,r_n_55__28_,r_n_55__27_,r_n_55__26_,
  r_n_55__25_,r_n_55__24_,r_n_55__23_,r_n_55__22_,r_n_55__21_,r_n_55__20_,
  r_n_55__19_,r_n_55__18_,r_n_55__17_,r_n_55__16_,r_n_55__15_,r_n_55__14_,r_n_55__13_,
  r_n_55__12_,r_n_55__11_,r_n_55__10_,r_n_55__9_,r_n_55__8_,r_n_55__7_,r_n_55__6_,
  r_n_55__5_,r_n_55__4_,r_n_55__3_,r_n_55__2_,r_n_55__1_,r_n_55__0_,r_n_54__31_,
  r_n_54__30_,r_n_54__29_,r_n_54__28_,r_n_54__27_,r_n_54__26_,r_n_54__25_,r_n_54__24_,
  r_n_54__23_,r_n_54__22_,r_n_54__21_,r_n_54__20_,r_n_54__19_,r_n_54__18_,
  r_n_54__17_,r_n_54__16_,r_n_54__15_,r_n_54__14_,r_n_54__13_,r_n_54__12_,r_n_54__11_,
  r_n_54__10_,r_n_54__9_,r_n_54__8_,r_n_54__7_,r_n_54__6_,r_n_54__5_,r_n_54__4_,
  r_n_54__3_,r_n_54__2_,r_n_54__1_,r_n_54__0_,r_n_53__31_,r_n_53__30_,r_n_53__29_,
  r_n_53__28_,r_n_53__27_,r_n_53__26_,r_n_53__25_,r_n_53__24_,r_n_53__23_,r_n_53__22_,
  r_n_53__21_,r_n_53__20_,r_n_53__19_,r_n_53__18_,r_n_53__17_,r_n_53__16_,r_n_53__15_,
  r_n_53__14_,r_n_53__13_,r_n_53__12_,r_n_53__11_,r_n_53__10_,r_n_53__9_,
  r_n_53__8_,r_n_53__7_,r_n_53__6_,r_n_53__5_,r_n_53__4_,r_n_53__3_,r_n_53__2_,r_n_53__1_,
  r_n_53__0_,r_n_52__31_,r_n_52__30_,r_n_52__29_,r_n_52__28_,r_n_52__27_,
  r_n_52__26_,r_n_52__25_,r_n_52__24_,r_n_52__23_,r_n_52__22_,r_n_52__21_,r_n_52__20_,
  r_n_52__19_,r_n_52__18_,r_n_52__17_,r_n_52__16_,r_n_52__15_,r_n_52__14_,r_n_52__13_,
  r_n_52__12_,r_n_52__11_,r_n_52__10_,r_n_52__9_,r_n_52__8_,r_n_52__7_,r_n_52__6_,
  r_n_52__5_,r_n_52__4_,r_n_52__3_,r_n_52__2_,r_n_52__1_,r_n_52__0_,r_n_51__31_,
  r_n_51__30_,r_n_51__29_,r_n_51__28_,r_n_51__27_,r_n_51__26_,r_n_51__25_,r_n_51__24_,
  r_n_51__23_,r_n_51__22_,r_n_51__21_,r_n_51__20_,r_n_51__19_,r_n_51__18_,
  r_n_51__17_,r_n_51__16_,r_n_51__15_,r_n_51__14_,r_n_51__13_,r_n_51__12_,r_n_51__11_,
  r_n_51__10_,r_n_51__9_,r_n_51__8_,r_n_51__7_,r_n_51__6_,r_n_51__5_,r_n_51__4_,
  r_n_51__3_,r_n_51__2_,r_n_51__1_,r_n_51__0_,r_n_50__31_,r_n_50__30_,r_n_50__29_,
  r_n_50__28_,r_n_50__27_,r_n_50__26_,r_n_50__25_,r_n_50__24_,r_n_50__23_,r_n_50__22_,
  r_n_50__21_,r_n_50__20_,r_n_50__19_,r_n_50__18_,r_n_50__17_,r_n_50__16_,
  r_n_50__15_,r_n_50__14_,r_n_50__13_,r_n_50__12_,r_n_50__11_,r_n_50__10_,r_n_50__9_,
  r_n_50__8_,r_n_50__7_,r_n_50__6_,r_n_50__5_,r_n_50__4_,r_n_50__3_,r_n_50__2_,r_n_50__1_,
  r_n_50__0_,r_n_49__31_,r_n_49__30_,r_n_49__29_,r_n_49__28_,r_n_49__27_,
  r_n_49__26_,r_n_49__25_,r_n_49__24_,r_n_49__23_,r_n_49__22_,r_n_49__21_,r_n_49__20_,
  r_n_49__19_,r_n_49__18_,r_n_49__17_,r_n_49__16_,r_n_49__15_,r_n_49__14_,r_n_49__13_,
  r_n_49__12_,r_n_49__11_,r_n_49__10_,r_n_49__9_,r_n_49__8_,r_n_49__7_,r_n_49__6_,
  r_n_49__5_,r_n_49__4_,r_n_49__3_,r_n_49__2_,r_n_49__1_,r_n_49__0_,r_n_80__31_,
  r_n_80__30_,r_n_80__29_,r_n_80__28_,r_n_80__27_,r_n_80__26_,r_n_80__25_,
  r_n_80__24_,r_n_80__23_,r_n_80__22_,r_n_80__21_,r_n_80__20_,r_n_80__19_,r_n_80__18_,
  r_n_80__17_,r_n_80__16_,r_n_80__15_,r_n_80__14_,r_n_80__13_,r_n_80__12_,r_n_80__11_,
  r_n_80__10_,r_n_80__9_,r_n_80__8_,r_n_80__7_,r_n_80__6_,r_n_80__5_,r_n_80__4_,
  r_n_80__3_,r_n_80__2_,r_n_80__1_,r_n_80__0_,r_n_79__31_,r_n_79__30_,r_n_79__29_,
  r_n_79__28_,r_n_79__27_,r_n_79__26_,r_n_79__25_,r_n_79__24_,r_n_79__23_,r_n_79__22_,
  r_n_79__21_,r_n_79__20_,r_n_79__19_,r_n_79__18_,r_n_79__17_,r_n_79__16_,
  r_n_79__15_,r_n_79__14_,r_n_79__13_,r_n_79__12_,r_n_79__11_,r_n_79__10_,r_n_79__9_,
  r_n_79__8_,r_n_79__7_,r_n_79__6_,r_n_79__5_,r_n_79__4_,r_n_79__3_,r_n_79__2_,
  r_n_79__1_,r_n_79__0_,r_n_78__31_,r_n_78__30_,r_n_78__29_,r_n_78__28_,r_n_78__27_,
  r_n_78__26_,r_n_78__25_,r_n_78__24_,r_n_78__23_,r_n_78__22_,r_n_78__21_,r_n_78__20_,
  r_n_78__19_,r_n_78__18_,r_n_78__17_,r_n_78__16_,r_n_78__15_,r_n_78__14_,
  r_n_78__13_,r_n_78__12_,r_n_78__11_,r_n_78__10_,r_n_78__9_,r_n_78__8_,r_n_78__7_,
  r_n_78__6_,r_n_78__5_,r_n_78__4_,r_n_78__3_,r_n_78__2_,r_n_78__1_,r_n_78__0_,r_n_77__31_,
  r_n_77__30_,r_n_77__29_,r_n_77__28_,r_n_77__27_,r_n_77__26_,r_n_77__25_,
  r_n_77__24_,r_n_77__23_,r_n_77__22_,r_n_77__21_,r_n_77__20_,r_n_77__19_,r_n_77__18_,
  r_n_77__17_,r_n_77__16_,r_n_77__15_,r_n_77__14_,r_n_77__13_,r_n_77__12_,r_n_77__11_,
  r_n_77__10_,r_n_77__9_,r_n_77__8_,r_n_77__7_,r_n_77__6_,r_n_77__5_,r_n_77__4_,
  r_n_77__3_,r_n_77__2_,r_n_77__1_,r_n_77__0_,r_n_76__31_,r_n_76__30_,r_n_76__29_,
  r_n_76__28_,r_n_76__27_,r_n_76__26_,r_n_76__25_,r_n_76__24_,r_n_76__23_,
  r_n_76__22_,r_n_76__21_,r_n_76__20_,r_n_76__19_,r_n_76__18_,r_n_76__17_,r_n_76__16_,
  r_n_76__15_,r_n_76__14_,r_n_76__13_,r_n_76__12_,r_n_76__11_,r_n_76__10_,r_n_76__9_,
  r_n_76__8_,r_n_76__7_,r_n_76__6_,r_n_76__5_,r_n_76__4_,r_n_76__3_,r_n_76__2_,
  r_n_76__1_,r_n_76__0_,r_n_75__31_,r_n_75__30_,r_n_75__29_,r_n_75__28_,r_n_75__27_,
  r_n_75__26_,r_n_75__25_,r_n_75__24_,r_n_75__23_,r_n_75__22_,r_n_75__21_,r_n_75__20_,
  r_n_75__19_,r_n_75__18_,r_n_75__17_,r_n_75__16_,r_n_75__15_,r_n_75__14_,
  r_n_75__13_,r_n_75__12_,r_n_75__11_,r_n_75__10_,r_n_75__9_,r_n_75__8_,r_n_75__7_,
  r_n_75__6_,r_n_75__5_,r_n_75__4_,r_n_75__3_,r_n_75__2_,r_n_75__1_,r_n_75__0_,
  r_n_74__31_,r_n_74__30_,r_n_74__29_,r_n_74__28_,r_n_74__27_,r_n_74__26_,r_n_74__25_,
  r_n_74__24_,r_n_74__23_,r_n_74__22_,r_n_74__21_,r_n_74__20_,r_n_74__19_,r_n_74__18_,
  r_n_74__17_,r_n_74__16_,r_n_74__15_,r_n_74__14_,r_n_74__13_,r_n_74__12_,
  r_n_74__11_,r_n_74__10_,r_n_74__9_,r_n_74__8_,r_n_74__7_,r_n_74__6_,r_n_74__5_,r_n_74__4_,
  r_n_74__3_,r_n_74__2_,r_n_74__1_,r_n_74__0_,r_n_73__31_,r_n_73__30_,r_n_73__29_,
  r_n_73__28_,r_n_73__27_,r_n_73__26_,r_n_73__25_,r_n_73__24_,r_n_73__23_,
  r_n_73__22_,r_n_73__21_,r_n_73__20_,r_n_73__19_,r_n_73__18_,r_n_73__17_,r_n_73__16_,
  r_n_73__15_,r_n_73__14_,r_n_73__13_,r_n_73__12_,r_n_73__11_,r_n_73__10_,r_n_73__9_,
  r_n_73__8_,r_n_73__7_,r_n_73__6_,r_n_73__5_,r_n_73__4_,r_n_73__3_,r_n_73__2_,
  r_n_73__1_,r_n_73__0_,r_n_72__31_,r_n_72__30_,r_n_72__29_,r_n_72__28_,r_n_72__27_,
  r_n_72__26_,r_n_72__25_,r_n_72__24_,r_n_72__23_,r_n_72__22_,r_n_72__21_,
  r_n_72__20_,r_n_72__19_,r_n_72__18_,r_n_72__17_,r_n_72__16_,r_n_72__15_,r_n_72__14_,
  r_n_72__13_,r_n_72__12_,r_n_72__11_,r_n_72__10_,r_n_72__9_,r_n_72__8_,r_n_72__7_,
  r_n_72__6_,r_n_72__5_,r_n_72__4_,r_n_72__3_,r_n_72__2_,r_n_72__1_,r_n_72__0_,
  r_n_71__31_,r_n_71__30_,r_n_71__29_,r_n_71__28_,r_n_71__27_,r_n_71__26_,r_n_71__25_,
  r_n_71__24_,r_n_71__23_,r_n_71__22_,r_n_71__21_,r_n_71__20_,r_n_71__19_,r_n_71__18_,
  r_n_71__17_,r_n_71__16_,r_n_71__15_,r_n_71__14_,r_n_71__13_,r_n_71__12_,
  r_n_71__11_,r_n_71__10_,r_n_71__9_,r_n_71__8_,r_n_71__7_,r_n_71__6_,r_n_71__5_,
  r_n_71__4_,r_n_71__3_,r_n_71__2_,r_n_71__1_,r_n_71__0_,r_n_70__31_,r_n_70__30_,
  r_n_70__29_,r_n_70__28_,r_n_70__27_,r_n_70__26_,r_n_70__25_,r_n_70__24_,r_n_70__23_,
  r_n_70__22_,r_n_70__21_,r_n_70__20_,r_n_70__19_,r_n_70__18_,r_n_70__17_,r_n_70__16_,
  r_n_70__15_,r_n_70__14_,r_n_70__13_,r_n_70__12_,r_n_70__11_,r_n_70__10_,r_n_70__9_,
  r_n_70__8_,r_n_70__7_,r_n_70__6_,r_n_70__5_,r_n_70__4_,r_n_70__3_,r_n_70__2_,
  r_n_70__1_,r_n_70__0_,r_n_69__31_,r_n_69__30_,r_n_69__29_,r_n_69__28_,r_n_69__27_,
  r_n_69__26_,r_n_69__25_,r_n_69__24_,r_n_69__23_,r_n_69__22_,r_n_69__21_,
  r_n_69__20_,r_n_69__19_,r_n_69__18_,r_n_69__17_,r_n_69__16_,r_n_69__15_,r_n_69__14_,
  r_n_69__13_,r_n_69__12_,r_n_69__11_,r_n_69__10_,r_n_69__9_,r_n_69__8_,r_n_69__7_,
  r_n_69__6_,r_n_69__5_,r_n_69__4_,r_n_69__3_,r_n_69__2_,r_n_69__1_,r_n_69__0_,
  r_n_68__31_,r_n_68__30_,r_n_68__29_,r_n_68__28_,r_n_68__27_,r_n_68__26_,r_n_68__25_,
  r_n_68__24_,r_n_68__23_,r_n_68__22_,r_n_68__21_,r_n_68__20_,r_n_68__19_,
  r_n_68__18_,r_n_68__17_,r_n_68__16_,r_n_68__15_,r_n_68__14_,r_n_68__13_,r_n_68__12_,
  r_n_68__11_,r_n_68__10_,r_n_68__9_,r_n_68__8_,r_n_68__7_,r_n_68__6_,r_n_68__5_,
  r_n_68__4_,r_n_68__3_,r_n_68__2_,r_n_68__1_,r_n_68__0_,r_n_67__31_,r_n_67__30_,
  r_n_67__29_,r_n_67__28_,r_n_67__27_,r_n_67__26_,r_n_67__25_,r_n_67__24_,r_n_67__23_,
  r_n_67__22_,r_n_67__21_,r_n_67__20_,r_n_67__19_,r_n_67__18_,r_n_67__17_,r_n_67__16_,
  r_n_67__15_,r_n_67__14_,r_n_67__13_,r_n_67__12_,r_n_67__11_,r_n_67__10_,
  r_n_67__9_,r_n_67__8_,r_n_67__7_,r_n_67__6_,r_n_67__5_,r_n_67__4_,r_n_67__3_,r_n_67__2_,
  r_n_67__1_,r_n_67__0_,r_n_66__31_,r_n_66__30_,r_n_66__29_,r_n_66__28_,
  r_n_66__27_,r_n_66__26_,r_n_66__25_,r_n_66__24_,r_n_66__23_,r_n_66__22_,r_n_66__21_,
  r_n_66__20_,r_n_66__19_,r_n_66__18_,r_n_66__17_,r_n_66__16_,r_n_66__15_,r_n_66__14_,
  r_n_66__13_,r_n_66__12_,r_n_66__11_,r_n_66__10_,r_n_66__9_,r_n_66__8_,r_n_66__7_,
  r_n_66__6_,r_n_66__5_,r_n_66__4_,r_n_66__3_,r_n_66__2_,r_n_66__1_,r_n_66__0_,
  r_n_65__31_,r_n_65__30_,r_n_65__29_,r_n_65__28_,r_n_65__27_,r_n_65__26_,r_n_65__25_,
  r_n_65__24_,r_n_65__23_,r_n_65__22_,r_n_65__21_,r_n_65__20_,r_n_65__19_,
  r_n_65__18_,r_n_65__17_,r_n_65__16_,r_n_65__15_,r_n_65__14_,r_n_65__13_,r_n_65__12_,
  r_n_65__11_,r_n_65__10_,r_n_65__9_,r_n_65__8_,r_n_65__7_,r_n_65__6_,r_n_65__5_,
  r_n_65__4_,r_n_65__3_,r_n_65__2_,r_n_65__1_,r_n_65__0_,r_n_96__31_,r_n_96__30_,
  r_n_96__29_,r_n_96__28_,r_n_96__27_,r_n_96__26_,r_n_96__25_,r_n_96__24_,r_n_96__23_,
  r_n_96__22_,r_n_96__21_,r_n_96__20_,r_n_96__19_,r_n_96__18_,r_n_96__17_,
  r_n_96__16_,r_n_96__15_,r_n_96__14_,r_n_96__13_,r_n_96__12_,r_n_96__11_,r_n_96__10_,
  r_n_96__9_,r_n_96__8_,r_n_96__7_,r_n_96__6_,r_n_96__5_,r_n_96__4_,r_n_96__3_,
  r_n_96__2_,r_n_96__1_,r_n_96__0_,r_n_95__31_,r_n_95__30_,r_n_95__29_,r_n_95__28_,
  r_n_95__27_,r_n_95__26_,r_n_95__25_,r_n_95__24_,r_n_95__23_,r_n_95__22_,r_n_95__21_,
  r_n_95__20_,r_n_95__19_,r_n_95__18_,r_n_95__17_,r_n_95__16_,r_n_95__15_,r_n_95__14_,
  r_n_95__13_,r_n_95__12_,r_n_95__11_,r_n_95__10_,r_n_95__9_,r_n_95__8_,r_n_95__7_,
  r_n_95__6_,r_n_95__5_,r_n_95__4_,r_n_95__3_,r_n_95__2_,r_n_95__1_,r_n_95__0_,
  r_n_94__31_,r_n_94__30_,r_n_94__29_,r_n_94__28_,r_n_94__27_,r_n_94__26_,
  r_n_94__25_,r_n_94__24_,r_n_94__23_,r_n_94__22_,r_n_94__21_,r_n_94__20_,r_n_94__19_,
  r_n_94__18_,r_n_94__17_,r_n_94__16_,r_n_94__15_,r_n_94__14_,r_n_94__13_,r_n_94__12_,
  r_n_94__11_,r_n_94__10_,r_n_94__9_,r_n_94__8_,r_n_94__7_,r_n_94__6_,r_n_94__5_,
  r_n_94__4_,r_n_94__3_,r_n_94__2_,r_n_94__1_,r_n_94__0_,r_n_93__31_,r_n_93__30_,
  r_n_93__29_,r_n_93__28_,r_n_93__27_,r_n_93__26_,r_n_93__25_,r_n_93__24_,r_n_93__23_,
  r_n_93__22_,r_n_93__21_,r_n_93__20_,r_n_93__19_,r_n_93__18_,r_n_93__17_,
  r_n_93__16_,r_n_93__15_,r_n_93__14_,r_n_93__13_,r_n_93__12_,r_n_93__11_,r_n_93__10_,
  r_n_93__9_,r_n_93__8_,r_n_93__7_,r_n_93__6_,r_n_93__5_,r_n_93__4_,r_n_93__3_,
  r_n_93__2_,r_n_93__1_,r_n_93__0_,r_n_92__31_,r_n_92__30_,r_n_92__29_,r_n_92__28_,
  r_n_92__27_,r_n_92__26_,r_n_92__25_,r_n_92__24_,r_n_92__23_,r_n_92__22_,r_n_92__21_,
  r_n_92__20_,r_n_92__19_,r_n_92__18_,r_n_92__17_,r_n_92__16_,r_n_92__15_,
  r_n_92__14_,r_n_92__13_,r_n_92__12_,r_n_92__11_,r_n_92__10_,r_n_92__9_,r_n_92__8_,
  r_n_92__7_,r_n_92__6_,r_n_92__5_,r_n_92__4_,r_n_92__3_,r_n_92__2_,r_n_92__1_,r_n_92__0_,
  r_n_91__31_,r_n_91__30_,r_n_91__29_,r_n_91__28_,r_n_91__27_,r_n_91__26_,
  r_n_91__25_,r_n_91__24_,r_n_91__23_,r_n_91__22_,r_n_91__21_,r_n_91__20_,r_n_91__19_,
  r_n_91__18_,r_n_91__17_,r_n_91__16_,r_n_91__15_,r_n_91__14_,r_n_91__13_,r_n_91__12_,
  r_n_91__11_,r_n_91__10_,r_n_91__9_,r_n_91__8_,r_n_91__7_,r_n_91__6_,r_n_91__5_,
  r_n_91__4_,r_n_91__3_,r_n_91__2_,r_n_91__1_,r_n_91__0_,r_n_90__31_,r_n_90__30_,
  r_n_90__29_,r_n_90__28_,r_n_90__27_,r_n_90__26_,r_n_90__25_,r_n_90__24_,
  r_n_90__23_,r_n_90__22_,r_n_90__21_,r_n_90__20_,r_n_90__19_,r_n_90__18_,r_n_90__17_,
  r_n_90__16_,r_n_90__15_,r_n_90__14_,r_n_90__13_,r_n_90__12_,r_n_90__11_,r_n_90__10_,
  r_n_90__9_,r_n_90__8_,r_n_90__7_,r_n_90__6_,r_n_90__5_,r_n_90__4_,r_n_90__3_,
  r_n_90__2_,r_n_90__1_,r_n_90__0_,r_n_89__31_,r_n_89__30_,r_n_89__29_,r_n_89__28_,
  r_n_89__27_,r_n_89__26_,r_n_89__25_,r_n_89__24_,r_n_89__23_,r_n_89__22_,r_n_89__21_,
  r_n_89__20_,r_n_89__19_,r_n_89__18_,r_n_89__17_,r_n_89__16_,r_n_89__15_,
  r_n_89__14_,r_n_89__13_,r_n_89__12_,r_n_89__11_,r_n_89__10_,r_n_89__9_,r_n_89__8_,
  r_n_89__7_,r_n_89__6_,r_n_89__5_,r_n_89__4_,r_n_89__3_,r_n_89__2_,r_n_89__1_,
  r_n_89__0_,r_n_88__31_,r_n_88__30_,r_n_88__29_,r_n_88__28_,r_n_88__27_,r_n_88__26_,
  r_n_88__25_,r_n_88__24_,r_n_88__23_,r_n_88__22_,r_n_88__21_,r_n_88__20_,r_n_88__19_,
  r_n_88__18_,r_n_88__17_,r_n_88__16_,r_n_88__15_,r_n_88__14_,r_n_88__13_,
  r_n_88__12_,r_n_88__11_,r_n_88__10_,r_n_88__9_,r_n_88__8_,r_n_88__7_,r_n_88__6_,r_n_88__5_,
  r_n_88__4_,r_n_88__3_,r_n_88__2_,r_n_88__1_,r_n_88__0_,r_n_87__31_,r_n_87__30_,
  r_n_87__29_,r_n_87__28_,r_n_87__27_,r_n_87__26_,r_n_87__25_,r_n_87__24_,
  r_n_87__23_,r_n_87__22_,r_n_87__21_,r_n_87__20_,r_n_87__19_,r_n_87__18_,r_n_87__17_,
  r_n_87__16_,r_n_87__15_,r_n_87__14_,r_n_87__13_,r_n_87__12_,r_n_87__11_,r_n_87__10_,
  r_n_87__9_,r_n_87__8_,r_n_87__7_,r_n_87__6_,r_n_87__5_,r_n_87__4_,r_n_87__3_,
  r_n_87__2_,r_n_87__1_,r_n_87__0_,r_n_86__31_,r_n_86__30_,r_n_86__29_,r_n_86__28_,
  r_n_86__27_,r_n_86__26_,r_n_86__25_,r_n_86__24_,r_n_86__23_,r_n_86__22_,
  r_n_86__21_,r_n_86__20_,r_n_86__19_,r_n_86__18_,r_n_86__17_,r_n_86__16_,r_n_86__15_,
  r_n_86__14_,r_n_86__13_,r_n_86__12_,r_n_86__11_,r_n_86__10_,r_n_86__9_,r_n_86__8_,
  r_n_86__7_,r_n_86__6_,r_n_86__5_,r_n_86__4_,r_n_86__3_,r_n_86__2_,r_n_86__1_,
  r_n_86__0_,r_n_85__31_,r_n_85__30_,r_n_85__29_,r_n_85__28_,r_n_85__27_,r_n_85__26_,
  r_n_85__25_,r_n_85__24_,r_n_85__23_,r_n_85__22_,r_n_85__21_,r_n_85__20_,r_n_85__19_,
  r_n_85__18_,r_n_85__17_,r_n_85__16_,r_n_85__15_,r_n_85__14_,r_n_85__13_,
  r_n_85__12_,r_n_85__11_,r_n_85__10_,r_n_85__9_,r_n_85__8_,r_n_85__7_,r_n_85__6_,
  r_n_85__5_,r_n_85__4_,r_n_85__3_,r_n_85__2_,r_n_85__1_,r_n_85__0_,r_n_84__31_,
  r_n_84__30_,r_n_84__29_,r_n_84__28_,r_n_84__27_,r_n_84__26_,r_n_84__25_,r_n_84__24_,
  r_n_84__23_,r_n_84__22_,r_n_84__21_,r_n_84__20_,r_n_84__19_,r_n_84__18_,r_n_84__17_,
  r_n_84__16_,r_n_84__15_,r_n_84__14_,r_n_84__13_,r_n_84__12_,r_n_84__11_,
  r_n_84__10_,r_n_84__9_,r_n_84__8_,r_n_84__7_,r_n_84__6_,r_n_84__5_,r_n_84__4_,r_n_84__3_,
  r_n_84__2_,r_n_84__1_,r_n_84__0_,r_n_83__31_,r_n_83__30_,r_n_83__29_,r_n_83__28_,
  r_n_83__27_,r_n_83__26_,r_n_83__25_,r_n_83__24_,r_n_83__23_,r_n_83__22_,
  r_n_83__21_,r_n_83__20_,r_n_83__19_,r_n_83__18_,r_n_83__17_,r_n_83__16_,r_n_83__15_,
  r_n_83__14_,r_n_83__13_,r_n_83__12_,r_n_83__11_,r_n_83__10_,r_n_83__9_,r_n_83__8_,
  r_n_83__7_,r_n_83__6_,r_n_83__5_,r_n_83__4_,r_n_83__3_,r_n_83__2_,r_n_83__1_,
  r_n_83__0_,r_n_82__31_,r_n_82__30_,r_n_82__29_,r_n_82__28_,r_n_82__27_,r_n_82__26_,
  r_n_82__25_,r_n_82__24_,r_n_82__23_,r_n_82__22_,r_n_82__21_,r_n_82__20_,
  r_n_82__19_,r_n_82__18_,r_n_82__17_,r_n_82__16_,r_n_82__15_,r_n_82__14_,r_n_82__13_,
  r_n_82__12_,r_n_82__11_,r_n_82__10_,r_n_82__9_,r_n_82__8_,r_n_82__7_,r_n_82__6_,
  r_n_82__5_,r_n_82__4_,r_n_82__3_,r_n_82__2_,r_n_82__1_,r_n_82__0_,r_n_81__31_,
  r_n_81__30_,r_n_81__29_,r_n_81__28_,r_n_81__27_,r_n_81__26_,r_n_81__25_,r_n_81__24_,
  r_n_81__23_,r_n_81__22_,r_n_81__21_,r_n_81__20_,r_n_81__19_,r_n_81__18_,r_n_81__17_,
  r_n_81__16_,r_n_81__15_,r_n_81__14_,r_n_81__13_,r_n_81__12_,r_n_81__11_,
  r_n_81__10_,r_n_81__9_,r_n_81__8_,r_n_81__7_,r_n_81__6_,r_n_81__5_,r_n_81__4_,r_n_81__3_,
  r_n_81__2_,r_n_81__1_,r_n_81__0_,r_n_112__31_,r_n_112__30_,r_n_112__29_,
  r_n_112__28_,r_n_112__27_,r_n_112__26_,r_n_112__25_,r_n_112__24_,r_n_112__23_,
  r_n_112__22_,r_n_112__21_,r_n_112__20_,r_n_112__19_,r_n_112__18_,r_n_112__17_,
  r_n_112__16_,r_n_112__15_,r_n_112__14_,r_n_112__13_,r_n_112__12_,r_n_112__11_,r_n_112__10_,
  r_n_112__9_,r_n_112__8_,r_n_112__7_,r_n_112__6_,r_n_112__5_,r_n_112__4_,
  r_n_112__3_,r_n_112__2_,r_n_112__1_,r_n_112__0_,r_n_111__31_,r_n_111__30_,r_n_111__29_,
  r_n_111__28_,r_n_111__27_,r_n_111__26_,r_n_111__25_,r_n_111__24_,r_n_111__23_,
  r_n_111__22_,r_n_111__21_,r_n_111__20_,r_n_111__19_,r_n_111__18_,r_n_111__17_,
  r_n_111__16_,r_n_111__15_,r_n_111__14_,r_n_111__13_,r_n_111__12_,r_n_111__11_,
  r_n_111__10_,r_n_111__9_,r_n_111__8_,r_n_111__7_,r_n_111__6_,r_n_111__5_,r_n_111__4_,
  r_n_111__3_,r_n_111__2_,r_n_111__1_,r_n_111__0_,r_n_110__31_,r_n_110__30_,
  r_n_110__29_,r_n_110__28_,r_n_110__27_,r_n_110__26_,r_n_110__25_,r_n_110__24_,
  r_n_110__23_,r_n_110__22_,r_n_110__21_,r_n_110__20_,r_n_110__19_,r_n_110__18_,r_n_110__17_,
  r_n_110__16_,r_n_110__15_,r_n_110__14_,r_n_110__13_,r_n_110__12_,r_n_110__11_,
  r_n_110__10_,r_n_110__9_,r_n_110__8_,r_n_110__7_,r_n_110__6_,r_n_110__5_,
  r_n_110__4_,r_n_110__3_,r_n_110__2_,r_n_110__1_,r_n_110__0_,r_n_109__31_,r_n_109__30_,
  r_n_109__29_,r_n_109__28_,r_n_109__27_,r_n_109__26_,r_n_109__25_,r_n_109__24_,
  r_n_109__23_,r_n_109__22_,r_n_109__21_,r_n_109__20_,r_n_109__19_,r_n_109__18_,
  r_n_109__17_,r_n_109__16_,r_n_109__15_,r_n_109__14_,r_n_109__13_,r_n_109__12_,
  r_n_109__11_,r_n_109__10_,r_n_109__9_,r_n_109__8_,r_n_109__7_,r_n_109__6_,r_n_109__5_,
  r_n_109__4_,r_n_109__3_,r_n_109__2_,r_n_109__1_,r_n_109__0_,r_n_108__31_,
  r_n_108__30_,r_n_108__29_,r_n_108__28_,r_n_108__27_,r_n_108__26_,r_n_108__25_,
  r_n_108__24_,r_n_108__23_,r_n_108__22_,r_n_108__21_,r_n_108__20_,r_n_108__19_,r_n_108__18_,
  r_n_108__17_,r_n_108__16_,r_n_108__15_,r_n_108__14_,r_n_108__13_,r_n_108__12_,
  r_n_108__11_,r_n_108__10_,r_n_108__9_,r_n_108__8_,r_n_108__7_,r_n_108__6_,
  r_n_108__5_,r_n_108__4_,r_n_108__3_,r_n_108__2_,r_n_108__1_,r_n_108__0_,r_n_107__31_,
  r_n_107__30_,r_n_107__29_,r_n_107__28_,r_n_107__27_,r_n_107__26_,r_n_107__25_,
  r_n_107__24_,r_n_107__23_,r_n_107__22_,r_n_107__21_,r_n_107__20_,r_n_107__19_,
  r_n_107__18_,r_n_107__17_,r_n_107__16_,r_n_107__15_,r_n_107__14_,r_n_107__13_,
  r_n_107__12_,r_n_107__11_,r_n_107__10_,r_n_107__9_,r_n_107__8_,r_n_107__7_,r_n_107__6_,
  r_n_107__5_,r_n_107__4_,r_n_107__3_,r_n_107__2_,r_n_107__1_,r_n_107__0_,
  r_n_106__31_,r_n_106__30_,r_n_106__29_,r_n_106__28_,r_n_106__27_,r_n_106__26_,r_n_106__25_,
  r_n_106__24_,r_n_106__23_,r_n_106__22_,r_n_106__21_,r_n_106__20_,r_n_106__19_,
  r_n_106__18_,r_n_106__17_,r_n_106__16_,r_n_106__15_,r_n_106__14_,r_n_106__13_,
  r_n_106__12_,r_n_106__11_,r_n_106__10_,r_n_106__9_,r_n_106__8_,r_n_106__7_,
  r_n_106__6_,r_n_106__5_,r_n_106__4_,r_n_106__3_,r_n_106__2_,r_n_106__1_,r_n_106__0_,
  r_n_105__31_,r_n_105__30_,r_n_105__29_,r_n_105__28_,r_n_105__27_,r_n_105__26_,
  r_n_105__25_,r_n_105__24_,r_n_105__23_,r_n_105__22_,r_n_105__21_,r_n_105__20_,
  r_n_105__19_,r_n_105__18_,r_n_105__17_,r_n_105__16_,r_n_105__15_,r_n_105__14_,
  r_n_105__13_,r_n_105__12_,r_n_105__11_,r_n_105__10_,r_n_105__9_,r_n_105__8_,r_n_105__7_,
  r_n_105__6_,r_n_105__5_,r_n_105__4_,r_n_105__3_,r_n_105__2_,r_n_105__1_,
  r_n_105__0_,r_n_104__31_,r_n_104__30_,r_n_104__29_,r_n_104__28_,r_n_104__27_,r_n_104__26_,
  r_n_104__25_,r_n_104__24_,r_n_104__23_,r_n_104__22_,r_n_104__21_,r_n_104__20_,
  r_n_104__19_,r_n_104__18_,r_n_104__17_,r_n_104__16_,r_n_104__15_,r_n_104__14_,
  r_n_104__13_,r_n_104__12_,r_n_104__11_,r_n_104__10_,r_n_104__9_,r_n_104__8_,
  r_n_104__7_,r_n_104__6_,r_n_104__5_,r_n_104__4_,r_n_104__3_,r_n_104__2_,r_n_104__1_,
  r_n_104__0_,r_n_103__31_,r_n_103__30_,r_n_103__29_,r_n_103__28_,r_n_103__27_,
  r_n_103__26_,r_n_103__25_,r_n_103__24_,r_n_103__23_,r_n_103__22_,r_n_103__21_,
  r_n_103__20_,r_n_103__19_,r_n_103__18_,r_n_103__17_,r_n_103__16_,r_n_103__15_,
  r_n_103__14_,r_n_103__13_,r_n_103__12_,r_n_103__11_,r_n_103__10_,r_n_103__9_,r_n_103__8_,
  r_n_103__7_,r_n_103__6_,r_n_103__5_,r_n_103__4_,r_n_103__3_,r_n_103__2_,
  r_n_103__1_,r_n_103__0_,r_n_102__31_,r_n_102__30_,r_n_102__29_,r_n_102__28_,r_n_102__27_,
  r_n_102__26_,r_n_102__25_,r_n_102__24_,r_n_102__23_,r_n_102__22_,r_n_102__21_,
  r_n_102__20_,r_n_102__19_,r_n_102__18_,r_n_102__17_,r_n_102__16_,r_n_102__15_,
  r_n_102__14_,r_n_102__13_,r_n_102__12_,r_n_102__11_,r_n_102__10_,r_n_102__9_,
  r_n_102__8_,r_n_102__7_,r_n_102__6_,r_n_102__5_,r_n_102__4_,r_n_102__3_,r_n_102__2_,
  r_n_102__1_,r_n_102__0_,r_n_101__31_,r_n_101__30_,r_n_101__29_,r_n_101__28_,
  r_n_101__27_,r_n_101__26_,r_n_101__25_,r_n_101__24_,r_n_101__23_,r_n_101__22_,
  r_n_101__21_,r_n_101__20_,r_n_101__19_,r_n_101__18_,r_n_101__17_,r_n_101__16_,r_n_101__15_,
  r_n_101__14_,r_n_101__13_,r_n_101__12_,r_n_101__11_,r_n_101__10_,r_n_101__9_,
  r_n_101__8_,r_n_101__7_,r_n_101__6_,r_n_101__5_,r_n_101__4_,r_n_101__3_,
  r_n_101__2_,r_n_101__1_,r_n_101__0_,r_n_100__31_,r_n_100__30_,r_n_100__29_,r_n_100__28_,
  r_n_100__27_,r_n_100__26_,r_n_100__25_,r_n_100__24_,r_n_100__23_,r_n_100__22_,
  r_n_100__21_,r_n_100__20_,r_n_100__19_,r_n_100__18_,r_n_100__17_,r_n_100__16_,
  r_n_100__15_,r_n_100__14_,r_n_100__13_,r_n_100__12_,r_n_100__11_,r_n_100__10_,
  r_n_100__9_,r_n_100__8_,r_n_100__7_,r_n_100__6_,r_n_100__5_,r_n_100__4_,r_n_100__3_,
  r_n_100__2_,r_n_100__1_,r_n_100__0_,r_n_99__31_,r_n_99__30_,r_n_99__29_,r_n_99__28_,
  r_n_99__27_,r_n_99__26_,r_n_99__25_,r_n_99__24_,r_n_99__23_,r_n_99__22_,
  r_n_99__21_,r_n_99__20_,r_n_99__19_,r_n_99__18_,r_n_99__17_,r_n_99__16_,r_n_99__15_,
  r_n_99__14_,r_n_99__13_,r_n_99__12_,r_n_99__11_,r_n_99__10_,r_n_99__9_,r_n_99__8_,
  r_n_99__7_,r_n_99__6_,r_n_99__5_,r_n_99__4_,r_n_99__3_,r_n_99__2_,r_n_99__1_,
  r_n_99__0_,r_n_98__31_,r_n_98__30_,r_n_98__29_,r_n_98__28_,r_n_98__27_,r_n_98__26_,
  r_n_98__25_,r_n_98__24_,r_n_98__23_,r_n_98__22_,r_n_98__21_,r_n_98__20_,
  r_n_98__19_,r_n_98__18_,r_n_98__17_,r_n_98__16_,r_n_98__15_,r_n_98__14_,r_n_98__13_,
  r_n_98__12_,r_n_98__11_,r_n_98__10_,r_n_98__9_,r_n_98__8_,r_n_98__7_,r_n_98__6_,
  r_n_98__5_,r_n_98__4_,r_n_98__3_,r_n_98__2_,r_n_98__1_,r_n_98__0_,r_n_97__31_,
  r_n_97__30_,r_n_97__29_,r_n_97__28_,r_n_97__27_,r_n_97__26_,r_n_97__25_,r_n_97__24_,
  r_n_97__23_,r_n_97__22_,r_n_97__21_,r_n_97__20_,r_n_97__19_,r_n_97__18_,r_n_97__17_,
  r_n_97__16_,r_n_97__15_,r_n_97__14_,r_n_97__13_,r_n_97__12_,r_n_97__11_,
  r_n_97__10_,r_n_97__9_,r_n_97__8_,r_n_97__7_,r_n_97__6_,r_n_97__5_,r_n_97__4_,r_n_97__3_,
  r_n_97__2_,r_n_97__1_,r_n_97__0_,r_n_128__31_,r_n_128__30_,r_n_128__29_,
  r_n_128__28_,r_n_128__27_,r_n_128__26_,r_n_128__25_,r_n_128__24_,r_n_128__23_,
  r_n_128__22_,r_n_128__21_,r_n_128__20_,r_n_128__19_,r_n_128__18_,r_n_128__17_,
  r_n_128__16_,r_n_128__15_,r_n_128__14_,r_n_128__13_,r_n_128__12_,r_n_128__11_,r_n_128__10_,
  r_n_128__9_,r_n_128__8_,r_n_128__7_,r_n_128__6_,r_n_128__5_,r_n_128__4_,
  r_n_128__3_,r_n_128__2_,r_n_128__1_,r_n_128__0_,r_n_127__31_,r_n_127__30_,r_n_127__29_,
  r_n_127__28_,r_n_127__27_,r_n_127__26_,r_n_127__25_,r_n_127__24_,r_n_127__23_,
  r_n_127__22_,r_n_127__21_,r_n_127__20_,r_n_127__19_,r_n_127__18_,r_n_127__17_,
  r_n_127__16_,r_n_127__15_,r_n_127__14_,r_n_127__13_,r_n_127__12_,r_n_127__11_,
  r_n_127__10_,r_n_127__9_,r_n_127__8_,r_n_127__7_,r_n_127__6_,r_n_127__5_,r_n_127__4_,
  r_n_127__3_,r_n_127__2_,r_n_127__1_,r_n_127__0_,r_n_126__31_,r_n_126__30_,
  r_n_126__29_,r_n_126__28_,r_n_126__27_,r_n_126__26_,r_n_126__25_,r_n_126__24_,
  r_n_126__23_,r_n_126__22_,r_n_126__21_,r_n_126__20_,r_n_126__19_,r_n_126__18_,r_n_126__17_,
  r_n_126__16_,r_n_126__15_,r_n_126__14_,r_n_126__13_,r_n_126__12_,r_n_126__11_,
  r_n_126__10_,r_n_126__9_,r_n_126__8_,r_n_126__7_,r_n_126__6_,r_n_126__5_,
  r_n_126__4_,r_n_126__3_,r_n_126__2_,r_n_126__1_,r_n_126__0_,r_n_125__31_,r_n_125__30_,
  r_n_125__29_,r_n_125__28_,r_n_125__27_,r_n_125__26_,r_n_125__25_,r_n_125__24_,
  r_n_125__23_,r_n_125__22_,r_n_125__21_,r_n_125__20_,r_n_125__19_,r_n_125__18_,
  r_n_125__17_,r_n_125__16_,r_n_125__15_,r_n_125__14_,r_n_125__13_,r_n_125__12_,
  r_n_125__11_,r_n_125__10_,r_n_125__9_,r_n_125__8_,r_n_125__7_,r_n_125__6_,r_n_125__5_,
  r_n_125__4_,r_n_125__3_,r_n_125__2_,r_n_125__1_,r_n_125__0_,r_n_124__31_,
  r_n_124__30_,r_n_124__29_,r_n_124__28_,r_n_124__27_,r_n_124__26_,r_n_124__25_,
  r_n_124__24_,r_n_124__23_,r_n_124__22_,r_n_124__21_,r_n_124__20_,r_n_124__19_,r_n_124__18_,
  r_n_124__17_,r_n_124__16_,r_n_124__15_,r_n_124__14_,r_n_124__13_,r_n_124__12_,
  r_n_124__11_,r_n_124__10_,r_n_124__9_,r_n_124__8_,r_n_124__7_,r_n_124__6_,
  r_n_124__5_,r_n_124__4_,r_n_124__3_,r_n_124__2_,r_n_124__1_,r_n_124__0_,r_n_123__31_,
  r_n_123__30_,r_n_123__29_,r_n_123__28_,r_n_123__27_,r_n_123__26_,r_n_123__25_,
  r_n_123__24_,r_n_123__23_,r_n_123__22_,r_n_123__21_,r_n_123__20_,r_n_123__19_,
  r_n_123__18_,r_n_123__17_,r_n_123__16_,r_n_123__15_,r_n_123__14_,r_n_123__13_,
  r_n_123__12_,r_n_123__11_,r_n_123__10_,r_n_123__9_,r_n_123__8_,r_n_123__7_,r_n_123__6_,
  r_n_123__5_,r_n_123__4_,r_n_123__3_,r_n_123__2_,r_n_123__1_,r_n_123__0_,
  r_n_122__31_,r_n_122__30_,r_n_122__29_,r_n_122__28_,r_n_122__27_,r_n_122__26_,r_n_122__25_,
  r_n_122__24_,r_n_122__23_,r_n_122__22_,r_n_122__21_,r_n_122__20_,r_n_122__19_,
  r_n_122__18_,r_n_122__17_,r_n_122__16_,r_n_122__15_,r_n_122__14_,r_n_122__13_,
  r_n_122__12_,r_n_122__11_,r_n_122__10_,r_n_122__9_,r_n_122__8_,r_n_122__7_,
  r_n_122__6_,r_n_122__5_,r_n_122__4_,r_n_122__3_,r_n_122__2_,r_n_122__1_,r_n_122__0_,
  r_n_121__31_,r_n_121__30_,r_n_121__29_,r_n_121__28_,r_n_121__27_,r_n_121__26_,
  r_n_121__25_,r_n_121__24_,r_n_121__23_,r_n_121__22_,r_n_121__21_,r_n_121__20_,
  r_n_121__19_,r_n_121__18_,r_n_121__17_,r_n_121__16_,r_n_121__15_,r_n_121__14_,
  r_n_121__13_,r_n_121__12_,r_n_121__11_,r_n_121__10_,r_n_121__9_,r_n_121__8_,r_n_121__7_,
  r_n_121__6_,r_n_121__5_,r_n_121__4_,r_n_121__3_,r_n_121__2_,r_n_121__1_,
  r_n_121__0_,r_n_120__31_,r_n_120__30_,r_n_120__29_,r_n_120__28_,r_n_120__27_,r_n_120__26_,
  r_n_120__25_,r_n_120__24_,r_n_120__23_,r_n_120__22_,r_n_120__21_,r_n_120__20_,
  r_n_120__19_,r_n_120__18_,r_n_120__17_,r_n_120__16_,r_n_120__15_,r_n_120__14_,
  r_n_120__13_,r_n_120__12_,r_n_120__11_,r_n_120__10_,r_n_120__9_,r_n_120__8_,
  r_n_120__7_,r_n_120__6_,r_n_120__5_,r_n_120__4_,r_n_120__3_,r_n_120__2_,r_n_120__1_,
  r_n_120__0_,r_n_119__31_,r_n_119__30_,r_n_119__29_,r_n_119__28_,r_n_119__27_,
  r_n_119__26_,r_n_119__25_,r_n_119__24_,r_n_119__23_,r_n_119__22_,r_n_119__21_,
  r_n_119__20_,r_n_119__19_,r_n_119__18_,r_n_119__17_,r_n_119__16_,r_n_119__15_,
  r_n_119__14_,r_n_119__13_,r_n_119__12_,r_n_119__11_,r_n_119__10_,r_n_119__9_,r_n_119__8_,
  r_n_119__7_,r_n_119__6_,r_n_119__5_,r_n_119__4_,r_n_119__3_,r_n_119__2_,
  r_n_119__1_,r_n_119__0_,r_n_118__31_,r_n_118__30_,r_n_118__29_,r_n_118__28_,r_n_118__27_,
  r_n_118__26_,r_n_118__25_,r_n_118__24_,r_n_118__23_,r_n_118__22_,r_n_118__21_,
  r_n_118__20_,r_n_118__19_,r_n_118__18_,r_n_118__17_,r_n_118__16_,r_n_118__15_,
  r_n_118__14_,r_n_118__13_,r_n_118__12_,r_n_118__11_,r_n_118__10_,r_n_118__9_,
  r_n_118__8_,r_n_118__7_,r_n_118__6_,r_n_118__5_,r_n_118__4_,r_n_118__3_,r_n_118__2_,
  r_n_118__1_,r_n_118__0_,r_n_117__31_,r_n_117__30_,r_n_117__29_,r_n_117__28_,
  r_n_117__27_,r_n_117__26_,r_n_117__25_,r_n_117__24_,r_n_117__23_,r_n_117__22_,
  r_n_117__21_,r_n_117__20_,r_n_117__19_,r_n_117__18_,r_n_117__17_,r_n_117__16_,r_n_117__15_,
  r_n_117__14_,r_n_117__13_,r_n_117__12_,r_n_117__11_,r_n_117__10_,r_n_117__9_,
  r_n_117__8_,r_n_117__7_,r_n_117__6_,r_n_117__5_,r_n_117__4_,r_n_117__3_,
  r_n_117__2_,r_n_117__1_,r_n_117__0_,r_n_116__31_,r_n_116__30_,r_n_116__29_,r_n_116__28_,
  r_n_116__27_,r_n_116__26_,r_n_116__25_,r_n_116__24_,r_n_116__23_,r_n_116__22_,
  r_n_116__21_,r_n_116__20_,r_n_116__19_,r_n_116__18_,r_n_116__17_,r_n_116__16_,
  r_n_116__15_,r_n_116__14_,r_n_116__13_,r_n_116__12_,r_n_116__11_,r_n_116__10_,
  r_n_116__9_,r_n_116__8_,r_n_116__7_,r_n_116__6_,r_n_116__5_,r_n_116__4_,r_n_116__3_,
  r_n_116__2_,r_n_116__1_,r_n_116__0_,r_n_115__31_,r_n_115__30_,r_n_115__29_,
  r_n_115__28_,r_n_115__27_,r_n_115__26_,r_n_115__25_,r_n_115__24_,r_n_115__23_,
  r_n_115__22_,r_n_115__21_,r_n_115__20_,r_n_115__19_,r_n_115__18_,r_n_115__17_,r_n_115__16_,
  r_n_115__15_,r_n_115__14_,r_n_115__13_,r_n_115__12_,r_n_115__11_,r_n_115__10_,
  r_n_115__9_,r_n_115__8_,r_n_115__7_,r_n_115__6_,r_n_115__5_,r_n_115__4_,
  r_n_115__3_,r_n_115__2_,r_n_115__1_,r_n_115__0_,r_n_114__31_,r_n_114__30_,r_n_114__29_,
  r_n_114__28_,r_n_114__27_,r_n_114__26_,r_n_114__25_,r_n_114__24_,r_n_114__23_,
  r_n_114__22_,r_n_114__21_,r_n_114__20_,r_n_114__19_,r_n_114__18_,r_n_114__17_,
  r_n_114__16_,r_n_114__15_,r_n_114__14_,r_n_114__13_,r_n_114__12_,r_n_114__11_,
  r_n_114__10_,r_n_114__9_,r_n_114__8_,r_n_114__7_,r_n_114__6_,r_n_114__5_,r_n_114__4_,
  r_n_114__3_,r_n_114__2_,r_n_114__1_,r_n_114__0_,r_n_113__31_,r_n_113__30_,
  r_n_113__29_,r_n_113__28_,r_n_113__27_,r_n_113__26_,r_n_113__25_,r_n_113__24_,r_n_113__23_,
  r_n_113__22_,r_n_113__21_,r_n_113__20_,r_n_113__19_,r_n_113__18_,r_n_113__17_,
  r_n_113__16_,r_n_113__15_,r_n_113__14_,r_n_113__13_,r_n_113__12_,r_n_113__11_,
  r_n_113__10_,r_n_113__9_,r_n_113__8_,r_n_113__7_,r_n_113__6_,r_n_113__5_,
  r_n_113__4_,r_n_113__3_,r_n_113__2_,r_n_113__1_,r_n_113__0_,r_n_144__31_,r_n_144__30_,
  r_n_144__29_,r_n_144__28_,r_n_144__27_,r_n_144__26_,r_n_144__25_,r_n_144__24_,
  r_n_144__23_,r_n_144__22_,r_n_144__21_,r_n_144__20_,r_n_144__19_,r_n_144__18_,
  r_n_144__17_,r_n_144__16_,r_n_144__15_,r_n_144__14_,r_n_144__13_,r_n_144__12_,
  r_n_144__11_,r_n_144__10_,r_n_144__9_,r_n_144__8_,r_n_144__7_,r_n_144__6_,r_n_144__5_,
  r_n_144__4_,r_n_144__3_,r_n_144__2_,r_n_144__1_,r_n_144__0_,r_n_143__31_,
  r_n_143__30_,r_n_143__29_,r_n_143__28_,r_n_143__27_,r_n_143__26_,r_n_143__25_,r_n_143__24_,
  r_n_143__23_,r_n_143__22_,r_n_143__21_,r_n_143__20_,r_n_143__19_,r_n_143__18_,
  r_n_143__17_,r_n_143__16_,r_n_143__15_,r_n_143__14_,r_n_143__13_,r_n_143__12_,
  r_n_143__11_,r_n_143__10_,r_n_143__9_,r_n_143__8_,r_n_143__7_,r_n_143__6_,
  r_n_143__5_,r_n_143__4_,r_n_143__3_,r_n_143__2_,r_n_143__1_,r_n_143__0_,r_n_142__31_,
  r_n_142__30_,r_n_142__29_,r_n_142__28_,r_n_142__27_,r_n_142__26_,r_n_142__25_,
  r_n_142__24_,r_n_142__23_,r_n_142__22_,r_n_142__21_,r_n_142__20_,r_n_142__19_,
  r_n_142__18_,r_n_142__17_,r_n_142__16_,r_n_142__15_,r_n_142__14_,r_n_142__13_,
  r_n_142__12_,r_n_142__11_,r_n_142__10_,r_n_142__9_,r_n_142__8_,r_n_142__7_,r_n_142__6_,
  r_n_142__5_,r_n_142__4_,r_n_142__3_,r_n_142__2_,r_n_142__1_,r_n_142__0_,r_n_141__31_,
  r_n_141__30_,r_n_141__29_,r_n_141__28_,r_n_141__27_,r_n_141__26_,r_n_141__25_,
  r_n_141__24_,r_n_141__23_,r_n_141__22_,r_n_141__21_,r_n_141__20_,r_n_141__19_,
  r_n_141__18_,r_n_141__17_,r_n_141__16_,r_n_141__15_,r_n_141__14_,r_n_141__13_,
  r_n_141__12_,r_n_141__11_,r_n_141__10_,r_n_141__9_,r_n_141__8_,r_n_141__7_,
  r_n_141__6_,r_n_141__5_,r_n_141__4_,r_n_141__3_,r_n_141__2_,r_n_141__1_,r_n_141__0_,
  r_n_140__31_,r_n_140__30_,r_n_140__29_,r_n_140__28_,r_n_140__27_,r_n_140__26_,
  r_n_140__25_,r_n_140__24_,r_n_140__23_,r_n_140__22_,r_n_140__21_,r_n_140__20_,
  r_n_140__19_,r_n_140__18_,r_n_140__17_,r_n_140__16_,r_n_140__15_,r_n_140__14_,r_n_140__13_,
  r_n_140__12_,r_n_140__11_,r_n_140__10_,r_n_140__9_,r_n_140__8_,r_n_140__7_,
  r_n_140__6_,r_n_140__5_,r_n_140__4_,r_n_140__3_,r_n_140__2_,r_n_140__1_,r_n_140__0_,
  r_n_139__31_,r_n_139__30_,r_n_139__29_,r_n_139__28_,r_n_139__27_,r_n_139__26_,
  r_n_139__25_,r_n_139__24_,r_n_139__23_,r_n_139__22_,r_n_139__21_,r_n_139__20_,
  r_n_139__19_,r_n_139__18_,r_n_139__17_,r_n_139__16_,r_n_139__15_,r_n_139__14_,
  r_n_139__13_,r_n_139__12_,r_n_139__11_,r_n_139__10_,r_n_139__9_,r_n_139__8_,
  r_n_139__7_,r_n_139__6_,r_n_139__5_,r_n_139__4_,r_n_139__3_,r_n_139__2_,r_n_139__1_,
  r_n_139__0_,r_n_138__31_,r_n_138__30_,r_n_138__29_,r_n_138__28_,r_n_138__27_,
  r_n_138__26_,r_n_138__25_,r_n_138__24_,r_n_138__23_,r_n_138__22_,r_n_138__21_,
  r_n_138__20_,r_n_138__19_,r_n_138__18_,r_n_138__17_,r_n_138__16_,r_n_138__15_,r_n_138__14_,
  r_n_138__13_,r_n_138__12_,r_n_138__11_,r_n_138__10_,r_n_138__9_,r_n_138__8_,
  r_n_138__7_,r_n_138__6_,r_n_138__5_,r_n_138__4_,r_n_138__3_,r_n_138__2_,r_n_138__1_,
  r_n_138__0_,r_n_137__31_,r_n_137__30_,r_n_137__29_,r_n_137__28_,r_n_137__27_,
  r_n_137__26_,r_n_137__25_,r_n_137__24_,r_n_137__23_,r_n_137__22_,r_n_137__21_,
  r_n_137__20_,r_n_137__19_,r_n_137__18_,r_n_137__17_,r_n_137__16_,r_n_137__15_,
  r_n_137__14_,r_n_137__13_,r_n_137__12_,r_n_137__11_,r_n_137__10_,r_n_137__9_,
  r_n_137__8_,r_n_137__7_,r_n_137__6_,r_n_137__5_,r_n_137__4_,r_n_137__3_,r_n_137__2_,
  r_n_137__1_,r_n_137__0_,r_n_136__31_,r_n_136__30_,r_n_136__29_,r_n_136__28_,
  r_n_136__27_,r_n_136__26_,r_n_136__25_,r_n_136__24_,r_n_136__23_,r_n_136__22_,r_n_136__21_,
  r_n_136__20_,r_n_136__19_,r_n_136__18_,r_n_136__17_,r_n_136__16_,r_n_136__15_,
  r_n_136__14_,r_n_136__13_,r_n_136__12_,r_n_136__11_,r_n_136__10_,r_n_136__9_,
  r_n_136__8_,r_n_136__7_,r_n_136__6_,r_n_136__5_,r_n_136__4_,r_n_136__3_,r_n_136__2_,
  r_n_136__1_,r_n_136__0_,r_n_135__31_,r_n_135__30_,r_n_135__29_,r_n_135__28_,
  r_n_135__27_,r_n_135__26_,r_n_135__25_,r_n_135__24_,r_n_135__23_,r_n_135__22_,
  r_n_135__21_,r_n_135__20_,r_n_135__19_,r_n_135__18_,r_n_135__17_,r_n_135__16_,
  r_n_135__15_,r_n_135__14_,r_n_135__13_,r_n_135__12_,r_n_135__11_,r_n_135__10_,
  r_n_135__9_,r_n_135__8_,r_n_135__7_,r_n_135__6_,r_n_135__5_,r_n_135__4_,r_n_135__3_,
  r_n_135__2_,r_n_135__1_,r_n_135__0_,r_n_134__31_,r_n_134__30_,r_n_134__29_,
  r_n_134__28_,r_n_134__27_,r_n_134__26_,r_n_134__25_,r_n_134__24_,r_n_134__23_,r_n_134__22_,
  r_n_134__21_,r_n_134__20_,r_n_134__19_,r_n_134__18_,r_n_134__17_,r_n_134__16_,
  r_n_134__15_,r_n_134__14_,r_n_134__13_,r_n_134__12_,r_n_134__11_,r_n_134__10_,
  r_n_134__9_,r_n_134__8_,r_n_134__7_,r_n_134__6_,r_n_134__5_,r_n_134__4_,r_n_134__3_,
  r_n_134__2_,r_n_134__1_,r_n_134__0_,r_n_133__31_,r_n_133__30_,r_n_133__29_,
  r_n_133__28_,r_n_133__27_,r_n_133__26_,r_n_133__25_,r_n_133__24_,r_n_133__23_,
  r_n_133__22_,r_n_133__21_,r_n_133__20_,r_n_133__19_,r_n_133__18_,r_n_133__17_,
  r_n_133__16_,r_n_133__15_,r_n_133__14_,r_n_133__13_,r_n_133__12_,r_n_133__11_,
  r_n_133__10_,r_n_133__9_,r_n_133__8_,r_n_133__7_,r_n_133__6_,r_n_133__5_,r_n_133__4_,
  r_n_133__3_,r_n_133__2_,r_n_133__1_,r_n_133__0_,r_n_132__31_,r_n_132__30_,r_n_132__29_,
  r_n_132__28_,r_n_132__27_,r_n_132__26_,r_n_132__25_,r_n_132__24_,r_n_132__23_,
  r_n_132__22_,r_n_132__21_,r_n_132__20_,r_n_132__19_,r_n_132__18_,r_n_132__17_,
  r_n_132__16_,r_n_132__15_,r_n_132__14_,r_n_132__13_,r_n_132__12_,r_n_132__11_,
  r_n_132__10_,r_n_132__9_,r_n_132__8_,r_n_132__7_,r_n_132__6_,r_n_132__5_,r_n_132__4_,
  r_n_132__3_,r_n_132__2_,r_n_132__1_,r_n_132__0_,r_n_131__31_,r_n_131__30_,
  r_n_131__29_,r_n_131__28_,r_n_131__27_,r_n_131__26_,r_n_131__25_,r_n_131__24_,
  r_n_131__23_,r_n_131__22_,r_n_131__21_,r_n_131__20_,r_n_131__19_,r_n_131__18_,
  r_n_131__17_,r_n_131__16_,r_n_131__15_,r_n_131__14_,r_n_131__13_,r_n_131__12_,r_n_131__11_,
  r_n_131__10_,r_n_131__9_,r_n_131__8_,r_n_131__7_,r_n_131__6_,r_n_131__5_,
  r_n_131__4_,r_n_131__3_,r_n_131__2_,r_n_131__1_,r_n_131__0_,r_n_130__31_,r_n_130__30_,
  r_n_130__29_,r_n_130__28_,r_n_130__27_,r_n_130__26_,r_n_130__25_,r_n_130__24_,
  r_n_130__23_,r_n_130__22_,r_n_130__21_,r_n_130__20_,r_n_130__19_,r_n_130__18_,
  r_n_130__17_,r_n_130__16_,r_n_130__15_,r_n_130__14_,r_n_130__13_,r_n_130__12_,
  r_n_130__11_,r_n_130__10_,r_n_130__9_,r_n_130__8_,r_n_130__7_,r_n_130__6_,r_n_130__5_,
  r_n_130__4_,r_n_130__3_,r_n_130__2_,r_n_130__1_,r_n_130__0_,r_n_129__31_,
  r_n_129__30_,r_n_129__29_,r_n_129__28_,r_n_129__27_,r_n_129__26_,r_n_129__25_,
  r_n_129__24_,r_n_129__23_,r_n_129__22_,r_n_129__21_,r_n_129__20_,r_n_129__19_,
  r_n_129__18_,r_n_129__17_,r_n_129__16_,r_n_129__15_,r_n_129__14_,r_n_129__13_,r_n_129__12_,
  r_n_129__11_,r_n_129__10_,r_n_129__9_,r_n_129__8_,r_n_129__7_,r_n_129__6_,
  r_n_129__5_,r_n_129__4_,r_n_129__3_,r_n_129__2_,r_n_129__1_,r_n_129__0_,r_n_160__31_,
  r_n_160__30_,r_n_160__29_,r_n_160__28_,r_n_160__27_,r_n_160__26_,r_n_160__25_,
  r_n_160__24_,r_n_160__23_,r_n_160__22_,r_n_160__21_,r_n_160__20_,r_n_160__19_,
  r_n_160__18_,r_n_160__17_,r_n_160__16_,r_n_160__15_,r_n_160__14_,r_n_160__13_,
  r_n_160__12_,r_n_160__11_,r_n_160__10_,r_n_160__9_,r_n_160__8_,r_n_160__7_,r_n_160__6_,
  r_n_160__5_,r_n_160__4_,r_n_160__3_,r_n_160__2_,r_n_160__1_,r_n_160__0_,
  r_n_159__31_,r_n_159__30_,r_n_159__29_,r_n_159__28_,r_n_159__27_,r_n_159__26_,
  r_n_159__25_,r_n_159__24_,r_n_159__23_,r_n_159__22_,r_n_159__21_,r_n_159__20_,r_n_159__19_,
  r_n_159__18_,r_n_159__17_,r_n_159__16_,r_n_159__15_,r_n_159__14_,r_n_159__13_,
  r_n_159__12_,r_n_159__11_,r_n_159__10_,r_n_159__9_,r_n_159__8_,r_n_159__7_,
  r_n_159__6_,r_n_159__5_,r_n_159__4_,r_n_159__3_,r_n_159__2_,r_n_159__1_,r_n_159__0_,
  r_n_158__31_,r_n_158__30_,r_n_158__29_,r_n_158__28_,r_n_158__27_,r_n_158__26_,
  r_n_158__25_,r_n_158__24_,r_n_158__23_,r_n_158__22_,r_n_158__21_,r_n_158__20_,
  r_n_158__19_,r_n_158__18_,r_n_158__17_,r_n_158__16_,r_n_158__15_,r_n_158__14_,
  r_n_158__13_,r_n_158__12_,r_n_158__11_,r_n_158__10_,r_n_158__9_,r_n_158__8_,r_n_158__7_,
  r_n_158__6_,r_n_158__5_,r_n_158__4_,r_n_158__3_,r_n_158__2_,r_n_158__1_,
  r_n_158__0_,r_n_157__31_,r_n_157__30_,r_n_157__29_,r_n_157__28_,r_n_157__27_,
  r_n_157__26_,r_n_157__25_,r_n_157__24_,r_n_157__23_,r_n_157__22_,r_n_157__21_,r_n_157__20_,
  r_n_157__19_,r_n_157__18_,r_n_157__17_,r_n_157__16_,r_n_157__15_,r_n_157__14_,
  r_n_157__13_,r_n_157__12_,r_n_157__11_,r_n_157__10_,r_n_157__9_,r_n_157__8_,
  r_n_157__7_,r_n_157__6_,r_n_157__5_,r_n_157__4_,r_n_157__3_,r_n_157__2_,r_n_157__1_,
  r_n_157__0_,r_n_156__31_,r_n_156__30_,r_n_156__29_,r_n_156__28_,r_n_156__27_,
  r_n_156__26_,r_n_156__25_,r_n_156__24_,r_n_156__23_,r_n_156__22_,r_n_156__21_,
  r_n_156__20_,r_n_156__19_,r_n_156__18_,r_n_156__17_,r_n_156__16_,r_n_156__15_,
  r_n_156__14_,r_n_156__13_,r_n_156__12_,r_n_156__11_,r_n_156__10_,r_n_156__9_,r_n_156__8_,
  r_n_156__7_,r_n_156__6_,r_n_156__5_,r_n_156__4_,r_n_156__3_,r_n_156__2_,
  r_n_156__1_,r_n_156__0_,r_n_155__31_,r_n_155__30_,r_n_155__29_,r_n_155__28_,r_n_155__27_,
  r_n_155__26_,r_n_155__25_,r_n_155__24_,r_n_155__23_,r_n_155__22_,r_n_155__21_,
  r_n_155__20_,r_n_155__19_,r_n_155__18_,r_n_155__17_,r_n_155__16_,r_n_155__15_,
  r_n_155__14_,r_n_155__13_,r_n_155__12_,r_n_155__11_,r_n_155__10_,r_n_155__9_,
  r_n_155__8_,r_n_155__7_,r_n_155__6_,r_n_155__5_,r_n_155__4_,r_n_155__3_,r_n_155__2_,
  r_n_155__1_,r_n_155__0_,r_n_154__31_,r_n_154__30_,r_n_154__29_,r_n_154__28_,
  r_n_154__27_,r_n_154__26_,r_n_154__25_,r_n_154__24_,r_n_154__23_,r_n_154__22_,
  r_n_154__21_,r_n_154__20_,r_n_154__19_,r_n_154__18_,r_n_154__17_,r_n_154__16_,
  r_n_154__15_,r_n_154__14_,r_n_154__13_,r_n_154__12_,r_n_154__11_,r_n_154__10_,r_n_154__9_,
  r_n_154__8_,r_n_154__7_,r_n_154__6_,r_n_154__5_,r_n_154__4_,r_n_154__3_,
  r_n_154__2_,r_n_154__1_,r_n_154__0_,r_n_153__31_,r_n_153__30_,r_n_153__29_,r_n_153__28_,
  r_n_153__27_,r_n_153__26_,r_n_153__25_,r_n_153__24_,r_n_153__23_,r_n_153__22_,
  r_n_153__21_,r_n_153__20_,r_n_153__19_,r_n_153__18_,r_n_153__17_,r_n_153__16_,
  r_n_153__15_,r_n_153__14_,r_n_153__13_,r_n_153__12_,r_n_153__11_,r_n_153__10_,
  r_n_153__9_,r_n_153__8_,r_n_153__7_,r_n_153__6_,r_n_153__5_,r_n_153__4_,r_n_153__3_,
  r_n_153__2_,r_n_153__1_,r_n_153__0_,r_n_152__31_,r_n_152__30_,r_n_152__29_,
  r_n_152__28_,r_n_152__27_,r_n_152__26_,r_n_152__25_,r_n_152__24_,r_n_152__23_,
  r_n_152__22_,r_n_152__21_,r_n_152__20_,r_n_152__19_,r_n_152__18_,r_n_152__17_,
  r_n_152__16_,r_n_152__15_,r_n_152__14_,r_n_152__13_,r_n_152__12_,r_n_152__11_,r_n_152__10_,
  r_n_152__9_,r_n_152__8_,r_n_152__7_,r_n_152__6_,r_n_152__5_,r_n_152__4_,
  r_n_152__3_,r_n_152__2_,r_n_152__1_,r_n_152__0_,r_n_151__31_,r_n_151__30_,r_n_151__29_,
  r_n_151__28_,r_n_151__27_,r_n_151__26_,r_n_151__25_,r_n_151__24_,r_n_151__23_,
  r_n_151__22_,r_n_151__21_,r_n_151__20_,r_n_151__19_,r_n_151__18_,r_n_151__17_,
  r_n_151__16_,r_n_151__15_,r_n_151__14_,r_n_151__13_,r_n_151__12_,r_n_151__11_,
  r_n_151__10_,r_n_151__9_,r_n_151__8_,r_n_151__7_,r_n_151__6_,r_n_151__5_,r_n_151__4_,
  r_n_151__3_,r_n_151__2_,r_n_151__1_,r_n_151__0_,r_n_150__31_,r_n_150__30_,
  r_n_150__29_,r_n_150__28_,r_n_150__27_,r_n_150__26_,r_n_150__25_,r_n_150__24_,
  r_n_150__23_,r_n_150__22_,r_n_150__21_,r_n_150__20_,r_n_150__19_,r_n_150__18_,r_n_150__17_,
  r_n_150__16_,r_n_150__15_,r_n_150__14_,r_n_150__13_,r_n_150__12_,r_n_150__11_,
  r_n_150__10_,r_n_150__9_,r_n_150__8_,r_n_150__7_,r_n_150__6_,r_n_150__5_,
  r_n_150__4_,r_n_150__3_,r_n_150__2_,r_n_150__1_,r_n_150__0_,r_n_149__31_,r_n_149__30_,
  r_n_149__29_,r_n_149__28_,r_n_149__27_,r_n_149__26_,r_n_149__25_,r_n_149__24_,
  r_n_149__23_,r_n_149__22_,r_n_149__21_,r_n_149__20_,r_n_149__19_,r_n_149__18_,
  r_n_149__17_,r_n_149__16_,r_n_149__15_,r_n_149__14_,r_n_149__13_,r_n_149__12_,
  r_n_149__11_,r_n_149__10_,r_n_149__9_,r_n_149__8_,r_n_149__7_,r_n_149__6_,r_n_149__5_,
  r_n_149__4_,r_n_149__3_,r_n_149__2_,r_n_149__1_,r_n_149__0_,r_n_148__31_,
  r_n_148__30_,r_n_148__29_,r_n_148__28_,r_n_148__27_,r_n_148__26_,r_n_148__25_,
  r_n_148__24_,r_n_148__23_,r_n_148__22_,r_n_148__21_,r_n_148__20_,r_n_148__19_,r_n_148__18_,
  r_n_148__17_,r_n_148__16_,r_n_148__15_,r_n_148__14_,r_n_148__13_,r_n_148__12_,
  r_n_148__11_,r_n_148__10_,r_n_148__9_,r_n_148__8_,r_n_148__7_,r_n_148__6_,
  r_n_148__5_,r_n_148__4_,r_n_148__3_,r_n_148__2_,r_n_148__1_,r_n_148__0_,r_n_147__31_,
  r_n_147__30_,r_n_147__29_,r_n_147__28_,r_n_147__27_,r_n_147__26_,r_n_147__25_,
  r_n_147__24_,r_n_147__23_,r_n_147__22_,r_n_147__21_,r_n_147__20_,r_n_147__19_,
  r_n_147__18_,r_n_147__17_,r_n_147__16_,r_n_147__15_,r_n_147__14_,r_n_147__13_,
  r_n_147__12_,r_n_147__11_,r_n_147__10_,r_n_147__9_,r_n_147__8_,r_n_147__7_,r_n_147__6_,
  r_n_147__5_,r_n_147__4_,r_n_147__3_,r_n_147__2_,r_n_147__1_,r_n_147__0_,
  r_n_146__31_,r_n_146__30_,r_n_146__29_,r_n_146__28_,r_n_146__27_,r_n_146__26_,r_n_146__25_,
  r_n_146__24_,r_n_146__23_,r_n_146__22_,r_n_146__21_,r_n_146__20_,r_n_146__19_,
  r_n_146__18_,r_n_146__17_,r_n_146__16_,r_n_146__15_,r_n_146__14_,r_n_146__13_,
  r_n_146__12_,r_n_146__11_,r_n_146__10_,r_n_146__9_,r_n_146__8_,r_n_146__7_,
  r_n_146__6_,r_n_146__5_,r_n_146__4_,r_n_146__3_,r_n_146__2_,r_n_146__1_,r_n_146__0_,
  r_n_145__31_,r_n_145__30_,r_n_145__29_,r_n_145__28_,r_n_145__27_,r_n_145__26_,
  r_n_145__25_,r_n_145__24_,r_n_145__23_,r_n_145__22_,r_n_145__21_,r_n_145__20_,
  r_n_145__19_,r_n_145__18_,r_n_145__17_,r_n_145__16_,r_n_145__15_,r_n_145__14_,
  r_n_145__13_,r_n_145__12_,r_n_145__11_,r_n_145__10_,r_n_145__9_,r_n_145__8_,r_n_145__7_,
  r_n_145__6_,r_n_145__5_,r_n_145__4_,r_n_145__3_,r_n_145__2_,r_n_145__1_,
  r_n_145__0_,r_n_176__31_,r_n_176__30_,r_n_176__29_,r_n_176__28_,r_n_176__27_,r_n_176__26_,
  r_n_176__25_,r_n_176__24_,r_n_176__23_,r_n_176__22_,r_n_176__21_,r_n_176__20_,
  r_n_176__19_,r_n_176__18_,r_n_176__17_,r_n_176__16_,r_n_176__15_,r_n_176__14_,
  r_n_176__13_,r_n_176__12_,r_n_176__11_,r_n_176__10_,r_n_176__9_,r_n_176__8_,
  r_n_176__7_,r_n_176__6_,r_n_176__5_,r_n_176__4_,r_n_176__3_,r_n_176__2_,r_n_176__1_,
  r_n_176__0_,r_n_175__31_,r_n_175__30_,r_n_175__29_,r_n_175__28_,r_n_175__27_,
  r_n_175__26_,r_n_175__25_,r_n_175__24_,r_n_175__23_,r_n_175__22_,r_n_175__21_,
  r_n_175__20_,r_n_175__19_,r_n_175__18_,r_n_175__17_,r_n_175__16_,r_n_175__15_,
  r_n_175__14_,r_n_175__13_,r_n_175__12_,r_n_175__11_,r_n_175__10_,r_n_175__9_,r_n_175__8_,
  r_n_175__7_,r_n_175__6_,r_n_175__5_,r_n_175__4_,r_n_175__3_,r_n_175__2_,
  r_n_175__1_,r_n_175__0_,r_n_174__31_,r_n_174__30_,r_n_174__29_,r_n_174__28_,r_n_174__27_,
  r_n_174__26_,r_n_174__25_,r_n_174__24_,r_n_174__23_,r_n_174__22_,r_n_174__21_,
  r_n_174__20_,r_n_174__19_,r_n_174__18_,r_n_174__17_,r_n_174__16_,r_n_174__15_,
  r_n_174__14_,r_n_174__13_,r_n_174__12_,r_n_174__11_,r_n_174__10_,r_n_174__9_,
  r_n_174__8_,r_n_174__7_,r_n_174__6_,r_n_174__5_,r_n_174__4_,r_n_174__3_,r_n_174__2_,
  r_n_174__1_,r_n_174__0_,r_n_173__31_,r_n_173__30_,r_n_173__29_,r_n_173__28_,
  r_n_173__27_,r_n_173__26_,r_n_173__25_,r_n_173__24_,r_n_173__23_,r_n_173__22_,
  r_n_173__21_,r_n_173__20_,r_n_173__19_,r_n_173__18_,r_n_173__17_,r_n_173__16_,r_n_173__15_,
  r_n_173__14_,r_n_173__13_,r_n_173__12_,r_n_173__11_,r_n_173__10_,r_n_173__9_,
  r_n_173__8_,r_n_173__7_,r_n_173__6_,r_n_173__5_,r_n_173__4_,r_n_173__3_,
  r_n_173__2_,r_n_173__1_,r_n_173__0_,r_n_172__31_,r_n_172__30_,r_n_172__29_,r_n_172__28_,
  r_n_172__27_,r_n_172__26_,r_n_172__25_,r_n_172__24_,r_n_172__23_,r_n_172__22_,
  r_n_172__21_,r_n_172__20_,r_n_172__19_,r_n_172__18_,r_n_172__17_,r_n_172__16_,
  r_n_172__15_,r_n_172__14_,r_n_172__13_,r_n_172__12_,r_n_172__11_,r_n_172__10_,
  r_n_172__9_,r_n_172__8_,r_n_172__7_,r_n_172__6_,r_n_172__5_,r_n_172__4_,r_n_172__3_,
  r_n_172__2_,r_n_172__1_,r_n_172__0_,r_n_171__31_,r_n_171__30_,r_n_171__29_,
  r_n_171__28_,r_n_171__27_,r_n_171__26_,r_n_171__25_,r_n_171__24_,r_n_171__23_,
  r_n_171__22_,r_n_171__21_,r_n_171__20_,r_n_171__19_,r_n_171__18_,r_n_171__17_,r_n_171__16_,
  r_n_171__15_,r_n_171__14_,r_n_171__13_,r_n_171__12_,r_n_171__11_,r_n_171__10_,
  r_n_171__9_,r_n_171__8_,r_n_171__7_,r_n_171__6_,r_n_171__5_,r_n_171__4_,
  r_n_171__3_,r_n_171__2_,r_n_171__1_,r_n_171__0_,r_n_170__31_,r_n_170__30_,r_n_170__29_,
  r_n_170__28_,r_n_170__27_,r_n_170__26_,r_n_170__25_,r_n_170__24_,r_n_170__23_,
  r_n_170__22_,r_n_170__21_,r_n_170__20_,r_n_170__19_,r_n_170__18_,r_n_170__17_,
  r_n_170__16_,r_n_170__15_,r_n_170__14_,r_n_170__13_,r_n_170__12_,r_n_170__11_,
  r_n_170__10_,r_n_170__9_,r_n_170__8_,r_n_170__7_,r_n_170__6_,r_n_170__5_,r_n_170__4_,
  r_n_170__3_,r_n_170__2_,r_n_170__1_,r_n_170__0_,r_n_169__31_,r_n_169__30_,
  r_n_169__29_,r_n_169__28_,r_n_169__27_,r_n_169__26_,r_n_169__25_,r_n_169__24_,r_n_169__23_,
  r_n_169__22_,r_n_169__21_,r_n_169__20_,r_n_169__19_,r_n_169__18_,r_n_169__17_,
  r_n_169__16_,r_n_169__15_,r_n_169__14_,r_n_169__13_,r_n_169__12_,r_n_169__11_,
  r_n_169__10_,r_n_169__9_,r_n_169__8_,r_n_169__7_,r_n_169__6_,r_n_169__5_,
  r_n_169__4_,r_n_169__3_,r_n_169__2_,r_n_169__1_,r_n_169__0_,r_n_168__31_,r_n_168__30_,
  r_n_168__29_,r_n_168__28_,r_n_168__27_,r_n_168__26_,r_n_168__25_,r_n_168__24_,
  r_n_168__23_,r_n_168__22_,r_n_168__21_,r_n_168__20_,r_n_168__19_,r_n_168__18_,
  r_n_168__17_,r_n_168__16_,r_n_168__15_,r_n_168__14_,r_n_168__13_,r_n_168__12_,
  r_n_168__11_,r_n_168__10_,r_n_168__9_,r_n_168__8_,r_n_168__7_,r_n_168__6_,r_n_168__5_,
  r_n_168__4_,r_n_168__3_,r_n_168__2_,r_n_168__1_,r_n_168__0_,r_n_167__31_,
  r_n_167__30_,r_n_167__29_,r_n_167__28_,r_n_167__27_,r_n_167__26_,r_n_167__25_,r_n_167__24_,
  r_n_167__23_,r_n_167__22_,r_n_167__21_,r_n_167__20_,r_n_167__19_,r_n_167__18_,
  r_n_167__17_,r_n_167__16_,r_n_167__15_,r_n_167__14_,r_n_167__13_,r_n_167__12_,
  r_n_167__11_,r_n_167__10_,r_n_167__9_,r_n_167__8_,r_n_167__7_,r_n_167__6_,
  r_n_167__5_,r_n_167__4_,r_n_167__3_,r_n_167__2_,r_n_167__1_,r_n_167__0_,r_n_166__31_,
  r_n_166__30_,r_n_166__29_,r_n_166__28_,r_n_166__27_,r_n_166__26_,r_n_166__25_,
  r_n_166__24_,r_n_166__23_,r_n_166__22_,r_n_166__21_,r_n_166__20_,r_n_166__19_,
  r_n_166__18_,r_n_166__17_,r_n_166__16_,r_n_166__15_,r_n_166__14_,r_n_166__13_,
  r_n_166__12_,r_n_166__11_,r_n_166__10_,r_n_166__9_,r_n_166__8_,r_n_166__7_,r_n_166__6_,
  r_n_166__5_,r_n_166__4_,r_n_166__3_,r_n_166__2_,r_n_166__1_,r_n_166__0_,r_n_165__31_,
  r_n_165__30_,r_n_165__29_,r_n_165__28_,r_n_165__27_,r_n_165__26_,r_n_165__25_,
  r_n_165__24_,r_n_165__23_,r_n_165__22_,r_n_165__21_,r_n_165__20_,r_n_165__19_,
  r_n_165__18_,r_n_165__17_,r_n_165__16_,r_n_165__15_,r_n_165__14_,r_n_165__13_,
  r_n_165__12_,r_n_165__11_,r_n_165__10_,r_n_165__9_,r_n_165__8_,r_n_165__7_,
  r_n_165__6_,r_n_165__5_,r_n_165__4_,r_n_165__3_,r_n_165__2_,r_n_165__1_,r_n_165__0_,
  r_n_164__31_,r_n_164__30_,r_n_164__29_,r_n_164__28_,r_n_164__27_,r_n_164__26_,
  r_n_164__25_,r_n_164__24_,r_n_164__23_,r_n_164__22_,r_n_164__21_,r_n_164__20_,
  r_n_164__19_,r_n_164__18_,r_n_164__17_,r_n_164__16_,r_n_164__15_,r_n_164__14_,r_n_164__13_,
  r_n_164__12_,r_n_164__11_,r_n_164__10_,r_n_164__9_,r_n_164__8_,r_n_164__7_,
  r_n_164__6_,r_n_164__5_,r_n_164__4_,r_n_164__3_,r_n_164__2_,r_n_164__1_,r_n_164__0_,
  r_n_163__31_,r_n_163__30_,r_n_163__29_,r_n_163__28_,r_n_163__27_,r_n_163__26_,
  r_n_163__25_,r_n_163__24_,r_n_163__23_,r_n_163__22_,r_n_163__21_,r_n_163__20_,
  r_n_163__19_,r_n_163__18_,r_n_163__17_,r_n_163__16_,r_n_163__15_,r_n_163__14_,
  r_n_163__13_,r_n_163__12_,r_n_163__11_,r_n_163__10_,r_n_163__9_,r_n_163__8_,
  r_n_163__7_,r_n_163__6_,r_n_163__5_,r_n_163__4_,r_n_163__3_,r_n_163__2_,r_n_163__1_,
  r_n_163__0_,r_n_162__31_,r_n_162__30_,r_n_162__29_,r_n_162__28_,r_n_162__27_,
  r_n_162__26_,r_n_162__25_,r_n_162__24_,r_n_162__23_,r_n_162__22_,r_n_162__21_,
  r_n_162__20_,r_n_162__19_,r_n_162__18_,r_n_162__17_,r_n_162__16_,r_n_162__15_,r_n_162__14_,
  r_n_162__13_,r_n_162__12_,r_n_162__11_,r_n_162__10_,r_n_162__9_,r_n_162__8_,
  r_n_162__7_,r_n_162__6_,r_n_162__5_,r_n_162__4_,r_n_162__3_,r_n_162__2_,r_n_162__1_,
  r_n_162__0_,r_n_161__31_,r_n_161__30_,r_n_161__29_,r_n_161__28_,r_n_161__27_,
  r_n_161__26_,r_n_161__25_,r_n_161__24_,r_n_161__23_,r_n_161__22_,r_n_161__21_,
  r_n_161__20_,r_n_161__19_,r_n_161__18_,r_n_161__17_,r_n_161__16_,r_n_161__15_,
  r_n_161__14_,r_n_161__13_,r_n_161__12_,r_n_161__11_,r_n_161__10_,r_n_161__9_,
  r_n_161__8_,r_n_161__7_,r_n_161__6_,r_n_161__5_,r_n_161__4_,r_n_161__3_,r_n_161__2_,
  r_n_161__1_,r_n_161__0_,r_n_192__31_,r_n_192__30_,r_n_192__29_,r_n_192__28_,
  r_n_192__27_,r_n_192__26_,r_n_192__25_,r_n_192__24_,r_n_192__23_,r_n_192__22_,r_n_192__21_,
  r_n_192__20_,r_n_192__19_,r_n_192__18_,r_n_192__17_,r_n_192__16_,r_n_192__15_,
  r_n_192__14_,r_n_192__13_,r_n_192__12_,r_n_192__11_,r_n_192__10_,r_n_192__9_,
  r_n_192__8_,r_n_192__7_,r_n_192__6_,r_n_192__5_,r_n_192__4_,r_n_192__3_,r_n_192__2_,
  r_n_192__1_,r_n_192__0_,r_n_191__31_,r_n_191__30_,r_n_191__29_,r_n_191__28_,
  r_n_191__27_,r_n_191__26_,r_n_191__25_,r_n_191__24_,r_n_191__23_,r_n_191__22_,
  r_n_191__21_,r_n_191__20_,r_n_191__19_,r_n_191__18_,r_n_191__17_,r_n_191__16_,
  r_n_191__15_,r_n_191__14_,r_n_191__13_,r_n_191__12_,r_n_191__11_,r_n_191__10_,
  r_n_191__9_,r_n_191__8_,r_n_191__7_,r_n_191__6_,r_n_191__5_,r_n_191__4_,r_n_191__3_,
  r_n_191__2_,r_n_191__1_,r_n_191__0_,r_n_190__31_,r_n_190__30_,r_n_190__29_,
  r_n_190__28_,r_n_190__27_,r_n_190__26_,r_n_190__25_,r_n_190__24_,r_n_190__23_,r_n_190__22_,
  r_n_190__21_,r_n_190__20_,r_n_190__19_,r_n_190__18_,r_n_190__17_,r_n_190__16_,
  r_n_190__15_,r_n_190__14_,r_n_190__13_,r_n_190__12_,r_n_190__11_,r_n_190__10_,
  r_n_190__9_,r_n_190__8_,r_n_190__7_,r_n_190__6_,r_n_190__5_,r_n_190__4_,r_n_190__3_,
  r_n_190__2_,r_n_190__1_,r_n_190__0_,r_n_189__31_,r_n_189__30_,r_n_189__29_,
  r_n_189__28_,r_n_189__27_,r_n_189__26_,r_n_189__25_,r_n_189__24_,r_n_189__23_,
  r_n_189__22_,r_n_189__21_,r_n_189__20_,r_n_189__19_,r_n_189__18_,r_n_189__17_,
  r_n_189__16_,r_n_189__15_,r_n_189__14_,r_n_189__13_,r_n_189__12_,r_n_189__11_,
  r_n_189__10_,r_n_189__9_,r_n_189__8_,r_n_189__7_,r_n_189__6_,r_n_189__5_,r_n_189__4_,
  r_n_189__3_,r_n_189__2_,r_n_189__1_,r_n_189__0_,r_n_188__31_,r_n_188__30_,r_n_188__29_,
  r_n_188__28_,r_n_188__27_,r_n_188__26_,r_n_188__25_,r_n_188__24_,r_n_188__23_,
  r_n_188__22_,r_n_188__21_,r_n_188__20_,r_n_188__19_,r_n_188__18_,r_n_188__17_,
  r_n_188__16_,r_n_188__15_,r_n_188__14_,r_n_188__13_,r_n_188__12_,r_n_188__11_,
  r_n_188__10_,r_n_188__9_,r_n_188__8_,r_n_188__7_,r_n_188__6_,r_n_188__5_,r_n_188__4_,
  r_n_188__3_,r_n_188__2_,r_n_188__1_,r_n_188__0_,r_n_187__31_,r_n_187__30_,
  r_n_187__29_,r_n_187__28_,r_n_187__27_,r_n_187__26_,r_n_187__25_,r_n_187__24_,
  r_n_187__23_,r_n_187__22_,r_n_187__21_,r_n_187__20_,r_n_187__19_,r_n_187__18_,
  r_n_187__17_,r_n_187__16_,r_n_187__15_,r_n_187__14_,r_n_187__13_,r_n_187__12_,r_n_187__11_,
  r_n_187__10_,r_n_187__9_,r_n_187__8_,r_n_187__7_,r_n_187__6_,r_n_187__5_,
  r_n_187__4_,r_n_187__3_,r_n_187__2_,r_n_187__1_,r_n_187__0_,r_n_186__31_,r_n_186__30_,
  r_n_186__29_,r_n_186__28_,r_n_186__27_,r_n_186__26_,r_n_186__25_,r_n_186__24_,
  r_n_186__23_,r_n_186__22_,r_n_186__21_,r_n_186__20_,r_n_186__19_,r_n_186__18_,
  r_n_186__17_,r_n_186__16_,r_n_186__15_,r_n_186__14_,r_n_186__13_,r_n_186__12_,
  r_n_186__11_,r_n_186__10_,r_n_186__9_,r_n_186__8_,r_n_186__7_,r_n_186__6_,r_n_186__5_,
  r_n_186__4_,r_n_186__3_,r_n_186__2_,r_n_186__1_,r_n_186__0_,r_n_185__31_,
  r_n_185__30_,r_n_185__29_,r_n_185__28_,r_n_185__27_,r_n_185__26_,r_n_185__25_,
  r_n_185__24_,r_n_185__23_,r_n_185__22_,r_n_185__21_,r_n_185__20_,r_n_185__19_,
  r_n_185__18_,r_n_185__17_,r_n_185__16_,r_n_185__15_,r_n_185__14_,r_n_185__13_,r_n_185__12_,
  r_n_185__11_,r_n_185__10_,r_n_185__9_,r_n_185__8_,r_n_185__7_,r_n_185__6_,
  r_n_185__5_,r_n_185__4_,r_n_185__3_,r_n_185__2_,r_n_185__1_,r_n_185__0_,r_n_184__31_,
  r_n_184__30_,r_n_184__29_,r_n_184__28_,r_n_184__27_,r_n_184__26_,r_n_184__25_,
  r_n_184__24_,r_n_184__23_,r_n_184__22_,r_n_184__21_,r_n_184__20_,r_n_184__19_,
  r_n_184__18_,r_n_184__17_,r_n_184__16_,r_n_184__15_,r_n_184__14_,r_n_184__13_,
  r_n_184__12_,r_n_184__11_,r_n_184__10_,r_n_184__9_,r_n_184__8_,r_n_184__7_,r_n_184__6_,
  r_n_184__5_,r_n_184__4_,r_n_184__3_,r_n_184__2_,r_n_184__1_,r_n_184__0_,
  r_n_183__31_,r_n_183__30_,r_n_183__29_,r_n_183__28_,r_n_183__27_,r_n_183__26_,
  r_n_183__25_,r_n_183__24_,r_n_183__23_,r_n_183__22_,r_n_183__21_,r_n_183__20_,r_n_183__19_,
  r_n_183__18_,r_n_183__17_,r_n_183__16_,r_n_183__15_,r_n_183__14_,r_n_183__13_,
  r_n_183__12_,r_n_183__11_,r_n_183__10_,r_n_183__9_,r_n_183__8_,r_n_183__7_,
  r_n_183__6_,r_n_183__5_,r_n_183__4_,r_n_183__3_,r_n_183__2_,r_n_183__1_,r_n_183__0_,
  r_n_182__31_,r_n_182__30_,r_n_182__29_,r_n_182__28_,r_n_182__27_,r_n_182__26_,
  r_n_182__25_,r_n_182__24_,r_n_182__23_,r_n_182__22_,r_n_182__21_,r_n_182__20_,
  r_n_182__19_,r_n_182__18_,r_n_182__17_,r_n_182__16_,r_n_182__15_,r_n_182__14_,
  r_n_182__13_,r_n_182__12_,r_n_182__11_,r_n_182__10_,r_n_182__9_,r_n_182__8_,r_n_182__7_,
  r_n_182__6_,r_n_182__5_,r_n_182__4_,r_n_182__3_,r_n_182__2_,r_n_182__1_,
  r_n_182__0_,r_n_181__31_,r_n_181__30_,r_n_181__29_,r_n_181__28_,r_n_181__27_,
  r_n_181__26_,r_n_181__25_,r_n_181__24_,r_n_181__23_,r_n_181__22_,r_n_181__21_,r_n_181__20_,
  r_n_181__19_,r_n_181__18_,r_n_181__17_,r_n_181__16_,r_n_181__15_,r_n_181__14_,
  r_n_181__13_,r_n_181__12_,r_n_181__11_,r_n_181__10_,r_n_181__9_,r_n_181__8_,
  r_n_181__7_,r_n_181__6_,r_n_181__5_,r_n_181__4_,r_n_181__3_,r_n_181__2_,r_n_181__1_,
  r_n_181__0_,r_n_180__31_,r_n_180__30_,r_n_180__29_,r_n_180__28_,r_n_180__27_,
  r_n_180__26_,r_n_180__25_,r_n_180__24_,r_n_180__23_,r_n_180__22_,r_n_180__21_,
  r_n_180__20_,r_n_180__19_,r_n_180__18_,r_n_180__17_,r_n_180__16_,r_n_180__15_,
  r_n_180__14_,r_n_180__13_,r_n_180__12_,r_n_180__11_,r_n_180__10_,r_n_180__9_,r_n_180__8_,
  r_n_180__7_,r_n_180__6_,r_n_180__5_,r_n_180__4_,r_n_180__3_,r_n_180__2_,
  r_n_180__1_,r_n_180__0_,r_n_179__31_,r_n_179__30_,r_n_179__29_,r_n_179__28_,r_n_179__27_,
  r_n_179__26_,r_n_179__25_,r_n_179__24_,r_n_179__23_,r_n_179__22_,r_n_179__21_,
  r_n_179__20_,r_n_179__19_,r_n_179__18_,r_n_179__17_,r_n_179__16_,r_n_179__15_,
  r_n_179__14_,r_n_179__13_,r_n_179__12_,r_n_179__11_,r_n_179__10_,r_n_179__9_,
  r_n_179__8_,r_n_179__7_,r_n_179__6_,r_n_179__5_,r_n_179__4_,r_n_179__3_,r_n_179__2_,
  r_n_179__1_,r_n_179__0_,r_n_178__31_,r_n_178__30_,r_n_178__29_,r_n_178__28_,
  r_n_178__27_,r_n_178__26_,r_n_178__25_,r_n_178__24_,r_n_178__23_,r_n_178__22_,
  r_n_178__21_,r_n_178__20_,r_n_178__19_,r_n_178__18_,r_n_178__17_,r_n_178__16_,
  r_n_178__15_,r_n_178__14_,r_n_178__13_,r_n_178__12_,r_n_178__11_,r_n_178__10_,r_n_178__9_,
  r_n_178__8_,r_n_178__7_,r_n_178__6_,r_n_178__5_,r_n_178__4_,r_n_178__3_,
  r_n_178__2_,r_n_178__1_,r_n_178__0_,r_n_177__31_,r_n_177__30_,r_n_177__29_,r_n_177__28_,
  r_n_177__27_,r_n_177__26_,r_n_177__25_,r_n_177__24_,r_n_177__23_,r_n_177__22_,
  r_n_177__21_,r_n_177__20_,r_n_177__19_,r_n_177__18_,r_n_177__17_,r_n_177__16_,
  r_n_177__15_,r_n_177__14_,r_n_177__13_,r_n_177__12_,r_n_177__11_,r_n_177__10_,
  r_n_177__9_,r_n_177__8_,r_n_177__7_,r_n_177__6_,r_n_177__5_,r_n_177__4_,r_n_177__3_,
  r_n_177__2_,r_n_177__1_,r_n_177__0_,r_n_208__31_,r_n_208__30_,r_n_208__29_,
  r_n_208__28_,r_n_208__27_,r_n_208__26_,r_n_208__25_,r_n_208__24_,r_n_208__23_,
  r_n_208__22_,r_n_208__21_,r_n_208__20_,r_n_208__19_,r_n_208__18_,r_n_208__17_,
  r_n_208__16_,r_n_208__15_,r_n_208__14_,r_n_208__13_,r_n_208__12_,r_n_208__11_,r_n_208__10_,
  r_n_208__9_,r_n_208__8_,r_n_208__7_,r_n_208__6_,r_n_208__5_,r_n_208__4_,
  r_n_208__3_,r_n_208__2_,r_n_208__1_,r_n_208__0_,r_n_207__31_,r_n_207__30_,r_n_207__29_,
  r_n_207__28_,r_n_207__27_,r_n_207__26_,r_n_207__25_,r_n_207__24_,r_n_207__23_,
  r_n_207__22_,r_n_207__21_,r_n_207__20_,r_n_207__19_,r_n_207__18_,r_n_207__17_,
  r_n_207__16_,r_n_207__15_,r_n_207__14_,r_n_207__13_,r_n_207__12_,r_n_207__11_,
  r_n_207__10_,r_n_207__9_,r_n_207__8_,r_n_207__7_,r_n_207__6_,r_n_207__5_,r_n_207__4_,
  r_n_207__3_,r_n_207__2_,r_n_207__1_,r_n_207__0_,r_n_206__31_,r_n_206__30_,
  r_n_206__29_,r_n_206__28_,r_n_206__27_,r_n_206__26_,r_n_206__25_,r_n_206__24_,
  r_n_206__23_,r_n_206__22_,r_n_206__21_,r_n_206__20_,r_n_206__19_,r_n_206__18_,r_n_206__17_,
  r_n_206__16_,r_n_206__15_,r_n_206__14_,r_n_206__13_,r_n_206__12_,r_n_206__11_,
  r_n_206__10_,r_n_206__9_,r_n_206__8_,r_n_206__7_,r_n_206__6_,r_n_206__5_,
  r_n_206__4_,r_n_206__3_,r_n_206__2_,r_n_206__1_,r_n_206__0_,r_n_205__31_,r_n_205__30_,
  r_n_205__29_,r_n_205__28_,r_n_205__27_,r_n_205__26_,r_n_205__25_,r_n_205__24_,
  r_n_205__23_,r_n_205__22_,r_n_205__21_,r_n_205__20_,r_n_205__19_,r_n_205__18_,
  r_n_205__17_,r_n_205__16_,r_n_205__15_,r_n_205__14_,r_n_205__13_,r_n_205__12_,
  r_n_205__11_,r_n_205__10_,r_n_205__9_,r_n_205__8_,r_n_205__7_,r_n_205__6_,r_n_205__5_,
  r_n_205__4_,r_n_205__3_,r_n_205__2_,r_n_205__1_,r_n_205__0_,r_n_204__31_,
  r_n_204__30_,r_n_204__29_,r_n_204__28_,r_n_204__27_,r_n_204__26_,r_n_204__25_,
  r_n_204__24_,r_n_204__23_,r_n_204__22_,r_n_204__21_,r_n_204__20_,r_n_204__19_,r_n_204__18_,
  r_n_204__17_,r_n_204__16_,r_n_204__15_,r_n_204__14_,r_n_204__13_,r_n_204__12_,
  r_n_204__11_,r_n_204__10_,r_n_204__9_,r_n_204__8_,r_n_204__7_,r_n_204__6_,
  r_n_204__5_,r_n_204__4_,r_n_204__3_,r_n_204__2_,r_n_204__1_,r_n_204__0_,r_n_203__31_,
  r_n_203__30_,r_n_203__29_,r_n_203__28_,r_n_203__27_,r_n_203__26_,r_n_203__25_,
  r_n_203__24_,r_n_203__23_,r_n_203__22_,r_n_203__21_,r_n_203__20_,r_n_203__19_,
  r_n_203__18_,r_n_203__17_,r_n_203__16_,r_n_203__15_,r_n_203__14_,r_n_203__13_,
  r_n_203__12_,r_n_203__11_,r_n_203__10_,r_n_203__9_,r_n_203__8_,r_n_203__7_,r_n_203__6_,
  r_n_203__5_,r_n_203__4_,r_n_203__3_,r_n_203__2_,r_n_203__1_,r_n_203__0_,
  r_n_202__31_,r_n_202__30_,r_n_202__29_,r_n_202__28_,r_n_202__27_,r_n_202__26_,r_n_202__25_,
  r_n_202__24_,r_n_202__23_,r_n_202__22_,r_n_202__21_,r_n_202__20_,r_n_202__19_,
  r_n_202__18_,r_n_202__17_,r_n_202__16_,r_n_202__15_,r_n_202__14_,r_n_202__13_,
  r_n_202__12_,r_n_202__11_,r_n_202__10_,r_n_202__9_,r_n_202__8_,r_n_202__7_,
  r_n_202__6_,r_n_202__5_,r_n_202__4_,r_n_202__3_,r_n_202__2_,r_n_202__1_,r_n_202__0_,
  r_n_201__31_,r_n_201__30_,r_n_201__29_,r_n_201__28_,r_n_201__27_,r_n_201__26_,
  r_n_201__25_,r_n_201__24_,r_n_201__23_,r_n_201__22_,r_n_201__21_,r_n_201__20_,
  r_n_201__19_,r_n_201__18_,r_n_201__17_,r_n_201__16_,r_n_201__15_,r_n_201__14_,
  r_n_201__13_,r_n_201__12_,r_n_201__11_,r_n_201__10_,r_n_201__9_,r_n_201__8_,r_n_201__7_,
  r_n_201__6_,r_n_201__5_,r_n_201__4_,r_n_201__3_,r_n_201__2_,r_n_201__1_,
  r_n_201__0_,r_n_200__31_,r_n_200__30_,r_n_200__29_,r_n_200__28_,r_n_200__27_,r_n_200__26_,
  r_n_200__25_,r_n_200__24_,r_n_200__23_,r_n_200__22_,r_n_200__21_,r_n_200__20_,
  r_n_200__19_,r_n_200__18_,r_n_200__17_,r_n_200__16_,r_n_200__15_,r_n_200__14_,
  r_n_200__13_,r_n_200__12_,r_n_200__11_,r_n_200__10_,r_n_200__9_,r_n_200__8_,
  r_n_200__7_,r_n_200__6_,r_n_200__5_,r_n_200__4_,r_n_200__3_,r_n_200__2_,r_n_200__1_,
  r_n_200__0_,r_n_199__31_,r_n_199__30_,r_n_199__29_,r_n_199__28_,r_n_199__27_,
  r_n_199__26_,r_n_199__25_,r_n_199__24_,r_n_199__23_,r_n_199__22_,r_n_199__21_,
  r_n_199__20_,r_n_199__19_,r_n_199__18_,r_n_199__17_,r_n_199__16_,r_n_199__15_,
  r_n_199__14_,r_n_199__13_,r_n_199__12_,r_n_199__11_,r_n_199__10_,r_n_199__9_,r_n_199__8_,
  r_n_199__7_,r_n_199__6_,r_n_199__5_,r_n_199__4_,r_n_199__3_,r_n_199__2_,
  r_n_199__1_,r_n_199__0_,r_n_198__31_,r_n_198__30_,r_n_198__29_,r_n_198__28_,r_n_198__27_,
  r_n_198__26_,r_n_198__25_,r_n_198__24_,r_n_198__23_,r_n_198__22_,r_n_198__21_,
  r_n_198__20_,r_n_198__19_,r_n_198__18_,r_n_198__17_,r_n_198__16_,r_n_198__15_,
  r_n_198__14_,r_n_198__13_,r_n_198__12_,r_n_198__11_,r_n_198__10_,r_n_198__9_,
  r_n_198__8_,r_n_198__7_,r_n_198__6_,r_n_198__5_,r_n_198__4_,r_n_198__3_,r_n_198__2_,
  r_n_198__1_,r_n_198__0_,r_n_197__31_,r_n_197__30_,r_n_197__29_,r_n_197__28_,
  r_n_197__27_,r_n_197__26_,r_n_197__25_,r_n_197__24_,r_n_197__23_,r_n_197__22_,
  r_n_197__21_,r_n_197__20_,r_n_197__19_,r_n_197__18_,r_n_197__17_,r_n_197__16_,r_n_197__15_,
  r_n_197__14_,r_n_197__13_,r_n_197__12_,r_n_197__11_,r_n_197__10_,r_n_197__9_,
  r_n_197__8_,r_n_197__7_,r_n_197__6_,r_n_197__5_,r_n_197__4_,r_n_197__3_,
  r_n_197__2_,r_n_197__1_,r_n_197__0_,r_n_196__31_,r_n_196__30_,r_n_196__29_,r_n_196__28_,
  r_n_196__27_,r_n_196__26_,r_n_196__25_,r_n_196__24_,r_n_196__23_,r_n_196__22_,
  r_n_196__21_,r_n_196__20_,r_n_196__19_,r_n_196__18_,r_n_196__17_,r_n_196__16_,
  r_n_196__15_,r_n_196__14_,r_n_196__13_,r_n_196__12_,r_n_196__11_,r_n_196__10_,
  r_n_196__9_,r_n_196__8_,r_n_196__7_,r_n_196__6_,r_n_196__5_,r_n_196__4_,r_n_196__3_,
  r_n_196__2_,r_n_196__1_,r_n_196__0_,r_n_195__31_,r_n_195__30_,r_n_195__29_,
  r_n_195__28_,r_n_195__27_,r_n_195__26_,r_n_195__25_,r_n_195__24_,r_n_195__23_,
  r_n_195__22_,r_n_195__21_,r_n_195__20_,r_n_195__19_,r_n_195__18_,r_n_195__17_,r_n_195__16_,
  r_n_195__15_,r_n_195__14_,r_n_195__13_,r_n_195__12_,r_n_195__11_,r_n_195__10_,
  r_n_195__9_,r_n_195__8_,r_n_195__7_,r_n_195__6_,r_n_195__5_,r_n_195__4_,
  r_n_195__3_,r_n_195__2_,r_n_195__1_,r_n_195__0_,r_n_194__31_,r_n_194__30_,r_n_194__29_,
  r_n_194__28_,r_n_194__27_,r_n_194__26_,r_n_194__25_,r_n_194__24_,r_n_194__23_,
  r_n_194__22_,r_n_194__21_,r_n_194__20_,r_n_194__19_,r_n_194__18_,r_n_194__17_,
  r_n_194__16_,r_n_194__15_,r_n_194__14_,r_n_194__13_,r_n_194__12_,r_n_194__11_,
  r_n_194__10_,r_n_194__9_,r_n_194__8_,r_n_194__7_,r_n_194__6_,r_n_194__5_,r_n_194__4_,
  r_n_194__3_,r_n_194__2_,r_n_194__1_,r_n_194__0_,r_n_193__31_,r_n_193__30_,
  r_n_193__29_,r_n_193__28_,r_n_193__27_,r_n_193__26_,r_n_193__25_,r_n_193__24_,r_n_193__23_,
  r_n_193__22_,r_n_193__21_,r_n_193__20_,r_n_193__19_,r_n_193__18_,r_n_193__17_,
  r_n_193__16_,r_n_193__15_,r_n_193__14_,r_n_193__13_,r_n_193__12_,r_n_193__11_,
  r_n_193__10_,r_n_193__9_,r_n_193__8_,r_n_193__7_,r_n_193__6_,r_n_193__5_,
  r_n_193__4_,r_n_193__3_,r_n_193__2_,r_n_193__1_,r_n_193__0_,r_n_224__31_,r_n_224__30_,
  r_n_224__29_,r_n_224__28_,r_n_224__27_,r_n_224__26_,r_n_224__25_,r_n_224__24_,
  r_n_224__23_,r_n_224__22_,r_n_224__21_,r_n_224__20_,r_n_224__19_,r_n_224__18_,
  r_n_224__17_,r_n_224__16_,r_n_224__15_,r_n_224__14_,r_n_224__13_,r_n_224__12_,
  r_n_224__11_,r_n_224__10_,r_n_224__9_,r_n_224__8_,r_n_224__7_,r_n_224__6_,r_n_224__5_,
  r_n_224__4_,r_n_224__3_,r_n_224__2_,r_n_224__1_,r_n_224__0_,r_n_223__31_,
  r_n_223__30_,r_n_223__29_,r_n_223__28_,r_n_223__27_,r_n_223__26_,r_n_223__25_,r_n_223__24_,
  r_n_223__23_,r_n_223__22_,r_n_223__21_,r_n_223__20_,r_n_223__19_,r_n_223__18_,
  r_n_223__17_,r_n_223__16_,r_n_223__15_,r_n_223__14_,r_n_223__13_,r_n_223__12_,
  r_n_223__11_,r_n_223__10_,r_n_223__9_,r_n_223__8_,r_n_223__7_,r_n_223__6_,
  r_n_223__5_,r_n_223__4_,r_n_223__3_,r_n_223__2_,r_n_223__1_,r_n_223__0_,r_n_222__31_,
  r_n_222__30_,r_n_222__29_,r_n_222__28_,r_n_222__27_,r_n_222__26_,r_n_222__25_,
  r_n_222__24_,r_n_222__23_,r_n_222__22_,r_n_222__21_,r_n_222__20_,r_n_222__19_,
  r_n_222__18_,r_n_222__17_,r_n_222__16_,r_n_222__15_,r_n_222__14_,r_n_222__13_,
  r_n_222__12_,r_n_222__11_,r_n_222__10_,r_n_222__9_,r_n_222__8_,r_n_222__7_,r_n_222__6_,
  r_n_222__5_,r_n_222__4_,r_n_222__3_,r_n_222__2_,r_n_222__1_,r_n_222__0_,r_n_221__31_,
  r_n_221__30_,r_n_221__29_,r_n_221__28_,r_n_221__27_,r_n_221__26_,r_n_221__25_,
  r_n_221__24_,r_n_221__23_,r_n_221__22_,r_n_221__21_,r_n_221__20_,r_n_221__19_,
  r_n_221__18_,r_n_221__17_,r_n_221__16_,r_n_221__15_,r_n_221__14_,r_n_221__13_,
  r_n_221__12_,r_n_221__11_,r_n_221__10_,r_n_221__9_,r_n_221__8_,r_n_221__7_,
  r_n_221__6_,r_n_221__5_,r_n_221__4_,r_n_221__3_,r_n_221__2_,r_n_221__1_,r_n_221__0_,
  r_n_220__31_,r_n_220__30_,r_n_220__29_,r_n_220__28_,r_n_220__27_,r_n_220__26_,
  r_n_220__25_,r_n_220__24_,r_n_220__23_,r_n_220__22_,r_n_220__21_,r_n_220__20_,
  r_n_220__19_,r_n_220__18_,r_n_220__17_,r_n_220__16_,r_n_220__15_,r_n_220__14_,r_n_220__13_,
  r_n_220__12_,r_n_220__11_,r_n_220__10_,r_n_220__9_,r_n_220__8_,r_n_220__7_,
  r_n_220__6_,r_n_220__5_,r_n_220__4_,r_n_220__3_,r_n_220__2_,r_n_220__1_,r_n_220__0_,
  r_n_219__31_,r_n_219__30_,r_n_219__29_,r_n_219__28_,r_n_219__27_,r_n_219__26_,
  r_n_219__25_,r_n_219__24_,r_n_219__23_,r_n_219__22_,r_n_219__21_,r_n_219__20_,
  r_n_219__19_,r_n_219__18_,r_n_219__17_,r_n_219__16_,r_n_219__15_,r_n_219__14_,
  r_n_219__13_,r_n_219__12_,r_n_219__11_,r_n_219__10_,r_n_219__9_,r_n_219__8_,
  r_n_219__7_,r_n_219__6_,r_n_219__5_,r_n_219__4_,r_n_219__3_,r_n_219__2_,r_n_219__1_,
  r_n_219__0_,r_n_218__31_,r_n_218__30_,r_n_218__29_,r_n_218__28_,r_n_218__27_,
  r_n_218__26_,r_n_218__25_,r_n_218__24_,r_n_218__23_,r_n_218__22_,r_n_218__21_,
  r_n_218__20_,r_n_218__19_,r_n_218__18_,r_n_218__17_,r_n_218__16_,r_n_218__15_,r_n_218__14_,
  r_n_218__13_,r_n_218__12_,r_n_218__11_,r_n_218__10_,r_n_218__9_,r_n_218__8_,
  r_n_218__7_,r_n_218__6_,r_n_218__5_,r_n_218__4_,r_n_218__3_,r_n_218__2_,r_n_218__1_,
  r_n_218__0_,r_n_217__31_,r_n_217__30_,r_n_217__29_,r_n_217__28_,r_n_217__27_,
  r_n_217__26_,r_n_217__25_,r_n_217__24_,r_n_217__23_,r_n_217__22_,r_n_217__21_,
  r_n_217__20_,r_n_217__19_,r_n_217__18_,r_n_217__17_,r_n_217__16_,r_n_217__15_,
  r_n_217__14_,r_n_217__13_,r_n_217__12_,r_n_217__11_,r_n_217__10_,r_n_217__9_,
  r_n_217__8_,r_n_217__7_,r_n_217__6_,r_n_217__5_,r_n_217__4_,r_n_217__3_,r_n_217__2_,
  r_n_217__1_,r_n_217__0_,r_n_216__31_,r_n_216__30_,r_n_216__29_,r_n_216__28_,
  r_n_216__27_,r_n_216__26_,r_n_216__25_,r_n_216__24_,r_n_216__23_,r_n_216__22_,r_n_216__21_,
  r_n_216__20_,r_n_216__19_,r_n_216__18_,r_n_216__17_,r_n_216__16_,r_n_216__15_,
  r_n_216__14_,r_n_216__13_,r_n_216__12_,r_n_216__11_,r_n_216__10_,r_n_216__9_,
  r_n_216__8_,r_n_216__7_,r_n_216__6_,r_n_216__5_,r_n_216__4_,r_n_216__3_,r_n_216__2_,
  r_n_216__1_,r_n_216__0_,r_n_215__31_,r_n_215__30_,r_n_215__29_,r_n_215__28_,
  r_n_215__27_,r_n_215__26_,r_n_215__25_,r_n_215__24_,r_n_215__23_,r_n_215__22_,
  r_n_215__21_,r_n_215__20_,r_n_215__19_,r_n_215__18_,r_n_215__17_,r_n_215__16_,
  r_n_215__15_,r_n_215__14_,r_n_215__13_,r_n_215__12_,r_n_215__11_,r_n_215__10_,
  r_n_215__9_,r_n_215__8_,r_n_215__7_,r_n_215__6_,r_n_215__5_,r_n_215__4_,r_n_215__3_,
  r_n_215__2_,r_n_215__1_,r_n_215__0_,r_n_214__31_,r_n_214__30_,r_n_214__29_,
  r_n_214__28_,r_n_214__27_,r_n_214__26_,r_n_214__25_,r_n_214__24_,r_n_214__23_,r_n_214__22_,
  r_n_214__21_,r_n_214__20_,r_n_214__19_,r_n_214__18_,r_n_214__17_,r_n_214__16_,
  r_n_214__15_,r_n_214__14_,r_n_214__13_,r_n_214__12_,r_n_214__11_,r_n_214__10_,
  r_n_214__9_,r_n_214__8_,r_n_214__7_,r_n_214__6_,r_n_214__5_,r_n_214__4_,r_n_214__3_,
  r_n_214__2_,r_n_214__1_,r_n_214__0_,r_n_213__31_,r_n_213__30_,r_n_213__29_,
  r_n_213__28_,r_n_213__27_,r_n_213__26_,r_n_213__25_,r_n_213__24_,r_n_213__23_,
  r_n_213__22_,r_n_213__21_,r_n_213__20_,r_n_213__19_,r_n_213__18_,r_n_213__17_,
  r_n_213__16_,r_n_213__15_,r_n_213__14_,r_n_213__13_,r_n_213__12_,r_n_213__11_,
  r_n_213__10_,r_n_213__9_,r_n_213__8_,r_n_213__7_,r_n_213__6_,r_n_213__5_,r_n_213__4_,
  r_n_213__3_,r_n_213__2_,r_n_213__1_,r_n_213__0_,r_n_212__31_,r_n_212__30_,r_n_212__29_,
  r_n_212__28_,r_n_212__27_,r_n_212__26_,r_n_212__25_,r_n_212__24_,r_n_212__23_,
  r_n_212__22_,r_n_212__21_,r_n_212__20_,r_n_212__19_,r_n_212__18_,r_n_212__17_,
  r_n_212__16_,r_n_212__15_,r_n_212__14_,r_n_212__13_,r_n_212__12_,r_n_212__11_,
  r_n_212__10_,r_n_212__9_,r_n_212__8_,r_n_212__7_,r_n_212__6_,r_n_212__5_,r_n_212__4_,
  r_n_212__3_,r_n_212__2_,r_n_212__1_,r_n_212__0_,r_n_211__31_,r_n_211__30_,
  r_n_211__29_,r_n_211__28_,r_n_211__27_,r_n_211__26_,r_n_211__25_,r_n_211__24_,
  r_n_211__23_,r_n_211__22_,r_n_211__21_,r_n_211__20_,r_n_211__19_,r_n_211__18_,
  r_n_211__17_,r_n_211__16_,r_n_211__15_,r_n_211__14_,r_n_211__13_,r_n_211__12_,r_n_211__11_,
  r_n_211__10_,r_n_211__9_,r_n_211__8_,r_n_211__7_,r_n_211__6_,r_n_211__5_,
  r_n_211__4_,r_n_211__3_,r_n_211__2_,r_n_211__1_,r_n_211__0_,r_n_210__31_,r_n_210__30_,
  r_n_210__29_,r_n_210__28_,r_n_210__27_,r_n_210__26_,r_n_210__25_,r_n_210__24_,
  r_n_210__23_,r_n_210__22_,r_n_210__21_,r_n_210__20_,r_n_210__19_,r_n_210__18_,
  r_n_210__17_,r_n_210__16_,r_n_210__15_,r_n_210__14_,r_n_210__13_,r_n_210__12_,
  r_n_210__11_,r_n_210__10_,r_n_210__9_,r_n_210__8_,r_n_210__7_,r_n_210__6_,r_n_210__5_,
  r_n_210__4_,r_n_210__3_,r_n_210__2_,r_n_210__1_,r_n_210__0_,r_n_209__31_,
  r_n_209__30_,r_n_209__29_,r_n_209__28_,r_n_209__27_,r_n_209__26_,r_n_209__25_,
  r_n_209__24_,r_n_209__23_,r_n_209__22_,r_n_209__21_,r_n_209__20_,r_n_209__19_,
  r_n_209__18_,r_n_209__17_,r_n_209__16_,r_n_209__15_,r_n_209__14_,r_n_209__13_,r_n_209__12_,
  r_n_209__11_,r_n_209__10_,r_n_209__9_,r_n_209__8_,r_n_209__7_,r_n_209__6_,
  r_n_209__5_,r_n_209__4_,r_n_209__3_,r_n_209__2_,r_n_209__1_,r_n_209__0_,r_n_240__31_,
  r_n_240__30_,r_n_240__29_,r_n_240__28_,r_n_240__27_,r_n_240__26_,r_n_240__25_,
  r_n_240__24_,r_n_240__23_,r_n_240__22_,r_n_240__21_,r_n_240__20_,r_n_240__19_,
  r_n_240__18_,r_n_240__17_,r_n_240__16_,r_n_240__15_,r_n_240__14_,r_n_240__13_,
  r_n_240__12_,r_n_240__11_,r_n_240__10_,r_n_240__9_,r_n_240__8_,r_n_240__7_,r_n_240__6_,
  r_n_240__5_,r_n_240__4_,r_n_240__3_,r_n_240__2_,r_n_240__1_,r_n_240__0_,
  r_n_239__31_,r_n_239__30_,r_n_239__29_,r_n_239__28_,r_n_239__27_,r_n_239__26_,
  r_n_239__25_,r_n_239__24_,r_n_239__23_,r_n_239__22_,r_n_239__21_,r_n_239__20_,r_n_239__19_,
  r_n_239__18_,r_n_239__17_,r_n_239__16_,r_n_239__15_,r_n_239__14_,r_n_239__13_,
  r_n_239__12_,r_n_239__11_,r_n_239__10_,r_n_239__9_,r_n_239__8_,r_n_239__7_,
  r_n_239__6_,r_n_239__5_,r_n_239__4_,r_n_239__3_,r_n_239__2_,r_n_239__1_,r_n_239__0_,
  r_n_238__31_,r_n_238__30_,r_n_238__29_,r_n_238__28_,r_n_238__27_,r_n_238__26_,
  r_n_238__25_,r_n_238__24_,r_n_238__23_,r_n_238__22_,r_n_238__21_,r_n_238__20_,
  r_n_238__19_,r_n_238__18_,r_n_238__17_,r_n_238__16_,r_n_238__15_,r_n_238__14_,
  r_n_238__13_,r_n_238__12_,r_n_238__11_,r_n_238__10_,r_n_238__9_,r_n_238__8_,r_n_238__7_,
  r_n_238__6_,r_n_238__5_,r_n_238__4_,r_n_238__3_,r_n_238__2_,r_n_238__1_,
  r_n_238__0_,r_n_237__31_,r_n_237__30_,r_n_237__29_,r_n_237__28_,r_n_237__27_,
  r_n_237__26_,r_n_237__25_,r_n_237__24_,r_n_237__23_,r_n_237__22_,r_n_237__21_,r_n_237__20_,
  r_n_237__19_,r_n_237__18_,r_n_237__17_,r_n_237__16_,r_n_237__15_,r_n_237__14_,
  r_n_237__13_,r_n_237__12_,r_n_237__11_,r_n_237__10_,r_n_237__9_,r_n_237__8_,
  r_n_237__7_,r_n_237__6_,r_n_237__5_,r_n_237__4_,r_n_237__3_,r_n_237__2_,r_n_237__1_,
  r_n_237__0_,r_n_236__31_,r_n_236__30_,r_n_236__29_,r_n_236__28_,r_n_236__27_,
  r_n_236__26_,r_n_236__25_,r_n_236__24_,r_n_236__23_,r_n_236__22_,r_n_236__21_,
  r_n_236__20_,r_n_236__19_,r_n_236__18_,r_n_236__17_,r_n_236__16_,r_n_236__15_,
  r_n_236__14_,r_n_236__13_,r_n_236__12_,r_n_236__11_,r_n_236__10_,r_n_236__9_,r_n_236__8_,
  r_n_236__7_,r_n_236__6_,r_n_236__5_,r_n_236__4_,r_n_236__3_,r_n_236__2_,
  r_n_236__1_,r_n_236__0_,r_n_235__31_,r_n_235__30_,r_n_235__29_,r_n_235__28_,r_n_235__27_,
  r_n_235__26_,r_n_235__25_,r_n_235__24_,r_n_235__23_,r_n_235__22_,r_n_235__21_,
  r_n_235__20_,r_n_235__19_,r_n_235__18_,r_n_235__17_,r_n_235__16_,r_n_235__15_,
  r_n_235__14_,r_n_235__13_,r_n_235__12_,r_n_235__11_,r_n_235__10_,r_n_235__9_,
  r_n_235__8_,r_n_235__7_,r_n_235__6_,r_n_235__5_,r_n_235__4_,r_n_235__3_,r_n_235__2_,
  r_n_235__1_,r_n_235__0_,r_n_234__31_,r_n_234__30_,r_n_234__29_,r_n_234__28_,
  r_n_234__27_,r_n_234__26_,r_n_234__25_,r_n_234__24_,r_n_234__23_,r_n_234__22_,
  r_n_234__21_,r_n_234__20_,r_n_234__19_,r_n_234__18_,r_n_234__17_,r_n_234__16_,
  r_n_234__15_,r_n_234__14_,r_n_234__13_,r_n_234__12_,r_n_234__11_,r_n_234__10_,r_n_234__9_,
  r_n_234__8_,r_n_234__7_,r_n_234__6_,r_n_234__5_,r_n_234__4_,r_n_234__3_,
  r_n_234__2_,r_n_234__1_,r_n_234__0_,r_n_233__31_,r_n_233__30_,r_n_233__29_,r_n_233__28_,
  r_n_233__27_,r_n_233__26_,r_n_233__25_,r_n_233__24_,r_n_233__23_,r_n_233__22_,
  r_n_233__21_,r_n_233__20_,r_n_233__19_,r_n_233__18_,r_n_233__17_,r_n_233__16_,
  r_n_233__15_,r_n_233__14_,r_n_233__13_,r_n_233__12_,r_n_233__11_,r_n_233__10_,
  r_n_233__9_,r_n_233__8_,r_n_233__7_,r_n_233__6_,r_n_233__5_,r_n_233__4_,r_n_233__3_,
  r_n_233__2_,r_n_233__1_,r_n_233__0_,r_n_232__31_,r_n_232__30_,r_n_232__29_,
  r_n_232__28_,r_n_232__27_,r_n_232__26_,r_n_232__25_,r_n_232__24_,r_n_232__23_,
  r_n_232__22_,r_n_232__21_,r_n_232__20_,r_n_232__19_,r_n_232__18_,r_n_232__17_,
  r_n_232__16_,r_n_232__15_,r_n_232__14_,r_n_232__13_,r_n_232__12_,r_n_232__11_,r_n_232__10_,
  r_n_232__9_,r_n_232__8_,r_n_232__7_,r_n_232__6_,r_n_232__5_,r_n_232__4_,
  r_n_232__3_,r_n_232__2_,r_n_232__1_,r_n_232__0_,r_n_231__31_,r_n_231__30_,r_n_231__29_,
  r_n_231__28_,r_n_231__27_,r_n_231__26_,r_n_231__25_,r_n_231__24_,r_n_231__23_,
  r_n_231__22_,r_n_231__21_,r_n_231__20_,r_n_231__19_,r_n_231__18_,r_n_231__17_,
  r_n_231__16_,r_n_231__15_,r_n_231__14_,r_n_231__13_,r_n_231__12_,r_n_231__11_,
  r_n_231__10_,r_n_231__9_,r_n_231__8_,r_n_231__7_,r_n_231__6_,r_n_231__5_,r_n_231__4_,
  r_n_231__3_,r_n_231__2_,r_n_231__1_,r_n_231__0_,r_n_230__31_,r_n_230__30_,
  r_n_230__29_,r_n_230__28_,r_n_230__27_,r_n_230__26_,r_n_230__25_,r_n_230__24_,
  r_n_230__23_,r_n_230__22_,r_n_230__21_,r_n_230__20_,r_n_230__19_,r_n_230__18_,r_n_230__17_,
  r_n_230__16_,r_n_230__15_,r_n_230__14_,r_n_230__13_,r_n_230__12_,r_n_230__11_,
  r_n_230__10_,r_n_230__9_,r_n_230__8_,r_n_230__7_,r_n_230__6_,r_n_230__5_,
  r_n_230__4_,r_n_230__3_,r_n_230__2_,r_n_230__1_,r_n_230__0_,r_n_229__31_,r_n_229__30_,
  r_n_229__29_,r_n_229__28_,r_n_229__27_,r_n_229__26_,r_n_229__25_,r_n_229__24_,
  r_n_229__23_,r_n_229__22_,r_n_229__21_,r_n_229__20_,r_n_229__19_,r_n_229__18_,
  r_n_229__17_,r_n_229__16_,r_n_229__15_,r_n_229__14_,r_n_229__13_,r_n_229__12_,
  r_n_229__11_,r_n_229__10_,r_n_229__9_,r_n_229__8_,r_n_229__7_,r_n_229__6_,r_n_229__5_,
  r_n_229__4_,r_n_229__3_,r_n_229__2_,r_n_229__1_,r_n_229__0_,r_n_228__31_,
  r_n_228__30_,r_n_228__29_,r_n_228__28_,r_n_228__27_,r_n_228__26_,r_n_228__25_,
  r_n_228__24_,r_n_228__23_,r_n_228__22_,r_n_228__21_,r_n_228__20_,r_n_228__19_,r_n_228__18_,
  r_n_228__17_,r_n_228__16_,r_n_228__15_,r_n_228__14_,r_n_228__13_,r_n_228__12_,
  r_n_228__11_,r_n_228__10_,r_n_228__9_,r_n_228__8_,r_n_228__7_,r_n_228__6_,
  r_n_228__5_,r_n_228__4_,r_n_228__3_,r_n_228__2_,r_n_228__1_,r_n_228__0_,r_n_227__31_,
  r_n_227__30_,r_n_227__29_,r_n_227__28_,r_n_227__27_,r_n_227__26_,r_n_227__25_,
  r_n_227__24_,r_n_227__23_,r_n_227__22_,r_n_227__21_,r_n_227__20_,r_n_227__19_,
  r_n_227__18_,r_n_227__17_,r_n_227__16_,r_n_227__15_,r_n_227__14_,r_n_227__13_,
  r_n_227__12_,r_n_227__11_,r_n_227__10_,r_n_227__9_,r_n_227__8_,r_n_227__7_,r_n_227__6_,
  r_n_227__5_,r_n_227__4_,r_n_227__3_,r_n_227__2_,r_n_227__1_,r_n_227__0_,
  r_n_226__31_,r_n_226__30_,r_n_226__29_,r_n_226__28_,r_n_226__27_,r_n_226__26_,r_n_226__25_,
  r_n_226__24_,r_n_226__23_,r_n_226__22_,r_n_226__21_,r_n_226__20_,r_n_226__19_,
  r_n_226__18_,r_n_226__17_,r_n_226__16_,r_n_226__15_,r_n_226__14_,r_n_226__13_,
  r_n_226__12_,r_n_226__11_,r_n_226__10_,r_n_226__9_,r_n_226__8_,r_n_226__7_,
  r_n_226__6_,r_n_226__5_,r_n_226__4_,r_n_226__3_,r_n_226__2_,r_n_226__1_,r_n_226__0_,
  r_n_225__31_,r_n_225__30_,r_n_225__29_,r_n_225__28_,r_n_225__27_,r_n_225__26_,
  r_n_225__25_,r_n_225__24_,r_n_225__23_,r_n_225__22_,r_n_225__21_,r_n_225__20_,
  r_n_225__19_,r_n_225__18_,r_n_225__17_,r_n_225__16_,r_n_225__15_,r_n_225__14_,
  r_n_225__13_,r_n_225__12_,r_n_225__11_,r_n_225__10_,r_n_225__9_,r_n_225__8_,r_n_225__7_,
  r_n_225__6_,r_n_225__5_,r_n_225__4_,r_n_225__3_,r_n_225__2_,r_n_225__1_,
  r_n_225__0_,r_n_255__31_,r_n_255__30_,r_n_255__29_,r_n_255__28_,r_n_255__27_,r_n_255__26_,
  r_n_255__25_,r_n_255__24_,r_n_255__23_,r_n_255__22_,r_n_255__21_,r_n_255__20_,
  r_n_255__19_,r_n_255__18_,r_n_255__17_,r_n_255__16_,r_n_255__15_,r_n_255__14_,
  r_n_255__13_,r_n_255__12_,r_n_255__11_,r_n_255__10_,r_n_255__9_,r_n_255__8_,
  r_n_255__7_,r_n_255__6_,r_n_255__5_,r_n_255__4_,r_n_255__3_,r_n_255__2_,r_n_255__1_,
  r_n_255__0_,r_n_254__31_,r_n_254__30_,r_n_254__29_,r_n_254__28_,r_n_254__27_,
  r_n_254__26_,r_n_254__25_,r_n_254__24_,r_n_254__23_,r_n_254__22_,r_n_254__21_,
  r_n_254__20_,r_n_254__19_,r_n_254__18_,r_n_254__17_,r_n_254__16_,r_n_254__15_,
  r_n_254__14_,r_n_254__13_,r_n_254__12_,r_n_254__11_,r_n_254__10_,r_n_254__9_,r_n_254__8_,
  r_n_254__7_,r_n_254__6_,r_n_254__5_,r_n_254__4_,r_n_254__3_,r_n_254__2_,
  r_n_254__1_,r_n_254__0_,r_n_253__31_,r_n_253__30_,r_n_253__29_,r_n_253__28_,r_n_253__27_,
  r_n_253__26_,r_n_253__25_,r_n_253__24_,r_n_253__23_,r_n_253__22_,r_n_253__21_,
  r_n_253__20_,r_n_253__19_,r_n_253__18_,r_n_253__17_,r_n_253__16_,r_n_253__15_,
  r_n_253__14_,r_n_253__13_,r_n_253__12_,r_n_253__11_,r_n_253__10_,r_n_253__9_,
  r_n_253__8_,r_n_253__7_,r_n_253__6_,r_n_253__5_,r_n_253__4_,r_n_253__3_,r_n_253__2_,
  r_n_253__1_,r_n_253__0_,r_n_252__31_,r_n_252__30_,r_n_252__29_,r_n_252__28_,
  r_n_252__27_,r_n_252__26_,r_n_252__25_,r_n_252__24_,r_n_252__23_,r_n_252__22_,
  r_n_252__21_,r_n_252__20_,r_n_252__19_,r_n_252__18_,r_n_252__17_,r_n_252__16_,r_n_252__15_,
  r_n_252__14_,r_n_252__13_,r_n_252__12_,r_n_252__11_,r_n_252__10_,r_n_252__9_,
  r_n_252__8_,r_n_252__7_,r_n_252__6_,r_n_252__5_,r_n_252__4_,r_n_252__3_,
  r_n_252__2_,r_n_252__1_,r_n_252__0_,r_n_251__31_,r_n_251__30_,r_n_251__29_,r_n_251__28_,
  r_n_251__27_,r_n_251__26_,r_n_251__25_,r_n_251__24_,r_n_251__23_,r_n_251__22_,
  r_n_251__21_,r_n_251__20_,r_n_251__19_,r_n_251__18_,r_n_251__17_,r_n_251__16_,
  r_n_251__15_,r_n_251__14_,r_n_251__13_,r_n_251__12_,r_n_251__11_,r_n_251__10_,
  r_n_251__9_,r_n_251__8_,r_n_251__7_,r_n_251__6_,r_n_251__5_,r_n_251__4_,r_n_251__3_,
  r_n_251__2_,r_n_251__1_,r_n_251__0_,r_n_250__31_,r_n_250__30_,r_n_250__29_,
  r_n_250__28_,r_n_250__27_,r_n_250__26_,r_n_250__25_,r_n_250__24_,r_n_250__23_,
  r_n_250__22_,r_n_250__21_,r_n_250__20_,r_n_250__19_,r_n_250__18_,r_n_250__17_,r_n_250__16_,
  r_n_250__15_,r_n_250__14_,r_n_250__13_,r_n_250__12_,r_n_250__11_,r_n_250__10_,
  r_n_250__9_,r_n_250__8_,r_n_250__7_,r_n_250__6_,r_n_250__5_,r_n_250__4_,
  r_n_250__3_,r_n_250__2_,r_n_250__1_,r_n_250__0_,r_n_249__31_,r_n_249__30_,r_n_249__29_,
  r_n_249__28_,r_n_249__27_,r_n_249__26_,r_n_249__25_,r_n_249__24_,r_n_249__23_,
  r_n_249__22_,r_n_249__21_,r_n_249__20_,r_n_249__19_,r_n_249__18_,r_n_249__17_,
  r_n_249__16_,r_n_249__15_,r_n_249__14_,r_n_249__13_,r_n_249__12_,r_n_249__11_,
  r_n_249__10_,r_n_249__9_,r_n_249__8_,r_n_249__7_,r_n_249__6_,r_n_249__5_,r_n_249__4_,
  r_n_249__3_,r_n_249__2_,r_n_249__1_,r_n_249__0_,r_n_248__31_,r_n_248__30_,
  r_n_248__29_,r_n_248__28_,r_n_248__27_,r_n_248__26_,r_n_248__25_,r_n_248__24_,r_n_248__23_,
  r_n_248__22_,r_n_248__21_,r_n_248__20_,r_n_248__19_,r_n_248__18_,r_n_248__17_,
  r_n_248__16_,r_n_248__15_,r_n_248__14_,r_n_248__13_,r_n_248__12_,r_n_248__11_,
  r_n_248__10_,r_n_248__9_,r_n_248__8_,r_n_248__7_,r_n_248__6_,r_n_248__5_,
  r_n_248__4_,r_n_248__3_,r_n_248__2_,r_n_248__1_,r_n_248__0_,r_n_247__31_,r_n_247__30_,
  r_n_247__29_,r_n_247__28_,r_n_247__27_,r_n_247__26_,r_n_247__25_,r_n_247__24_,
  r_n_247__23_,r_n_247__22_,r_n_247__21_,r_n_247__20_,r_n_247__19_,r_n_247__18_,
  r_n_247__17_,r_n_247__16_,r_n_247__15_,r_n_247__14_,r_n_247__13_,r_n_247__12_,
  r_n_247__11_,r_n_247__10_,r_n_247__9_,r_n_247__8_,r_n_247__7_,r_n_247__6_,r_n_247__5_,
  r_n_247__4_,r_n_247__3_,r_n_247__2_,r_n_247__1_,r_n_247__0_,r_n_246__31_,
  r_n_246__30_,r_n_246__29_,r_n_246__28_,r_n_246__27_,r_n_246__26_,r_n_246__25_,r_n_246__24_,
  r_n_246__23_,r_n_246__22_,r_n_246__21_,r_n_246__20_,r_n_246__19_,r_n_246__18_,
  r_n_246__17_,r_n_246__16_,r_n_246__15_,r_n_246__14_,r_n_246__13_,r_n_246__12_,
  r_n_246__11_,r_n_246__10_,r_n_246__9_,r_n_246__8_,r_n_246__7_,r_n_246__6_,
  r_n_246__5_,r_n_246__4_,r_n_246__3_,r_n_246__2_,r_n_246__1_,r_n_246__0_,r_n_245__31_,
  r_n_245__30_,r_n_245__29_,r_n_245__28_,r_n_245__27_,r_n_245__26_,r_n_245__25_,
  r_n_245__24_,r_n_245__23_,r_n_245__22_,r_n_245__21_,r_n_245__20_,r_n_245__19_,
  r_n_245__18_,r_n_245__17_,r_n_245__16_,r_n_245__15_,r_n_245__14_,r_n_245__13_,
  r_n_245__12_,r_n_245__11_,r_n_245__10_,r_n_245__9_,r_n_245__8_,r_n_245__7_,r_n_245__6_,
  r_n_245__5_,r_n_245__4_,r_n_245__3_,r_n_245__2_,r_n_245__1_,r_n_245__0_,r_n_244__31_,
  r_n_244__30_,r_n_244__29_,r_n_244__28_,r_n_244__27_,r_n_244__26_,r_n_244__25_,
  r_n_244__24_,r_n_244__23_,r_n_244__22_,r_n_244__21_,r_n_244__20_,r_n_244__19_,
  r_n_244__18_,r_n_244__17_,r_n_244__16_,r_n_244__15_,r_n_244__14_,r_n_244__13_,
  r_n_244__12_,r_n_244__11_,r_n_244__10_,r_n_244__9_,r_n_244__8_,r_n_244__7_,
  r_n_244__6_,r_n_244__5_,r_n_244__4_,r_n_244__3_,r_n_244__2_,r_n_244__1_,r_n_244__0_,
  r_n_243__31_,r_n_243__30_,r_n_243__29_,r_n_243__28_,r_n_243__27_,r_n_243__26_,
  r_n_243__25_,r_n_243__24_,r_n_243__23_,r_n_243__22_,r_n_243__21_,r_n_243__20_,
  r_n_243__19_,r_n_243__18_,r_n_243__17_,r_n_243__16_,r_n_243__15_,r_n_243__14_,r_n_243__13_,
  r_n_243__12_,r_n_243__11_,r_n_243__10_,r_n_243__9_,r_n_243__8_,r_n_243__7_,
  r_n_243__6_,r_n_243__5_,r_n_243__4_,r_n_243__3_,r_n_243__2_,r_n_243__1_,r_n_243__0_,
  r_n_242__31_,r_n_242__30_,r_n_242__29_,r_n_242__28_,r_n_242__27_,r_n_242__26_,
  r_n_242__25_,r_n_242__24_,r_n_242__23_,r_n_242__22_,r_n_242__21_,r_n_242__20_,
  r_n_242__19_,r_n_242__18_,r_n_242__17_,r_n_242__16_,r_n_242__15_,r_n_242__14_,
  r_n_242__13_,r_n_242__12_,r_n_242__11_,r_n_242__10_,r_n_242__9_,r_n_242__8_,
  r_n_242__7_,r_n_242__6_,r_n_242__5_,r_n_242__4_,r_n_242__3_,r_n_242__2_,r_n_242__1_,
  r_n_242__0_,r_n_241__31_,r_n_241__30_,r_n_241__29_,r_n_241__28_,r_n_241__27_,
  r_n_241__26_,r_n_241__25_,r_n_241__24_,r_n_241__23_,r_n_241__22_,r_n_241__21_,
  r_n_241__20_,r_n_241__19_,r_n_241__18_,r_n_241__17_,r_n_241__16_,r_n_241__15_,r_n_241__14_,
  r_n_241__13_,r_n_241__12_,r_n_241__11_,r_n_241__10_,r_n_241__9_,r_n_241__8_,
  r_n_241__7_,r_n_241__6_,r_n_241__5_,r_n_241__4_,r_n_241__3_,r_n_241__2_,r_n_241__1_,
  r_n_241__0_,N517,N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
  N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,
  N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,
  N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,
  N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
  N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,
  N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,
  N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,
  N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,
  N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,
  N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,
  N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,
  N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,
  N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,
  N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
  N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,
  N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,
  N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,
  N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,
  N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,
  N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,
  N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,
  N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,
  N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,
  N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,
  N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,
  N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,
  N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,
  N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,
  N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,
  N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,
  N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,
  N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,
  N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,
  N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,
  N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,
  N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,
  N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,
  N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,
  N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,
  N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,
  N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,
  N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,
  N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,
  N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,
  N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,
  N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,
  N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,
  N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,
  N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,
  N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,
  N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,
  N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,
  N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,
  N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,
  N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,
  N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,
  N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,
  N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,
  N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,
  N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,
  N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,
  N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,
  N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,
  N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,
  N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,
  N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,
  N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,
  N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,
  N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,
  N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,
  N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,
  N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,
  N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,
  N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,
  N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,
  N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,
  N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,
  N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,
  N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,
  N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,
  N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,
  N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,
  N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,
  N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,
  N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,
  N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,
  N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,
  N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,
  N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,
  N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,
  N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,
  N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,
  N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,
  N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,
  N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,
  N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,
  N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,
  N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,
  N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,
  N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,
  N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,
  N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,
  N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,
  N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,
  N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,
  N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,
  N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,
  N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047;
  reg [31:0] data_o;
  reg r_1__31_,r_1__30_,r_1__29_,r_1__28_,r_1__27_,r_1__26_,r_1__25_,r_1__24_,
  r_1__23_,r_1__22_,r_1__21_,r_1__20_,r_1__19_,r_1__18_,r_1__17_,r_1__16_,r_1__15_,
  r_1__14_,r_1__13_,r_1__12_,r_1__11_,r_1__10_,r_1__9_,r_1__8_,r_1__7_,r_1__6_,r_1__5_,
  r_1__4_,r_1__3_,r_1__2_,r_1__1_,r_1__0_,r_2__31_,r_2__30_,r_2__29_,r_2__28_,
  r_2__27_,r_2__26_,r_2__25_,r_2__24_,r_2__23_,r_2__22_,r_2__21_,r_2__20_,r_2__19_,
  r_2__18_,r_2__17_,r_2__16_,r_2__15_,r_2__14_,r_2__13_,r_2__12_,r_2__11_,r_2__10_,
  r_2__9_,r_2__8_,r_2__7_,r_2__6_,r_2__5_,r_2__4_,r_2__3_,r_2__2_,r_2__1_,r_2__0_,
  r_3__31_,r_3__30_,r_3__29_,r_3__28_,r_3__27_,r_3__26_,r_3__25_,r_3__24_,r_3__23_,
  r_3__22_,r_3__21_,r_3__20_,r_3__19_,r_3__18_,r_3__17_,r_3__16_,r_3__15_,r_3__14_,
  r_3__13_,r_3__12_,r_3__11_,r_3__10_,r_3__9_,r_3__8_,r_3__7_,r_3__6_,r_3__5_,
  r_3__4_,r_3__3_,r_3__2_,r_3__1_,r_3__0_,r_4__31_,r_4__30_,r_4__29_,r_4__28_,r_4__27_,
  r_4__26_,r_4__25_,r_4__24_,r_4__23_,r_4__22_,r_4__21_,r_4__20_,r_4__19_,r_4__18_,
  r_4__17_,r_4__16_,r_4__15_,r_4__14_,r_4__13_,r_4__12_,r_4__11_,r_4__10_,r_4__9_,
  r_4__8_,r_4__7_,r_4__6_,r_4__5_,r_4__4_,r_4__3_,r_4__2_,r_4__1_,r_4__0_,
  r_5__31_,r_5__30_,r_5__29_,r_5__28_,r_5__27_,r_5__26_,r_5__25_,r_5__24_,r_5__23_,
  r_5__22_,r_5__21_,r_5__20_,r_5__19_,r_5__18_,r_5__17_,r_5__16_,r_5__15_,r_5__14_,
  r_5__13_,r_5__12_,r_5__11_,r_5__10_,r_5__9_,r_5__8_,r_5__7_,r_5__6_,r_5__5_,r_5__4_,
  r_5__3_,r_5__2_,r_5__1_,r_5__0_,r_6__31_,r_6__30_,r_6__29_,r_6__28_,r_6__27_,
  r_6__26_,r_6__25_,r_6__24_,r_6__23_,r_6__22_,r_6__21_,r_6__20_,r_6__19_,r_6__18_,
  r_6__17_,r_6__16_,r_6__15_,r_6__14_,r_6__13_,r_6__12_,r_6__11_,r_6__10_,r_6__9_,
  r_6__8_,r_6__7_,r_6__6_,r_6__5_,r_6__4_,r_6__3_,r_6__2_,r_6__1_,r_6__0_,r_7__31_,
  r_7__30_,r_7__29_,r_7__28_,r_7__27_,r_7__26_,r_7__25_,r_7__24_,r_7__23_,r_7__22_,
  r_7__21_,r_7__20_,r_7__19_,r_7__18_,r_7__17_,r_7__16_,r_7__15_,r_7__14_,r_7__13_,
  r_7__12_,r_7__11_,r_7__10_,r_7__9_,r_7__8_,r_7__7_,r_7__6_,r_7__5_,r_7__4_,
  r_7__3_,r_7__2_,r_7__1_,r_7__0_,r_8__31_,r_8__30_,r_8__29_,r_8__28_,r_8__27_,r_8__26_,
  r_8__25_,r_8__24_,r_8__23_,r_8__22_,r_8__21_,r_8__20_,r_8__19_,r_8__18_,
  r_8__17_,r_8__16_,r_8__15_,r_8__14_,r_8__13_,r_8__12_,r_8__11_,r_8__10_,r_8__9_,r_8__8_,
  r_8__7_,r_8__6_,r_8__5_,r_8__4_,r_8__3_,r_8__2_,r_8__1_,r_8__0_,r_9__31_,
  r_9__30_,r_9__29_,r_9__28_,r_9__27_,r_9__26_,r_9__25_,r_9__24_,r_9__23_,r_9__22_,
  r_9__21_,r_9__20_,r_9__19_,r_9__18_,r_9__17_,r_9__16_,r_9__15_,r_9__14_,r_9__13_,
  r_9__12_,r_9__11_,r_9__10_,r_9__9_,r_9__8_,r_9__7_,r_9__6_,r_9__5_,r_9__4_,r_9__3_,
  r_9__2_,r_9__1_,r_9__0_,r_10__31_,r_10__30_,r_10__29_,r_10__28_,r_10__27_,
  r_10__26_,r_10__25_,r_10__24_,r_10__23_,r_10__22_,r_10__21_,r_10__20_,r_10__19_,
  r_10__18_,r_10__17_,r_10__16_,r_10__15_,r_10__14_,r_10__13_,r_10__12_,r_10__11_,
  r_10__10_,r_10__9_,r_10__8_,r_10__7_,r_10__6_,r_10__5_,r_10__4_,r_10__3_,r_10__2_,
  r_10__1_,r_10__0_,r_11__31_,r_11__30_,r_11__29_,r_11__28_,r_11__27_,r_11__26_,
  r_11__25_,r_11__24_,r_11__23_,r_11__22_,r_11__21_,r_11__20_,r_11__19_,r_11__18_,
  r_11__17_,r_11__16_,r_11__15_,r_11__14_,r_11__13_,r_11__12_,r_11__11_,r_11__10_,
  r_11__9_,r_11__8_,r_11__7_,r_11__6_,r_11__5_,r_11__4_,r_11__3_,r_11__2_,r_11__1_,
  r_11__0_,r_12__31_,r_12__30_,r_12__29_,r_12__28_,r_12__27_,r_12__26_,r_12__25_,
  r_12__24_,r_12__23_,r_12__22_,r_12__21_,r_12__20_,r_12__19_,r_12__18_,r_12__17_,
  r_12__16_,r_12__15_,r_12__14_,r_12__13_,r_12__12_,r_12__11_,r_12__10_,r_12__9_,r_12__8_,
  r_12__7_,r_12__6_,r_12__5_,r_12__4_,r_12__3_,r_12__2_,r_12__1_,r_12__0_,
  r_13__31_,r_13__30_,r_13__29_,r_13__28_,r_13__27_,r_13__26_,r_13__25_,r_13__24_,
  r_13__23_,r_13__22_,r_13__21_,r_13__20_,r_13__19_,r_13__18_,r_13__17_,r_13__16_,
  r_13__15_,r_13__14_,r_13__13_,r_13__12_,r_13__11_,r_13__10_,r_13__9_,r_13__8_,r_13__7_,
  r_13__6_,r_13__5_,r_13__4_,r_13__3_,r_13__2_,r_13__1_,r_13__0_,r_14__31_,
  r_14__30_,r_14__29_,r_14__28_,r_14__27_,r_14__26_,r_14__25_,r_14__24_,r_14__23_,
  r_14__22_,r_14__21_,r_14__20_,r_14__19_,r_14__18_,r_14__17_,r_14__16_,r_14__15_,
  r_14__14_,r_14__13_,r_14__12_,r_14__11_,r_14__10_,r_14__9_,r_14__8_,r_14__7_,r_14__6_,
  r_14__5_,r_14__4_,r_14__3_,r_14__2_,r_14__1_,r_14__0_,r_15__31_,r_15__30_,
  r_15__29_,r_15__28_,r_15__27_,r_15__26_,r_15__25_,r_15__24_,r_15__23_,r_15__22_,
  r_15__21_,r_15__20_,r_15__19_,r_15__18_,r_15__17_,r_15__16_,r_15__15_,r_15__14_,
  r_15__13_,r_15__12_,r_15__11_,r_15__10_,r_15__9_,r_15__8_,r_15__7_,r_15__6_,r_15__5_,
  r_15__4_,r_15__3_,r_15__2_,r_15__1_,r_15__0_,r_16__31_,r_16__30_,r_16__29_,
  r_16__28_,r_16__27_,r_16__26_,r_16__25_,r_16__24_,r_16__23_,r_16__22_,r_16__21_,
  r_16__20_,r_16__19_,r_16__18_,r_16__17_,r_16__16_,r_16__15_,r_16__14_,r_16__13_,
  r_16__12_,r_16__11_,r_16__10_,r_16__9_,r_16__8_,r_16__7_,r_16__6_,r_16__5_,r_16__4_,
  r_16__3_,r_16__2_,r_16__1_,r_16__0_,r_17__31_,r_17__30_,r_17__29_,r_17__28_,
  r_17__27_,r_17__26_,r_17__25_,r_17__24_,r_17__23_,r_17__22_,r_17__21_,r_17__20_,
  r_17__19_,r_17__18_,r_17__17_,r_17__16_,r_17__15_,r_17__14_,r_17__13_,r_17__12_,
  r_17__11_,r_17__10_,r_17__9_,r_17__8_,r_17__7_,r_17__6_,r_17__5_,r_17__4_,r_17__3_,
  r_17__2_,r_17__1_,r_17__0_,r_18__31_,r_18__30_,r_18__29_,r_18__28_,r_18__27_,
  r_18__26_,r_18__25_,r_18__24_,r_18__23_,r_18__22_,r_18__21_,r_18__20_,r_18__19_,
  r_18__18_,r_18__17_,r_18__16_,r_18__15_,r_18__14_,r_18__13_,r_18__12_,r_18__11_,
  r_18__10_,r_18__9_,r_18__8_,r_18__7_,r_18__6_,r_18__5_,r_18__4_,r_18__3_,r_18__2_,
  r_18__1_,r_18__0_,r_19__31_,r_19__30_,r_19__29_,r_19__28_,r_19__27_,r_19__26_,
  r_19__25_,r_19__24_,r_19__23_,r_19__22_,r_19__21_,r_19__20_,r_19__19_,r_19__18_,
  r_19__17_,r_19__16_,r_19__15_,r_19__14_,r_19__13_,r_19__12_,r_19__11_,r_19__10_,
  r_19__9_,r_19__8_,r_19__7_,r_19__6_,r_19__5_,r_19__4_,r_19__3_,r_19__2_,r_19__1_,
  r_19__0_,r_20__31_,r_20__30_,r_20__29_,r_20__28_,r_20__27_,r_20__26_,r_20__25_,
  r_20__24_,r_20__23_,r_20__22_,r_20__21_,r_20__20_,r_20__19_,r_20__18_,r_20__17_,
  r_20__16_,r_20__15_,r_20__14_,r_20__13_,r_20__12_,r_20__11_,r_20__10_,r_20__9_,r_20__8_,
  r_20__7_,r_20__6_,r_20__5_,r_20__4_,r_20__3_,r_20__2_,r_20__1_,r_20__0_,
  r_21__31_,r_21__30_,r_21__29_,r_21__28_,r_21__27_,r_21__26_,r_21__25_,r_21__24_,
  r_21__23_,r_21__22_,r_21__21_,r_21__20_,r_21__19_,r_21__18_,r_21__17_,r_21__16_,
  r_21__15_,r_21__14_,r_21__13_,r_21__12_,r_21__11_,r_21__10_,r_21__9_,r_21__8_,r_21__7_,
  r_21__6_,r_21__5_,r_21__4_,r_21__3_,r_21__2_,r_21__1_,r_21__0_,r_22__31_,
  r_22__30_,r_22__29_,r_22__28_,r_22__27_,r_22__26_,r_22__25_,r_22__24_,r_22__23_,
  r_22__22_,r_22__21_,r_22__20_,r_22__19_,r_22__18_,r_22__17_,r_22__16_,r_22__15_,
  r_22__14_,r_22__13_,r_22__12_,r_22__11_,r_22__10_,r_22__9_,r_22__8_,r_22__7_,r_22__6_,
  r_22__5_,r_22__4_,r_22__3_,r_22__2_,r_22__1_,r_22__0_,r_23__31_,r_23__30_,
  r_23__29_,r_23__28_,r_23__27_,r_23__26_,r_23__25_,r_23__24_,r_23__23_,r_23__22_,
  r_23__21_,r_23__20_,r_23__19_,r_23__18_,r_23__17_,r_23__16_,r_23__15_,r_23__14_,
  r_23__13_,r_23__12_,r_23__11_,r_23__10_,r_23__9_,r_23__8_,r_23__7_,r_23__6_,r_23__5_,
  r_23__4_,r_23__3_,r_23__2_,r_23__1_,r_23__0_,r_24__31_,r_24__30_,r_24__29_,
  r_24__28_,r_24__27_,r_24__26_,r_24__25_,r_24__24_,r_24__23_,r_24__22_,r_24__21_,
  r_24__20_,r_24__19_,r_24__18_,r_24__17_,r_24__16_,r_24__15_,r_24__14_,r_24__13_,
  r_24__12_,r_24__11_,r_24__10_,r_24__9_,r_24__8_,r_24__7_,r_24__6_,r_24__5_,r_24__4_,
  r_24__3_,r_24__2_,r_24__1_,r_24__0_,r_25__31_,r_25__30_,r_25__29_,r_25__28_,
  r_25__27_,r_25__26_,r_25__25_,r_25__24_,r_25__23_,r_25__22_,r_25__21_,r_25__20_,
  r_25__19_,r_25__18_,r_25__17_,r_25__16_,r_25__15_,r_25__14_,r_25__13_,r_25__12_,
  r_25__11_,r_25__10_,r_25__9_,r_25__8_,r_25__7_,r_25__6_,r_25__5_,r_25__4_,r_25__3_,
  r_25__2_,r_25__1_,r_25__0_,r_26__31_,r_26__30_,r_26__29_,r_26__28_,r_26__27_,
  r_26__26_,r_26__25_,r_26__24_,r_26__23_,r_26__22_,r_26__21_,r_26__20_,r_26__19_,
  r_26__18_,r_26__17_,r_26__16_,r_26__15_,r_26__14_,r_26__13_,r_26__12_,r_26__11_,
  r_26__10_,r_26__9_,r_26__8_,r_26__7_,r_26__6_,r_26__5_,r_26__4_,r_26__3_,r_26__2_,
  r_26__1_,r_26__0_,r_27__31_,r_27__30_,r_27__29_,r_27__28_,r_27__27_,r_27__26_,
  r_27__25_,r_27__24_,r_27__23_,r_27__22_,r_27__21_,r_27__20_,r_27__19_,r_27__18_,
  r_27__17_,r_27__16_,r_27__15_,r_27__14_,r_27__13_,r_27__12_,r_27__11_,r_27__10_,
  r_27__9_,r_27__8_,r_27__7_,r_27__6_,r_27__5_,r_27__4_,r_27__3_,r_27__2_,r_27__1_,
  r_27__0_,r_28__31_,r_28__30_,r_28__29_,r_28__28_,r_28__27_,r_28__26_,r_28__25_,
  r_28__24_,r_28__23_,r_28__22_,r_28__21_,r_28__20_,r_28__19_,r_28__18_,r_28__17_,
  r_28__16_,r_28__15_,r_28__14_,r_28__13_,r_28__12_,r_28__11_,r_28__10_,r_28__9_,r_28__8_,
  r_28__7_,r_28__6_,r_28__5_,r_28__4_,r_28__3_,r_28__2_,r_28__1_,r_28__0_,
  r_29__31_,r_29__30_,r_29__29_,r_29__28_,r_29__27_,r_29__26_,r_29__25_,r_29__24_,
  r_29__23_,r_29__22_,r_29__21_,r_29__20_,r_29__19_,r_29__18_,r_29__17_,r_29__16_,
  r_29__15_,r_29__14_,r_29__13_,r_29__12_,r_29__11_,r_29__10_,r_29__9_,r_29__8_,r_29__7_,
  r_29__6_,r_29__5_,r_29__4_,r_29__3_,r_29__2_,r_29__1_,r_29__0_,r_30__31_,
  r_30__30_,r_30__29_,r_30__28_,r_30__27_,r_30__26_,r_30__25_,r_30__24_,r_30__23_,
  r_30__22_,r_30__21_,r_30__20_,r_30__19_,r_30__18_,r_30__17_,r_30__16_,r_30__15_,
  r_30__14_,r_30__13_,r_30__12_,r_30__11_,r_30__10_,r_30__9_,r_30__8_,r_30__7_,r_30__6_,
  r_30__5_,r_30__4_,r_30__3_,r_30__2_,r_30__1_,r_30__0_,r_31__31_,r_31__30_,
  r_31__29_,r_31__28_,r_31__27_,r_31__26_,r_31__25_,r_31__24_,r_31__23_,r_31__22_,
  r_31__21_,r_31__20_,r_31__19_,r_31__18_,r_31__17_,r_31__16_,r_31__15_,r_31__14_,
  r_31__13_,r_31__12_,r_31__11_,r_31__10_,r_31__9_,r_31__8_,r_31__7_,r_31__6_,r_31__5_,
  r_31__4_,r_31__3_,r_31__2_,r_31__1_,r_31__0_,r_32__31_,r_32__30_,r_32__29_,
  r_32__28_,r_32__27_,r_32__26_,r_32__25_,r_32__24_,r_32__23_,r_32__22_,r_32__21_,
  r_32__20_,r_32__19_,r_32__18_,r_32__17_,r_32__16_,r_32__15_,r_32__14_,r_32__13_,
  r_32__12_,r_32__11_,r_32__10_,r_32__9_,r_32__8_,r_32__7_,r_32__6_,r_32__5_,r_32__4_,
  r_32__3_,r_32__2_,r_32__1_,r_32__0_,r_33__31_,r_33__30_,r_33__29_,r_33__28_,
  r_33__27_,r_33__26_,r_33__25_,r_33__24_,r_33__23_,r_33__22_,r_33__21_,r_33__20_,
  r_33__19_,r_33__18_,r_33__17_,r_33__16_,r_33__15_,r_33__14_,r_33__13_,r_33__12_,
  r_33__11_,r_33__10_,r_33__9_,r_33__8_,r_33__7_,r_33__6_,r_33__5_,r_33__4_,r_33__3_,
  r_33__2_,r_33__1_,r_33__0_,r_34__31_,r_34__30_,r_34__29_,r_34__28_,r_34__27_,
  r_34__26_,r_34__25_,r_34__24_,r_34__23_,r_34__22_,r_34__21_,r_34__20_,r_34__19_,
  r_34__18_,r_34__17_,r_34__16_,r_34__15_,r_34__14_,r_34__13_,r_34__12_,r_34__11_,
  r_34__10_,r_34__9_,r_34__8_,r_34__7_,r_34__6_,r_34__5_,r_34__4_,r_34__3_,r_34__2_,
  r_34__1_,r_34__0_,r_35__31_,r_35__30_,r_35__29_,r_35__28_,r_35__27_,r_35__26_,
  r_35__25_,r_35__24_,r_35__23_,r_35__22_,r_35__21_,r_35__20_,r_35__19_,r_35__18_,
  r_35__17_,r_35__16_,r_35__15_,r_35__14_,r_35__13_,r_35__12_,r_35__11_,r_35__10_,
  r_35__9_,r_35__8_,r_35__7_,r_35__6_,r_35__5_,r_35__4_,r_35__3_,r_35__2_,r_35__1_,
  r_35__0_,r_36__31_,r_36__30_,r_36__29_,r_36__28_,r_36__27_,r_36__26_,r_36__25_,
  r_36__24_,r_36__23_,r_36__22_,r_36__21_,r_36__20_,r_36__19_,r_36__18_,r_36__17_,
  r_36__16_,r_36__15_,r_36__14_,r_36__13_,r_36__12_,r_36__11_,r_36__10_,r_36__9_,r_36__8_,
  r_36__7_,r_36__6_,r_36__5_,r_36__4_,r_36__3_,r_36__2_,r_36__1_,r_36__0_,
  r_37__31_,r_37__30_,r_37__29_,r_37__28_,r_37__27_,r_37__26_,r_37__25_,r_37__24_,
  r_37__23_,r_37__22_,r_37__21_,r_37__20_,r_37__19_,r_37__18_,r_37__17_,r_37__16_,
  r_37__15_,r_37__14_,r_37__13_,r_37__12_,r_37__11_,r_37__10_,r_37__9_,r_37__8_,r_37__7_,
  r_37__6_,r_37__5_,r_37__4_,r_37__3_,r_37__2_,r_37__1_,r_37__0_,r_38__31_,
  r_38__30_,r_38__29_,r_38__28_,r_38__27_,r_38__26_,r_38__25_,r_38__24_,r_38__23_,
  r_38__22_,r_38__21_,r_38__20_,r_38__19_,r_38__18_,r_38__17_,r_38__16_,r_38__15_,
  r_38__14_,r_38__13_,r_38__12_,r_38__11_,r_38__10_,r_38__9_,r_38__8_,r_38__7_,r_38__6_,
  r_38__5_,r_38__4_,r_38__3_,r_38__2_,r_38__1_,r_38__0_,r_39__31_,r_39__30_,
  r_39__29_,r_39__28_,r_39__27_,r_39__26_,r_39__25_,r_39__24_,r_39__23_,r_39__22_,
  r_39__21_,r_39__20_,r_39__19_,r_39__18_,r_39__17_,r_39__16_,r_39__15_,r_39__14_,
  r_39__13_,r_39__12_,r_39__11_,r_39__10_,r_39__9_,r_39__8_,r_39__7_,r_39__6_,r_39__5_,
  r_39__4_,r_39__3_,r_39__2_,r_39__1_,r_39__0_,r_40__31_,r_40__30_,r_40__29_,
  r_40__28_,r_40__27_,r_40__26_,r_40__25_,r_40__24_,r_40__23_,r_40__22_,r_40__21_,
  r_40__20_,r_40__19_,r_40__18_,r_40__17_,r_40__16_,r_40__15_,r_40__14_,r_40__13_,
  r_40__12_,r_40__11_,r_40__10_,r_40__9_,r_40__8_,r_40__7_,r_40__6_,r_40__5_,r_40__4_,
  r_40__3_,r_40__2_,r_40__1_,r_40__0_,r_41__31_,r_41__30_,r_41__29_,r_41__28_,
  r_41__27_,r_41__26_,r_41__25_,r_41__24_,r_41__23_,r_41__22_,r_41__21_,r_41__20_,
  r_41__19_,r_41__18_,r_41__17_,r_41__16_,r_41__15_,r_41__14_,r_41__13_,r_41__12_,
  r_41__11_,r_41__10_,r_41__9_,r_41__8_,r_41__7_,r_41__6_,r_41__5_,r_41__4_,r_41__3_,
  r_41__2_,r_41__1_,r_41__0_,r_42__31_,r_42__30_,r_42__29_,r_42__28_,r_42__27_,
  r_42__26_,r_42__25_,r_42__24_,r_42__23_,r_42__22_,r_42__21_,r_42__20_,r_42__19_,
  r_42__18_,r_42__17_,r_42__16_,r_42__15_,r_42__14_,r_42__13_,r_42__12_,r_42__11_,
  r_42__10_,r_42__9_,r_42__8_,r_42__7_,r_42__6_,r_42__5_,r_42__4_,r_42__3_,r_42__2_,
  r_42__1_,r_42__0_,r_43__31_,r_43__30_,r_43__29_,r_43__28_,r_43__27_,r_43__26_,
  r_43__25_,r_43__24_,r_43__23_,r_43__22_,r_43__21_,r_43__20_,r_43__19_,r_43__18_,
  r_43__17_,r_43__16_,r_43__15_,r_43__14_,r_43__13_,r_43__12_,r_43__11_,r_43__10_,
  r_43__9_,r_43__8_,r_43__7_,r_43__6_,r_43__5_,r_43__4_,r_43__3_,r_43__2_,r_43__1_,
  r_43__0_,r_44__31_,r_44__30_,r_44__29_,r_44__28_,r_44__27_,r_44__26_,r_44__25_,
  r_44__24_,r_44__23_,r_44__22_,r_44__21_,r_44__20_,r_44__19_,r_44__18_,r_44__17_,
  r_44__16_,r_44__15_,r_44__14_,r_44__13_,r_44__12_,r_44__11_,r_44__10_,r_44__9_,r_44__8_,
  r_44__7_,r_44__6_,r_44__5_,r_44__4_,r_44__3_,r_44__2_,r_44__1_,r_44__0_,
  r_45__31_,r_45__30_,r_45__29_,r_45__28_,r_45__27_,r_45__26_,r_45__25_,r_45__24_,
  r_45__23_,r_45__22_,r_45__21_,r_45__20_,r_45__19_,r_45__18_,r_45__17_,r_45__16_,
  r_45__15_,r_45__14_,r_45__13_,r_45__12_,r_45__11_,r_45__10_,r_45__9_,r_45__8_,r_45__7_,
  r_45__6_,r_45__5_,r_45__4_,r_45__3_,r_45__2_,r_45__1_,r_45__0_,r_46__31_,
  r_46__30_,r_46__29_,r_46__28_,r_46__27_,r_46__26_,r_46__25_,r_46__24_,r_46__23_,
  r_46__22_,r_46__21_,r_46__20_,r_46__19_,r_46__18_,r_46__17_,r_46__16_,r_46__15_,
  r_46__14_,r_46__13_,r_46__12_,r_46__11_,r_46__10_,r_46__9_,r_46__8_,r_46__7_,r_46__6_,
  r_46__5_,r_46__4_,r_46__3_,r_46__2_,r_46__1_,r_46__0_,r_47__31_,r_47__30_,
  r_47__29_,r_47__28_,r_47__27_,r_47__26_,r_47__25_,r_47__24_,r_47__23_,r_47__22_,
  r_47__21_,r_47__20_,r_47__19_,r_47__18_,r_47__17_,r_47__16_,r_47__15_,r_47__14_,
  r_47__13_,r_47__12_,r_47__11_,r_47__10_,r_47__9_,r_47__8_,r_47__7_,r_47__6_,r_47__5_,
  r_47__4_,r_47__3_,r_47__2_,r_47__1_,r_47__0_,r_48__31_,r_48__30_,r_48__29_,
  r_48__28_,r_48__27_,r_48__26_,r_48__25_,r_48__24_,r_48__23_,r_48__22_,r_48__21_,
  r_48__20_,r_48__19_,r_48__18_,r_48__17_,r_48__16_,r_48__15_,r_48__14_,r_48__13_,
  r_48__12_,r_48__11_,r_48__10_,r_48__9_,r_48__8_,r_48__7_,r_48__6_,r_48__5_,r_48__4_,
  r_48__3_,r_48__2_,r_48__1_,r_48__0_,r_49__31_,r_49__30_,r_49__29_,r_49__28_,
  r_49__27_,r_49__26_,r_49__25_,r_49__24_,r_49__23_,r_49__22_,r_49__21_,r_49__20_,
  r_49__19_,r_49__18_,r_49__17_,r_49__16_,r_49__15_,r_49__14_,r_49__13_,r_49__12_,
  r_49__11_,r_49__10_,r_49__9_,r_49__8_,r_49__7_,r_49__6_,r_49__5_,r_49__4_,r_49__3_,
  r_49__2_,r_49__1_,r_49__0_,r_50__31_,r_50__30_,r_50__29_,r_50__28_,r_50__27_,
  r_50__26_,r_50__25_,r_50__24_,r_50__23_,r_50__22_,r_50__21_,r_50__20_,r_50__19_,
  r_50__18_,r_50__17_,r_50__16_,r_50__15_,r_50__14_,r_50__13_,r_50__12_,r_50__11_,
  r_50__10_,r_50__9_,r_50__8_,r_50__7_,r_50__6_,r_50__5_,r_50__4_,r_50__3_,r_50__2_,
  r_50__1_,r_50__0_,r_51__31_,r_51__30_,r_51__29_,r_51__28_,r_51__27_,r_51__26_,
  r_51__25_,r_51__24_,r_51__23_,r_51__22_,r_51__21_,r_51__20_,r_51__19_,r_51__18_,
  r_51__17_,r_51__16_,r_51__15_,r_51__14_,r_51__13_,r_51__12_,r_51__11_,r_51__10_,
  r_51__9_,r_51__8_,r_51__7_,r_51__6_,r_51__5_,r_51__4_,r_51__3_,r_51__2_,r_51__1_,
  r_51__0_,r_52__31_,r_52__30_,r_52__29_,r_52__28_,r_52__27_,r_52__26_,r_52__25_,
  r_52__24_,r_52__23_,r_52__22_,r_52__21_,r_52__20_,r_52__19_,r_52__18_,r_52__17_,
  r_52__16_,r_52__15_,r_52__14_,r_52__13_,r_52__12_,r_52__11_,r_52__10_,r_52__9_,r_52__8_,
  r_52__7_,r_52__6_,r_52__5_,r_52__4_,r_52__3_,r_52__2_,r_52__1_,r_52__0_,
  r_53__31_,r_53__30_,r_53__29_,r_53__28_,r_53__27_,r_53__26_,r_53__25_,r_53__24_,
  r_53__23_,r_53__22_,r_53__21_,r_53__20_,r_53__19_,r_53__18_,r_53__17_,r_53__16_,
  r_53__15_,r_53__14_,r_53__13_,r_53__12_,r_53__11_,r_53__10_,r_53__9_,r_53__8_,r_53__7_,
  r_53__6_,r_53__5_,r_53__4_,r_53__3_,r_53__2_,r_53__1_,r_53__0_,r_54__31_,
  r_54__30_,r_54__29_,r_54__28_,r_54__27_,r_54__26_,r_54__25_,r_54__24_,r_54__23_,
  r_54__22_,r_54__21_,r_54__20_,r_54__19_,r_54__18_,r_54__17_,r_54__16_,r_54__15_,
  r_54__14_,r_54__13_,r_54__12_,r_54__11_,r_54__10_,r_54__9_,r_54__8_,r_54__7_,r_54__6_,
  r_54__5_,r_54__4_,r_54__3_,r_54__2_,r_54__1_,r_54__0_,r_55__31_,r_55__30_,
  r_55__29_,r_55__28_,r_55__27_,r_55__26_,r_55__25_,r_55__24_,r_55__23_,r_55__22_,
  r_55__21_,r_55__20_,r_55__19_,r_55__18_,r_55__17_,r_55__16_,r_55__15_,r_55__14_,
  r_55__13_,r_55__12_,r_55__11_,r_55__10_,r_55__9_,r_55__8_,r_55__7_,r_55__6_,r_55__5_,
  r_55__4_,r_55__3_,r_55__2_,r_55__1_,r_55__0_,r_56__31_,r_56__30_,r_56__29_,
  r_56__28_,r_56__27_,r_56__26_,r_56__25_,r_56__24_,r_56__23_,r_56__22_,r_56__21_,
  r_56__20_,r_56__19_,r_56__18_,r_56__17_,r_56__16_,r_56__15_,r_56__14_,r_56__13_,
  r_56__12_,r_56__11_,r_56__10_,r_56__9_,r_56__8_,r_56__7_,r_56__6_,r_56__5_,r_56__4_,
  r_56__3_,r_56__2_,r_56__1_,r_56__0_,r_57__31_,r_57__30_,r_57__29_,r_57__28_,
  r_57__27_,r_57__26_,r_57__25_,r_57__24_,r_57__23_,r_57__22_,r_57__21_,r_57__20_,
  r_57__19_,r_57__18_,r_57__17_,r_57__16_,r_57__15_,r_57__14_,r_57__13_,r_57__12_,
  r_57__11_,r_57__10_,r_57__9_,r_57__8_,r_57__7_,r_57__6_,r_57__5_,r_57__4_,r_57__3_,
  r_57__2_,r_57__1_,r_57__0_,r_58__31_,r_58__30_,r_58__29_,r_58__28_,r_58__27_,
  r_58__26_,r_58__25_,r_58__24_,r_58__23_,r_58__22_,r_58__21_,r_58__20_,r_58__19_,
  r_58__18_,r_58__17_,r_58__16_,r_58__15_,r_58__14_,r_58__13_,r_58__12_,r_58__11_,
  r_58__10_,r_58__9_,r_58__8_,r_58__7_,r_58__6_,r_58__5_,r_58__4_,r_58__3_,r_58__2_,
  r_58__1_,r_58__0_,r_59__31_,r_59__30_,r_59__29_,r_59__28_,r_59__27_,r_59__26_,
  r_59__25_,r_59__24_,r_59__23_,r_59__22_,r_59__21_,r_59__20_,r_59__19_,r_59__18_,
  r_59__17_,r_59__16_,r_59__15_,r_59__14_,r_59__13_,r_59__12_,r_59__11_,r_59__10_,
  r_59__9_,r_59__8_,r_59__7_,r_59__6_,r_59__5_,r_59__4_,r_59__3_,r_59__2_,r_59__1_,
  r_59__0_,r_60__31_,r_60__30_,r_60__29_,r_60__28_,r_60__27_,r_60__26_,r_60__25_,
  r_60__24_,r_60__23_,r_60__22_,r_60__21_,r_60__20_,r_60__19_,r_60__18_,r_60__17_,
  r_60__16_,r_60__15_,r_60__14_,r_60__13_,r_60__12_,r_60__11_,r_60__10_,r_60__9_,r_60__8_,
  r_60__7_,r_60__6_,r_60__5_,r_60__4_,r_60__3_,r_60__2_,r_60__1_,r_60__0_,
  r_61__31_,r_61__30_,r_61__29_,r_61__28_,r_61__27_,r_61__26_,r_61__25_,r_61__24_,
  r_61__23_,r_61__22_,r_61__21_,r_61__20_,r_61__19_,r_61__18_,r_61__17_,r_61__16_,
  r_61__15_,r_61__14_,r_61__13_,r_61__12_,r_61__11_,r_61__10_,r_61__9_,r_61__8_,r_61__7_,
  r_61__6_,r_61__5_,r_61__4_,r_61__3_,r_61__2_,r_61__1_,r_61__0_,r_62__31_,
  r_62__30_,r_62__29_,r_62__28_,r_62__27_,r_62__26_,r_62__25_,r_62__24_,r_62__23_,
  r_62__22_,r_62__21_,r_62__20_,r_62__19_,r_62__18_,r_62__17_,r_62__16_,r_62__15_,
  r_62__14_,r_62__13_,r_62__12_,r_62__11_,r_62__10_,r_62__9_,r_62__8_,r_62__7_,r_62__6_,
  r_62__5_,r_62__4_,r_62__3_,r_62__2_,r_62__1_,r_62__0_,r_63__31_,r_63__30_,
  r_63__29_,r_63__28_,r_63__27_,r_63__26_,r_63__25_,r_63__24_,r_63__23_,r_63__22_,
  r_63__21_,r_63__20_,r_63__19_,r_63__18_,r_63__17_,r_63__16_,r_63__15_,r_63__14_,
  r_63__13_,r_63__12_,r_63__11_,r_63__10_,r_63__9_,r_63__8_,r_63__7_,r_63__6_,r_63__5_,
  r_63__4_,r_63__3_,r_63__2_,r_63__1_,r_63__0_,r_64__31_,r_64__30_,r_64__29_,
  r_64__28_,r_64__27_,r_64__26_,r_64__25_,r_64__24_,r_64__23_,r_64__22_,r_64__21_,
  r_64__20_,r_64__19_,r_64__18_,r_64__17_,r_64__16_,r_64__15_,r_64__14_,r_64__13_,
  r_64__12_,r_64__11_,r_64__10_,r_64__9_,r_64__8_,r_64__7_,r_64__6_,r_64__5_,r_64__4_,
  r_64__3_,r_64__2_,r_64__1_,r_64__0_,r_65__31_,r_65__30_,r_65__29_,r_65__28_,
  r_65__27_,r_65__26_,r_65__25_,r_65__24_,r_65__23_,r_65__22_,r_65__21_,r_65__20_,
  r_65__19_,r_65__18_,r_65__17_,r_65__16_,r_65__15_,r_65__14_,r_65__13_,r_65__12_,
  r_65__11_,r_65__10_,r_65__9_,r_65__8_,r_65__7_,r_65__6_,r_65__5_,r_65__4_,r_65__3_,
  r_65__2_,r_65__1_,r_65__0_,r_66__31_,r_66__30_,r_66__29_,r_66__28_,r_66__27_,
  r_66__26_,r_66__25_,r_66__24_,r_66__23_,r_66__22_,r_66__21_,r_66__20_,r_66__19_,
  r_66__18_,r_66__17_,r_66__16_,r_66__15_,r_66__14_,r_66__13_,r_66__12_,r_66__11_,
  r_66__10_,r_66__9_,r_66__8_,r_66__7_,r_66__6_,r_66__5_,r_66__4_,r_66__3_,r_66__2_,
  r_66__1_,r_66__0_,r_67__31_,r_67__30_,r_67__29_,r_67__28_,r_67__27_,r_67__26_,
  r_67__25_,r_67__24_,r_67__23_,r_67__22_,r_67__21_,r_67__20_,r_67__19_,r_67__18_,
  r_67__17_,r_67__16_,r_67__15_,r_67__14_,r_67__13_,r_67__12_,r_67__11_,r_67__10_,
  r_67__9_,r_67__8_,r_67__7_,r_67__6_,r_67__5_,r_67__4_,r_67__3_,r_67__2_,r_67__1_,
  r_67__0_,r_68__31_,r_68__30_,r_68__29_,r_68__28_,r_68__27_,r_68__26_,r_68__25_,
  r_68__24_,r_68__23_,r_68__22_,r_68__21_,r_68__20_,r_68__19_,r_68__18_,r_68__17_,
  r_68__16_,r_68__15_,r_68__14_,r_68__13_,r_68__12_,r_68__11_,r_68__10_,r_68__9_,r_68__8_,
  r_68__7_,r_68__6_,r_68__5_,r_68__4_,r_68__3_,r_68__2_,r_68__1_,r_68__0_,
  r_69__31_,r_69__30_,r_69__29_,r_69__28_,r_69__27_,r_69__26_,r_69__25_,r_69__24_,
  r_69__23_,r_69__22_,r_69__21_,r_69__20_,r_69__19_,r_69__18_,r_69__17_,r_69__16_,
  r_69__15_,r_69__14_,r_69__13_,r_69__12_,r_69__11_,r_69__10_,r_69__9_,r_69__8_,r_69__7_,
  r_69__6_,r_69__5_,r_69__4_,r_69__3_,r_69__2_,r_69__1_,r_69__0_,r_70__31_,
  r_70__30_,r_70__29_,r_70__28_,r_70__27_,r_70__26_,r_70__25_,r_70__24_,r_70__23_,
  r_70__22_,r_70__21_,r_70__20_,r_70__19_,r_70__18_,r_70__17_,r_70__16_,r_70__15_,
  r_70__14_,r_70__13_,r_70__12_,r_70__11_,r_70__10_,r_70__9_,r_70__8_,r_70__7_,r_70__6_,
  r_70__5_,r_70__4_,r_70__3_,r_70__2_,r_70__1_,r_70__0_,r_71__31_,r_71__30_,
  r_71__29_,r_71__28_,r_71__27_,r_71__26_,r_71__25_,r_71__24_,r_71__23_,r_71__22_,
  r_71__21_,r_71__20_,r_71__19_,r_71__18_,r_71__17_,r_71__16_,r_71__15_,r_71__14_,
  r_71__13_,r_71__12_,r_71__11_,r_71__10_,r_71__9_,r_71__8_,r_71__7_,r_71__6_,r_71__5_,
  r_71__4_,r_71__3_,r_71__2_,r_71__1_,r_71__0_,r_72__31_,r_72__30_,r_72__29_,
  r_72__28_,r_72__27_,r_72__26_,r_72__25_,r_72__24_,r_72__23_,r_72__22_,r_72__21_,
  r_72__20_,r_72__19_,r_72__18_,r_72__17_,r_72__16_,r_72__15_,r_72__14_,r_72__13_,
  r_72__12_,r_72__11_,r_72__10_,r_72__9_,r_72__8_,r_72__7_,r_72__6_,r_72__5_,r_72__4_,
  r_72__3_,r_72__2_,r_72__1_,r_72__0_,r_73__31_,r_73__30_,r_73__29_,r_73__28_,
  r_73__27_,r_73__26_,r_73__25_,r_73__24_,r_73__23_,r_73__22_,r_73__21_,r_73__20_,
  r_73__19_,r_73__18_,r_73__17_,r_73__16_,r_73__15_,r_73__14_,r_73__13_,r_73__12_,
  r_73__11_,r_73__10_,r_73__9_,r_73__8_,r_73__7_,r_73__6_,r_73__5_,r_73__4_,r_73__3_,
  r_73__2_,r_73__1_,r_73__0_,r_74__31_,r_74__30_,r_74__29_,r_74__28_,r_74__27_,
  r_74__26_,r_74__25_,r_74__24_,r_74__23_,r_74__22_,r_74__21_,r_74__20_,r_74__19_,
  r_74__18_,r_74__17_,r_74__16_,r_74__15_,r_74__14_,r_74__13_,r_74__12_,r_74__11_,
  r_74__10_,r_74__9_,r_74__8_,r_74__7_,r_74__6_,r_74__5_,r_74__4_,r_74__3_,r_74__2_,
  r_74__1_,r_74__0_,r_75__31_,r_75__30_,r_75__29_,r_75__28_,r_75__27_,r_75__26_,
  r_75__25_,r_75__24_,r_75__23_,r_75__22_,r_75__21_,r_75__20_,r_75__19_,r_75__18_,
  r_75__17_,r_75__16_,r_75__15_,r_75__14_,r_75__13_,r_75__12_,r_75__11_,r_75__10_,
  r_75__9_,r_75__8_,r_75__7_,r_75__6_,r_75__5_,r_75__4_,r_75__3_,r_75__2_,r_75__1_,
  r_75__0_,r_76__31_,r_76__30_,r_76__29_,r_76__28_,r_76__27_,r_76__26_,r_76__25_,
  r_76__24_,r_76__23_,r_76__22_,r_76__21_,r_76__20_,r_76__19_,r_76__18_,r_76__17_,
  r_76__16_,r_76__15_,r_76__14_,r_76__13_,r_76__12_,r_76__11_,r_76__10_,r_76__9_,r_76__8_,
  r_76__7_,r_76__6_,r_76__5_,r_76__4_,r_76__3_,r_76__2_,r_76__1_,r_76__0_,
  r_77__31_,r_77__30_,r_77__29_,r_77__28_,r_77__27_,r_77__26_,r_77__25_,r_77__24_,
  r_77__23_,r_77__22_,r_77__21_,r_77__20_,r_77__19_,r_77__18_,r_77__17_,r_77__16_,
  r_77__15_,r_77__14_,r_77__13_,r_77__12_,r_77__11_,r_77__10_,r_77__9_,r_77__8_,r_77__7_,
  r_77__6_,r_77__5_,r_77__4_,r_77__3_,r_77__2_,r_77__1_,r_77__0_,r_78__31_,
  r_78__30_,r_78__29_,r_78__28_,r_78__27_,r_78__26_,r_78__25_,r_78__24_,r_78__23_,
  r_78__22_,r_78__21_,r_78__20_,r_78__19_,r_78__18_,r_78__17_,r_78__16_,r_78__15_,
  r_78__14_,r_78__13_,r_78__12_,r_78__11_,r_78__10_,r_78__9_,r_78__8_,r_78__7_,r_78__6_,
  r_78__5_,r_78__4_,r_78__3_,r_78__2_,r_78__1_,r_78__0_,r_79__31_,r_79__30_,
  r_79__29_,r_79__28_,r_79__27_,r_79__26_,r_79__25_,r_79__24_,r_79__23_,r_79__22_,
  r_79__21_,r_79__20_,r_79__19_,r_79__18_,r_79__17_,r_79__16_,r_79__15_,r_79__14_,
  r_79__13_,r_79__12_,r_79__11_,r_79__10_,r_79__9_,r_79__8_,r_79__7_,r_79__6_,r_79__5_,
  r_79__4_,r_79__3_,r_79__2_,r_79__1_,r_79__0_,r_80__31_,r_80__30_,r_80__29_,
  r_80__28_,r_80__27_,r_80__26_,r_80__25_,r_80__24_,r_80__23_,r_80__22_,r_80__21_,
  r_80__20_,r_80__19_,r_80__18_,r_80__17_,r_80__16_,r_80__15_,r_80__14_,r_80__13_,
  r_80__12_,r_80__11_,r_80__10_,r_80__9_,r_80__8_,r_80__7_,r_80__6_,r_80__5_,r_80__4_,
  r_80__3_,r_80__2_,r_80__1_,r_80__0_,r_81__31_,r_81__30_,r_81__29_,r_81__28_,
  r_81__27_,r_81__26_,r_81__25_,r_81__24_,r_81__23_,r_81__22_,r_81__21_,r_81__20_,
  r_81__19_,r_81__18_,r_81__17_,r_81__16_,r_81__15_,r_81__14_,r_81__13_,r_81__12_,
  r_81__11_,r_81__10_,r_81__9_,r_81__8_,r_81__7_,r_81__6_,r_81__5_,r_81__4_,r_81__3_,
  r_81__2_,r_81__1_,r_81__0_,r_82__31_,r_82__30_,r_82__29_,r_82__28_,r_82__27_,
  r_82__26_,r_82__25_,r_82__24_,r_82__23_,r_82__22_,r_82__21_,r_82__20_,r_82__19_,
  r_82__18_,r_82__17_,r_82__16_,r_82__15_,r_82__14_,r_82__13_,r_82__12_,r_82__11_,
  r_82__10_,r_82__9_,r_82__8_,r_82__7_,r_82__6_,r_82__5_,r_82__4_,r_82__3_,r_82__2_,
  r_82__1_,r_82__0_,r_83__31_,r_83__30_,r_83__29_,r_83__28_,r_83__27_,r_83__26_,
  r_83__25_,r_83__24_,r_83__23_,r_83__22_,r_83__21_,r_83__20_,r_83__19_,r_83__18_,
  r_83__17_,r_83__16_,r_83__15_,r_83__14_,r_83__13_,r_83__12_,r_83__11_,r_83__10_,
  r_83__9_,r_83__8_,r_83__7_,r_83__6_,r_83__5_,r_83__4_,r_83__3_,r_83__2_,r_83__1_,
  r_83__0_,r_84__31_,r_84__30_,r_84__29_,r_84__28_,r_84__27_,r_84__26_,r_84__25_,
  r_84__24_,r_84__23_,r_84__22_,r_84__21_,r_84__20_,r_84__19_,r_84__18_,r_84__17_,
  r_84__16_,r_84__15_,r_84__14_,r_84__13_,r_84__12_,r_84__11_,r_84__10_,r_84__9_,r_84__8_,
  r_84__7_,r_84__6_,r_84__5_,r_84__4_,r_84__3_,r_84__2_,r_84__1_,r_84__0_,
  r_85__31_,r_85__30_,r_85__29_,r_85__28_,r_85__27_,r_85__26_,r_85__25_,r_85__24_,
  r_85__23_,r_85__22_,r_85__21_,r_85__20_,r_85__19_,r_85__18_,r_85__17_,r_85__16_,
  r_85__15_,r_85__14_,r_85__13_,r_85__12_,r_85__11_,r_85__10_,r_85__9_,r_85__8_,r_85__7_,
  r_85__6_,r_85__5_,r_85__4_,r_85__3_,r_85__2_,r_85__1_,r_85__0_,r_86__31_,
  r_86__30_,r_86__29_,r_86__28_,r_86__27_,r_86__26_,r_86__25_,r_86__24_,r_86__23_,
  r_86__22_,r_86__21_,r_86__20_,r_86__19_,r_86__18_,r_86__17_,r_86__16_,r_86__15_,
  r_86__14_,r_86__13_,r_86__12_,r_86__11_,r_86__10_,r_86__9_,r_86__8_,r_86__7_,r_86__6_,
  r_86__5_,r_86__4_,r_86__3_,r_86__2_,r_86__1_,r_86__0_,r_87__31_,r_87__30_,
  r_87__29_,r_87__28_,r_87__27_,r_87__26_,r_87__25_,r_87__24_,r_87__23_,r_87__22_,
  r_87__21_,r_87__20_,r_87__19_,r_87__18_,r_87__17_,r_87__16_,r_87__15_,r_87__14_,
  r_87__13_,r_87__12_,r_87__11_,r_87__10_,r_87__9_,r_87__8_,r_87__7_,r_87__6_,r_87__5_,
  r_87__4_,r_87__3_,r_87__2_,r_87__1_,r_87__0_,r_88__31_,r_88__30_,r_88__29_,
  r_88__28_,r_88__27_,r_88__26_,r_88__25_,r_88__24_,r_88__23_,r_88__22_,r_88__21_,
  r_88__20_,r_88__19_,r_88__18_,r_88__17_,r_88__16_,r_88__15_,r_88__14_,r_88__13_,
  r_88__12_,r_88__11_,r_88__10_,r_88__9_,r_88__8_,r_88__7_,r_88__6_,r_88__5_,r_88__4_,
  r_88__3_,r_88__2_,r_88__1_,r_88__0_,r_89__31_,r_89__30_,r_89__29_,r_89__28_,
  r_89__27_,r_89__26_,r_89__25_,r_89__24_,r_89__23_,r_89__22_,r_89__21_,r_89__20_,
  r_89__19_,r_89__18_,r_89__17_,r_89__16_,r_89__15_,r_89__14_,r_89__13_,r_89__12_,
  r_89__11_,r_89__10_,r_89__9_,r_89__8_,r_89__7_,r_89__6_,r_89__5_,r_89__4_,r_89__3_,
  r_89__2_,r_89__1_,r_89__0_,r_90__31_,r_90__30_,r_90__29_,r_90__28_,r_90__27_,
  r_90__26_,r_90__25_,r_90__24_,r_90__23_,r_90__22_,r_90__21_,r_90__20_,r_90__19_,
  r_90__18_,r_90__17_,r_90__16_,r_90__15_,r_90__14_,r_90__13_,r_90__12_,r_90__11_,
  r_90__10_,r_90__9_,r_90__8_,r_90__7_,r_90__6_,r_90__5_,r_90__4_,r_90__3_,r_90__2_,
  r_90__1_,r_90__0_,r_91__31_,r_91__30_,r_91__29_,r_91__28_,r_91__27_,r_91__26_,
  r_91__25_,r_91__24_,r_91__23_,r_91__22_,r_91__21_,r_91__20_,r_91__19_,r_91__18_,
  r_91__17_,r_91__16_,r_91__15_,r_91__14_,r_91__13_,r_91__12_,r_91__11_,r_91__10_,
  r_91__9_,r_91__8_,r_91__7_,r_91__6_,r_91__5_,r_91__4_,r_91__3_,r_91__2_,r_91__1_,
  r_91__0_,r_92__31_,r_92__30_,r_92__29_,r_92__28_,r_92__27_,r_92__26_,r_92__25_,
  r_92__24_,r_92__23_,r_92__22_,r_92__21_,r_92__20_,r_92__19_,r_92__18_,r_92__17_,
  r_92__16_,r_92__15_,r_92__14_,r_92__13_,r_92__12_,r_92__11_,r_92__10_,r_92__9_,r_92__8_,
  r_92__7_,r_92__6_,r_92__5_,r_92__4_,r_92__3_,r_92__2_,r_92__1_,r_92__0_,
  r_93__31_,r_93__30_,r_93__29_,r_93__28_,r_93__27_,r_93__26_,r_93__25_,r_93__24_,
  r_93__23_,r_93__22_,r_93__21_,r_93__20_,r_93__19_,r_93__18_,r_93__17_,r_93__16_,
  r_93__15_,r_93__14_,r_93__13_,r_93__12_,r_93__11_,r_93__10_,r_93__9_,r_93__8_,r_93__7_,
  r_93__6_,r_93__5_,r_93__4_,r_93__3_,r_93__2_,r_93__1_,r_93__0_,r_94__31_,
  r_94__30_,r_94__29_,r_94__28_,r_94__27_,r_94__26_,r_94__25_,r_94__24_,r_94__23_,
  r_94__22_,r_94__21_,r_94__20_,r_94__19_,r_94__18_,r_94__17_,r_94__16_,r_94__15_,
  r_94__14_,r_94__13_,r_94__12_,r_94__11_,r_94__10_,r_94__9_,r_94__8_,r_94__7_,r_94__6_,
  r_94__5_,r_94__4_,r_94__3_,r_94__2_,r_94__1_,r_94__0_,r_95__31_,r_95__30_,
  r_95__29_,r_95__28_,r_95__27_,r_95__26_,r_95__25_,r_95__24_,r_95__23_,r_95__22_,
  r_95__21_,r_95__20_,r_95__19_,r_95__18_,r_95__17_,r_95__16_,r_95__15_,r_95__14_,
  r_95__13_,r_95__12_,r_95__11_,r_95__10_,r_95__9_,r_95__8_,r_95__7_,r_95__6_,r_95__5_,
  r_95__4_,r_95__3_,r_95__2_,r_95__1_,r_95__0_,r_96__31_,r_96__30_,r_96__29_,
  r_96__28_,r_96__27_,r_96__26_,r_96__25_,r_96__24_,r_96__23_,r_96__22_,r_96__21_,
  r_96__20_,r_96__19_,r_96__18_,r_96__17_,r_96__16_,r_96__15_,r_96__14_,r_96__13_,
  r_96__12_,r_96__11_,r_96__10_,r_96__9_,r_96__8_,r_96__7_,r_96__6_,r_96__5_,r_96__4_,
  r_96__3_,r_96__2_,r_96__1_,r_96__0_,r_97__31_,r_97__30_,r_97__29_,r_97__28_,
  r_97__27_,r_97__26_,r_97__25_,r_97__24_,r_97__23_,r_97__22_,r_97__21_,r_97__20_,
  r_97__19_,r_97__18_,r_97__17_,r_97__16_,r_97__15_,r_97__14_,r_97__13_,r_97__12_,
  r_97__11_,r_97__10_,r_97__9_,r_97__8_,r_97__7_,r_97__6_,r_97__5_,r_97__4_,r_97__3_,
  r_97__2_,r_97__1_,r_97__0_,r_98__31_,r_98__30_,r_98__29_,r_98__28_,r_98__27_,
  r_98__26_,r_98__25_,r_98__24_,r_98__23_,r_98__22_,r_98__21_,r_98__20_,r_98__19_,
  r_98__18_,r_98__17_,r_98__16_,r_98__15_,r_98__14_,r_98__13_,r_98__12_,r_98__11_,
  r_98__10_,r_98__9_,r_98__8_,r_98__7_,r_98__6_,r_98__5_,r_98__4_,r_98__3_,r_98__2_,
  r_98__1_,r_98__0_,r_99__31_,r_99__30_,r_99__29_,r_99__28_,r_99__27_,r_99__26_,
  r_99__25_,r_99__24_,r_99__23_,r_99__22_,r_99__21_,r_99__20_,r_99__19_,r_99__18_,
  r_99__17_,r_99__16_,r_99__15_,r_99__14_,r_99__13_,r_99__12_,r_99__11_,r_99__10_,
  r_99__9_,r_99__8_,r_99__7_,r_99__6_,r_99__5_,r_99__4_,r_99__3_,r_99__2_,r_99__1_,
  r_99__0_,r_100__31_,r_100__30_,r_100__29_,r_100__28_,r_100__27_,r_100__26_,r_100__25_,
  r_100__24_,r_100__23_,r_100__22_,r_100__21_,r_100__20_,r_100__19_,r_100__18_,
  r_100__17_,r_100__16_,r_100__15_,r_100__14_,r_100__13_,r_100__12_,r_100__11_,
  r_100__10_,r_100__9_,r_100__8_,r_100__7_,r_100__6_,r_100__5_,r_100__4_,r_100__3_,
  r_100__2_,r_100__1_,r_100__0_,r_101__31_,r_101__30_,r_101__29_,r_101__28_,r_101__27_,
  r_101__26_,r_101__25_,r_101__24_,r_101__23_,r_101__22_,r_101__21_,r_101__20_,
  r_101__19_,r_101__18_,r_101__17_,r_101__16_,r_101__15_,r_101__14_,r_101__13_,
  r_101__12_,r_101__11_,r_101__10_,r_101__9_,r_101__8_,r_101__7_,r_101__6_,r_101__5_,
  r_101__4_,r_101__3_,r_101__2_,r_101__1_,r_101__0_,r_102__31_,r_102__30_,r_102__29_,
  r_102__28_,r_102__27_,r_102__26_,r_102__25_,r_102__24_,r_102__23_,r_102__22_,
  r_102__21_,r_102__20_,r_102__19_,r_102__18_,r_102__17_,r_102__16_,r_102__15_,
  r_102__14_,r_102__13_,r_102__12_,r_102__11_,r_102__10_,r_102__9_,r_102__8_,r_102__7_,
  r_102__6_,r_102__5_,r_102__4_,r_102__3_,r_102__2_,r_102__1_,r_102__0_,r_103__31_,
  r_103__30_,r_103__29_,r_103__28_,r_103__27_,r_103__26_,r_103__25_,r_103__24_,
  r_103__23_,r_103__22_,r_103__21_,r_103__20_,r_103__19_,r_103__18_,r_103__17_,
  r_103__16_,r_103__15_,r_103__14_,r_103__13_,r_103__12_,r_103__11_,r_103__10_,r_103__9_,
  r_103__8_,r_103__7_,r_103__6_,r_103__5_,r_103__4_,r_103__3_,r_103__2_,r_103__1_,
  r_103__0_,r_104__31_,r_104__30_,r_104__29_,r_104__28_,r_104__27_,r_104__26_,
  r_104__25_,r_104__24_,r_104__23_,r_104__22_,r_104__21_,r_104__20_,r_104__19_,
  r_104__18_,r_104__17_,r_104__16_,r_104__15_,r_104__14_,r_104__13_,r_104__12_,
  r_104__11_,r_104__10_,r_104__9_,r_104__8_,r_104__7_,r_104__6_,r_104__5_,r_104__4_,
  r_104__3_,r_104__2_,r_104__1_,r_104__0_,r_105__31_,r_105__30_,r_105__29_,r_105__28_,
  r_105__27_,r_105__26_,r_105__25_,r_105__24_,r_105__23_,r_105__22_,r_105__21_,
  r_105__20_,r_105__19_,r_105__18_,r_105__17_,r_105__16_,r_105__15_,r_105__14_,
  r_105__13_,r_105__12_,r_105__11_,r_105__10_,r_105__9_,r_105__8_,r_105__7_,r_105__6_,
  r_105__5_,r_105__4_,r_105__3_,r_105__2_,r_105__1_,r_105__0_,r_106__31_,r_106__30_,
  r_106__29_,r_106__28_,r_106__27_,r_106__26_,r_106__25_,r_106__24_,r_106__23_,
  r_106__22_,r_106__21_,r_106__20_,r_106__19_,r_106__18_,r_106__17_,r_106__16_,
  r_106__15_,r_106__14_,r_106__13_,r_106__12_,r_106__11_,r_106__10_,r_106__9_,r_106__8_,
  r_106__7_,r_106__6_,r_106__5_,r_106__4_,r_106__3_,r_106__2_,r_106__1_,r_106__0_,
  r_107__31_,r_107__30_,r_107__29_,r_107__28_,r_107__27_,r_107__26_,r_107__25_,
  r_107__24_,r_107__23_,r_107__22_,r_107__21_,r_107__20_,r_107__19_,r_107__18_,
  r_107__17_,r_107__16_,r_107__15_,r_107__14_,r_107__13_,r_107__12_,r_107__11_,r_107__10_,
  r_107__9_,r_107__8_,r_107__7_,r_107__6_,r_107__5_,r_107__4_,r_107__3_,r_107__2_,
  r_107__1_,r_107__0_,r_108__31_,r_108__30_,r_108__29_,r_108__28_,r_108__27_,
  r_108__26_,r_108__25_,r_108__24_,r_108__23_,r_108__22_,r_108__21_,r_108__20_,
  r_108__19_,r_108__18_,r_108__17_,r_108__16_,r_108__15_,r_108__14_,r_108__13_,r_108__12_,
  r_108__11_,r_108__10_,r_108__9_,r_108__8_,r_108__7_,r_108__6_,r_108__5_,r_108__4_,
  r_108__3_,r_108__2_,r_108__1_,r_108__0_,r_109__31_,r_109__30_,r_109__29_,
  r_109__28_,r_109__27_,r_109__26_,r_109__25_,r_109__24_,r_109__23_,r_109__22_,
  r_109__21_,r_109__20_,r_109__19_,r_109__18_,r_109__17_,r_109__16_,r_109__15_,r_109__14_,
  r_109__13_,r_109__12_,r_109__11_,r_109__10_,r_109__9_,r_109__8_,r_109__7_,
  r_109__6_,r_109__5_,r_109__4_,r_109__3_,r_109__2_,r_109__1_,r_109__0_,r_110__31_,
  r_110__30_,r_110__29_,r_110__28_,r_110__27_,r_110__26_,r_110__25_,r_110__24_,
  r_110__23_,r_110__22_,r_110__21_,r_110__20_,r_110__19_,r_110__18_,r_110__17_,r_110__16_,
  r_110__15_,r_110__14_,r_110__13_,r_110__12_,r_110__11_,r_110__10_,r_110__9_,
  r_110__8_,r_110__7_,r_110__6_,r_110__5_,r_110__4_,r_110__3_,r_110__2_,r_110__1_,
  r_110__0_,r_111__31_,r_111__30_,r_111__29_,r_111__28_,r_111__27_,r_111__26_,
  r_111__25_,r_111__24_,r_111__23_,r_111__22_,r_111__21_,r_111__20_,r_111__19_,r_111__18_,
  r_111__17_,r_111__16_,r_111__15_,r_111__14_,r_111__13_,r_111__12_,r_111__11_,
  r_111__10_,r_111__9_,r_111__8_,r_111__7_,r_111__6_,r_111__5_,r_111__4_,r_111__3_,
  r_111__2_,r_111__1_,r_111__0_,r_112__31_,r_112__30_,r_112__29_,r_112__28_,
  r_112__27_,r_112__26_,r_112__25_,r_112__24_,r_112__23_,r_112__22_,r_112__21_,r_112__20_,
  r_112__19_,r_112__18_,r_112__17_,r_112__16_,r_112__15_,r_112__14_,r_112__13_,
  r_112__12_,r_112__11_,r_112__10_,r_112__9_,r_112__8_,r_112__7_,r_112__6_,r_112__5_,
  r_112__4_,r_112__3_,r_112__2_,r_112__1_,r_112__0_,r_113__31_,r_113__30_,
  r_113__29_,r_113__28_,r_113__27_,r_113__26_,r_113__25_,r_113__24_,r_113__23_,r_113__22_,
  r_113__21_,r_113__20_,r_113__19_,r_113__18_,r_113__17_,r_113__16_,r_113__15_,
  r_113__14_,r_113__13_,r_113__12_,r_113__11_,r_113__10_,r_113__9_,r_113__8_,r_113__7_,
  r_113__6_,r_113__5_,r_113__4_,r_113__3_,r_113__2_,r_113__1_,r_113__0_,
  r_114__31_,r_114__30_,r_114__29_,r_114__28_,r_114__27_,r_114__26_,r_114__25_,r_114__24_,
  r_114__23_,r_114__22_,r_114__21_,r_114__20_,r_114__19_,r_114__18_,r_114__17_,
  r_114__16_,r_114__15_,r_114__14_,r_114__13_,r_114__12_,r_114__11_,r_114__10_,
  r_114__9_,r_114__8_,r_114__7_,r_114__6_,r_114__5_,r_114__4_,r_114__3_,r_114__2_,
  r_114__1_,r_114__0_,r_115__31_,r_115__30_,r_115__29_,r_115__28_,r_115__27_,r_115__26_,
  r_115__25_,r_115__24_,r_115__23_,r_115__22_,r_115__21_,r_115__20_,r_115__19_,
  r_115__18_,r_115__17_,r_115__16_,r_115__15_,r_115__14_,r_115__13_,r_115__12_,
  r_115__11_,r_115__10_,r_115__9_,r_115__8_,r_115__7_,r_115__6_,r_115__5_,r_115__4_,
  r_115__3_,r_115__2_,r_115__1_,r_115__0_,r_116__31_,r_116__30_,r_116__29_,r_116__28_,
  r_116__27_,r_116__26_,r_116__25_,r_116__24_,r_116__23_,r_116__22_,r_116__21_,
  r_116__20_,r_116__19_,r_116__18_,r_116__17_,r_116__16_,r_116__15_,r_116__14_,
  r_116__13_,r_116__12_,r_116__11_,r_116__10_,r_116__9_,r_116__8_,r_116__7_,r_116__6_,
  r_116__5_,r_116__4_,r_116__3_,r_116__2_,r_116__1_,r_116__0_,r_117__31_,r_117__30_,
  r_117__29_,r_117__28_,r_117__27_,r_117__26_,r_117__25_,r_117__24_,r_117__23_,
  r_117__22_,r_117__21_,r_117__20_,r_117__19_,r_117__18_,r_117__17_,r_117__16_,
  r_117__15_,r_117__14_,r_117__13_,r_117__12_,r_117__11_,r_117__10_,r_117__9_,r_117__8_,
  r_117__7_,r_117__6_,r_117__5_,r_117__4_,r_117__3_,r_117__2_,r_117__1_,r_117__0_,
  r_118__31_,r_118__30_,r_118__29_,r_118__28_,r_118__27_,r_118__26_,r_118__25_,
  r_118__24_,r_118__23_,r_118__22_,r_118__21_,r_118__20_,r_118__19_,r_118__18_,
  r_118__17_,r_118__16_,r_118__15_,r_118__14_,r_118__13_,r_118__12_,r_118__11_,r_118__10_,
  r_118__9_,r_118__8_,r_118__7_,r_118__6_,r_118__5_,r_118__4_,r_118__3_,r_118__2_,
  r_118__1_,r_118__0_,r_119__31_,r_119__30_,r_119__29_,r_119__28_,r_119__27_,
  r_119__26_,r_119__25_,r_119__24_,r_119__23_,r_119__22_,r_119__21_,r_119__20_,
  r_119__19_,r_119__18_,r_119__17_,r_119__16_,r_119__15_,r_119__14_,r_119__13_,r_119__12_,
  r_119__11_,r_119__10_,r_119__9_,r_119__8_,r_119__7_,r_119__6_,r_119__5_,
  r_119__4_,r_119__3_,r_119__2_,r_119__1_,r_119__0_,r_120__31_,r_120__30_,r_120__29_,
  r_120__28_,r_120__27_,r_120__26_,r_120__25_,r_120__24_,r_120__23_,r_120__22_,
  r_120__21_,r_120__20_,r_120__19_,r_120__18_,r_120__17_,r_120__16_,r_120__15_,r_120__14_,
  r_120__13_,r_120__12_,r_120__11_,r_120__10_,r_120__9_,r_120__8_,r_120__7_,
  r_120__6_,r_120__5_,r_120__4_,r_120__3_,r_120__2_,r_120__1_,r_120__0_,r_121__31_,
  r_121__30_,r_121__29_,r_121__28_,r_121__27_,r_121__26_,r_121__25_,r_121__24_,
  r_121__23_,r_121__22_,r_121__21_,r_121__20_,r_121__19_,r_121__18_,r_121__17_,r_121__16_,
  r_121__15_,r_121__14_,r_121__13_,r_121__12_,r_121__11_,r_121__10_,r_121__9_,
  r_121__8_,r_121__7_,r_121__6_,r_121__5_,r_121__4_,r_121__3_,r_121__2_,r_121__1_,
  r_121__0_,r_122__31_,r_122__30_,r_122__29_,r_122__28_,r_122__27_,r_122__26_,
  r_122__25_,r_122__24_,r_122__23_,r_122__22_,r_122__21_,r_122__20_,r_122__19_,r_122__18_,
  r_122__17_,r_122__16_,r_122__15_,r_122__14_,r_122__13_,r_122__12_,r_122__11_,
  r_122__10_,r_122__9_,r_122__8_,r_122__7_,r_122__6_,r_122__5_,r_122__4_,r_122__3_,
  r_122__2_,r_122__1_,r_122__0_,r_123__31_,r_123__30_,r_123__29_,r_123__28_,
  r_123__27_,r_123__26_,r_123__25_,r_123__24_,r_123__23_,r_123__22_,r_123__21_,r_123__20_,
  r_123__19_,r_123__18_,r_123__17_,r_123__16_,r_123__15_,r_123__14_,r_123__13_,
  r_123__12_,r_123__11_,r_123__10_,r_123__9_,r_123__8_,r_123__7_,r_123__6_,r_123__5_,
  r_123__4_,r_123__3_,r_123__2_,r_123__1_,r_123__0_,r_124__31_,r_124__30_,
  r_124__29_,r_124__28_,r_124__27_,r_124__26_,r_124__25_,r_124__24_,r_124__23_,r_124__22_,
  r_124__21_,r_124__20_,r_124__19_,r_124__18_,r_124__17_,r_124__16_,r_124__15_,
  r_124__14_,r_124__13_,r_124__12_,r_124__11_,r_124__10_,r_124__9_,r_124__8_,
  r_124__7_,r_124__6_,r_124__5_,r_124__4_,r_124__3_,r_124__2_,r_124__1_,r_124__0_,
  r_125__31_,r_125__30_,r_125__29_,r_125__28_,r_125__27_,r_125__26_,r_125__25_,r_125__24_,
  r_125__23_,r_125__22_,r_125__21_,r_125__20_,r_125__19_,r_125__18_,r_125__17_,
  r_125__16_,r_125__15_,r_125__14_,r_125__13_,r_125__12_,r_125__11_,r_125__10_,
  r_125__9_,r_125__8_,r_125__7_,r_125__6_,r_125__5_,r_125__4_,r_125__3_,r_125__2_,
  r_125__1_,r_125__0_,r_126__31_,r_126__30_,r_126__29_,r_126__28_,r_126__27_,r_126__26_,
  r_126__25_,r_126__24_,r_126__23_,r_126__22_,r_126__21_,r_126__20_,r_126__19_,
  r_126__18_,r_126__17_,r_126__16_,r_126__15_,r_126__14_,r_126__13_,r_126__12_,
  r_126__11_,r_126__10_,r_126__9_,r_126__8_,r_126__7_,r_126__6_,r_126__5_,r_126__4_,
  r_126__3_,r_126__2_,r_126__1_,r_126__0_,r_127__31_,r_127__30_,r_127__29_,r_127__28_,
  r_127__27_,r_127__26_,r_127__25_,r_127__24_,r_127__23_,r_127__22_,r_127__21_,
  r_127__20_,r_127__19_,r_127__18_,r_127__17_,r_127__16_,r_127__15_,r_127__14_,
  r_127__13_,r_127__12_,r_127__11_,r_127__10_,r_127__9_,r_127__8_,r_127__7_,r_127__6_,
  r_127__5_,r_127__4_,r_127__3_,r_127__2_,r_127__1_,r_127__0_,r_128__31_,r_128__30_,
  r_128__29_,r_128__28_,r_128__27_,r_128__26_,r_128__25_,r_128__24_,r_128__23_,
  r_128__22_,r_128__21_,r_128__20_,r_128__19_,r_128__18_,r_128__17_,r_128__16_,
  r_128__15_,r_128__14_,r_128__13_,r_128__12_,r_128__11_,r_128__10_,r_128__9_,r_128__8_,
  r_128__7_,r_128__6_,r_128__5_,r_128__4_,r_128__3_,r_128__2_,r_128__1_,r_128__0_,
  r_129__31_,r_129__30_,r_129__29_,r_129__28_,r_129__27_,r_129__26_,r_129__25_,
  r_129__24_,r_129__23_,r_129__22_,r_129__21_,r_129__20_,r_129__19_,r_129__18_,
  r_129__17_,r_129__16_,r_129__15_,r_129__14_,r_129__13_,r_129__12_,r_129__11_,
  r_129__10_,r_129__9_,r_129__8_,r_129__7_,r_129__6_,r_129__5_,r_129__4_,r_129__3_,
  r_129__2_,r_129__1_,r_129__0_,r_130__31_,r_130__30_,r_130__29_,r_130__28_,r_130__27_,
  r_130__26_,r_130__25_,r_130__24_,r_130__23_,r_130__22_,r_130__21_,r_130__20_,
  r_130__19_,r_130__18_,r_130__17_,r_130__16_,r_130__15_,r_130__14_,r_130__13_,
  r_130__12_,r_130__11_,r_130__10_,r_130__9_,r_130__8_,r_130__7_,r_130__6_,r_130__5_,
  r_130__4_,r_130__3_,r_130__2_,r_130__1_,r_130__0_,r_131__31_,r_131__30_,r_131__29_,
  r_131__28_,r_131__27_,r_131__26_,r_131__25_,r_131__24_,r_131__23_,r_131__22_,
  r_131__21_,r_131__20_,r_131__19_,r_131__18_,r_131__17_,r_131__16_,r_131__15_,
  r_131__14_,r_131__13_,r_131__12_,r_131__11_,r_131__10_,r_131__9_,r_131__8_,r_131__7_,
  r_131__6_,r_131__5_,r_131__4_,r_131__3_,r_131__2_,r_131__1_,r_131__0_,r_132__31_,
  r_132__30_,r_132__29_,r_132__28_,r_132__27_,r_132__26_,r_132__25_,r_132__24_,
  r_132__23_,r_132__22_,r_132__21_,r_132__20_,r_132__19_,r_132__18_,r_132__17_,
  r_132__16_,r_132__15_,r_132__14_,r_132__13_,r_132__12_,r_132__11_,r_132__10_,r_132__9_,
  r_132__8_,r_132__7_,r_132__6_,r_132__5_,r_132__4_,r_132__3_,r_132__2_,r_132__1_,
  r_132__0_,r_133__31_,r_133__30_,r_133__29_,r_133__28_,r_133__27_,r_133__26_,
  r_133__25_,r_133__24_,r_133__23_,r_133__22_,r_133__21_,r_133__20_,r_133__19_,
  r_133__18_,r_133__17_,r_133__16_,r_133__15_,r_133__14_,r_133__13_,r_133__12_,r_133__11_,
  r_133__10_,r_133__9_,r_133__8_,r_133__7_,r_133__6_,r_133__5_,r_133__4_,r_133__3_,
  r_133__2_,r_133__1_,r_133__0_,r_134__31_,r_134__30_,r_134__29_,r_134__28_,
  r_134__27_,r_134__26_,r_134__25_,r_134__24_,r_134__23_,r_134__22_,r_134__21_,
  r_134__20_,r_134__19_,r_134__18_,r_134__17_,r_134__16_,r_134__15_,r_134__14_,r_134__13_,
  r_134__12_,r_134__11_,r_134__10_,r_134__9_,r_134__8_,r_134__7_,r_134__6_,
  r_134__5_,r_134__4_,r_134__3_,r_134__2_,r_134__1_,r_134__0_,r_135__31_,r_135__30_,
  r_135__29_,r_135__28_,r_135__27_,r_135__26_,r_135__25_,r_135__24_,r_135__23_,
  r_135__22_,r_135__21_,r_135__20_,r_135__19_,r_135__18_,r_135__17_,r_135__16_,r_135__15_,
  r_135__14_,r_135__13_,r_135__12_,r_135__11_,r_135__10_,r_135__9_,r_135__8_,
  r_135__7_,r_135__6_,r_135__5_,r_135__4_,r_135__3_,r_135__2_,r_135__1_,r_135__0_,
  r_136__31_,r_136__30_,r_136__29_,r_136__28_,r_136__27_,r_136__26_,r_136__25_,
  r_136__24_,r_136__23_,r_136__22_,r_136__21_,r_136__20_,r_136__19_,r_136__18_,r_136__17_,
  r_136__16_,r_136__15_,r_136__14_,r_136__13_,r_136__12_,r_136__11_,r_136__10_,
  r_136__9_,r_136__8_,r_136__7_,r_136__6_,r_136__5_,r_136__4_,r_136__3_,r_136__2_,
  r_136__1_,r_136__0_,r_137__31_,r_137__30_,r_137__29_,r_137__28_,r_137__27_,
  r_137__26_,r_137__25_,r_137__24_,r_137__23_,r_137__22_,r_137__21_,r_137__20_,r_137__19_,
  r_137__18_,r_137__17_,r_137__16_,r_137__15_,r_137__14_,r_137__13_,r_137__12_,
  r_137__11_,r_137__10_,r_137__9_,r_137__8_,r_137__7_,r_137__6_,r_137__5_,r_137__4_,
  r_137__3_,r_137__2_,r_137__1_,r_137__0_,r_138__31_,r_138__30_,r_138__29_,
  r_138__28_,r_138__27_,r_138__26_,r_138__25_,r_138__24_,r_138__23_,r_138__22_,r_138__21_,
  r_138__20_,r_138__19_,r_138__18_,r_138__17_,r_138__16_,r_138__15_,r_138__14_,
  r_138__13_,r_138__12_,r_138__11_,r_138__10_,r_138__9_,r_138__8_,r_138__7_,r_138__6_,
  r_138__5_,r_138__4_,r_138__3_,r_138__2_,r_138__1_,r_138__0_,r_139__31_,
  r_139__30_,r_139__29_,r_139__28_,r_139__27_,r_139__26_,r_139__25_,r_139__24_,r_139__23_,
  r_139__22_,r_139__21_,r_139__20_,r_139__19_,r_139__18_,r_139__17_,r_139__16_,
  r_139__15_,r_139__14_,r_139__13_,r_139__12_,r_139__11_,r_139__10_,r_139__9_,
  r_139__8_,r_139__7_,r_139__6_,r_139__5_,r_139__4_,r_139__3_,r_139__2_,r_139__1_,
  r_139__0_,r_140__31_,r_140__30_,r_140__29_,r_140__28_,r_140__27_,r_140__26_,r_140__25_,
  r_140__24_,r_140__23_,r_140__22_,r_140__21_,r_140__20_,r_140__19_,r_140__18_,
  r_140__17_,r_140__16_,r_140__15_,r_140__14_,r_140__13_,r_140__12_,r_140__11_,
  r_140__10_,r_140__9_,r_140__8_,r_140__7_,r_140__6_,r_140__5_,r_140__4_,r_140__3_,
  r_140__2_,r_140__1_,r_140__0_,r_141__31_,r_141__30_,r_141__29_,r_141__28_,r_141__27_,
  r_141__26_,r_141__25_,r_141__24_,r_141__23_,r_141__22_,r_141__21_,r_141__20_,
  r_141__19_,r_141__18_,r_141__17_,r_141__16_,r_141__15_,r_141__14_,r_141__13_,
  r_141__12_,r_141__11_,r_141__10_,r_141__9_,r_141__8_,r_141__7_,r_141__6_,r_141__5_,
  r_141__4_,r_141__3_,r_141__2_,r_141__1_,r_141__0_,r_142__31_,r_142__30_,r_142__29_,
  r_142__28_,r_142__27_,r_142__26_,r_142__25_,r_142__24_,r_142__23_,r_142__22_,
  r_142__21_,r_142__20_,r_142__19_,r_142__18_,r_142__17_,r_142__16_,r_142__15_,
  r_142__14_,r_142__13_,r_142__12_,r_142__11_,r_142__10_,r_142__9_,r_142__8_,r_142__7_,
  r_142__6_,r_142__5_,r_142__4_,r_142__3_,r_142__2_,r_142__1_,r_142__0_,r_143__31_,
  r_143__30_,r_143__29_,r_143__28_,r_143__27_,r_143__26_,r_143__25_,r_143__24_,
  r_143__23_,r_143__22_,r_143__21_,r_143__20_,r_143__19_,r_143__18_,r_143__17_,
  r_143__16_,r_143__15_,r_143__14_,r_143__13_,r_143__12_,r_143__11_,r_143__10_,r_143__9_,
  r_143__8_,r_143__7_,r_143__6_,r_143__5_,r_143__4_,r_143__3_,r_143__2_,r_143__1_,
  r_143__0_,r_144__31_,r_144__30_,r_144__29_,r_144__28_,r_144__27_,r_144__26_,
  r_144__25_,r_144__24_,r_144__23_,r_144__22_,r_144__21_,r_144__20_,r_144__19_,
  r_144__18_,r_144__17_,r_144__16_,r_144__15_,r_144__14_,r_144__13_,r_144__12_,
  r_144__11_,r_144__10_,r_144__9_,r_144__8_,r_144__7_,r_144__6_,r_144__5_,r_144__4_,
  r_144__3_,r_144__2_,r_144__1_,r_144__0_,r_145__31_,r_145__30_,r_145__29_,r_145__28_,
  r_145__27_,r_145__26_,r_145__25_,r_145__24_,r_145__23_,r_145__22_,r_145__21_,
  r_145__20_,r_145__19_,r_145__18_,r_145__17_,r_145__16_,r_145__15_,r_145__14_,
  r_145__13_,r_145__12_,r_145__11_,r_145__10_,r_145__9_,r_145__8_,r_145__7_,r_145__6_,
  r_145__5_,r_145__4_,r_145__3_,r_145__2_,r_145__1_,r_145__0_,r_146__31_,r_146__30_,
  r_146__29_,r_146__28_,r_146__27_,r_146__26_,r_146__25_,r_146__24_,r_146__23_,
  r_146__22_,r_146__21_,r_146__20_,r_146__19_,r_146__18_,r_146__17_,r_146__16_,
  r_146__15_,r_146__14_,r_146__13_,r_146__12_,r_146__11_,r_146__10_,r_146__9_,r_146__8_,
  r_146__7_,r_146__6_,r_146__5_,r_146__4_,r_146__3_,r_146__2_,r_146__1_,r_146__0_,
  r_147__31_,r_147__30_,r_147__29_,r_147__28_,r_147__27_,r_147__26_,r_147__25_,
  r_147__24_,r_147__23_,r_147__22_,r_147__21_,r_147__20_,r_147__19_,r_147__18_,
  r_147__17_,r_147__16_,r_147__15_,r_147__14_,r_147__13_,r_147__12_,r_147__11_,r_147__10_,
  r_147__9_,r_147__8_,r_147__7_,r_147__6_,r_147__5_,r_147__4_,r_147__3_,r_147__2_,
  r_147__1_,r_147__0_,r_148__31_,r_148__30_,r_148__29_,r_148__28_,r_148__27_,
  r_148__26_,r_148__25_,r_148__24_,r_148__23_,r_148__22_,r_148__21_,r_148__20_,
  r_148__19_,r_148__18_,r_148__17_,r_148__16_,r_148__15_,r_148__14_,r_148__13_,r_148__12_,
  r_148__11_,r_148__10_,r_148__9_,r_148__8_,r_148__7_,r_148__6_,r_148__5_,r_148__4_,
  r_148__3_,r_148__2_,r_148__1_,r_148__0_,r_149__31_,r_149__30_,r_149__29_,
  r_149__28_,r_149__27_,r_149__26_,r_149__25_,r_149__24_,r_149__23_,r_149__22_,
  r_149__21_,r_149__20_,r_149__19_,r_149__18_,r_149__17_,r_149__16_,r_149__15_,r_149__14_,
  r_149__13_,r_149__12_,r_149__11_,r_149__10_,r_149__9_,r_149__8_,r_149__7_,
  r_149__6_,r_149__5_,r_149__4_,r_149__3_,r_149__2_,r_149__1_,r_149__0_,r_150__31_,
  r_150__30_,r_150__29_,r_150__28_,r_150__27_,r_150__26_,r_150__25_,r_150__24_,
  r_150__23_,r_150__22_,r_150__21_,r_150__20_,r_150__19_,r_150__18_,r_150__17_,r_150__16_,
  r_150__15_,r_150__14_,r_150__13_,r_150__12_,r_150__11_,r_150__10_,r_150__9_,
  r_150__8_,r_150__7_,r_150__6_,r_150__5_,r_150__4_,r_150__3_,r_150__2_,r_150__1_,
  r_150__0_,r_151__31_,r_151__30_,r_151__29_,r_151__28_,r_151__27_,r_151__26_,
  r_151__25_,r_151__24_,r_151__23_,r_151__22_,r_151__21_,r_151__20_,r_151__19_,r_151__18_,
  r_151__17_,r_151__16_,r_151__15_,r_151__14_,r_151__13_,r_151__12_,r_151__11_,
  r_151__10_,r_151__9_,r_151__8_,r_151__7_,r_151__6_,r_151__5_,r_151__4_,r_151__3_,
  r_151__2_,r_151__1_,r_151__0_,r_152__31_,r_152__30_,r_152__29_,r_152__28_,
  r_152__27_,r_152__26_,r_152__25_,r_152__24_,r_152__23_,r_152__22_,r_152__21_,r_152__20_,
  r_152__19_,r_152__18_,r_152__17_,r_152__16_,r_152__15_,r_152__14_,r_152__13_,
  r_152__12_,r_152__11_,r_152__10_,r_152__9_,r_152__8_,r_152__7_,r_152__6_,r_152__5_,
  r_152__4_,r_152__3_,r_152__2_,r_152__1_,r_152__0_,r_153__31_,r_153__30_,
  r_153__29_,r_153__28_,r_153__27_,r_153__26_,r_153__25_,r_153__24_,r_153__23_,r_153__22_,
  r_153__21_,r_153__20_,r_153__19_,r_153__18_,r_153__17_,r_153__16_,r_153__15_,
  r_153__14_,r_153__13_,r_153__12_,r_153__11_,r_153__10_,r_153__9_,r_153__8_,r_153__7_,
  r_153__6_,r_153__5_,r_153__4_,r_153__3_,r_153__2_,r_153__1_,r_153__0_,
  r_154__31_,r_154__30_,r_154__29_,r_154__28_,r_154__27_,r_154__26_,r_154__25_,r_154__24_,
  r_154__23_,r_154__22_,r_154__21_,r_154__20_,r_154__19_,r_154__18_,r_154__17_,
  r_154__16_,r_154__15_,r_154__14_,r_154__13_,r_154__12_,r_154__11_,r_154__10_,
  r_154__9_,r_154__8_,r_154__7_,r_154__6_,r_154__5_,r_154__4_,r_154__3_,r_154__2_,
  r_154__1_,r_154__0_,r_155__31_,r_155__30_,r_155__29_,r_155__28_,r_155__27_,r_155__26_,
  r_155__25_,r_155__24_,r_155__23_,r_155__22_,r_155__21_,r_155__20_,r_155__19_,
  r_155__18_,r_155__17_,r_155__16_,r_155__15_,r_155__14_,r_155__13_,r_155__12_,
  r_155__11_,r_155__10_,r_155__9_,r_155__8_,r_155__7_,r_155__6_,r_155__5_,r_155__4_,
  r_155__3_,r_155__2_,r_155__1_,r_155__0_,r_156__31_,r_156__30_,r_156__29_,r_156__28_,
  r_156__27_,r_156__26_,r_156__25_,r_156__24_,r_156__23_,r_156__22_,r_156__21_,
  r_156__20_,r_156__19_,r_156__18_,r_156__17_,r_156__16_,r_156__15_,r_156__14_,
  r_156__13_,r_156__12_,r_156__11_,r_156__10_,r_156__9_,r_156__8_,r_156__7_,r_156__6_,
  r_156__5_,r_156__4_,r_156__3_,r_156__2_,r_156__1_,r_156__0_,r_157__31_,r_157__30_,
  r_157__29_,r_157__28_,r_157__27_,r_157__26_,r_157__25_,r_157__24_,r_157__23_,
  r_157__22_,r_157__21_,r_157__20_,r_157__19_,r_157__18_,r_157__17_,r_157__16_,
  r_157__15_,r_157__14_,r_157__13_,r_157__12_,r_157__11_,r_157__10_,r_157__9_,r_157__8_,
  r_157__7_,r_157__6_,r_157__5_,r_157__4_,r_157__3_,r_157__2_,r_157__1_,r_157__0_,
  r_158__31_,r_158__30_,r_158__29_,r_158__28_,r_158__27_,r_158__26_,r_158__25_,
  r_158__24_,r_158__23_,r_158__22_,r_158__21_,r_158__20_,r_158__19_,r_158__18_,
  r_158__17_,r_158__16_,r_158__15_,r_158__14_,r_158__13_,r_158__12_,r_158__11_,r_158__10_,
  r_158__9_,r_158__8_,r_158__7_,r_158__6_,r_158__5_,r_158__4_,r_158__3_,r_158__2_,
  r_158__1_,r_158__0_,r_159__31_,r_159__30_,r_159__29_,r_159__28_,r_159__27_,
  r_159__26_,r_159__25_,r_159__24_,r_159__23_,r_159__22_,r_159__21_,r_159__20_,
  r_159__19_,r_159__18_,r_159__17_,r_159__16_,r_159__15_,r_159__14_,r_159__13_,r_159__12_,
  r_159__11_,r_159__10_,r_159__9_,r_159__8_,r_159__7_,r_159__6_,r_159__5_,
  r_159__4_,r_159__3_,r_159__2_,r_159__1_,r_159__0_,r_160__31_,r_160__30_,r_160__29_,
  r_160__28_,r_160__27_,r_160__26_,r_160__25_,r_160__24_,r_160__23_,r_160__22_,
  r_160__21_,r_160__20_,r_160__19_,r_160__18_,r_160__17_,r_160__16_,r_160__15_,r_160__14_,
  r_160__13_,r_160__12_,r_160__11_,r_160__10_,r_160__9_,r_160__8_,r_160__7_,
  r_160__6_,r_160__5_,r_160__4_,r_160__3_,r_160__2_,r_160__1_,r_160__0_,r_161__31_,
  r_161__30_,r_161__29_,r_161__28_,r_161__27_,r_161__26_,r_161__25_,r_161__24_,
  r_161__23_,r_161__22_,r_161__21_,r_161__20_,r_161__19_,r_161__18_,r_161__17_,r_161__16_,
  r_161__15_,r_161__14_,r_161__13_,r_161__12_,r_161__11_,r_161__10_,r_161__9_,
  r_161__8_,r_161__7_,r_161__6_,r_161__5_,r_161__4_,r_161__3_,r_161__2_,r_161__1_,
  r_161__0_,r_162__31_,r_162__30_,r_162__29_,r_162__28_,r_162__27_,r_162__26_,
  r_162__25_,r_162__24_,r_162__23_,r_162__22_,r_162__21_,r_162__20_,r_162__19_,r_162__18_,
  r_162__17_,r_162__16_,r_162__15_,r_162__14_,r_162__13_,r_162__12_,r_162__11_,
  r_162__10_,r_162__9_,r_162__8_,r_162__7_,r_162__6_,r_162__5_,r_162__4_,r_162__3_,
  r_162__2_,r_162__1_,r_162__0_,r_163__31_,r_163__30_,r_163__29_,r_163__28_,
  r_163__27_,r_163__26_,r_163__25_,r_163__24_,r_163__23_,r_163__22_,r_163__21_,r_163__20_,
  r_163__19_,r_163__18_,r_163__17_,r_163__16_,r_163__15_,r_163__14_,r_163__13_,
  r_163__12_,r_163__11_,r_163__10_,r_163__9_,r_163__8_,r_163__7_,r_163__6_,r_163__5_,
  r_163__4_,r_163__3_,r_163__2_,r_163__1_,r_163__0_,r_164__31_,r_164__30_,
  r_164__29_,r_164__28_,r_164__27_,r_164__26_,r_164__25_,r_164__24_,r_164__23_,r_164__22_,
  r_164__21_,r_164__20_,r_164__19_,r_164__18_,r_164__17_,r_164__16_,r_164__15_,
  r_164__14_,r_164__13_,r_164__12_,r_164__11_,r_164__10_,r_164__9_,r_164__8_,
  r_164__7_,r_164__6_,r_164__5_,r_164__4_,r_164__3_,r_164__2_,r_164__1_,r_164__0_,
  r_165__31_,r_165__30_,r_165__29_,r_165__28_,r_165__27_,r_165__26_,r_165__25_,r_165__24_,
  r_165__23_,r_165__22_,r_165__21_,r_165__20_,r_165__19_,r_165__18_,r_165__17_,
  r_165__16_,r_165__15_,r_165__14_,r_165__13_,r_165__12_,r_165__11_,r_165__10_,
  r_165__9_,r_165__8_,r_165__7_,r_165__6_,r_165__5_,r_165__4_,r_165__3_,r_165__2_,
  r_165__1_,r_165__0_,r_166__31_,r_166__30_,r_166__29_,r_166__28_,r_166__27_,r_166__26_,
  r_166__25_,r_166__24_,r_166__23_,r_166__22_,r_166__21_,r_166__20_,r_166__19_,
  r_166__18_,r_166__17_,r_166__16_,r_166__15_,r_166__14_,r_166__13_,r_166__12_,
  r_166__11_,r_166__10_,r_166__9_,r_166__8_,r_166__7_,r_166__6_,r_166__5_,r_166__4_,
  r_166__3_,r_166__2_,r_166__1_,r_166__0_,r_167__31_,r_167__30_,r_167__29_,r_167__28_,
  r_167__27_,r_167__26_,r_167__25_,r_167__24_,r_167__23_,r_167__22_,r_167__21_,
  r_167__20_,r_167__19_,r_167__18_,r_167__17_,r_167__16_,r_167__15_,r_167__14_,
  r_167__13_,r_167__12_,r_167__11_,r_167__10_,r_167__9_,r_167__8_,r_167__7_,r_167__6_,
  r_167__5_,r_167__4_,r_167__3_,r_167__2_,r_167__1_,r_167__0_,r_168__31_,r_168__30_,
  r_168__29_,r_168__28_,r_168__27_,r_168__26_,r_168__25_,r_168__24_,r_168__23_,
  r_168__22_,r_168__21_,r_168__20_,r_168__19_,r_168__18_,r_168__17_,r_168__16_,
  r_168__15_,r_168__14_,r_168__13_,r_168__12_,r_168__11_,r_168__10_,r_168__9_,r_168__8_,
  r_168__7_,r_168__6_,r_168__5_,r_168__4_,r_168__3_,r_168__2_,r_168__1_,r_168__0_,
  r_169__31_,r_169__30_,r_169__29_,r_169__28_,r_169__27_,r_169__26_,r_169__25_,
  r_169__24_,r_169__23_,r_169__22_,r_169__21_,r_169__20_,r_169__19_,r_169__18_,
  r_169__17_,r_169__16_,r_169__15_,r_169__14_,r_169__13_,r_169__12_,r_169__11_,
  r_169__10_,r_169__9_,r_169__8_,r_169__7_,r_169__6_,r_169__5_,r_169__4_,r_169__3_,
  r_169__2_,r_169__1_,r_169__0_,r_170__31_,r_170__30_,r_170__29_,r_170__28_,r_170__27_,
  r_170__26_,r_170__25_,r_170__24_,r_170__23_,r_170__22_,r_170__21_,r_170__20_,
  r_170__19_,r_170__18_,r_170__17_,r_170__16_,r_170__15_,r_170__14_,r_170__13_,
  r_170__12_,r_170__11_,r_170__10_,r_170__9_,r_170__8_,r_170__7_,r_170__6_,r_170__5_,
  r_170__4_,r_170__3_,r_170__2_,r_170__1_,r_170__0_,r_171__31_,r_171__30_,r_171__29_,
  r_171__28_,r_171__27_,r_171__26_,r_171__25_,r_171__24_,r_171__23_,r_171__22_,
  r_171__21_,r_171__20_,r_171__19_,r_171__18_,r_171__17_,r_171__16_,r_171__15_,
  r_171__14_,r_171__13_,r_171__12_,r_171__11_,r_171__10_,r_171__9_,r_171__8_,r_171__7_,
  r_171__6_,r_171__5_,r_171__4_,r_171__3_,r_171__2_,r_171__1_,r_171__0_,r_172__31_,
  r_172__30_,r_172__29_,r_172__28_,r_172__27_,r_172__26_,r_172__25_,r_172__24_,
  r_172__23_,r_172__22_,r_172__21_,r_172__20_,r_172__19_,r_172__18_,r_172__17_,
  r_172__16_,r_172__15_,r_172__14_,r_172__13_,r_172__12_,r_172__11_,r_172__10_,r_172__9_,
  r_172__8_,r_172__7_,r_172__6_,r_172__5_,r_172__4_,r_172__3_,r_172__2_,r_172__1_,
  r_172__0_,r_173__31_,r_173__30_,r_173__29_,r_173__28_,r_173__27_,r_173__26_,
  r_173__25_,r_173__24_,r_173__23_,r_173__22_,r_173__21_,r_173__20_,r_173__19_,
  r_173__18_,r_173__17_,r_173__16_,r_173__15_,r_173__14_,r_173__13_,r_173__12_,r_173__11_,
  r_173__10_,r_173__9_,r_173__8_,r_173__7_,r_173__6_,r_173__5_,r_173__4_,r_173__3_,
  r_173__2_,r_173__1_,r_173__0_,r_174__31_,r_174__30_,r_174__29_,r_174__28_,
  r_174__27_,r_174__26_,r_174__25_,r_174__24_,r_174__23_,r_174__22_,r_174__21_,
  r_174__20_,r_174__19_,r_174__18_,r_174__17_,r_174__16_,r_174__15_,r_174__14_,r_174__13_,
  r_174__12_,r_174__11_,r_174__10_,r_174__9_,r_174__8_,r_174__7_,r_174__6_,
  r_174__5_,r_174__4_,r_174__3_,r_174__2_,r_174__1_,r_174__0_,r_175__31_,r_175__30_,
  r_175__29_,r_175__28_,r_175__27_,r_175__26_,r_175__25_,r_175__24_,r_175__23_,
  r_175__22_,r_175__21_,r_175__20_,r_175__19_,r_175__18_,r_175__17_,r_175__16_,r_175__15_,
  r_175__14_,r_175__13_,r_175__12_,r_175__11_,r_175__10_,r_175__9_,r_175__8_,
  r_175__7_,r_175__6_,r_175__5_,r_175__4_,r_175__3_,r_175__2_,r_175__1_,r_175__0_,
  r_176__31_,r_176__30_,r_176__29_,r_176__28_,r_176__27_,r_176__26_,r_176__25_,
  r_176__24_,r_176__23_,r_176__22_,r_176__21_,r_176__20_,r_176__19_,r_176__18_,r_176__17_,
  r_176__16_,r_176__15_,r_176__14_,r_176__13_,r_176__12_,r_176__11_,r_176__10_,
  r_176__9_,r_176__8_,r_176__7_,r_176__6_,r_176__5_,r_176__4_,r_176__3_,r_176__2_,
  r_176__1_,r_176__0_,r_177__31_,r_177__30_,r_177__29_,r_177__28_,r_177__27_,
  r_177__26_,r_177__25_,r_177__24_,r_177__23_,r_177__22_,r_177__21_,r_177__20_,r_177__19_,
  r_177__18_,r_177__17_,r_177__16_,r_177__15_,r_177__14_,r_177__13_,r_177__12_,
  r_177__11_,r_177__10_,r_177__9_,r_177__8_,r_177__7_,r_177__6_,r_177__5_,r_177__4_,
  r_177__3_,r_177__2_,r_177__1_,r_177__0_,r_178__31_,r_178__30_,r_178__29_,
  r_178__28_,r_178__27_,r_178__26_,r_178__25_,r_178__24_,r_178__23_,r_178__22_,r_178__21_,
  r_178__20_,r_178__19_,r_178__18_,r_178__17_,r_178__16_,r_178__15_,r_178__14_,
  r_178__13_,r_178__12_,r_178__11_,r_178__10_,r_178__9_,r_178__8_,r_178__7_,r_178__6_,
  r_178__5_,r_178__4_,r_178__3_,r_178__2_,r_178__1_,r_178__0_,r_179__31_,
  r_179__30_,r_179__29_,r_179__28_,r_179__27_,r_179__26_,r_179__25_,r_179__24_,r_179__23_,
  r_179__22_,r_179__21_,r_179__20_,r_179__19_,r_179__18_,r_179__17_,r_179__16_,
  r_179__15_,r_179__14_,r_179__13_,r_179__12_,r_179__11_,r_179__10_,r_179__9_,
  r_179__8_,r_179__7_,r_179__6_,r_179__5_,r_179__4_,r_179__3_,r_179__2_,r_179__1_,
  r_179__0_,r_180__31_,r_180__30_,r_180__29_,r_180__28_,r_180__27_,r_180__26_,r_180__25_,
  r_180__24_,r_180__23_,r_180__22_,r_180__21_,r_180__20_,r_180__19_,r_180__18_,
  r_180__17_,r_180__16_,r_180__15_,r_180__14_,r_180__13_,r_180__12_,r_180__11_,
  r_180__10_,r_180__9_,r_180__8_,r_180__7_,r_180__6_,r_180__5_,r_180__4_,r_180__3_,
  r_180__2_,r_180__1_,r_180__0_,r_181__31_,r_181__30_,r_181__29_,r_181__28_,r_181__27_,
  r_181__26_,r_181__25_,r_181__24_,r_181__23_,r_181__22_,r_181__21_,r_181__20_,
  r_181__19_,r_181__18_,r_181__17_,r_181__16_,r_181__15_,r_181__14_,r_181__13_,
  r_181__12_,r_181__11_,r_181__10_,r_181__9_,r_181__8_,r_181__7_,r_181__6_,r_181__5_,
  r_181__4_,r_181__3_,r_181__2_,r_181__1_,r_181__0_,r_182__31_,r_182__30_,r_182__29_,
  r_182__28_,r_182__27_,r_182__26_,r_182__25_,r_182__24_,r_182__23_,r_182__22_,
  r_182__21_,r_182__20_,r_182__19_,r_182__18_,r_182__17_,r_182__16_,r_182__15_,
  r_182__14_,r_182__13_,r_182__12_,r_182__11_,r_182__10_,r_182__9_,r_182__8_,r_182__7_,
  r_182__6_,r_182__5_,r_182__4_,r_182__3_,r_182__2_,r_182__1_,r_182__0_,r_183__31_,
  r_183__30_,r_183__29_,r_183__28_,r_183__27_,r_183__26_,r_183__25_,r_183__24_,
  r_183__23_,r_183__22_,r_183__21_,r_183__20_,r_183__19_,r_183__18_,r_183__17_,
  r_183__16_,r_183__15_,r_183__14_,r_183__13_,r_183__12_,r_183__11_,r_183__10_,r_183__9_,
  r_183__8_,r_183__7_,r_183__6_,r_183__5_,r_183__4_,r_183__3_,r_183__2_,r_183__1_,
  r_183__0_,r_184__31_,r_184__30_,r_184__29_,r_184__28_,r_184__27_,r_184__26_,
  r_184__25_,r_184__24_,r_184__23_,r_184__22_,r_184__21_,r_184__20_,r_184__19_,
  r_184__18_,r_184__17_,r_184__16_,r_184__15_,r_184__14_,r_184__13_,r_184__12_,
  r_184__11_,r_184__10_,r_184__9_,r_184__8_,r_184__7_,r_184__6_,r_184__5_,r_184__4_,
  r_184__3_,r_184__2_,r_184__1_,r_184__0_,r_185__31_,r_185__30_,r_185__29_,r_185__28_,
  r_185__27_,r_185__26_,r_185__25_,r_185__24_,r_185__23_,r_185__22_,r_185__21_,
  r_185__20_,r_185__19_,r_185__18_,r_185__17_,r_185__16_,r_185__15_,r_185__14_,
  r_185__13_,r_185__12_,r_185__11_,r_185__10_,r_185__9_,r_185__8_,r_185__7_,r_185__6_,
  r_185__5_,r_185__4_,r_185__3_,r_185__2_,r_185__1_,r_185__0_,r_186__31_,r_186__30_,
  r_186__29_,r_186__28_,r_186__27_,r_186__26_,r_186__25_,r_186__24_,r_186__23_,
  r_186__22_,r_186__21_,r_186__20_,r_186__19_,r_186__18_,r_186__17_,r_186__16_,
  r_186__15_,r_186__14_,r_186__13_,r_186__12_,r_186__11_,r_186__10_,r_186__9_,r_186__8_,
  r_186__7_,r_186__6_,r_186__5_,r_186__4_,r_186__3_,r_186__2_,r_186__1_,r_186__0_,
  r_187__31_,r_187__30_,r_187__29_,r_187__28_,r_187__27_,r_187__26_,r_187__25_,
  r_187__24_,r_187__23_,r_187__22_,r_187__21_,r_187__20_,r_187__19_,r_187__18_,
  r_187__17_,r_187__16_,r_187__15_,r_187__14_,r_187__13_,r_187__12_,r_187__11_,r_187__10_,
  r_187__9_,r_187__8_,r_187__7_,r_187__6_,r_187__5_,r_187__4_,r_187__3_,r_187__2_,
  r_187__1_,r_187__0_,r_188__31_,r_188__30_,r_188__29_,r_188__28_,r_188__27_,
  r_188__26_,r_188__25_,r_188__24_,r_188__23_,r_188__22_,r_188__21_,r_188__20_,
  r_188__19_,r_188__18_,r_188__17_,r_188__16_,r_188__15_,r_188__14_,r_188__13_,r_188__12_,
  r_188__11_,r_188__10_,r_188__9_,r_188__8_,r_188__7_,r_188__6_,r_188__5_,r_188__4_,
  r_188__3_,r_188__2_,r_188__1_,r_188__0_,r_189__31_,r_189__30_,r_189__29_,
  r_189__28_,r_189__27_,r_189__26_,r_189__25_,r_189__24_,r_189__23_,r_189__22_,
  r_189__21_,r_189__20_,r_189__19_,r_189__18_,r_189__17_,r_189__16_,r_189__15_,r_189__14_,
  r_189__13_,r_189__12_,r_189__11_,r_189__10_,r_189__9_,r_189__8_,r_189__7_,
  r_189__6_,r_189__5_,r_189__4_,r_189__3_,r_189__2_,r_189__1_,r_189__0_,r_190__31_,
  r_190__30_,r_190__29_,r_190__28_,r_190__27_,r_190__26_,r_190__25_,r_190__24_,
  r_190__23_,r_190__22_,r_190__21_,r_190__20_,r_190__19_,r_190__18_,r_190__17_,r_190__16_,
  r_190__15_,r_190__14_,r_190__13_,r_190__12_,r_190__11_,r_190__10_,r_190__9_,
  r_190__8_,r_190__7_,r_190__6_,r_190__5_,r_190__4_,r_190__3_,r_190__2_,r_190__1_,
  r_190__0_,r_191__31_,r_191__30_,r_191__29_,r_191__28_,r_191__27_,r_191__26_,
  r_191__25_,r_191__24_,r_191__23_,r_191__22_,r_191__21_,r_191__20_,r_191__19_,r_191__18_,
  r_191__17_,r_191__16_,r_191__15_,r_191__14_,r_191__13_,r_191__12_,r_191__11_,
  r_191__10_,r_191__9_,r_191__8_,r_191__7_,r_191__6_,r_191__5_,r_191__4_,r_191__3_,
  r_191__2_,r_191__1_,r_191__0_,r_192__31_,r_192__30_,r_192__29_,r_192__28_,
  r_192__27_,r_192__26_,r_192__25_,r_192__24_,r_192__23_,r_192__22_,r_192__21_,r_192__20_,
  r_192__19_,r_192__18_,r_192__17_,r_192__16_,r_192__15_,r_192__14_,r_192__13_,
  r_192__12_,r_192__11_,r_192__10_,r_192__9_,r_192__8_,r_192__7_,r_192__6_,r_192__5_,
  r_192__4_,r_192__3_,r_192__2_,r_192__1_,r_192__0_,r_193__31_,r_193__30_,
  r_193__29_,r_193__28_,r_193__27_,r_193__26_,r_193__25_,r_193__24_,r_193__23_,r_193__22_,
  r_193__21_,r_193__20_,r_193__19_,r_193__18_,r_193__17_,r_193__16_,r_193__15_,
  r_193__14_,r_193__13_,r_193__12_,r_193__11_,r_193__10_,r_193__9_,r_193__8_,r_193__7_,
  r_193__6_,r_193__5_,r_193__4_,r_193__3_,r_193__2_,r_193__1_,r_193__0_,
  r_194__31_,r_194__30_,r_194__29_,r_194__28_,r_194__27_,r_194__26_,r_194__25_,r_194__24_,
  r_194__23_,r_194__22_,r_194__21_,r_194__20_,r_194__19_,r_194__18_,r_194__17_,
  r_194__16_,r_194__15_,r_194__14_,r_194__13_,r_194__12_,r_194__11_,r_194__10_,
  r_194__9_,r_194__8_,r_194__7_,r_194__6_,r_194__5_,r_194__4_,r_194__3_,r_194__2_,
  r_194__1_,r_194__0_,r_195__31_,r_195__30_,r_195__29_,r_195__28_,r_195__27_,r_195__26_,
  r_195__25_,r_195__24_,r_195__23_,r_195__22_,r_195__21_,r_195__20_,r_195__19_,
  r_195__18_,r_195__17_,r_195__16_,r_195__15_,r_195__14_,r_195__13_,r_195__12_,
  r_195__11_,r_195__10_,r_195__9_,r_195__8_,r_195__7_,r_195__6_,r_195__5_,r_195__4_,
  r_195__3_,r_195__2_,r_195__1_,r_195__0_,r_196__31_,r_196__30_,r_196__29_,r_196__28_,
  r_196__27_,r_196__26_,r_196__25_,r_196__24_,r_196__23_,r_196__22_,r_196__21_,
  r_196__20_,r_196__19_,r_196__18_,r_196__17_,r_196__16_,r_196__15_,r_196__14_,
  r_196__13_,r_196__12_,r_196__11_,r_196__10_,r_196__9_,r_196__8_,r_196__7_,r_196__6_,
  r_196__5_,r_196__4_,r_196__3_,r_196__2_,r_196__1_,r_196__0_,r_197__31_,r_197__30_,
  r_197__29_,r_197__28_,r_197__27_,r_197__26_,r_197__25_,r_197__24_,r_197__23_,
  r_197__22_,r_197__21_,r_197__20_,r_197__19_,r_197__18_,r_197__17_,r_197__16_,
  r_197__15_,r_197__14_,r_197__13_,r_197__12_,r_197__11_,r_197__10_,r_197__9_,r_197__8_,
  r_197__7_,r_197__6_,r_197__5_,r_197__4_,r_197__3_,r_197__2_,r_197__1_,r_197__0_,
  r_198__31_,r_198__30_,r_198__29_,r_198__28_,r_198__27_,r_198__26_,r_198__25_,
  r_198__24_,r_198__23_,r_198__22_,r_198__21_,r_198__20_,r_198__19_,r_198__18_,
  r_198__17_,r_198__16_,r_198__15_,r_198__14_,r_198__13_,r_198__12_,r_198__11_,r_198__10_,
  r_198__9_,r_198__8_,r_198__7_,r_198__6_,r_198__5_,r_198__4_,r_198__3_,r_198__2_,
  r_198__1_,r_198__0_,r_199__31_,r_199__30_,r_199__29_,r_199__28_,r_199__27_,
  r_199__26_,r_199__25_,r_199__24_,r_199__23_,r_199__22_,r_199__21_,r_199__20_,
  r_199__19_,r_199__18_,r_199__17_,r_199__16_,r_199__15_,r_199__14_,r_199__13_,r_199__12_,
  r_199__11_,r_199__10_,r_199__9_,r_199__8_,r_199__7_,r_199__6_,r_199__5_,
  r_199__4_,r_199__3_,r_199__2_,r_199__1_,r_199__0_,r_200__31_,r_200__30_,r_200__29_,
  r_200__28_,r_200__27_,r_200__26_,r_200__25_,r_200__24_,r_200__23_,r_200__22_,
  r_200__21_,r_200__20_,r_200__19_,r_200__18_,r_200__17_,r_200__16_,r_200__15_,r_200__14_,
  r_200__13_,r_200__12_,r_200__11_,r_200__10_,r_200__9_,r_200__8_,r_200__7_,
  r_200__6_,r_200__5_,r_200__4_,r_200__3_,r_200__2_,r_200__1_,r_200__0_,r_201__31_,
  r_201__30_,r_201__29_,r_201__28_,r_201__27_,r_201__26_,r_201__25_,r_201__24_,
  r_201__23_,r_201__22_,r_201__21_,r_201__20_,r_201__19_,r_201__18_,r_201__17_,r_201__16_,
  r_201__15_,r_201__14_,r_201__13_,r_201__12_,r_201__11_,r_201__10_,r_201__9_,
  r_201__8_,r_201__7_,r_201__6_,r_201__5_,r_201__4_,r_201__3_,r_201__2_,r_201__1_,
  r_201__0_,r_202__31_,r_202__30_,r_202__29_,r_202__28_,r_202__27_,r_202__26_,
  r_202__25_,r_202__24_,r_202__23_,r_202__22_,r_202__21_,r_202__20_,r_202__19_,r_202__18_,
  r_202__17_,r_202__16_,r_202__15_,r_202__14_,r_202__13_,r_202__12_,r_202__11_,
  r_202__10_,r_202__9_,r_202__8_,r_202__7_,r_202__6_,r_202__5_,r_202__4_,r_202__3_,
  r_202__2_,r_202__1_,r_202__0_,r_203__31_,r_203__30_,r_203__29_,r_203__28_,
  r_203__27_,r_203__26_,r_203__25_,r_203__24_,r_203__23_,r_203__22_,r_203__21_,r_203__20_,
  r_203__19_,r_203__18_,r_203__17_,r_203__16_,r_203__15_,r_203__14_,r_203__13_,
  r_203__12_,r_203__11_,r_203__10_,r_203__9_,r_203__8_,r_203__7_,r_203__6_,r_203__5_,
  r_203__4_,r_203__3_,r_203__2_,r_203__1_,r_203__0_,r_204__31_,r_204__30_,
  r_204__29_,r_204__28_,r_204__27_,r_204__26_,r_204__25_,r_204__24_,r_204__23_,r_204__22_,
  r_204__21_,r_204__20_,r_204__19_,r_204__18_,r_204__17_,r_204__16_,r_204__15_,
  r_204__14_,r_204__13_,r_204__12_,r_204__11_,r_204__10_,r_204__9_,r_204__8_,
  r_204__7_,r_204__6_,r_204__5_,r_204__4_,r_204__3_,r_204__2_,r_204__1_,r_204__0_,
  r_205__31_,r_205__30_,r_205__29_,r_205__28_,r_205__27_,r_205__26_,r_205__25_,r_205__24_,
  r_205__23_,r_205__22_,r_205__21_,r_205__20_,r_205__19_,r_205__18_,r_205__17_,
  r_205__16_,r_205__15_,r_205__14_,r_205__13_,r_205__12_,r_205__11_,r_205__10_,
  r_205__9_,r_205__8_,r_205__7_,r_205__6_,r_205__5_,r_205__4_,r_205__3_,r_205__2_,
  r_205__1_,r_205__0_,r_206__31_,r_206__30_,r_206__29_,r_206__28_,r_206__27_,r_206__26_,
  r_206__25_,r_206__24_,r_206__23_,r_206__22_,r_206__21_,r_206__20_,r_206__19_,
  r_206__18_,r_206__17_,r_206__16_,r_206__15_,r_206__14_,r_206__13_,r_206__12_,
  r_206__11_,r_206__10_,r_206__9_,r_206__8_,r_206__7_,r_206__6_,r_206__5_,r_206__4_,
  r_206__3_,r_206__2_,r_206__1_,r_206__0_,r_207__31_,r_207__30_,r_207__29_,r_207__28_,
  r_207__27_,r_207__26_,r_207__25_,r_207__24_,r_207__23_,r_207__22_,r_207__21_,
  r_207__20_,r_207__19_,r_207__18_,r_207__17_,r_207__16_,r_207__15_,r_207__14_,
  r_207__13_,r_207__12_,r_207__11_,r_207__10_,r_207__9_,r_207__8_,r_207__7_,r_207__6_,
  r_207__5_,r_207__4_,r_207__3_,r_207__2_,r_207__1_,r_207__0_,r_208__31_,r_208__30_,
  r_208__29_,r_208__28_,r_208__27_,r_208__26_,r_208__25_,r_208__24_,r_208__23_,
  r_208__22_,r_208__21_,r_208__20_,r_208__19_,r_208__18_,r_208__17_,r_208__16_,
  r_208__15_,r_208__14_,r_208__13_,r_208__12_,r_208__11_,r_208__10_,r_208__9_,r_208__8_,
  r_208__7_,r_208__6_,r_208__5_,r_208__4_,r_208__3_,r_208__2_,r_208__1_,r_208__0_,
  r_209__31_,r_209__30_,r_209__29_,r_209__28_,r_209__27_,r_209__26_,r_209__25_,
  r_209__24_,r_209__23_,r_209__22_,r_209__21_,r_209__20_,r_209__19_,r_209__18_,
  r_209__17_,r_209__16_,r_209__15_,r_209__14_,r_209__13_,r_209__12_,r_209__11_,
  r_209__10_,r_209__9_,r_209__8_,r_209__7_,r_209__6_,r_209__5_,r_209__4_,r_209__3_,
  r_209__2_,r_209__1_,r_209__0_,r_210__31_,r_210__30_,r_210__29_,r_210__28_,r_210__27_,
  r_210__26_,r_210__25_,r_210__24_,r_210__23_,r_210__22_,r_210__21_,r_210__20_,
  r_210__19_,r_210__18_,r_210__17_,r_210__16_,r_210__15_,r_210__14_,r_210__13_,
  r_210__12_,r_210__11_,r_210__10_,r_210__9_,r_210__8_,r_210__7_,r_210__6_,r_210__5_,
  r_210__4_,r_210__3_,r_210__2_,r_210__1_,r_210__0_,r_211__31_,r_211__30_,r_211__29_,
  r_211__28_,r_211__27_,r_211__26_,r_211__25_,r_211__24_,r_211__23_,r_211__22_,
  r_211__21_,r_211__20_,r_211__19_,r_211__18_,r_211__17_,r_211__16_,r_211__15_,
  r_211__14_,r_211__13_,r_211__12_,r_211__11_,r_211__10_,r_211__9_,r_211__8_,r_211__7_,
  r_211__6_,r_211__5_,r_211__4_,r_211__3_,r_211__2_,r_211__1_,r_211__0_,r_212__31_,
  r_212__30_,r_212__29_,r_212__28_,r_212__27_,r_212__26_,r_212__25_,r_212__24_,
  r_212__23_,r_212__22_,r_212__21_,r_212__20_,r_212__19_,r_212__18_,r_212__17_,
  r_212__16_,r_212__15_,r_212__14_,r_212__13_,r_212__12_,r_212__11_,r_212__10_,r_212__9_,
  r_212__8_,r_212__7_,r_212__6_,r_212__5_,r_212__4_,r_212__3_,r_212__2_,r_212__1_,
  r_212__0_,r_213__31_,r_213__30_,r_213__29_,r_213__28_,r_213__27_,r_213__26_,
  r_213__25_,r_213__24_,r_213__23_,r_213__22_,r_213__21_,r_213__20_,r_213__19_,
  r_213__18_,r_213__17_,r_213__16_,r_213__15_,r_213__14_,r_213__13_,r_213__12_,r_213__11_,
  r_213__10_,r_213__9_,r_213__8_,r_213__7_,r_213__6_,r_213__5_,r_213__4_,r_213__3_,
  r_213__2_,r_213__1_,r_213__0_,r_214__31_,r_214__30_,r_214__29_,r_214__28_,
  r_214__27_,r_214__26_,r_214__25_,r_214__24_,r_214__23_,r_214__22_,r_214__21_,
  r_214__20_,r_214__19_,r_214__18_,r_214__17_,r_214__16_,r_214__15_,r_214__14_,r_214__13_,
  r_214__12_,r_214__11_,r_214__10_,r_214__9_,r_214__8_,r_214__7_,r_214__6_,
  r_214__5_,r_214__4_,r_214__3_,r_214__2_,r_214__1_,r_214__0_,r_215__31_,r_215__30_,
  r_215__29_,r_215__28_,r_215__27_,r_215__26_,r_215__25_,r_215__24_,r_215__23_,
  r_215__22_,r_215__21_,r_215__20_,r_215__19_,r_215__18_,r_215__17_,r_215__16_,r_215__15_,
  r_215__14_,r_215__13_,r_215__12_,r_215__11_,r_215__10_,r_215__9_,r_215__8_,
  r_215__7_,r_215__6_,r_215__5_,r_215__4_,r_215__3_,r_215__2_,r_215__1_,r_215__0_,
  r_216__31_,r_216__30_,r_216__29_,r_216__28_,r_216__27_,r_216__26_,r_216__25_,
  r_216__24_,r_216__23_,r_216__22_,r_216__21_,r_216__20_,r_216__19_,r_216__18_,r_216__17_,
  r_216__16_,r_216__15_,r_216__14_,r_216__13_,r_216__12_,r_216__11_,r_216__10_,
  r_216__9_,r_216__8_,r_216__7_,r_216__6_,r_216__5_,r_216__4_,r_216__3_,r_216__2_,
  r_216__1_,r_216__0_,r_217__31_,r_217__30_,r_217__29_,r_217__28_,r_217__27_,
  r_217__26_,r_217__25_,r_217__24_,r_217__23_,r_217__22_,r_217__21_,r_217__20_,r_217__19_,
  r_217__18_,r_217__17_,r_217__16_,r_217__15_,r_217__14_,r_217__13_,r_217__12_,
  r_217__11_,r_217__10_,r_217__9_,r_217__8_,r_217__7_,r_217__6_,r_217__5_,r_217__4_,
  r_217__3_,r_217__2_,r_217__1_,r_217__0_,r_218__31_,r_218__30_,r_218__29_,
  r_218__28_,r_218__27_,r_218__26_,r_218__25_,r_218__24_,r_218__23_,r_218__22_,r_218__21_,
  r_218__20_,r_218__19_,r_218__18_,r_218__17_,r_218__16_,r_218__15_,r_218__14_,
  r_218__13_,r_218__12_,r_218__11_,r_218__10_,r_218__9_,r_218__8_,r_218__7_,r_218__6_,
  r_218__5_,r_218__4_,r_218__3_,r_218__2_,r_218__1_,r_218__0_,r_219__31_,
  r_219__30_,r_219__29_,r_219__28_,r_219__27_,r_219__26_,r_219__25_,r_219__24_,r_219__23_,
  r_219__22_,r_219__21_,r_219__20_,r_219__19_,r_219__18_,r_219__17_,r_219__16_,
  r_219__15_,r_219__14_,r_219__13_,r_219__12_,r_219__11_,r_219__10_,r_219__9_,
  r_219__8_,r_219__7_,r_219__6_,r_219__5_,r_219__4_,r_219__3_,r_219__2_,r_219__1_,
  r_219__0_,r_220__31_,r_220__30_,r_220__29_,r_220__28_,r_220__27_,r_220__26_,r_220__25_,
  r_220__24_,r_220__23_,r_220__22_,r_220__21_,r_220__20_,r_220__19_,r_220__18_,
  r_220__17_,r_220__16_,r_220__15_,r_220__14_,r_220__13_,r_220__12_,r_220__11_,
  r_220__10_,r_220__9_,r_220__8_,r_220__7_,r_220__6_,r_220__5_,r_220__4_,r_220__3_,
  r_220__2_,r_220__1_,r_220__0_,r_221__31_,r_221__30_,r_221__29_,r_221__28_,r_221__27_,
  r_221__26_,r_221__25_,r_221__24_,r_221__23_,r_221__22_,r_221__21_,r_221__20_,
  r_221__19_,r_221__18_,r_221__17_,r_221__16_,r_221__15_,r_221__14_,r_221__13_,
  r_221__12_,r_221__11_,r_221__10_,r_221__9_,r_221__8_,r_221__7_,r_221__6_,r_221__5_,
  r_221__4_,r_221__3_,r_221__2_,r_221__1_,r_221__0_,r_222__31_,r_222__30_,r_222__29_,
  r_222__28_,r_222__27_,r_222__26_,r_222__25_,r_222__24_,r_222__23_,r_222__22_,
  r_222__21_,r_222__20_,r_222__19_,r_222__18_,r_222__17_,r_222__16_,r_222__15_,
  r_222__14_,r_222__13_,r_222__12_,r_222__11_,r_222__10_,r_222__9_,r_222__8_,r_222__7_,
  r_222__6_,r_222__5_,r_222__4_,r_222__3_,r_222__2_,r_222__1_,r_222__0_,r_223__31_,
  r_223__30_,r_223__29_,r_223__28_,r_223__27_,r_223__26_,r_223__25_,r_223__24_,
  r_223__23_,r_223__22_,r_223__21_,r_223__20_,r_223__19_,r_223__18_,r_223__17_,
  r_223__16_,r_223__15_,r_223__14_,r_223__13_,r_223__12_,r_223__11_,r_223__10_,r_223__9_,
  r_223__8_,r_223__7_,r_223__6_,r_223__5_,r_223__4_,r_223__3_,r_223__2_,r_223__1_,
  r_223__0_,r_224__31_,r_224__30_,r_224__29_,r_224__28_,r_224__27_,r_224__26_,
  r_224__25_,r_224__24_,r_224__23_,r_224__22_,r_224__21_,r_224__20_,r_224__19_,
  r_224__18_,r_224__17_,r_224__16_,r_224__15_,r_224__14_,r_224__13_,r_224__12_,
  r_224__11_,r_224__10_,r_224__9_,r_224__8_,r_224__7_,r_224__6_,r_224__5_,r_224__4_,
  r_224__3_,r_224__2_,r_224__1_,r_224__0_,r_225__31_,r_225__30_,r_225__29_,r_225__28_,
  r_225__27_,r_225__26_,r_225__25_,r_225__24_,r_225__23_,r_225__22_,r_225__21_,
  r_225__20_,r_225__19_,r_225__18_,r_225__17_,r_225__16_,r_225__15_,r_225__14_,
  r_225__13_,r_225__12_,r_225__11_,r_225__10_,r_225__9_,r_225__8_,r_225__7_,r_225__6_,
  r_225__5_,r_225__4_,r_225__3_,r_225__2_,r_225__1_,r_225__0_,r_226__31_,r_226__30_,
  r_226__29_,r_226__28_,r_226__27_,r_226__26_,r_226__25_,r_226__24_,r_226__23_,
  r_226__22_,r_226__21_,r_226__20_,r_226__19_,r_226__18_,r_226__17_,r_226__16_,
  r_226__15_,r_226__14_,r_226__13_,r_226__12_,r_226__11_,r_226__10_,r_226__9_,r_226__8_,
  r_226__7_,r_226__6_,r_226__5_,r_226__4_,r_226__3_,r_226__2_,r_226__1_,r_226__0_,
  r_227__31_,r_227__30_,r_227__29_,r_227__28_,r_227__27_,r_227__26_,r_227__25_,
  r_227__24_,r_227__23_,r_227__22_,r_227__21_,r_227__20_,r_227__19_,r_227__18_,
  r_227__17_,r_227__16_,r_227__15_,r_227__14_,r_227__13_,r_227__12_,r_227__11_,r_227__10_,
  r_227__9_,r_227__8_,r_227__7_,r_227__6_,r_227__5_,r_227__4_,r_227__3_,r_227__2_,
  r_227__1_,r_227__0_,r_228__31_,r_228__30_,r_228__29_,r_228__28_,r_228__27_,
  r_228__26_,r_228__25_,r_228__24_,r_228__23_,r_228__22_,r_228__21_,r_228__20_,
  r_228__19_,r_228__18_,r_228__17_,r_228__16_,r_228__15_,r_228__14_,r_228__13_,r_228__12_,
  r_228__11_,r_228__10_,r_228__9_,r_228__8_,r_228__7_,r_228__6_,r_228__5_,r_228__4_,
  r_228__3_,r_228__2_,r_228__1_,r_228__0_,r_229__31_,r_229__30_,r_229__29_,
  r_229__28_,r_229__27_,r_229__26_,r_229__25_,r_229__24_,r_229__23_,r_229__22_,
  r_229__21_,r_229__20_,r_229__19_,r_229__18_,r_229__17_,r_229__16_,r_229__15_,r_229__14_,
  r_229__13_,r_229__12_,r_229__11_,r_229__10_,r_229__9_,r_229__8_,r_229__7_,
  r_229__6_,r_229__5_,r_229__4_,r_229__3_,r_229__2_,r_229__1_,r_229__0_,r_230__31_,
  r_230__30_,r_230__29_,r_230__28_,r_230__27_,r_230__26_,r_230__25_,r_230__24_,
  r_230__23_,r_230__22_,r_230__21_,r_230__20_,r_230__19_,r_230__18_,r_230__17_,r_230__16_,
  r_230__15_,r_230__14_,r_230__13_,r_230__12_,r_230__11_,r_230__10_,r_230__9_,
  r_230__8_,r_230__7_,r_230__6_,r_230__5_,r_230__4_,r_230__3_,r_230__2_,r_230__1_,
  r_230__0_,r_231__31_,r_231__30_,r_231__29_,r_231__28_,r_231__27_,r_231__26_,
  r_231__25_,r_231__24_,r_231__23_,r_231__22_,r_231__21_,r_231__20_,r_231__19_,r_231__18_,
  r_231__17_,r_231__16_,r_231__15_,r_231__14_,r_231__13_,r_231__12_,r_231__11_,
  r_231__10_,r_231__9_,r_231__8_,r_231__7_,r_231__6_,r_231__5_,r_231__4_,r_231__3_,
  r_231__2_,r_231__1_,r_231__0_,r_232__31_,r_232__30_,r_232__29_,r_232__28_,
  r_232__27_,r_232__26_,r_232__25_,r_232__24_,r_232__23_,r_232__22_,r_232__21_,r_232__20_,
  r_232__19_,r_232__18_,r_232__17_,r_232__16_,r_232__15_,r_232__14_,r_232__13_,
  r_232__12_,r_232__11_,r_232__10_,r_232__9_,r_232__8_,r_232__7_,r_232__6_,r_232__5_,
  r_232__4_,r_232__3_,r_232__2_,r_232__1_,r_232__0_,r_233__31_,r_233__30_,
  r_233__29_,r_233__28_,r_233__27_,r_233__26_,r_233__25_,r_233__24_,r_233__23_,r_233__22_,
  r_233__21_,r_233__20_,r_233__19_,r_233__18_,r_233__17_,r_233__16_,r_233__15_,
  r_233__14_,r_233__13_,r_233__12_,r_233__11_,r_233__10_,r_233__9_,r_233__8_,r_233__7_,
  r_233__6_,r_233__5_,r_233__4_,r_233__3_,r_233__2_,r_233__1_,r_233__0_,
  r_234__31_,r_234__30_,r_234__29_,r_234__28_,r_234__27_,r_234__26_,r_234__25_,r_234__24_,
  r_234__23_,r_234__22_,r_234__21_,r_234__20_,r_234__19_,r_234__18_,r_234__17_,
  r_234__16_,r_234__15_,r_234__14_,r_234__13_,r_234__12_,r_234__11_,r_234__10_,
  r_234__9_,r_234__8_,r_234__7_,r_234__6_,r_234__5_,r_234__4_,r_234__3_,r_234__2_,
  r_234__1_,r_234__0_,r_235__31_,r_235__30_,r_235__29_,r_235__28_,r_235__27_,r_235__26_,
  r_235__25_,r_235__24_,r_235__23_,r_235__22_,r_235__21_,r_235__20_,r_235__19_,
  r_235__18_,r_235__17_,r_235__16_,r_235__15_,r_235__14_,r_235__13_,r_235__12_,
  r_235__11_,r_235__10_,r_235__9_,r_235__8_,r_235__7_,r_235__6_,r_235__5_,r_235__4_,
  r_235__3_,r_235__2_,r_235__1_,r_235__0_,r_236__31_,r_236__30_,r_236__29_,r_236__28_,
  r_236__27_,r_236__26_,r_236__25_,r_236__24_,r_236__23_,r_236__22_,r_236__21_,
  r_236__20_,r_236__19_,r_236__18_,r_236__17_,r_236__16_,r_236__15_,r_236__14_,
  r_236__13_,r_236__12_,r_236__11_,r_236__10_,r_236__9_,r_236__8_,r_236__7_,r_236__6_,
  r_236__5_,r_236__4_,r_236__3_,r_236__2_,r_236__1_,r_236__0_,r_237__31_,r_237__30_,
  r_237__29_,r_237__28_,r_237__27_,r_237__26_,r_237__25_,r_237__24_,r_237__23_,
  r_237__22_,r_237__21_,r_237__20_,r_237__19_,r_237__18_,r_237__17_,r_237__16_,
  r_237__15_,r_237__14_,r_237__13_,r_237__12_,r_237__11_,r_237__10_,r_237__9_,r_237__8_,
  r_237__7_,r_237__6_,r_237__5_,r_237__4_,r_237__3_,r_237__2_,r_237__1_,r_237__0_,
  r_238__31_,r_238__30_,r_238__29_,r_238__28_,r_238__27_,r_238__26_,r_238__25_,
  r_238__24_,r_238__23_,r_238__22_,r_238__21_,r_238__20_,r_238__19_,r_238__18_,
  r_238__17_,r_238__16_,r_238__15_,r_238__14_,r_238__13_,r_238__12_,r_238__11_,r_238__10_,
  r_238__9_,r_238__8_,r_238__7_,r_238__6_,r_238__5_,r_238__4_,r_238__3_,r_238__2_,
  r_238__1_,r_238__0_,r_239__31_,r_239__30_,r_239__29_,r_239__28_,r_239__27_,
  r_239__26_,r_239__25_,r_239__24_,r_239__23_,r_239__22_,r_239__21_,r_239__20_,
  r_239__19_,r_239__18_,r_239__17_,r_239__16_,r_239__15_,r_239__14_,r_239__13_,r_239__12_,
  r_239__11_,r_239__10_,r_239__9_,r_239__8_,r_239__7_,r_239__6_,r_239__5_,
  r_239__4_,r_239__3_,r_239__2_,r_239__1_,r_239__0_,r_240__31_,r_240__30_,r_240__29_,
  r_240__28_,r_240__27_,r_240__26_,r_240__25_,r_240__24_,r_240__23_,r_240__22_,
  r_240__21_,r_240__20_,r_240__19_,r_240__18_,r_240__17_,r_240__16_,r_240__15_,r_240__14_,
  r_240__13_,r_240__12_,r_240__11_,r_240__10_,r_240__9_,r_240__8_,r_240__7_,
  r_240__6_,r_240__5_,r_240__4_,r_240__3_,r_240__2_,r_240__1_,r_240__0_,r_241__31_,
  r_241__30_,r_241__29_,r_241__28_,r_241__27_,r_241__26_,r_241__25_,r_241__24_,
  r_241__23_,r_241__22_,r_241__21_,r_241__20_,r_241__19_,r_241__18_,r_241__17_,r_241__16_,
  r_241__15_,r_241__14_,r_241__13_,r_241__12_,r_241__11_,r_241__10_,r_241__9_,
  r_241__8_,r_241__7_,r_241__6_,r_241__5_,r_241__4_,r_241__3_,r_241__2_,r_241__1_,
  r_241__0_,r_242__31_,r_242__30_,r_242__29_,r_242__28_,r_242__27_,r_242__26_,
  r_242__25_,r_242__24_,r_242__23_,r_242__22_,r_242__21_,r_242__20_,r_242__19_,r_242__18_,
  r_242__17_,r_242__16_,r_242__15_,r_242__14_,r_242__13_,r_242__12_,r_242__11_,
  r_242__10_,r_242__9_,r_242__8_,r_242__7_,r_242__6_,r_242__5_,r_242__4_,r_242__3_,
  r_242__2_,r_242__1_,r_242__0_,r_243__31_,r_243__30_,r_243__29_,r_243__28_,
  r_243__27_,r_243__26_,r_243__25_,r_243__24_,r_243__23_,r_243__22_,r_243__21_,r_243__20_,
  r_243__19_,r_243__18_,r_243__17_,r_243__16_,r_243__15_,r_243__14_,r_243__13_,
  r_243__12_,r_243__11_,r_243__10_,r_243__9_,r_243__8_,r_243__7_,r_243__6_,r_243__5_,
  r_243__4_,r_243__3_,r_243__2_,r_243__1_,r_243__0_,r_244__31_,r_244__30_,
  r_244__29_,r_244__28_,r_244__27_,r_244__26_,r_244__25_,r_244__24_,r_244__23_,r_244__22_,
  r_244__21_,r_244__20_,r_244__19_,r_244__18_,r_244__17_,r_244__16_,r_244__15_,
  r_244__14_,r_244__13_,r_244__12_,r_244__11_,r_244__10_,r_244__9_,r_244__8_,
  r_244__7_,r_244__6_,r_244__5_,r_244__4_,r_244__3_,r_244__2_,r_244__1_,r_244__0_,
  r_245__31_,r_245__30_,r_245__29_,r_245__28_,r_245__27_,r_245__26_,r_245__25_,r_245__24_,
  r_245__23_,r_245__22_,r_245__21_,r_245__20_,r_245__19_,r_245__18_,r_245__17_,
  r_245__16_,r_245__15_,r_245__14_,r_245__13_,r_245__12_,r_245__11_,r_245__10_,
  r_245__9_,r_245__8_,r_245__7_,r_245__6_,r_245__5_,r_245__4_,r_245__3_,r_245__2_,
  r_245__1_,r_245__0_,r_246__31_,r_246__30_,r_246__29_,r_246__28_,r_246__27_,r_246__26_,
  r_246__25_,r_246__24_,r_246__23_,r_246__22_,r_246__21_,r_246__20_,r_246__19_,
  r_246__18_,r_246__17_,r_246__16_,r_246__15_,r_246__14_,r_246__13_,r_246__12_,
  r_246__11_,r_246__10_,r_246__9_,r_246__8_,r_246__7_,r_246__6_,r_246__5_,r_246__4_,
  r_246__3_,r_246__2_,r_246__1_,r_246__0_,r_247__31_,r_247__30_,r_247__29_,r_247__28_,
  r_247__27_,r_247__26_,r_247__25_,r_247__24_,r_247__23_,r_247__22_,r_247__21_,
  r_247__20_,r_247__19_,r_247__18_,r_247__17_,r_247__16_,r_247__15_,r_247__14_,
  r_247__13_,r_247__12_,r_247__11_,r_247__10_,r_247__9_,r_247__8_,r_247__7_,r_247__6_,
  r_247__5_,r_247__4_,r_247__3_,r_247__2_,r_247__1_,r_247__0_,r_248__31_,r_248__30_,
  r_248__29_,r_248__28_,r_248__27_,r_248__26_,r_248__25_,r_248__24_,r_248__23_,
  r_248__22_,r_248__21_,r_248__20_,r_248__19_,r_248__18_,r_248__17_,r_248__16_,
  r_248__15_,r_248__14_,r_248__13_,r_248__12_,r_248__11_,r_248__10_,r_248__9_,r_248__8_,
  r_248__7_,r_248__6_,r_248__5_,r_248__4_,r_248__3_,r_248__2_,r_248__1_,r_248__0_,
  r_249__31_,r_249__30_,r_249__29_,r_249__28_,r_249__27_,r_249__26_,r_249__25_,
  r_249__24_,r_249__23_,r_249__22_,r_249__21_,r_249__20_,r_249__19_,r_249__18_,
  r_249__17_,r_249__16_,r_249__15_,r_249__14_,r_249__13_,r_249__12_,r_249__11_,
  r_249__10_,r_249__9_,r_249__8_,r_249__7_,r_249__6_,r_249__5_,r_249__4_,r_249__3_,
  r_249__2_,r_249__1_,r_249__0_,r_250__31_,r_250__30_,r_250__29_,r_250__28_,r_250__27_,
  r_250__26_,r_250__25_,r_250__24_,r_250__23_,r_250__22_,r_250__21_,r_250__20_,
  r_250__19_,r_250__18_,r_250__17_,r_250__16_,r_250__15_,r_250__14_,r_250__13_,
  r_250__12_,r_250__11_,r_250__10_,r_250__9_,r_250__8_,r_250__7_,r_250__6_,r_250__5_,
  r_250__4_,r_250__3_,r_250__2_,r_250__1_,r_250__0_,r_251__31_,r_251__30_,r_251__29_,
  r_251__28_,r_251__27_,r_251__26_,r_251__25_,r_251__24_,r_251__23_,r_251__22_,
  r_251__21_,r_251__20_,r_251__19_,r_251__18_,r_251__17_,r_251__16_,r_251__15_,
  r_251__14_,r_251__13_,r_251__12_,r_251__11_,r_251__10_,r_251__9_,r_251__8_,r_251__7_,
  r_251__6_,r_251__5_,r_251__4_,r_251__3_,r_251__2_,r_251__1_,r_251__0_,r_252__31_,
  r_252__30_,r_252__29_,r_252__28_,r_252__27_,r_252__26_,r_252__25_,r_252__24_,
  r_252__23_,r_252__22_,r_252__21_,r_252__20_,r_252__19_,r_252__18_,r_252__17_,
  r_252__16_,r_252__15_,r_252__14_,r_252__13_,r_252__12_,r_252__11_,r_252__10_,r_252__9_,
  r_252__8_,r_252__7_,r_252__6_,r_252__5_,r_252__4_,r_252__3_,r_252__2_,r_252__1_,
  r_252__0_,r_253__31_,r_253__30_,r_253__29_,r_253__28_,r_253__27_,r_253__26_,
  r_253__25_,r_253__24_,r_253__23_,r_253__22_,r_253__21_,r_253__20_,r_253__19_,
  r_253__18_,r_253__17_,r_253__16_,r_253__15_,r_253__14_,r_253__13_,r_253__12_,r_253__11_,
  r_253__10_,r_253__9_,r_253__8_,r_253__7_,r_253__6_,r_253__5_,r_253__4_,r_253__3_,
  r_253__2_,r_253__1_,r_253__0_,r_254__31_,r_254__30_,r_254__29_,r_254__28_,
  r_254__27_,r_254__26_,r_254__25_,r_254__24_,r_254__23_,r_254__22_,r_254__21_,
  r_254__20_,r_254__19_,r_254__18_,r_254__17_,r_254__16_,r_254__15_,r_254__14_,r_254__13_,
  r_254__12_,r_254__11_,r_254__10_,r_254__9_,r_254__8_,r_254__7_,r_254__6_,
  r_254__5_,r_254__4_,r_254__3_,r_254__2_,r_254__1_,r_254__0_,r_255__31_,r_255__30_,
  r_255__29_,r_255__28_,r_255__27_,r_255__26_,r_255__25_,r_255__24_,r_255__23_,
  r_255__22_,r_255__21_,r_255__20_,r_255__19_,r_255__18_,r_255__17_,r_255__16_,r_255__15_,
  r_255__14_,r_255__13_,r_255__12_,r_255__11_,r_255__10_,r_255__9_,r_255__8_,
  r_255__7_,r_255__6_,r_255__5_,r_255__4_,r_255__3_,r_255__2_,r_255__1_,r_255__0_;
  assign N512 = sel_i[1] & sel_i[0];
  assign N514 = N513 & N516;
  assign N517 = sel_i[3] & sel_i[2];
  assign N519 = N518 & N521;
  assign N522 = sel_i[5] & sel_i[4];
  assign N524 = N523 & N526;
  assign N527 = sel_i[7] & sel_i[6];
  assign N529 = N528 & N531;
  assign N532 = sel_i[9] & sel_i[8];
  assign N534 = N533 & N536;
  assign N537 = sel_i[11] & sel_i[10];
  assign N539 = N538 & N541;
  assign N542 = sel_i[13] & sel_i[12];
  assign N544 = N543 & N546;
  assign N547 = sel_i[15] & sel_i[14];
  assign N549 = N548 & N551;
  assign N552 = sel_i[17] & sel_i[16];
  assign N554 = N553 & N556;
  assign N557 = sel_i[19] & sel_i[18];
  assign N559 = N558 & N561;
  assign N562 = sel_i[21] & sel_i[20];
  assign N564 = N563 & N566;
  assign N567 = sel_i[23] & sel_i[22];
  assign N569 = N568 & N571;
  assign N572 = sel_i[25] & sel_i[24];
  assign N574 = N573 & N576;
  assign N577 = sel_i[27] & sel_i[26];
  assign N579 = N578 & N581;
  assign N582 = sel_i[29] & sel_i[28];
  assign N584 = N583 & N586;
  assign N587 = sel_i[31] & sel_i[30];
  assign N589 = N588 & N591;
  assign N592 = sel_i[33] & sel_i[32];
  assign N594 = N593 & N596;
  assign N597 = sel_i[35] & sel_i[34];
  assign N599 = N598 & N601;
  assign N602 = sel_i[37] & sel_i[36];
  assign N604 = N603 & N606;
  assign N607 = sel_i[39] & sel_i[38];
  assign N609 = N608 & N611;
  assign N612 = sel_i[41] & sel_i[40];
  assign N614 = N613 & N616;
  assign N617 = sel_i[43] & sel_i[42];
  assign N619 = N618 & N621;
  assign N622 = sel_i[45] & sel_i[44];
  assign N624 = N623 & N626;
  assign N627 = sel_i[47] & sel_i[46];
  assign N629 = N628 & N631;
  assign N632 = sel_i[49] & sel_i[48];
  assign N634 = N633 & N636;
  assign N637 = sel_i[51] & sel_i[50];
  assign N639 = N638 & N641;
  assign N642 = sel_i[53] & sel_i[52];
  assign N644 = N643 & N646;
  assign N647 = sel_i[55] & sel_i[54];
  assign N649 = N648 & N651;
  assign N652 = sel_i[57] & sel_i[56];
  assign N654 = N653 & N656;
  assign N657 = sel_i[59] & sel_i[58];
  assign N659 = N658 & N661;
  assign N662 = sel_i[61] & sel_i[60];
  assign N664 = N663 & N666;
  assign N667 = sel_i[63] & sel_i[62];
  assign N669 = N668 & N671;
  assign N672 = sel_i[65] & sel_i[64];
  assign N674 = N673 & N676;
  assign N677 = sel_i[67] & sel_i[66];
  assign N679 = N678 & N681;
  assign N682 = sel_i[69] & sel_i[68];
  assign N684 = N683 & N686;
  assign N687 = sel_i[71] & sel_i[70];
  assign N689 = N688 & N691;
  assign N692 = sel_i[73] & sel_i[72];
  assign N694 = N693 & N696;
  assign N697 = sel_i[75] & sel_i[74];
  assign N699 = N698 & N701;
  assign N702 = sel_i[77] & sel_i[76];
  assign N704 = N703 & N706;
  assign N707 = sel_i[79] & sel_i[78];
  assign N709 = N708 & N711;
  assign N712 = sel_i[81] & sel_i[80];
  assign N714 = N713 & N716;
  assign N717 = sel_i[83] & sel_i[82];
  assign N719 = N718 & N721;
  assign N722 = sel_i[85] & sel_i[84];
  assign N724 = N723 & N726;
  assign N727 = sel_i[87] & sel_i[86];
  assign N729 = N728 & N731;
  assign N732 = sel_i[89] & sel_i[88];
  assign N734 = N733 & N736;
  assign N737 = sel_i[91] & sel_i[90];
  assign N739 = N738 & N741;
  assign N742 = sel_i[93] & sel_i[92];
  assign N744 = N743 & N746;
  assign N747 = sel_i[95] & sel_i[94];
  assign N749 = N748 & N751;
  assign N752 = sel_i[97] & sel_i[96];
  assign N754 = N753 & N756;
  assign N757 = sel_i[99] & sel_i[98];
  assign N759 = N758 & N761;
  assign N762 = sel_i[101] & sel_i[100];
  assign N764 = N763 & N766;
  assign N767 = sel_i[103] & sel_i[102];
  assign N769 = N768 & N771;
  assign N772 = sel_i[105] & sel_i[104];
  assign N774 = N773 & N776;
  assign N777 = sel_i[107] & sel_i[106];
  assign N779 = N778 & N781;
  assign N782 = sel_i[109] & sel_i[108];
  assign N784 = N783 & N786;
  assign N787 = sel_i[111] & sel_i[110];
  assign N789 = N788 & N791;
  assign N792 = sel_i[113] & sel_i[112];
  assign N794 = N793 & N796;
  assign N797 = sel_i[115] & sel_i[114];
  assign N799 = N798 & N801;
  assign N802 = sel_i[117] & sel_i[116];
  assign N804 = N803 & N806;
  assign N807 = sel_i[119] & sel_i[118];
  assign N809 = N808 & N811;
  assign N812 = sel_i[121] & sel_i[120];
  assign N814 = N813 & N816;
  assign N817 = sel_i[123] & sel_i[122];
  assign N819 = N818 & N821;
  assign N822 = sel_i[125] & sel_i[124];
  assign N824 = N823 & N826;
  assign N827 = sel_i[127] & sel_i[126];
  assign N829 = N828 & N831;
  assign N832 = sel_i[129] & sel_i[128];
  assign N834 = N833 & N836;
  assign N837 = sel_i[131] & sel_i[130];
  assign N839 = N838 & N841;
  assign N842 = sel_i[133] & sel_i[132];
  assign N844 = N843 & N846;
  assign N847 = sel_i[135] & sel_i[134];
  assign N849 = N848 & N851;
  assign N852 = sel_i[137] & sel_i[136];
  assign N854 = N853 & N856;
  assign N857 = sel_i[139] & sel_i[138];
  assign N859 = N858 & N861;
  assign N862 = sel_i[141] & sel_i[140];
  assign N864 = N863 & N866;
  assign N867 = sel_i[143] & sel_i[142];
  assign N869 = N868 & N871;
  assign N872 = sel_i[145] & sel_i[144];
  assign N874 = N873 & N876;
  assign N877 = sel_i[147] & sel_i[146];
  assign N879 = N878 & N881;
  assign N882 = sel_i[149] & sel_i[148];
  assign N884 = N883 & N886;
  assign N887 = sel_i[151] & sel_i[150];
  assign N889 = N888 & N891;
  assign N892 = sel_i[153] & sel_i[152];
  assign N894 = N893 & N896;
  assign N897 = sel_i[155] & sel_i[154];
  assign N899 = N898 & N901;
  assign N902 = sel_i[157] & sel_i[156];
  assign N904 = N903 & N906;
  assign N907 = sel_i[159] & sel_i[158];
  assign N909 = N908 & N911;
  assign N912 = sel_i[161] & sel_i[160];
  assign N914 = N913 & N916;
  assign N917 = sel_i[163] & sel_i[162];
  assign N919 = N918 & N921;
  assign N922 = sel_i[165] & sel_i[164];
  assign N924 = N923 & N926;
  assign N927 = sel_i[167] & sel_i[166];
  assign N929 = N928 & N931;
  assign N932 = sel_i[169] & sel_i[168];
  assign N934 = N933 & N936;
  assign N937 = sel_i[171] & sel_i[170];
  assign N939 = N938 & N941;
  assign N942 = sel_i[173] & sel_i[172];
  assign N944 = N943 & N946;
  assign N947 = sel_i[175] & sel_i[174];
  assign N949 = N948 & N951;
  assign N952 = sel_i[177] & sel_i[176];
  assign N954 = N953 & N956;
  assign N957 = sel_i[179] & sel_i[178];
  assign N959 = N958 & N961;
  assign N962 = sel_i[181] & sel_i[180];
  assign N964 = N963 & N966;
  assign N967 = sel_i[183] & sel_i[182];
  assign N969 = N968 & N971;
  assign N972 = sel_i[185] & sel_i[184];
  assign N974 = N973 & N976;
  assign N977 = sel_i[187] & sel_i[186];
  assign N979 = N978 & N981;
  assign N982 = sel_i[189] & sel_i[188];
  assign N984 = N983 & N986;
  assign N987 = sel_i[191] & sel_i[190];
  assign N989 = N988 & N991;
  assign N992 = sel_i[193] & sel_i[192];
  assign N994 = N993 & N996;
  assign N997 = sel_i[195] & sel_i[194];
  assign N999 = N998 & N1001;
  assign N1002 = sel_i[197] & sel_i[196];
  assign N1004 = N1003 & N1006;
  assign N1007 = sel_i[199] & sel_i[198];
  assign N1009 = N1008 & N1011;
  assign N1012 = sel_i[201] & sel_i[200];
  assign N1014 = N1013 & N1016;
  assign N1017 = sel_i[203] & sel_i[202];
  assign N1019 = N1018 & N1021;
  assign N1022 = sel_i[205] & sel_i[204];
  assign N1024 = N1023 & N1026;
  assign N1027 = sel_i[207] & sel_i[206];
  assign N1029 = N1028 & N1031;
  assign N1032 = sel_i[209] & sel_i[208];
  assign N1034 = N1033 & N1036;
  assign N1037 = sel_i[211] & sel_i[210];
  assign N1039 = N1038 & N1041;
  assign N1042 = sel_i[213] & sel_i[212];
  assign N1044 = N1043 & N1046;
  assign N1047 = sel_i[215] & sel_i[214];
  assign N1049 = N1048 & N1051;
  assign N1052 = sel_i[217] & sel_i[216];
  assign N1054 = N1053 & N1056;
  assign N1057 = sel_i[219] & sel_i[218];
  assign N1059 = N1058 & N1061;
  assign N1062 = sel_i[221] & sel_i[220];
  assign N1064 = N1063 & N1066;
  assign N1067 = sel_i[223] & sel_i[222];
  assign N1069 = N1068 & N1071;
  assign N1072 = sel_i[225] & sel_i[224];
  assign N1074 = N1073 & N1076;
  assign N1077 = sel_i[227] & sel_i[226];
  assign N1079 = N1078 & N1081;
  assign N1082 = sel_i[229] & sel_i[228];
  assign N1084 = N1083 & N1086;
  assign N1087 = sel_i[231] & sel_i[230];
  assign N1089 = N1088 & N1091;
  assign N1092 = sel_i[233] & sel_i[232];
  assign N1094 = N1093 & N1096;
  assign N1097 = sel_i[235] & sel_i[234];
  assign N1099 = N1098 & N1101;
  assign N1102 = sel_i[237] & sel_i[236];
  assign N1104 = N1103 & N1106;
  assign N1107 = sel_i[239] & sel_i[238];
  assign N1109 = N1108 & N1111;
  assign N1112 = sel_i[241] & sel_i[240];
  assign N1114 = N1113 & N1116;
  assign N1117 = sel_i[243] & sel_i[242];
  assign N1119 = N1118 & N1121;
  assign N1122 = sel_i[245] & sel_i[244];
  assign N1124 = N1123 & N1126;
  assign N1127 = sel_i[247] & sel_i[246];
  assign N1129 = N1128 & N1131;
  assign N1132 = sel_i[249] & sel_i[248];
  assign N1134 = N1133 & N1136;
  assign N1137 = sel_i[251] & sel_i[250];
  assign N1139 = N1138 & N1141;
  assign N1142 = sel_i[253] & sel_i[252];
  assign N1144 = N1143 & N1146;
  assign N1147 = sel_i[255] & sel_i[254];
  assign N1149 = N1148 & N1151;
  assign N1152 = sel_i[257] & sel_i[256];
  assign N1154 = N1153 & N1156;
  assign N1157 = sel_i[259] & sel_i[258];
  assign N1159 = N1158 & N1161;
  assign N1162 = sel_i[261] & sel_i[260];
  assign N1164 = N1163 & N1166;
  assign N1167 = sel_i[263] & sel_i[262];
  assign N1169 = N1168 & N1171;
  assign N1172 = sel_i[265] & sel_i[264];
  assign N1174 = N1173 & N1176;
  assign N1177 = sel_i[267] & sel_i[266];
  assign N1179 = N1178 & N1181;
  assign N1182 = sel_i[269] & sel_i[268];
  assign N1184 = N1183 & N1186;
  assign N1187 = sel_i[271] & sel_i[270];
  assign N1189 = N1188 & N1191;
  assign N1192 = sel_i[273] & sel_i[272];
  assign N1194 = N1193 & N1196;
  assign N1197 = sel_i[275] & sel_i[274];
  assign N1199 = N1198 & N1201;
  assign N1202 = sel_i[277] & sel_i[276];
  assign N1204 = N1203 & N1206;
  assign N1207 = sel_i[279] & sel_i[278];
  assign N1209 = N1208 & N1211;
  assign N1212 = sel_i[281] & sel_i[280];
  assign N1214 = N1213 & N1216;
  assign N1217 = sel_i[283] & sel_i[282];
  assign N1219 = N1218 & N1221;
  assign N1222 = sel_i[285] & sel_i[284];
  assign N1224 = N1223 & N1226;
  assign N1227 = sel_i[287] & sel_i[286];
  assign N1229 = N1228 & N1231;
  assign N1232 = sel_i[289] & sel_i[288];
  assign N1234 = N1233 & N1236;
  assign N1237 = sel_i[291] & sel_i[290];
  assign N1239 = N1238 & N1241;
  assign N1242 = sel_i[293] & sel_i[292];
  assign N1244 = N1243 & N1246;
  assign N1247 = sel_i[295] & sel_i[294];
  assign N1249 = N1248 & N1251;
  assign N1252 = sel_i[297] & sel_i[296];
  assign N1254 = N1253 & N1256;
  assign N1257 = sel_i[299] & sel_i[298];
  assign N1259 = N1258 & N1261;
  assign N1262 = sel_i[301] & sel_i[300];
  assign N1264 = N1263 & N1266;
  assign N1267 = sel_i[303] & sel_i[302];
  assign N1269 = N1268 & N1271;
  assign N1272 = sel_i[305] & sel_i[304];
  assign N1274 = N1273 & N1276;
  assign N1277 = sel_i[307] & sel_i[306];
  assign N1279 = N1278 & N1281;
  assign N1282 = sel_i[309] & sel_i[308];
  assign N1284 = N1283 & N1286;
  assign N1287 = sel_i[311] & sel_i[310];
  assign N1289 = N1288 & N1291;
  assign N1292 = sel_i[313] & sel_i[312];
  assign N1294 = N1293 & N1296;
  assign N1297 = sel_i[315] & sel_i[314];
  assign N1299 = N1298 & N1301;
  assign N1302 = sel_i[317] & sel_i[316];
  assign N1304 = N1303 & N1306;
  assign N1307 = sel_i[319] & sel_i[318];
  assign N1309 = N1308 & N1311;
  assign N1312 = sel_i[321] & sel_i[320];
  assign N1314 = N1313 & N1316;
  assign N1317 = sel_i[323] & sel_i[322];
  assign N1319 = N1318 & N1321;
  assign N1322 = sel_i[325] & sel_i[324];
  assign N1324 = N1323 & N1326;
  assign N1327 = sel_i[327] & sel_i[326];
  assign N1329 = N1328 & N1331;
  assign N1332 = sel_i[329] & sel_i[328];
  assign N1334 = N1333 & N1336;
  assign N1337 = sel_i[331] & sel_i[330];
  assign N1339 = N1338 & N1341;
  assign N1342 = sel_i[333] & sel_i[332];
  assign N1344 = N1343 & N1346;
  assign N1347 = sel_i[335] & sel_i[334];
  assign N1349 = N1348 & N1351;
  assign N1352 = sel_i[337] & sel_i[336];
  assign N1354 = N1353 & N1356;
  assign N1357 = sel_i[339] & sel_i[338];
  assign N1359 = N1358 & N1361;
  assign N1362 = sel_i[341] & sel_i[340];
  assign N1364 = N1363 & N1366;
  assign N1367 = sel_i[343] & sel_i[342];
  assign N1369 = N1368 & N1371;
  assign N1372 = sel_i[345] & sel_i[344];
  assign N1374 = N1373 & N1376;
  assign N1377 = sel_i[347] & sel_i[346];
  assign N1379 = N1378 & N1381;
  assign N1382 = sel_i[349] & sel_i[348];
  assign N1384 = N1383 & N1386;
  assign N1387 = sel_i[351] & sel_i[350];
  assign N1389 = N1388 & N1391;
  assign N1392 = sel_i[353] & sel_i[352];
  assign N1394 = N1393 & N1396;
  assign N1397 = sel_i[355] & sel_i[354];
  assign N1399 = N1398 & N1401;
  assign N1402 = sel_i[357] & sel_i[356];
  assign N1404 = N1403 & N1406;
  assign N1407 = sel_i[359] & sel_i[358];
  assign N1409 = N1408 & N1411;
  assign N1412 = sel_i[361] & sel_i[360];
  assign N1414 = N1413 & N1416;
  assign N1417 = sel_i[363] & sel_i[362];
  assign N1419 = N1418 & N1421;
  assign N1422 = sel_i[365] & sel_i[364];
  assign N1424 = N1423 & N1426;
  assign N1427 = sel_i[367] & sel_i[366];
  assign N1429 = N1428 & N1431;
  assign N1432 = sel_i[369] & sel_i[368];
  assign N1434 = N1433 & N1436;
  assign N1437 = sel_i[371] & sel_i[370];
  assign N1439 = N1438 & N1441;
  assign N1442 = sel_i[373] & sel_i[372];
  assign N1444 = N1443 & N1446;
  assign N1447 = sel_i[375] & sel_i[374];
  assign N1449 = N1448 & N1451;
  assign N1452 = sel_i[377] & sel_i[376];
  assign N1454 = N1453 & N1456;
  assign N1457 = sel_i[379] & sel_i[378];
  assign N1459 = N1458 & N1461;
  assign N1462 = sel_i[381] & sel_i[380];
  assign N1464 = N1463 & N1466;
  assign N1467 = sel_i[383] & sel_i[382];
  assign N1469 = N1468 & N1471;
  assign N1472 = sel_i[385] & sel_i[384];
  assign N1474 = N1473 & N1476;
  assign N1477 = sel_i[387] & sel_i[386];
  assign N1479 = N1478 & N1481;
  assign N1482 = sel_i[389] & sel_i[388];
  assign N1484 = N1483 & N1486;
  assign N1487 = sel_i[391] & sel_i[390];
  assign N1489 = N1488 & N1491;
  assign N1492 = sel_i[393] & sel_i[392];
  assign N1494 = N1493 & N1496;
  assign N1497 = sel_i[395] & sel_i[394];
  assign N1499 = N1498 & N1501;
  assign N1502 = sel_i[397] & sel_i[396];
  assign N1504 = N1503 & N1506;
  assign N1507 = sel_i[399] & sel_i[398];
  assign N1509 = N1508 & N1511;
  assign N1512 = sel_i[401] & sel_i[400];
  assign N1514 = N1513 & N1516;
  assign N1517 = sel_i[403] & sel_i[402];
  assign N1519 = N1518 & N1521;
  assign N1522 = sel_i[405] & sel_i[404];
  assign N1524 = N1523 & N1526;
  assign N1527 = sel_i[407] & sel_i[406];
  assign N1529 = N1528 & N1531;
  assign N1532 = sel_i[409] & sel_i[408];
  assign N1534 = N1533 & N1536;
  assign N1537 = sel_i[411] & sel_i[410];
  assign N1539 = N1538 & N1541;
  assign N1542 = sel_i[413] & sel_i[412];
  assign N1544 = N1543 & N1546;
  assign N1547 = sel_i[415] & sel_i[414];
  assign N1549 = N1548 & N1551;
  assign N1552 = sel_i[417] & sel_i[416];
  assign N1554 = N1553 & N1556;
  assign N1557 = sel_i[419] & sel_i[418];
  assign N1559 = N1558 & N1561;
  assign N1562 = sel_i[421] & sel_i[420];
  assign N1564 = N1563 & N1566;
  assign N1567 = sel_i[423] & sel_i[422];
  assign N1569 = N1568 & N1571;
  assign N1572 = sel_i[425] & sel_i[424];
  assign N1574 = N1573 & N1576;
  assign N1577 = sel_i[427] & sel_i[426];
  assign N1579 = N1578 & N1581;
  assign N1582 = sel_i[429] & sel_i[428];
  assign N1584 = N1583 & N1586;
  assign N1587 = sel_i[431] & sel_i[430];
  assign N1589 = N1588 & N1591;
  assign N1592 = sel_i[433] & sel_i[432];
  assign N1594 = N1593 & N1596;
  assign N1597 = sel_i[435] & sel_i[434];
  assign N1599 = N1598 & N1601;
  assign N1602 = sel_i[437] & sel_i[436];
  assign N1604 = N1603 & N1606;
  assign N1607 = sel_i[439] & sel_i[438];
  assign N1609 = N1608 & N1611;
  assign N1612 = sel_i[441] & sel_i[440];
  assign N1614 = N1613 & N1616;
  assign N1617 = sel_i[443] & sel_i[442];
  assign N1619 = N1618 & N1621;
  assign N1622 = sel_i[445] & sel_i[444];
  assign N1624 = N1623 & N1626;
  assign N1627 = sel_i[447] & sel_i[446];
  assign N1629 = N1628 & N1631;
  assign N1632 = sel_i[449] & sel_i[448];
  assign N1634 = N1633 & N1636;
  assign N1637 = sel_i[451] & sel_i[450];
  assign N1639 = N1638 & N1641;
  assign N1642 = sel_i[453] & sel_i[452];
  assign N1644 = N1643 & N1646;
  assign N1647 = sel_i[455] & sel_i[454];
  assign N1649 = N1648 & N1651;
  assign N1652 = sel_i[457] & sel_i[456];
  assign N1654 = N1653 & N1656;
  assign N1657 = sel_i[459] & sel_i[458];
  assign N1659 = N1658 & N1661;
  assign N1662 = sel_i[461] & sel_i[460];
  assign N1664 = N1663 & N1666;
  assign N1667 = sel_i[463] & sel_i[462];
  assign N1669 = N1668 & N1671;
  assign N1672 = sel_i[465] & sel_i[464];
  assign N1674 = N1673 & N1676;
  assign N1677 = sel_i[467] & sel_i[466];
  assign N1679 = N1678 & N1681;
  assign N1682 = sel_i[469] & sel_i[468];
  assign N1684 = N1683 & N1686;
  assign N1687 = sel_i[471] & sel_i[470];
  assign N1689 = N1688 & N1691;
  assign N1692 = sel_i[473] & sel_i[472];
  assign N1694 = N1693 & N1696;
  assign N1697 = sel_i[475] & sel_i[474];
  assign N1699 = N1698 & N1701;
  assign N1702 = sel_i[477] & sel_i[476];
  assign N1704 = N1703 & N1706;
  assign N1707 = sel_i[479] & sel_i[478];
  assign N1709 = N1708 & N1711;
  assign N1712 = sel_i[481] & sel_i[480];
  assign N1714 = N1713 & N1716;
  assign N1717 = sel_i[483] & sel_i[482];
  assign N1719 = N1718 & N1721;
  assign N1722 = sel_i[485] & sel_i[484];
  assign N1724 = N1723 & N1726;
  assign N1727 = sel_i[487] & sel_i[486];
  assign N1729 = N1728 & N1731;
  assign N1732 = sel_i[489] & sel_i[488];
  assign N1734 = N1733 & N1736;
  assign N1737 = sel_i[491] & sel_i[490];
  assign N1739 = N1738 & N1741;
  assign N1742 = sel_i[493] & sel_i[492];
  assign N1744 = N1743 & N1746;
  assign N1747 = sel_i[495] & sel_i[494];
  assign N1749 = N1748 & N1751;
  assign N1752 = sel_i[497] & sel_i[496];
  assign N1754 = N1753 & N1756;
  assign N1757 = sel_i[499] & sel_i[498];
  assign N1759 = N1758 & N1761;
  assign N1762 = sel_i[501] & sel_i[500];
  assign N1764 = N1763 & N1766;
  assign N1767 = sel_i[503] & sel_i[502];
  assign N1769 = N1768 & N1771;
  assign N1772 = sel_i[505] & sel_i[504];
  assign N1774 = N1773 & N1776;
  assign N1777 = sel_i[507] & sel_i[506];
  assign N1779 = N1778 & N1781;
  assign N1782 = sel_i[509] & sel_i[508];
  assign N1784 = N1783 & N1786;
  assign N1787 = sel_i[511] & sel_i[510];
  assign N1789 = N1788 & N1791;
  assign N516 = ~sel_i[0];
  assign N521 = ~sel_i[2];
  assign N526 = ~sel_i[4];
  assign N531 = ~sel_i[6];
  assign N536 = ~sel_i[8];
  assign N541 = ~sel_i[10];
  assign N546 = ~sel_i[12];
  assign N551 = ~sel_i[14];
  assign N556 = ~sel_i[16];
  assign N561 = ~sel_i[18];
  assign N566 = ~sel_i[20];
  assign N571 = ~sel_i[22];
  assign N576 = ~sel_i[24];
  assign N581 = ~sel_i[26];
  assign N586 = ~sel_i[28];
  assign N591 = ~sel_i[30];
  assign N596 = ~sel_i[32];
  assign N601 = ~sel_i[34];
  assign N606 = ~sel_i[36];
  assign N611 = ~sel_i[38];
  assign N616 = ~sel_i[40];
  assign N621 = ~sel_i[42];
  assign N626 = ~sel_i[44];
  assign N631 = ~sel_i[46];
  assign N636 = ~sel_i[48];
  assign N641 = ~sel_i[50];
  assign N646 = ~sel_i[52];
  assign N651 = ~sel_i[54];
  assign N656 = ~sel_i[56];
  assign N661 = ~sel_i[58];
  assign N666 = ~sel_i[60];
  assign N671 = ~sel_i[62];
  assign N676 = ~sel_i[64];
  assign N681 = ~sel_i[66];
  assign N686 = ~sel_i[68];
  assign N691 = ~sel_i[70];
  assign N696 = ~sel_i[72];
  assign N701 = ~sel_i[74];
  assign N706 = ~sel_i[76];
  assign N711 = ~sel_i[78];
  assign N716 = ~sel_i[80];
  assign N721 = ~sel_i[82];
  assign N726 = ~sel_i[84];
  assign N731 = ~sel_i[86];
  assign N736 = ~sel_i[88];
  assign N741 = ~sel_i[90];
  assign N746 = ~sel_i[92];
  assign N751 = ~sel_i[94];
  assign N756 = ~sel_i[96];
  assign N761 = ~sel_i[98];
  assign N766 = ~sel_i[100];
  assign N771 = ~sel_i[102];
  assign N776 = ~sel_i[104];
  assign N781 = ~sel_i[106];
  assign N786 = ~sel_i[108];
  assign N791 = ~sel_i[110];
  assign N796 = ~sel_i[112];
  assign N801 = ~sel_i[114];
  assign N806 = ~sel_i[116];
  assign N811 = ~sel_i[118];
  assign N816 = ~sel_i[120];
  assign N821 = ~sel_i[122];
  assign N826 = ~sel_i[124];
  assign N831 = ~sel_i[126];
  assign N836 = ~sel_i[128];
  assign N841 = ~sel_i[130];
  assign N846 = ~sel_i[132];
  assign N851 = ~sel_i[134];
  assign N856 = ~sel_i[136];
  assign N861 = ~sel_i[138];
  assign N866 = ~sel_i[140];
  assign N871 = ~sel_i[142];
  assign N876 = ~sel_i[144];
  assign N881 = ~sel_i[146];
  assign N886 = ~sel_i[148];
  assign N891 = ~sel_i[150];
  assign N896 = ~sel_i[152];
  assign N901 = ~sel_i[154];
  assign N906 = ~sel_i[156];
  assign N911 = ~sel_i[158];
  assign N916 = ~sel_i[160];
  assign N921 = ~sel_i[162];
  assign N926 = ~sel_i[164];
  assign N931 = ~sel_i[166];
  assign N936 = ~sel_i[168];
  assign N941 = ~sel_i[170];
  assign N946 = ~sel_i[172];
  assign N951 = ~sel_i[174];
  assign N956 = ~sel_i[176];
  assign N961 = ~sel_i[178];
  assign N966 = ~sel_i[180];
  assign N971 = ~sel_i[182];
  assign N976 = ~sel_i[184];
  assign N981 = ~sel_i[186];
  assign N986 = ~sel_i[188];
  assign N991 = ~sel_i[190];
  assign N996 = ~sel_i[192];
  assign N1001 = ~sel_i[194];
  assign N1006 = ~sel_i[196];
  assign N1011 = ~sel_i[198];
  assign N1016 = ~sel_i[200];
  assign N1021 = ~sel_i[202];
  assign N1026 = ~sel_i[204];
  assign N1031 = ~sel_i[206];
  assign N1036 = ~sel_i[208];
  assign N1041 = ~sel_i[210];
  assign N1046 = ~sel_i[212];
  assign N1051 = ~sel_i[214];
  assign N1056 = ~sel_i[216];
  assign N1061 = ~sel_i[218];
  assign N1066 = ~sel_i[220];
  assign N1071 = ~sel_i[222];
  assign N1076 = ~sel_i[224];
  assign N1081 = ~sel_i[226];
  assign N1086 = ~sel_i[228];
  assign N1091 = ~sel_i[230];
  assign N1096 = ~sel_i[232];
  assign N1101 = ~sel_i[234];
  assign N1106 = ~sel_i[236];
  assign N1111 = ~sel_i[238];
  assign N1116 = ~sel_i[240];
  assign N1121 = ~sel_i[242];
  assign N1126 = ~sel_i[244];
  assign N1131 = ~sel_i[246];
  assign N1136 = ~sel_i[248];
  assign N1141 = ~sel_i[250];
  assign N1146 = ~sel_i[252];
  assign N1151 = ~sel_i[254];
  assign N1156 = ~sel_i[256];
  assign N1161 = ~sel_i[258];
  assign N1166 = ~sel_i[260];
  assign N1171 = ~sel_i[262];
  assign N1176 = ~sel_i[264];
  assign N1181 = ~sel_i[266];
  assign N1186 = ~sel_i[268];
  assign N1191 = ~sel_i[270];
  assign N1196 = ~sel_i[272];
  assign N1201 = ~sel_i[274];
  assign N1206 = ~sel_i[276];
  assign N1211 = ~sel_i[278];
  assign N1216 = ~sel_i[280];
  assign N1221 = ~sel_i[282];
  assign N1226 = ~sel_i[284];
  assign N1231 = ~sel_i[286];
  assign N1236 = ~sel_i[288];
  assign N1241 = ~sel_i[290];
  assign N1246 = ~sel_i[292];
  assign N1251 = ~sel_i[294];
  assign N1256 = ~sel_i[296];
  assign N1261 = ~sel_i[298];
  assign N1266 = ~sel_i[300];
  assign N1271 = ~sel_i[302];
  assign N1276 = ~sel_i[304];
  assign N1281 = ~sel_i[306];
  assign N1286 = ~sel_i[308];
  assign N1291 = ~sel_i[310];
  assign N1296 = ~sel_i[312];
  assign N1301 = ~sel_i[314];
  assign N1306 = ~sel_i[316];
  assign N1311 = ~sel_i[318];
  assign N1316 = ~sel_i[320];
  assign N1321 = ~sel_i[322];
  assign N1326 = ~sel_i[324];
  assign N1331 = ~sel_i[326];
  assign N1336 = ~sel_i[328];
  assign N1341 = ~sel_i[330];
  assign N1346 = ~sel_i[332];
  assign N1351 = ~sel_i[334];
  assign N1356 = ~sel_i[336];
  assign N1361 = ~sel_i[338];
  assign N1366 = ~sel_i[340];
  assign N1371 = ~sel_i[342];
  assign N1376 = ~sel_i[344];
  assign N1381 = ~sel_i[346];
  assign N1386 = ~sel_i[348];
  assign N1391 = ~sel_i[350];
  assign N1396 = ~sel_i[352];
  assign N1401 = ~sel_i[354];
  assign N1406 = ~sel_i[356];
  assign N1411 = ~sel_i[358];
  assign N1416 = ~sel_i[360];
  assign N1421 = ~sel_i[362];
  assign N1426 = ~sel_i[364];
  assign N1431 = ~sel_i[366];
  assign N1436 = ~sel_i[368];
  assign N1441 = ~sel_i[370];
  assign N1446 = ~sel_i[372];
  assign N1451 = ~sel_i[374];
  assign N1456 = ~sel_i[376];
  assign N1461 = ~sel_i[378];
  assign N1466 = ~sel_i[380];
  assign N1471 = ~sel_i[382];
  assign N1476 = ~sel_i[384];
  assign N1481 = ~sel_i[386];
  assign N1486 = ~sel_i[388];
  assign N1491 = ~sel_i[390];
  assign N1496 = ~sel_i[392];
  assign N1501 = ~sel_i[394];
  assign N1506 = ~sel_i[396];
  assign N1511 = ~sel_i[398];
  assign N1516 = ~sel_i[400];
  assign N1521 = ~sel_i[402];
  assign N1526 = ~sel_i[404];
  assign N1531 = ~sel_i[406];
  assign N1536 = ~sel_i[408];
  assign N1541 = ~sel_i[410];
  assign N1546 = ~sel_i[412];
  assign N1551 = ~sel_i[414];
  assign N1556 = ~sel_i[416];
  assign N1561 = ~sel_i[418];
  assign N1566 = ~sel_i[420];
  assign N1571 = ~sel_i[422];
  assign N1576 = ~sel_i[424];
  assign N1581 = ~sel_i[426];
  assign N1586 = ~sel_i[428];
  assign N1591 = ~sel_i[430];
  assign N1596 = ~sel_i[432];
  assign N1601 = ~sel_i[434];
  assign N1606 = ~sel_i[436];
  assign N1611 = ~sel_i[438];
  assign N1616 = ~sel_i[440];
  assign N1621 = ~sel_i[442];
  assign N1626 = ~sel_i[444];
  assign N1631 = ~sel_i[446];
  assign N1636 = ~sel_i[448];
  assign N1641 = ~sel_i[450];
  assign N1646 = ~sel_i[452];
  assign N1651 = ~sel_i[454];
  assign N1656 = ~sel_i[456];
  assign N1661 = ~sel_i[458];
  assign N1666 = ~sel_i[460];
  assign N1671 = ~sel_i[462];
  assign N1676 = ~sel_i[464];
  assign N1681 = ~sel_i[466];
  assign N1686 = ~sel_i[468];
  assign N1691 = ~sel_i[470];
  assign N1696 = ~sel_i[472];
  assign N1701 = ~sel_i[474];
  assign N1706 = ~sel_i[476];
  assign N1711 = ~sel_i[478];
  assign N1716 = ~sel_i[480];
  assign N1721 = ~sel_i[482];
  assign N1726 = ~sel_i[484];
  assign N1731 = ~sel_i[486];
  assign N1736 = ~sel_i[488];
  assign N1741 = ~sel_i[490];
  assign N1746 = ~sel_i[492];
  assign N1751 = ~sel_i[494];
  assign N1756 = ~sel_i[496];
  assign N1761 = ~sel_i[498];
  assign N1766 = ~sel_i[500];
  assign N1771 = ~sel_i[502];
  assign N1776 = ~sel_i[504];
  assign N1781 = ~sel_i[506];
  assign N1786 = ~sel_i[508];
  assign N1791 = ~sel_i[510];
  assign { r_n_0__31_, r_n_0__30_, r_n_0__29_, r_n_0__28_, r_n_0__27_, r_n_0__26_, r_n_0__25_, r_n_0__24_, r_n_0__23_, r_n_0__22_, r_n_0__21_, r_n_0__20_, r_n_0__19_, r_n_0__18_, r_n_0__17_, r_n_0__16_, r_n_0__15_, r_n_0__14_, r_n_0__13_, r_n_0__12_, r_n_0__11_, r_n_0__10_, r_n_0__9_, r_n_0__8_, r_n_0__7_, r_n_0__6_, r_n_0__5_, r_n_0__4_, r_n_0__3_, r_n_0__2_, r_n_0__1_, r_n_0__0_ } = (N0)? { r_1__31_, r_1__30_, r_1__29_, r_1__28_, r_1__27_, r_1__26_, r_1__25_, r_1__24_, r_1__23_, r_1__22_, r_1__21_, r_1__20_, r_1__19_, r_1__18_, r_1__17_, r_1__16_, r_1__15_, r_1__14_, r_1__13_, r_1__12_, r_1__11_, r_1__10_, r_1__9_, r_1__8_, r_1__7_, r_1__6_, r_1__5_, r_1__4_, r_1__3_, r_1__2_, r_1__1_, r_1__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                    (N1)? data_i : 1'b0;
  assign N0 = sel_i[0];
  assign N1 = N516;
  assign { r_n_1__31_, r_n_1__30_, r_n_1__29_, r_n_1__28_, r_n_1__27_, r_n_1__26_, r_n_1__25_, r_n_1__24_, r_n_1__23_, r_n_1__22_, r_n_1__21_, r_n_1__20_, r_n_1__19_, r_n_1__18_, r_n_1__17_, r_n_1__16_, r_n_1__15_, r_n_1__14_, r_n_1__13_, r_n_1__12_, r_n_1__11_, r_n_1__10_, r_n_1__9_, r_n_1__8_, r_n_1__7_, r_n_1__6_, r_n_1__5_, r_n_1__4_, r_n_1__3_, r_n_1__2_, r_n_1__1_, r_n_1__0_ } = (N2)? { r_2__31_, r_2__30_, r_2__29_, r_2__28_, r_2__27_, r_2__26_, r_2__25_, r_2__24_, r_2__23_, r_2__22_, r_2__21_, r_2__20_, r_2__19_, r_2__18_, r_2__17_, r_2__16_, r_2__15_, r_2__14_, r_2__13_, r_2__12_, r_2__11_, r_2__10_, r_2__9_, r_2__8_, r_2__7_, r_2__6_, r_2__5_, r_2__4_, r_2__3_, r_2__2_, r_2__1_, r_2__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                    (N3)? data_i : 1'b0;
  assign N2 = sel_i[2];
  assign N3 = N521;
  assign { r_n_2__31_, r_n_2__30_, r_n_2__29_, r_n_2__28_, r_n_2__27_, r_n_2__26_, r_n_2__25_, r_n_2__24_, r_n_2__23_, r_n_2__22_, r_n_2__21_, r_n_2__20_, r_n_2__19_, r_n_2__18_, r_n_2__17_, r_n_2__16_, r_n_2__15_, r_n_2__14_, r_n_2__13_, r_n_2__12_, r_n_2__11_, r_n_2__10_, r_n_2__9_, r_n_2__8_, r_n_2__7_, r_n_2__6_, r_n_2__5_, r_n_2__4_, r_n_2__3_, r_n_2__2_, r_n_2__1_, r_n_2__0_ } = (N4)? { r_3__31_, r_3__30_, r_3__29_, r_3__28_, r_3__27_, r_3__26_, r_3__25_, r_3__24_, r_3__23_, r_3__22_, r_3__21_, r_3__20_, r_3__19_, r_3__18_, r_3__17_, r_3__16_, r_3__15_, r_3__14_, r_3__13_, r_3__12_, r_3__11_, r_3__10_, r_3__9_, r_3__8_, r_3__7_, r_3__6_, r_3__5_, r_3__4_, r_3__3_, r_3__2_, r_3__1_, r_3__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                    (N5)? data_i : 1'b0;
  assign N4 = sel_i[4];
  assign N5 = N526;
  assign { r_n_3__31_, r_n_3__30_, r_n_3__29_, r_n_3__28_, r_n_3__27_, r_n_3__26_, r_n_3__25_, r_n_3__24_, r_n_3__23_, r_n_3__22_, r_n_3__21_, r_n_3__20_, r_n_3__19_, r_n_3__18_, r_n_3__17_, r_n_3__16_, r_n_3__15_, r_n_3__14_, r_n_3__13_, r_n_3__12_, r_n_3__11_, r_n_3__10_, r_n_3__9_, r_n_3__8_, r_n_3__7_, r_n_3__6_, r_n_3__5_, r_n_3__4_, r_n_3__3_, r_n_3__2_, r_n_3__1_, r_n_3__0_ } = (N6)? { r_4__31_, r_4__30_, r_4__29_, r_4__28_, r_4__27_, r_4__26_, r_4__25_, r_4__24_, r_4__23_, r_4__22_, r_4__21_, r_4__20_, r_4__19_, r_4__18_, r_4__17_, r_4__16_, r_4__15_, r_4__14_, r_4__13_, r_4__12_, r_4__11_, r_4__10_, r_4__9_, r_4__8_, r_4__7_, r_4__6_, r_4__5_, r_4__4_, r_4__3_, r_4__2_, r_4__1_, r_4__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                    (N7)? data_i : 1'b0;
  assign N6 = sel_i[6];
  assign N7 = N531;
  assign { r_n_4__31_, r_n_4__30_, r_n_4__29_, r_n_4__28_, r_n_4__27_, r_n_4__26_, r_n_4__25_, r_n_4__24_, r_n_4__23_, r_n_4__22_, r_n_4__21_, r_n_4__20_, r_n_4__19_, r_n_4__18_, r_n_4__17_, r_n_4__16_, r_n_4__15_, r_n_4__14_, r_n_4__13_, r_n_4__12_, r_n_4__11_, r_n_4__10_, r_n_4__9_, r_n_4__8_, r_n_4__7_, r_n_4__6_, r_n_4__5_, r_n_4__4_, r_n_4__3_, r_n_4__2_, r_n_4__1_, r_n_4__0_ } = (N8)? { r_5__31_, r_5__30_, r_5__29_, r_5__28_, r_5__27_, r_5__26_, r_5__25_, r_5__24_, r_5__23_, r_5__22_, r_5__21_, r_5__20_, r_5__19_, r_5__18_, r_5__17_, r_5__16_, r_5__15_, r_5__14_, r_5__13_, r_5__12_, r_5__11_, r_5__10_, r_5__9_, r_5__8_, r_5__7_, r_5__6_, r_5__5_, r_5__4_, r_5__3_, r_5__2_, r_5__1_, r_5__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                    (N9)? data_i : 1'b0;
  assign N8 = sel_i[8];
  assign N9 = N536;
  assign { r_n_5__31_, r_n_5__30_, r_n_5__29_, r_n_5__28_, r_n_5__27_, r_n_5__26_, r_n_5__25_, r_n_5__24_, r_n_5__23_, r_n_5__22_, r_n_5__21_, r_n_5__20_, r_n_5__19_, r_n_5__18_, r_n_5__17_, r_n_5__16_, r_n_5__15_, r_n_5__14_, r_n_5__13_, r_n_5__12_, r_n_5__11_, r_n_5__10_, r_n_5__9_, r_n_5__8_, r_n_5__7_, r_n_5__6_, r_n_5__5_, r_n_5__4_, r_n_5__3_, r_n_5__2_, r_n_5__1_, r_n_5__0_ } = (N10)? { r_6__31_, r_6__30_, r_6__29_, r_6__28_, r_6__27_, r_6__26_, r_6__25_, r_6__24_, r_6__23_, r_6__22_, r_6__21_, r_6__20_, r_6__19_, r_6__18_, r_6__17_, r_6__16_, r_6__15_, r_6__14_, r_6__13_, r_6__12_, r_6__11_, r_6__10_, r_6__9_, r_6__8_, r_6__7_, r_6__6_, r_6__5_, r_6__4_, r_6__3_, r_6__2_, r_6__1_, r_6__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                    (N11)? data_i : 1'b0;
  assign N10 = sel_i[10];
  assign N11 = N541;
  assign { r_n_6__31_, r_n_6__30_, r_n_6__29_, r_n_6__28_, r_n_6__27_, r_n_6__26_, r_n_6__25_, r_n_6__24_, r_n_6__23_, r_n_6__22_, r_n_6__21_, r_n_6__20_, r_n_6__19_, r_n_6__18_, r_n_6__17_, r_n_6__16_, r_n_6__15_, r_n_6__14_, r_n_6__13_, r_n_6__12_, r_n_6__11_, r_n_6__10_, r_n_6__9_, r_n_6__8_, r_n_6__7_, r_n_6__6_, r_n_6__5_, r_n_6__4_, r_n_6__3_, r_n_6__2_, r_n_6__1_, r_n_6__0_ } = (N12)? { r_7__31_, r_7__30_, r_7__29_, r_7__28_, r_7__27_, r_7__26_, r_7__25_, r_7__24_, r_7__23_, r_7__22_, r_7__21_, r_7__20_, r_7__19_, r_7__18_, r_7__17_, r_7__16_, r_7__15_, r_7__14_, r_7__13_, r_7__12_, r_7__11_, r_7__10_, r_7__9_, r_7__8_, r_7__7_, r_7__6_, r_7__5_, r_7__4_, r_7__3_, r_7__2_, r_7__1_, r_7__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                    (N13)? data_i : 1'b0;
  assign N12 = sel_i[12];
  assign N13 = N546;
  assign { r_n_7__31_, r_n_7__30_, r_n_7__29_, r_n_7__28_, r_n_7__27_, r_n_7__26_, r_n_7__25_, r_n_7__24_, r_n_7__23_, r_n_7__22_, r_n_7__21_, r_n_7__20_, r_n_7__19_, r_n_7__18_, r_n_7__17_, r_n_7__16_, r_n_7__15_, r_n_7__14_, r_n_7__13_, r_n_7__12_, r_n_7__11_, r_n_7__10_, r_n_7__9_, r_n_7__8_, r_n_7__7_, r_n_7__6_, r_n_7__5_, r_n_7__4_, r_n_7__3_, r_n_7__2_, r_n_7__1_, r_n_7__0_ } = (N14)? { r_8__31_, r_8__30_, r_8__29_, r_8__28_, r_8__27_, r_8__26_, r_8__25_, r_8__24_, r_8__23_, r_8__22_, r_8__21_, r_8__20_, r_8__19_, r_8__18_, r_8__17_, r_8__16_, r_8__15_, r_8__14_, r_8__13_, r_8__12_, r_8__11_, r_8__10_, r_8__9_, r_8__8_, r_8__7_, r_8__6_, r_8__5_, r_8__4_, r_8__3_, r_8__2_, r_8__1_, r_8__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                    (N15)? data_i : 1'b0;
  assign N14 = sel_i[14];
  assign N15 = N551;
  assign { r_n_8__31_, r_n_8__30_, r_n_8__29_, r_n_8__28_, r_n_8__27_, r_n_8__26_, r_n_8__25_, r_n_8__24_, r_n_8__23_, r_n_8__22_, r_n_8__21_, r_n_8__20_, r_n_8__19_, r_n_8__18_, r_n_8__17_, r_n_8__16_, r_n_8__15_, r_n_8__14_, r_n_8__13_, r_n_8__12_, r_n_8__11_, r_n_8__10_, r_n_8__9_, r_n_8__8_, r_n_8__7_, r_n_8__6_, r_n_8__5_, r_n_8__4_, r_n_8__3_, r_n_8__2_, r_n_8__1_, r_n_8__0_ } = (N16)? { r_9__31_, r_9__30_, r_9__29_, r_9__28_, r_9__27_, r_9__26_, r_9__25_, r_9__24_, r_9__23_, r_9__22_, r_9__21_, r_9__20_, r_9__19_, r_9__18_, r_9__17_, r_9__16_, r_9__15_, r_9__14_, r_9__13_, r_9__12_, r_9__11_, r_9__10_, r_9__9_, r_9__8_, r_9__7_, r_9__6_, r_9__5_, r_9__4_, r_9__3_, r_9__2_, r_9__1_, r_9__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                    (N17)? data_i : 1'b0;
  assign N16 = sel_i[16];
  assign N17 = N556;
  assign { r_n_9__31_, r_n_9__30_, r_n_9__29_, r_n_9__28_, r_n_9__27_, r_n_9__26_, r_n_9__25_, r_n_9__24_, r_n_9__23_, r_n_9__22_, r_n_9__21_, r_n_9__20_, r_n_9__19_, r_n_9__18_, r_n_9__17_, r_n_9__16_, r_n_9__15_, r_n_9__14_, r_n_9__13_, r_n_9__12_, r_n_9__11_, r_n_9__10_, r_n_9__9_, r_n_9__8_, r_n_9__7_, r_n_9__6_, r_n_9__5_, r_n_9__4_, r_n_9__3_, r_n_9__2_, r_n_9__1_, r_n_9__0_ } = (N18)? { r_10__31_, r_10__30_, r_10__29_, r_10__28_, r_10__27_, r_10__26_, r_10__25_, r_10__24_, r_10__23_, r_10__22_, r_10__21_, r_10__20_, r_10__19_, r_10__18_, r_10__17_, r_10__16_, r_10__15_, r_10__14_, r_10__13_, r_10__12_, r_10__11_, r_10__10_, r_10__9_, r_10__8_, r_10__7_, r_10__6_, r_10__5_, r_10__4_, r_10__3_, r_10__2_, r_10__1_, r_10__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                    (N19)? data_i : 1'b0;
  assign N18 = sel_i[18];
  assign N19 = N561;
  assign { r_n_10__31_, r_n_10__30_, r_n_10__29_, r_n_10__28_, r_n_10__27_, r_n_10__26_, r_n_10__25_, r_n_10__24_, r_n_10__23_, r_n_10__22_, r_n_10__21_, r_n_10__20_, r_n_10__19_, r_n_10__18_, r_n_10__17_, r_n_10__16_, r_n_10__15_, r_n_10__14_, r_n_10__13_, r_n_10__12_, r_n_10__11_, r_n_10__10_, r_n_10__9_, r_n_10__8_, r_n_10__7_, r_n_10__6_, r_n_10__5_, r_n_10__4_, r_n_10__3_, r_n_10__2_, r_n_10__1_, r_n_10__0_ } = (N20)? { r_11__31_, r_11__30_, r_11__29_, r_11__28_, r_11__27_, r_11__26_, r_11__25_, r_11__24_, r_11__23_, r_11__22_, r_11__21_, r_11__20_, r_11__19_, r_11__18_, r_11__17_, r_11__16_, r_11__15_, r_11__14_, r_11__13_, r_11__12_, r_11__11_, r_11__10_, r_11__9_, r_11__8_, r_11__7_, r_11__6_, r_11__5_, r_11__4_, r_11__3_, r_11__2_, r_11__1_, r_11__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N21)? data_i : 1'b0;
  assign N20 = sel_i[20];
  assign N21 = N566;
  assign { r_n_11__31_, r_n_11__30_, r_n_11__29_, r_n_11__28_, r_n_11__27_, r_n_11__26_, r_n_11__25_, r_n_11__24_, r_n_11__23_, r_n_11__22_, r_n_11__21_, r_n_11__20_, r_n_11__19_, r_n_11__18_, r_n_11__17_, r_n_11__16_, r_n_11__15_, r_n_11__14_, r_n_11__13_, r_n_11__12_, r_n_11__11_, r_n_11__10_, r_n_11__9_, r_n_11__8_, r_n_11__7_, r_n_11__6_, r_n_11__5_, r_n_11__4_, r_n_11__3_, r_n_11__2_, r_n_11__1_, r_n_11__0_ } = (N22)? { r_12__31_, r_12__30_, r_12__29_, r_12__28_, r_12__27_, r_12__26_, r_12__25_, r_12__24_, r_12__23_, r_12__22_, r_12__21_, r_12__20_, r_12__19_, r_12__18_, r_12__17_, r_12__16_, r_12__15_, r_12__14_, r_12__13_, r_12__12_, r_12__11_, r_12__10_, r_12__9_, r_12__8_, r_12__7_, r_12__6_, r_12__5_, r_12__4_, r_12__3_, r_12__2_, r_12__1_, r_12__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N23)? data_i : 1'b0;
  assign N22 = sel_i[22];
  assign N23 = N571;
  assign { r_n_12__31_, r_n_12__30_, r_n_12__29_, r_n_12__28_, r_n_12__27_, r_n_12__26_, r_n_12__25_, r_n_12__24_, r_n_12__23_, r_n_12__22_, r_n_12__21_, r_n_12__20_, r_n_12__19_, r_n_12__18_, r_n_12__17_, r_n_12__16_, r_n_12__15_, r_n_12__14_, r_n_12__13_, r_n_12__12_, r_n_12__11_, r_n_12__10_, r_n_12__9_, r_n_12__8_, r_n_12__7_, r_n_12__6_, r_n_12__5_, r_n_12__4_, r_n_12__3_, r_n_12__2_, r_n_12__1_, r_n_12__0_ } = (N24)? { r_13__31_, r_13__30_, r_13__29_, r_13__28_, r_13__27_, r_13__26_, r_13__25_, r_13__24_, r_13__23_, r_13__22_, r_13__21_, r_13__20_, r_13__19_, r_13__18_, r_13__17_, r_13__16_, r_13__15_, r_13__14_, r_13__13_, r_13__12_, r_13__11_, r_13__10_, r_13__9_, r_13__8_, r_13__7_, r_13__6_, r_13__5_, r_13__4_, r_13__3_, r_13__2_, r_13__1_, r_13__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N25)? data_i : 1'b0;
  assign N24 = sel_i[24];
  assign N25 = N576;
  assign { r_n_13__31_, r_n_13__30_, r_n_13__29_, r_n_13__28_, r_n_13__27_, r_n_13__26_, r_n_13__25_, r_n_13__24_, r_n_13__23_, r_n_13__22_, r_n_13__21_, r_n_13__20_, r_n_13__19_, r_n_13__18_, r_n_13__17_, r_n_13__16_, r_n_13__15_, r_n_13__14_, r_n_13__13_, r_n_13__12_, r_n_13__11_, r_n_13__10_, r_n_13__9_, r_n_13__8_, r_n_13__7_, r_n_13__6_, r_n_13__5_, r_n_13__4_, r_n_13__3_, r_n_13__2_, r_n_13__1_, r_n_13__0_ } = (N26)? { r_14__31_, r_14__30_, r_14__29_, r_14__28_, r_14__27_, r_14__26_, r_14__25_, r_14__24_, r_14__23_, r_14__22_, r_14__21_, r_14__20_, r_14__19_, r_14__18_, r_14__17_, r_14__16_, r_14__15_, r_14__14_, r_14__13_, r_14__12_, r_14__11_, r_14__10_, r_14__9_, r_14__8_, r_14__7_, r_14__6_, r_14__5_, r_14__4_, r_14__3_, r_14__2_, r_14__1_, r_14__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N27)? data_i : 1'b0;
  assign N26 = sel_i[26];
  assign N27 = N581;
  assign { r_n_14__31_, r_n_14__30_, r_n_14__29_, r_n_14__28_, r_n_14__27_, r_n_14__26_, r_n_14__25_, r_n_14__24_, r_n_14__23_, r_n_14__22_, r_n_14__21_, r_n_14__20_, r_n_14__19_, r_n_14__18_, r_n_14__17_, r_n_14__16_, r_n_14__15_, r_n_14__14_, r_n_14__13_, r_n_14__12_, r_n_14__11_, r_n_14__10_, r_n_14__9_, r_n_14__8_, r_n_14__7_, r_n_14__6_, r_n_14__5_, r_n_14__4_, r_n_14__3_, r_n_14__2_, r_n_14__1_, r_n_14__0_ } = (N28)? { r_15__31_, r_15__30_, r_15__29_, r_15__28_, r_15__27_, r_15__26_, r_15__25_, r_15__24_, r_15__23_, r_15__22_, r_15__21_, r_15__20_, r_15__19_, r_15__18_, r_15__17_, r_15__16_, r_15__15_, r_15__14_, r_15__13_, r_15__12_, r_15__11_, r_15__10_, r_15__9_, r_15__8_, r_15__7_, r_15__6_, r_15__5_, r_15__4_, r_15__3_, r_15__2_, r_15__1_, r_15__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N29)? data_i : 1'b0;
  assign N28 = sel_i[28];
  assign N29 = N586;
  assign { r_n_15__31_, r_n_15__30_, r_n_15__29_, r_n_15__28_, r_n_15__27_, r_n_15__26_, r_n_15__25_, r_n_15__24_, r_n_15__23_, r_n_15__22_, r_n_15__21_, r_n_15__20_, r_n_15__19_, r_n_15__18_, r_n_15__17_, r_n_15__16_, r_n_15__15_, r_n_15__14_, r_n_15__13_, r_n_15__12_, r_n_15__11_, r_n_15__10_, r_n_15__9_, r_n_15__8_, r_n_15__7_, r_n_15__6_, r_n_15__5_, r_n_15__4_, r_n_15__3_, r_n_15__2_, r_n_15__1_, r_n_15__0_ } = (N30)? { r_16__31_, r_16__30_, r_16__29_, r_16__28_, r_16__27_, r_16__26_, r_16__25_, r_16__24_, r_16__23_, r_16__22_, r_16__21_, r_16__20_, r_16__19_, r_16__18_, r_16__17_, r_16__16_, r_16__15_, r_16__14_, r_16__13_, r_16__12_, r_16__11_, r_16__10_, r_16__9_, r_16__8_, r_16__7_, r_16__6_, r_16__5_, r_16__4_, r_16__3_, r_16__2_, r_16__1_, r_16__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N31)? data_i : 1'b0;
  assign N30 = sel_i[30];
  assign N31 = N591;
  assign { r_n_16__31_, r_n_16__30_, r_n_16__29_, r_n_16__28_, r_n_16__27_, r_n_16__26_, r_n_16__25_, r_n_16__24_, r_n_16__23_, r_n_16__22_, r_n_16__21_, r_n_16__20_, r_n_16__19_, r_n_16__18_, r_n_16__17_, r_n_16__16_, r_n_16__15_, r_n_16__14_, r_n_16__13_, r_n_16__12_, r_n_16__11_, r_n_16__10_, r_n_16__9_, r_n_16__8_, r_n_16__7_, r_n_16__6_, r_n_16__5_, r_n_16__4_, r_n_16__3_, r_n_16__2_, r_n_16__1_, r_n_16__0_ } = (N32)? { r_17__31_, r_17__30_, r_17__29_, r_17__28_, r_17__27_, r_17__26_, r_17__25_, r_17__24_, r_17__23_, r_17__22_, r_17__21_, r_17__20_, r_17__19_, r_17__18_, r_17__17_, r_17__16_, r_17__15_, r_17__14_, r_17__13_, r_17__12_, r_17__11_, r_17__10_, r_17__9_, r_17__8_, r_17__7_, r_17__6_, r_17__5_, r_17__4_, r_17__3_, r_17__2_, r_17__1_, r_17__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N33)? data_i : 1'b0;
  assign N32 = sel_i[32];
  assign N33 = N596;
  assign { r_n_17__31_, r_n_17__30_, r_n_17__29_, r_n_17__28_, r_n_17__27_, r_n_17__26_, r_n_17__25_, r_n_17__24_, r_n_17__23_, r_n_17__22_, r_n_17__21_, r_n_17__20_, r_n_17__19_, r_n_17__18_, r_n_17__17_, r_n_17__16_, r_n_17__15_, r_n_17__14_, r_n_17__13_, r_n_17__12_, r_n_17__11_, r_n_17__10_, r_n_17__9_, r_n_17__8_, r_n_17__7_, r_n_17__6_, r_n_17__5_, r_n_17__4_, r_n_17__3_, r_n_17__2_, r_n_17__1_, r_n_17__0_ } = (N34)? { r_18__31_, r_18__30_, r_18__29_, r_18__28_, r_18__27_, r_18__26_, r_18__25_, r_18__24_, r_18__23_, r_18__22_, r_18__21_, r_18__20_, r_18__19_, r_18__18_, r_18__17_, r_18__16_, r_18__15_, r_18__14_, r_18__13_, r_18__12_, r_18__11_, r_18__10_, r_18__9_, r_18__8_, r_18__7_, r_18__6_, r_18__5_, r_18__4_, r_18__3_, r_18__2_, r_18__1_, r_18__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N35)? data_i : 1'b0;
  assign N34 = sel_i[34];
  assign N35 = N601;
  assign { r_n_18__31_, r_n_18__30_, r_n_18__29_, r_n_18__28_, r_n_18__27_, r_n_18__26_, r_n_18__25_, r_n_18__24_, r_n_18__23_, r_n_18__22_, r_n_18__21_, r_n_18__20_, r_n_18__19_, r_n_18__18_, r_n_18__17_, r_n_18__16_, r_n_18__15_, r_n_18__14_, r_n_18__13_, r_n_18__12_, r_n_18__11_, r_n_18__10_, r_n_18__9_, r_n_18__8_, r_n_18__7_, r_n_18__6_, r_n_18__5_, r_n_18__4_, r_n_18__3_, r_n_18__2_, r_n_18__1_, r_n_18__0_ } = (N36)? { r_19__31_, r_19__30_, r_19__29_, r_19__28_, r_19__27_, r_19__26_, r_19__25_, r_19__24_, r_19__23_, r_19__22_, r_19__21_, r_19__20_, r_19__19_, r_19__18_, r_19__17_, r_19__16_, r_19__15_, r_19__14_, r_19__13_, r_19__12_, r_19__11_, r_19__10_, r_19__9_, r_19__8_, r_19__7_, r_19__6_, r_19__5_, r_19__4_, r_19__3_, r_19__2_, r_19__1_, r_19__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N37)? data_i : 1'b0;
  assign N36 = sel_i[36];
  assign N37 = N606;
  assign { r_n_19__31_, r_n_19__30_, r_n_19__29_, r_n_19__28_, r_n_19__27_, r_n_19__26_, r_n_19__25_, r_n_19__24_, r_n_19__23_, r_n_19__22_, r_n_19__21_, r_n_19__20_, r_n_19__19_, r_n_19__18_, r_n_19__17_, r_n_19__16_, r_n_19__15_, r_n_19__14_, r_n_19__13_, r_n_19__12_, r_n_19__11_, r_n_19__10_, r_n_19__9_, r_n_19__8_, r_n_19__7_, r_n_19__6_, r_n_19__5_, r_n_19__4_, r_n_19__3_, r_n_19__2_, r_n_19__1_, r_n_19__0_ } = (N38)? { r_20__31_, r_20__30_, r_20__29_, r_20__28_, r_20__27_, r_20__26_, r_20__25_, r_20__24_, r_20__23_, r_20__22_, r_20__21_, r_20__20_, r_20__19_, r_20__18_, r_20__17_, r_20__16_, r_20__15_, r_20__14_, r_20__13_, r_20__12_, r_20__11_, r_20__10_, r_20__9_, r_20__8_, r_20__7_, r_20__6_, r_20__5_, r_20__4_, r_20__3_, r_20__2_, r_20__1_, r_20__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N39)? data_i : 1'b0;
  assign N38 = sel_i[38];
  assign N39 = N611;
  assign { r_n_20__31_, r_n_20__30_, r_n_20__29_, r_n_20__28_, r_n_20__27_, r_n_20__26_, r_n_20__25_, r_n_20__24_, r_n_20__23_, r_n_20__22_, r_n_20__21_, r_n_20__20_, r_n_20__19_, r_n_20__18_, r_n_20__17_, r_n_20__16_, r_n_20__15_, r_n_20__14_, r_n_20__13_, r_n_20__12_, r_n_20__11_, r_n_20__10_, r_n_20__9_, r_n_20__8_, r_n_20__7_, r_n_20__6_, r_n_20__5_, r_n_20__4_, r_n_20__3_, r_n_20__2_, r_n_20__1_, r_n_20__0_ } = (N40)? { r_21__31_, r_21__30_, r_21__29_, r_21__28_, r_21__27_, r_21__26_, r_21__25_, r_21__24_, r_21__23_, r_21__22_, r_21__21_, r_21__20_, r_21__19_, r_21__18_, r_21__17_, r_21__16_, r_21__15_, r_21__14_, r_21__13_, r_21__12_, r_21__11_, r_21__10_, r_21__9_, r_21__8_, r_21__7_, r_21__6_, r_21__5_, r_21__4_, r_21__3_, r_21__2_, r_21__1_, r_21__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N41)? data_i : 1'b0;
  assign N40 = sel_i[40];
  assign N41 = N616;
  assign { r_n_21__31_, r_n_21__30_, r_n_21__29_, r_n_21__28_, r_n_21__27_, r_n_21__26_, r_n_21__25_, r_n_21__24_, r_n_21__23_, r_n_21__22_, r_n_21__21_, r_n_21__20_, r_n_21__19_, r_n_21__18_, r_n_21__17_, r_n_21__16_, r_n_21__15_, r_n_21__14_, r_n_21__13_, r_n_21__12_, r_n_21__11_, r_n_21__10_, r_n_21__9_, r_n_21__8_, r_n_21__7_, r_n_21__6_, r_n_21__5_, r_n_21__4_, r_n_21__3_, r_n_21__2_, r_n_21__1_, r_n_21__0_ } = (N42)? { r_22__31_, r_22__30_, r_22__29_, r_22__28_, r_22__27_, r_22__26_, r_22__25_, r_22__24_, r_22__23_, r_22__22_, r_22__21_, r_22__20_, r_22__19_, r_22__18_, r_22__17_, r_22__16_, r_22__15_, r_22__14_, r_22__13_, r_22__12_, r_22__11_, r_22__10_, r_22__9_, r_22__8_, r_22__7_, r_22__6_, r_22__5_, r_22__4_, r_22__3_, r_22__2_, r_22__1_, r_22__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N43)? data_i : 1'b0;
  assign N42 = sel_i[42];
  assign N43 = N621;
  assign { r_n_22__31_, r_n_22__30_, r_n_22__29_, r_n_22__28_, r_n_22__27_, r_n_22__26_, r_n_22__25_, r_n_22__24_, r_n_22__23_, r_n_22__22_, r_n_22__21_, r_n_22__20_, r_n_22__19_, r_n_22__18_, r_n_22__17_, r_n_22__16_, r_n_22__15_, r_n_22__14_, r_n_22__13_, r_n_22__12_, r_n_22__11_, r_n_22__10_, r_n_22__9_, r_n_22__8_, r_n_22__7_, r_n_22__6_, r_n_22__5_, r_n_22__4_, r_n_22__3_, r_n_22__2_, r_n_22__1_, r_n_22__0_ } = (N44)? { r_23__31_, r_23__30_, r_23__29_, r_23__28_, r_23__27_, r_23__26_, r_23__25_, r_23__24_, r_23__23_, r_23__22_, r_23__21_, r_23__20_, r_23__19_, r_23__18_, r_23__17_, r_23__16_, r_23__15_, r_23__14_, r_23__13_, r_23__12_, r_23__11_, r_23__10_, r_23__9_, r_23__8_, r_23__7_, r_23__6_, r_23__5_, r_23__4_, r_23__3_, r_23__2_, r_23__1_, r_23__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N45)? data_i : 1'b0;
  assign N44 = sel_i[44];
  assign N45 = N626;
  assign { r_n_23__31_, r_n_23__30_, r_n_23__29_, r_n_23__28_, r_n_23__27_, r_n_23__26_, r_n_23__25_, r_n_23__24_, r_n_23__23_, r_n_23__22_, r_n_23__21_, r_n_23__20_, r_n_23__19_, r_n_23__18_, r_n_23__17_, r_n_23__16_, r_n_23__15_, r_n_23__14_, r_n_23__13_, r_n_23__12_, r_n_23__11_, r_n_23__10_, r_n_23__9_, r_n_23__8_, r_n_23__7_, r_n_23__6_, r_n_23__5_, r_n_23__4_, r_n_23__3_, r_n_23__2_, r_n_23__1_, r_n_23__0_ } = (N46)? { r_24__31_, r_24__30_, r_24__29_, r_24__28_, r_24__27_, r_24__26_, r_24__25_, r_24__24_, r_24__23_, r_24__22_, r_24__21_, r_24__20_, r_24__19_, r_24__18_, r_24__17_, r_24__16_, r_24__15_, r_24__14_, r_24__13_, r_24__12_, r_24__11_, r_24__10_, r_24__9_, r_24__8_, r_24__7_, r_24__6_, r_24__5_, r_24__4_, r_24__3_, r_24__2_, r_24__1_, r_24__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N47)? data_i : 1'b0;
  assign N46 = sel_i[46];
  assign N47 = N631;
  assign { r_n_24__31_, r_n_24__30_, r_n_24__29_, r_n_24__28_, r_n_24__27_, r_n_24__26_, r_n_24__25_, r_n_24__24_, r_n_24__23_, r_n_24__22_, r_n_24__21_, r_n_24__20_, r_n_24__19_, r_n_24__18_, r_n_24__17_, r_n_24__16_, r_n_24__15_, r_n_24__14_, r_n_24__13_, r_n_24__12_, r_n_24__11_, r_n_24__10_, r_n_24__9_, r_n_24__8_, r_n_24__7_, r_n_24__6_, r_n_24__5_, r_n_24__4_, r_n_24__3_, r_n_24__2_, r_n_24__1_, r_n_24__0_ } = (N48)? { r_25__31_, r_25__30_, r_25__29_, r_25__28_, r_25__27_, r_25__26_, r_25__25_, r_25__24_, r_25__23_, r_25__22_, r_25__21_, r_25__20_, r_25__19_, r_25__18_, r_25__17_, r_25__16_, r_25__15_, r_25__14_, r_25__13_, r_25__12_, r_25__11_, r_25__10_, r_25__9_, r_25__8_, r_25__7_, r_25__6_, r_25__5_, r_25__4_, r_25__3_, r_25__2_, r_25__1_, r_25__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N49)? data_i : 1'b0;
  assign N48 = sel_i[48];
  assign N49 = N636;
  assign { r_n_25__31_, r_n_25__30_, r_n_25__29_, r_n_25__28_, r_n_25__27_, r_n_25__26_, r_n_25__25_, r_n_25__24_, r_n_25__23_, r_n_25__22_, r_n_25__21_, r_n_25__20_, r_n_25__19_, r_n_25__18_, r_n_25__17_, r_n_25__16_, r_n_25__15_, r_n_25__14_, r_n_25__13_, r_n_25__12_, r_n_25__11_, r_n_25__10_, r_n_25__9_, r_n_25__8_, r_n_25__7_, r_n_25__6_, r_n_25__5_, r_n_25__4_, r_n_25__3_, r_n_25__2_, r_n_25__1_, r_n_25__0_ } = (N50)? { r_26__31_, r_26__30_, r_26__29_, r_26__28_, r_26__27_, r_26__26_, r_26__25_, r_26__24_, r_26__23_, r_26__22_, r_26__21_, r_26__20_, r_26__19_, r_26__18_, r_26__17_, r_26__16_, r_26__15_, r_26__14_, r_26__13_, r_26__12_, r_26__11_, r_26__10_, r_26__9_, r_26__8_, r_26__7_, r_26__6_, r_26__5_, r_26__4_, r_26__3_, r_26__2_, r_26__1_, r_26__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N51)? data_i : 1'b0;
  assign N50 = sel_i[50];
  assign N51 = N641;
  assign { r_n_26__31_, r_n_26__30_, r_n_26__29_, r_n_26__28_, r_n_26__27_, r_n_26__26_, r_n_26__25_, r_n_26__24_, r_n_26__23_, r_n_26__22_, r_n_26__21_, r_n_26__20_, r_n_26__19_, r_n_26__18_, r_n_26__17_, r_n_26__16_, r_n_26__15_, r_n_26__14_, r_n_26__13_, r_n_26__12_, r_n_26__11_, r_n_26__10_, r_n_26__9_, r_n_26__8_, r_n_26__7_, r_n_26__6_, r_n_26__5_, r_n_26__4_, r_n_26__3_, r_n_26__2_, r_n_26__1_, r_n_26__0_ } = (N52)? { r_27__31_, r_27__30_, r_27__29_, r_27__28_, r_27__27_, r_27__26_, r_27__25_, r_27__24_, r_27__23_, r_27__22_, r_27__21_, r_27__20_, r_27__19_, r_27__18_, r_27__17_, r_27__16_, r_27__15_, r_27__14_, r_27__13_, r_27__12_, r_27__11_, r_27__10_, r_27__9_, r_27__8_, r_27__7_, r_27__6_, r_27__5_, r_27__4_, r_27__3_, r_27__2_, r_27__1_, r_27__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N53)? data_i : 1'b0;
  assign N52 = sel_i[52];
  assign N53 = N646;
  assign { r_n_27__31_, r_n_27__30_, r_n_27__29_, r_n_27__28_, r_n_27__27_, r_n_27__26_, r_n_27__25_, r_n_27__24_, r_n_27__23_, r_n_27__22_, r_n_27__21_, r_n_27__20_, r_n_27__19_, r_n_27__18_, r_n_27__17_, r_n_27__16_, r_n_27__15_, r_n_27__14_, r_n_27__13_, r_n_27__12_, r_n_27__11_, r_n_27__10_, r_n_27__9_, r_n_27__8_, r_n_27__7_, r_n_27__6_, r_n_27__5_, r_n_27__4_, r_n_27__3_, r_n_27__2_, r_n_27__1_, r_n_27__0_ } = (N54)? { r_28__31_, r_28__30_, r_28__29_, r_28__28_, r_28__27_, r_28__26_, r_28__25_, r_28__24_, r_28__23_, r_28__22_, r_28__21_, r_28__20_, r_28__19_, r_28__18_, r_28__17_, r_28__16_, r_28__15_, r_28__14_, r_28__13_, r_28__12_, r_28__11_, r_28__10_, r_28__9_, r_28__8_, r_28__7_, r_28__6_, r_28__5_, r_28__4_, r_28__3_, r_28__2_, r_28__1_, r_28__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N55)? data_i : 1'b0;
  assign N54 = sel_i[54];
  assign N55 = N651;
  assign { r_n_28__31_, r_n_28__30_, r_n_28__29_, r_n_28__28_, r_n_28__27_, r_n_28__26_, r_n_28__25_, r_n_28__24_, r_n_28__23_, r_n_28__22_, r_n_28__21_, r_n_28__20_, r_n_28__19_, r_n_28__18_, r_n_28__17_, r_n_28__16_, r_n_28__15_, r_n_28__14_, r_n_28__13_, r_n_28__12_, r_n_28__11_, r_n_28__10_, r_n_28__9_, r_n_28__8_, r_n_28__7_, r_n_28__6_, r_n_28__5_, r_n_28__4_, r_n_28__3_, r_n_28__2_, r_n_28__1_, r_n_28__0_ } = (N56)? { r_29__31_, r_29__30_, r_29__29_, r_29__28_, r_29__27_, r_29__26_, r_29__25_, r_29__24_, r_29__23_, r_29__22_, r_29__21_, r_29__20_, r_29__19_, r_29__18_, r_29__17_, r_29__16_, r_29__15_, r_29__14_, r_29__13_, r_29__12_, r_29__11_, r_29__10_, r_29__9_, r_29__8_, r_29__7_, r_29__6_, r_29__5_, r_29__4_, r_29__3_, r_29__2_, r_29__1_, r_29__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N57)? data_i : 1'b0;
  assign N56 = sel_i[56];
  assign N57 = N656;
  assign { r_n_29__31_, r_n_29__30_, r_n_29__29_, r_n_29__28_, r_n_29__27_, r_n_29__26_, r_n_29__25_, r_n_29__24_, r_n_29__23_, r_n_29__22_, r_n_29__21_, r_n_29__20_, r_n_29__19_, r_n_29__18_, r_n_29__17_, r_n_29__16_, r_n_29__15_, r_n_29__14_, r_n_29__13_, r_n_29__12_, r_n_29__11_, r_n_29__10_, r_n_29__9_, r_n_29__8_, r_n_29__7_, r_n_29__6_, r_n_29__5_, r_n_29__4_, r_n_29__3_, r_n_29__2_, r_n_29__1_, r_n_29__0_ } = (N58)? { r_30__31_, r_30__30_, r_30__29_, r_30__28_, r_30__27_, r_30__26_, r_30__25_, r_30__24_, r_30__23_, r_30__22_, r_30__21_, r_30__20_, r_30__19_, r_30__18_, r_30__17_, r_30__16_, r_30__15_, r_30__14_, r_30__13_, r_30__12_, r_30__11_, r_30__10_, r_30__9_, r_30__8_, r_30__7_, r_30__6_, r_30__5_, r_30__4_, r_30__3_, r_30__2_, r_30__1_, r_30__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N59)? data_i : 1'b0;
  assign N58 = sel_i[58];
  assign N59 = N661;
  assign { r_n_30__31_, r_n_30__30_, r_n_30__29_, r_n_30__28_, r_n_30__27_, r_n_30__26_, r_n_30__25_, r_n_30__24_, r_n_30__23_, r_n_30__22_, r_n_30__21_, r_n_30__20_, r_n_30__19_, r_n_30__18_, r_n_30__17_, r_n_30__16_, r_n_30__15_, r_n_30__14_, r_n_30__13_, r_n_30__12_, r_n_30__11_, r_n_30__10_, r_n_30__9_, r_n_30__8_, r_n_30__7_, r_n_30__6_, r_n_30__5_, r_n_30__4_, r_n_30__3_, r_n_30__2_, r_n_30__1_, r_n_30__0_ } = (N60)? { r_31__31_, r_31__30_, r_31__29_, r_31__28_, r_31__27_, r_31__26_, r_31__25_, r_31__24_, r_31__23_, r_31__22_, r_31__21_, r_31__20_, r_31__19_, r_31__18_, r_31__17_, r_31__16_, r_31__15_, r_31__14_, r_31__13_, r_31__12_, r_31__11_, r_31__10_, r_31__9_, r_31__8_, r_31__7_, r_31__6_, r_31__5_, r_31__4_, r_31__3_, r_31__2_, r_31__1_, r_31__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N61)? data_i : 1'b0;
  assign N60 = sel_i[60];
  assign N61 = N666;
  assign { r_n_31__31_, r_n_31__30_, r_n_31__29_, r_n_31__28_, r_n_31__27_, r_n_31__26_, r_n_31__25_, r_n_31__24_, r_n_31__23_, r_n_31__22_, r_n_31__21_, r_n_31__20_, r_n_31__19_, r_n_31__18_, r_n_31__17_, r_n_31__16_, r_n_31__15_, r_n_31__14_, r_n_31__13_, r_n_31__12_, r_n_31__11_, r_n_31__10_, r_n_31__9_, r_n_31__8_, r_n_31__7_, r_n_31__6_, r_n_31__5_, r_n_31__4_, r_n_31__3_, r_n_31__2_, r_n_31__1_, r_n_31__0_ } = (N62)? { r_32__31_, r_32__30_, r_32__29_, r_32__28_, r_32__27_, r_32__26_, r_32__25_, r_32__24_, r_32__23_, r_32__22_, r_32__21_, r_32__20_, r_32__19_, r_32__18_, r_32__17_, r_32__16_, r_32__15_, r_32__14_, r_32__13_, r_32__12_, r_32__11_, r_32__10_, r_32__9_, r_32__8_, r_32__7_, r_32__6_, r_32__5_, r_32__4_, r_32__3_, r_32__2_, r_32__1_, r_32__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N63)? data_i : 1'b0;
  assign N62 = sel_i[62];
  assign N63 = N671;
  assign { r_n_32__31_, r_n_32__30_, r_n_32__29_, r_n_32__28_, r_n_32__27_, r_n_32__26_, r_n_32__25_, r_n_32__24_, r_n_32__23_, r_n_32__22_, r_n_32__21_, r_n_32__20_, r_n_32__19_, r_n_32__18_, r_n_32__17_, r_n_32__16_, r_n_32__15_, r_n_32__14_, r_n_32__13_, r_n_32__12_, r_n_32__11_, r_n_32__10_, r_n_32__9_, r_n_32__8_, r_n_32__7_, r_n_32__6_, r_n_32__5_, r_n_32__4_, r_n_32__3_, r_n_32__2_, r_n_32__1_, r_n_32__0_ } = (N64)? { r_33__31_, r_33__30_, r_33__29_, r_33__28_, r_33__27_, r_33__26_, r_33__25_, r_33__24_, r_33__23_, r_33__22_, r_33__21_, r_33__20_, r_33__19_, r_33__18_, r_33__17_, r_33__16_, r_33__15_, r_33__14_, r_33__13_, r_33__12_, r_33__11_, r_33__10_, r_33__9_, r_33__8_, r_33__7_, r_33__6_, r_33__5_, r_33__4_, r_33__3_, r_33__2_, r_33__1_, r_33__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N65)? data_i : 1'b0;
  assign N64 = sel_i[64];
  assign N65 = N676;
  assign { r_n_33__31_, r_n_33__30_, r_n_33__29_, r_n_33__28_, r_n_33__27_, r_n_33__26_, r_n_33__25_, r_n_33__24_, r_n_33__23_, r_n_33__22_, r_n_33__21_, r_n_33__20_, r_n_33__19_, r_n_33__18_, r_n_33__17_, r_n_33__16_, r_n_33__15_, r_n_33__14_, r_n_33__13_, r_n_33__12_, r_n_33__11_, r_n_33__10_, r_n_33__9_, r_n_33__8_, r_n_33__7_, r_n_33__6_, r_n_33__5_, r_n_33__4_, r_n_33__3_, r_n_33__2_, r_n_33__1_, r_n_33__0_ } = (N66)? { r_34__31_, r_34__30_, r_34__29_, r_34__28_, r_34__27_, r_34__26_, r_34__25_, r_34__24_, r_34__23_, r_34__22_, r_34__21_, r_34__20_, r_34__19_, r_34__18_, r_34__17_, r_34__16_, r_34__15_, r_34__14_, r_34__13_, r_34__12_, r_34__11_, r_34__10_, r_34__9_, r_34__8_, r_34__7_, r_34__6_, r_34__5_, r_34__4_, r_34__3_, r_34__2_, r_34__1_, r_34__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N67)? data_i : 1'b0;
  assign N66 = sel_i[66];
  assign N67 = N681;
  assign { r_n_34__31_, r_n_34__30_, r_n_34__29_, r_n_34__28_, r_n_34__27_, r_n_34__26_, r_n_34__25_, r_n_34__24_, r_n_34__23_, r_n_34__22_, r_n_34__21_, r_n_34__20_, r_n_34__19_, r_n_34__18_, r_n_34__17_, r_n_34__16_, r_n_34__15_, r_n_34__14_, r_n_34__13_, r_n_34__12_, r_n_34__11_, r_n_34__10_, r_n_34__9_, r_n_34__8_, r_n_34__7_, r_n_34__6_, r_n_34__5_, r_n_34__4_, r_n_34__3_, r_n_34__2_, r_n_34__1_, r_n_34__0_ } = (N68)? { r_35__31_, r_35__30_, r_35__29_, r_35__28_, r_35__27_, r_35__26_, r_35__25_, r_35__24_, r_35__23_, r_35__22_, r_35__21_, r_35__20_, r_35__19_, r_35__18_, r_35__17_, r_35__16_, r_35__15_, r_35__14_, r_35__13_, r_35__12_, r_35__11_, r_35__10_, r_35__9_, r_35__8_, r_35__7_, r_35__6_, r_35__5_, r_35__4_, r_35__3_, r_35__2_, r_35__1_, r_35__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N69)? data_i : 1'b0;
  assign N68 = sel_i[68];
  assign N69 = N686;
  assign { r_n_35__31_, r_n_35__30_, r_n_35__29_, r_n_35__28_, r_n_35__27_, r_n_35__26_, r_n_35__25_, r_n_35__24_, r_n_35__23_, r_n_35__22_, r_n_35__21_, r_n_35__20_, r_n_35__19_, r_n_35__18_, r_n_35__17_, r_n_35__16_, r_n_35__15_, r_n_35__14_, r_n_35__13_, r_n_35__12_, r_n_35__11_, r_n_35__10_, r_n_35__9_, r_n_35__8_, r_n_35__7_, r_n_35__6_, r_n_35__5_, r_n_35__4_, r_n_35__3_, r_n_35__2_, r_n_35__1_, r_n_35__0_ } = (N70)? { r_36__31_, r_36__30_, r_36__29_, r_36__28_, r_36__27_, r_36__26_, r_36__25_, r_36__24_, r_36__23_, r_36__22_, r_36__21_, r_36__20_, r_36__19_, r_36__18_, r_36__17_, r_36__16_, r_36__15_, r_36__14_, r_36__13_, r_36__12_, r_36__11_, r_36__10_, r_36__9_, r_36__8_, r_36__7_, r_36__6_, r_36__5_, r_36__4_, r_36__3_, r_36__2_, r_36__1_, r_36__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N71)? data_i : 1'b0;
  assign N70 = sel_i[70];
  assign N71 = N691;
  assign { r_n_36__31_, r_n_36__30_, r_n_36__29_, r_n_36__28_, r_n_36__27_, r_n_36__26_, r_n_36__25_, r_n_36__24_, r_n_36__23_, r_n_36__22_, r_n_36__21_, r_n_36__20_, r_n_36__19_, r_n_36__18_, r_n_36__17_, r_n_36__16_, r_n_36__15_, r_n_36__14_, r_n_36__13_, r_n_36__12_, r_n_36__11_, r_n_36__10_, r_n_36__9_, r_n_36__8_, r_n_36__7_, r_n_36__6_, r_n_36__5_, r_n_36__4_, r_n_36__3_, r_n_36__2_, r_n_36__1_, r_n_36__0_ } = (N72)? { r_37__31_, r_37__30_, r_37__29_, r_37__28_, r_37__27_, r_37__26_, r_37__25_, r_37__24_, r_37__23_, r_37__22_, r_37__21_, r_37__20_, r_37__19_, r_37__18_, r_37__17_, r_37__16_, r_37__15_, r_37__14_, r_37__13_, r_37__12_, r_37__11_, r_37__10_, r_37__9_, r_37__8_, r_37__7_, r_37__6_, r_37__5_, r_37__4_, r_37__3_, r_37__2_, r_37__1_, r_37__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N73)? data_i : 1'b0;
  assign N72 = sel_i[72];
  assign N73 = N696;
  assign { r_n_37__31_, r_n_37__30_, r_n_37__29_, r_n_37__28_, r_n_37__27_, r_n_37__26_, r_n_37__25_, r_n_37__24_, r_n_37__23_, r_n_37__22_, r_n_37__21_, r_n_37__20_, r_n_37__19_, r_n_37__18_, r_n_37__17_, r_n_37__16_, r_n_37__15_, r_n_37__14_, r_n_37__13_, r_n_37__12_, r_n_37__11_, r_n_37__10_, r_n_37__9_, r_n_37__8_, r_n_37__7_, r_n_37__6_, r_n_37__5_, r_n_37__4_, r_n_37__3_, r_n_37__2_, r_n_37__1_, r_n_37__0_ } = (N74)? { r_38__31_, r_38__30_, r_38__29_, r_38__28_, r_38__27_, r_38__26_, r_38__25_, r_38__24_, r_38__23_, r_38__22_, r_38__21_, r_38__20_, r_38__19_, r_38__18_, r_38__17_, r_38__16_, r_38__15_, r_38__14_, r_38__13_, r_38__12_, r_38__11_, r_38__10_, r_38__9_, r_38__8_, r_38__7_, r_38__6_, r_38__5_, r_38__4_, r_38__3_, r_38__2_, r_38__1_, r_38__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N75)? data_i : 1'b0;
  assign N74 = sel_i[74];
  assign N75 = N701;
  assign { r_n_38__31_, r_n_38__30_, r_n_38__29_, r_n_38__28_, r_n_38__27_, r_n_38__26_, r_n_38__25_, r_n_38__24_, r_n_38__23_, r_n_38__22_, r_n_38__21_, r_n_38__20_, r_n_38__19_, r_n_38__18_, r_n_38__17_, r_n_38__16_, r_n_38__15_, r_n_38__14_, r_n_38__13_, r_n_38__12_, r_n_38__11_, r_n_38__10_, r_n_38__9_, r_n_38__8_, r_n_38__7_, r_n_38__6_, r_n_38__5_, r_n_38__4_, r_n_38__3_, r_n_38__2_, r_n_38__1_, r_n_38__0_ } = (N76)? { r_39__31_, r_39__30_, r_39__29_, r_39__28_, r_39__27_, r_39__26_, r_39__25_, r_39__24_, r_39__23_, r_39__22_, r_39__21_, r_39__20_, r_39__19_, r_39__18_, r_39__17_, r_39__16_, r_39__15_, r_39__14_, r_39__13_, r_39__12_, r_39__11_, r_39__10_, r_39__9_, r_39__8_, r_39__7_, r_39__6_, r_39__5_, r_39__4_, r_39__3_, r_39__2_, r_39__1_, r_39__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N77)? data_i : 1'b0;
  assign N76 = sel_i[76];
  assign N77 = N706;
  assign { r_n_39__31_, r_n_39__30_, r_n_39__29_, r_n_39__28_, r_n_39__27_, r_n_39__26_, r_n_39__25_, r_n_39__24_, r_n_39__23_, r_n_39__22_, r_n_39__21_, r_n_39__20_, r_n_39__19_, r_n_39__18_, r_n_39__17_, r_n_39__16_, r_n_39__15_, r_n_39__14_, r_n_39__13_, r_n_39__12_, r_n_39__11_, r_n_39__10_, r_n_39__9_, r_n_39__8_, r_n_39__7_, r_n_39__6_, r_n_39__5_, r_n_39__4_, r_n_39__3_, r_n_39__2_, r_n_39__1_, r_n_39__0_ } = (N78)? { r_40__31_, r_40__30_, r_40__29_, r_40__28_, r_40__27_, r_40__26_, r_40__25_, r_40__24_, r_40__23_, r_40__22_, r_40__21_, r_40__20_, r_40__19_, r_40__18_, r_40__17_, r_40__16_, r_40__15_, r_40__14_, r_40__13_, r_40__12_, r_40__11_, r_40__10_, r_40__9_, r_40__8_, r_40__7_, r_40__6_, r_40__5_, r_40__4_, r_40__3_, r_40__2_, r_40__1_, r_40__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N79)? data_i : 1'b0;
  assign N78 = sel_i[78];
  assign N79 = N711;
  assign { r_n_40__31_, r_n_40__30_, r_n_40__29_, r_n_40__28_, r_n_40__27_, r_n_40__26_, r_n_40__25_, r_n_40__24_, r_n_40__23_, r_n_40__22_, r_n_40__21_, r_n_40__20_, r_n_40__19_, r_n_40__18_, r_n_40__17_, r_n_40__16_, r_n_40__15_, r_n_40__14_, r_n_40__13_, r_n_40__12_, r_n_40__11_, r_n_40__10_, r_n_40__9_, r_n_40__8_, r_n_40__7_, r_n_40__6_, r_n_40__5_, r_n_40__4_, r_n_40__3_, r_n_40__2_, r_n_40__1_, r_n_40__0_ } = (N80)? { r_41__31_, r_41__30_, r_41__29_, r_41__28_, r_41__27_, r_41__26_, r_41__25_, r_41__24_, r_41__23_, r_41__22_, r_41__21_, r_41__20_, r_41__19_, r_41__18_, r_41__17_, r_41__16_, r_41__15_, r_41__14_, r_41__13_, r_41__12_, r_41__11_, r_41__10_, r_41__9_, r_41__8_, r_41__7_, r_41__6_, r_41__5_, r_41__4_, r_41__3_, r_41__2_, r_41__1_, r_41__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N81)? data_i : 1'b0;
  assign N80 = sel_i[80];
  assign N81 = N716;
  assign { r_n_41__31_, r_n_41__30_, r_n_41__29_, r_n_41__28_, r_n_41__27_, r_n_41__26_, r_n_41__25_, r_n_41__24_, r_n_41__23_, r_n_41__22_, r_n_41__21_, r_n_41__20_, r_n_41__19_, r_n_41__18_, r_n_41__17_, r_n_41__16_, r_n_41__15_, r_n_41__14_, r_n_41__13_, r_n_41__12_, r_n_41__11_, r_n_41__10_, r_n_41__9_, r_n_41__8_, r_n_41__7_, r_n_41__6_, r_n_41__5_, r_n_41__4_, r_n_41__3_, r_n_41__2_, r_n_41__1_, r_n_41__0_ } = (N82)? { r_42__31_, r_42__30_, r_42__29_, r_42__28_, r_42__27_, r_42__26_, r_42__25_, r_42__24_, r_42__23_, r_42__22_, r_42__21_, r_42__20_, r_42__19_, r_42__18_, r_42__17_, r_42__16_, r_42__15_, r_42__14_, r_42__13_, r_42__12_, r_42__11_, r_42__10_, r_42__9_, r_42__8_, r_42__7_, r_42__6_, r_42__5_, r_42__4_, r_42__3_, r_42__2_, r_42__1_, r_42__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N83)? data_i : 1'b0;
  assign N82 = sel_i[82];
  assign N83 = N721;
  assign { r_n_42__31_, r_n_42__30_, r_n_42__29_, r_n_42__28_, r_n_42__27_, r_n_42__26_, r_n_42__25_, r_n_42__24_, r_n_42__23_, r_n_42__22_, r_n_42__21_, r_n_42__20_, r_n_42__19_, r_n_42__18_, r_n_42__17_, r_n_42__16_, r_n_42__15_, r_n_42__14_, r_n_42__13_, r_n_42__12_, r_n_42__11_, r_n_42__10_, r_n_42__9_, r_n_42__8_, r_n_42__7_, r_n_42__6_, r_n_42__5_, r_n_42__4_, r_n_42__3_, r_n_42__2_, r_n_42__1_, r_n_42__0_ } = (N84)? { r_43__31_, r_43__30_, r_43__29_, r_43__28_, r_43__27_, r_43__26_, r_43__25_, r_43__24_, r_43__23_, r_43__22_, r_43__21_, r_43__20_, r_43__19_, r_43__18_, r_43__17_, r_43__16_, r_43__15_, r_43__14_, r_43__13_, r_43__12_, r_43__11_, r_43__10_, r_43__9_, r_43__8_, r_43__7_, r_43__6_, r_43__5_, r_43__4_, r_43__3_, r_43__2_, r_43__1_, r_43__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N85)? data_i : 1'b0;
  assign N84 = sel_i[84];
  assign N85 = N726;
  assign { r_n_43__31_, r_n_43__30_, r_n_43__29_, r_n_43__28_, r_n_43__27_, r_n_43__26_, r_n_43__25_, r_n_43__24_, r_n_43__23_, r_n_43__22_, r_n_43__21_, r_n_43__20_, r_n_43__19_, r_n_43__18_, r_n_43__17_, r_n_43__16_, r_n_43__15_, r_n_43__14_, r_n_43__13_, r_n_43__12_, r_n_43__11_, r_n_43__10_, r_n_43__9_, r_n_43__8_, r_n_43__7_, r_n_43__6_, r_n_43__5_, r_n_43__4_, r_n_43__3_, r_n_43__2_, r_n_43__1_, r_n_43__0_ } = (N86)? { r_44__31_, r_44__30_, r_44__29_, r_44__28_, r_44__27_, r_44__26_, r_44__25_, r_44__24_, r_44__23_, r_44__22_, r_44__21_, r_44__20_, r_44__19_, r_44__18_, r_44__17_, r_44__16_, r_44__15_, r_44__14_, r_44__13_, r_44__12_, r_44__11_, r_44__10_, r_44__9_, r_44__8_, r_44__7_, r_44__6_, r_44__5_, r_44__4_, r_44__3_, r_44__2_, r_44__1_, r_44__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N87)? data_i : 1'b0;
  assign N86 = sel_i[86];
  assign N87 = N731;
  assign { r_n_44__31_, r_n_44__30_, r_n_44__29_, r_n_44__28_, r_n_44__27_, r_n_44__26_, r_n_44__25_, r_n_44__24_, r_n_44__23_, r_n_44__22_, r_n_44__21_, r_n_44__20_, r_n_44__19_, r_n_44__18_, r_n_44__17_, r_n_44__16_, r_n_44__15_, r_n_44__14_, r_n_44__13_, r_n_44__12_, r_n_44__11_, r_n_44__10_, r_n_44__9_, r_n_44__8_, r_n_44__7_, r_n_44__6_, r_n_44__5_, r_n_44__4_, r_n_44__3_, r_n_44__2_, r_n_44__1_, r_n_44__0_ } = (N88)? { r_45__31_, r_45__30_, r_45__29_, r_45__28_, r_45__27_, r_45__26_, r_45__25_, r_45__24_, r_45__23_, r_45__22_, r_45__21_, r_45__20_, r_45__19_, r_45__18_, r_45__17_, r_45__16_, r_45__15_, r_45__14_, r_45__13_, r_45__12_, r_45__11_, r_45__10_, r_45__9_, r_45__8_, r_45__7_, r_45__6_, r_45__5_, r_45__4_, r_45__3_, r_45__2_, r_45__1_, r_45__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N89)? data_i : 1'b0;
  assign N88 = sel_i[88];
  assign N89 = N736;
  assign { r_n_45__31_, r_n_45__30_, r_n_45__29_, r_n_45__28_, r_n_45__27_, r_n_45__26_, r_n_45__25_, r_n_45__24_, r_n_45__23_, r_n_45__22_, r_n_45__21_, r_n_45__20_, r_n_45__19_, r_n_45__18_, r_n_45__17_, r_n_45__16_, r_n_45__15_, r_n_45__14_, r_n_45__13_, r_n_45__12_, r_n_45__11_, r_n_45__10_, r_n_45__9_, r_n_45__8_, r_n_45__7_, r_n_45__6_, r_n_45__5_, r_n_45__4_, r_n_45__3_, r_n_45__2_, r_n_45__1_, r_n_45__0_ } = (N90)? { r_46__31_, r_46__30_, r_46__29_, r_46__28_, r_46__27_, r_46__26_, r_46__25_, r_46__24_, r_46__23_, r_46__22_, r_46__21_, r_46__20_, r_46__19_, r_46__18_, r_46__17_, r_46__16_, r_46__15_, r_46__14_, r_46__13_, r_46__12_, r_46__11_, r_46__10_, r_46__9_, r_46__8_, r_46__7_, r_46__6_, r_46__5_, r_46__4_, r_46__3_, r_46__2_, r_46__1_, r_46__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N91)? data_i : 1'b0;
  assign N90 = sel_i[90];
  assign N91 = N741;
  assign { r_n_46__31_, r_n_46__30_, r_n_46__29_, r_n_46__28_, r_n_46__27_, r_n_46__26_, r_n_46__25_, r_n_46__24_, r_n_46__23_, r_n_46__22_, r_n_46__21_, r_n_46__20_, r_n_46__19_, r_n_46__18_, r_n_46__17_, r_n_46__16_, r_n_46__15_, r_n_46__14_, r_n_46__13_, r_n_46__12_, r_n_46__11_, r_n_46__10_, r_n_46__9_, r_n_46__8_, r_n_46__7_, r_n_46__6_, r_n_46__5_, r_n_46__4_, r_n_46__3_, r_n_46__2_, r_n_46__1_, r_n_46__0_ } = (N92)? { r_47__31_, r_47__30_, r_47__29_, r_47__28_, r_47__27_, r_47__26_, r_47__25_, r_47__24_, r_47__23_, r_47__22_, r_47__21_, r_47__20_, r_47__19_, r_47__18_, r_47__17_, r_47__16_, r_47__15_, r_47__14_, r_47__13_, r_47__12_, r_47__11_, r_47__10_, r_47__9_, r_47__8_, r_47__7_, r_47__6_, r_47__5_, r_47__4_, r_47__3_, r_47__2_, r_47__1_, r_47__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N93)? data_i : 1'b0;
  assign N92 = sel_i[92];
  assign N93 = N746;
  assign { r_n_47__31_, r_n_47__30_, r_n_47__29_, r_n_47__28_, r_n_47__27_, r_n_47__26_, r_n_47__25_, r_n_47__24_, r_n_47__23_, r_n_47__22_, r_n_47__21_, r_n_47__20_, r_n_47__19_, r_n_47__18_, r_n_47__17_, r_n_47__16_, r_n_47__15_, r_n_47__14_, r_n_47__13_, r_n_47__12_, r_n_47__11_, r_n_47__10_, r_n_47__9_, r_n_47__8_, r_n_47__7_, r_n_47__6_, r_n_47__5_, r_n_47__4_, r_n_47__3_, r_n_47__2_, r_n_47__1_, r_n_47__0_ } = (N94)? { r_48__31_, r_48__30_, r_48__29_, r_48__28_, r_48__27_, r_48__26_, r_48__25_, r_48__24_, r_48__23_, r_48__22_, r_48__21_, r_48__20_, r_48__19_, r_48__18_, r_48__17_, r_48__16_, r_48__15_, r_48__14_, r_48__13_, r_48__12_, r_48__11_, r_48__10_, r_48__9_, r_48__8_, r_48__7_, r_48__6_, r_48__5_, r_48__4_, r_48__3_, r_48__2_, r_48__1_, r_48__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N95)? data_i : 1'b0;
  assign N94 = sel_i[94];
  assign N95 = N751;
  assign { r_n_48__31_, r_n_48__30_, r_n_48__29_, r_n_48__28_, r_n_48__27_, r_n_48__26_, r_n_48__25_, r_n_48__24_, r_n_48__23_, r_n_48__22_, r_n_48__21_, r_n_48__20_, r_n_48__19_, r_n_48__18_, r_n_48__17_, r_n_48__16_, r_n_48__15_, r_n_48__14_, r_n_48__13_, r_n_48__12_, r_n_48__11_, r_n_48__10_, r_n_48__9_, r_n_48__8_, r_n_48__7_, r_n_48__6_, r_n_48__5_, r_n_48__4_, r_n_48__3_, r_n_48__2_, r_n_48__1_, r_n_48__0_ } = (N96)? { r_49__31_, r_49__30_, r_49__29_, r_49__28_, r_49__27_, r_49__26_, r_49__25_, r_49__24_, r_49__23_, r_49__22_, r_49__21_, r_49__20_, r_49__19_, r_49__18_, r_49__17_, r_49__16_, r_49__15_, r_49__14_, r_49__13_, r_49__12_, r_49__11_, r_49__10_, r_49__9_, r_49__8_, r_49__7_, r_49__6_, r_49__5_, r_49__4_, r_49__3_, r_49__2_, r_49__1_, r_49__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N97)? data_i : 1'b0;
  assign N96 = sel_i[96];
  assign N97 = N756;
  assign { r_n_49__31_, r_n_49__30_, r_n_49__29_, r_n_49__28_, r_n_49__27_, r_n_49__26_, r_n_49__25_, r_n_49__24_, r_n_49__23_, r_n_49__22_, r_n_49__21_, r_n_49__20_, r_n_49__19_, r_n_49__18_, r_n_49__17_, r_n_49__16_, r_n_49__15_, r_n_49__14_, r_n_49__13_, r_n_49__12_, r_n_49__11_, r_n_49__10_, r_n_49__9_, r_n_49__8_, r_n_49__7_, r_n_49__6_, r_n_49__5_, r_n_49__4_, r_n_49__3_, r_n_49__2_, r_n_49__1_, r_n_49__0_ } = (N98)? { r_50__31_, r_50__30_, r_50__29_, r_50__28_, r_50__27_, r_50__26_, r_50__25_, r_50__24_, r_50__23_, r_50__22_, r_50__21_, r_50__20_, r_50__19_, r_50__18_, r_50__17_, r_50__16_, r_50__15_, r_50__14_, r_50__13_, r_50__12_, r_50__11_, r_50__10_, r_50__9_, r_50__8_, r_50__7_, r_50__6_, r_50__5_, r_50__4_, r_50__3_, r_50__2_, r_50__1_, r_50__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N99)? data_i : 1'b0;
  assign N98 = sel_i[98];
  assign N99 = N761;
  assign { r_n_50__31_, r_n_50__30_, r_n_50__29_, r_n_50__28_, r_n_50__27_, r_n_50__26_, r_n_50__25_, r_n_50__24_, r_n_50__23_, r_n_50__22_, r_n_50__21_, r_n_50__20_, r_n_50__19_, r_n_50__18_, r_n_50__17_, r_n_50__16_, r_n_50__15_, r_n_50__14_, r_n_50__13_, r_n_50__12_, r_n_50__11_, r_n_50__10_, r_n_50__9_, r_n_50__8_, r_n_50__7_, r_n_50__6_, r_n_50__5_, r_n_50__4_, r_n_50__3_, r_n_50__2_, r_n_50__1_, r_n_50__0_ } = (N100)? { r_51__31_, r_51__30_, r_51__29_, r_51__28_, r_51__27_, r_51__26_, r_51__25_, r_51__24_, r_51__23_, r_51__22_, r_51__21_, r_51__20_, r_51__19_, r_51__18_, r_51__17_, r_51__16_, r_51__15_, r_51__14_, r_51__13_, r_51__12_, r_51__11_, r_51__10_, r_51__9_, r_51__8_, r_51__7_, r_51__6_, r_51__5_, r_51__4_, r_51__3_, r_51__2_, r_51__1_, r_51__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N101)? data_i : 1'b0;
  assign N100 = sel_i[100];
  assign N101 = N766;
  assign { r_n_51__31_, r_n_51__30_, r_n_51__29_, r_n_51__28_, r_n_51__27_, r_n_51__26_, r_n_51__25_, r_n_51__24_, r_n_51__23_, r_n_51__22_, r_n_51__21_, r_n_51__20_, r_n_51__19_, r_n_51__18_, r_n_51__17_, r_n_51__16_, r_n_51__15_, r_n_51__14_, r_n_51__13_, r_n_51__12_, r_n_51__11_, r_n_51__10_, r_n_51__9_, r_n_51__8_, r_n_51__7_, r_n_51__6_, r_n_51__5_, r_n_51__4_, r_n_51__3_, r_n_51__2_, r_n_51__1_, r_n_51__0_ } = (N102)? { r_52__31_, r_52__30_, r_52__29_, r_52__28_, r_52__27_, r_52__26_, r_52__25_, r_52__24_, r_52__23_, r_52__22_, r_52__21_, r_52__20_, r_52__19_, r_52__18_, r_52__17_, r_52__16_, r_52__15_, r_52__14_, r_52__13_, r_52__12_, r_52__11_, r_52__10_, r_52__9_, r_52__8_, r_52__7_, r_52__6_, r_52__5_, r_52__4_, r_52__3_, r_52__2_, r_52__1_, r_52__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N103)? data_i : 1'b0;
  assign N102 = sel_i[102];
  assign N103 = N771;
  assign { r_n_52__31_, r_n_52__30_, r_n_52__29_, r_n_52__28_, r_n_52__27_, r_n_52__26_, r_n_52__25_, r_n_52__24_, r_n_52__23_, r_n_52__22_, r_n_52__21_, r_n_52__20_, r_n_52__19_, r_n_52__18_, r_n_52__17_, r_n_52__16_, r_n_52__15_, r_n_52__14_, r_n_52__13_, r_n_52__12_, r_n_52__11_, r_n_52__10_, r_n_52__9_, r_n_52__8_, r_n_52__7_, r_n_52__6_, r_n_52__5_, r_n_52__4_, r_n_52__3_, r_n_52__2_, r_n_52__1_, r_n_52__0_ } = (N104)? { r_53__31_, r_53__30_, r_53__29_, r_53__28_, r_53__27_, r_53__26_, r_53__25_, r_53__24_, r_53__23_, r_53__22_, r_53__21_, r_53__20_, r_53__19_, r_53__18_, r_53__17_, r_53__16_, r_53__15_, r_53__14_, r_53__13_, r_53__12_, r_53__11_, r_53__10_, r_53__9_, r_53__8_, r_53__7_, r_53__6_, r_53__5_, r_53__4_, r_53__3_, r_53__2_, r_53__1_, r_53__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N105)? data_i : 1'b0;
  assign N104 = sel_i[104];
  assign N105 = N776;
  assign { r_n_53__31_, r_n_53__30_, r_n_53__29_, r_n_53__28_, r_n_53__27_, r_n_53__26_, r_n_53__25_, r_n_53__24_, r_n_53__23_, r_n_53__22_, r_n_53__21_, r_n_53__20_, r_n_53__19_, r_n_53__18_, r_n_53__17_, r_n_53__16_, r_n_53__15_, r_n_53__14_, r_n_53__13_, r_n_53__12_, r_n_53__11_, r_n_53__10_, r_n_53__9_, r_n_53__8_, r_n_53__7_, r_n_53__6_, r_n_53__5_, r_n_53__4_, r_n_53__3_, r_n_53__2_, r_n_53__1_, r_n_53__0_ } = (N106)? { r_54__31_, r_54__30_, r_54__29_, r_54__28_, r_54__27_, r_54__26_, r_54__25_, r_54__24_, r_54__23_, r_54__22_, r_54__21_, r_54__20_, r_54__19_, r_54__18_, r_54__17_, r_54__16_, r_54__15_, r_54__14_, r_54__13_, r_54__12_, r_54__11_, r_54__10_, r_54__9_, r_54__8_, r_54__7_, r_54__6_, r_54__5_, r_54__4_, r_54__3_, r_54__2_, r_54__1_, r_54__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N107)? data_i : 1'b0;
  assign N106 = sel_i[106];
  assign N107 = N781;
  assign { r_n_54__31_, r_n_54__30_, r_n_54__29_, r_n_54__28_, r_n_54__27_, r_n_54__26_, r_n_54__25_, r_n_54__24_, r_n_54__23_, r_n_54__22_, r_n_54__21_, r_n_54__20_, r_n_54__19_, r_n_54__18_, r_n_54__17_, r_n_54__16_, r_n_54__15_, r_n_54__14_, r_n_54__13_, r_n_54__12_, r_n_54__11_, r_n_54__10_, r_n_54__9_, r_n_54__8_, r_n_54__7_, r_n_54__6_, r_n_54__5_, r_n_54__4_, r_n_54__3_, r_n_54__2_, r_n_54__1_, r_n_54__0_ } = (N108)? { r_55__31_, r_55__30_, r_55__29_, r_55__28_, r_55__27_, r_55__26_, r_55__25_, r_55__24_, r_55__23_, r_55__22_, r_55__21_, r_55__20_, r_55__19_, r_55__18_, r_55__17_, r_55__16_, r_55__15_, r_55__14_, r_55__13_, r_55__12_, r_55__11_, r_55__10_, r_55__9_, r_55__8_, r_55__7_, r_55__6_, r_55__5_, r_55__4_, r_55__3_, r_55__2_, r_55__1_, r_55__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N109)? data_i : 1'b0;
  assign N108 = sel_i[108];
  assign N109 = N786;
  assign { r_n_55__31_, r_n_55__30_, r_n_55__29_, r_n_55__28_, r_n_55__27_, r_n_55__26_, r_n_55__25_, r_n_55__24_, r_n_55__23_, r_n_55__22_, r_n_55__21_, r_n_55__20_, r_n_55__19_, r_n_55__18_, r_n_55__17_, r_n_55__16_, r_n_55__15_, r_n_55__14_, r_n_55__13_, r_n_55__12_, r_n_55__11_, r_n_55__10_, r_n_55__9_, r_n_55__8_, r_n_55__7_, r_n_55__6_, r_n_55__5_, r_n_55__4_, r_n_55__3_, r_n_55__2_, r_n_55__1_, r_n_55__0_ } = (N110)? { r_56__31_, r_56__30_, r_56__29_, r_56__28_, r_56__27_, r_56__26_, r_56__25_, r_56__24_, r_56__23_, r_56__22_, r_56__21_, r_56__20_, r_56__19_, r_56__18_, r_56__17_, r_56__16_, r_56__15_, r_56__14_, r_56__13_, r_56__12_, r_56__11_, r_56__10_, r_56__9_, r_56__8_, r_56__7_, r_56__6_, r_56__5_, r_56__4_, r_56__3_, r_56__2_, r_56__1_, r_56__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N111)? data_i : 1'b0;
  assign N110 = sel_i[110];
  assign N111 = N791;
  assign { r_n_56__31_, r_n_56__30_, r_n_56__29_, r_n_56__28_, r_n_56__27_, r_n_56__26_, r_n_56__25_, r_n_56__24_, r_n_56__23_, r_n_56__22_, r_n_56__21_, r_n_56__20_, r_n_56__19_, r_n_56__18_, r_n_56__17_, r_n_56__16_, r_n_56__15_, r_n_56__14_, r_n_56__13_, r_n_56__12_, r_n_56__11_, r_n_56__10_, r_n_56__9_, r_n_56__8_, r_n_56__7_, r_n_56__6_, r_n_56__5_, r_n_56__4_, r_n_56__3_, r_n_56__2_, r_n_56__1_, r_n_56__0_ } = (N112)? { r_57__31_, r_57__30_, r_57__29_, r_57__28_, r_57__27_, r_57__26_, r_57__25_, r_57__24_, r_57__23_, r_57__22_, r_57__21_, r_57__20_, r_57__19_, r_57__18_, r_57__17_, r_57__16_, r_57__15_, r_57__14_, r_57__13_, r_57__12_, r_57__11_, r_57__10_, r_57__9_, r_57__8_, r_57__7_, r_57__6_, r_57__5_, r_57__4_, r_57__3_, r_57__2_, r_57__1_, r_57__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N113)? data_i : 1'b0;
  assign N112 = sel_i[112];
  assign N113 = N796;
  assign { r_n_57__31_, r_n_57__30_, r_n_57__29_, r_n_57__28_, r_n_57__27_, r_n_57__26_, r_n_57__25_, r_n_57__24_, r_n_57__23_, r_n_57__22_, r_n_57__21_, r_n_57__20_, r_n_57__19_, r_n_57__18_, r_n_57__17_, r_n_57__16_, r_n_57__15_, r_n_57__14_, r_n_57__13_, r_n_57__12_, r_n_57__11_, r_n_57__10_, r_n_57__9_, r_n_57__8_, r_n_57__7_, r_n_57__6_, r_n_57__5_, r_n_57__4_, r_n_57__3_, r_n_57__2_, r_n_57__1_, r_n_57__0_ } = (N114)? { r_58__31_, r_58__30_, r_58__29_, r_58__28_, r_58__27_, r_58__26_, r_58__25_, r_58__24_, r_58__23_, r_58__22_, r_58__21_, r_58__20_, r_58__19_, r_58__18_, r_58__17_, r_58__16_, r_58__15_, r_58__14_, r_58__13_, r_58__12_, r_58__11_, r_58__10_, r_58__9_, r_58__8_, r_58__7_, r_58__6_, r_58__5_, r_58__4_, r_58__3_, r_58__2_, r_58__1_, r_58__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N115)? data_i : 1'b0;
  assign N114 = sel_i[114];
  assign N115 = N801;
  assign { r_n_58__31_, r_n_58__30_, r_n_58__29_, r_n_58__28_, r_n_58__27_, r_n_58__26_, r_n_58__25_, r_n_58__24_, r_n_58__23_, r_n_58__22_, r_n_58__21_, r_n_58__20_, r_n_58__19_, r_n_58__18_, r_n_58__17_, r_n_58__16_, r_n_58__15_, r_n_58__14_, r_n_58__13_, r_n_58__12_, r_n_58__11_, r_n_58__10_, r_n_58__9_, r_n_58__8_, r_n_58__7_, r_n_58__6_, r_n_58__5_, r_n_58__4_, r_n_58__3_, r_n_58__2_, r_n_58__1_, r_n_58__0_ } = (N116)? { r_59__31_, r_59__30_, r_59__29_, r_59__28_, r_59__27_, r_59__26_, r_59__25_, r_59__24_, r_59__23_, r_59__22_, r_59__21_, r_59__20_, r_59__19_, r_59__18_, r_59__17_, r_59__16_, r_59__15_, r_59__14_, r_59__13_, r_59__12_, r_59__11_, r_59__10_, r_59__9_, r_59__8_, r_59__7_, r_59__6_, r_59__5_, r_59__4_, r_59__3_, r_59__2_, r_59__1_, r_59__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N117)? data_i : 1'b0;
  assign N116 = sel_i[116];
  assign N117 = N806;
  assign { r_n_59__31_, r_n_59__30_, r_n_59__29_, r_n_59__28_, r_n_59__27_, r_n_59__26_, r_n_59__25_, r_n_59__24_, r_n_59__23_, r_n_59__22_, r_n_59__21_, r_n_59__20_, r_n_59__19_, r_n_59__18_, r_n_59__17_, r_n_59__16_, r_n_59__15_, r_n_59__14_, r_n_59__13_, r_n_59__12_, r_n_59__11_, r_n_59__10_, r_n_59__9_, r_n_59__8_, r_n_59__7_, r_n_59__6_, r_n_59__5_, r_n_59__4_, r_n_59__3_, r_n_59__2_, r_n_59__1_, r_n_59__0_ } = (N118)? { r_60__31_, r_60__30_, r_60__29_, r_60__28_, r_60__27_, r_60__26_, r_60__25_, r_60__24_, r_60__23_, r_60__22_, r_60__21_, r_60__20_, r_60__19_, r_60__18_, r_60__17_, r_60__16_, r_60__15_, r_60__14_, r_60__13_, r_60__12_, r_60__11_, r_60__10_, r_60__9_, r_60__8_, r_60__7_, r_60__6_, r_60__5_, r_60__4_, r_60__3_, r_60__2_, r_60__1_, r_60__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N119)? data_i : 1'b0;
  assign N118 = sel_i[118];
  assign N119 = N811;
  assign { r_n_60__31_, r_n_60__30_, r_n_60__29_, r_n_60__28_, r_n_60__27_, r_n_60__26_, r_n_60__25_, r_n_60__24_, r_n_60__23_, r_n_60__22_, r_n_60__21_, r_n_60__20_, r_n_60__19_, r_n_60__18_, r_n_60__17_, r_n_60__16_, r_n_60__15_, r_n_60__14_, r_n_60__13_, r_n_60__12_, r_n_60__11_, r_n_60__10_, r_n_60__9_, r_n_60__8_, r_n_60__7_, r_n_60__6_, r_n_60__5_, r_n_60__4_, r_n_60__3_, r_n_60__2_, r_n_60__1_, r_n_60__0_ } = (N120)? { r_61__31_, r_61__30_, r_61__29_, r_61__28_, r_61__27_, r_61__26_, r_61__25_, r_61__24_, r_61__23_, r_61__22_, r_61__21_, r_61__20_, r_61__19_, r_61__18_, r_61__17_, r_61__16_, r_61__15_, r_61__14_, r_61__13_, r_61__12_, r_61__11_, r_61__10_, r_61__9_, r_61__8_, r_61__7_, r_61__6_, r_61__5_, r_61__4_, r_61__3_, r_61__2_, r_61__1_, r_61__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N121)? data_i : 1'b0;
  assign N120 = sel_i[120];
  assign N121 = N816;
  assign { r_n_61__31_, r_n_61__30_, r_n_61__29_, r_n_61__28_, r_n_61__27_, r_n_61__26_, r_n_61__25_, r_n_61__24_, r_n_61__23_, r_n_61__22_, r_n_61__21_, r_n_61__20_, r_n_61__19_, r_n_61__18_, r_n_61__17_, r_n_61__16_, r_n_61__15_, r_n_61__14_, r_n_61__13_, r_n_61__12_, r_n_61__11_, r_n_61__10_, r_n_61__9_, r_n_61__8_, r_n_61__7_, r_n_61__6_, r_n_61__5_, r_n_61__4_, r_n_61__3_, r_n_61__2_, r_n_61__1_, r_n_61__0_ } = (N122)? { r_62__31_, r_62__30_, r_62__29_, r_62__28_, r_62__27_, r_62__26_, r_62__25_, r_62__24_, r_62__23_, r_62__22_, r_62__21_, r_62__20_, r_62__19_, r_62__18_, r_62__17_, r_62__16_, r_62__15_, r_62__14_, r_62__13_, r_62__12_, r_62__11_, r_62__10_, r_62__9_, r_62__8_, r_62__7_, r_62__6_, r_62__5_, r_62__4_, r_62__3_, r_62__2_, r_62__1_, r_62__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N123)? data_i : 1'b0;
  assign N122 = sel_i[122];
  assign N123 = N821;
  assign { r_n_62__31_, r_n_62__30_, r_n_62__29_, r_n_62__28_, r_n_62__27_, r_n_62__26_, r_n_62__25_, r_n_62__24_, r_n_62__23_, r_n_62__22_, r_n_62__21_, r_n_62__20_, r_n_62__19_, r_n_62__18_, r_n_62__17_, r_n_62__16_, r_n_62__15_, r_n_62__14_, r_n_62__13_, r_n_62__12_, r_n_62__11_, r_n_62__10_, r_n_62__9_, r_n_62__8_, r_n_62__7_, r_n_62__6_, r_n_62__5_, r_n_62__4_, r_n_62__3_, r_n_62__2_, r_n_62__1_, r_n_62__0_ } = (N124)? { r_63__31_, r_63__30_, r_63__29_, r_63__28_, r_63__27_, r_63__26_, r_63__25_, r_63__24_, r_63__23_, r_63__22_, r_63__21_, r_63__20_, r_63__19_, r_63__18_, r_63__17_, r_63__16_, r_63__15_, r_63__14_, r_63__13_, r_63__12_, r_63__11_, r_63__10_, r_63__9_, r_63__8_, r_63__7_, r_63__6_, r_63__5_, r_63__4_, r_63__3_, r_63__2_, r_63__1_, r_63__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N125)? data_i : 1'b0;
  assign N124 = sel_i[124];
  assign N125 = N826;
  assign { r_n_63__31_, r_n_63__30_, r_n_63__29_, r_n_63__28_, r_n_63__27_, r_n_63__26_, r_n_63__25_, r_n_63__24_, r_n_63__23_, r_n_63__22_, r_n_63__21_, r_n_63__20_, r_n_63__19_, r_n_63__18_, r_n_63__17_, r_n_63__16_, r_n_63__15_, r_n_63__14_, r_n_63__13_, r_n_63__12_, r_n_63__11_, r_n_63__10_, r_n_63__9_, r_n_63__8_, r_n_63__7_, r_n_63__6_, r_n_63__5_, r_n_63__4_, r_n_63__3_, r_n_63__2_, r_n_63__1_, r_n_63__0_ } = (N126)? { r_64__31_, r_64__30_, r_64__29_, r_64__28_, r_64__27_, r_64__26_, r_64__25_, r_64__24_, r_64__23_, r_64__22_, r_64__21_, r_64__20_, r_64__19_, r_64__18_, r_64__17_, r_64__16_, r_64__15_, r_64__14_, r_64__13_, r_64__12_, r_64__11_, r_64__10_, r_64__9_, r_64__8_, r_64__7_, r_64__6_, r_64__5_, r_64__4_, r_64__3_, r_64__2_, r_64__1_, r_64__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N127)? data_i : 1'b0;
  assign N126 = sel_i[126];
  assign N127 = N831;
  assign { r_n_64__31_, r_n_64__30_, r_n_64__29_, r_n_64__28_, r_n_64__27_, r_n_64__26_, r_n_64__25_, r_n_64__24_, r_n_64__23_, r_n_64__22_, r_n_64__21_, r_n_64__20_, r_n_64__19_, r_n_64__18_, r_n_64__17_, r_n_64__16_, r_n_64__15_, r_n_64__14_, r_n_64__13_, r_n_64__12_, r_n_64__11_, r_n_64__10_, r_n_64__9_, r_n_64__8_, r_n_64__7_, r_n_64__6_, r_n_64__5_, r_n_64__4_, r_n_64__3_, r_n_64__2_, r_n_64__1_, r_n_64__0_ } = (N128)? { r_65__31_, r_65__30_, r_65__29_, r_65__28_, r_65__27_, r_65__26_, r_65__25_, r_65__24_, r_65__23_, r_65__22_, r_65__21_, r_65__20_, r_65__19_, r_65__18_, r_65__17_, r_65__16_, r_65__15_, r_65__14_, r_65__13_, r_65__12_, r_65__11_, r_65__10_, r_65__9_, r_65__8_, r_65__7_, r_65__6_, r_65__5_, r_65__4_, r_65__3_, r_65__2_, r_65__1_, r_65__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N129)? data_i : 1'b0;
  assign N128 = sel_i[128];
  assign N129 = N836;
  assign { r_n_65__31_, r_n_65__30_, r_n_65__29_, r_n_65__28_, r_n_65__27_, r_n_65__26_, r_n_65__25_, r_n_65__24_, r_n_65__23_, r_n_65__22_, r_n_65__21_, r_n_65__20_, r_n_65__19_, r_n_65__18_, r_n_65__17_, r_n_65__16_, r_n_65__15_, r_n_65__14_, r_n_65__13_, r_n_65__12_, r_n_65__11_, r_n_65__10_, r_n_65__9_, r_n_65__8_, r_n_65__7_, r_n_65__6_, r_n_65__5_, r_n_65__4_, r_n_65__3_, r_n_65__2_, r_n_65__1_, r_n_65__0_ } = (N130)? { r_66__31_, r_66__30_, r_66__29_, r_66__28_, r_66__27_, r_66__26_, r_66__25_, r_66__24_, r_66__23_, r_66__22_, r_66__21_, r_66__20_, r_66__19_, r_66__18_, r_66__17_, r_66__16_, r_66__15_, r_66__14_, r_66__13_, r_66__12_, r_66__11_, r_66__10_, r_66__9_, r_66__8_, r_66__7_, r_66__6_, r_66__5_, r_66__4_, r_66__3_, r_66__2_, r_66__1_, r_66__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N131)? data_i : 1'b0;
  assign N130 = sel_i[130];
  assign N131 = N841;
  assign { r_n_66__31_, r_n_66__30_, r_n_66__29_, r_n_66__28_, r_n_66__27_, r_n_66__26_, r_n_66__25_, r_n_66__24_, r_n_66__23_, r_n_66__22_, r_n_66__21_, r_n_66__20_, r_n_66__19_, r_n_66__18_, r_n_66__17_, r_n_66__16_, r_n_66__15_, r_n_66__14_, r_n_66__13_, r_n_66__12_, r_n_66__11_, r_n_66__10_, r_n_66__9_, r_n_66__8_, r_n_66__7_, r_n_66__6_, r_n_66__5_, r_n_66__4_, r_n_66__3_, r_n_66__2_, r_n_66__1_, r_n_66__0_ } = (N132)? { r_67__31_, r_67__30_, r_67__29_, r_67__28_, r_67__27_, r_67__26_, r_67__25_, r_67__24_, r_67__23_, r_67__22_, r_67__21_, r_67__20_, r_67__19_, r_67__18_, r_67__17_, r_67__16_, r_67__15_, r_67__14_, r_67__13_, r_67__12_, r_67__11_, r_67__10_, r_67__9_, r_67__8_, r_67__7_, r_67__6_, r_67__5_, r_67__4_, r_67__3_, r_67__2_, r_67__1_, r_67__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N133)? data_i : 1'b0;
  assign N132 = sel_i[132];
  assign N133 = N846;
  assign { r_n_67__31_, r_n_67__30_, r_n_67__29_, r_n_67__28_, r_n_67__27_, r_n_67__26_, r_n_67__25_, r_n_67__24_, r_n_67__23_, r_n_67__22_, r_n_67__21_, r_n_67__20_, r_n_67__19_, r_n_67__18_, r_n_67__17_, r_n_67__16_, r_n_67__15_, r_n_67__14_, r_n_67__13_, r_n_67__12_, r_n_67__11_, r_n_67__10_, r_n_67__9_, r_n_67__8_, r_n_67__7_, r_n_67__6_, r_n_67__5_, r_n_67__4_, r_n_67__3_, r_n_67__2_, r_n_67__1_, r_n_67__0_ } = (N134)? { r_68__31_, r_68__30_, r_68__29_, r_68__28_, r_68__27_, r_68__26_, r_68__25_, r_68__24_, r_68__23_, r_68__22_, r_68__21_, r_68__20_, r_68__19_, r_68__18_, r_68__17_, r_68__16_, r_68__15_, r_68__14_, r_68__13_, r_68__12_, r_68__11_, r_68__10_, r_68__9_, r_68__8_, r_68__7_, r_68__6_, r_68__5_, r_68__4_, r_68__3_, r_68__2_, r_68__1_, r_68__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N135)? data_i : 1'b0;
  assign N134 = sel_i[134];
  assign N135 = N851;
  assign { r_n_68__31_, r_n_68__30_, r_n_68__29_, r_n_68__28_, r_n_68__27_, r_n_68__26_, r_n_68__25_, r_n_68__24_, r_n_68__23_, r_n_68__22_, r_n_68__21_, r_n_68__20_, r_n_68__19_, r_n_68__18_, r_n_68__17_, r_n_68__16_, r_n_68__15_, r_n_68__14_, r_n_68__13_, r_n_68__12_, r_n_68__11_, r_n_68__10_, r_n_68__9_, r_n_68__8_, r_n_68__7_, r_n_68__6_, r_n_68__5_, r_n_68__4_, r_n_68__3_, r_n_68__2_, r_n_68__1_, r_n_68__0_ } = (N136)? { r_69__31_, r_69__30_, r_69__29_, r_69__28_, r_69__27_, r_69__26_, r_69__25_, r_69__24_, r_69__23_, r_69__22_, r_69__21_, r_69__20_, r_69__19_, r_69__18_, r_69__17_, r_69__16_, r_69__15_, r_69__14_, r_69__13_, r_69__12_, r_69__11_, r_69__10_, r_69__9_, r_69__8_, r_69__7_, r_69__6_, r_69__5_, r_69__4_, r_69__3_, r_69__2_, r_69__1_, r_69__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N137)? data_i : 1'b0;
  assign N136 = sel_i[136];
  assign N137 = N856;
  assign { r_n_69__31_, r_n_69__30_, r_n_69__29_, r_n_69__28_, r_n_69__27_, r_n_69__26_, r_n_69__25_, r_n_69__24_, r_n_69__23_, r_n_69__22_, r_n_69__21_, r_n_69__20_, r_n_69__19_, r_n_69__18_, r_n_69__17_, r_n_69__16_, r_n_69__15_, r_n_69__14_, r_n_69__13_, r_n_69__12_, r_n_69__11_, r_n_69__10_, r_n_69__9_, r_n_69__8_, r_n_69__7_, r_n_69__6_, r_n_69__5_, r_n_69__4_, r_n_69__3_, r_n_69__2_, r_n_69__1_, r_n_69__0_ } = (N138)? { r_70__31_, r_70__30_, r_70__29_, r_70__28_, r_70__27_, r_70__26_, r_70__25_, r_70__24_, r_70__23_, r_70__22_, r_70__21_, r_70__20_, r_70__19_, r_70__18_, r_70__17_, r_70__16_, r_70__15_, r_70__14_, r_70__13_, r_70__12_, r_70__11_, r_70__10_, r_70__9_, r_70__8_, r_70__7_, r_70__6_, r_70__5_, r_70__4_, r_70__3_, r_70__2_, r_70__1_, r_70__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N139)? data_i : 1'b0;
  assign N138 = sel_i[138];
  assign N139 = N861;
  assign { r_n_70__31_, r_n_70__30_, r_n_70__29_, r_n_70__28_, r_n_70__27_, r_n_70__26_, r_n_70__25_, r_n_70__24_, r_n_70__23_, r_n_70__22_, r_n_70__21_, r_n_70__20_, r_n_70__19_, r_n_70__18_, r_n_70__17_, r_n_70__16_, r_n_70__15_, r_n_70__14_, r_n_70__13_, r_n_70__12_, r_n_70__11_, r_n_70__10_, r_n_70__9_, r_n_70__8_, r_n_70__7_, r_n_70__6_, r_n_70__5_, r_n_70__4_, r_n_70__3_, r_n_70__2_, r_n_70__1_, r_n_70__0_ } = (N140)? { r_71__31_, r_71__30_, r_71__29_, r_71__28_, r_71__27_, r_71__26_, r_71__25_, r_71__24_, r_71__23_, r_71__22_, r_71__21_, r_71__20_, r_71__19_, r_71__18_, r_71__17_, r_71__16_, r_71__15_, r_71__14_, r_71__13_, r_71__12_, r_71__11_, r_71__10_, r_71__9_, r_71__8_, r_71__7_, r_71__6_, r_71__5_, r_71__4_, r_71__3_, r_71__2_, r_71__1_, r_71__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N141)? data_i : 1'b0;
  assign N140 = sel_i[140];
  assign N141 = N866;
  assign { r_n_71__31_, r_n_71__30_, r_n_71__29_, r_n_71__28_, r_n_71__27_, r_n_71__26_, r_n_71__25_, r_n_71__24_, r_n_71__23_, r_n_71__22_, r_n_71__21_, r_n_71__20_, r_n_71__19_, r_n_71__18_, r_n_71__17_, r_n_71__16_, r_n_71__15_, r_n_71__14_, r_n_71__13_, r_n_71__12_, r_n_71__11_, r_n_71__10_, r_n_71__9_, r_n_71__8_, r_n_71__7_, r_n_71__6_, r_n_71__5_, r_n_71__4_, r_n_71__3_, r_n_71__2_, r_n_71__1_, r_n_71__0_ } = (N142)? { r_72__31_, r_72__30_, r_72__29_, r_72__28_, r_72__27_, r_72__26_, r_72__25_, r_72__24_, r_72__23_, r_72__22_, r_72__21_, r_72__20_, r_72__19_, r_72__18_, r_72__17_, r_72__16_, r_72__15_, r_72__14_, r_72__13_, r_72__12_, r_72__11_, r_72__10_, r_72__9_, r_72__8_, r_72__7_, r_72__6_, r_72__5_, r_72__4_, r_72__3_, r_72__2_, r_72__1_, r_72__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N143)? data_i : 1'b0;
  assign N142 = sel_i[142];
  assign N143 = N871;
  assign { r_n_72__31_, r_n_72__30_, r_n_72__29_, r_n_72__28_, r_n_72__27_, r_n_72__26_, r_n_72__25_, r_n_72__24_, r_n_72__23_, r_n_72__22_, r_n_72__21_, r_n_72__20_, r_n_72__19_, r_n_72__18_, r_n_72__17_, r_n_72__16_, r_n_72__15_, r_n_72__14_, r_n_72__13_, r_n_72__12_, r_n_72__11_, r_n_72__10_, r_n_72__9_, r_n_72__8_, r_n_72__7_, r_n_72__6_, r_n_72__5_, r_n_72__4_, r_n_72__3_, r_n_72__2_, r_n_72__1_, r_n_72__0_ } = (N144)? { r_73__31_, r_73__30_, r_73__29_, r_73__28_, r_73__27_, r_73__26_, r_73__25_, r_73__24_, r_73__23_, r_73__22_, r_73__21_, r_73__20_, r_73__19_, r_73__18_, r_73__17_, r_73__16_, r_73__15_, r_73__14_, r_73__13_, r_73__12_, r_73__11_, r_73__10_, r_73__9_, r_73__8_, r_73__7_, r_73__6_, r_73__5_, r_73__4_, r_73__3_, r_73__2_, r_73__1_, r_73__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N145)? data_i : 1'b0;
  assign N144 = sel_i[144];
  assign N145 = N876;
  assign { r_n_73__31_, r_n_73__30_, r_n_73__29_, r_n_73__28_, r_n_73__27_, r_n_73__26_, r_n_73__25_, r_n_73__24_, r_n_73__23_, r_n_73__22_, r_n_73__21_, r_n_73__20_, r_n_73__19_, r_n_73__18_, r_n_73__17_, r_n_73__16_, r_n_73__15_, r_n_73__14_, r_n_73__13_, r_n_73__12_, r_n_73__11_, r_n_73__10_, r_n_73__9_, r_n_73__8_, r_n_73__7_, r_n_73__6_, r_n_73__5_, r_n_73__4_, r_n_73__3_, r_n_73__2_, r_n_73__1_, r_n_73__0_ } = (N146)? { r_74__31_, r_74__30_, r_74__29_, r_74__28_, r_74__27_, r_74__26_, r_74__25_, r_74__24_, r_74__23_, r_74__22_, r_74__21_, r_74__20_, r_74__19_, r_74__18_, r_74__17_, r_74__16_, r_74__15_, r_74__14_, r_74__13_, r_74__12_, r_74__11_, r_74__10_, r_74__9_, r_74__8_, r_74__7_, r_74__6_, r_74__5_, r_74__4_, r_74__3_, r_74__2_, r_74__1_, r_74__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N147)? data_i : 1'b0;
  assign N146 = sel_i[146];
  assign N147 = N881;
  assign { r_n_74__31_, r_n_74__30_, r_n_74__29_, r_n_74__28_, r_n_74__27_, r_n_74__26_, r_n_74__25_, r_n_74__24_, r_n_74__23_, r_n_74__22_, r_n_74__21_, r_n_74__20_, r_n_74__19_, r_n_74__18_, r_n_74__17_, r_n_74__16_, r_n_74__15_, r_n_74__14_, r_n_74__13_, r_n_74__12_, r_n_74__11_, r_n_74__10_, r_n_74__9_, r_n_74__8_, r_n_74__7_, r_n_74__6_, r_n_74__5_, r_n_74__4_, r_n_74__3_, r_n_74__2_, r_n_74__1_, r_n_74__0_ } = (N148)? { r_75__31_, r_75__30_, r_75__29_, r_75__28_, r_75__27_, r_75__26_, r_75__25_, r_75__24_, r_75__23_, r_75__22_, r_75__21_, r_75__20_, r_75__19_, r_75__18_, r_75__17_, r_75__16_, r_75__15_, r_75__14_, r_75__13_, r_75__12_, r_75__11_, r_75__10_, r_75__9_, r_75__8_, r_75__7_, r_75__6_, r_75__5_, r_75__4_, r_75__3_, r_75__2_, r_75__1_, r_75__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N149)? data_i : 1'b0;
  assign N148 = sel_i[148];
  assign N149 = N886;
  assign { r_n_75__31_, r_n_75__30_, r_n_75__29_, r_n_75__28_, r_n_75__27_, r_n_75__26_, r_n_75__25_, r_n_75__24_, r_n_75__23_, r_n_75__22_, r_n_75__21_, r_n_75__20_, r_n_75__19_, r_n_75__18_, r_n_75__17_, r_n_75__16_, r_n_75__15_, r_n_75__14_, r_n_75__13_, r_n_75__12_, r_n_75__11_, r_n_75__10_, r_n_75__9_, r_n_75__8_, r_n_75__7_, r_n_75__6_, r_n_75__5_, r_n_75__4_, r_n_75__3_, r_n_75__2_, r_n_75__1_, r_n_75__0_ } = (N150)? { r_76__31_, r_76__30_, r_76__29_, r_76__28_, r_76__27_, r_76__26_, r_76__25_, r_76__24_, r_76__23_, r_76__22_, r_76__21_, r_76__20_, r_76__19_, r_76__18_, r_76__17_, r_76__16_, r_76__15_, r_76__14_, r_76__13_, r_76__12_, r_76__11_, r_76__10_, r_76__9_, r_76__8_, r_76__7_, r_76__6_, r_76__5_, r_76__4_, r_76__3_, r_76__2_, r_76__1_, r_76__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N151)? data_i : 1'b0;
  assign N150 = sel_i[150];
  assign N151 = N891;
  assign { r_n_76__31_, r_n_76__30_, r_n_76__29_, r_n_76__28_, r_n_76__27_, r_n_76__26_, r_n_76__25_, r_n_76__24_, r_n_76__23_, r_n_76__22_, r_n_76__21_, r_n_76__20_, r_n_76__19_, r_n_76__18_, r_n_76__17_, r_n_76__16_, r_n_76__15_, r_n_76__14_, r_n_76__13_, r_n_76__12_, r_n_76__11_, r_n_76__10_, r_n_76__9_, r_n_76__8_, r_n_76__7_, r_n_76__6_, r_n_76__5_, r_n_76__4_, r_n_76__3_, r_n_76__2_, r_n_76__1_, r_n_76__0_ } = (N152)? { r_77__31_, r_77__30_, r_77__29_, r_77__28_, r_77__27_, r_77__26_, r_77__25_, r_77__24_, r_77__23_, r_77__22_, r_77__21_, r_77__20_, r_77__19_, r_77__18_, r_77__17_, r_77__16_, r_77__15_, r_77__14_, r_77__13_, r_77__12_, r_77__11_, r_77__10_, r_77__9_, r_77__8_, r_77__7_, r_77__6_, r_77__5_, r_77__4_, r_77__3_, r_77__2_, r_77__1_, r_77__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N153)? data_i : 1'b0;
  assign N152 = sel_i[152];
  assign N153 = N896;
  assign { r_n_77__31_, r_n_77__30_, r_n_77__29_, r_n_77__28_, r_n_77__27_, r_n_77__26_, r_n_77__25_, r_n_77__24_, r_n_77__23_, r_n_77__22_, r_n_77__21_, r_n_77__20_, r_n_77__19_, r_n_77__18_, r_n_77__17_, r_n_77__16_, r_n_77__15_, r_n_77__14_, r_n_77__13_, r_n_77__12_, r_n_77__11_, r_n_77__10_, r_n_77__9_, r_n_77__8_, r_n_77__7_, r_n_77__6_, r_n_77__5_, r_n_77__4_, r_n_77__3_, r_n_77__2_, r_n_77__1_, r_n_77__0_ } = (N154)? { r_78__31_, r_78__30_, r_78__29_, r_78__28_, r_78__27_, r_78__26_, r_78__25_, r_78__24_, r_78__23_, r_78__22_, r_78__21_, r_78__20_, r_78__19_, r_78__18_, r_78__17_, r_78__16_, r_78__15_, r_78__14_, r_78__13_, r_78__12_, r_78__11_, r_78__10_, r_78__9_, r_78__8_, r_78__7_, r_78__6_, r_78__5_, r_78__4_, r_78__3_, r_78__2_, r_78__1_, r_78__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N155)? data_i : 1'b0;
  assign N154 = sel_i[154];
  assign N155 = N901;
  assign { r_n_78__31_, r_n_78__30_, r_n_78__29_, r_n_78__28_, r_n_78__27_, r_n_78__26_, r_n_78__25_, r_n_78__24_, r_n_78__23_, r_n_78__22_, r_n_78__21_, r_n_78__20_, r_n_78__19_, r_n_78__18_, r_n_78__17_, r_n_78__16_, r_n_78__15_, r_n_78__14_, r_n_78__13_, r_n_78__12_, r_n_78__11_, r_n_78__10_, r_n_78__9_, r_n_78__8_, r_n_78__7_, r_n_78__6_, r_n_78__5_, r_n_78__4_, r_n_78__3_, r_n_78__2_, r_n_78__1_, r_n_78__0_ } = (N156)? { r_79__31_, r_79__30_, r_79__29_, r_79__28_, r_79__27_, r_79__26_, r_79__25_, r_79__24_, r_79__23_, r_79__22_, r_79__21_, r_79__20_, r_79__19_, r_79__18_, r_79__17_, r_79__16_, r_79__15_, r_79__14_, r_79__13_, r_79__12_, r_79__11_, r_79__10_, r_79__9_, r_79__8_, r_79__7_, r_79__6_, r_79__5_, r_79__4_, r_79__3_, r_79__2_, r_79__1_, r_79__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N157)? data_i : 1'b0;
  assign N156 = sel_i[156];
  assign N157 = N906;
  assign { r_n_79__31_, r_n_79__30_, r_n_79__29_, r_n_79__28_, r_n_79__27_, r_n_79__26_, r_n_79__25_, r_n_79__24_, r_n_79__23_, r_n_79__22_, r_n_79__21_, r_n_79__20_, r_n_79__19_, r_n_79__18_, r_n_79__17_, r_n_79__16_, r_n_79__15_, r_n_79__14_, r_n_79__13_, r_n_79__12_, r_n_79__11_, r_n_79__10_, r_n_79__9_, r_n_79__8_, r_n_79__7_, r_n_79__6_, r_n_79__5_, r_n_79__4_, r_n_79__3_, r_n_79__2_, r_n_79__1_, r_n_79__0_ } = (N158)? { r_80__31_, r_80__30_, r_80__29_, r_80__28_, r_80__27_, r_80__26_, r_80__25_, r_80__24_, r_80__23_, r_80__22_, r_80__21_, r_80__20_, r_80__19_, r_80__18_, r_80__17_, r_80__16_, r_80__15_, r_80__14_, r_80__13_, r_80__12_, r_80__11_, r_80__10_, r_80__9_, r_80__8_, r_80__7_, r_80__6_, r_80__5_, r_80__4_, r_80__3_, r_80__2_, r_80__1_, r_80__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N159)? data_i : 1'b0;
  assign N158 = sel_i[158];
  assign N159 = N911;
  assign { r_n_80__31_, r_n_80__30_, r_n_80__29_, r_n_80__28_, r_n_80__27_, r_n_80__26_, r_n_80__25_, r_n_80__24_, r_n_80__23_, r_n_80__22_, r_n_80__21_, r_n_80__20_, r_n_80__19_, r_n_80__18_, r_n_80__17_, r_n_80__16_, r_n_80__15_, r_n_80__14_, r_n_80__13_, r_n_80__12_, r_n_80__11_, r_n_80__10_, r_n_80__9_, r_n_80__8_, r_n_80__7_, r_n_80__6_, r_n_80__5_, r_n_80__4_, r_n_80__3_, r_n_80__2_, r_n_80__1_, r_n_80__0_ } = (N160)? { r_81__31_, r_81__30_, r_81__29_, r_81__28_, r_81__27_, r_81__26_, r_81__25_, r_81__24_, r_81__23_, r_81__22_, r_81__21_, r_81__20_, r_81__19_, r_81__18_, r_81__17_, r_81__16_, r_81__15_, r_81__14_, r_81__13_, r_81__12_, r_81__11_, r_81__10_, r_81__9_, r_81__8_, r_81__7_, r_81__6_, r_81__5_, r_81__4_, r_81__3_, r_81__2_, r_81__1_, r_81__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N161)? data_i : 1'b0;
  assign N160 = sel_i[160];
  assign N161 = N916;
  assign { r_n_81__31_, r_n_81__30_, r_n_81__29_, r_n_81__28_, r_n_81__27_, r_n_81__26_, r_n_81__25_, r_n_81__24_, r_n_81__23_, r_n_81__22_, r_n_81__21_, r_n_81__20_, r_n_81__19_, r_n_81__18_, r_n_81__17_, r_n_81__16_, r_n_81__15_, r_n_81__14_, r_n_81__13_, r_n_81__12_, r_n_81__11_, r_n_81__10_, r_n_81__9_, r_n_81__8_, r_n_81__7_, r_n_81__6_, r_n_81__5_, r_n_81__4_, r_n_81__3_, r_n_81__2_, r_n_81__1_, r_n_81__0_ } = (N162)? { r_82__31_, r_82__30_, r_82__29_, r_82__28_, r_82__27_, r_82__26_, r_82__25_, r_82__24_, r_82__23_, r_82__22_, r_82__21_, r_82__20_, r_82__19_, r_82__18_, r_82__17_, r_82__16_, r_82__15_, r_82__14_, r_82__13_, r_82__12_, r_82__11_, r_82__10_, r_82__9_, r_82__8_, r_82__7_, r_82__6_, r_82__5_, r_82__4_, r_82__3_, r_82__2_, r_82__1_, r_82__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N163)? data_i : 1'b0;
  assign N162 = sel_i[162];
  assign N163 = N921;
  assign { r_n_82__31_, r_n_82__30_, r_n_82__29_, r_n_82__28_, r_n_82__27_, r_n_82__26_, r_n_82__25_, r_n_82__24_, r_n_82__23_, r_n_82__22_, r_n_82__21_, r_n_82__20_, r_n_82__19_, r_n_82__18_, r_n_82__17_, r_n_82__16_, r_n_82__15_, r_n_82__14_, r_n_82__13_, r_n_82__12_, r_n_82__11_, r_n_82__10_, r_n_82__9_, r_n_82__8_, r_n_82__7_, r_n_82__6_, r_n_82__5_, r_n_82__4_, r_n_82__3_, r_n_82__2_, r_n_82__1_, r_n_82__0_ } = (N164)? { r_83__31_, r_83__30_, r_83__29_, r_83__28_, r_83__27_, r_83__26_, r_83__25_, r_83__24_, r_83__23_, r_83__22_, r_83__21_, r_83__20_, r_83__19_, r_83__18_, r_83__17_, r_83__16_, r_83__15_, r_83__14_, r_83__13_, r_83__12_, r_83__11_, r_83__10_, r_83__9_, r_83__8_, r_83__7_, r_83__6_, r_83__5_, r_83__4_, r_83__3_, r_83__2_, r_83__1_, r_83__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N165)? data_i : 1'b0;
  assign N164 = sel_i[164];
  assign N165 = N926;
  assign { r_n_83__31_, r_n_83__30_, r_n_83__29_, r_n_83__28_, r_n_83__27_, r_n_83__26_, r_n_83__25_, r_n_83__24_, r_n_83__23_, r_n_83__22_, r_n_83__21_, r_n_83__20_, r_n_83__19_, r_n_83__18_, r_n_83__17_, r_n_83__16_, r_n_83__15_, r_n_83__14_, r_n_83__13_, r_n_83__12_, r_n_83__11_, r_n_83__10_, r_n_83__9_, r_n_83__8_, r_n_83__7_, r_n_83__6_, r_n_83__5_, r_n_83__4_, r_n_83__3_, r_n_83__2_, r_n_83__1_, r_n_83__0_ } = (N166)? { r_84__31_, r_84__30_, r_84__29_, r_84__28_, r_84__27_, r_84__26_, r_84__25_, r_84__24_, r_84__23_, r_84__22_, r_84__21_, r_84__20_, r_84__19_, r_84__18_, r_84__17_, r_84__16_, r_84__15_, r_84__14_, r_84__13_, r_84__12_, r_84__11_, r_84__10_, r_84__9_, r_84__8_, r_84__7_, r_84__6_, r_84__5_, r_84__4_, r_84__3_, r_84__2_, r_84__1_, r_84__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N167)? data_i : 1'b0;
  assign N166 = sel_i[166];
  assign N167 = N931;
  assign { r_n_84__31_, r_n_84__30_, r_n_84__29_, r_n_84__28_, r_n_84__27_, r_n_84__26_, r_n_84__25_, r_n_84__24_, r_n_84__23_, r_n_84__22_, r_n_84__21_, r_n_84__20_, r_n_84__19_, r_n_84__18_, r_n_84__17_, r_n_84__16_, r_n_84__15_, r_n_84__14_, r_n_84__13_, r_n_84__12_, r_n_84__11_, r_n_84__10_, r_n_84__9_, r_n_84__8_, r_n_84__7_, r_n_84__6_, r_n_84__5_, r_n_84__4_, r_n_84__3_, r_n_84__2_, r_n_84__1_, r_n_84__0_ } = (N168)? { r_85__31_, r_85__30_, r_85__29_, r_85__28_, r_85__27_, r_85__26_, r_85__25_, r_85__24_, r_85__23_, r_85__22_, r_85__21_, r_85__20_, r_85__19_, r_85__18_, r_85__17_, r_85__16_, r_85__15_, r_85__14_, r_85__13_, r_85__12_, r_85__11_, r_85__10_, r_85__9_, r_85__8_, r_85__7_, r_85__6_, r_85__5_, r_85__4_, r_85__3_, r_85__2_, r_85__1_, r_85__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N169)? data_i : 1'b0;
  assign N168 = sel_i[168];
  assign N169 = N936;
  assign { r_n_85__31_, r_n_85__30_, r_n_85__29_, r_n_85__28_, r_n_85__27_, r_n_85__26_, r_n_85__25_, r_n_85__24_, r_n_85__23_, r_n_85__22_, r_n_85__21_, r_n_85__20_, r_n_85__19_, r_n_85__18_, r_n_85__17_, r_n_85__16_, r_n_85__15_, r_n_85__14_, r_n_85__13_, r_n_85__12_, r_n_85__11_, r_n_85__10_, r_n_85__9_, r_n_85__8_, r_n_85__7_, r_n_85__6_, r_n_85__5_, r_n_85__4_, r_n_85__3_, r_n_85__2_, r_n_85__1_, r_n_85__0_ } = (N170)? { r_86__31_, r_86__30_, r_86__29_, r_86__28_, r_86__27_, r_86__26_, r_86__25_, r_86__24_, r_86__23_, r_86__22_, r_86__21_, r_86__20_, r_86__19_, r_86__18_, r_86__17_, r_86__16_, r_86__15_, r_86__14_, r_86__13_, r_86__12_, r_86__11_, r_86__10_, r_86__9_, r_86__8_, r_86__7_, r_86__6_, r_86__5_, r_86__4_, r_86__3_, r_86__2_, r_86__1_, r_86__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N171)? data_i : 1'b0;
  assign N170 = sel_i[170];
  assign N171 = N941;
  assign { r_n_86__31_, r_n_86__30_, r_n_86__29_, r_n_86__28_, r_n_86__27_, r_n_86__26_, r_n_86__25_, r_n_86__24_, r_n_86__23_, r_n_86__22_, r_n_86__21_, r_n_86__20_, r_n_86__19_, r_n_86__18_, r_n_86__17_, r_n_86__16_, r_n_86__15_, r_n_86__14_, r_n_86__13_, r_n_86__12_, r_n_86__11_, r_n_86__10_, r_n_86__9_, r_n_86__8_, r_n_86__7_, r_n_86__6_, r_n_86__5_, r_n_86__4_, r_n_86__3_, r_n_86__2_, r_n_86__1_, r_n_86__0_ } = (N172)? { r_87__31_, r_87__30_, r_87__29_, r_87__28_, r_87__27_, r_87__26_, r_87__25_, r_87__24_, r_87__23_, r_87__22_, r_87__21_, r_87__20_, r_87__19_, r_87__18_, r_87__17_, r_87__16_, r_87__15_, r_87__14_, r_87__13_, r_87__12_, r_87__11_, r_87__10_, r_87__9_, r_87__8_, r_87__7_, r_87__6_, r_87__5_, r_87__4_, r_87__3_, r_87__2_, r_87__1_, r_87__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N173)? data_i : 1'b0;
  assign N172 = sel_i[172];
  assign N173 = N946;
  assign { r_n_87__31_, r_n_87__30_, r_n_87__29_, r_n_87__28_, r_n_87__27_, r_n_87__26_, r_n_87__25_, r_n_87__24_, r_n_87__23_, r_n_87__22_, r_n_87__21_, r_n_87__20_, r_n_87__19_, r_n_87__18_, r_n_87__17_, r_n_87__16_, r_n_87__15_, r_n_87__14_, r_n_87__13_, r_n_87__12_, r_n_87__11_, r_n_87__10_, r_n_87__9_, r_n_87__8_, r_n_87__7_, r_n_87__6_, r_n_87__5_, r_n_87__4_, r_n_87__3_, r_n_87__2_, r_n_87__1_, r_n_87__0_ } = (N174)? { r_88__31_, r_88__30_, r_88__29_, r_88__28_, r_88__27_, r_88__26_, r_88__25_, r_88__24_, r_88__23_, r_88__22_, r_88__21_, r_88__20_, r_88__19_, r_88__18_, r_88__17_, r_88__16_, r_88__15_, r_88__14_, r_88__13_, r_88__12_, r_88__11_, r_88__10_, r_88__9_, r_88__8_, r_88__7_, r_88__6_, r_88__5_, r_88__4_, r_88__3_, r_88__2_, r_88__1_, r_88__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N175)? data_i : 1'b0;
  assign N174 = sel_i[174];
  assign N175 = N951;
  assign { r_n_88__31_, r_n_88__30_, r_n_88__29_, r_n_88__28_, r_n_88__27_, r_n_88__26_, r_n_88__25_, r_n_88__24_, r_n_88__23_, r_n_88__22_, r_n_88__21_, r_n_88__20_, r_n_88__19_, r_n_88__18_, r_n_88__17_, r_n_88__16_, r_n_88__15_, r_n_88__14_, r_n_88__13_, r_n_88__12_, r_n_88__11_, r_n_88__10_, r_n_88__9_, r_n_88__8_, r_n_88__7_, r_n_88__6_, r_n_88__5_, r_n_88__4_, r_n_88__3_, r_n_88__2_, r_n_88__1_, r_n_88__0_ } = (N176)? { r_89__31_, r_89__30_, r_89__29_, r_89__28_, r_89__27_, r_89__26_, r_89__25_, r_89__24_, r_89__23_, r_89__22_, r_89__21_, r_89__20_, r_89__19_, r_89__18_, r_89__17_, r_89__16_, r_89__15_, r_89__14_, r_89__13_, r_89__12_, r_89__11_, r_89__10_, r_89__9_, r_89__8_, r_89__7_, r_89__6_, r_89__5_, r_89__4_, r_89__3_, r_89__2_, r_89__1_, r_89__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N177)? data_i : 1'b0;
  assign N176 = sel_i[176];
  assign N177 = N956;
  assign { r_n_89__31_, r_n_89__30_, r_n_89__29_, r_n_89__28_, r_n_89__27_, r_n_89__26_, r_n_89__25_, r_n_89__24_, r_n_89__23_, r_n_89__22_, r_n_89__21_, r_n_89__20_, r_n_89__19_, r_n_89__18_, r_n_89__17_, r_n_89__16_, r_n_89__15_, r_n_89__14_, r_n_89__13_, r_n_89__12_, r_n_89__11_, r_n_89__10_, r_n_89__9_, r_n_89__8_, r_n_89__7_, r_n_89__6_, r_n_89__5_, r_n_89__4_, r_n_89__3_, r_n_89__2_, r_n_89__1_, r_n_89__0_ } = (N178)? { r_90__31_, r_90__30_, r_90__29_, r_90__28_, r_90__27_, r_90__26_, r_90__25_, r_90__24_, r_90__23_, r_90__22_, r_90__21_, r_90__20_, r_90__19_, r_90__18_, r_90__17_, r_90__16_, r_90__15_, r_90__14_, r_90__13_, r_90__12_, r_90__11_, r_90__10_, r_90__9_, r_90__8_, r_90__7_, r_90__6_, r_90__5_, r_90__4_, r_90__3_, r_90__2_, r_90__1_, r_90__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N179)? data_i : 1'b0;
  assign N178 = sel_i[178];
  assign N179 = N961;
  assign { r_n_90__31_, r_n_90__30_, r_n_90__29_, r_n_90__28_, r_n_90__27_, r_n_90__26_, r_n_90__25_, r_n_90__24_, r_n_90__23_, r_n_90__22_, r_n_90__21_, r_n_90__20_, r_n_90__19_, r_n_90__18_, r_n_90__17_, r_n_90__16_, r_n_90__15_, r_n_90__14_, r_n_90__13_, r_n_90__12_, r_n_90__11_, r_n_90__10_, r_n_90__9_, r_n_90__8_, r_n_90__7_, r_n_90__6_, r_n_90__5_, r_n_90__4_, r_n_90__3_, r_n_90__2_, r_n_90__1_, r_n_90__0_ } = (N180)? { r_91__31_, r_91__30_, r_91__29_, r_91__28_, r_91__27_, r_91__26_, r_91__25_, r_91__24_, r_91__23_, r_91__22_, r_91__21_, r_91__20_, r_91__19_, r_91__18_, r_91__17_, r_91__16_, r_91__15_, r_91__14_, r_91__13_, r_91__12_, r_91__11_, r_91__10_, r_91__9_, r_91__8_, r_91__7_, r_91__6_, r_91__5_, r_91__4_, r_91__3_, r_91__2_, r_91__1_, r_91__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N181)? data_i : 1'b0;
  assign N180 = sel_i[180];
  assign N181 = N966;
  assign { r_n_91__31_, r_n_91__30_, r_n_91__29_, r_n_91__28_, r_n_91__27_, r_n_91__26_, r_n_91__25_, r_n_91__24_, r_n_91__23_, r_n_91__22_, r_n_91__21_, r_n_91__20_, r_n_91__19_, r_n_91__18_, r_n_91__17_, r_n_91__16_, r_n_91__15_, r_n_91__14_, r_n_91__13_, r_n_91__12_, r_n_91__11_, r_n_91__10_, r_n_91__9_, r_n_91__8_, r_n_91__7_, r_n_91__6_, r_n_91__5_, r_n_91__4_, r_n_91__3_, r_n_91__2_, r_n_91__1_, r_n_91__0_ } = (N182)? { r_92__31_, r_92__30_, r_92__29_, r_92__28_, r_92__27_, r_92__26_, r_92__25_, r_92__24_, r_92__23_, r_92__22_, r_92__21_, r_92__20_, r_92__19_, r_92__18_, r_92__17_, r_92__16_, r_92__15_, r_92__14_, r_92__13_, r_92__12_, r_92__11_, r_92__10_, r_92__9_, r_92__8_, r_92__7_, r_92__6_, r_92__5_, r_92__4_, r_92__3_, r_92__2_, r_92__1_, r_92__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N183)? data_i : 1'b0;
  assign N182 = sel_i[182];
  assign N183 = N971;
  assign { r_n_92__31_, r_n_92__30_, r_n_92__29_, r_n_92__28_, r_n_92__27_, r_n_92__26_, r_n_92__25_, r_n_92__24_, r_n_92__23_, r_n_92__22_, r_n_92__21_, r_n_92__20_, r_n_92__19_, r_n_92__18_, r_n_92__17_, r_n_92__16_, r_n_92__15_, r_n_92__14_, r_n_92__13_, r_n_92__12_, r_n_92__11_, r_n_92__10_, r_n_92__9_, r_n_92__8_, r_n_92__7_, r_n_92__6_, r_n_92__5_, r_n_92__4_, r_n_92__3_, r_n_92__2_, r_n_92__1_, r_n_92__0_ } = (N184)? { r_93__31_, r_93__30_, r_93__29_, r_93__28_, r_93__27_, r_93__26_, r_93__25_, r_93__24_, r_93__23_, r_93__22_, r_93__21_, r_93__20_, r_93__19_, r_93__18_, r_93__17_, r_93__16_, r_93__15_, r_93__14_, r_93__13_, r_93__12_, r_93__11_, r_93__10_, r_93__9_, r_93__8_, r_93__7_, r_93__6_, r_93__5_, r_93__4_, r_93__3_, r_93__2_, r_93__1_, r_93__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N185)? data_i : 1'b0;
  assign N184 = sel_i[184];
  assign N185 = N976;
  assign { r_n_93__31_, r_n_93__30_, r_n_93__29_, r_n_93__28_, r_n_93__27_, r_n_93__26_, r_n_93__25_, r_n_93__24_, r_n_93__23_, r_n_93__22_, r_n_93__21_, r_n_93__20_, r_n_93__19_, r_n_93__18_, r_n_93__17_, r_n_93__16_, r_n_93__15_, r_n_93__14_, r_n_93__13_, r_n_93__12_, r_n_93__11_, r_n_93__10_, r_n_93__9_, r_n_93__8_, r_n_93__7_, r_n_93__6_, r_n_93__5_, r_n_93__4_, r_n_93__3_, r_n_93__2_, r_n_93__1_, r_n_93__0_ } = (N186)? { r_94__31_, r_94__30_, r_94__29_, r_94__28_, r_94__27_, r_94__26_, r_94__25_, r_94__24_, r_94__23_, r_94__22_, r_94__21_, r_94__20_, r_94__19_, r_94__18_, r_94__17_, r_94__16_, r_94__15_, r_94__14_, r_94__13_, r_94__12_, r_94__11_, r_94__10_, r_94__9_, r_94__8_, r_94__7_, r_94__6_, r_94__5_, r_94__4_, r_94__3_, r_94__2_, r_94__1_, r_94__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N187)? data_i : 1'b0;
  assign N186 = sel_i[186];
  assign N187 = N981;
  assign { r_n_94__31_, r_n_94__30_, r_n_94__29_, r_n_94__28_, r_n_94__27_, r_n_94__26_, r_n_94__25_, r_n_94__24_, r_n_94__23_, r_n_94__22_, r_n_94__21_, r_n_94__20_, r_n_94__19_, r_n_94__18_, r_n_94__17_, r_n_94__16_, r_n_94__15_, r_n_94__14_, r_n_94__13_, r_n_94__12_, r_n_94__11_, r_n_94__10_, r_n_94__9_, r_n_94__8_, r_n_94__7_, r_n_94__6_, r_n_94__5_, r_n_94__4_, r_n_94__3_, r_n_94__2_, r_n_94__1_, r_n_94__0_ } = (N188)? { r_95__31_, r_95__30_, r_95__29_, r_95__28_, r_95__27_, r_95__26_, r_95__25_, r_95__24_, r_95__23_, r_95__22_, r_95__21_, r_95__20_, r_95__19_, r_95__18_, r_95__17_, r_95__16_, r_95__15_, r_95__14_, r_95__13_, r_95__12_, r_95__11_, r_95__10_, r_95__9_, r_95__8_, r_95__7_, r_95__6_, r_95__5_, r_95__4_, r_95__3_, r_95__2_, r_95__1_, r_95__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N189)? data_i : 1'b0;
  assign N188 = sel_i[188];
  assign N189 = N986;
  assign { r_n_95__31_, r_n_95__30_, r_n_95__29_, r_n_95__28_, r_n_95__27_, r_n_95__26_, r_n_95__25_, r_n_95__24_, r_n_95__23_, r_n_95__22_, r_n_95__21_, r_n_95__20_, r_n_95__19_, r_n_95__18_, r_n_95__17_, r_n_95__16_, r_n_95__15_, r_n_95__14_, r_n_95__13_, r_n_95__12_, r_n_95__11_, r_n_95__10_, r_n_95__9_, r_n_95__8_, r_n_95__7_, r_n_95__6_, r_n_95__5_, r_n_95__4_, r_n_95__3_, r_n_95__2_, r_n_95__1_, r_n_95__0_ } = (N190)? { r_96__31_, r_96__30_, r_96__29_, r_96__28_, r_96__27_, r_96__26_, r_96__25_, r_96__24_, r_96__23_, r_96__22_, r_96__21_, r_96__20_, r_96__19_, r_96__18_, r_96__17_, r_96__16_, r_96__15_, r_96__14_, r_96__13_, r_96__12_, r_96__11_, r_96__10_, r_96__9_, r_96__8_, r_96__7_, r_96__6_, r_96__5_, r_96__4_, r_96__3_, r_96__2_, r_96__1_, r_96__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N191)? data_i : 1'b0;
  assign N190 = sel_i[190];
  assign N191 = N991;
  assign { r_n_96__31_, r_n_96__30_, r_n_96__29_, r_n_96__28_, r_n_96__27_, r_n_96__26_, r_n_96__25_, r_n_96__24_, r_n_96__23_, r_n_96__22_, r_n_96__21_, r_n_96__20_, r_n_96__19_, r_n_96__18_, r_n_96__17_, r_n_96__16_, r_n_96__15_, r_n_96__14_, r_n_96__13_, r_n_96__12_, r_n_96__11_, r_n_96__10_, r_n_96__9_, r_n_96__8_, r_n_96__7_, r_n_96__6_, r_n_96__5_, r_n_96__4_, r_n_96__3_, r_n_96__2_, r_n_96__1_, r_n_96__0_ } = (N192)? { r_97__31_, r_97__30_, r_97__29_, r_97__28_, r_97__27_, r_97__26_, r_97__25_, r_97__24_, r_97__23_, r_97__22_, r_97__21_, r_97__20_, r_97__19_, r_97__18_, r_97__17_, r_97__16_, r_97__15_, r_97__14_, r_97__13_, r_97__12_, r_97__11_, r_97__10_, r_97__9_, r_97__8_, r_97__7_, r_97__6_, r_97__5_, r_97__4_, r_97__3_, r_97__2_, r_97__1_, r_97__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N193)? data_i : 1'b0;
  assign N192 = sel_i[192];
  assign N193 = N996;
  assign { r_n_97__31_, r_n_97__30_, r_n_97__29_, r_n_97__28_, r_n_97__27_, r_n_97__26_, r_n_97__25_, r_n_97__24_, r_n_97__23_, r_n_97__22_, r_n_97__21_, r_n_97__20_, r_n_97__19_, r_n_97__18_, r_n_97__17_, r_n_97__16_, r_n_97__15_, r_n_97__14_, r_n_97__13_, r_n_97__12_, r_n_97__11_, r_n_97__10_, r_n_97__9_, r_n_97__8_, r_n_97__7_, r_n_97__6_, r_n_97__5_, r_n_97__4_, r_n_97__3_, r_n_97__2_, r_n_97__1_, r_n_97__0_ } = (N194)? { r_98__31_, r_98__30_, r_98__29_, r_98__28_, r_98__27_, r_98__26_, r_98__25_, r_98__24_, r_98__23_, r_98__22_, r_98__21_, r_98__20_, r_98__19_, r_98__18_, r_98__17_, r_98__16_, r_98__15_, r_98__14_, r_98__13_, r_98__12_, r_98__11_, r_98__10_, r_98__9_, r_98__8_, r_98__7_, r_98__6_, r_98__5_, r_98__4_, r_98__3_, r_98__2_, r_98__1_, r_98__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N195)? data_i : 1'b0;
  assign N194 = sel_i[194];
  assign N195 = N1001;
  assign { r_n_98__31_, r_n_98__30_, r_n_98__29_, r_n_98__28_, r_n_98__27_, r_n_98__26_, r_n_98__25_, r_n_98__24_, r_n_98__23_, r_n_98__22_, r_n_98__21_, r_n_98__20_, r_n_98__19_, r_n_98__18_, r_n_98__17_, r_n_98__16_, r_n_98__15_, r_n_98__14_, r_n_98__13_, r_n_98__12_, r_n_98__11_, r_n_98__10_, r_n_98__9_, r_n_98__8_, r_n_98__7_, r_n_98__6_, r_n_98__5_, r_n_98__4_, r_n_98__3_, r_n_98__2_, r_n_98__1_, r_n_98__0_ } = (N196)? { r_99__31_, r_99__30_, r_99__29_, r_99__28_, r_99__27_, r_99__26_, r_99__25_, r_99__24_, r_99__23_, r_99__22_, r_99__21_, r_99__20_, r_99__19_, r_99__18_, r_99__17_, r_99__16_, r_99__15_, r_99__14_, r_99__13_, r_99__12_, r_99__11_, r_99__10_, r_99__9_, r_99__8_, r_99__7_, r_99__6_, r_99__5_, r_99__4_, r_99__3_, r_99__2_, r_99__1_, r_99__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N197)? data_i : 1'b0;
  assign N196 = sel_i[196];
  assign N197 = N1006;
  assign { r_n_99__31_, r_n_99__30_, r_n_99__29_, r_n_99__28_, r_n_99__27_, r_n_99__26_, r_n_99__25_, r_n_99__24_, r_n_99__23_, r_n_99__22_, r_n_99__21_, r_n_99__20_, r_n_99__19_, r_n_99__18_, r_n_99__17_, r_n_99__16_, r_n_99__15_, r_n_99__14_, r_n_99__13_, r_n_99__12_, r_n_99__11_, r_n_99__10_, r_n_99__9_, r_n_99__8_, r_n_99__7_, r_n_99__6_, r_n_99__5_, r_n_99__4_, r_n_99__3_, r_n_99__2_, r_n_99__1_, r_n_99__0_ } = (N198)? { r_100__31_, r_100__30_, r_100__29_, r_100__28_, r_100__27_, r_100__26_, r_100__25_, r_100__24_, r_100__23_, r_100__22_, r_100__21_, r_100__20_, r_100__19_, r_100__18_, r_100__17_, r_100__16_, r_100__15_, r_100__14_, r_100__13_, r_100__12_, r_100__11_, r_100__10_, r_100__9_, r_100__8_, r_100__7_, r_100__6_, r_100__5_, r_100__4_, r_100__3_, r_100__2_, r_100__1_, r_100__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                    (N199)? data_i : 1'b0;
  assign N198 = sel_i[198];
  assign N199 = N1011;
  assign { r_n_100__31_, r_n_100__30_, r_n_100__29_, r_n_100__28_, r_n_100__27_, r_n_100__26_, r_n_100__25_, r_n_100__24_, r_n_100__23_, r_n_100__22_, r_n_100__21_, r_n_100__20_, r_n_100__19_, r_n_100__18_, r_n_100__17_, r_n_100__16_, r_n_100__15_, r_n_100__14_, r_n_100__13_, r_n_100__12_, r_n_100__11_, r_n_100__10_, r_n_100__9_, r_n_100__8_, r_n_100__7_, r_n_100__6_, r_n_100__5_, r_n_100__4_, r_n_100__3_, r_n_100__2_, r_n_100__1_, r_n_100__0_ } = (N200)? { r_101__31_, r_101__30_, r_101__29_, r_101__28_, r_101__27_, r_101__26_, r_101__25_, r_101__24_, r_101__23_, r_101__22_, r_101__21_, r_101__20_, r_101__19_, r_101__18_, r_101__17_, r_101__16_, r_101__15_, r_101__14_, r_101__13_, r_101__12_, r_101__11_, r_101__10_, r_101__9_, r_101__8_, r_101__7_, r_101__6_, r_101__5_, r_101__4_, r_101__3_, r_101__2_, r_101__1_, r_101__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N201)? data_i : 1'b0;
  assign N200 = sel_i[200];
  assign N201 = N1016;
  assign { r_n_101__31_, r_n_101__30_, r_n_101__29_, r_n_101__28_, r_n_101__27_, r_n_101__26_, r_n_101__25_, r_n_101__24_, r_n_101__23_, r_n_101__22_, r_n_101__21_, r_n_101__20_, r_n_101__19_, r_n_101__18_, r_n_101__17_, r_n_101__16_, r_n_101__15_, r_n_101__14_, r_n_101__13_, r_n_101__12_, r_n_101__11_, r_n_101__10_, r_n_101__9_, r_n_101__8_, r_n_101__7_, r_n_101__6_, r_n_101__5_, r_n_101__4_, r_n_101__3_, r_n_101__2_, r_n_101__1_, r_n_101__0_ } = (N202)? { r_102__31_, r_102__30_, r_102__29_, r_102__28_, r_102__27_, r_102__26_, r_102__25_, r_102__24_, r_102__23_, r_102__22_, r_102__21_, r_102__20_, r_102__19_, r_102__18_, r_102__17_, r_102__16_, r_102__15_, r_102__14_, r_102__13_, r_102__12_, r_102__11_, r_102__10_, r_102__9_, r_102__8_, r_102__7_, r_102__6_, r_102__5_, r_102__4_, r_102__3_, r_102__2_, r_102__1_, r_102__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N203)? data_i : 1'b0;
  assign N202 = sel_i[202];
  assign N203 = N1021;
  assign { r_n_102__31_, r_n_102__30_, r_n_102__29_, r_n_102__28_, r_n_102__27_, r_n_102__26_, r_n_102__25_, r_n_102__24_, r_n_102__23_, r_n_102__22_, r_n_102__21_, r_n_102__20_, r_n_102__19_, r_n_102__18_, r_n_102__17_, r_n_102__16_, r_n_102__15_, r_n_102__14_, r_n_102__13_, r_n_102__12_, r_n_102__11_, r_n_102__10_, r_n_102__9_, r_n_102__8_, r_n_102__7_, r_n_102__6_, r_n_102__5_, r_n_102__4_, r_n_102__3_, r_n_102__2_, r_n_102__1_, r_n_102__0_ } = (N204)? { r_103__31_, r_103__30_, r_103__29_, r_103__28_, r_103__27_, r_103__26_, r_103__25_, r_103__24_, r_103__23_, r_103__22_, r_103__21_, r_103__20_, r_103__19_, r_103__18_, r_103__17_, r_103__16_, r_103__15_, r_103__14_, r_103__13_, r_103__12_, r_103__11_, r_103__10_, r_103__9_, r_103__8_, r_103__7_, r_103__6_, r_103__5_, r_103__4_, r_103__3_, r_103__2_, r_103__1_, r_103__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N205)? data_i : 1'b0;
  assign N204 = sel_i[204];
  assign N205 = N1026;
  assign { r_n_103__31_, r_n_103__30_, r_n_103__29_, r_n_103__28_, r_n_103__27_, r_n_103__26_, r_n_103__25_, r_n_103__24_, r_n_103__23_, r_n_103__22_, r_n_103__21_, r_n_103__20_, r_n_103__19_, r_n_103__18_, r_n_103__17_, r_n_103__16_, r_n_103__15_, r_n_103__14_, r_n_103__13_, r_n_103__12_, r_n_103__11_, r_n_103__10_, r_n_103__9_, r_n_103__8_, r_n_103__7_, r_n_103__6_, r_n_103__5_, r_n_103__4_, r_n_103__3_, r_n_103__2_, r_n_103__1_, r_n_103__0_ } = (N206)? { r_104__31_, r_104__30_, r_104__29_, r_104__28_, r_104__27_, r_104__26_, r_104__25_, r_104__24_, r_104__23_, r_104__22_, r_104__21_, r_104__20_, r_104__19_, r_104__18_, r_104__17_, r_104__16_, r_104__15_, r_104__14_, r_104__13_, r_104__12_, r_104__11_, r_104__10_, r_104__9_, r_104__8_, r_104__7_, r_104__6_, r_104__5_, r_104__4_, r_104__3_, r_104__2_, r_104__1_, r_104__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N207)? data_i : 1'b0;
  assign N206 = sel_i[206];
  assign N207 = N1031;
  assign { r_n_104__31_, r_n_104__30_, r_n_104__29_, r_n_104__28_, r_n_104__27_, r_n_104__26_, r_n_104__25_, r_n_104__24_, r_n_104__23_, r_n_104__22_, r_n_104__21_, r_n_104__20_, r_n_104__19_, r_n_104__18_, r_n_104__17_, r_n_104__16_, r_n_104__15_, r_n_104__14_, r_n_104__13_, r_n_104__12_, r_n_104__11_, r_n_104__10_, r_n_104__9_, r_n_104__8_, r_n_104__7_, r_n_104__6_, r_n_104__5_, r_n_104__4_, r_n_104__3_, r_n_104__2_, r_n_104__1_, r_n_104__0_ } = (N208)? { r_105__31_, r_105__30_, r_105__29_, r_105__28_, r_105__27_, r_105__26_, r_105__25_, r_105__24_, r_105__23_, r_105__22_, r_105__21_, r_105__20_, r_105__19_, r_105__18_, r_105__17_, r_105__16_, r_105__15_, r_105__14_, r_105__13_, r_105__12_, r_105__11_, r_105__10_, r_105__9_, r_105__8_, r_105__7_, r_105__6_, r_105__5_, r_105__4_, r_105__3_, r_105__2_, r_105__1_, r_105__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N209)? data_i : 1'b0;
  assign N208 = sel_i[208];
  assign N209 = N1036;
  assign { r_n_105__31_, r_n_105__30_, r_n_105__29_, r_n_105__28_, r_n_105__27_, r_n_105__26_, r_n_105__25_, r_n_105__24_, r_n_105__23_, r_n_105__22_, r_n_105__21_, r_n_105__20_, r_n_105__19_, r_n_105__18_, r_n_105__17_, r_n_105__16_, r_n_105__15_, r_n_105__14_, r_n_105__13_, r_n_105__12_, r_n_105__11_, r_n_105__10_, r_n_105__9_, r_n_105__8_, r_n_105__7_, r_n_105__6_, r_n_105__5_, r_n_105__4_, r_n_105__3_, r_n_105__2_, r_n_105__1_, r_n_105__0_ } = (N210)? { r_106__31_, r_106__30_, r_106__29_, r_106__28_, r_106__27_, r_106__26_, r_106__25_, r_106__24_, r_106__23_, r_106__22_, r_106__21_, r_106__20_, r_106__19_, r_106__18_, r_106__17_, r_106__16_, r_106__15_, r_106__14_, r_106__13_, r_106__12_, r_106__11_, r_106__10_, r_106__9_, r_106__8_, r_106__7_, r_106__6_, r_106__5_, r_106__4_, r_106__3_, r_106__2_, r_106__1_, r_106__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N211)? data_i : 1'b0;
  assign N210 = sel_i[210];
  assign N211 = N1041;
  assign { r_n_106__31_, r_n_106__30_, r_n_106__29_, r_n_106__28_, r_n_106__27_, r_n_106__26_, r_n_106__25_, r_n_106__24_, r_n_106__23_, r_n_106__22_, r_n_106__21_, r_n_106__20_, r_n_106__19_, r_n_106__18_, r_n_106__17_, r_n_106__16_, r_n_106__15_, r_n_106__14_, r_n_106__13_, r_n_106__12_, r_n_106__11_, r_n_106__10_, r_n_106__9_, r_n_106__8_, r_n_106__7_, r_n_106__6_, r_n_106__5_, r_n_106__4_, r_n_106__3_, r_n_106__2_, r_n_106__1_, r_n_106__0_ } = (N212)? { r_107__31_, r_107__30_, r_107__29_, r_107__28_, r_107__27_, r_107__26_, r_107__25_, r_107__24_, r_107__23_, r_107__22_, r_107__21_, r_107__20_, r_107__19_, r_107__18_, r_107__17_, r_107__16_, r_107__15_, r_107__14_, r_107__13_, r_107__12_, r_107__11_, r_107__10_, r_107__9_, r_107__8_, r_107__7_, r_107__6_, r_107__5_, r_107__4_, r_107__3_, r_107__2_, r_107__1_, r_107__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N213)? data_i : 1'b0;
  assign N212 = sel_i[212];
  assign N213 = N1046;
  assign { r_n_107__31_, r_n_107__30_, r_n_107__29_, r_n_107__28_, r_n_107__27_, r_n_107__26_, r_n_107__25_, r_n_107__24_, r_n_107__23_, r_n_107__22_, r_n_107__21_, r_n_107__20_, r_n_107__19_, r_n_107__18_, r_n_107__17_, r_n_107__16_, r_n_107__15_, r_n_107__14_, r_n_107__13_, r_n_107__12_, r_n_107__11_, r_n_107__10_, r_n_107__9_, r_n_107__8_, r_n_107__7_, r_n_107__6_, r_n_107__5_, r_n_107__4_, r_n_107__3_, r_n_107__2_, r_n_107__1_, r_n_107__0_ } = (N214)? { r_108__31_, r_108__30_, r_108__29_, r_108__28_, r_108__27_, r_108__26_, r_108__25_, r_108__24_, r_108__23_, r_108__22_, r_108__21_, r_108__20_, r_108__19_, r_108__18_, r_108__17_, r_108__16_, r_108__15_, r_108__14_, r_108__13_, r_108__12_, r_108__11_, r_108__10_, r_108__9_, r_108__8_, r_108__7_, r_108__6_, r_108__5_, r_108__4_, r_108__3_, r_108__2_, r_108__1_, r_108__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N215)? data_i : 1'b0;
  assign N214 = sel_i[214];
  assign N215 = N1051;
  assign { r_n_108__31_, r_n_108__30_, r_n_108__29_, r_n_108__28_, r_n_108__27_, r_n_108__26_, r_n_108__25_, r_n_108__24_, r_n_108__23_, r_n_108__22_, r_n_108__21_, r_n_108__20_, r_n_108__19_, r_n_108__18_, r_n_108__17_, r_n_108__16_, r_n_108__15_, r_n_108__14_, r_n_108__13_, r_n_108__12_, r_n_108__11_, r_n_108__10_, r_n_108__9_, r_n_108__8_, r_n_108__7_, r_n_108__6_, r_n_108__5_, r_n_108__4_, r_n_108__3_, r_n_108__2_, r_n_108__1_, r_n_108__0_ } = (N216)? { r_109__31_, r_109__30_, r_109__29_, r_109__28_, r_109__27_, r_109__26_, r_109__25_, r_109__24_, r_109__23_, r_109__22_, r_109__21_, r_109__20_, r_109__19_, r_109__18_, r_109__17_, r_109__16_, r_109__15_, r_109__14_, r_109__13_, r_109__12_, r_109__11_, r_109__10_, r_109__9_, r_109__8_, r_109__7_, r_109__6_, r_109__5_, r_109__4_, r_109__3_, r_109__2_, r_109__1_, r_109__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N217)? data_i : 1'b0;
  assign N216 = sel_i[216];
  assign N217 = N1056;
  assign { r_n_109__31_, r_n_109__30_, r_n_109__29_, r_n_109__28_, r_n_109__27_, r_n_109__26_, r_n_109__25_, r_n_109__24_, r_n_109__23_, r_n_109__22_, r_n_109__21_, r_n_109__20_, r_n_109__19_, r_n_109__18_, r_n_109__17_, r_n_109__16_, r_n_109__15_, r_n_109__14_, r_n_109__13_, r_n_109__12_, r_n_109__11_, r_n_109__10_, r_n_109__9_, r_n_109__8_, r_n_109__7_, r_n_109__6_, r_n_109__5_, r_n_109__4_, r_n_109__3_, r_n_109__2_, r_n_109__1_, r_n_109__0_ } = (N218)? { r_110__31_, r_110__30_, r_110__29_, r_110__28_, r_110__27_, r_110__26_, r_110__25_, r_110__24_, r_110__23_, r_110__22_, r_110__21_, r_110__20_, r_110__19_, r_110__18_, r_110__17_, r_110__16_, r_110__15_, r_110__14_, r_110__13_, r_110__12_, r_110__11_, r_110__10_, r_110__9_, r_110__8_, r_110__7_, r_110__6_, r_110__5_, r_110__4_, r_110__3_, r_110__2_, r_110__1_, r_110__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N219)? data_i : 1'b0;
  assign N218 = sel_i[218];
  assign N219 = N1061;
  assign { r_n_110__31_, r_n_110__30_, r_n_110__29_, r_n_110__28_, r_n_110__27_, r_n_110__26_, r_n_110__25_, r_n_110__24_, r_n_110__23_, r_n_110__22_, r_n_110__21_, r_n_110__20_, r_n_110__19_, r_n_110__18_, r_n_110__17_, r_n_110__16_, r_n_110__15_, r_n_110__14_, r_n_110__13_, r_n_110__12_, r_n_110__11_, r_n_110__10_, r_n_110__9_, r_n_110__8_, r_n_110__7_, r_n_110__6_, r_n_110__5_, r_n_110__4_, r_n_110__3_, r_n_110__2_, r_n_110__1_, r_n_110__0_ } = (N220)? { r_111__31_, r_111__30_, r_111__29_, r_111__28_, r_111__27_, r_111__26_, r_111__25_, r_111__24_, r_111__23_, r_111__22_, r_111__21_, r_111__20_, r_111__19_, r_111__18_, r_111__17_, r_111__16_, r_111__15_, r_111__14_, r_111__13_, r_111__12_, r_111__11_, r_111__10_, r_111__9_, r_111__8_, r_111__7_, r_111__6_, r_111__5_, r_111__4_, r_111__3_, r_111__2_, r_111__1_, r_111__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N221)? data_i : 1'b0;
  assign N220 = sel_i[220];
  assign N221 = N1066;
  assign { r_n_111__31_, r_n_111__30_, r_n_111__29_, r_n_111__28_, r_n_111__27_, r_n_111__26_, r_n_111__25_, r_n_111__24_, r_n_111__23_, r_n_111__22_, r_n_111__21_, r_n_111__20_, r_n_111__19_, r_n_111__18_, r_n_111__17_, r_n_111__16_, r_n_111__15_, r_n_111__14_, r_n_111__13_, r_n_111__12_, r_n_111__11_, r_n_111__10_, r_n_111__9_, r_n_111__8_, r_n_111__7_, r_n_111__6_, r_n_111__5_, r_n_111__4_, r_n_111__3_, r_n_111__2_, r_n_111__1_, r_n_111__0_ } = (N222)? { r_112__31_, r_112__30_, r_112__29_, r_112__28_, r_112__27_, r_112__26_, r_112__25_, r_112__24_, r_112__23_, r_112__22_, r_112__21_, r_112__20_, r_112__19_, r_112__18_, r_112__17_, r_112__16_, r_112__15_, r_112__14_, r_112__13_, r_112__12_, r_112__11_, r_112__10_, r_112__9_, r_112__8_, r_112__7_, r_112__6_, r_112__5_, r_112__4_, r_112__3_, r_112__2_, r_112__1_, r_112__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N223)? data_i : 1'b0;
  assign N222 = sel_i[222];
  assign N223 = N1071;
  assign { r_n_112__31_, r_n_112__30_, r_n_112__29_, r_n_112__28_, r_n_112__27_, r_n_112__26_, r_n_112__25_, r_n_112__24_, r_n_112__23_, r_n_112__22_, r_n_112__21_, r_n_112__20_, r_n_112__19_, r_n_112__18_, r_n_112__17_, r_n_112__16_, r_n_112__15_, r_n_112__14_, r_n_112__13_, r_n_112__12_, r_n_112__11_, r_n_112__10_, r_n_112__9_, r_n_112__8_, r_n_112__7_, r_n_112__6_, r_n_112__5_, r_n_112__4_, r_n_112__3_, r_n_112__2_, r_n_112__1_, r_n_112__0_ } = (N224)? { r_113__31_, r_113__30_, r_113__29_, r_113__28_, r_113__27_, r_113__26_, r_113__25_, r_113__24_, r_113__23_, r_113__22_, r_113__21_, r_113__20_, r_113__19_, r_113__18_, r_113__17_, r_113__16_, r_113__15_, r_113__14_, r_113__13_, r_113__12_, r_113__11_, r_113__10_, r_113__9_, r_113__8_, r_113__7_, r_113__6_, r_113__5_, r_113__4_, r_113__3_, r_113__2_, r_113__1_, r_113__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N225)? data_i : 1'b0;
  assign N224 = sel_i[224];
  assign N225 = N1076;
  assign { r_n_113__31_, r_n_113__30_, r_n_113__29_, r_n_113__28_, r_n_113__27_, r_n_113__26_, r_n_113__25_, r_n_113__24_, r_n_113__23_, r_n_113__22_, r_n_113__21_, r_n_113__20_, r_n_113__19_, r_n_113__18_, r_n_113__17_, r_n_113__16_, r_n_113__15_, r_n_113__14_, r_n_113__13_, r_n_113__12_, r_n_113__11_, r_n_113__10_, r_n_113__9_, r_n_113__8_, r_n_113__7_, r_n_113__6_, r_n_113__5_, r_n_113__4_, r_n_113__3_, r_n_113__2_, r_n_113__1_, r_n_113__0_ } = (N226)? { r_114__31_, r_114__30_, r_114__29_, r_114__28_, r_114__27_, r_114__26_, r_114__25_, r_114__24_, r_114__23_, r_114__22_, r_114__21_, r_114__20_, r_114__19_, r_114__18_, r_114__17_, r_114__16_, r_114__15_, r_114__14_, r_114__13_, r_114__12_, r_114__11_, r_114__10_, r_114__9_, r_114__8_, r_114__7_, r_114__6_, r_114__5_, r_114__4_, r_114__3_, r_114__2_, r_114__1_, r_114__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N227)? data_i : 1'b0;
  assign N226 = sel_i[226];
  assign N227 = N1081;
  assign { r_n_114__31_, r_n_114__30_, r_n_114__29_, r_n_114__28_, r_n_114__27_, r_n_114__26_, r_n_114__25_, r_n_114__24_, r_n_114__23_, r_n_114__22_, r_n_114__21_, r_n_114__20_, r_n_114__19_, r_n_114__18_, r_n_114__17_, r_n_114__16_, r_n_114__15_, r_n_114__14_, r_n_114__13_, r_n_114__12_, r_n_114__11_, r_n_114__10_, r_n_114__9_, r_n_114__8_, r_n_114__7_, r_n_114__6_, r_n_114__5_, r_n_114__4_, r_n_114__3_, r_n_114__2_, r_n_114__1_, r_n_114__0_ } = (N228)? { r_115__31_, r_115__30_, r_115__29_, r_115__28_, r_115__27_, r_115__26_, r_115__25_, r_115__24_, r_115__23_, r_115__22_, r_115__21_, r_115__20_, r_115__19_, r_115__18_, r_115__17_, r_115__16_, r_115__15_, r_115__14_, r_115__13_, r_115__12_, r_115__11_, r_115__10_, r_115__9_, r_115__8_, r_115__7_, r_115__6_, r_115__5_, r_115__4_, r_115__3_, r_115__2_, r_115__1_, r_115__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N229)? data_i : 1'b0;
  assign N228 = sel_i[228];
  assign N229 = N1086;
  assign { r_n_115__31_, r_n_115__30_, r_n_115__29_, r_n_115__28_, r_n_115__27_, r_n_115__26_, r_n_115__25_, r_n_115__24_, r_n_115__23_, r_n_115__22_, r_n_115__21_, r_n_115__20_, r_n_115__19_, r_n_115__18_, r_n_115__17_, r_n_115__16_, r_n_115__15_, r_n_115__14_, r_n_115__13_, r_n_115__12_, r_n_115__11_, r_n_115__10_, r_n_115__9_, r_n_115__8_, r_n_115__7_, r_n_115__6_, r_n_115__5_, r_n_115__4_, r_n_115__3_, r_n_115__2_, r_n_115__1_, r_n_115__0_ } = (N230)? { r_116__31_, r_116__30_, r_116__29_, r_116__28_, r_116__27_, r_116__26_, r_116__25_, r_116__24_, r_116__23_, r_116__22_, r_116__21_, r_116__20_, r_116__19_, r_116__18_, r_116__17_, r_116__16_, r_116__15_, r_116__14_, r_116__13_, r_116__12_, r_116__11_, r_116__10_, r_116__9_, r_116__8_, r_116__7_, r_116__6_, r_116__5_, r_116__4_, r_116__3_, r_116__2_, r_116__1_, r_116__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N231)? data_i : 1'b0;
  assign N230 = sel_i[230];
  assign N231 = N1091;
  assign { r_n_116__31_, r_n_116__30_, r_n_116__29_, r_n_116__28_, r_n_116__27_, r_n_116__26_, r_n_116__25_, r_n_116__24_, r_n_116__23_, r_n_116__22_, r_n_116__21_, r_n_116__20_, r_n_116__19_, r_n_116__18_, r_n_116__17_, r_n_116__16_, r_n_116__15_, r_n_116__14_, r_n_116__13_, r_n_116__12_, r_n_116__11_, r_n_116__10_, r_n_116__9_, r_n_116__8_, r_n_116__7_, r_n_116__6_, r_n_116__5_, r_n_116__4_, r_n_116__3_, r_n_116__2_, r_n_116__1_, r_n_116__0_ } = (N232)? { r_117__31_, r_117__30_, r_117__29_, r_117__28_, r_117__27_, r_117__26_, r_117__25_, r_117__24_, r_117__23_, r_117__22_, r_117__21_, r_117__20_, r_117__19_, r_117__18_, r_117__17_, r_117__16_, r_117__15_, r_117__14_, r_117__13_, r_117__12_, r_117__11_, r_117__10_, r_117__9_, r_117__8_, r_117__7_, r_117__6_, r_117__5_, r_117__4_, r_117__3_, r_117__2_, r_117__1_, r_117__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N233)? data_i : 1'b0;
  assign N232 = sel_i[232];
  assign N233 = N1096;
  assign { r_n_117__31_, r_n_117__30_, r_n_117__29_, r_n_117__28_, r_n_117__27_, r_n_117__26_, r_n_117__25_, r_n_117__24_, r_n_117__23_, r_n_117__22_, r_n_117__21_, r_n_117__20_, r_n_117__19_, r_n_117__18_, r_n_117__17_, r_n_117__16_, r_n_117__15_, r_n_117__14_, r_n_117__13_, r_n_117__12_, r_n_117__11_, r_n_117__10_, r_n_117__9_, r_n_117__8_, r_n_117__7_, r_n_117__6_, r_n_117__5_, r_n_117__4_, r_n_117__3_, r_n_117__2_, r_n_117__1_, r_n_117__0_ } = (N234)? { r_118__31_, r_118__30_, r_118__29_, r_118__28_, r_118__27_, r_118__26_, r_118__25_, r_118__24_, r_118__23_, r_118__22_, r_118__21_, r_118__20_, r_118__19_, r_118__18_, r_118__17_, r_118__16_, r_118__15_, r_118__14_, r_118__13_, r_118__12_, r_118__11_, r_118__10_, r_118__9_, r_118__8_, r_118__7_, r_118__6_, r_118__5_, r_118__4_, r_118__3_, r_118__2_, r_118__1_, r_118__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N235)? data_i : 1'b0;
  assign N234 = sel_i[234];
  assign N235 = N1101;
  assign { r_n_118__31_, r_n_118__30_, r_n_118__29_, r_n_118__28_, r_n_118__27_, r_n_118__26_, r_n_118__25_, r_n_118__24_, r_n_118__23_, r_n_118__22_, r_n_118__21_, r_n_118__20_, r_n_118__19_, r_n_118__18_, r_n_118__17_, r_n_118__16_, r_n_118__15_, r_n_118__14_, r_n_118__13_, r_n_118__12_, r_n_118__11_, r_n_118__10_, r_n_118__9_, r_n_118__8_, r_n_118__7_, r_n_118__6_, r_n_118__5_, r_n_118__4_, r_n_118__3_, r_n_118__2_, r_n_118__1_, r_n_118__0_ } = (N236)? { r_119__31_, r_119__30_, r_119__29_, r_119__28_, r_119__27_, r_119__26_, r_119__25_, r_119__24_, r_119__23_, r_119__22_, r_119__21_, r_119__20_, r_119__19_, r_119__18_, r_119__17_, r_119__16_, r_119__15_, r_119__14_, r_119__13_, r_119__12_, r_119__11_, r_119__10_, r_119__9_, r_119__8_, r_119__7_, r_119__6_, r_119__5_, r_119__4_, r_119__3_, r_119__2_, r_119__1_, r_119__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N237)? data_i : 1'b0;
  assign N236 = sel_i[236];
  assign N237 = N1106;
  assign { r_n_119__31_, r_n_119__30_, r_n_119__29_, r_n_119__28_, r_n_119__27_, r_n_119__26_, r_n_119__25_, r_n_119__24_, r_n_119__23_, r_n_119__22_, r_n_119__21_, r_n_119__20_, r_n_119__19_, r_n_119__18_, r_n_119__17_, r_n_119__16_, r_n_119__15_, r_n_119__14_, r_n_119__13_, r_n_119__12_, r_n_119__11_, r_n_119__10_, r_n_119__9_, r_n_119__8_, r_n_119__7_, r_n_119__6_, r_n_119__5_, r_n_119__4_, r_n_119__3_, r_n_119__2_, r_n_119__1_, r_n_119__0_ } = (N238)? { r_120__31_, r_120__30_, r_120__29_, r_120__28_, r_120__27_, r_120__26_, r_120__25_, r_120__24_, r_120__23_, r_120__22_, r_120__21_, r_120__20_, r_120__19_, r_120__18_, r_120__17_, r_120__16_, r_120__15_, r_120__14_, r_120__13_, r_120__12_, r_120__11_, r_120__10_, r_120__9_, r_120__8_, r_120__7_, r_120__6_, r_120__5_, r_120__4_, r_120__3_, r_120__2_, r_120__1_, r_120__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N239)? data_i : 1'b0;
  assign N238 = sel_i[238];
  assign N239 = N1111;
  assign { r_n_120__31_, r_n_120__30_, r_n_120__29_, r_n_120__28_, r_n_120__27_, r_n_120__26_, r_n_120__25_, r_n_120__24_, r_n_120__23_, r_n_120__22_, r_n_120__21_, r_n_120__20_, r_n_120__19_, r_n_120__18_, r_n_120__17_, r_n_120__16_, r_n_120__15_, r_n_120__14_, r_n_120__13_, r_n_120__12_, r_n_120__11_, r_n_120__10_, r_n_120__9_, r_n_120__8_, r_n_120__7_, r_n_120__6_, r_n_120__5_, r_n_120__4_, r_n_120__3_, r_n_120__2_, r_n_120__1_, r_n_120__0_ } = (N240)? { r_121__31_, r_121__30_, r_121__29_, r_121__28_, r_121__27_, r_121__26_, r_121__25_, r_121__24_, r_121__23_, r_121__22_, r_121__21_, r_121__20_, r_121__19_, r_121__18_, r_121__17_, r_121__16_, r_121__15_, r_121__14_, r_121__13_, r_121__12_, r_121__11_, r_121__10_, r_121__9_, r_121__8_, r_121__7_, r_121__6_, r_121__5_, r_121__4_, r_121__3_, r_121__2_, r_121__1_, r_121__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N241)? data_i : 1'b0;
  assign N240 = sel_i[240];
  assign N241 = N1116;
  assign { r_n_121__31_, r_n_121__30_, r_n_121__29_, r_n_121__28_, r_n_121__27_, r_n_121__26_, r_n_121__25_, r_n_121__24_, r_n_121__23_, r_n_121__22_, r_n_121__21_, r_n_121__20_, r_n_121__19_, r_n_121__18_, r_n_121__17_, r_n_121__16_, r_n_121__15_, r_n_121__14_, r_n_121__13_, r_n_121__12_, r_n_121__11_, r_n_121__10_, r_n_121__9_, r_n_121__8_, r_n_121__7_, r_n_121__6_, r_n_121__5_, r_n_121__4_, r_n_121__3_, r_n_121__2_, r_n_121__1_, r_n_121__0_ } = (N242)? { r_122__31_, r_122__30_, r_122__29_, r_122__28_, r_122__27_, r_122__26_, r_122__25_, r_122__24_, r_122__23_, r_122__22_, r_122__21_, r_122__20_, r_122__19_, r_122__18_, r_122__17_, r_122__16_, r_122__15_, r_122__14_, r_122__13_, r_122__12_, r_122__11_, r_122__10_, r_122__9_, r_122__8_, r_122__7_, r_122__6_, r_122__5_, r_122__4_, r_122__3_, r_122__2_, r_122__1_, r_122__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N243)? data_i : 1'b0;
  assign N242 = sel_i[242];
  assign N243 = N1121;
  assign { r_n_122__31_, r_n_122__30_, r_n_122__29_, r_n_122__28_, r_n_122__27_, r_n_122__26_, r_n_122__25_, r_n_122__24_, r_n_122__23_, r_n_122__22_, r_n_122__21_, r_n_122__20_, r_n_122__19_, r_n_122__18_, r_n_122__17_, r_n_122__16_, r_n_122__15_, r_n_122__14_, r_n_122__13_, r_n_122__12_, r_n_122__11_, r_n_122__10_, r_n_122__9_, r_n_122__8_, r_n_122__7_, r_n_122__6_, r_n_122__5_, r_n_122__4_, r_n_122__3_, r_n_122__2_, r_n_122__1_, r_n_122__0_ } = (N244)? { r_123__31_, r_123__30_, r_123__29_, r_123__28_, r_123__27_, r_123__26_, r_123__25_, r_123__24_, r_123__23_, r_123__22_, r_123__21_, r_123__20_, r_123__19_, r_123__18_, r_123__17_, r_123__16_, r_123__15_, r_123__14_, r_123__13_, r_123__12_, r_123__11_, r_123__10_, r_123__9_, r_123__8_, r_123__7_, r_123__6_, r_123__5_, r_123__4_, r_123__3_, r_123__2_, r_123__1_, r_123__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N245)? data_i : 1'b0;
  assign N244 = sel_i[244];
  assign N245 = N1126;
  assign { r_n_123__31_, r_n_123__30_, r_n_123__29_, r_n_123__28_, r_n_123__27_, r_n_123__26_, r_n_123__25_, r_n_123__24_, r_n_123__23_, r_n_123__22_, r_n_123__21_, r_n_123__20_, r_n_123__19_, r_n_123__18_, r_n_123__17_, r_n_123__16_, r_n_123__15_, r_n_123__14_, r_n_123__13_, r_n_123__12_, r_n_123__11_, r_n_123__10_, r_n_123__9_, r_n_123__8_, r_n_123__7_, r_n_123__6_, r_n_123__5_, r_n_123__4_, r_n_123__3_, r_n_123__2_, r_n_123__1_, r_n_123__0_ } = (N246)? { r_124__31_, r_124__30_, r_124__29_, r_124__28_, r_124__27_, r_124__26_, r_124__25_, r_124__24_, r_124__23_, r_124__22_, r_124__21_, r_124__20_, r_124__19_, r_124__18_, r_124__17_, r_124__16_, r_124__15_, r_124__14_, r_124__13_, r_124__12_, r_124__11_, r_124__10_, r_124__9_, r_124__8_, r_124__7_, r_124__6_, r_124__5_, r_124__4_, r_124__3_, r_124__2_, r_124__1_, r_124__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N247)? data_i : 1'b0;
  assign N246 = sel_i[246];
  assign N247 = N1131;
  assign { r_n_124__31_, r_n_124__30_, r_n_124__29_, r_n_124__28_, r_n_124__27_, r_n_124__26_, r_n_124__25_, r_n_124__24_, r_n_124__23_, r_n_124__22_, r_n_124__21_, r_n_124__20_, r_n_124__19_, r_n_124__18_, r_n_124__17_, r_n_124__16_, r_n_124__15_, r_n_124__14_, r_n_124__13_, r_n_124__12_, r_n_124__11_, r_n_124__10_, r_n_124__9_, r_n_124__8_, r_n_124__7_, r_n_124__6_, r_n_124__5_, r_n_124__4_, r_n_124__3_, r_n_124__2_, r_n_124__1_, r_n_124__0_ } = (N248)? { r_125__31_, r_125__30_, r_125__29_, r_125__28_, r_125__27_, r_125__26_, r_125__25_, r_125__24_, r_125__23_, r_125__22_, r_125__21_, r_125__20_, r_125__19_, r_125__18_, r_125__17_, r_125__16_, r_125__15_, r_125__14_, r_125__13_, r_125__12_, r_125__11_, r_125__10_, r_125__9_, r_125__8_, r_125__7_, r_125__6_, r_125__5_, r_125__4_, r_125__3_, r_125__2_, r_125__1_, r_125__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N249)? data_i : 1'b0;
  assign N248 = sel_i[248];
  assign N249 = N1136;
  assign { r_n_125__31_, r_n_125__30_, r_n_125__29_, r_n_125__28_, r_n_125__27_, r_n_125__26_, r_n_125__25_, r_n_125__24_, r_n_125__23_, r_n_125__22_, r_n_125__21_, r_n_125__20_, r_n_125__19_, r_n_125__18_, r_n_125__17_, r_n_125__16_, r_n_125__15_, r_n_125__14_, r_n_125__13_, r_n_125__12_, r_n_125__11_, r_n_125__10_, r_n_125__9_, r_n_125__8_, r_n_125__7_, r_n_125__6_, r_n_125__5_, r_n_125__4_, r_n_125__3_, r_n_125__2_, r_n_125__1_, r_n_125__0_ } = (N250)? { r_126__31_, r_126__30_, r_126__29_, r_126__28_, r_126__27_, r_126__26_, r_126__25_, r_126__24_, r_126__23_, r_126__22_, r_126__21_, r_126__20_, r_126__19_, r_126__18_, r_126__17_, r_126__16_, r_126__15_, r_126__14_, r_126__13_, r_126__12_, r_126__11_, r_126__10_, r_126__9_, r_126__8_, r_126__7_, r_126__6_, r_126__5_, r_126__4_, r_126__3_, r_126__2_, r_126__1_, r_126__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N251)? data_i : 1'b0;
  assign N250 = sel_i[250];
  assign N251 = N1141;
  assign { r_n_126__31_, r_n_126__30_, r_n_126__29_, r_n_126__28_, r_n_126__27_, r_n_126__26_, r_n_126__25_, r_n_126__24_, r_n_126__23_, r_n_126__22_, r_n_126__21_, r_n_126__20_, r_n_126__19_, r_n_126__18_, r_n_126__17_, r_n_126__16_, r_n_126__15_, r_n_126__14_, r_n_126__13_, r_n_126__12_, r_n_126__11_, r_n_126__10_, r_n_126__9_, r_n_126__8_, r_n_126__7_, r_n_126__6_, r_n_126__5_, r_n_126__4_, r_n_126__3_, r_n_126__2_, r_n_126__1_, r_n_126__0_ } = (N252)? { r_127__31_, r_127__30_, r_127__29_, r_127__28_, r_127__27_, r_127__26_, r_127__25_, r_127__24_, r_127__23_, r_127__22_, r_127__21_, r_127__20_, r_127__19_, r_127__18_, r_127__17_, r_127__16_, r_127__15_, r_127__14_, r_127__13_, r_127__12_, r_127__11_, r_127__10_, r_127__9_, r_127__8_, r_127__7_, r_127__6_, r_127__5_, r_127__4_, r_127__3_, r_127__2_, r_127__1_, r_127__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N253)? data_i : 1'b0;
  assign N252 = sel_i[252];
  assign N253 = N1146;
  assign { r_n_127__31_, r_n_127__30_, r_n_127__29_, r_n_127__28_, r_n_127__27_, r_n_127__26_, r_n_127__25_, r_n_127__24_, r_n_127__23_, r_n_127__22_, r_n_127__21_, r_n_127__20_, r_n_127__19_, r_n_127__18_, r_n_127__17_, r_n_127__16_, r_n_127__15_, r_n_127__14_, r_n_127__13_, r_n_127__12_, r_n_127__11_, r_n_127__10_, r_n_127__9_, r_n_127__8_, r_n_127__7_, r_n_127__6_, r_n_127__5_, r_n_127__4_, r_n_127__3_, r_n_127__2_, r_n_127__1_, r_n_127__0_ } = (N254)? { r_128__31_, r_128__30_, r_128__29_, r_128__28_, r_128__27_, r_128__26_, r_128__25_, r_128__24_, r_128__23_, r_128__22_, r_128__21_, r_128__20_, r_128__19_, r_128__18_, r_128__17_, r_128__16_, r_128__15_, r_128__14_, r_128__13_, r_128__12_, r_128__11_, r_128__10_, r_128__9_, r_128__8_, r_128__7_, r_128__6_, r_128__5_, r_128__4_, r_128__3_, r_128__2_, r_128__1_, r_128__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N255)? data_i : 1'b0;
  assign N254 = sel_i[254];
  assign N255 = N1151;
  assign { r_n_128__31_, r_n_128__30_, r_n_128__29_, r_n_128__28_, r_n_128__27_, r_n_128__26_, r_n_128__25_, r_n_128__24_, r_n_128__23_, r_n_128__22_, r_n_128__21_, r_n_128__20_, r_n_128__19_, r_n_128__18_, r_n_128__17_, r_n_128__16_, r_n_128__15_, r_n_128__14_, r_n_128__13_, r_n_128__12_, r_n_128__11_, r_n_128__10_, r_n_128__9_, r_n_128__8_, r_n_128__7_, r_n_128__6_, r_n_128__5_, r_n_128__4_, r_n_128__3_, r_n_128__2_, r_n_128__1_, r_n_128__0_ } = (N256)? { r_129__31_, r_129__30_, r_129__29_, r_129__28_, r_129__27_, r_129__26_, r_129__25_, r_129__24_, r_129__23_, r_129__22_, r_129__21_, r_129__20_, r_129__19_, r_129__18_, r_129__17_, r_129__16_, r_129__15_, r_129__14_, r_129__13_, r_129__12_, r_129__11_, r_129__10_, r_129__9_, r_129__8_, r_129__7_, r_129__6_, r_129__5_, r_129__4_, r_129__3_, r_129__2_, r_129__1_, r_129__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N257)? data_i : 1'b0;
  assign N256 = sel_i[256];
  assign N257 = N1156;
  assign { r_n_129__31_, r_n_129__30_, r_n_129__29_, r_n_129__28_, r_n_129__27_, r_n_129__26_, r_n_129__25_, r_n_129__24_, r_n_129__23_, r_n_129__22_, r_n_129__21_, r_n_129__20_, r_n_129__19_, r_n_129__18_, r_n_129__17_, r_n_129__16_, r_n_129__15_, r_n_129__14_, r_n_129__13_, r_n_129__12_, r_n_129__11_, r_n_129__10_, r_n_129__9_, r_n_129__8_, r_n_129__7_, r_n_129__6_, r_n_129__5_, r_n_129__4_, r_n_129__3_, r_n_129__2_, r_n_129__1_, r_n_129__0_ } = (N258)? { r_130__31_, r_130__30_, r_130__29_, r_130__28_, r_130__27_, r_130__26_, r_130__25_, r_130__24_, r_130__23_, r_130__22_, r_130__21_, r_130__20_, r_130__19_, r_130__18_, r_130__17_, r_130__16_, r_130__15_, r_130__14_, r_130__13_, r_130__12_, r_130__11_, r_130__10_, r_130__9_, r_130__8_, r_130__7_, r_130__6_, r_130__5_, r_130__4_, r_130__3_, r_130__2_, r_130__1_, r_130__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N259)? data_i : 1'b0;
  assign N258 = sel_i[258];
  assign N259 = N1161;
  assign { r_n_130__31_, r_n_130__30_, r_n_130__29_, r_n_130__28_, r_n_130__27_, r_n_130__26_, r_n_130__25_, r_n_130__24_, r_n_130__23_, r_n_130__22_, r_n_130__21_, r_n_130__20_, r_n_130__19_, r_n_130__18_, r_n_130__17_, r_n_130__16_, r_n_130__15_, r_n_130__14_, r_n_130__13_, r_n_130__12_, r_n_130__11_, r_n_130__10_, r_n_130__9_, r_n_130__8_, r_n_130__7_, r_n_130__6_, r_n_130__5_, r_n_130__4_, r_n_130__3_, r_n_130__2_, r_n_130__1_, r_n_130__0_ } = (N260)? { r_131__31_, r_131__30_, r_131__29_, r_131__28_, r_131__27_, r_131__26_, r_131__25_, r_131__24_, r_131__23_, r_131__22_, r_131__21_, r_131__20_, r_131__19_, r_131__18_, r_131__17_, r_131__16_, r_131__15_, r_131__14_, r_131__13_, r_131__12_, r_131__11_, r_131__10_, r_131__9_, r_131__8_, r_131__7_, r_131__6_, r_131__5_, r_131__4_, r_131__3_, r_131__2_, r_131__1_, r_131__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N261)? data_i : 1'b0;
  assign N260 = sel_i[260];
  assign N261 = N1166;
  assign { r_n_131__31_, r_n_131__30_, r_n_131__29_, r_n_131__28_, r_n_131__27_, r_n_131__26_, r_n_131__25_, r_n_131__24_, r_n_131__23_, r_n_131__22_, r_n_131__21_, r_n_131__20_, r_n_131__19_, r_n_131__18_, r_n_131__17_, r_n_131__16_, r_n_131__15_, r_n_131__14_, r_n_131__13_, r_n_131__12_, r_n_131__11_, r_n_131__10_, r_n_131__9_, r_n_131__8_, r_n_131__7_, r_n_131__6_, r_n_131__5_, r_n_131__4_, r_n_131__3_, r_n_131__2_, r_n_131__1_, r_n_131__0_ } = (N262)? { r_132__31_, r_132__30_, r_132__29_, r_132__28_, r_132__27_, r_132__26_, r_132__25_, r_132__24_, r_132__23_, r_132__22_, r_132__21_, r_132__20_, r_132__19_, r_132__18_, r_132__17_, r_132__16_, r_132__15_, r_132__14_, r_132__13_, r_132__12_, r_132__11_, r_132__10_, r_132__9_, r_132__8_, r_132__7_, r_132__6_, r_132__5_, r_132__4_, r_132__3_, r_132__2_, r_132__1_, r_132__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N263)? data_i : 1'b0;
  assign N262 = sel_i[262];
  assign N263 = N1171;
  assign { r_n_132__31_, r_n_132__30_, r_n_132__29_, r_n_132__28_, r_n_132__27_, r_n_132__26_, r_n_132__25_, r_n_132__24_, r_n_132__23_, r_n_132__22_, r_n_132__21_, r_n_132__20_, r_n_132__19_, r_n_132__18_, r_n_132__17_, r_n_132__16_, r_n_132__15_, r_n_132__14_, r_n_132__13_, r_n_132__12_, r_n_132__11_, r_n_132__10_, r_n_132__9_, r_n_132__8_, r_n_132__7_, r_n_132__6_, r_n_132__5_, r_n_132__4_, r_n_132__3_, r_n_132__2_, r_n_132__1_, r_n_132__0_ } = (N264)? { r_133__31_, r_133__30_, r_133__29_, r_133__28_, r_133__27_, r_133__26_, r_133__25_, r_133__24_, r_133__23_, r_133__22_, r_133__21_, r_133__20_, r_133__19_, r_133__18_, r_133__17_, r_133__16_, r_133__15_, r_133__14_, r_133__13_, r_133__12_, r_133__11_, r_133__10_, r_133__9_, r_133__8_, r_133__7_, r_133__6_, r_133__5_, r_133__4_, r_133__3_, r_133__2_, r_133__1_, r_133__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N265)? data_i : 1'b0;
  assign N264 = sel_i[264];
  assign N265 = N1176;
  assign { r_n_133__31_, r_n_133__30_, r_n_133__29_, r_n_133__28_, r_n_133__27_, r_n_133__26_, r_n_133__25_, r_n_133__24_, r_n_133__23_, r_n_133__22_, r_n_133__21_, r_n_133__20_, r_n_133__19_, r_n_133__18_, r_n_133__17_, r_n_133__16_, r_n_133__15_, r_n_133__14_, r_n_133__13_, r_n_133__12_, r_n_133__11_, r_n_133__10_, r_n_133__9_, r_n_133__8_, r_n_133__7_, r_n_133__6_, r_n_133__5_, r_n_133__4_, r_n_133__3_, r_n_133__2_, r_n_133__1_, r_n_133__0_ } = (N266)? { r_134__31_, r_134__30_, r_134__29_, r_134__28_, r_134__27_, r_134__26_, r_134__25_, r_134__24_, r_134__23_, r_134__22_, r_134__21_, r_134__20_, r_134__19_, r_134__18_, r_134__17_, r_134__16_, r_134__15_, r_134__14_, r_134__13_, r_134__12_, r_134__11_, r_134__10_, r_134__9_, r_134__8_, r_134__7_, r_134__6_, r_134__5_, r_134__4_, r_134__3_, r_134__2_, r_134__1_, r_134__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N267)? data_i : 1'b0;
  assign N266 = sel_i[266];
  assign N267 = N1181;
  assign { r_n_134__31_, r_n_134__30_, r_n_134__29_, r_n_134__28_, r_n_134__27_, r_n_134__26_, r_n_134__25_, r_n_134__24_, r_n_134__23_, r_n_134__22_, r_n_134__21_, r_n_134__20_, r_n_134__19_, r_n_134__18_, r_n_134__17_, r_n_134__16_, r_n_134__15_, r_n_134__14_, r_n_134__13_, r_n_134__12_, r_n_134__11_, r_n_134__10_, r_n_134__9_, r_n_134__8_, r_n_134__7_, r_n_134__6_, r_n_134__5_, r_n_134__4_, r_n_134__3_, r_n_134__2_, r_n_134__1_, r_n_134__0_ } = (N268)? { r_135__31_, r_135__30_, r_135__29_, r_135__28_, r_135__27_, r_135__26_, r_135__25_, r_135__24_, r_135__23_, r_135__22_, r_135__21_, r_135__20_, r_135__19_, r_135__18_, r_135__17_, r_135__16_, r_135__15_, r_135__14_, r_135__13_, r_135__12_, r_135__11_, r_135__10_, r_135__9_, r_135__8_, r_135__7_, r_135__6_, r_135__5_, r_135__4_, r_135__3_, r_135__2_, r_135__1_, r_135__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N269)? data_i : 1'b0;
  assign N268 = sel_i[268];
  assign N269 = N1186;
  assign { r_n_135__31_, r_n_135__30_, r_n_135__29_, r_n_135__28_, r_n_135__27_, r_n_135__26_, r_n_135__25_, r_n_135__24_, r_n_135__23_, r_n_135__22_, r_n_135__21_, r_n_135__20_, r_n_135__19_, r_n_135__18_, r_n_135__17_, r_n_135__16_, r_n_135__15_, r_n_135__14_, r_n_135__13_, r_n_135__12_, r_n_135__11_, r_n_135__10_, r_n_135__9_, r_n_135__8_, r_n_135__7_, r_n_135__6_, r_n_135__5_, r_n_135__4_, r_n_135__3_, r_n_135__2_, r_n_135__1_, r_n_135__0_ } = (N270)? { r_136__31_, r_136__30_, r_136__29_, r_136__28_, r_136__27_, r_136__26_, r_136__25_, r_136__24_, r_136__23_, r_136__22_, r_136__21_, r_136__20_, r_136__19_, r_136__18_, r_136__17_, r_136__16_, r_136__15_, r_136__14_, r_136__13_, r_136__12_, r_136__11_, r_136__10_, r_136__9_, r_136__8_, r_136__7_, r_136__6_, r_136__5_, r_136__4_, r_136__3_, r_136__2_, r_136__1_, r_136__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N271)? data_i : 1'b0;
  assign N270 = sel_i[270];
  assign N271 = N1191;
  assign { r_n_136__31_, r_n_136__30_, r_n_136__29_, r_n_136__28_, r_n_136__27_, r_n_136__26_, r_n_136__25_, r_n_136__24_, r_n_136__23_, r_n_136__22_, r_n_136__21_, r_n_136__20_, r_n_136__19_, r_n_136__18_, r_n_136__17_, r_n_136__16_, r_n_136__15_, r_n_136__14_, r_n_136__13_, r_n_136__12_, r_n_136__11_, r_n_136__10_, r_n_136__9_, r_n_136__8_, r_n_136__7_, r_n_136__6_, r_n_136__5_, r_n_136__4_, r_n_136__3_, r_n_136__2_, r_n_136__1_, r_n_136__0_ } = (N272)? { r_137__31_, r_137__30_, r_137__29_, r_137__28_, r_137__27_, r_137__26_, r_137__25_, r_137__24_, r_137__23_, r_137__22_, r_137__21_, r_137__20_, r_137__19_, r_137__18_, r_137__17_, r_137__16_, r_137__15_, r_137__14_, r_137__13_, r_137__12_, r_137__11_, r_137__10_, r_137__9_, r_137__8_, r_137__7_, r_137__6_, r_137__5_, r_137__4_, r_137__3_, r_137__2_, r_137__1_, r_137__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N273)? data_i : 1'b0;
  assign N272 = sel_i[272];
  assign N273 = N1196;
  assign { r_n_137__31_, r_n_137__30_, r_n_137__29_, r_n_137__28_, r_n_137__27_, r_n_137__26_, r_n_137__25_, r_n_137__24_, r_n_137__23_, r_n_137__22_, r_n_137__21_, r_n_137__20_, r_n_137__19_, r_n_137__18_, r_n_137__17_, r_n_137__16_, r_n_137__15_, r_n_137__14_, r_n_137__13_, r_n_137__12_, r_n_137__11_, r_n_137__10_, r_n_137__9_, r_n_137__8_, r_n_137__7_, r_n_137__6_, r_n_137__5_, r_n_137__4_, r_n_137__3_, r_n_137__2_, r_n_137__1_, r_n_137__0_ } = (N274)? { r_138__31_, r_138__30_, r_138__29_, r_138__28_, r_138__27_, r_138__26_, r_138__25_, r_138__24_, r_138__23_, r_138__22_, r_138__21_, r_138__20_, r_138__19_, r_138__18_, r_138__17_, r_138__16_, r_138__15_, r_138__14_, r_138__13_, r_138__12_, r_138__11_, r_138__10_, r_138__9_, r_138__8_, r_138__7_, r_138__6_, r_138__5_, r_138__4_, r_138__3_, r_138__2_, r_138__1_, r_138__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N275)? data_i : 1'b0;
  assign N274 = sel_i[274];
  assign N275 = N1201;
  assign { r_n_138__31_, r_n_138__30_, r_n_138__29_, r_n_138__28_, r_n_138__27_, r_n_138__26_, r_n_138__25_, r_n_138__24_, r_n_138__23_, r_n_138__22_, r_n_138__21_, r_n_138__20_, r_n_138__19_, r_n_138__18_, r_n_138__17_, r_n_138__16_, r_n_138__15_, r_n_138__14_, r_n_138__13_, r_n_138__12_, r_n_138__11_, r_n_138__10_, r_n_138__9_, r_n_138__8_, r_n_138__7_, r_n_138__6_, r_n_138__5_, r_n_138__4_, r_n_138__3_, r_n_138__2_, r_n_138__1_, r_n_138__0_ } = (N276)? { r_139__31_, r_139__30_, r_139__29_, r_139__28_, r_139__27_, r_139__26_, r_139__25_, r_139__24_, r_139__23_, r_139__22_, r_139__21_, r_139__20_, r_139__19_, r_139__18_, r_139__17_, r_139__16_, r_139__15_, r_139__14_, r_139__13_, r_139__12_, r_139__11_, r_139__10_, r_139__9_, r_139__8_, r_139__7_, r_139__6_, r_139__5_, r_139__4_, r_139__3_, r_139__2_, r_139__1_, r_139__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N277)? data_i : 1'b0;
  assign N276 = sel_i[276];
  assign N277 = N1206;
  assign { r_n_139__31_, r_n_139__30_, r_n_139__29_, r_n_139__28_, r_n_139__27_, r_n_139__26_, r_n_139__25_, r_n_139__24_, r_n_139__23_, r_n_139__22_, r_n_139__21_, r_n_139__20_, r_n_139__19_, r_n_139__18_, r_n_139__17_, r_n_139__16_, r_n_139__15_, r_n_139__14_, r_n_139__13_, r_n_139__12_, r_n_139__11_, r_n_139__10_, r_n_139__9_, r_n_139__8_, r_n_139__7_, r_n_139__6_, r_n_139__5_, r_n_139__4_, r_n_139__3_, r_n_139__2_, r_n_139__1_, r_n_139__0_ } = (N278)? { r_140__31_, r_140__30_, r_140__29_, r_140__28_, r_140__27_, r_140__26_, r_140__25_, r_140__24_, r_140__23_, r_140__22_, r_140__21_, r_140__20_, r_140__19_, r_140__18_, r_140__17_, r_140__16_, r_140__15_, r_140__14_, r_140__13_, r_140__12_, r_140__11_, r_140__10_, r_140__9_, r_140__8_, r_140__7_, r_140__6_, r_140__5_, r_140__4_, r_140__3_, r_140__2_, r_140__1_, r_140__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N279)? data_i : 1'b0;
  assign N278 = sel_i[278];
  assign N279 = N1211;
  assign { r_n_140__31_, r_n_140__30_, r_n_140__29_, r_n_140__28_, r_n_140__27_, r_n_140__26_, r_n_140__25_, r_n_140__24_, r_n_140__23_, r_n_140__22_, r_n_140__21_, r_n_140__20_, r_n_140__19_, r_n_140__18_, r_n_140__17_, r_n_140__16_, r_n_140__15_, r_n_140__14_, r_n_140__13_, r_n_140__12_, r_n_140__11_, r_n_140__10_, r_n_140__9_, r_n_140__8_, r_n_140__7_, r_n_140__6_, r_n_140__5_, r_n_140__4_, r_n_140__3_, r_n_140__2_, r_n_140__1_, r_n_140__0_ } = (N280)? { r_141__31_, r_141__30_, r_141__29_, r_141__28_, r_141__27_, r_141__26_, r_141__25_, r_141__24_, r_141__23_, r_141__22_, r_141__21_, r_141__20_, r_141__19_, r_141__18_, r_141__17_, r_141__16_, r_141__15_, r_141__14_, r_141__13_, r_141__12_, r_141__11_, r_141__10_, r_141__9_, r_141__8_, r_141__7_, r_141__6_, r_141__5_, r_141__4_, r_141__3_, r_141__2_, r_141__1_, r_141__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N281)? data_i : 1'b0;
  assign N280 = sel_i[280];
  assign N281 = N1216;
  assign { r_n_141__31_, r_n_141__30_, r_n_141__29_, r_n_141__28_, r_n_141__27_, r_n_141__26_, r_n_141__25_, r_n_141__24_, r_n_141__23_, r_n_141__22_, r_n_141__21_, r_n_141__20_, r_n_141__19_, r_n_141__18_, r_n_141__17_, r_n_141__16_, r_n_141__15_, r_n_141__14_, r_n_141__13_, r_n_141__12_, r_n_141__11_, r_n_141__10_, r_n_141__9_, r_n_141__8_, r_n_141__7_, r_n_141__6_, r_n_141__5_, r_n_141__4_, r_n_141__3_, r_n_141__2_, r_n_141__1_, r_n_141__0_ } = (N282)? { r_142__31_, r_142__30_, r_142__29_, r_142__28_, r_142__27_, r_142__26_, r_142__25_, r_142__24_, r_142__23_, r_142__22_, r_142__21_, r_142__20_, r_142__19_, r_142__18_, r_142__17_, r_142__16_, r_142__15_, r_142__14_, r_142__13_, r_142__12_, r_142__11_, r_142__10_, r_142__9_, r_142__8_, r_142__7_, r_142__6_, r_142__5_, r_142__4_, r_142__3_, r_142__2_, r_142__1_, r_142__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N283)? data_i : 1'b0;
  assign N282 = sel_i[282];
  assign N283 = N1221;
  assign { r_n_142__31_, r_n_142__30_, r_n_142__29_, r_n_142__28_, r_n_142__27_, r_n_142__26_, r_n_142__25_, r_n_142__24_, r_n_142__23_, r_n_142__22_, r_n_142__21_, r_n_142__20_, r_n_142__19_, r_n_142__18_, r_n_142__17_, r_n_142__16_, r_n_142__15_, r_n_142__14_, r_n_142__13_, r_n_142__12_, r_n_142__11_, r_n_142__10_, r_n_142__9_, r_n_142__8_, r_n_142__7_, r_n_142__6_, r_n_142__5_, r_n_142__4_, r_n_142__3_, r_n_142__2_, r_n_142__1_, r_n_142__0_ } = (N284)? { r_143__31_, r_143__30_, r_143__29_, r_143__28_, r_143__27_, r_143__26_, r_143__25_, r_143__24_, r_143__23_, r_143__22_, r_143__21_, r_143__20_, r_143__19_, r_143__18_, r_143__17_, r_143__16_, r_143__15_, r_143__14_, r_143__13_, r_143__12_, r_143__11_, r_143__10_, r_143__9_, r_143__8_, r_143__7_, r_143__6_, r_143__5_, r_143__4_, r_143__3_, r_143__2_, r_143__1_, r_143__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N285)? data_i : 1'b0;
  assign N284 = sel_i[284];
  assign N285 = N1226;
  assign { r_n_143__31_, r_n_143__30_, r_n_143__29_, r_n_143__28_, r_n_143__27_, r_n_143__26_, r_n_143__25_, r_n_143__24_, r_n_143__23_, r_n_143__22_, r_n_143__21_, r_n_143__20_, r_n_143__19_, r_n_143__18_, r_n_143__17_, r_n_143__16_, r_n_143__15_, r_n_143__14_, r_n_143__13_, r_n_143__12_, r_n_143__11_, r_n_143__10_, r_n_143__9_, r_n_143__8_, r_n_143__7_, r_n_143__6_, r_n_143__5_, r_n_143__4_, r_n_143__3_, r_n_143__2_, r_n_143__1_, r_n_143__0_ } = (N286)? { r_144__31_, r_144__30_, r_144__29_, r_144__28_, r_144__27_, r_144__26_, r_144__25_, r_144__24_, r_144__23_, r_144__22_, r_144__21_, r_144__20_, r_144__19_, r_144__18_, r_144__17_, r_144__16_, r_144__15_, r_144__14_, r_144__13_, r_144__12_, r_144__11_, r_144__10_, r_144__9_, r_144__8_, r_144__7_, r_144__6_, r_144__5_, r_144__4_, r_144__3_, r_144__2_, r_144__1_, r_144__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N287)? data_i : 1'b0;
  assign N286 = sel_i[286];
  assign N287 = N1231;
  assign { r_n_144__31_, r_n_144__30_, r_n_144__29_, r_n_144__28_, r_n_144__27_, r_n_144__26_, r_n_144__25_, r_n_144__24_, r_n_144__23_, r_n_144__22_, r_n_144__21_, r_n_144__20_, r_n_144__19_, r_n_144__18_, r_n_144__17_, r_n_144__16_, r_n_144__15_, r_n_144__14_, r_n_144__13_, r_n_144__12_, r_n_144__11_, r_n_144__10_, r_n_144__9_, r_n_144__8_, r_n_144__7_, r_n_144__6_, r_n_144__5_, r_n_144__4_, r_n_144__3_, r_n_144__2_, r_n_144__1_, r_n_144__0_ } = (N288)? { r_145__31_, r_145__30_, r_145__29_, r_145__28_, r_145__27_, r_145__26_, r_145__25_, r_145__24_, r_145__23_, r_145__22_, r_145__21_, r_145__20_, r_145__19_, r_145__18_, r_145__17_, r_145__16_, r_145__15_, r_145__14_, r_145__13_, r_145__12_, r_145__11_, r_145__10_, r_145__9_, r_145__8_, r_145__7_, r_145__6_, r_145__5_, r_145__4_, r_145__3_, r_145__2_, r_145__1_, r_145__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N289)? data_i : 1'b0;
  assign N288 = sel_i[288];
  assign N289 = N1236;
  assign { r_n_145__31_, r_n_145__30_, r_n_145__29_, r_n_145__28_, r_n_145__27_, r_n_145__26_, r_n_145__25_, r_n_145__24_, r_n_145__23_, r_n_145__22_, r_n_145__21_, r_n_145__20_, r_n_145__19_, r_n_145__18_, r_n_145__17_, r_n_145__16_, r_n_145__15_, r_n_145__14_, r_n_145__13_, r_n_145__12_, r_n_145__11_, r_n_145__10_, r_n_145__9_, r_n_145__8_, r_n_145__7_, r_n_145__6_, r_n_145__5_, r_n_145__4_, r_n_145__3_, r_n_145__2_, r_n_145__1_, r_n_145__0_ } = (N290)? { r_146__31_, r_146__30_, r_146__29_, r_146__28_, r_146__27_, r_146__26_, r_146__25_, r_146__24_, r_146__23_, r_146__22_, r_146__21_, r_146__20_, r_146__19_, r_146__18_, r_146__17_, r_146__16_, r_146__15_, r_146__14_, r_146__13_, r_146__12_, r_146__11_, r_146__10_, r_146__9_, r_146__8_, r_146__7_, r_146__6_, r_146__5_, r_146__4_, r_146__3_, r_146__2_, r_146__1_, r_146__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N291)? data_i : 1'b0;
  assign N290 = sel_i[290];
  assign N291 = N1241;
  assign { r_n_146__31_, r_n_146__30_, r_n_146__29_, r_n_146__28_, r_n_146__27_, r_n_146__26_, r_n_146__25_, r_n_146__24_, r_n_146__23_, r_n_146__22_, r_n_146__21_, r_n_146__20_, r_n_146__19_, r_n_146__18_, r_n_146__17_, r_n_146__16_, r_n_146__15_, r_n_146__14_, r_n_146__13_, r_n_146__12_, r_n_146__11_, r_n_146__10_, r_n_146__9_, r_n_146__8_, r_n_146__7_, r_n_146__6_, r_n_146__5_, r_n_146__4_, r_n_146__3_, r_n_146__2_, r_n_146__1_, r_n_146__0_ } = (N292)? { r_147__31_, r_147__30_, r_147__29_, r_147__28_, r_147__27_, r_147__26_, r_147__25_, r_147__24_, r_147__23_, r_147__22_, r_147__21_, r_147__20_, r_147__19_, r_147__18_, r_147__17_, r_147__16_, r_147__15_, r_147__14_, r_147__13_, r_147__12_, r_147__11_, r_147__10_, r_147__9_, r_147__8_, r_147__7_, r_147__6_, r_147__5_, r_147__4_, r_147__3_, r_147__2_, r_147__1_, r_147__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N293)? data_i : 1'b0;
  assign N292 = sel_i[292];
  assign N293 = N1246;
  assign { r_n_147__31_, r_n_147__30_, r_n_147__29_, r_n_147__28_, r_n_147__27_, r_n_147__26_, r_n_147__25_, r_n_147__24_, r_n_147__23_, r_n_147__22_, r_n_147__21_, r_n_147__20_, r_n_147__19_, r_n_147__18_, r_n_147__17_, r_n_147__16_, r_n_147__15_, r_n_147__14_, r_n_147__13_, r_n_147__12_, r_n_147__11_, r_n_147__10_, r_n_147__9_, r_n_147__8_, r_n_147__7_, r_n_147__6_, r_n_147__5_, r_n_147__4_, r_n_147__3_, r_n_147__2_, r_n_147__1_, r_n_147__0_ } = (N294)? { r_148__31_, r_148__30_, r_148__29_, r_148__28_, r_148__27_, r_148__26_, r_148__25_, r_148__24_, r_148__23_, r_148__22_, r_148__21_, r_148__20_, r_148__19_, r_148__18_, r_148__17_, r_148__16_, r_148__15_, r_148__14_, r_148__13_, r_148__12_, r_148__11_, r_148__10_, r_148__9_, r_148__8_, r_148__7_, r_148__6_, r_148__5_, r_148__4_, r_148__3_, r_148__2_, r_148__1_, r_148__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N295)? data_i : 1'b0;
  assign N294 = sel_i[294];
  assign N295 = N1251;
  assign { r_n_148__31_, r_n_148__30_, r_n_148__29_, r_n_148__28_, r_n_148__27_, r_n_148__26_, r_n_148__25_, r_n_148__24_, r_n_148__23_, r_n_148__22_, r_n_148__21_, r_n_148__20_, r_n_148__19_, r_n_148__18_, r_n_148__17_, r_n_148__16_, r_n_148__15_, r_n_148__14_, r_n_148__13_, r_n_148__12_, r_n_148__11_, r_n_148__10_, r_n_148__9_, r_n_148__8_, r_n_148__7_, r_n_148__6_, r_n_148__5_, r_n_148__4_, r_n_148__3_, r_n_148__2_, r_n_148__1_, r_n_148__0_ } = (N296)? { r_149__31_, r_149__30_, r_149__29_, r_149__28_, r_149__27_, r_149__26_, r_149__25_, r_149__24_, r_149__23_, r_149__22_, r_149__21_, r_149__20_, r_149__19_, r_149__18_, r_149__17_, r_149__16_, r_149__15_, r_149__14_, r_149__13_, r_149__12_, r_149__11_, r_149__10_, r_149__9_, r_149__8_, r_149__7_, r_149__6_, r_149__5_, r_149__4_, r_149__3_, r_149__2_, r_149__1_, r_149__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N297)? data_i : 1'b0;
  assign N296 = sel_i[296];
  assign N297 = N1256;
  assign { r_n_149__31_, r_n_149__30_, r_n_149__29_, r_n_149__28_, r_n_149__27_, r_n_149__26_, r_n_149__25_, r_n_149__24_, r_n_149__23_, r_n_149__22_, r_n_149__21_, r_n_149__20_, r_n_149__19_, r_n_149__18_, r_n_149__17_, r_n_149__16_, r_n_149__15_, r_n_149__14_, r_n_149__13_, r_n_149__12_, r_n_149__11_, r_n_149__10_, r_n_149__9_, r_n_149__8_, r_n_149__7_, r_n_149__6_, r_n_149__5_, r_n_149__4_, r_n_149__3_, r_n_149__2_, r_n_149__1_, r_n_149__0_ } = (N298)? { r_150__31_, r_150__30_, r_150__29_, r_150__28_, r_150__27_, r_150__26_, r_150__25_, r_150__24_, r_150__23_, r_150__22_, r_150__21_, r_150__20_, r_150__19_, r_150__18_, r_150__17_, r_150__16_, r_150__15_, r_150__14_, r_150__13_, r_150__12_, r_150__11_, r_150__10_, r_150__9_, r_150__8_, r_150__7_, r_150__6_, r_150__5_, r_150__4_, r_150__3_, r_150__2_, r_150__1_, r_150__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N299)? data_i : 1'b0;
  assign N298 = sel_i[298];
  assign N299 = N1261;
  assign { r_n_150__31_, r_n_150__30_, r_n_150__29_, r_n_150__28_, r_n_150__27_, r_n_150__26_, r_n_150__25_, r_n_150__24_, r_n_150__23_, r_n_150__22_, r_n_150__21_, r_n_150__20_, r_n_150__19_, r_n_150__18_, r_n_150__17_, r_n_150__16_, r_n_150__15_, r_n_150__14_, r_n_150__13_, r_n_150__12_, r_n_150__11_, r_n_150__10_, r_n_150__9_, r_n_150__8_, r_n_150__7_, r_n_150__6_, r_n_150__5_, r_n_150__4_, r_n_150__3_, r_n_150__2_, r_n_150__1_, r_n_150__0_ } = (N300)? { r_151__31_, r_151__30_, r_151__29_, r_151__28_, r_151__27_, r_151__26_, r_151__25_, r_151__24_, r_151__23_, r_151__22_, r_151__21_, r_151__20_, r_151__19_, r_151__18_, r_151__17_, r_151__16_, r_151__15_, r_151__14_, r_151__13_, r_151__12_, r_151__11_, r_151__10_, r_151__9_, r_151__8_, r_151__7_, r_151__6_, r_151__5_, r_151__4_, r_151__3_, r_151__2_, r_151__1_, r_151__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N301)? data_i : 1'b0;
  assign N300 = sel_i[300];
  assign N301 = N1266;
  assign { r_n_151__31_, r_n_151__30_, r_n_151__29_, r_n_151__28_, r_n_151__27_, r_n_151__26_, r_n_151__25_, r_n_151__24_, r_n_151__23_, r_n_151__22_, r_n_151__21_, r_n_151__20_, r_n_151__19_, r_n_151__18_, r_n_151__17_, r_n_151__16_, r_n_151__15_, r_n_151__14_, r_n_151__13_, r_n_151__12_, r_n_151__11_, r_n_151__10_, r_n_151__9_, r_n_151__8_, r_n_151__7_, r_n_151__6_, r_n_151__5_, r_n_151__4_, r_n_151__3_, r_n_151__2_, r_n_151__1_, r_n_151__0_ } = (N302)? { r_152__31_, r_152__30_, r_152__29_, r_152__28_, r_152__27_, r_152__26_, r_152__25_, r_152__24_, r_152__23_, r_152__22_, r_152__21_, r_152__20_, r_152__19_, r_152__18_, r_152__17_, r_152__16_, r_152__15_, r_152__14_, r_152__13_, r_152__12_, r_152__11_, r_152__10_, r_152__9_, r_152__8_, r_152__7_, r_152__6_, r_152__5_, r_152__4_, r_152__3_, r_152__2_, r_152__1_, r_152__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N303)? data_i : 1'b0;
  assign N302 = sel_i[302];
  assign N303 = N1271;
  assign { r_n_152__31_, r_n_152__30_, r_n_152__29_, r_n_152__28_, r_n_152__27_, r_n_152__26_, r_n_152__25_, r_n_152__24_, r_n_152__23_, r_n_152__22_, r_n_152__21_, r_n_152__20_, r_n_152__19_, r_n_152__18_, r_n_152__17_, r_n_152__16_, r_n_152__15_, r_n_152__14_, r_n_152__13_, r_n_152__12_, r_n_152__11_, r_n_152__10_, r_n_152__9_, r_n_152__8_, r_n_152__7_, r_n_152__6_, r_n_152__5_, r_n_152__4_, r_n_152__3_, r_n_152__2_, r_n_152__1_, r_n_152__0_ } = (N304)? { r_153__31_, r_153__30_, r_153__29_, r_153__28_, r_153__27_, r_153__26_, r_153__25_, r_153__24_, r_153__23_, r_153__22_, r_153__21_, r_153__20_, r_153__19_, r_153__18_, r_153__17_, r_153__16_, r_153__15_, r_153__14_, r_153__13_, r_153__12_, r_153__11_, r_153__10_, r_153__9_, r_153__8_, r_153__7_, r_153__6_, r_153__5_, r_153__4_, r_153__3_, r_153__2_, r_153__1_, r_153__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N305)? data_i : 1'b0;
  assign N304 = sel_i[304];
  assign N305 = N1276;
  assign { r_n_153__31_, r_n_153__30_, r_n_153__29_, r_n_153__28_, r_n_153__27_, r_n_153__26_, r_n_153__25_, r_n_153__24_, r_n_153__23_, r_n_153__22_, r_n_153__21_, r_n_153__20_, r_n_153__19_, r_n_153__18_, r_n_153__17_, r_n_153__16_, r_n_153__15_, r_n_153__14_, r_n_153__13_, r_n_153__12_, r_n_153__11_, r_n_153__10_, r_n_153__9_, r_n_153__8_, r_n_153__7_, r_n_153__6_, r_n_153__5_, r_n_153__4_, r_n_153__3_, r_n_153__2_, r_n_153__1_, r_n_153__0_ } = (N306)? { r_154__31_, r_154__30_, r_154__29_, r_154__28_, r_154__27_, r_154__26_, r_154__25_, r_154__24_, r_154__23_, r_154__22_, r_154__21_, r_154__20_, r_154__19_, r_154__18_, r_154__17_, r_154__16_, r_154__15_, r_154__14_, r_154__13_, r_154__12_, r_154__11_, r_154__10_, r_154__9_, r_154__8_, r_154__7_, r_154__6_, r_154__5_, r_154__4_, r_154__3_, r_154__2_, r_154__1_, r_154__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N307)? data_i : 1'b0;
  assign N306 = sel_i[306];
  assign N307 = N1281;
  assign { r_n_154__31_, r_n_154__30_, r_n_154__29_, r_n_154__28_, r_n_154__27_, r_n_154__26_, r_n_154__25_, r_n_154__24_, r_n_154__23_, r_n_154__22_, r_n_154__21_, r_n_154__20_, r_n_154__19_, r_n_154__18_, r_n_154__17_, r_n_154__16_, r_n_154__15_, r_n_154__14_, r_n_154__13_, r_n_154__12_, r_n_154__11_, r_n_154__10_, r_n_154__9_, r_n_154__8_, r_n_154__7_, r_n_154__6_, r_n_154__5_, r_n_154__4_, r_n_154__3_, r_n_154__2_, r_n_154__1_, r_n_154__0_ } = (N308)? { r_155__31_, r_155__30_, r_155__29_, r_155__28_, r_155__27_, r_155__26_, r_155__25_, r_155__24_, r_155__23_, r_155__22_, r_155__21_, r_155__20_, r_155__19_, r_155__18_, r_155__17_, r_155__16_, r_155__15_, r_155__14_, r_155__13_, r_155__12_, r_155__11_, r_155__10_, r_155__9_, r_155__8_, r_155__7_, r_155__6_, r_155__5_, r_155__4_, r_155__3_, r_155__2_, r_155__1_, r_155__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N309)? data_i : 1'b0;
  assign N308 = sel_i[308];
  assign N309 = N1286;
  assign { r_n_155__31_, r_n_155__30_, r_n_155__29_, r_n_155__28_, r_n_155__27_, r_n_155__26_, r_n_155__25_, r_n_155__24_, r_n_155__23_, r_n_155__22_, r_n_155__21_, r_n_155__20_, r_n_155__19_, r_n_155__18_, r_n_155__17_, r_n_155__16_, r_n_155__15_, r_n_155__14_, r_n_155__13_, r_n_155__12_, r_n_155__11_, r_n_155__10_, r_n_155__9_, r_n_155__8_, r_n_155__7_, r_n_155__6_, r_n_155__5_, r_n_155__4_, r_n_155__3_, r_n_155__2_, r_n_155__1_, r_n_155__0_ } = (N310)? { r_156__31_, r_156__30_, r_156__29_, r_156__28_, r_156__27_, r_156__26_, r_156__25_, r_156__24_, r_156__23_, r_156__22_, r_156__21_, r_156__20_, r_156__19_, r_156__18_, r_156__17_, r_156__16_, r_156__15_, r_156__14_, r_156__13_, r_156__12_, r_156__11_, r_156__10_, r_156__9_, r_156__8_, r_156__7_, r_156__6_, r_156__5_, r_156__4_, r_156__3_, r_156__2_, r_156__1_, r_156__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N311)? data_i : 1'b0;
  assign N310 = sel_i[310];
  assign N311 = N1291;
  assign { r_n_156__31_, r_n_156__30_, r_n_156__29_, r_n_156__28_, r_n_156__27_, r_n_156__26_, r_n_156__25_, r_n_156__24_, r_n_156__23_, r_n_156__22_, r_n_156__21_, r_n_156__20_, r_n_156__19_, r_n_156__18_, r_n_156__17_, r_n_156__16_, r_n_156__15_, r_n_156__14_, r_n_156__13_, r_n_156__12_, r_n_156__11_, r_n_156__10_, r_n_156__9_, r_n_156__8_, r_n_156__7_, r_n_156__6_, r_n_156__5_, r_n_156__4_, r_n_156__3_, r_n_156__2_, r_n_156__1_, r_n_156__0_ } = (N312)? { r_157__31_, r_157__30_, r_157__29_, r_157__28_, r_157__27_, r_157__26_, r_157__25_, r_157__24_, r_157__23_, r_157__22_, r_157__21_, r_157__20_, r_157__19_, r_157__18_, r_157__17_, r_157__16_, r_157__15_, r_157__14_, r_157__13_, r_157__12_, r_157__11_, r_157__10_, r_157__9_, r_157__8_, r_157__7_, r_157__6_, r_157__5_, r_157__4_, r_157__3_, r_157__2_, r_157__1_, r_157__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N313)? data_i : 1'b0;
  assign N312 = sel_i[312];
  assign N313 = N1296;
  assign { r_n_157__31_, r_n_157__30_, r_n_157__29_, r_n_157__28_, r_n_157__27_, r_n_157__26_, r_n_157__25_, r_n_157__24_, r_n_157__23_, r_n_157__22_, r_n_157__21_, r_n_157__20_, r_n_157__19_, r_n_157__18_, r_n_157__17_, r_n_157__16_, r_n_157__15_, r_n_157__14_, r_n_157__13_, r_n_157__12_, r_n_157__11_, r_n_157__10_, r_n_157__9_, r_n_157__8_, r_n_157__7_, r_n_157__6_, r_n_157__5_, r_n_157__4_, r_n_157__3_, r_n_157__2_, r_n_157__1_, r_n_157__0_ } = (N314)? { r_158__31_, r_158__30_, r_158__29_, r_158__28_, r_158__27_, r_158__26_, r_158__25_, r_158__24_, r_158__23_, r_158__22_, r_158__21_, r_158__20_, r_158__19_, r_158__18_, r_158__17_, r_158__16_, r_158__15_, r_158__14_, r_158__13_, r_158__12_, r_158__11_, r_158__10_, r_158__9_, r_158__8_, r_158__7_, r_158__6_, r_158__5_, r_158__4_, r_158__3_, r_158__2_, r_158__1_, r_158__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N315)? data_i : 1'b0;
  assign N314 = sel_i[314];
  assign N315 = N1301;
  assign { r_n_158__31_, r_n_158__30_, r_n_158__29_, r_n_158__28_, r_n_158__27_, r_n_158__26_, r_n_158__25_, r_n_158__24_, r_n_158__23_, r_n_158__22_, r_n_158__21_, r_n_158__20_, r_n_158__19_, r_n_158__18_, r_n_158__17_, r_n_158__16_, r_n_158__15_, r_n_158__14_, r_n_158__13_, r_n_158__12_, r_n_158__11_, r_n_158__10_, r_n_158__9_, r_n_158__8_, r_n_158__7_, r_n_158__6_, r_n_158__5_, r_n_158__4_, r_n_158__3_, r_n_158__2_, r_n_158__1_, r_n_158__0_ } = (N316)? { r_159__31_, r_159__30_, r_159__29_, r_159__28_, r_159__27_, r_159__26_, r_159__25_, r_159__24_, r_159__23_, r_159__22_, r_159__21_, r_159__20_, r_159__19_, r_159__18_, r_159__17_, r_159__16_, r_159__15_, r_159__14_, r_159__13_, r_159__12_, r_159__11_, r_159__10_, r_159__9_, r_159__8_, r_159__7_, r_159__6_, r_159__5_, r_159__4_, r_159__3_, r_159__2_, r_159__1_, r_159__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N317)? data_i : 1'b0;
  assign N316 = sel_i[316];
  assign N317 = N1306;
  assign { r_n_159__31_, r_n_159__30_, r_n_159__29_, r_n_159__28_, r_n_159__27_, r_n_159__26_, r_n_159__25_, r_n_159__24_, r_n_159__23_, r_n_159__22_, r_n_159__21_, r_n_159__20_, r_n_159__19_, r_n_159__18_, r_n_159__17_, r_n_159__16_, r_n_159__15_, r_n_159__14_, r_n_159__13_, r_n_159__12_, r_n_159__11_, r_n_159__10_, r_n_159__9_, r_n_159__8_, r_n_159__7_, r_n_159__6_, r_n_159__5_, r_n_159__4_, r_n_159__3_, r_n_159__2_, r_n_159__1_, r_n_159__0_ } = (N318)? { r_160__31_, r_160__30_, r_160__29_, r_160__28_, r_160__27_, r_160__26_, r_160__25_, r_160__24_, r_160__23_, r_160__22_, r_160__21_, r_160__20_, r_160__19_, r_160__18_, r_160__17_, r_160__16_, r_160__15_, r_160__14_, r_160__13_, r_160__12_, r_160__11_, r_160__10_, r_160__9_, r_160__8_, r_160__7_, r_160__6_, r_160__5_, r_160__4_, r_160__3_, r_160__2_, r_160__1_, r_160__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N319)? data_i : 1'b0;
  assign N318 = sel_i[318];
  assign N319 = N1311;
  assign { r_n_160__31_, r_n_160__30_, r_n_160__29_, r_n_160__28_, r_n_160__27_, r_n_160__26_, r_n_160__25_, r_n_160__24_, r_n_160__23_, r_n_160__22_, r_n_160__21_, r_n_160__20_, r_n_160__19_, r_n_160__18_, r_n_160__17_, r_n_160__16_, r_n_160__15_, r_n_160__14_, r_n_160__13_, r_n_160__12_, r_n_160__11_, r_n_160__10_, r_n_160__9_, r_n_160__8_, r_n_160__7_, r_n_160__6_, r_n_160__5_, r_n_160__4_, r_n_160__3_, r_n_160__2_, r_n_160__1_, r_n_160__0_ } = (N320)? { r_161__31_, r_161__30_, r_161__29_, r_161__28_, r_161__27_, r_161__26_, r_161__25_, r_161__24_, r_161__23_, r_161__22_, r_161__21_, r_161__20_, r_161__19_, r_161__18_, r_161__17_, r_161__16_, r_161__15_, r_161__14_, r_161__13_, r_161__12_, r_161__11_, r_161__10_, r_161__9_, r_161__8_, r_161__7_, r_161__6_, r_161__5_, r_161__4_, r_161__3_, r_161__2_, r_161__1_, r_161__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N321)? data_i : 1'b0;
  assign N320 = sel_i[320];
  assign N321 = N1316;
  assign { r_n_161__31_, r_n_161__30_, r_n_161__29_, r_n_161__28_, r_n_161__27_, r_n_161__26_, r_n_161__25_, r_n_161__24_, r_n_161__23_, r_n_161__22_, r_n_161__21_, r_n_161__20_, r_n_161__19_, r_n_161__18_, r_n_161__17_, r_n_161__16_, r_n_161__15_, r_n_161__14_, r_n_161__13_, r_n_161__12_, r_n_161__11_, r_n_161__10_, r_n_161__9_, r_n_161__8_, r_n_161__7_, r_n_161__6_, r_n_161__5_, r_n_161__4_, r_n_161__3_, r_n_161__2_, r_n_161__1_, r_n_161__0_ } = (N322)? { r_162__31_, r_162__30_, r_162__29_, r_162__28_, r_162__27_, r_162__26_, r_162__25_, r_162__24_, r_162__23_, r_162__22_, r_162__21_, r_162__20_, r_162__19_, r_162__18_, r_162__17_, r_162__16_, r_162__15_, r_162__14_, r_162__13_, r_162__12_, r_162__11_, r_162__10_, r_162__9_, r_162__8_, r_162__7_, r_162__6_, r_162__5_, r_162__4_, r_162__3_, r_162__2_, r_162__1_, r_162__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N323)? data_i : 1'b0;
  assign N322 = sel_i[322];
  assign N323 = N1321;
  assign { r_n_162__31_, r_n_162__30_, r_n_162__29_, r_n_162__28_, r_n_162__27_, r_n_162__26_, r_n_162__25_, r_n_162__24_, r_n_162__23_, r_n_162__22_, r_n_162__21_, r_n_162__20_, r_n_162__19_, r_n_162__18_, r_n_162__17_, r_n_162__16_, r_n_162__15_, r_n_162__14_, r_n_162__13_, r_n_162__12_, r_n_162__11_, r_n_162__10_, r_n_162__9_, r_n_162__8_, r_n_162__7_, r_n_162__6_, r_n_162__5_, r_n_162__4_, r_n_162__3_, r_n_162__2_, r_n_162__1_, r_n_162__0_ } = (N324)? { r_163__31_, r_163__30_, r_163__29_, r_163__28_, r_163__27_, r_163__26_, r_163__25_, r_163__24_, r_163__23_, r_163__22_, r_163__21_, r_163__20_, r_163__19_, r_163__18_, r_163__17_, r_163__16_, r_163__15_, r_163__14_, r_163__13_, r_163__12_, r_163__11_, r_163__10_, r_163__9_, r_163__8_, r_163__7_, r_163__6_, r_163__5_, r_163__4_, r_163__3_, r_163__2_, r_163__1_, r_163__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N325)? data_i : 1'b0;
  assign N324 = sel_i[324];
  assign N325 = N1326;
  assign { r_n_163__31_, r_n_163__30_, r_n_163__29_, r_n_163__28_, r_n_163__27_, r_n_163__26_, r_n_163__25_, r_n_163__24_, r_n_163__23_, r_n_163__22_, r_n_163__21_, r_n_163__20_, r_n_163__19_, r_n_163__18_, r_n_163__17_, r_n_163__16_, r_n_163__15_, r_n_163__14_, r_n_163__13_, r_n_163__12_, r_n_163__11_, r_n_163__10_, r_n_163__9_, r_n_163__8_, r_n_163__7_, r_n_163__6_, r_n_163__5_, r_n_163__4_, r_n_163__3_, r_n_163__2_, r_n_163__1_, r_n_163__0_ } = (N326)? { r_164__31_, r_164__30_, r_164__29_, r_164__28_, r_164__27_, r_164__26_, r_164__25_, r_164__24_, r_164__23_, r_164__22_, r_164__21_, r_164__20_, r_164__19_, r_164__18_, r_164__17_, r_164__16_, r_164__15_, r_164__14_, r_164__13_, r_164__12_, r_164__11_, r_164__10_, r_164__9_, r_164__8_, r_164__7_, r_164__6_, r_164__5_, r_164__4_, r_164__3_, r_164__2_, r_164__1_, r_164__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N327)? data_i : 1'b0;
  assign N326 = sel_i[326];
  assign N327 = N1331;
  assign { r_n_164__31_, r_n_164__30_, r_n_164__29_, r_n_164__28_, r_n_164__27_, r_n_164__26_, r_n_164__25_, r_n_164__24_, r_n_164__23_, r_n_164__22_, r_n_164__21_, r_n_164__20_, r_n_164__19_, r_n_164__18_, r_n_164__17_, r_n_164__16_, r_n_164__15_, r_n_164__14_, r_n_164__13_, r_n_164__12_, r_n_164__11_, r_n_164__10_, r_n_164__9_, r_n_164__8_, r_n_164__7_, r_n_164__6_, r_n_164__5_, r_n_164__4_, r_n_164__3_, r_n_164__2_, r_n_164__1_, r_n_164__0_ } = (N328)? { r_165__31_, r_165__30_, r_165__29_, r_165__28_, r_165__27_, r_165__26_, r_165__25_, r_165__24_, r_165__23_, r_165__22_, r_165__21_, r_165__20_, r_165__19_, r_165__18_, r_165__17_, r_165__16_, r_165__15_, r_165__14_, r_165__13_, r_165__12_, r_165__11_, r_165__10_, r_165__9_, r_165__8_, r_165__7_, r_165__6_, r_165__5_, r_165__4_, r_165__3_, r_165__2_, r_165__1_, r_165__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N329)? data_i : 1'b0;
  assign N328 = sel_i[328];
  assign N329 = N1336;
  assign { r_n_165__31_, r_n_165__30_, r_n_165__29_, r_n_165__28_, r_n_165__27_, r_n_165__26_, r_n_165__25_, r_n_165__24_, r_n_165__23_, r_n_165__22_, r_n_165__21_, r_n_165__20_, r_n_165__19_, r_n_165__18_, r_n_165__17_, r_n_165__16_, r_n_165__15_, r_n_165__14_, r_n_165__13_, r_n_165__12_, r_n_165__11_, r_n_165__10_, r_n_165__9_, r_n_165__8_, r_n_165__7_, r_n_165__6_, r_n_165__5_, r_n_165__4_, r_n_165__3_, r_n_165__2_, r_n_165__1_, r_n_165__0_ } = (N330)? { r_166__31_, r_166__30_, r_166__29_, r_166__28_, r_166__27_, r_166__26_, r_166__25_, r_166__24_, r_166__23_, r_166__22_, r_166__21_, r_166__20_, r_166__19_, r_166__18_, r_166__17_, r_166__16_, r_166__15_, r_166__14_, r_166__13_, r_166__12_, r_166__11_, r_166__10_, r_166__9_, r_166__8_, r_166__7_, r_166__6_, r_166__5_, r_166__4_, r_166__3_, r_166__2_, r_166__1_, r_166__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N331)? data_i : 1'b0;
  assign N330 = sel_i[330];
  assign N331 = N1341;
  assign { r_n_166__31_, r_n_166__30_, r_n_166__29_, r_n_166__28_, r_n_166__27_, r_n_166__26_, r_n_166__25_, r_n_166__24_, r_n_166__23_, r_n_166__22_, r_n_166__21_, r_n_166__20_, r_n_166__19_, r_n_166__18_, r_n_166__17_, r_n_166__16_, r_n_166__15_, r_n_166__14_, r_n_166__13_, r_n_166__12_, r_n_166__11_, r_n_166__10_, r_n_166__9_, r_n_166__8_, r_n_166__7_, r_n_166__6_, r_n_166__5_, r_n_166__4_, r_n_166__3_, r_n_166__2_, r_n_166__1_, r_n_166__0_ } = (N332)? { r_167__31_, r_167__30_, r_167__29_, r_167__28_, r_167__27_, r_167__26_, r_167__25_, r_167__24_, r_167__23_, r_167__22_, r_167__21_, r_167__20_, r_167__19_, r_167__18_, r_167__17_, r_167__16_, r_167__15_, r_167__14_, r_167__13_, r_167__12_, r_167__11_, r_167__10_, r_167__9_, r_167__8_, r_167__7_, r_167__6_, r_167__5_, r_167__4_, r_167__3_, r_167__2_, r_167__1_, r_167__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N333)? data_i : 1'b0;
  assign N332 = sel_i[332];
  assign N333 = N1346;
  assign { r_n_167__31_, r_n_167__30_, r_n_167__29_, r_n_167__28_, r_n_167__27_, r_n_167__26_, r_n_167__25_, r_n_167__24_, r_n_167__23_, r_n_167__22_, r_n_167__21_, r_n_167__20_, r_n_167__19_, r_n_167__18_, r_n_167__17_, r_n_167__16_, r_n_167__15_, r_n_167__14_, r_n_167__13_, r_n_167__12_, r_n_167__11_, r_n_167__10_, r_n_167__9_, r_n_167__8_, r_n_167__7_, r_n_167__6_, r_n_167__5_, r_n_167__4_, r_n_167__3_, r_n_167__2_, r_n_167__1_, r_n_167__0_ } = (N334)? { r_168__31_, r_168__30_, r_168__29_, r_168__28_, r_168__27_, r_168__26_, r_168__25_, r_168__24_, r_168__23_, r_168__22_, r_168__21_, r_168__20_, r_168__19_, r_168__18_, r_168__17_, r_168__16_, r_168__15_, r_168__14_, r_168__13_, r_168__12_, r_168__11_, r_168__10_, r_168__9_, r_168__8_, r_168__7_, r_168__6_, r_168__5_, r_168__4_, r_168__3_, r_168__2_, r_168__1_, r_168__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N335)? data_i : 1'b0;
  assign N334 = sel_i[334];
  assign N335 = N1351;
  assign { r_n_168__31_, r_n_168__30_, r_n_168__29_, r_n_168__28_, r_n_168__27_, r_n_168__26_, r_n_168__25_, r_n_168__24_, r_n_168__23_, r_n_168__22_, r_n_168__21_, r_n_168__20_, r_n_168__19_, r_n_168__18_, r_n_168__17_, r_n_168__16_, r_n_168__15_, r_n_168__14_, r_n_168__13_, r_n_168__12_, r_n_168__11_, r_n_168__10_, r_n_168__9_, r_n_168__8_, r_n_168__7_, r_n_168__6_, r_n_168__5_, r_n_168__4_, r_n_168__3_, r_n_168__2_, r_n_168__1_, r_n_168__0_ } = (N336)? { r_169__31_, r_169__30_, r_169__29_, r_169__28_, r_169__27_, r_169__26_, r_169__25_, r_169__24_, r_169__23_, r_169__22_, r_169__21_, r_169__20_, r_169__19_, r_169__18_, r_169__17_, r_169__16_, r_169__15_, r_169__14_, r_169__13_, r_169__12_, r_169__11_, r_169__10_, r_169__9_, r_169__8_, r_169__7_, r_169__6_, r_169__5_, r_169__4_, r_169__3_, r_169__2_, r_169__1_, r_169__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N337)? data_i : 1'b0;
  assign N336 = sel_i[336];
  assign N337 = N1356;
  assign { r_n_169__31_, r_n_169__30_, r_n_169__29_, r_n_169__28_, r_n_169__27_, r_n_169__26_, r_n_169__25_, r_n_169__24_, r_n_169__23_, r_n_169__22_, r_n_169__21_, r_n_169__20_, r_n_169__19_, r_n_169__18_, r_n_169__17_, r_n_169__16_, r_n_169__15_, r_n_169__14_, r_n_169__13_, r_n_169__12_, r_n_169__11_, r_n_169__10_, r_n_169__9_, r_n_169__8_, r_n_169__7_, r_n_169__6_, r_n_169__5_, r_n_169__4_, r_n_169__3_, r_n_169__2_, r_n_169__1_, r_n_169__0_ } = (N338)? { r_170__31_, r_170__30_, r_170__29_, r_170__28_, r_170__27_, r_170__26_, r_170__25_, r_170__24_, r_170__23_, r_170__22_, r_170__21_, r_170__20_, r_170__19_, r_170__18_, r_170__17_, r_170__16_, r_170__15_, r_170__14_, r_170__13_, r_170__12_, r_170__11_, r_170__10_, r_170__9_, r_170__8_, r_170__7_, r_170__6_, r_170__5_, r_170__4_, r_170__3_, r_170__2_, r_170__1_, r_170__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N339)? data_i : 1'b0;
  assign N338 = sel_i[338];
  assign N339 = N1361;
  assign { r_n_170__31_, r_n_170__30_, r_n_170__29_, r_n_170__28_, r_n_170__27_, r_n_170__26_, r_n_170__25_, r_n_170__24_, r_n_170__23_, r_n_170__22_, r_n_170__21_, r_n_170__20_, r_n_170__19_, r_n_170__18_, r_n_170__17_, r_n_170__16_, r_n_170__15_, r_n_170__14_, r_n_170__13_, r_n_170__12_, r_n_170__11_, r_n_170__10_, r_n_170__9_, r_n_170__8_, r_n_170__7_, r_n_170__6_, r_n_170__5_, r_n_170__4_, r_n_170__3_, r_n_170__2_, r_n_170__1_, r_n_170__0_ } = (N340)? { r_171__31_, r_171__30_, r_171__29_, r_171__28_, r_171__27_, r_171__26_, r_171__25_, r_171__24_, r_171__23_, r_171__22_, r_171__21_, r_171__20_, r_171__19_, r_171__18_, r_171__17_, r_171__16_, r_171__15_, r_171__14_, r_171__13_, r_171__12_, r_171__11_, r_171__10_, r_171__9_, r_171__8_, r_171__7_, r_171__6_, r_171__5_, r_171__4_, r_171__3_, r_171__2_, r_171__1_, r_171__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N341)? data_i : 1'b0;
  assign N340 = sel_i[340];
  assign N341 = N1366;
  assign { r_n_171__31_, r_n_171__30_, r_n_171__29_, r_n_171__28_, r_n_171__27_, r_n_171__26_, r_n_171__25_, r_n_171__24_, r_n_171__23_, r_n_171__22_, r_n_171__21_, r_n_171__20_, r_n_171__19_, r_n_171__18_, r_n_171__17_, r_n_171__16_, r_n_171__15_, r_n_171__14_, r_n_171__13_, r_n_171__12_, r_n_171__11_, r_n_171__10_, r_n_171__9_, r_n_171__8_, r_n_171__7_, r_n_171__6_, r_n_171__5_, r_n_171__4_, r_n_171__3_, r_n_171__2_, r_n_171__1_, r_n_171__0_ } = (N342)? { r_172__31_, r_172__30_, r_172__29_, r_172__28_, r_172__27_, r_172__26_, r_172__25_, r_172__24_, r_172__23_, r_172__22_, r_172__21_, r_172__20_, r_172__19_, r_172__18_, r_172__17_, r_172__16_, r_172__15_, r_172__14_, r_172__13_, r_172__12_, r_172__11_, r_172__10_, r_172__9_, r_172__8_, r_172__7_, r_172__6_, r_172__5_, r_172__4_, r_172__3_, r_172__2_, r_172__1_, r_172__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N343)? data_i : 1'b0;
  assign N342 = sel_i[342];
  assign N343 = N1371;
  assign { r_n_172__31_, r_n_172__30_, r_n_172__29_, r_n_172__28_, r_n_172__27_, r_n_172__26_, r_n_172__25_, r_n_172__24_, r_n_172__23_, r_n_172__22_, r_n_172__21_, r_n_172__20_, r_n_172__19_, r_n_172__18_, r_n_172__17_, r_n_172__16_, r_n_172__15_, r_n_172__14_, r_n_172__13_, r_n_172__12_, r_n_172__11_, r_n_172__10_, r_n_172__9_, r_n_172__8_, r_n_172__7_, r_n_172__6_, r_n_172__5_, r_n_172__4_, r_n_172__3_, r_n_172__2_, r_n_172__1_, r_n_172__0_ } = (N344)? { r_173__31_, r_173__30_, r_173__29_, r_173__28_, r_173__27_, r_173__26_, r_173__25_, r_173__24_, r_173__23_, r_173__22_, r_173__21_, r_173__20_, r_173__19_, r_173__18_, r_173__17_, r_173__16_, r_173__15_, r_173__14_, r_173__13_, r_173__12_, r_173__11_, r_173__10_, r_173__9_, r_173__8_, r_173__7_, r_173__6_, r_173__5_, r_173__4_, r_173__3_, r_173__2_, r_173__1_, r_173__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N345)? data_i : 1'b0;
  assign N344 = sel_i[344];
  assign N345 = N1376;
  assign { r_n_173__31_, r_n_173__30_, r_n_173__29_, r_n_173__28_, r_n_173__27_, r_n_173__26_, r_n_173__25_, r_n_173__24_, r_n_173__23_, r_n_173__22_, r_n_173__21_, r_n_173__20_, r_n_173__19_, r_n_173__18_, r_n_173__17_, r_n_173__16_, r_n_173__15_, r_n_173__14_, r_n_173__13_, r_n_173__12_, r_n_173__11_, r_n_173__10_, r_n_173__9_, r_n_173__8_, r_n_173__7_, r_n_173__6_, r_n_173__5_, r_n_173__4_, r_n_173__3_, r_n_173__2_, r_n_173__1_, r_n_173__0_ } = (N346)? { r_174__31_, r_174__30_, r_174__29_, r_174__28_, r_174__27_, r_174__26_, r_174__25_, r_174__24_, r_174__23_, r_174__22_, r_174__21_, r_174__20_, r_174__19_, r_174__18_, r_174__17_, r_174__16_, r_174__15_, r_174__14_, r_174__13_, r_174__12_, r_174__11_, r_174__10_, r_174__9_, r_174__8_, r_174__7_, r_174__6_, r_174__5_, r_174__4_, r_174__3_, r_174__2_, r_174__1_, r_174__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N347)? data_i : 1'b0;
  assign N346 = sel_i[346];
  assign N347 = N1381;
  assign { r_n_174__31_, r_n_174__30_, r_n_174__29_, r_n_174__28_, r_n_174__27_, r_n_174__26_, r_n_174__25_, r_n_174__24_, r_n_174__23_, r_n_174__22_, r_n_174__21_, r_n_174__20_, r_n_174__19_, r_n_174__18_, r_n_174__17_, r_n_174__16_, r_n_174__15_, r_n_174__14_, r_n_174__13_, r_n_174__12_, r_n_174__11_, r_n_174__10_, r_n_174__9_, r_n_174__8_, r_n_174__7_, r_n_174__6_, r_n_174__5_, r_n_174__4_, r_n_174__3_, r_n_174__2_, r_n_174__1_, r_n_174__0_ } = (N348)? { r_175__31_, r_175__30_, r_175__29_, r_175__28_, r_175__27_, r_175__26_, r_175__25_, r_175__24_, r_175__23_, r_175__22_, r_175__21_, r_175__20_, r_175__19_, r_175__18_, r_175__17_, r_175__16_, r_175__15_, r_175__14_, r_175__13_, r_175__12_, r_175__11_, r_175__10_, r_175__9_, r_175__8_, r_175__7_, r_175__6_, r_175__5_, r_175__4_, r_175__3_, r_175__2_, r_175__1_, r_175__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N349)? data_i : 1'b0;
  assign N348 = sel_i[348];
  assign N349 = N1386;
  assign { r_n_175__31_, r_n_175__30_, r_n_175__29_, r_n_175__28_, r_n_175__27_, r_n_175__26_, r_n_175__25_, r_n_175__24_, r_n_175__23_, r_n_175__22_, r_n_175__21_, r_n_175__20_, r_n_175__19_, r_n_175__18_, r_n_175__17_, r_n_175__16_, r_n_175__15_, r_n_175__14_, r_n_175__13_, r_n_175__12_, r_n_175__11_, r_n_175__10_, r_n_175__9_, r_n_175__8_, r_n_175__7_, r_n_175__6_, r_n_175__5_, r_n_175__4_, r_n_175__3_, r_n_175__2_, r_n_175__1_, r_n_175__0_ } = (N350)? { r_176__31_, r_176__30_, r_176__29_, r_176__28_, r_176__27_, r_176__26_, r_176__25_, r_176__24_, r_176__23_, r_176__22_, r_176__21_, r_176__20_, r_176__19_, r_176__18_, r_176__17_, r_176__16_, r_176__15_, r_176__14_, r_176__13_, r_176__12_, r_176__11_, r_176__10_, r_176__9_, r_176__8_, r_176__7_, r_176__6_, r_176__5_, r_176__4_, r_176__3_, r_176__2_, r_176__1_, r_176__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N351)? data_i : 1'b0;
  assign N350 = sel_i[350];
  assign N351 = N1391;
  assign { r_n_176__31_, r_n_176__30_, r_n_176__29_, r_n_176__28_, r_n_176__27_, r_n_176__26_, r_n_176__25_, r_n_176__24_, r_n_176__23_, r_n_176__22_, r_n_176__21_, r_n_176__20_, r_n_176__19_, r_n_176__18_, r_n_176__17_, r_n_176__16_, r_n_176__15_, r_n_176__14_, r_n_176__13_, r_n_176__12_, r_n_176__11_, r_n_176__10_, r_n_176__9_, r_n_176__8_, r_n_176__7_, r_n_176__6_, r_n_176__5_, r_n_176__4_, r_n_176__3_, r_n_176__2_, r_n_176__1_, r_n_176__0_ } = (N352)? { r_177__31_, r_177__30_, r_177__29_, r_177__28_, r_177__27_, r_177__26_, r_177__25_, r_177__24_, r_177__23_, r_177__22_, r_177__21_, r_177__20_, r_177__19_, r_177__18_, r_177__17_, r_177__16_, r_177__15_, r_177__14_, r_177__13_, r_177__12_, r_177__11_, r_177__10_, r_177__9_, r_177__8_, r_177__7_, r_177__6_, r_177__5_, r_177__4_, r_177__3_, r_177__2_, r_177__1_, r_177__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N353)? data_i : 1'b0;
  assign N352 = sel_i[352];
  assign N353 = N1396;
  assign { r_n_177__31_, r_n_177__30_, r_n_177__29_, r_n_177__28_, r_n_177__27_, r_n_177__26_, r_n_177__25_, r_n_177__24_, r_n_177__23_, r_n_177__22_, r_n_177__21_, r_n_177__20_, r_n_177__19_, r_n_177__18_, r_n_177__17_, r_n_177__16_, r_n_177__15_, r_n_177__14_, r_n_177__13_, r_n_177__12_, r_n_177__11_, r_n_177__10_, r_n_177__9_, r_n_177__8_, r_n_177__7_, r_n_177__6_, r_n_177__5_, r_n_177__4_, r_n_177__3_, r_n_177__2_, r_n_177__1_, r_n_177__0_ } = (N354)? { r_178__31_, r_178__30_, r_178__29_, r_178__28_, r_178__27_, r_178__26_, r_178__25_, r_178__24_, r_178__23_, r_178__22_, r_178__21_, r_178__20_, r_178__19_, r_178__18_, r_178__17_, r_178__16_, r_178__15_, r_178__14_, r_178__13_, r_178__12_, r_178__11_, r_178__10_, r_178__9_, r_178__8_, r_178__7_, r_178__6_, r_178__5_, r_178__4_, r_178__3_, r_178__2_, r_178__1_, r_178__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N355)? data_i : 1'b0;
  assign N354 = sel_i[354];
  assign N355 = N1401;
  assign { r_n_178__31_, r_n_178__30_, r_n_178__29_, r_n_178__28_, r_n_178__27_, r_n_178__26_, r_n_178__25_, r_n_178__24_, r_n_178__23_, r_n_178__22_, r_n_178__21_, r_n_178__20_, r_n_178__19_, r_n_178__18_, r_n_178__17_, r_n_178__16_, r_n_178__15_, r_n_178__14_, r_n_178__13_, r_n_178__12_, r_n_178__11_, r_n_178__10_, r_n_178__9_, r_n_178__8_, r_n_178__7_, r_n_178__6_, r_n_178__5_, r_n_178__4_, r_n_178__3_, r_n_178__2_, r_n_178__1_, r_n_178__0_ } = (N356)? { r_179__31_, r_179__30_, r_179__29_, r_179__28_, r_179__27_, r_179__26_, r_179__25_, r_179__24_, r_179__23_, r_179__22_, r_179__21_, r_179__20_, r_179__19_, r_179__18_, r_179__17_, r_179__16_, r_179__15_, r_179__14_, r_179__13_, r_179__12_, r_179__11_, r_179__10_, r_179__9_, r_179__8_, r_179__7_, r_179__6_, r_179__5_, r_179__4_, r_179__3_, r_179__2_, r_179__1_, r_179__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N357)? data_i : 1'b0;
  assign N356 = sel_i[356];
  assign N357 = N1406;
  assign { r_n_179__31_, r_n_179__30_, r_n_179__29_, r_n_179__28_, r_n_179__27_, r_n_179__26_, r_n_179__25_, r_n_179__24_, r_n_179__23_, r_n_179__22_, r_n_179__21_, r_n_179__20_, r_n_179__19_, r_n_179__18_, r_n_179__17_, r_n_179__16_, r_n_179__15_, r_n_179__14_, r_n_179__13_, r_n_179__12_, r_n_179__11_, r_n_179__10_, r_n_179__9_, r_n_179__8_, r_n_179__7_, r_n_179__6_, r_n_179__5_, r_n_179__4_, r_n_179__3_, r_n_179__2_, r_n_179__1_, r_n_179__0_ } = (N358)? { r_180__31_, r_180__30_, r_180__29_, r_180__28_, r_180__27_, r_180__26_, r_180__25_, r_180__24_, r_180__23_, r_180__22_, r_180__21_, r_180__20_, r_180__19_, r_180__18_, r_180__17_, r_180__16_, r_180__15_, r_180__14_, r_180__13_, r_180__12_, r_180__11_, r_180__10_, r_180__9_, r_180__8_, r_180__7_, r_180__6_, r_180__5_, r_180__4_, r_180__3_, r_180__2_, r_180__1_, r_180__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N359)? data_i : 1'b0;
  assign N358 = sel_i[358];
  assign N359 = N1411;
  assign { r_n_180__31_, r_n_180__30_, r_n_180__29_, r_n_180__28_, r_n_180__27_, r_n_180__26_, r_n_180__25_, r_n_180__24_, r_n_180__23_, r_n_180__22_, r_n_180__21_, r_n_180__20_, r_n_180__19_, r_n_180__18_, r_n_180__17_, r_n_180__16_, r_n_180__15_, r_n_180__14_, r_n_180__13_, r_n_180__12_, r_n_180__11_, r_n_180__10_, r_n_180__9_, r_n_180__8_, r_n_180__7_, r_n_180__6_, r_n_180__5_, r_n_180__4_, r_n_180__3_, r_n_180__2_, r_n_180__1_, r_n_180__0_ } = (N360)? { r_181__31_, r_181__30_, r_181__29_, r_181__28_, r_181__27_, r_181__26_, r_181__25_, r_181__24_, r_181__23_, r_181__22_, r_181__21_, r_181__20_, r_181__19_, r_181__18_, r_181__17_, r_181__16_, r_181__15_, r_181__14_, r_181__13_, r_181__12_, r_181__11_, r_181__10_, r_181__9_, r_181__8_, r_181__7_, r_181__6_, r_181__5_, r_181__4_, r_181__3_, r_181__2_, r_181__1_, r_181__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N361)? data_i : 1'b0;
  assign N360 = sel_i[360];
  assign N361 = N1416;
  assign { r_n_181__31_, r_n_181__30_, r_n_181__29_, r_n_181__28_, r_n_181__27_, r_n_181__26_, r_n_181__25_, r_n_181__24_, r_n_181__23_, r_n_181__22_, r_n_181__21_, r_n_181__20_, r_n_181__19_, r_n_181__18_, r_n_181__17_, r_n_181__16_, r_n_181__15_, r_n_181__14_, r_n_181__13_, r_n_181__12_, r_n_181__11_, r_n_181__10_, r_n_181__9_, r_n_181__8_, r_n_181__7_, r_n_181__6_, r_n_181__5_, r_n_181__4_, r_n_181__3_, r_n_181__2_, r_n_181__1_, r_n_181__0_ } = (N362)? { r_182__31_, r_182__30_, r_182__29_, r_182__28_, r_182__27_, r_182__26_, r_182__25_, r_182__24_, r_182__23_, r_182__22_, r_182__21_, r_182__20_, r_182__19_, r_182__18_, r_182__17_, r_182__16_, r_182__15_, r_182__14_, r_182__13_, r_182__12_, r_182__11_, r_182__10_, r_182__9_, r_182__8_, r_182__7_, r_182__6_, r_182__5_, r_182__4_, r_182__3_, r_182__2_, r_182__1_, r_182__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N363)? data_i : 1'b0;
  assign N362 = sel_i[362];
  assign N363 = N1421;
  assign { r_n_182__31_, r_n_182__30_, r_n_182__29_, r_n_182__28_, r_n_182__27_, r_n_182__26_, r_n_182__25_, r_n_182__24_, r_n_182__23_, r_n_182__22_, r_n_182__21_, r_n_182__20_, r_n_182__19_, r_n_182__18_, r_n_182__17_, r_n_182__16_, r_n_182__15_, r_n_182__14_, r_n_182__13_, r_n_182__12_, r_n_182__11_, r_n_182__10_, r_n_182__9_, r_n_182__8_, r_n_182__7_, r_n_182__6_, r_n_182__5_, r_n_182__4_, r_n_182__3_, r_n_182__2_, r_n_182__1_, r_n_182__0_ } = (N364)? { r_183__31_, r_183__30_, r_183__29_, r_183__28_, r_183__27_, r_183__26_, r_183__25_, r_183__24_, r_183__23_, r_183__22_, r_183__21_, r_183__20_, r_183__19_, r_183__18_, r_183__17_, r_183__16_, r_183__15_, r_183__14_, r_183__13_, r_183__12_, r_183__11_, r_183__10_, r_183__9_, r_183__8_, r_183__7_, r_183__6_, r_183__5_, r_183__4_, r_183__3_, r_183__2_, r_183__1_, r_183__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N365)? data_i : 1'b0;
  assign N364 = sel_i[364];
  assign N365 = N1426;
  assign { r_n_183__31_, r_n_183__30_, r_n_183__29_, r_n_183__28_, r_n_183__27_, r_n_183__26_, r_n_183__25_, r_n_183__24_, r_n_183__23_, r_n_183__22_, r_n_183__21_, r_n_183__20_, r_n_183__19_, r_n_183__18_, r_n_183__17_, r_n_183__16_, r_n_183__15_, r_n_183__14_, r_n_183__13_, r_n_183__12_, r_n_183__11_, r_n_183__10_, r_n_183__9_, r_n_183__8_, r_n_183__7_, r_n_183__6_, r_n_183__5_, r_n_183__4_, r_n_183__3_, r_n_183__2_, r_n_183__1_, r_n_183__0_ } = (N366)? { r_184__31_, r_184__30_, r_184__29_, r_184__28_, r_184__27_, r_184__26_, r_184__25_, r_184__24_, r_184__23_, r_184__22_, r_184__21_, r_184__20_, r_184__19_, r_184__18_, r_184__17_, r_184__16_, r_184__15_, r_184__14_, r_184__13_, r_184__12_, r_184__11_, r_184__10_, r_184__9_, r_184__8_, r_184__7_, r_184__6_, r_184__5_, r_184__4_, r_184__3_, r_184__2_, r_184__1_, r_184__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N367)? data_i : 1'b0;
  assign N366 = sel_i[366];
  assign N367 = N1431;
  assign { r_n_184__31_, r_n_184__30_, r_n_184__29_, r_n_184__28_, r_n_184__27_, r_n_184__26_, r_n_184__25_, r_n_184__24_, r_n_184__23_, r_n_184__22_, r_n_184__21_, r_n_184__20_, r_n_184__19_, r_n_184__18_, r_n_184__17_, r_n_184__16_, r_n_184__15_, r_n_184__14_, r_n_184__13_, r_n_184__12_, r_n_184__11_, r_n_184__10_, r_n_184__9_, r_n_184__8_, r_n_184__7_, r_n_184__6_, r_n_184__5_, r_n_184__4_, r_n_184__3_, r_n_184__2_, r_n_184__1_, r_n_184__0_ } = (N368)? { r_185__31_, r_185__30_, r_185__29_, r_185__28_, r_185__27_, r_185__26_, r_185__25_, r_185__24_, r_185__23_, r_185__22_, r_185__21_, r_185__20_, r_185__19_, r_185__18_, r_185__17_, r_185__16_, r_185__15_, r_185__14_, r_185__13_, r_185__12_, r_185__11_, r_185__10_, r_185__9_, r_185__8_, r_185__7_, r_185__6_, r_185__5_, r_185__4_, r_185__3_, r_185__2_, r_185__1_, r_185__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N369)? data_i : 1'b0;
  assign N368 = sel_i[368];
  assign N369 = N1436;
  assign { r_n_185__31_, r_n_185__30_, r_n_185__29_, r_n_185__28_, r_n_185__27_, r_n_185__26_, r_n_185__25_, r_n_185__24_, r_n_185__23_, r_n_185__22_, r_n_185__21_, r_n_185__20_, r_n_185__19_, r_n_185__18_, r_n_185__17_, r_n_185__16_, r_n_185__15_, r_n_185__14_, r_n_185__13_, r_n_185__12_, r_n_185__11_, r_n_185__10_, r_n_185__9_, r_n_185__8_, r_n_185__7_, r_n_185__6_, r_n_185__5_, r_n_185__4_, r_n_185__3_, r_n_185__2_, r_n_185__1_, r_n_185__0_ } = (N370)? { r_186__31_, r_186__30_, r_186__29_, r_186__28_, r_186__27_, r_186__26_, r_186__25_, r_186__24_, r_186__23_, r_186__22_, r_186__21_, r_186__20_, r_186__19_, r_186__18_, r_186__17_, r_186__16_, r_186__15_, r_186__14_, r_186__13_, r_186__12_, r_186__11_, r_186__10_, r_186__9_, r_186__8_, r_186__7_, r_186__6_, r_186__5_, r_186__4_, r_186__3_, r_186__2_, r_186__1_, r_186__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N371)? data_i : 1'b0;
  assign N370 = sel_i[370];
  assign N371 = N1441;
  assign { r_n_186__31_, r_n_186__30_, r_n_186__29_, r_n_186__28_, r_n_186__27_, r_n_186__26_, r_n_186__25_, r_n_186__24_, r_n_186__23_, r_n_186__22_, r_n_186__21_, r_n_186__20_, r_n_186__19_, r_n_186__18_, r_n_186__17_, r_n_186__16_, r_n_186__15_, r_n_186__14_, r_n_186__13_, r_n_186__12_, r_n_186__11_, r_n_186__10_, r_n_186__9_, r_n_186__8_, r_n_186__7_, r_n_186__6_, r_n_186__5_, r_n_186__4_, r_n_186__3_, r_n_186__2_, r_n_186__1_, r_n_186__0_ } = (N372)? { r_187__31_, r_187__30_, r_187__29_, r_187__28_, r_187__27_, r_187__26_, r_187__25_, r_187__24_, r_187__23_, r_187__22_, r_187__21_, r_187__20_, r_187__19_, r_187__18_, r_187__17_, r_187__16_, r_187__15_, r_187__14_, r_187__13_, r_187__12_, r_187__11_, r_187__10_, r_187__9_, r_187__8_, r_187__7_, r_187__6_, r_187__5_, r_187__4_, r_187__3_, r_187__2_, r_187__1_, r_187__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N373)? data_i : 1'b0;
  assign N372 = sel_i[372];
  assign N373 = N1446;
  assign { r_n_187__31_, r_n_187__30_, r_n_187__29_, r_n_187__28_, r_n_187__27_, r_n_187__26_, r_n_187__25_, r_n_187__24_, r_n_187__23_, r_n_187__22_, r_n_187__21_, r_n_187__20_, r_n_187__19_, r_n_187__18_, r_n_187__17_, r_n_187__16_, r_n_187__15_, r_n_187__14_, r_n_187__13_, r_n_187__12_, r_n_187__11_, r_n_187__10_, r_n_187__9_, r_n_187__8_, r_n_187__7_, r_n_187__6_, r_n_187__5_, r_n_187__4_, r_n_187__3_, r_n_187__2_, r_n_187__1_, r_n_187__0_ } = (N374)? { r_188__31_, r_188__30_, r_188__29_, r_188__28_, r_188__27_, r_188__26_, r_188__25_, r_188__24_, r_188__23_, r_188__22_, r_188__21_, r_188__20_, r_188__19_, r_188__18_, r_188__17_, r_188__16_, r_188__15_, r_188__14_, r_188__13_, r_188__12_, r_188__11_, r_188__10_, r_188__9_, r_188__8_, r_188__7_, r_188__6_, r_188__5_, r_188__4_, r_188__3_, r_188__2_, r_188__1_, r_188__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N375)? data_i : 1'b0;
  assign N374 = sel_i[374];
  assign N375 = N1451;
  assign { r_n_188__31_, r_n_188__30_, r_n_188__29_, r_n_188__28_, r_n_188__27_, r_n_188__26_, r_n_188__25_, r_n_188__24_, r_n_188__23_, r_n_188__22_, r_n_188__21_, r_n_188__20_, r_n_188__19_, r_n_188__18_, r_n_188__17_, r_n_188__16_, r_n_188__15_, r_n_188__14_, r_n_188__13_, r_n_188__12_, r_n_188__11_, r_n_188__10_, r_n_188__9_, r_n_188__8_, r_n_188__7_, r_n_188__6_, r_n_188__5_, r_n_188__4_, r_n_188__3_, r_n_188__2_, r_n_188__1_, r_n_188__0_ } = (N376)? { r_189__31_, r_189__30_, r_189__29_, r_189__28_, r_189__27_, r_189__26_, r_189__25_, r_189__24_, r_189__23_, r_189__22_, r_189__21_, r_189__20_, r_189__19_, r_189__18_, r_189__17_, r_189__16_, r_189__15_, r_189__14_, r_189__13_, r_189__12_, r_189__11_, r_189__10_, r_189__9_, r_189__8_, r_189__7_, r_189__6_, r_189__5_, r_189__4_, r_189__3_, r_189__2_, r_189__1_, r_189__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N377)? data_i : 1'b0;
  assign N376 = sel_i[376];
  assign N377 = N1456;
  assign { r_n_189__31_, r_n_189__30_, r_n_189__29_, r_n_189__28_, r_n_189__27_, r_n_189__26_, r_n_189__25_, r_n_189__24_, r_n_189__23_, r_n_189__22_, r_n_189__21_, r_n_189__20_, r_n_189__19_, r_n_189__18_, r_n_189__17_, r_n_189__16_, r_n_189__15_, r_n_189__14_, r_n_189__13_, r_n_189__12_, r_n_189__11_, r_n_189__10_, r_n_189__9_, r_n_189__8_, r_n_189__7_, r_n_189__6_, r_n_189__5_, r_n_189__4_, r_n_189__3_, r_n_189__2_, r_n_189__1_, r_n_189__0_ } = (N378)? { r_190__31_, r_190__30_, r_190__29_, r_190__28_, r_190__27_, r_190__26_, r_190__25_, r_190__24_, r_190__23_, r_190__22_, r_190__21_, r_190__20_, r_190__19_, r_190__18_, r_190__17_, r_190__16_, r_190__15_, r_190__14_, r_190__13_, r_190__12_, r_190__11_, r_190__10_, r_190__9_, r_190__8_, r_190__7_, r_190__6_, r_190__5_, r_190__4_, r_190__3_, r_190__2_, r_190__1_, r_190__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N379)? data_i : 1'b0;
  assign N378 = sel_i[378];
  assign N379 = N1461;
  assign { r_n_190__31_, r_n_190__30_, r_n_190__29_, r_n_190__28_, r_n_190__27_, r_n_190__26_, r_n_190__25_, r_n_190__24_, r_n_190__23_, r_n_190__22_, r_n_190__21_, r_n_190__20_, r_n_190__19_, r_n_190__18_, r_n_190__17_, r_n_190__16_, r_n_190__15_, r_n_190__14_, r_n_190__13_, r_n_190__12_, r_n_190__11_, r_n_190__10_, r_n_190__9_, r_n_190__8_, r_n_190__7_, r_n_190__6_, r_n_190__5_, r_n_190__4_, r_n_190__3_, r_n_190__2_, r_n_190__1_, r_n_190__0_ } = (N380)? { r_191__31_, r_191__30_, r_191__29_, r_191__28_, r_191__27_, r_191__26_, r_191__25_, r_191__24_, r_191__23_, r_191__22_, r_191__21_, r_191__20_, r_191__19_, r_191__18_, r_191__17_, r_191__16_, r_191__15_, r_191__14_, r_191__13_, r_191__12_, r_191__11_, r_191__10_, r_191__9_, r_191__8_, r_191__7_, r_191__6_, r_191__5_, r_191__4_, r_191__3_, r_191__2_, r_191__1_, r_191__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N381)? data_i : 1'b0;
  assign N380 = sel_i[380];
  assign N381 = N1466;
  assign { r_n_191__31_, r_n_191__30_, r_n_191__29_, r_n_191__28_, r_n_191__27_, r_n_191__26_, r_n_191__25_, r_n_191__24_, r_n_191__23_, r_n_191__22_, r_n_191__21_, r_n_191__20_, r_n_191__19_, r_n_191__18_, r_n_191__17_, r_n_191__16_, r_n_191__15_, r_n_191__14_, r_n_191__13_, r_n_191__12_, r_n_191__11_, r_n_191__10_, r_n_191__9_, r_n_191__8_, r_n_191__7_, r_n_191__6_, r_n_191__5_, r_n_191__4_, r_n_191__3_, r_n_191__2_, r_n_191__1_, r_n_191__0_ } = (N382)? { r_192__31_, r_192__30_, r_192__29_, r_192__28_, r_192__27_, r_192__26_, r_192__25_, r_192__24_, r_192__23_, r_192__22_, r_192__21_, r_192__20_, r_192__19_, r_192__18_, r_192__17_, r_192__16_, r_192__15_, r_192__14_, r_192__13_, r_192__12_, r_192__11_, r_192__10_, r_192__9_, r_192__8_, r_192__7_, r_192__6_, r_192__5_, r_192__4_, r_192__3_, r_192__2_, r_192__1_, r_192__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N383)? data_i : 1'b0;
  assign N382 = sel_i[382];
  assign N383 = N1471;
  assign { r_n_192__31_, r_n_192__30_, r_n_192__29_, r_n_192__28_, r_n_192__27_, r_n_192__26_, r_n_192__25_, r_n_192__24_, r_n_192__23_, r_n_192__22_, r_n_192__21_, r_n_192__20_, r_n_192__19_, r_n_192__18_, r_n_192__17_, r_n_192__16_, r_n_192__15_, r_n_192__14_, r_n_192__13_, r_n_192__12_, r_n_192__11_, r_n_192__10_, r_n_192__9_, r_n_192__8_, r_n_192__7_, r_n_192__6_, r_n_192__5_, r_n_192__4_, r_n_192__3_, r_n_192__2_, r_n_192__1_, r_n_192__0_ } = (N384)? { r_193__31_, r_193__30_, r_193__29_, r_193__28_, r_193__27_, r_193__26_, r_193__25_, r_193__24_, r_193__23_, r_193__22_, r_193__21_, r_193__20_, r_193__19_, r_193__18_, r_193__17_, r_193__16_, r_193__15_, r_193__14_, r_193__13_, r_193__12_, r_193__11_, r_193__10_, r_193__9_, r_193__8_, r_193__7_, r_193__6_, r_193__5_, r_193__4_, r_193__3_, r_193__2_, r_193__1_, r_193__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N385)? data_i : 1'b0;
  assign N384 = sel_i[384];
  assign N385 = N1476;
  assign { r_n_193__31_, r_n_193__30_, r_n_193__29_, r_n_193__28_, r_n_193__27_, r_n_193__26_, r_n_193__25_, r_n_193__24_, r_n_193__23_, r_n_193__22_, r_n_193__21_, r_n_193__20_, r_n_193__19_, r_n_193__18_, r_n_193__17_, r_n_193__16_, r_n_193__15_, r_n_193__14_, r_n_193__13_, r_n_193__12_, r_n_193__11_, r_n_193__10_, r_n_193__9_, r_n_193__8_, r_n_193__7_, r_n_193__6_, r_n_193__5_, r_n_193__4_, r_n_193__3_, r_n_193__2_, r_n_193__1_, r_n_193__0_ } = (N386)? { r_194__31_, r_194__30_, r_194__29_, r_194__28_, r_194__27_, r_194__26_, r_194__25_, r_194__24_, r_194__23_, r_194__22_, r_194__21_, r_194__20_, r_194__19_, r_194__18_, r_194__17_, r_194__16_, r_194__15_, r_194__14_, r_194__13_, r_194__12_, r_194__11_, r_194__10_, r_194__9_, r_194__8_, r_194__7_, r_194__6_, r_194__5_, r_194__4_, r_194__3_, r_194__2_, r_194__1_, r_194__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N387)? data_i : 1'b0;
  assign N386 = sel_i[386];
  assign N387 = N1481;
  assign { r_n_194__31_, r_n_194__30_, r_n_194__29_, r_n_194__28_, r_n_194__27_, r_n_194__26_, r_n_194__25_, r_n_194__24_, r_n_194__23_, r_n_194__22_, r_n_194__21_, r_n_194__20_, r_n_194__19_, r_n_194__18_, r_n_194__17_, r_n_194__16_, r_n_194__15_, r_n_194__14_, r_n_194__13_, r_n_194__12_, r_n_194__11_, r_n_194__10_, r_n_194__9_, r_n_194__8_, r_n_194__7_, r_n_194__6_, r_n_194__5_, r_n_194__4_, r_n_194__3_, r_n_194__2_, r_n_194__1_, r_n_194__0_ } = (N388)? { r_195__31_, r_195__30_, r_195__29_, r_195__28_, r_195__27_, r_195__26_, r_195__25_, r_195__24_, r_195__23_, r_195__22_, r_195__21_, r_195__20_, r_195__19_, r_195__18_, r_195__17_, r_195__16_, r_195__15_, r_195__14_, r_195__13_, r_195__12_, r_195__11_, r_195__10_, r_195__9_, r_195__8_, r_195__7_, r_195__6_, r_195__5_, r_195__4_, r_195__3_, r_195__2_, r_195__1_, r_195__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N389)? data_i : 1'b0;
  assign N388 = sel_i[388];
  assign N389 = N1486;
  assign { r_n_195__31_, r_n_195__30_, r_n_195__29_, r_n_195__28_, r_n_195__27_, r_n_195__26_, r_n_195__25_, r_n_195__24_, r_n_195__23_, r_n_195__22_, r_n_195__21_, r_n_195__20_, r_n_195__19_, r_n_195__18_, r_n_195__17_, r_n_195__16_, r_n_195__15_, r_n_195__14_, r_n_195__13_, r_n_195__12_, r_n_195__11_, r_n_195__10_, r_n_195__9_, r_n_195__8_, r_n_195__7_, r_n_195__6_, r_n_195__5_, r_n_195__4_, r_n_195__3_, r_n_195__2_, r_n_195__1_, r_n_195__0_ } = (N390)? { r_196__31_, r_196__30_, r_196__29_, r_196__28_, r_196__27_, r_196__26_, r_196__25_, r_196__24_, r_196__23_, r_196__22_, r_196__21_, r_196__20_, r_196__19_, r_196__18_, r_196__17_, r_196__16_, r_196__15_, r_196__14_, r_196__13_, r_196__12_, r_196__11_, r_196__10_, r_196__9_, r_196__8_, r_196__7_, r_196__6_, r_196__5_, r_196__4_, r_196__3_, r_196__2_, r_196__1_, r_196__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N391)? data_i : 1'b0;
  assign N390 = sel_i[390];
  assign N391 = N1491;
  assign { r_n_196__31_, r_n_196__30_, r_n_196__29_, r_n_196__28_, r_n_196__27_, r_n_196__26_, r_n_196__25_, r_n_196__24_, r_n_196__23_, r_n_196__22_, r_n_196__21_, r_n_196__20_, r_n_196__19_, r_n_196__18_, r_n_196__17_, r_n_196__16_, r_n_196__15_, r_n_196__14_, r_n_196__13_, r_n_196__12_, r_n_196__11_, r_n_196__10_, r_n_196__9_, r_n_196__8_, r_n_196__7_, r_n_196__6_, r_n_196__5_, r_n_196__4_, r_n_196__3_, r_n_196__2_, r_n_196__1_, r_n_196__0_ } = (N392)? { r_197__31_, r_197__30_, r_197__29_, r_197__28_, r_197__27_, r_197__26_, r_197__25_, r_197__24_, r_197__23_, r_197__22_, r_197__21_, r_197__20_, r_197__19_, r_197__18_, r_197__17_, r_197__16_, r_197__15_, r_197__14_, r_197__13_, r_197__12_, r_197__11_, r_197__10_, r_197__9_, r_197__8_, r_197__7_, r_197__6_, r_197__5_, r_197__4_, r_197__3_, r_197__2_, r_197__1_, r_197__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N393)? data_i : 1'b0;
  assign N392 = sel_i[392];
  assign N393 = N1496;
  assign { r_n_197__31_, r_n_197__30_, r_n_197__29_, r_n_197__28_, r_n_197__27_, r_n_197__26_, r_n_197__25_, r_n_197__24_, r_n_197__23_, r_n_197__22_, r_n_197__21_, r_n_197__20_, r_n_197__19_, r_n_197__18_, r_n_197__17_, r_n_197__16_, r_n_197__15_, r_n_197__14_, r_n_197__13_, r_n_197__12_, r_n_197__11_, r_n_197__10_, r_n_197__9_, r_n_197__8_, r_n_197__7_, r_n_197__6_, r_n_197__5_, r_n_197__4_, r_n_197__3_, r_n_197__2_, r_n_197__1_, r_n_197__0_ } = (N394)? { r_198__31_, r_198__30_, r_198__29_, r_198__28_, r_198__27_, r_198__26_, r_198__25_, r_198__24_, r_198__23_, r_198__22_, r_198__21_, r_198__20_, r_198__19_, r_198__18_, r_198__17_, r_198__16_, r_198__15_, r_198__14_, r_198__13_, r_198__12_, r_198__11_, r_198__10_, r_198__9_, r_198__8_, r_198__7_, r_198__6_, r_198__5_, r_198__4_, r_198__3_, r_198__2_, r_198__1_, r_198__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N395)? data_i : 1'b0;
  assign N394 = sel_i[394];
  assign N395 = N1501;
  assign { r_n_198__31_, r_n_198__30_, r_n_198__29_, r_n_198__28_, r_n_198__27_, r_n_198__26_, r_n_198__25_, r_n_198__24_, r_n_198__23_, r_n_198__22_, r_n_198__21_, r_n_198__20_, r_n_198__19_, r_n_198__18_, r_n_198__17_, r_n_198__16_, r_n_198__15_, r_n_198__14_, r_n_198__13_, r_n_198__12_, r_n_198__11_, r_n_198__10_, r_n_198__9_, r_n_198__8_, r_n_198__7_, r_n_198__6_, r_n_198__5_, r_n_198__4_, r_n_198__3_, r_n_198__2_, r_n_198__1_, r_n_198__0_ } = (N396)? { r_199__31_, r_199__30_, r_199__29_, r_199__28_, r_199__27_, r_199__26_, r_199__25_, r_199__24_, r_199__23_, r_199__22_, r_199__21_, r_199__20_, r_199__19_, r_199__18_, r_199__17_, r_199__16_, r_199__15_, r_199__14_, r_199__13_, r_199__12_, r_199__11_, r_199__10_, r_199__9_, r_199__8_, r_199__7_, r_199__6_, r_199__5_, r_199__4_, r_199__3_, r_199__2_, r_199__1_, r_199__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N397)? data_i : 1'b0;
  assign N396 = sel_i[396];
  assign N397 = N1506;
  assign { r_n_199__31_, r_n_199__30_, r_n_199__29_, r_n_199__28_, r_n_199__27_, r_n_199__26_, r_n_199__25_, r_n_199__24_, r_n_199__23_, r_n_199__22_, r_n_199__21_, r_n_199__20_, r_n_199__19_, r_n_199__18_, r_n_199__17_, r_n_199__16_, r_n_199__15_, r_n_199__14_, r_n_199__13_, r_n_199__12_, r_n_199__11_, r_n_199__10_, r_n_199__9_, r_n_199__8_, r_n_199__7_, r_n_199__6_, r_n_199__5_, r_n_199__4_, r_n_199__3_, r_n_199__2_, r_n_199__1_, r_n_199__0_ } = (N398)? { r_200__31_, r_200__30_, r_200__29_, r_200__28_, r_200__27_, r_200__26_, r_200__25_, r_200__24_, r_200__23_, r_200__22_, r_200__21_, r_200__20_, r_200__19_, r_200__18_, r_200__17_, r_200__16_, r_200__15_, r_200__14_, r_200__13_, r_200__12_, r_200__11_, r_200__10_, r_200__9_, r_200__8_, r_200__7_, r_200__6_, r_200__5_, r_200__4_, r_200__3_, r_200__2_, r_200__1_, r_200__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N399)? data_i : 1'b0;
  assign N398 = sel_i[398];
  assign N399 = N1511;
  assign { r_n_200__31_, r_n_200__30_, r_n_200__29_, r_n_200__28_, r_n_200__27_, r_n_200__26_, r_n_200__25_, r_n_200__24_, r_n_200__23_, r_n_200__22_, r_n_200__21_, r_n_200__20_, r_n_200__19_, r_n_200__18_, r_n_200__17_, r_n_200__16_, r_n_200__15_, r_n_200__14_, r_n_200__13_, r_n_200__12_, r_n_200__11_, r_n_200__10_, r_n_200__9_, r_n_200__8_, r_n_200__7_, r_n_200__6_, r_n_200__5_, r_n_200__4_, r_n_200__3_, r_n_200__2_, r_n_200__1_, r_n_200__0_ } = (N400)? { r_201__31_, r_201__30_, r_201__29_, r_201__28_, r_201__27_, r_201__26_, r_201__25_, r_201__24_, r_201__23_, r_201__22_, r_201__21_, r_201__20_, r_201__19_, r_201__18_, r_201__17_, r_201__16_, r_201__15_, r_201__14_, r_201__13_, r_201__12_, r_201__11_, r_201__10_, r_201__9_, r_201__8_, r_201__7_, r_201__6_, r_201__5_, r_201__4_, r_201__3_, r_201__2_, r_201__1_, r_201__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N401)? data_i : 1'b0;
  assign N400 = sel_i[400];
  assign N401 = N1516;
  assign { r_n_201__31_, r_n_201__30_, r_n_201__29_, r_n_201__28_, r_n_201__27_, r_n_201__26_, r_n_201__25_, r_n_201__24_, r_n_201__23_, r_n_201__22_, r_n_201__21_, r_n_201__20_, r_n_201__19_, r_n_201__18_, r_n_201__17_, r_n_201__16_, r_n_201__15_, r_n_201__14_, r_n_201__13_, r_n_201__12_, r_n_201__11_, r_n_201__10_, r_n_201__9_, r_n_201__8_, r_n_201__7_, r_n_201__6_, r_n_201__5_, r_n_201__4_, r_n_201__3_, r_n_201__2_, r_n_201__1_, r_n_201__0_ } = (N402)? { r_202__31_, r_202__30_, r_202__29_, r_202__28_, r_202__27_, r_202__26_, r_202__25_, r_202__24_, r_202__23_, r_202__22_, r_202__21_, r_202__20_, r_202__19_, r_202__18_, r_202__17_, r_202__16_, r_202__15_, r_202__14_, r_202__13_, r_202__12_, r_202__11_, r_202__10_, r_202__9_, r_202__8_, r_202__7_, r_202__6_, r_202__5_, r_202__4_, r_202__3_, r_202__2_, r_202__1_, r_202__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N403)? data_i : 1'b0;
  assign N402 = sel_i[402];
  assign N403 = N1521;
  assign { r_n_202__31_, r_n_202__30_, r_n_202__29_, r_n_202__28_, r_n_202__27_, r_n_202__26_, r_n_202__25_, r_n_202__24_, r_n_202__23_, r_n_202__22_, r_n_202__21_, r_n_202__20_, r_n_202__19_, r_n_202__18_, r_n_202__17_, r_n_202__16_, r_n_202__15_, r_n_202__14_, r_n_202__13_, r_n_202__12_, r_n_202__11_, r_n_202__10_, r_n_202__9_, r_n_202__8_, r_n_202__7_, r_n_202__6_, r_n_202__5_, r_n_202__4_, r_n_202__3_, r_n_202__2_, r_n_202__1_, r_n_202__0_ } = (N404)? { r_203__31_, r_203__30_, r_203__29_, r_203__28_, r_203__27_, r_203__26_, r_203__25_, r_203__24_, r_203__23_, r_203__22_, r_203__21_, r_203__20_, r_203__19_, r_203__18_, r_203__17_, r_203__16_, r_203__15_, r_203__14_, r_203__13_, r_203__12_, r_203__11_, r_203__10_, r_203__9_, r_203__8_, r_203__7_, r_203__6_, r_203__5_, r_203__4_, r_203__3_, r_203__2_, r_203__1_, r_203__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N405)? data_i : 1'b0;
  assign N404 = sel_i[404];
  assign N405 = N1526;
  assign { r_n_203__31_, r_n_203__30_, r_n_203__29_, r_n_203__28_, r_n_203__27_, r_n_203__26_, r_n_203__25_, r_n_203__24_, r_n_203__23_, r_n_203__22_, r_n_203__21_, r_n_203__20_, r_n_203__19_, r_n_203__18_, r_n_203__17_, r_n_203__16_, r_n_203__15_, r_n_203__14_, r_n_203__13_, r_n_203__12_, r_n_203__11_, r_n_203__10_, r_n_203__9_, r_n_203__8_, r_n_203__7_, r_n_203__6_, r_n_203__5_, r_n_203__4_, r_n_203__3_, r_n_203__2_, r_n_203__1_, r_n_203__0_ } = (N406)? { r_204__31_, r_204__30_, r_204__29_, r_204__28_, r_204__27_, r_204__26_, r_204__25_, r_204__24_, r_204__23_, r_204__22_, r_204__21_, r_204__20_, r_204__19_, r_204__18_, r_204__17_, r_204__16_, r_204__15_, r_204__14_, r_204__13_, r_204__12_, r_204__11_, r_204__10_, r_204__9_, r_204__8_, r_204__7_, r_204__6_, r_204__5_, r_204__4_, r_204__3_, r_204__2_, r_204__1_, r_204__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N407)? data_i : 1'b0;
  assign N406 = sel_i[406];
  assign N407 = N1531;
  assign { r_n_204__31_, r_n_204__30_, r_n_204__29_, r_n_204__28_, r_n_204__27_, r_n_204__26_, r_n_204__25_, r_n_204__24_, r_n_204__23_, r_n_204__22_, r_n_204__21_, r_n_204__20_, r_n_204__19_, r_n_204__18_, r_n_204__17_, r_n_204__16_, r_n_204__15_, r_n_204__14_, r_n_204__13_, r_n_204__12_, r_n_204__11_, r_n_204__10_, r_n_204__9_, r_n_204__8_, r_n_204__7_, r_n_204__6_, r_n_204__5_, r_n_204__4_, r_n_204__3_, r_n_204__2_, r_n_204__1_, r_n_204__0_ } = (N408)? { r_205__31_, r_205__30_, r_205__29_, r_205__28_, r_205__27_, r_205__26_, r_205__25_, r_205__24_, r_205__23_, r_205__22_, r_205__21_, r_205__20_, r_205__19_, r_205__18_, r_205__17_, r_205__16_, r_205__15_, r_205__14_, r_205__13_, r_205__12_, r_205__11_, r_205__10_, r_205__9_, r_205__8_, r_205__7_, r_205__6_, r_205__5_, r_205__4_, r_205__3_, r_205__2_, r_205__1_, r_205__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N409)? data_i : 1'b0;
  assign N408 = sel_i[408];
  assign N409 = N1536;
  assign { r_n_205__31_, r_n_205__30_, r_n_205__29_, r_n_205__28_, r_n_205__27_, r_n_205__26_, r_n_205__25_, r_n_205__24_, r_n_205__23_, r_n_205__22_, r_n_205__21_, r_n_205__20_, r_n_205__19_, r_n_205__18_, r_n_205__17_, r_n_205__16_, r_n_205__15_, r_n_205__14_, r_n_205__13_, r_n_205__12_, r_n_205__11_, r_n_205__10_, r_n_205__9_, r_n_205__8_, r_n_205__7_, r_n_205__6_, r_n_205__5_, r_n_205__4_, r_n_205__3_, r_n_205__2_, r_n_205__1_, r_n_205__0_ } = (N410)? { r_206__31_, r_206__30_, r_206__29_, r_206__28_, r_206__27_, r_206__26_, r_206__25_, r_206__24_, r_206__23_, r_206__22_, r_206__21_, r_206__20_, r_206__19_, r_206__18_, r_206__17_, r_206__16_, r_206__15_, r_206__14_, r_206__13_, r_206__12_, r_206__11_, r_206__10_, r_206__9_, r_206__8_, r_206__7_, r_206__6_, r_206__5_, r_206__4_, r_206__3_, r_206__2_, r_206__1_, r_206__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N411)? data_i : 1'b0;
  assign N410 = sel_i[410];
  assign N411 = N1541;
  assign { r_n_206__31_, r_n_206__30_, r_n_206__29_, r_n_206__28_, r_n_206__27_, r_n_206__26_, r_n_206__25_, r_n_206__24_, r_n_206__23_, r_n_206__22_, r_n_206__21_, r_n_206__20_, r_n_206__19_, r_n_206__18_, r_n_206__17_, r_n_206__16_, r_n_206__15_, r_n_206__14_, r_n_206__13_, r_n_206__12_, r_n_206__11_, r_n_206__10_, r_n_206__9_, r_n_206__8_, r_n_206__7_, r_n_206__6_, r_n_206__5_, r_n_206__4_, r_n_206__3_, r_n_206__2_, r_n_206__1_, r_n_206__0_ } = (N412)? { r_207__31_, r_207__30_, r_207__29_, r_207__28_, r_207__27_, r_207__26_, r_207__25_, r_207__24_, r_207__23_, r_207__22_, r_207__21_, r_207__20_, r_207__19_, r_207__18_, r_207__17_, r_207__16_, r_207__15_, r_207__14_, r_207__13_, r_207__12_, r_207__11_, r_207__10_, r_207__9_, r_207__8_, r_207__7_, r_207__6_, r_207__5_, r_207__4_, r_207__3_, r_207__2_, r_207__1_, r_207__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N413)? data_i : 1'b0;
  assign N412 = sel_i[412];
  assign N413 = N1546;
  assign { r_n_207__31_, r_n_207__30_, r_n_207__29_, r_n_207__28_, r_n_207__27_, r_n_207__26_, r_n_207__25_, r_n_207__24_, r_n_207__23_, r_n_207__22_, r_n_207__21_, r_n_207__20_, r_n_207__19_, r_n_207__18_, r_n_207__17_, r_n_207__16_, r_n_207__15_, r_n_207__14_, r_n_207__13_, r_n_207__12_, r_n_207__11_, r_n_207__10_, r_n_207__9_, r_n_207__8_, r_n_207__7_, r_n_207__6_, r_n_207__5_, r_n_207__4_, r_n_207__3_, r_n_207__2_, r_n_207__1_, r_n_207__0_ } = (N414)? { r_208__31_, r_208__30_, r_208__29_, r_208__28_, r_208__27_, r_208__26_, r_208__25_, r_208__24_, r_208__23_, r_208__22_, r_208__21_, r_208__20_, r_208__19_, r_208__18_, r_208__17_, r_208__16_, r_208__15_, r_208__14_, r_208__13_, r_208__12_, r_208__11_, r_208__10_, r_208__9_, r_208__8_, r_208__7_, r_208__6_, r_208__5_, r_208__4_, r_208__3_, r_208__2_, r_208__1_, r_208__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N415)? data_i : 1'b0;
  assign N414 = sel_i[414];
  assign N415 = N1551;
  assign { r_n_208__31_, r_n_208__30_, r_n_208__29_, r_n_208__28_, r_n_208__27_, r_n_208__26_, r_n_208__25_, r_n_208__24_, r_n_208__23_, r_n_208__22_, r_n_208__21_, r_n_208__20_, r_n_208__19_, r_n_208__18_, r_n_208__17_, r_n_208__16_, r_n_208__15_, r_n_208__14_, r_n_208__13_, r_n_208__12_, r_n_208__11_, r_n_208__10_, r_n_208__9_, r_n_208__8_, r_n_208__7_, r_n_208__6_, r_n_208__5_, r_n_208__4_, r_n_208__3_, r_n_208__2_, r_n_208__1_, r_n_208__0_ } = (N416)? { r_209__31_, r_209__30_, r_209__29_, r_209__28_, r_209__27_, r_209__26_, r_209__25_, r_209__24_, r_209__23_, r_209__22_, r_209__21_, r_209__20_, r_209__19_, r_209__18_, r_209__17_, r_209__16_, r_209__15_, r_209__14_, r_209__13_, r_209__12_, r_209__11_, r_209__10_, r_209__9_, r_209__8_, r_209__7_, r_209__6_, r_209__5_, r_209__4_, r_209__3_, r_209__2_, r_209__1_, r_209__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N417)? data_i : 1'b0;
  assign N416 = sel_i[416];
  assign N417 = N1556;
  assign { r_n_209__31_, r_n_209__30_, r_n_209__29_, r_n_209__28_, r_n_209__27_, r_n_209__26_, r_n_209__25_, r_n_209__24_, r_n_209__23_, r_n_209__22_, r_n_209__21_, r_n_209__20_, r_n_209__19_, r_n_209__18_, r_n_209__17_, r_n_209__16_, r_n_209__15_, r_n_209__14_, r_n_209__13_, r_n_209__12_, r_n_209__11_, r_n_209__10_, r_n_209__9_, r_n_209__8_, r_n_209__7_, r_n_209__6_, r_n_209__5_, r_n_209__4_, r_n_209__3_, r_n_209__2_, r_n_209__1_, r_n_209__0_ } = (N418)? { r_210__31_, r_210__30_, r_210__29_, r_210__28_, r_210__27_, r_210__26_, r_210__25_, r_210__24_, r_210__23_, r_210__22_, r_210__21_, r_210__20_, r_210__19_, r_210__18_, r_210__17_, r_210__16_, r_210__15_, r_210__14_, r_210__13_, r_210__12_, r_210__11_, r_210__10_, r_210__9_, r_210__8_, r_210__7_, r_210__6_, r_210__5_, r_210__4_, r_210__3_, r_210__2_, r_210__1_, r_210__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N419)? data_i : 1'b0;
  assign N418 = sel_i[418];
  assign N419 = N1561;
  assign { r_n_210__31_, r_n_210__30_, r_n_210__29_, r_n_210__28_, r_n_210__27_, r_n_210__26_, r_n_210__25_, r_n_210__24_, r_n_210__23_, r_n_210__22_, r_n_210__21_, r_n_210__20_, r_n_210__19_, r_n_210__18_, r_n_210__17_, r_n_210__16_, r_n_210__15_, r_n_210__14_, r_n_210__13_, r_n_210__12_, r_n_210__11_, r_n_210__10_, r_n_210__9_, r_n_210__8_, r_n_210__7_, r_n_210__6_, r_n_210__5_, r_n_210__4_, r_n_210__3_, r_n_210__2_, r_n_210__1_, r_n_210__0_ } = (N420)? { r_211__31_, r_211__30_, r_211__29_, r_211__28_, r_211__27_, r_211__26_, r_211__25_, r_211__24_, r_211__23_, r_211__22_, r_211__21_, r_211__20_, r_211__19_, r_211__18_, r_211__17_, r_211__16_, r_211__15_, r_211__14_, r_211__13_, r_211__12_, r_211__11_, r_211__10_, r_211__9_, r_211__8_, r_211__7_, r_211__6_, r_211__5_, r_211__4_, r_211__3_, r_211__2_, r_211__1_, r_211__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N421)? data_i : 1'b0;
  assign N420 = sel_i[420];
  assign N421 = N1566;
  assign { r_n_211__31_, r_n_211__30_, r_n_211__29_, r_n_211__28_, r_n_211__27_, r_n_211__26_, r_n_211__25_, r_n_211__24_, r_n_211__23_, r_n_211__22_, r_n_211__21_, r_n_211__20_, r_n_211__19_, r_n_211__18_, r_n_211__17_, r_n_211__16_, r_n_211__15_, r_n_211__14_, r_n_211__13_, r_n_211__12_, r_n_211__11_, r_n_211__10_, r_n_211__9_, r_n_211__8_, r_n_211__7_, r_n_211__6_, r_n_211__5_, r_n_211__4_, r_n_211__3_, r_n_211__2_, r_n_211__1_, r_n_211__0_ } = (N422)? { r_212__31_, r_212__30_, r_212__29_, r_212__28_, r_212__27_, r_212__26_, r_212__25_, r_212__24_, r_212__23_, r_212__22_, r_212__21_, r_212__20_, r_212__19_, r_212__18_, r_212__17_, r_212__16_, r_212__15_, r_212__14_, r_212__13_, r_212__12_, r_212__11_, r_212__10_, r_212__9_, r_212__8_, r_212__7_, r_212__6_, r_212__5_, r_212__4_, r_212__3_, r_212__2_, r_212__1_, r_212__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N423)? data_i : 1'b0;
  assign N422 = sel_i[422];
  assign N423 = N1571;
  assign { r_n_212__31_, r_n_212__30_, r_n_212__29_, r_n_212__28_, r_n_212__27_, r_n_212__26_, r_n_212__25_, r_n_212__24_, r_n_212__23_, r_n_212__22_, r_n_212__21_, r_n_212__20_, r_n_212__19_, r_n_212__18_, r_n_212__17_, r_n_212__16_, r_n_212__15_, r_n_212__14_, r_n_212__13_, r_n_212__12_, r_n_212__11_, r_n_212__10_, r_n_212__9_, r_n_212__8_, r_n_212__7_, r_n_212__6_, r_n_212__5_, r_n_212__4_, r_n_212__3_, r_n_212__2_, r_n_212__1_, r_n_212__0_ } = (N424)? { r_213__31_, r_213__30_, r_213__29_, r_213__28_, r_213__27_, r_213__26_, r_213__25_, r_213__24_, r_213__23_, r_213__22_, r_213__21_, r_213__20_, r_213__19_, r_213__18_, r_213__17_, r_213__16_, r_213__15_, r_213__14_, r_213__13_, r_213__12_, r_213__11_, r_213__10_, r_213__9_, r_213__8_, r_213__7_, r_213__6_, r_213__5_, r_213__4_, r_213__3_, r_213__2_, r_213__1_, r_213__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N425)? data_i : 1'b0;
  assign N424 = sel_i[424];
  assign N425 = N1576;
  assign { r_n_213__31_, r_n_213__30_, r_n_213__29_, r_n_213__28_, r_n_213__27_, r_n_213__26_, r_n_213__25_, r_n_213__24_, r_n_213__23_, r_n_213__22_, r_n_213__21_, r_n_213__20_, r_n_213__19_, r_n_213__18_, r_n_213__17_, r_n_213__16_, r_n_213__15_, r_n_213__14_, r_n_213__13_, r_n_213__12_, r_n_213__11_, r_n_213__10_, r_n_213__9_, r_n_213__8_, r_n_213__7_, r_n_213__6_, r_n_213__5_, r_n_213__4_, r_n_213__3_, r_n_213__2_, r_n_213__1_, r_n_213__0_ } = (N426)? { r_214__31_, r_214__30_, r_214__29_, r_214__28_, r_214__27_, r_214__26_, r_214__25_, r_214__24_, r_214__23_, r_214__22_, r_214__21_, r_214__20_, r_214__19_, r_214__18_, r_214__17_, r_214__16_, r_214__15_, r_214__14_, r_214__13_, r_214__12_, r_214__11_, r_214__10_, r_214__9_, r_214__8_, r_214__7_, r_214__6_, r_214__5_, r_214__4_, r_214__3_, r_214__2_, r_214__1_, r_214__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N427)? data_i : 1'b0;
  assign N426 = sel_i[426];
  assign N427 = N1581;
  assign { r_n_214__31_, r_n_214__30_, r_n_214__29_, r_n_214__28_, r_n_214__27_, r_n_214__26_, r_n_214__25_, r_n_214__24_, r_n_214__23_, r_n_214__22_, r_n_214__21_, r_n_214__20_, r_n_214__19_, r_n_214__18_, r_n_214__17_, r_n_214__16_, r_n_214__15_, r_n_214__14_, r_n_214__13_, r_n_214__12_, r_n_214__11_, r_n_214__10_, r_n_214__9_, r_n_214__8_, r_n_214__7_, r_n_214__6_, r_n_214__5_, r_n_214__4_, r_n_214__3_, r_n_214__2_, r_n_214__1_, r_n_214__0_ } = (N428)? { r_215__31_, r_215__30_, r_215__29_, r_215__28_, r_215__27_, r_215__26_, r_215__25_, r_215__24_, r_215__23_, r_215__22_, r_215__21_, r_215__20_, r_215__19_, r_215__18_, r_215__17_, r_215__16_, r_215__15_, r_215__14_, r_215__13_, r_215__12_, r_215__11_, r_215__10_, r_215__9_, r_215__8_, r_215__7_, r_215__6_, r_215__5_, r_215__4_, r_215__3_, r_215__2_, r_215__1_, r_215__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N429)? data_i : 1'b0;
  assign N428 = sel_i[428];
  assign N429 = N1586;
  assign { r_n_215__31_, r_n_215__30_, r_n_215__29_, r_n_215__28_, r_n_215__27_, r_n_215__26_, r_n_215__25_, r_n_215__24_, r_n_215__23_, r_n_215__22_, r_n_215__21_, r_n_215__20_, r_n_215__19_, r_n_215__18_, r_n_215__17_, r_n_215__16_, r_n_215__15_, r_n_215__14_, r_n_215__13_, r_n_215__12_, r_n_215__11_, r_n_215__10_, r_n_215__9_, r_n_215__8_, r_n_215__7_, r_n_215__6_, r_n_215__5_, r_n_215__4_, r_n_215__3_, r_n_215__2_, r_n_215__1_, r_n_215__0_ } = (N430)? { r_216__31_, r_216__30_, r_216__29_, r_216__28_, r_216__27_, r_216__26_, r_216__25_, r_216__24_, r_216__23_, r_216__22_, r_216__21_, r_216__20_, r_216__19_, r_216__18_, r_216__17_, r_216__16_, r_216__15_, r_216__14_, r_216__13_, r_216__12_, r_216__11_, r_216__10_, r_216__9_, r_216__8_, r_216__7_, r_216__6_, r_216__5_, r_216__4_, r_216__3_, r_216__2_, r_216__1_, r_216__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N431)? data_i : 1'b0;
  assign N430 = sel_i[430];
  assign N431 = N1591;
  assign { r_n_216__31_, r_n_216__30_, r_n_216__29_, r_n_216__28_, r_n_216__27_, r_n_216__26_, r_n_216__25_, r_n_216__24_, r_n_216__23_, r_n_216__22_, r_n_216__21_, r_n_216__20_, r_n_216__19_, r_n_216__18_, r_n_216__17_, r_n_216__16_, r_n_216__15_, r_n_216__14_, r_n_216__13_, r_n_216__12_, r_n_216__11_, r_n_216__10_, r_n_216__9_, r_n_216__8_, r_n_216__7_, r_n_216__6_, r_n_216__5_, r_n_216__4_, r_n_216__3_, r_n_216__2_, r_n_216__1_, r_n_216__0_ } = (N432)? { r_217__31_, r_217__30_, r_217__29_, r_217__28_, r_217__27_, r_217__26_, r_217__25_, r_217__24_, r_217__23_, r_217__22_, r_217__21_, r_217__20_, r_217__19_, r_217__18_, r_217__17_, r_217__16_, r_217__15_, r_217__14_, r_217__13_, r_217__12_, r_217__11_, r_217__10_, r_217__9_, r_217__8_, r_217__7_, r_217__6_, r_217__5_, r_217__4_, r_217__3_, r_217__2_, r_217__1_, r_217__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N433)? data_i : 1'b0;
  assign N432 = sel_i[432];
  assign N433 = N1596;
  assign { r_n_217__31_, r_n_217__30_, r_n_217__29_, r_n_217__28_, r_n_217__27_, r_n_217__26_, r_n_217__25_, r_n_217__24_, r_n_217__23_, r_n_217__22_, r_n_217__21_, r_n_217__20_, r_n_217__19_, r_n_217__18_, r_n_217__17_, r_n_217__16_, r_n_217__15_, r_n_217__14_, r_n_217__13_, r_n_217__12_, r_n_217__11_, r_n_217__10_, r_n_217__9_, r_n_217__8_, r_n_217__7_, r_n_217__6_, r_n_217__5_, r_n_217__4_, r_n_217__3_, r_n_217__2_, r_n_217__1_, r_n_217__0_ } = (N434)? { r_218__31_, r_218__30_, r_218__29_, r_218__28_, r_218__27_, r_218__26_, r_218__25_, r_218__24_, r_218__23_, r_218__22_, r_218__21_, r_218__20_, r_218__19_, r_218__18_, r_218__17_, r_218__16_, r_218__15_, r_218__14_, r_218__13_, r_218__12_, r_218__11_, r_218__10_, r_218__9_, r_218__8_, r_218__7_, r_218__6_, r_218__5_, r_218__4_, r_218__3_, r_218__2_, r_218__1_, r_218__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N435)? data_i : 1'b0;
  assign N434 = sel_i[434];
  assign N435 = N1601;
  assign { r_n_218__31_, r_n_218__30_, r_n_218__29_, r_n_218__28_, r_n_218__27_, r_n_218__26_, r_n_218__25_, r_n_218__24_, r_n_218__23_, r_n_218__22_, r_n_218__21_, r_n_218__20_, r_n_218__19_, r_n_218__18_, r_n_218__17_, r_n_218__16_, r_n_218__15_, r_n_218__14_, r_n_218__13_, r_n_218__12_, r_n_218__11_, r_n_218__10_, r_n_218__9_, r_n_218__8_, r_n_218__7_, r_n_218__6_, r_n_218__5_, r_n_218__4_, r_n_218__3_, r_n_218__2_, r_n_218__1_, r_n_218__0_ } = (N436)? { r_219__31_, r_219__30_, r_219__29_, r_219__28_, r_219__27_, r_219__26_, r_219__25_, r_219__24_, r_219__23_, r_219__22_, r_219__21_, r_219__20_, r_219__19_, r_219__18_, r_219__17_, r_219__16_, r_219__15_, r_219__14_, r_219__13_, r_219__12_, r_219__11_, r_219__10_, r_219__9_, r_219__8_, r_219__7_, r_219__6_, r_219__5_, r_219__4_, r_219__3_, r_219__2_, r_219__1_, r_219__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N437)? data_i : 1'b0;
  assign N436 = sel_i[436];
  assign N437 = N1606;
  assign { r_n_219__31_, r_n_219__30_, r_n_219__29_, r_n_219__28_, r_n_219__27_, r_n_219__26_, r_n_219__25_, r_n_219__24_, r_n_219__23_, r_n_219__22_, r_n_219__21_, r_n_219__20_, r_n_219__19_, r_n_219__18_, r_n_219__17_, r_n_219__16_, r_n_219__15_, r_n_219__14_, r_n_219__13_, r_n_219__12_, r_n_219__11_, r_n_219__10_, r_n_219__9_, r_n_219__8_, r_n_219__7_, r_n_219__6_, r_n_219__5_, r_n_219__4_, r_n_219__3_, r_n_219__2_, r_n_219__1_, r_n_219__0_ } = (N438)? { r_220__31_, r_220__30_, r_220__29_, r_220__28_, r_220__27_, r_220__26_, r_220__25_, r_220__24_, r_220__23_, r_220__22_, r_220__21_, r_220__20_, r_220__19_, r_220__18_, r_220__17_, r_220__16_, r_220__15_, r_220__14_, r_220__13_, r_220__12_, r_220__11_, r_220__10_, r_220__9_, r_220__8_, r_220__7_, r_220__6_, r_220__5_, r_220__4_, r_220__3_, r_220__2_, r_220__1_, r_220__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N439)? data_i : 1'b0;
  assign N438 = sel_i[438];
  assign N439 = N1611;
  assign { r_n_220__31_, r_n_220__30_, r_n_220__29_, r_n_220__28_, r_n_220__27_, r_n_220__26_, r_n_220__25_, r_n_220__24_, r_n_220__23_, r_n_220__22_, r_n_220__21_, r_n_220__20_, r_n_220__19_, r_n_220__18_, r_n_220__17_, r_n_220__16_, r_n_220__15_, r_n_220__14_, r_n_220__13_, r_n_220__12_, r_n_220__11_, r_n_220__10_, r_n_220__9_, r_n_220__8_, r_n_220__7_, r_n_220__6_, r_n_220__5_, r_n_220__4_, r_n_220__3_, r_n_220__2_, r_n_220__1_, r_n_220__0_ } = (N440)? { r_221__31_, r_221__30_, r_221__29_, r_221__28_, r_221__27_, r_221__26_, r_221__25_, r_221__24_, r_221__23_, r_221__22_, r_221__21_, r_221__20_, r_221__19_, r_221__18_, r_221__17_, r_221__16_, r_221__15_, r_221__14_, r_221__13_, r_221__12_, r_221__11_, r_221__10_, r_221__9_, r_221__8_, r_221__7_, r_221__6_, r_221__5_, r_221__4_, r_221__3_, r_221__2_, r_221__1_, r_221__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N441)? data_i : 1'b0;
  assign N440 = sel_i[440];
  assign N441 = N1616;
  assign { r_n_221__31_, r_n_221__30_, r_n_221__29_, r_n_221__28_, r_n_221__27_, r_n_221__26_, r_n_221__25_, r_n_221__24_, r_n_221__23_, r_n_221__22_, r_n_221__21_, r_n_221__20_, r_n_221__19_, r_n_221__18_, r_n_221__17_, r_n_221__16_, r_n_221__15_, r_n_221__14_, r_n_221__13_, r_n_221__12_, r_n_221__11_, r_n_221__10_, r_n_221__9_, r_n_221__8_, r_n_221__7_, r_n_221__6_, r_n_221__5_, r_n_221__4_, r_n_221__3_, r_n_221__2_, r_n_221__1_, r_n_221__0_ } = (N442)? { r_222__31_, r_222__30_, r_222__29_, r_222__28_, r_222__27_, r_222__26_, r_222__25_, r_222__24_, r_222__23_, r_222__22_, r_222__21_, r_222__20_, r_222__19_, r_222__18_, r_222__17_, r_222__16_, r_222__15_, r_222__14_, r_222__13_, r_222__12_, r_222__11_, r_222__10_, r_222__9_, r_222__8_, r_222__7_, r_222__6_, r_222__5_, r_222__4_, r_222__3_, r_222__2_, r_222__1_, r_222__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N443)? data_i : 1'b0;
  assign N442 = sel_i[442];
  assign N443 = N1621;
  assign { r_n_222__31_, r_n_222__30_, r_n_222__29_, r_n_222__28_, r_n_222__27_, r_n_222__26_, r_n_222__25_, r_n_222__24_, r_n_222__23_, r_n_222__22_, r_n_222__21_, r_n_222__20_, r_n_222__19_, r_n_222__18_, r_n_222__17_, r_n_222__16_, r_n_222__15_, r_n_222__14_, r_n_222__13_, r_n_222__12_, r_n_222__11_, r_n_222__10_, r_n_222__9_, r_n_222__8_, r_n_222__7_, r_n_222__6_, r_n_222__5_, r_n_222__4_, r_n_222__3_, r_n_222__2_, r_n_222__1_, r_n_222__0_ } = (N444)? { r_223__31_, r_223__30_, r_223__29_, r_223__28_, r_223__27_, r_223__26_, r_223__25_, r_223__24_, r_223__23_, r_223__22_, r_223__21_, r_223__20_, r_223__19_, r_223__18_, r_223__17_, r_223__16_, r_223__15_, r_223__14_, r_223__13_, r_223__12_, r_223__11_, r_223__10_, r_223__9_, r_223__8_, r_223__7_, r_223__6_, r_223__5_, r_223__4_, r_223__3_, r_223__2_, r_223__1_, r_223__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N445)? data_i : 1'b0;
  assign N444 = sel_i[444];
  assign N445 = N1626;
  assign { r_n_223__31_, r_n_223__30_, r_n_223__29_, r_n_223__28_, r_n_223__27_, r_n_223__26_, r_n_223__25_, r_n_223__24_, r_n_223__23_, r_n_223__22_, r_n_223__21_, r_n_223__20_, r_n_223__19_, r_n_223__18_, r_n_223__17_, r_n_223__16_, r_n_223__15_, r_n_223__14_, r_n_223__13_, r_n_223__12_, r_n_223__11_, r_n_223__10_, r_n_223__9_, r_n_223__8_, r_n_223__7_, r_n_223__6_, r_n_223__5_, r_n_223__4_, r_n_223__3_, r_n_223__2_, r_n_223__1_, r_n_223__0_ } = (N446)? { r_224__31_, r_224__30_, r_224__29_, r_224__28_, r_224__27_, r_224__26_, r_224__25_, r_224__24_, r_224__23_, r_224__22_, r_224__21_, r_224__20_, r_224__19_, r_224__18_, r_224__17_, r_224__16_, r_224__15_, r_224__14_, r_224__13_, r_224__12_, r_224__11_, r_224__10_, r_224__9_, r_224__8_, r_224__7_, r_224__6_, r_224__5_, r_224__4_, r_224__3_, r_224__2_, r_224__1_, r_224__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N447)? data_i : 1'b0;
  assign N446 = sel_i[446];
  assign N447 = N1631;
  assign { r_n_224__31_, r_n_224__30_, r_n_224__29_, r_n_224__28_, r_n_224__27_, r_n_224__26_, r_n_224__25_, r_n_224__24_, r_n_224__23_, r_n_224__22_, r_n_224__21_, r_n_224__20_, r_n_224__19_, r_n_224__18_, r_n_224__17_, r_n_224__16_, r_n_224__15_, r_n_224__14_, r_n_224__13_, r_n_224__12_, r_n_224__11_, r_n_224__10_, r_n_224__9_, r_n_224__8_, r_n_224__7_, r_n_224__6_, r_n_224__5_, r_n_224__4_, r_n_224__3_, r_n_224__2_, r_n_224__1_, r_n_224__0_ } = (N448)? { r_225__31_, r_225__30_, r_225__29_, r_225__28_, r_225__27_, r_225__26_, r_225__25_, r_225__24_, r_225__23_, r_225__22_, r_225__21_, r_225__20_, r_225__19_, r_225__18_, r_225__17_, r_225__16_, r_225__15_, r_225__14_, r_225__13_, r_225__12_, r_225__11_, r_225__10_, r_225__9_, r_225__8_, r_225__7_, r_225__6_, r_225__5_, r_225__4_, r_225__3_, r_225__2_, r_225__1_, r_225__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N449)? data_i : 1'b0;
  assign N448 = sel_i[448];
  assign N449 = N1636;
  assign { r_n_225__31_, r_n_225__30_, r_n_225__29_, r_n_225__28_, r_n_225__27_, r_n_225__26_, r_n_225__25_, r_n_225__24_, r_n_225__23_, r_n_225__22_, r_n_225__21_, r_n_225__20_, r_n_225__19_, r_n_225__18_, r_n_225__17_, r_n_225__16_, r_n_225__15_, r_n_225__14_, r_n_225__13_, r_n_225__12_, r_n_225__11_, r_n_225__10_, r_n_225__9_, r_n_225__8_, r_n_225__7_, r_n_225__6_, r_n_225__5_, r_n_225__4_, r_n_225__3_, r_n_225__2_, r_n_225__1_, r_n_225__0_ } = (N450)? { r_226__31_, r_226__30_, r_226__29_, r_226__28_, r_226__27_, r_226__26_, r_226__25_, r_226__24_, r_226__23_, r_226__22_, r_226__21_, r_226__20_, r_226__19_, r_226__18_, r_226__17_, r_226__16_, r_226__15_, r_226__14_, r_226__13_, r_226__12_, r_226__11_, r_226__10_, r_226__9_, r_226__8_, r_226__7_, r_226__6_, r_226__5_, r_226__4_, r_226__3_, r_226__2_, r_226__1_, r_226__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N451)? data_i : 1'b0;
  assign N450 = sel_i[450];
  assign N451 = N1641;
  assign { r_n_226__31_, r_n_226__30_, r_n_226__29_, r_n_226__28_, r_n_226__27_, r_n_226__26_, r_n_226__25_, r_n_226__24_, r_n_226__23_, r_n_226__22_, r_n_226__21_, r_n_226__20_, r_n_226__19_, r_n_226__18_, r_n_226__17_, r_n_226__16_, r_n_226__15_, r_n_226__14_, r_n_226__13_, r_n_226__12_, r_n_226__11_, r_n_226__10_, r_n_226__9_, r_n_226__8_, r_n_226__7_, r_n_226__6_, r_n_226__5_, r_n_226__4_, r_n_226__3_, r_n_226__2_, r_n_226__1_, r_n_226__0_ } = (N452)? { r_227__31_, r_227__30_, r_227__29_, r_227__28_, r_227__27_, r_227__26_, r_227__25_, r_227__24_, r_227__23_, r_227__22_, r_227__21_, r_227__20_, r_227__19_, r_227__18_, r_227__17_, r_227__16_, r_227__15_, r_227__14_, r_227__13_, r_227__12_, r_227__11_, r_227__10_, r_227__9_, r_227__8_, r_227__7_, r_227__6_, r_227__5_, r_227__4_, r_227__3_, r_227__2_, r_227__1_, r_227__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N453)? data_i : 1'b0;
  assign N452 = sel_i[452];
  assign N453 = N1646;
  assign { r_n_227__31_, r_n_227__30_, r_n_227__29_, r_n_227__28_, r_n_227__27_, r_n_227__26_, r_n_227__25_, r_n_227__24_, r_n_227__23_, r_n_227__22_, r_n_227__21_, r_n_227__20_, r_n_227__19_, r_n_227__18_, r_n_227__17_, r_n_227__16_, r_n_227__15_, r_n_227__14_, r_n_227__13_, r_n_227__12_, r_n_227__11_, r_n_227__10_, r_n_227__9_, r_n_227__8_, r_n_227__7_, r_n_227__6_, r_n_227__5_, r_n_227__4_, r_n_227__3_, r_n_227__2_, r_n_227__1_, r_n_227__0_ } = (N454)? { r_228__31_, r_228__30_, r_228__29_, r_228__28_, r_228__27_, r_228__26_, r_228__25_, r_228__24_, r_228__23_, r_228__22_, r_228__21_, r_228__20_, r_228__19_, r_228__18_, r_228__17_, r_228__16_, r_228__15_, r_228__14_, r_228__13_, r_228__12_, r_228__11_, r_228__10_, r_228__9_, r_228__8_, r_228__7_, r_228__6_, r_228__5_, r_228__4_, r_228__3_, r_228__2_, r_228__1_, r_228__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N455)? data_i : 1'b0;
  assign N454 = sel_i[454];
  assign N455 = N1651;
  assign { r_n_228__31_, r_n_228__30_, r_n_228__29_, r_n_228__28_, r_n_228__27_, r_n_228__26_, r_n_228__25_, r_n_228__24_, r_n_228__23_, r_n_228__22_, r_n_228__21_, r_n_228__20_, r_n_228__19_, r_n_228__18_, r_n_228__17_, r_n_228__16_, r_n_228__15_, r_n_228__14_, r_n_228__13_, r_n_228__12_, r_n_228__11_, r_n_228__10_, r_n_228__9_, r_n_228__8_, r_n_228__7_, r_n_228__6_, r_n_228__5_, r_n_228__4_, r_n_228__3_, r_n_228__2_, r_n_228__1_, r_n_228__0_ } = (N456)? { r_229__31_, r_229__30_, r_229__29_, r_229__28_, r_229__27_, r_229__26_, r_229__25_, r_229__24_, r_229__23_, r_229__22_, r_229__21_, r_229__20_, r_229__19_, r_229__18_, r_229__17_, r_229__16_, r_229__15_, r_229__14_, r_229__13_, r_229__12_, r_229__11_, r_229__10_, r_229__9_, r_229__8_, r_229__7_, r_229__6_, r_229__5_, r_229__4_, r_229__3_, r_229__2_, r_229__1_, r_229__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N457)? data_i : 1'b0;
  assign N456 = sel_i[456];
  assign N457 = N1656;
  assign { r_n_229__31_, r_n_229__30_, r_n_229__29_, r_n_229__28_, r_n_229__27_, r_n_229__26_, r_n_229__25_, r_n_229__24_, r_n_229__23_, r_n_229__22_, r_n_229__21_, r_n_229__20_, r_n_229__19_, r_n_229__18_, r_n_229__17_, r_n_229__16_, r_n_229__15_, r_n_229__14_, r_n_229__13_, r_n_229__12_, r_n_229__11_, r_n_229__10_, r_n_229__9_, r_n_229__8_, r_n_229__7_, r_n_229__6_, r_n_229__5_, r_n_229__4_, r_n_229__3_, r_n_229__2_, r_n_229__1_, r_n_229__0_ } = (N458)? { r_230__31_, r_230__30_, r_230__29_, r_230__28_, r_230__27_, r_230__26_, r_230__25_, r_230__24_, r_230__23_, r_230__22_, r_230__21_, r_230__20_, r_230__19_, r_230__18_, r_230__17_, r_230__16_, r_230__15_, r_230__14_, r_230__13_, r_230__12_, r_230__11_, r_230__10_, r_230__9_, r_230__8_, r_230__7_, r_230__6_, r_230__5_, r_230__4_, r_230__3_, r_230__2_, r_230__1_, r_230__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N459)? data_i : 1'b0;
  assign N458 = sel_i[458];
  assign N459 = N1661;
  assign { r_n_230__31_, r_n_230__30_, r_n_230__29_, r_n_230__28_, r_n_230__27_, r_n_230__26_, r_n_230__25_, r_n_230__24_, r_n_230__23_, r_n_230__22_, r_n_230__21_, r_n_230__20_, r_n_230__19_, r_n_230__18_, r_n_230__17_, r_n_230__16_, r_n_230__15_, r_n_230__14_, r_n_230__13_, r_n_230__12_, r_n_230__11_, r_n_230__10_, r_n_230__9_, r_n_230__8_, r_n_230__7_, r_n_230__6_, r_n_230__5_, r_n_230__4_, r_n_230__3_, r_n_230__2_, r_n_230__1_, r_n_230__0_ } = (N460)? { r_231__31_, r_231__30_, r_231__29_, r_231__28_, r_231__27_, r_231__26_, r_231__25_, r_231__24_, r_231__23_, r_231__22_, r_231__21_, r_231__20_, r_231__19_, r_231__18_, r_231__17_, r_231__16_, r_231__15_, r_231__14_, r_231__13_, r_231__12_, r_231__11_, r_231__10_, r_231__9_, r_231__8_, r_231__7_, r_231__6_, r_231__5_, r_231__4_, r_231__3_, r_231__2_, r_231__1_, r_231__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N461)? data_i : 1'b0;
  assign N460 = sel_i[460];
  assign N461 = N1666;
  assign { r_n_231__31_, r_n_231__30_, r_n_231__29_, r_n_231__28_, r_n_231__27_, r_n_231__26_, r_n_231__25_, r_n_231__24_, r_n_231__23_, r_n_231__22_, r_n_231__21_, r_n_231__20_, r_n_231__19_, r_n_231__18_, r_n_231__17_, r_n_231__16_, r_n_231__15_, r_n_231__14_, r_n_231__13_, r_n_231__12_, r_n_231__11_, r_n_231__10_, r_n_231__9_, r_n_231__8_, r_n_231__7_, r_n_231__6_, r_n_231__5_, r_n_231__4_, r_n_231__3_, r_n_231__2_, r_n_231__1_, r_n_231__0_ } = (N462)? { r_232__31_, r_232__30_, r_232__29_, r_232__28_, r_232__27_, r_232__26_, r_232__25_, r_232__24_, r_232__23_, r_232__22_, r_232__21_, r_232__20_, r_232__19_, r_232__18_, r_232__17_, r_232__16_, r_232__15_, r_232__14_, r_232__13_, r_232__12_, r_232__11_, r_232__10_, r_232__9_, r_232__8_, r_232__7_, r_232__6_, r_232__5_, r_232__4_, r_232__3_, r_232__2_, r_232__1_, r_232__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N463)? data_i : 1'b0;
  assign N462 = sel_i[462];
  assign N463 = N1671;
  assign { r_n_232__31_, r_n_232__30_, r_n_232__29_, r_n_232__28_, r_n_232__27_, r_n_232__26_, r_n_232__25_, r_n_232__24_, r_n_232__23_, r_n_232__22_, r_n_232__21_, r_n_232__20_, r_n_232__19_, r_n_232__18_, r_n_232__17_, r_n_232__16_, r_n_232__15_, r_n_232__14_, r_n_232__13_, r_n_232__12_, r_n_232__11_, r_n_232__10_, r_n_232__9_, r_n_232__8_, r_n_232__7_, r_n_232__6_, r_n_232__5_, r_n_232__4_, r_n_232__3_, r_n_232__2_, r_n_232__1_, r_n_232__0_ } = (N464)? { r_233__31_, r_233__30_, r_233__29_, r_233__28_, r_233__27_, r_233__26_, r_233__25_, r_233__24_, r_233__23_, r_233__22_, r_233__21_, r_233__20_, r_233__19_, r_233__18_, r_233__17_, r_233__16_, r_233__15_, r_233__14_, r_233__13_, r_233__12_, r_233__11_, r_233__10_, r_233__9_, r_233__8_, r_233__7_, r_233__6_, r_233__5_, r_233__4_, r_233__3_, r_233__2_, r_233__1_, r_233__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N465)? data_i : 1'b0;
  assign N464 = sel_i[464];
  assign N465 = N1676;
  assign { r_n_233__31_, r_n_233__30_, r_n_233__29_, r_n_233__28_, r_n_233__27_, r_n_233__26_, r_n_233__25_, r_n_233__24_, r_n_233__23_, r_n_233__22_, r_n_233__21_, r_n_233__20_, r_n_233__19_, r_n_233__18_, r_n_233__17_, r_n_233__16_, r_n_233__15_, r_n_233__14_, r_n_233__13_, r_n_233__12_, r_n_233__11_, r_n_233__10_, r_n_233__9_, r_n_233__8_, r_n_233__7_, r_n_233__6_, r_n_233__5_, r_n_233__4_, r_n_233__3_, r_n_233__2_, r_n_233__1_, r_n_233__0_ } = (N466)? { r_234__31_, r_234__30_, r_234__29_, r_234__28_, r_234__27_, r_234__26_, r_234__25_, r_234__24_, r_234__23_, r_234__22_, r_234__21_, r_234__20_, r_234__19_, r_234__18_, r_234__17_, r_234__16_, r_234__15_, r_234__14_, r_234__13_, r_234__12_, r_234__11_, r_234__10_, r_234__9_, r_234__8_, r_234__7_, r_234__6_, r_234__5_, r_234__4_, r_234__3_, r_234__2_, r_234__1_, r_234__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N467)? data_i : 1'b0;
  assign N466 = sel_i[466];
  assign N467 = N1681;
  assign { r_n_234__31_, r_n_234__30_, r_n_234__29_, r_n_234__28_, r_n_234__27_, r_n_234__26_, r_n_234__25_, r_n_234__24_, r_n_234__23_, r_n_234__22_, r_n_234__21_, r_n_234__20_, r_n_234__19_, r_n_234__18_, r_n_234__17_, r_n_234__16_, r_n_234__15_, r_n_234__14_, r_n_234__13_, r_n_234__12_, r_n_234__11_, r_n_234__10_, r_n_234__9_, r_n_234__8_, r_n_234__7_, r_n_234__6_, r_n_234__5_, r_n_234__4_, r_n_234__3_, r_n_234__2_, r_n_234__1_, r_n_234__0_ } = (N468)? { r_235__31_, r_235__30_, r_235__29_, r_235__28_, r_235__27_, r_235__26_, r_235__25_, r_235__24_, r_235__23_, r_235__22_, r_235__21_, r_235__20_, r_235__19_, r_235__18_, r_235__17_, r_235__16_, r_235__15_, r_235__14_, r_235__13_, r_235__12_, r_235__11_, r_235__10_, r_235__9_, r_235__8_, r_235__7_, r_235__6_, r_235__5_, r_235__4_, r_235__3_, r_235__2_, r_235__1_, r_235__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N469)? data_i : 1'b0;
  assign N468 = sel_i[468];
  assign N469 = N1686;
  assign { r_n_235__31_, r_n_235__30_, r_n_235__29_, r_n_235__28_, r_n_235__27_, r_n_235__26_, r_n_235__25_, r_n_235__24_, r_n_235__23_, r_n_235__22_, r_n_235__21_, r_n_235__20_, r_n_235__19_, r_n_235__18_, r_n_235__17_, r_n_235__16_, r_n_235__15_, r_n_235__14_, r_n_235__13_, r_n_235__12_, r_n_235__11_, r_n_235__10_, r_n_235__9_, r_n_235__8_, r_n_235__7_, r_n_235__6_, r_n_235__5_, r_n_235__4_, r_n_235__3_, r_n_235__2_, r_n_235__1_, r_n_235__0_ } = (N470)? { r_236__31_, r_236__30_, r_236__29_, r_236__28_, r_236__27_, r_236__26_, r_236__25_, r_236__24_, r_236__23_, r_236__22_, r_236__21_, r_236__20_, r_236__19_, r_236__18_, r_236__17_, r_236__16_, r_236__15_, r_236__14_, r_236__13_, r_236__12_, r_236__11_, r_236__10_, r_236__9_, r_236__8_, r_236__7_, r_236__6_, r_236__5_, r_236__4_, r_236__3_, r_236__2_, r_236__1_, r_236__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N471)? data_i : 1'b0;
  assign N470 = sel_i[470];
  assign N471 = N1691;
  assign { r_n_236__31_, r_n_236__30_, r_n_236__29_, r_n_236__28_, r_n_236__27_, r_n_236__26_, r_n_236__25_, r_n_236__24_, r_n_236__23_, r_n_236__22_, r_n_236__21_, r_n_236__20_, r_n_236__19_, r_n_236__18_, r_n_236__17_, r_n_236__16_, r_n_236__15_, r_n_236__14_, r_n_236__13_, r_n_236__12_, r_n_236__11_, r_n_236__10_, r_n_236__9_, r_n_236__8_, r_n_236__7_, r_n_236__6_, r_n_236__5_, r_n_236__4_, r_n_236__3_, r_n_236__2_, r_n_236__1_, r_n_236__0_ } = (N472)? { r_237__31_, r_237__30_, r_237__29_, r_237__28_, r_237__27_, r_237__26_, r_237__25_, r_237__24_, r_237__23_, r_237__22_, r_237__21_, r_237__20_, r_237__19_, r_237__18_, r_237__17_, r_237__16_, r_237__15_, r_237__14_, r_237__13_, r_237__12_, r_237__11_, r_237__10_, r_237__9_, r_237__8_, r_237__7_, r_237__6_, r_237__5_, r_237__4_, r_237__3_, r_237__2_, r_237__1_, r_237__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N473)? data_i : 1'b0;
  assign N472 = sel_i[472];
  assign N473 = N1696;
  assign { r_n_237__31_, r_n_237__30_, r_n_237__29_, r_n_237__28_, r_n_237__27_, r_n_237__26_, r_n_237__25_, r_n_237__24_, r_n_237__23_, r_n_237__22_, r_n_237__21_, r_n_237__20_, r_n_237__19_, r_n_237__18_, r_n_237__17_, r_n_237__16_, r_n_237__15_, r_n_237__14_, r_n_237__13_, r_n_237__12_, r_n_237__11_, r_n_237__10_, r_n_237__9_, r_n_237__8_, r_n_237__7_, r_n_237__6_, r_n_237__5_, r_n_237__4_, r_n_237__3_, r_n_237__2_, r_n_237__1_, r_n_237__0_ } = (N474)? { r_238__31_, r_238__30_, r_238__29_, r_238__28_, r_238__27_, r_238__26_, r_238__25_, r_238__24_, r_238__23_, r_238__22_, r_238__21_, r_238__20_, r_238__19_, r_238__18_, r_238__17_, r_238__16_, r_238__15_, r_238__14_, r_238__13_, r_238__12_, r_238__11_, r_238__10_, r_238__9_, r_238__8_, r_238__7_, r_238__6_, r_238__5_, r_238__4_, r_238__3_, r_238__2_, r_238__1_, r_238__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N475)? data_i : 1'b0;
  assign N474 = sel_i[474];
  assign N475 = N1701;
  assign { r_n_238__31_, r_n_238__30_, r_n_238__29_, r_n_238__28_, r_n_238__27_, r_n_238__26_, r_n_238__25_, r_n_238__24_, r_n_238__23_, r_n_238__22_, r_n_238__21_, r_n_238__20_, r_n_238__19_, r_n_238__18_, r_n_238__17_, r_n_238__16_, r_n_238__15_, r_n_238__14_, r_n_238__13_, r_n_238__12_, r_n_238__11_, r_n_238__10_, r_n_238__9_, r_n_238__8_, r_n_238__7_, r_n_238__6_, r_n_238__5_, r_n_238__4_, r_n_238__3_, r_n_238__2_, r_n_238__1_, r_n_238__0_ } = (N476)? { r_239__31_, r_239__30_, r_239__29_, r_239__28_, r_239__27_, r_239__26_, r_239__25_, r_239__24_, r_239__23_, r_239__22_, r_239__21_, r_239__20_, r_239__19_, r_239__18_, r_239__17_, r_239__16_, r_239__15_, r_239__14_, r_239__13_, r_239__12_, r_239__11_, r_239__10_, r_239__9_, r_239__8_, r_239__7_, r_239__6_, r_239__5_, r_239__4_, r_239__3_, r_239__2_, r_239__1_, r_239__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N477)? data_i : 1'b0;
  assign N476 = sel_i[476];
  assign N477 = N1706;
  assign { r_n_239__31_, r_n_239__30_, r_n_239__29_, r_n_239__28_, r_n_239__27_, r_n_239__26_, r_n_239__25_, r_n_239__24_, r_n_239__23_, r_n_239__22_, r_n_239__21_, r_n_239__20_, r_n_239__19_, r_n_239__18_, r_n_239__17_, r_n_239__16_, r_n_239__15_, r_n_239__14_, r_n_239__13_, r_n_239__12_, r_n_239__11_, r_n_239__10_, r_n_239__9_, r_n_239__8_, r_n_239__7_, r_n_239__6_, r_n_239__5_, r_n_239__4_, r_n_239__3_, r_n_239__2_, r_n_239__1_, r_n_239__0_ } = (N478)? { r_240__31_, r_240__30_, r_240__29_, r_240__28_, r_240__27_, r_240__26_, r_240__25_, r_240__24_, r_240__23_, r_240__22_, r_240__21_, r_240__20_, r_240__19_, r_240__18_, r_240__17_, r_240__16_, r_240__15_, r_240__14_, r_240__13_, r_240__12_, r_240__11_, r_240__10_, r_240__9_, r_240__8_, r_240__7_, r_240__6_, r_240__5_, r_240__4_, r_240__3_, r_240__2_, r_240__1_, r_240__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N479)? data_i : 1'b0;
  assign N478 = sel_i[478];
  assign N479 = N1711;
  assign { r_n_240__31_, r_n_240__30_, r_n_240__29_, r_n_240__28_, r_n_240__27_, r_n_240__26_, r_n_240__25_, r_n_240__24_, r_n_240__23_, r_n_240__22_, r_n_240__21_, r_n_240__20_, r_n_240__19_, r_n_240__18_, r_n_240__17_, r_n_240__16_, r_n_240__15_, r_n_240__14_, r_n_240__13_, r_n_240__12_, r_n_240__11_, r_n_240__10_, r_n_240__9_, r_n_240__8_, r_n_240__7_, r_n_240__6_, r_n_240__5_, r_n_240__4_, r_n_240__3_, r_n_240__2_, r_n_240__1_, r_n_240__0_ } = (N480)? { r_241__31_, r_241__30_, r_241__29_, r_241__28_, r_241__27_, r_241__26_, r_241__25_, r_241__24_, r_241__23_, r_241__22_, r_241__21_, r_241__20_, r_241__19_, r_241__18_, r_241__17_, r_241__16_, r_241__15_, r_241__14_, r_241__13_, r_241__12_, r_241__11_, r_241__10_, r_241__9_, r_241__8_, r_241__7_, r_241__6_, r_241__5_, r_241__4_, r_241__3_, r_241__2_, r_241__1_, r_241__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N481)? data_i : 1'b0;
  assign N480 = sel_i[480];
  assign N481 = N1716;
  assign { r_n_241__31_, r_n_241__30_, r_n_241__29_, r_n_241__28_, r_n_241__27_, r_n_241__26_, r_n_241__25_, r_n_241__24_, r_n_241__23_, r_n_241__22_, r_n_241__21_, r_n_241__20_, r_n_241__19_, r_n_241__18_, r_n_241__17_, r_n_241__16_, r_n_241__15_, r_n_241__14_, r_n_241__13_, r_n_241__12_, r_n_241__11_, r_n_241__10_, r_n_241__9_, r_n_241__8_, r_n_241__7_, r_n_241__6_, r_n_241__5_, r_n_241__4_, r_n_241__3_, r_n_241__2_, r_n_241__1_, r_n_241__0_ } = (N482)? { r_242__31_, r_242__30_, r_242__29_, r_242__28_, r_242__27_, r_242__26_, r_242__25_, r_242__24_, r_242__23_, r_242__22_, r_242__21_, r_242__20_, r_242__19_, r_242__18_, r_242__17_, r_242__16_, r_242__15_, r_242__14_, r_242__13_, r_242__12_, r_242__11_, r_242__10_, r_242__9_, r_242__8_, r_242__7_, r_242__6_, r_242__5_, r_242__4_, r_242__3_, r_242__2_, r_242__1_, r_242__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N483)? data_i : 1'b0;
  assign N482 = sel_i[482];
  assign N483 = N1721;
  assign { r_n_242__31_, r_n_242__30_, r_n_242__29_, r_n_242__28_, r_n_242__27_, r_n_242__26_, r_n_242__25_, r_n_242__24_, r_n_242__23_, r_n_242__22_, r_n_242__21_, r_n_242__20_, r_n_242__19_, r_n_242__18_, r_n_242__17_, r_n_242__16_, r_n_242__15_, r_n_242__14_, r_n_242__13_, r_n_242__12_, r_n_242__11_, r_n_242__10_, r_n_242__9_, r_n_242__8_, r_n_242__7_, r_n_242__6_, r_n_242__5_, r_n_242__4_, r_n_242__3_, r_n_242__2_, r_n_242__1_, r_n_242__0_ } = (N484)? { r_243__31_, r_243__30_, r_243__29_, r_243__28_, r_243__27_, r_243__26_, r_243__25_, r_243__24_, r_243__23_, r_243__22_, r_243__21_, r_243__20_, r_243__19_, r_243__18_, r_243__17_, r_243__16_, r_243__15_, r_243__14_, r_243__13_, r_243__12_, r_243__11_, r_243__10_, r_243__9_, r_243__8_, r_243__7_, r_243__6_, r_243__5_, r_243__4_, r_243__3_, r_243__2_, r_243__1_, r_243__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N485)? data_i : 1'b0;
  assign N484 = sel_i[484];
  assign N485 = N1726;
  assign { r_n_243__31_, r_n_243__30_, r_n_243__29_, r_n_243__28_, r_n_243__27_, r_n_243__26_, r_n_243__25_, r_n_243__24_, r_n_243__23_, r_n_243__22_, r_n_243__21_, r_n_243__20_, r_n_243__19_, r_n_243__18_, r_n_243__17_, r_n_243__16_, r_n_243__15_, r_n_243__14_, r_n_243__13_, r_n_243__12_, r_n_243__11_, r_n_243__10_, r_n_243__9_, r_n_243__8_, r_n_243__7_, r_n_243__6_, r_n_243__5_, r_n_243__4_, r_n_243__3_, r_n_243__2_, r_n_243__1_, r_n_243__0_ } = (N486)? { r_244__31_, r_244__30_, r_244__29_, r_244__28_, r_244__27_, r_244__26_, r_244__25_, r_244__24_, r_244__23_, r_244__22_, r_244__21_, r_244__20_, r_244__19_, r_244__18_, r_244__17_, r_244__16_, r_244__15_, r_244__14_, r_244__13_, r_244__12_, r_244__11_, r_244__10_, r_244__9_, r_244__8_, r_244__7_, r_244__6_, r_244__5_, r_244__4_, r_244__3_, r_244__2_, r_244__1_, r_244__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N487)? data_i : 1'b0;
  assign N486 = sel_i[486];
  assign N487 = N1731;
  assign { r_n_244__31_, r_n_244__30_, r_n_244__29_, r_n_244__28_, r_n_244__27_, r_n_244__26_, r_n_244__25_, r_n_244__24_, r_n_244__23_, r_n_244__22_, r_n_244__21_, r_n_244__20_, r_n_244__19_, r_n_244__18_, r_n_244__17_, r_n_244__16_, r_n_244__15_, r_n_244__14_, r_n_244__13_, r_n_244__12_, r_n_244__11_, r_n_244__10_, r_n_244__9_, r_n_244__8_, r_n_244__7_, r_n_244__6_, r_n_244__5_, r_n_244__4_, r_n_244__3_, r_n_244__2_, r_n_244__1_, r_n_244__0_ } = (N488)? { r_245__31_, r_245__30_, r_245__29_, r_245__28_, r_245__27_, r_245__26_, r_245__25_, r_245__24_, r_245__23_, r_245__22_, r_245__21_, r_245__20_, r_245__19_, r_245__18_, r_245__17_, r_245__16_, r_245__15_, r_245__14_, r_245__13_, r_245__12_, r_245__11_, r_245__10_, r_245__9_, r_245__8_, r_245__7_, r_245__6_, r_245__5_, r_245__4_, r_245__3_, r_245__2_, r_245__1_, r_245__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N489)? data_i : 1'b0;
  assign N488 = sel_i[488];
  assign N489 = N1736;
  assign { r_n_245__31_, r_n_245__30_, r_n_245__29_, r_n_245__28_, r_n_245__27_, r_n_245__26_, r_n_245__25_, r_n_245__24_, r_n_245__23_, r_n_245__22_, r_n_245__21_, r_n_245__20_, r_n_245__19_, r_n_245__18_, r_n_245__17_, r_n_245__16_, r_n_245__15_, r_n_245__14_, r_n_245__13_, r_n_245__12_, r_n_245__11_, r_n_245__10_, r_n_245__9_, r_n_245__8_, r_n_245__7_, r_n_245__6_, r_n_245__5_, r_n_245__4_, r_n_245__3_, r_n_245__2_, r_n_245__1_, r_n_245__0_ } = (N490)? { r_246__31_, r_246__30_, r_246__29_, r_246__28_, r_246__27_, r_246__26_, r_246__25_, r_246__24_, r_246__23_, r_246__22_, r_246__21_, r_246__20_, r_246__19_, r_246__18_, r_246__17_, r_246__16_, r_246__15_, r_246__14_, r_246__13_, r_246__12_, r_246__11_, r_246__10_, r_246__9_, r_246__8_, r_246__7_, r_246__6_, r_246__5_, r_246__4_, r_246__3_, r_246__2_, r_246__1_, r_246__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N491)? data_i : 1'b0;
  assign N490 = sel_i[490];
  assign N491 = N1741;
  assign { r_n_246__31_, r_n_246__30_, r_n_246__29_, r_n_246__28_, r_n_246__27_, r_n_246__26_, r_n_246__25_, r_n_246__24_, r_n_246__23_, r_n_246__22_, r_n_246__21_, r_n_246__20_, r_n_246__19_, r_n_246__18_, r_n_246__17_, r_n_246__16_, r_n_246__15_, r_n_246__14_, r_n_246__13_, r_n_246__12_, r_n_246__11_, r_n_246__10_, r_n_246__9_, r_n_246__8_, r_n_246__7_, r_n_246__6_, r_n_246__5_, r_n_246__4_, r_n_246__3_, r_n_246__2_, r_n_246__1_, r_n_246__0_ } = (N492)? { r_247__31_, r_247__30_, r_247__29_, r_247__28_, r_247__27_, r_247__26_, r_247__25_, r_247__24_, r_247__23_, r_247__22_, r_247__21_, r_247__20_, r_247__19_, r_247__18_, r_247__17_, r_247__16_, r_247__15_, r_247__14_, r_247__13_, r_247__12_, r_247__11_, r_247__10_, r_247__9_, r_247__8_, r_247__7_, r_247__6_, r_247__5_, r_247__4_, r_247__3_, r_247__2_, r_247__1_, r_247__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N493)? data_i : 1'b0;
  assign N492 = sel_i[492];
  assign N493 = N1746;
  assign { r_n_247__31_, r_n_247__30_, r_n_247__29_, r_n_247__28_, r_n_247__27_, r_n_247__26_, r_n_247__25_, r_n_247__24_, r_n_247__23_, r_n_247__22_, r_n_247__21_, r_n_247__20_, r_n_247__19_, r_n_247__18_, r_n_247__17_, r_n_247__16_, r_n_247__15_, r_n_247__14_, r_n_247__13_, r_n_247__12_, r_n_247__11_, r_n_247__10_, r_n_247__9_, r_n_247__8_, r_n_247__7_, r_n_247__6_, r_n_247__5_, r_n_247__4_, r_n_247__3_, r_n_247__2_, r_n_247__1_, r_n_247__0_ } = (N494)? { r_248__31_, r_248__30_, r_248__29_, r_248__28_, r_248__27_, r_248__26_, r_248__25_, r_248__24_, r_248__23_, r_248__22_, r_248__21_, r_248__20_, r_248__19_, r_248__18_, r_248__17_, r_248__16_, r_248__15_, r_248__14_, r_248__13_, r_248__12_, r_248__11_, r_248__10_, r_248__9_, r_248__8_, r_248__7_, r_248__6_, r_248__5_, r_248__4_, r_248__3_, r_248__2_, r_248__1_, r_248__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N495)? data_i : 1'b0;
  assign N494 = sel_i[494];
  assign N495 = N1751;
  assign { r_n_248__31_, r_n_248__30_, r_n_248__29_, r_n_248__28_, r_n_248__27_, r_n_248__26_, r_n_248__25_, r_n_248__24_, r_n_248__23_, r_n_248__22_, r_n_248__21_, r_n_248__20_, r_n_248__19_, r_n_248__18_, r_n_248__17_, r_n_248__16_, r_n_248__15_, r_n_248__14_, r_n_248__13_, r_n_248__12_, r_n_248__11_, r_n_248__10_, r_n_248__9_, r_n_248__8_, r_n_248__7_, r_n_248__6_, r_n_248__5_, r_n_248__4_, r_n_248__3_, r_n_248__2_, r_n_248__1_, r_n_248__0_ } = (N496)? { r_249__31_, r_249__30_, r_249__29_, r_249__28_, r_249__27_, r_249__26_, r_249__25_, r_249__24_, r_249__23_, r_249__22_, r_249__21_, r_249__20_, r_249__19_, r_249__18_, r_249__17_, r_249__16_, r_249__15_, r_249__14_, r_249__13_, r_249__12_, r_249__11_, r_249__10_, r_249__9_, r_249__8_, r_249__7_, r_249__6_, r_249__5_, r_249__4_, r_249__3_, r_249__2_, r_249__1_, r_249__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N497)? data_i : 1'b0;
  assign N496 = sel_i[496];
  assign N497 = N1756;
  assign { r_n_249__31_, r_n_249__30_, r_n_249__29_, r_n_249__28_, r_n_249__27_, r_n_249__26_, r_n_249__25_, r_n_249__24_, r_n_249__23_, r_n_249__22_, r_n_249__21_, r_n_249__20_, r_n_249__19_, r_n_249__18_, r_n_249__17_, r_n_249__16_, r_n_249__15_, r_n_249__14_, r_n_249__13_, r_n_249__12_, r_n_249__11_, r_n_249__10_, r_n_249__9_, r_n_249__8_, r_n_249__7_, r_n_249__6_, r_n_249__5_, r_n_249__4_, r_n_249__3_, r_n_249__2_, r_n_249__1_, r_n_249__0_ } = (N498)? { r_250__31_, r_250__30_, r_250__29_, r_250__28_, r_250__27_, r_250__26_, r_250__25_, r_250__24_, r_250__23_, r_250__22_, r_250__21_, r_250__20_, r_250__19_, r_250__18_, r_250__17_, r_250__16_, r_250__15_, r_250__14_, r_250__13_, r_250__12_, r_250__11_, r_250__10_, r_250__9_, r_250__8_, r_250__7_, r_250__6_, r_250__5_, r_250__4_, r_250__3_, r_250__2_, r_250__1_, r_250__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N499)? data_i : 1'b0;
  assign N498 = sel_i[498];
  assign N499 = N1761;
  assign { r_n_250__31_, r_n_250__30_, r_n_250__29_, r_n_250__28_, r_n_250__27_, r_n_250__26_, r_n_250__25_, r_n_250__24_, r_n_250__23_, r_n_250__22_, r_n_250__21_, r_n_250__20_, r_n_250__19_, r_n_250__18_, r_n_250__17_, r_n_250__16_, r_n_250__15_, r_n_250__14_, r_n_250__13_, r_n_250__12_, r_n_250__11_, r_n_250__10_, r_n_250__9_, r_n_250__8_, r_n_250__7_, r_n_250__6_, r_n_250__5_, r_n_250__4_, r_n_250__3_, r_n_250__2_, r_n_250__1_, r_n_250__0_ } = (N500)? { r_251__31_, r_251__30_, r_251__29_, r_251__28_, r_251__27_, r_251__26_, r_251__25_, r_251__24_, r_251__23_, r_251__22_, r_251__21_, r_251__20_, r_251__19_, r_251__18_, r_251__17_, r_251__16_, r_251__15_, r_251__14_, r_251__13_, r_251__12_, r_251__11_, r_251__10_, r_251__9_, r_251__8_, r_251__7_, r_251__6_, r_251__5_, r_251__4_, r_251__3_, r_251__2_, r_251__1_, r_251__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N501)? data_i : 1'b0;
  assign N500 = sel_i[500];
  assign N501 = N1766;
  assign { r_n_251__31_, r_n_251__30_, r_n_251__29_, r_n_251__28_, r_n_251__27_, r_n_251__26_, r_n_251__25_, r_n_251__24_, r_n_251__23_, r_n_251__22_, r_n_251__21_, r_n_251__20_, r_n_251__19_, r_n_251__18_, r_n_251__17_, r_n_251__16_, r_n_251__15_, r_n_251__14_, r_n_251__13_, r_n_251__12_, r_n_251__11_, r_n_251__10_, r_n_251__9_, r_n_251__8_, r_n_251__7_, r_n_251__6_, r_n_251__5_, r_n_251__4_, r_n_251__3_, r_n_251__2_, r_n_251__1_, r_n_251__0_ } = (N502)? { r_252__31_, r_252__30_, r_252__29_, r_252__28_, r_252__27_, r_252__26_, r_252__25_, r_252__24_, r_252__23_, r_252__22_, r_252__21_, r_252__20_, r_252__19_, r_252__18_, r_252__17_, r_252__16_, r_252__15_, r_252__14_, r_252__13_, r_252__12_, r_252__11_, r_252__10_, r_252__9_, r_252__8_, r_252__7_, r_252__6_, r_252__5_, r_252__4_, r_252__3_, r_252__2_, r_252__1_, r_252__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N503)? data_i : 1'b0;
  assign N502 = sel_i[502];
  assign N503 = N1771;
  assign { r_n_252__31_, r_n_252__30_, r_n_252__29_, r_n_252__28_, r_n_252__27_, r_n_252__26_, r_n_252__25_, r_n_252__24_, r_n_252__23_, r_n_252__22_, r_n_252__21_, r_n_252__20_, r_n_252__19_, r_n_252__18_, r_n_252__17_, r_n_252__16_, r_n_252__15_, r_n_252__14_, r_n_252__13_, r_n_252__12_, r_n_252__11_, r_n_252__10_, r_n_252__9_, r_n_252__8_, r_n_252__7_, r_n_252__6_, r_n_252__5_, r_n_252__4_, r_n_252__3_, r_n_252__2_, r_n_252__1_, r_n_252__0_ } = (N504)? { r_253__31_, r_253__30_, r_253__29_, r_253__28_, r_253__27_, r_253__26_, r_253__25_, r_253__24_, r_253__23_, r_253__22_, r_253__21_, r_253__20_, r_253__19_, r_253__18_, r_253__17_, r_253__16_, r_253__15_, r_253__14_, r_253__13_, r_253__12_, r_253__11_, r_253__10_, r_253__9_, r_253__8_, r_253__7_, r_253__6_, r_253__5_, r_253__4_, r_253__3_, r_253__2_, r_253__1_, r_253__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N505)? data_i : 1'b0;
  assign N504 = sel_i[504];
  assign N505 = N1776;
  assign { r_n_253__31_, r_n_253__30_, r_n_253__29_, r_n_253__28_, r_n_253__27_, r_n_253__26_, r_n_253__25_, r_n_253__24_, r_n_253__23_, r_n_253__22_, r_n_253__21_, r_n_253__20_, r_n_253__19_, r_n_253__18_, r_n_253__17_, r_n_253__16_, r_n_253__15_, r_n_253__14_, r_n_253__13_, r_n_253__12_, r_n_253__11_, r_n_253__10_, r_n_253__9_, r_n_253__8_, r_n_253__7_, r_n_253__6_, r_n_253__5_, r_n_253__4_, r_n_253__3_, r_n_253__2_, r_n_253__1_, r_n_253__0_ } = (N506)? { r_254__31_, r_254__30_, r_254__29_, r_254__28_, r_254__27_, r_254__26_, r_254__25_, r_254__24_, r_254__23_, r_254__22_, r_254__21_, r_254__20_, r_254__19_, r_254__18_, r_254__17_, r_254__16_, r_254__15_, r_254__14_, r_254__13_, r_254__12_, r_254__11_, r_254__10_, r_254__9_, r_254__8_, r_254__7_, r_254__6_, r_254__5_, r_254__4_, r_254__3_, r_254__2_, r_254__1_, r_254__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N507)? data_i : 1'b0;
  assign N506 = sel_i[506];
  assign N507 = N1781;
  assign { r_n_254__31_, r_n_254__30_, r_n_254__29_, r_n_254__28_, r_n_254__27_, r_n_254__26_, r_n_254__25_, r_n_254__24_, r_n_254__23_, r_n_254__22_, r_n_254__21_, r_n_254__20_, r_n_254__19_, r_n_254__18_, r_n_254__17_, r_n_254__16_, r_n_254__15_, r_n_254__14_, r_n_254__13_, r_n_254__12_, r_n_254__11_, r_n_254__10_, r_n_254__9_, r_n_254__8_, r_n_254__7_, r_n_254__6_, r_n_254__5_, r_n_254__4_, r_n_254__3_, r_n_254__2_, r_n_254__1_, r_n_254__0_ } = (N508)? { r_255__31_, r_255__30_, r_255__29_, r_255__28_, r_255__27_, r_255__26_, r_255__25_, r_255__24_, r_255__23_, r_255__22_, r_255__21_, r_255__20_, r_255__19_, r_255__18_, r_255__17_, r_255__16_, r_255__15_, r_255__14_, r_255__13_, r_255__12_, r_255__11_, r_255__10_, r_255__9_, r_255__8_, r_255__7_, r_255__6_, r_255__5_, r_255__4_, r_255__3_, r_255__2_, r_255__1_, r_255__0_ } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N509)? data_i : 1'b0;
  assign N508 = sel_i[508];
  assign N509 = N1786;
  assign { r_n_255__31_, r_n_255__30_, r_n_255__29_, r_n_255__28_, r_n_255__27_, r_n_255__26_, r_n_255__25_, r_n_255__24_, r_n_255__23_, r_n_255__22_, r_n_255__21_, r_n_255__20_, r_n_255__19_, r_n_255__18_, r_n_255__17_, r_n_255__16_, r_n_255__15_, r_n_255__14_, r_n_255__13_, r_n_255__12_, r_n_255__11_, r_n_255__10_, r_n_255__9_, r_n_255__8_, r_n_255__7_, r_n_255__6_, r_n_255__5_, r_n_255__4_, r_n_255__3_, r_n_255__2_, r_n_255__1_, r_n_255__0_ } = (N510)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    (N511)? data_i : 1'b0;
  assign N510 = sel_i[510];
  assign N511 = N1791;
  assign N513 = ~sel_i[1];
  assign N515 = N512 | N514;
  assign N518 = ~sel_i[3];
  assign N520 = N517 | N519;
  assign N523 = ~sel_i[5];
  assign N525 = N522 | N524;
  assign N528 = ~sel_i[7];
  assign N530 = N527 | N529;
  assign N533 = ~sel_i[9];
  assign N535 = N532 | N534;
  assign N538 = ~sel_i[11];
  assign N540 = N537 | N539;
  assign N543 = ~sel_i[13];
  assign N545 = N542 | N544;
  assign N548 = ~sel_i[15];
  assign N550 = N547 | N549;
  assign N553 = ~sel_i[17];
  assign N555 = N552 | N554;
  assign N558 = ~sel_i[19];
  assign N560 = N557 | N559;
  assign N563 = ~sel_i[21];
  assign N565 = N562 | N564;
  assign N568 = ~sel_i[23];
  assign N570 = N567 | N569;
  assign N573 = ~sel_i[25];
  assign N575 = N572 | N574;
  assign N578 = ~sel_i[27];
  assign N580 = N577 | N579;
  assign N583 = ~sel_i[29];
  assign N585 = N582 | N584;
  assign N588 = ~sel_i[31];
  assign N590 = N587 | N589;
  assign N593 = ~sel_i[33];
  assign N595 = N592 | N594;
  assign N598 = ~sel_i[35];
  assign N600 = N597 | N599;
  assign N603 = ~sel_i[37];
  assign N605 = N602 | N604;
  assign N608 = ~sel_i[39];
  assign N610 = N607 | N609;
  assign N613 = ~sel_i[41];
  assign N615 = N612 | N614;
  assign N618 = ~sel_i[43];
  assign N620 = N617 | N619;
  assign N623 = ~sel_i[45];
  assign N625 = N622 | N624;
  assign N628 = ~sel_i[47];
  assign N630 = N627 | N629;
  assign N633 = ~sel_i[49];
  assign N635 = N632 | N634;
  assign N638 = ~sel_i[51];
  assign N640 = N637 | N639;
  assign N643 = ~sel_i[53];
  assign N645 = N642 | N644;
  assign N648 = ~sel_i[55];
  assign N650 = N647 | N649;
  assign N653 = ~sel_i[57];
  assign N655 = N652 | N654;
  assign N658 = ~sel_i[59];
  assign N660 = N657 | N659;
  assign N663 = ~sel_i[61];
  assign N665 = N662 | N664;
  assign N668 = ~sel_i[63];
  assign N670 = N667 | N669;
  assign N673 = ~sel_i[65];
  assign N675 = N672 | N674;
  assign N678 = ~sel_i[67];
  assign N680 = N677 | N679;
  assign N683 = ~sel_i[69];
  assign N685 = N682 | N684;
  assign N688 = ~sel_i[71];
  assign N690 = N687 | N689;
  assign N693 = ~sel_i[73];
  assign N695 = N692 | N694;
  assign N698 = ~sel_i[75];
  assign N700 = N697 | N699;
  assign N703 = ~sel_i[77];
  assign N705 = N702 | N704;
  assign N708 = ~sel_i[79];
  assign N710 = N707 | N709;
  assign N713 = ~sel_i[81];
  assign N715 = N712 | N714;
  assign N718 = ~sel_i[83];
  assign N720 = N717 | N719;
  assign N723 = ~sel_i[85];
  assign N725 = N722 | N724;
  assign N728 = ~sel_i[87];
  assign N730 = N727 | N729;
  assign N733 = ~sel_i[89];
  assign N735 = N732 | N734;
  assign N738 = ~sel_i[91];
  assign N740 = N737 | N739;
  assign N743 = ~sel_i[93];
  assign N745 = N742 | N744;
  assign N748 = ~sel_i[95];
  assign N750 = N747 | N749;
  assign N753 = ~sel_i[97];
  assign N755 = N752 | N754;
  assign N758 = ~sel_i[99];
  assign N760 = N757 | N759;
  assign N763 = ~sel_i[101];
  assign N765 = N762 | N764;
  assign N768 = ~sel_i[103];
  assign N770 = N767 | N769;
  assign N773 = ~sel_i[105];
  assign N775 = N772 | N774;
  assign N778 = ~sel_i[107];
  assign N780 = N777 | N779;
  assign N783 = ~sel_i[109];
  assign N785 = N782 | N784;
  assign N788 = ~sel_i[111];
  assign N790 = N787 | N789;
  assign N793 = ~sel_i[113];
  assign N795 = N792 | N794;
  assign N798 = ~sel_i[115];
  assign N800 = N797 | N799;
  assign N803 = ~sel_i[117];
  assign N805 = N802 | N804;
  assign N808 = ~sel_i[119];
  assign N810 = N807 | N809;
  assign N813 = ~sel_i[121];
  assign N815 = N812 | N814;
  assign N818 = ~sel_i[123];
  assign N820 = N817 | N819;
  assign N823 = ~sel_i[125];
  assign N825 = N822 | N824;
  assign N828 = ~sel_i[127];
  assign N830 = N827 | N829;
  assign N833 = ~sel_i[129];
  assign N835 = N832 | N834;
  assign N838 = ~sel_i[131];
  assign N840 = N837 | N839;
  assign N843 = ~sel_i[133];
  assign N845 = N842 | N844;
  assign N848 = ~sel_i[135];
  assign N850 = N847 | N849;
  assign N853 = ~sel_i[137];
  assign N855 = N852 | N854;
  assign N858 = ~sel_i[139];
  assign N860 = N857 | N859;
  assign N863 = ~sel_i[141];
  assign N865 = N862 | N864;
  assign N868 = ~sel_i[143];
  assign N870 = N867 | N869;
  assign N873 = ~sel_i[145];
  assign N875 = N872 | N874;
  assign N878 = ~sel_i[147];
  assign N880 = N877 | N879;
  assign N883 = ~sel_i[149];
  assign N885 = N882 | N884;
  assign N888 = ~sel_i[151];
  assign N890 = N887 | N889;
  assign N893 = ~sel_i[153];
  assign N895 = N892 | N894;
  assign N898 = ~sel_i[155];
  assign N900 = N897 | N899;
  assign N903 = ~sel_i[157];
  assign N905 = N902 | N904;
  assign N908 = ~sel_i[159];
  assign N910 = N907 | N909;
  assign N913 = ~sel_i[161];
  assign N915 = N912 | N914;
  assign N918 = ~sel_i[163];
  assign N920 = N917 | N919;
  assign N923 = ~sel_i[165];
  assign N925 = N922 | N924;
  assign N928 = ~sel_i[167];
  assign N930 = N927 | N929;
  assign N933 = ~sel_i[169];
  assign N935 = N932 | N934;
  assign N938 = ~sel_i[171];
  assign N940 = N937 | N939;
  assign N943 = ~sel_i[173];
  assign N945 = N942 | N944;
  assign N948 = ~sel_i[175];
  assign N950 = N947 | N949;
  assign N953 = ~sel_i[177];
  assign N955 = N952 | N954;
  assign N958 = ~sel_i[179];
  assign N960 = N957 | N959;
  assign N963 = ~sel_i[181];
  assign N965 = N962 | N964;
  assign N968 = ~sel_i[183];
  assign N970 = N967 | N969;
  assign N973 = ~sel_i[185];
  assign N975 = N972 | N974;
  assign N978 = ~sel_i[187];
  assign N980 = N977 | N979;
  assign N983 = ~sel_i[189];
  assign N985 = N982 | N984;
  assign N988 = ~sel_i[191];
  assign N990 = N987 | N989;
  assign N993 = ~sel_i[193];
  assign N995 = N992 | N994;
  assign N998 = ~sel_i[195];
  assign N1000 = N997 | N999;
  assign N1003 = ~sel_i[197];
  assign N1005 = N1002 | N1004;
  assign N1008 = ~sel_i[199];
  assign N1010 = N1007 | N1009;
  assign N1013 = ~sel_i[201];
  assign N1015 = N1012 | N1014;
  assign N1018 = ~sel_i[203];
  assign N1020 = N1017 | N1019;
  assign N1023 = ~sel_i[205];
  assign N1025 = N1022 | N1024;
  assign N1028 = ~sel_i[207];
  assign N1030 = N1027 | N1029;
  assign N1033 = ~sel_i[209];
  assign N1035 = N1032 | N1034;
  assign N1038 = ~sel_i[211];
  assign N1040 = N1037 | N1039;
  assign N1043 = ~sel_i[213];
  assign N1045 = N1042 | N1044;
  assign N1048 = ~sel_i[215];
  assign N1050 = N1047 | N1049;
  assign N1053 = ~sel_i[217];
  assign N1055 = N1052 | N1054;
  assign N1058 = ~sel_i[219];
  assign N1060 = N1057 | N1059;
  assign N1063 = ~sel_i[221];
  assign N1065 = N1062 | N1064;
  assign N1068 = ~sel_i[223];
  assign N1070 = N1067 | N1069;
  assign N1073 = ~sel_i[225];
  assign N1075 = N1072 | N1074;
  assign N1078 = ~sel_i[227];
  assign N1080 = N1077 | N1079;
  assign N1083 = ~sel_i[229];
  assign N1085 = N1082 | N1084;
  assign N1088 = ~sel_i[231];
  assign N1090 = N1087 | N1089;
  assign N1093 = ~sel_i[233];
  assign N1095 = N1092 | N1094;
  assign N1098 = ~sel_i[235];
  assign N1100 = N1097 | N1099;
  assign N1103 = ~sel_i[237];
  assign N1105 = N1102 | N1104;
  assign N1108 = ~sel_i[239];
  assign N1110 = N1107 | N1109;
  assign N1113 = ~sel_i[241];
  assign N1115 = N1112 | N1114;
  assign N1118 = ~sel_i[243];
  assign N1120 = N1117 | N1119;
  assign N1123 = ~sel_i[245];
  assign N1125 = N1122 | N1124;
  assign N1128 = ~sel_i[247];
  assign N1130 = N1127 | N1129;
  assign N1133 = ~sel_i[249];
  assign N1135 = N1132 | N1134;
  assign N1138 = ~sel_i[251];
  assign N1140 = N1137 | N1139;
  assign N1143 = ~sel_i[253];
  assign N1145 = N1142 | N1144;
  assign N1148 = ~sel_i[255];
  assign N1150 = N1147 | N1149;
  assign N1153 = ~sel_i[257];
  assign N1155 = N1152 | N1154;
  assign N1158 = ~sel_i[259];
  assign N1160 = N1157 | N1159;
  assign N1163 = ~sel_i[261];
  assign N1165 = N1162 | N1164;
  assign N1168 = ~sel_i[263];
  assign N1170 = N1167 | N1169;
  assign N1173 = ~sel_i[265];
  assign N1175 = N1172 | N1174;
  assign N1178 = ~sel_i[267];
  assign N1180 = N1177 | N1179;
  assign N1183 = ~sel_i[269];
  assign N1185 = N1182 | N1184;
  assign N1188 = ~sel_i[271];
  assign N1190 = N1187 | N1189;
  assign N1193 = ~sel_i[273];
  assign N1195 = N1192 | N1194;
  assign N1198 = ~sel_i[275];
  assign N1200 = N1197 | N1199;
  assign N1203 = ~sel_i[277];
  assign N1205 = N1202 | N1204;
  assign N1208 = ~sel_i[279];
  assign N1210 = N1207 | N1209;
  assign N1213 = ~sel_i[281];
  assign N1215 = N1212 | N1214;
  assign N1218 = ~sel_i[283];
  assign N1220 = N1217 | N1219;
  assign N1223 = ~sel_i[285];
  assign N1225 = N1222 | N1224;
  assign N1228 = ~sel_i[287];
  assign N1230 = N1227 | N1229;
  assign N1233 = ~sel_i[289];
  assign N1235 = N1232 | N1234;
  assign N1238 = ~sel_i[291];
  assign N1240 = N1237 | N1239;
  assign N1243 = ~sel_i[293];
  assign N1245 = N1242 | N1244;
  assign N1248 = ~sel_i[295];
  assign N1250 = N1247 | N1249;
  assign N1253 = ~sel_i[297];
  assign N1255 = N1252 | N1254;
  assign N1258 = ~sel_i[299];
  assign N1260 = N1257 | N1259;
  assign N1263 = ~sel_i[301];
  assign N1265 = N1262 | N1264;
  assign N1268 = ~sel_i[303];
  assign N1270 = N1267 | N1269;
  assign N1273 = ~sel_i[305];
  assign N1275 = N1272 | N1274;
  assign N1278 = ~sel_i[307];
  assign N1280 = N1277 | N1279;
  assign N1283 = ~sel_i[309];
  assign N1285 = N1282 | N1284;
  assign N1288 = ~sel_i[311];
  assign N1290 = N1287 | N1289;
  assign N1293 = ~sel_i[313];
  assign N1295 = N1292 | N1294;
  assign N1298 = ~sel_i[315];
  assign N1300 = N1297 | N1299;
  assign N1303 = ~sel_i[317];
  assign N1305 = N1302 | N1304;
  assign N1308 = ~sel_i[319];
  assign N1310 = N1307 | N1309;
  assign N1313 = ~sel_i[321];
  assign N1315 = N1312 | N1314;
  assign N1318 = ~sel_i[323];
  assign N1320 = N1317 | N1319;
  assign N1323 = ~sel_i[325];
  assign N1325 = N1322 | N1324;
  assign N1328 = ~sel_i[327];
  assign N1330 = N1327 | N1329;
  assign N1333 = ~sel_i[329];
  assign N1335 = N1332 | N1334;
  assign N1338 = ~sel_i[331];
  assign N1340 = N1337 | N1339;
  assign N1343 = ~sel_i[333];
  assign N1345 = N1342 | N1344;
  assign N1348 = ~sel_i[335];
  assign N1350 = N1347 | N1349;
  assign N1353 = ~sel_i[337];
  assign N1355 = N1352 | N1354;
  assign N1358 = ~sel_i[339];
  assign N1360 = N1357 | N1359;
  assign N1363 = ~sel_i[341];
  assign N1365 = N1362 | N1364;
  assign N1368 = ~sel_i[343];
  assign N1370 = N1367 | N1369;
  assign N1373 = ~sel_i[345];
  assign N1375 = N1372 | N1374;
  assign N1378 = ~sel_i[347];
  assign N1380 = N1377 | N1379;
  assign N1383 = ~sel_i[349];
  assign N1385 = N1382 | N1384;
  assign N1388 = ~sel_i[351];
  assign N1390 = N1387 | N1389;
  assign N1393 = ~sel_i[353];
  assign N1395 = N1392 | N1394;
  assign N1398 = ~sel_i[355];
  assign N1400 = N1397 | N1399;
  assign N1403 = ~sel_i[357];
  assign N1405 = N1402 | N1404;
  assign N1408 = ~sel_i[359];
  assign N1410 = N1407 | N1409;
  assign N1413 = ~sel_i[361];
  assign N1415 = N1412 | N1414;
  assign N1418 = ~sel_i[363];
  assign N1420 = N1417 | N1419;
  assign N1423 = ~sel_i[365];
  assign N1425 = N1422 | N1424;
  assign N1428 = ~sel_i[367];
  assign N1430 = N1427 | N1429;
  assign N1433 = ~sel_i[369];
  assign N1435 = N1432 | N1434;
  assign N1438 = ~sel_i[371];
  assign N1440 = N1437 | N1439;
  assign N1443 = ~sel_i[373];
  assign N1445 = N1442 | N1444;
  assign N1448 = ~sel_i[375];
  assign N1450 = N1447 | N1449;
  assign N1453 = ~sel_i[377];
  assign N1455 = N1452 | N1454;
  assign N1458 = ~sel_i[379];
  assign N1460 = N1457 | N1459;
  assign N1463 = ~sel_i[381];
  assign N1465 = N1462 | N1464;
  assign N1468 = ~sel_i[383];
  assign N1470 = N1467 | N1469;
  assign N1473 = ~sel_i[385];
  assign N1475 = N1472 | N1474;
  assign N1478 = ~sel_i[387];
  assign N1480 = N1477 | N1479;
  assign N1483 = ~sel_i[389];
  assign N1485 = N1482 | N1484;
  assign N1488 = ~sel_i[391];
  assign N1490 = N1487 | N1489;
  assign N1493 = ~sel_i[393];
  assign N1495 = N1492 | N1494;
  assign N1498 = ~sel_i[395];
  assign N1500 = N1497 | N1499;
  assign N1503 = ~sel_i[397];
  assign N1505 = N1502 | N1504;
  assign N1508 = ~sel_i[399];
  assign N1510 = N1507 | N1509;
  assign N1513 = ~sel_i[401];
  assign N1515 = N1512 | N1514;
  assign N1518 = ~sel_i[403];
  assign N1520 = N1517 | N1519;
  assign N1523 = ~sel_i[405];
  assign N1525 = N1522 | N1524;
  assign N1528 = ~sel_i[407];
  assign N1530 = N1527 | N1529;
  assign N1533 = ~sel_i[409];
  assign N1535 = N1532 | N1534;
  assign N1538 = ~sel_i[411];
  assign N1540 = N1537 | N1539;
  assign N1543 = ~sel_i[413];
  assign N1545 = N1542 | N1544;
  assign N1548 = ~sel_i[415];
  assign N1550 = N1547 | N1549;
  assign N1553 = ~sel_i[417];
  assign N1555 = N1552 | N1554;
  assign N1558 = ~sel_i[419];
  assign N1560 = N1557 | N1559;
  assign N1563 = ~sel_i[421];
  assign N1565 = N1562 | N1564;
  assign N1568 = ~sel_i[423];
  assign N1570 = N1567 | N1569;
  assign N1573 = ~sel_i[425];
  assign N1575 = N1572 | N1574;
  assign N1578 = ~sel_i[427];
  assign N1580 = N1577 | N1579;
  assign N1583 = ~sel_i[429];
  assign N1585 = N1582 | N1584;
  assign N1588 = ~sel_i[431];
  assign N1590 = N1587 | N1589;
  assign N1593 = ~sel_i[433];
  assign N1595 = N1592 | N1594;
  assign N1598 = ~sel_i[435];
  assign N1600 = N1597 | N1599;
  assign N1603 = ~sel_i[437];
  assign N1605 = N1602 | N1604;
  assign N1608 = ~sel_i[439];
  assign N1610 = N1607 | N1609;
  assign N1613 = ~sel_i[441];
  assign N1615 = N1612 | N1614;
  assign N1618 = ~sel_i[443];
  assign N1620 = N1617 | N1619;
  assign N1623 = ~sel_i[445];
  assign N1625 = N1622 | N1624;
  assign N1628 = ~sel_i[447];
  assign N1630 = N1627 | N1629;
  assign N1633 = ~sel_i[449];
  assign N1635 = N1632 | N1634;
  assign N1638 = ~sel_i[451];
  assign N1640 = N1637 | N1639;
  assign N1643 = ~sel_i[453];
  assign N1645 = N1642 | N1644;
  assign N1648 = ~sel_i[455];
  assign N1650 = N1647 | N1649;
  assign N1653 = ~sel_i[457];
  assign N1655 = N1652 | N1654;
  assign N1658 = ~sel_i[459];
  assign N1660 = N1657 | N1659;
  assign N1663 = ~sel_i[461];
  assign N1665 = N1662 | N1664;
  assign N1668 = ~sel_i[463];
  assign N1670 = N1667 | N1669;
  assign N1673 = ~sel_i[465];
  assign N1675 = N1672 | N1674;
  assign N1678 = ~sel_i[467];
  assign N1680 = N1677 | N1679;
  assign N1683 = ~sel_i[469];
  assign N1685 = N1682 | N1684;
  assign N1688 = ~sel_i[471];
  assign N1690 = N1687 | N1689;
  assign N1693 = ~sel_i[473];
  assign N1695 = N1692 | N1694;
  assign N1698 = ~sel_i[475];
  assign N1700 = N1697 | N1699;
  assign N1703 = ~sel_i[477];
  assign N1705 = N1702 | N1704;
  assign N1708 = ~sel_i[479];
  assign N1710 = N1707 | N1709;
  assign N1713 = ~sel_i[481];
  assign N1715 = N1712 | N1714;
  assign N1718 = ~sel_i[483];
  assign N1720 = N1717 | N1719;
  assign N1723 = ~sel_i[485];
  assign N1725 = N1722 | N1724;
  assign N1728 = ~sel_i[487];
  assign N1730 = N1727 | N1729;
  assign N1733 = ~sel_i[489];
  assign N1735 = N1732 | N1734;
  assign N1738 = ~sel_i[491];
  assign N1740 = N1737 | N1739;
  assign N1743 = ~sel_i[493];
  assign N1745 = N1742 | N1744;
  assign N1748 = ~sel_i[495];
  assign N1750 = N1747 | N1749;
  assign N1753 = ~sel_i[497];
  assign N1755 = N1752 | N1754;
  assign N1758 = ~sel_i[499];
  assign N1760 = N1757 | N1759;
  assign N1763 = ~sel_i[501];
  assign N1765 = N1762 | N1764;
  assign N1768 = ~sel_i[503];
  assign N1770 = N1767 | N1769;
  assign N1773 = ~sel_i[505];
  assign N1775 = N1772 | N1774;
  assign N1778 = ~sel_i[507];
  assign N1780 = N1777 | N1779;
  assign N1783 = ~sel_i[509];
  assign N1785 = N1782 | N1784;
  assign N1788 = ~sel_i[511];
  assign N1790 = N1787 | N1789;
  assign N1792 = ~N515;
  assign N1793 = ~N520;
  assign N1794 = ~N525;
  assign N1795 = ~N530;
  assign N1796 = ~N535;
  assign N1797 = ~N540;
  assign N1798 = ~N545;
  assign N1799 = ~N550;
  assign N1800 = ~N555;
  assign N1801 = ~N560;
  assign N1802 = ~N565;
  assign N1803 = ~N570;
  assign N1804 = ~N575;
  assign N1805 = ~N580;
  assign N1806 = ~N585;
  assign N1807 = ~N590;
  assign N1808 = ~N595;
  assign N1809 = ~N600;
  assign N1810 = ~N605;
  assign N1811 = ~N610;
  assign N1812 = ~N615;
  assign N1813 = ~N620;
  assign N1814 = ~N625;
  assign N1815 = ~N630;
  assign N1816 = ~N635;
  assign N1817 = ~N640;
  assign N1818 = ~N645;
  assign N1819 = ~N650;
  assign N1820 = ~N655;
  assign N1821 = ~N660;
  assign N1822 = ~N665;
  assign N1823 = ~N670;
  assign N1824 = ~N675;
  assign N1825 = ~N680;
  assign N1826 = ~N685;
  assign N1827 = ~N690;
  assign N1828 = ~N695;
  assign N1829 = ~N700;
  assign N1830 = ~N705;
  assign N1831 = ~N710;
  assign N1832 = ~N715;
  assign N1833 = ~N720;
  assign N1834 = ~N725;
  assign N1835 = ~N730;
  assign N1836 = ~N735;
  assign N1837 = ~N740;
  assign N1838 = ~N745;
  assign N1839 = ~N750;
  assign N1840 = ~N755;
  assign N1841 = ~N760;
  assign N1842 = ~N765;
  assign N1843 = ~N770;
  assign N1844 = ~N775;
  assign N1845 = ~N780;
  assign N1846 = ~N785;
  assign N1847 = ~N790;
  assign N1848 = ~N795;
  assign N1849 = ~N800;
  assign N1850 = ~N805;
  assign N1851 = ~N810;
  assign N1852 = ~N815;
  assign N1853 = ~N820;
  assign N1854 = ~N825;
  assign N1855 = ~N830;
  assign N1856 = ~N835;
  assign N1857 = ~N840;
  assign N1858 = ~N845;
  assign N1859 = ~N850;
  assign N1860 = ~N855;
  assign N1861 = ~N860;
  assign N1862 = ~N865;
  assign N1863 = ~N870;
  assign N1864 = ~N875;
  assign N1865 = ~N880;
  assign N1866 = ~N885;
  assign N1867 = ~N890;
  assign N1868 = ~N895;
  assign N1869 = ~N900;
  assign N1870 = ~N905;
  assign N1871 = ~N910;
  assign N1872 = ~N915;
  assign N1873 = ~N920;
  assign N1874 = ~N925;
  assign N1875 = ~N930;
  assign N1876 = ~N935;
  assign N1877 = ~N940;
  assign N1878 = ~N945;
  assign N1879 = ~N950;
  assign N1880 = ~N955;
  assign N1881 = ~N960;
  assign N1882 = ~N965;
  assign N1883 = ~N970;
  assign N1884 = ~N975;
  assign N1885 = ~N980;
  assign N1886 = ~N985;
  assign N1887 = ~N990;
  assign N1888 = ~N995;
  assign N1889 = ~N1000;
  assign N1890 = ~N1005;
  assign N1891 = ~N1010;
  assign N1892 = ~N1015;
  assign N1893 = ~N1020;
  assign N1894 = ~N1025;
  assign N1895 = ~N1030;
  assign N1896 = ~N1035;
  assign N1897 = ~N1040;
  assign N1898 = ~N1045;
  assign N1899 = ~N1050;
  assign N1900 = ~N1055;
  assign N1901 = ~N1060;
  assign N1902 = ~N1065;
  assign N1903 = ~N1070;
  assign N1904 = ~N1075;
  assign N1905 = ~N1080;
  assign N1906 = ~N1085;
  assign N1907 = ~N1090;
  assign N1908 = ~N1095;
  assign N1909 = ~N1100;
  assign N1910 = ~N1105;
  assign N1911 = ~N1110;
  assign N1912 = ~N1115;
  assign N1913 = ~N1120;
  assign N1914 = ~N1125;
  assign N1915 = ~N1130;
  assign N1916 = ~N1135;
  assign N1917 = ~N1140;
  assign N1918 = ~N1145;
  assign N1919 = ~N1150;
  assign N1920 = ~N1155;
  assign N1921 = ~N1160;
  assign N1922 = ~N1165;
  assign N1923 = ~N1170;
  assign N1924 = ~N1175;
  assign N1925 = ~N1180;
  assign N1926 = ~N1185;
  assign N1927 = ~N1190;
  assign N1928 = ~N1195;
  assign N1929 = ~N1200;
  assign N1930 = ~N1205;
  assign N1931 = ~N1210;
  assign N1932 = ~N1215;
  assign N1933 = ~N1220;
  assign N1934 = ~N1225;
  assign N1935 = ~N1230;
  assign N1936 = ~N1235;
  assign N1937 = ~N1240;
  assign N1938 = ~N1245;
  assign N1939 = ~N1250;
  assign N1940 = ~N1255;
  assign N1941 = ~N1260;
  assign N1942 = ~N1265;
  assign N1943 = ~N1270;
  assign N1944 = ~N1275;
  assign N1945 = ~N1280;
  assign N1946 = ~N1285;
  assign N1947 = ~N1290;
  assign N1948 = ~N1295;
  assign N1949 = ~N1300;
  assign N1950 = ~N1305;
  assign N1951 = ~N1310;
  assign N1952 = ~N1315;
  assign N1953 = ~N1320;
  assign N1954 = ~N1325;
  assign N1955 = ~N1330;
  assign N1956 = ~N1335;
  assign N1957 = ~N1340;
  assign N1958 = ~N1345;
  assign N1959 = ~N1350;
  assign N1960 = ~N1355;
  assign N1961 = ~N1360;
  assign N1962 = ~N1365;
  assign N1963 = ~N1370;
  assign N1964 = ~N1375;
  assign N1965 = ~N1380;
  assign N1966 = ~N1385;
  assign N1967 = ~N1390;
  assign N1968 = ~N1395;
  assign N1969 = ~N1400;
  assign N1970 = ~N1405;
  assign N1971 = ~N1410;
  assign N1972 = ~N1415;
  assign N1973 = ~N1420;
  assign N1974 = ~N1425;
  assign N1975 = ~N1430;
  assign N1976 = ~N1435;
  assign N1977 = ~N1440;
  assign N1978 = ~N1445;
  assign N1979 = ~N1450;
  assign N1980 = ~N1455;
  assign N1981 = ~N1460;
  assign N1982 = ~N1465;
  assign N1983 = ~N1470;
  assign N1984 = ~N1475;
  assign N1985 = ~N1480;
  assign N1986 = ~N1485;
  assign N1987 = ~N1490;
  assign N1988 = ~N1495;
  assign N1989 = ~N1500;
  assign N1990 = ~N1505;
  assign N1991 = ~N1510;
  assign N1992 = ~N1515;
  assign N1993 = ~N1520;
  assign N1994 = ~N1525;
  assign N1995 = ~N1530;
  assign N1996 = ~N1535;
  assign N1997 = ~N1540;
  assign N1998 = ~N1545;
  assign N1999 = ~N1550;
  assign N2000 = ~N1555;
  assign N2001 = ~N1560;
  assign N2002 = ~N1565;
  assign N2003 = ~N1570;
  assign N2004 = ~N1575;
  assign N2005 = ~N1580;
  assign N2006 = ~N1585;
  assign N2007 = ~N1590;
  assign N2008 = ~N1595;
  assign N2009 = ~N1600;
  assign N2010 = ~N1605;
  assign N2011 = ~N1610;
  assign N2012 = ~N1615;
  assign N2013 = ~N1620;
  assign N2014 = ~N1625;
  assign N2015 = ~N1630;
  assign N2016 = ~N1635;
  assign N2017 = ~N1640;
  assign N2018 = ~N1645;
  assign N2019 = ~N1650;
  assign N2020 = ~N1655;
  assign N2021 = ~N1660;
  assign N2022 = ~N1665;
  assign N2023 = ~N1670;
  assign N2024 = ~N1675;
  assign N2025 = ~N1680;
  assign N2026 = ~N1685;
  assign N2027 = ~N1690;
  assign N2028 = ~N1695;
  assign N2029 = ~N1700;
  assign N2030 = ~N1705;
  assign N2031 = ~N1710;
  assign N2032 = ~N1715;
  assign N2033 = ~N1720;
  assign N2034 = ~N1725;
  assign N2035 = ~N1730;
  assign N2036 = ~N1735;
  assign N2037 = ~N1740;
  assign N2038 = ~N1745;
  assign N2039 = ~N1750;
  assign N2040 = ~N1755;
  assign N2041 = ~N1760;
  assign N2042 = ~N1765;
  assign N2043 = ~N1770;
  assign N2044 = ~N1775;
  assign N2045 = ~N1780;
  assign N2046 = ~N1785;
  assign N2047 = ~N1790;

  always @(posedge clk_i) begin
    if(N1792) begin
      { data_o[31:0] } <= { r_n_0__31_, r_n_0__30_, r_n_0__29_, r_n_0__28_, r_n_0__27_, r_n_0__26_, r_n_0__25_, r_n_0__24_, r_n_0__23_, r_n_0__22_, r_n_0__21_, r_n_0__20_, r_n_0__19_, r_n_0__18_, r_n_0__17_, r_n_0__16_, r_n_0__15_, r_n_0__14_, r_n_0__13_, r_n_0__12_, r_n_0__11_, r_n_0__10_, r_n_0__9_, r_n_0__8_, r_n_0__7_, r_n_0__6_, r_n_0__5_, r_n_0__4_, r_n_0__3_, r_n_0__2_, r_n_0__1_, r_n_0__0_ };
    end 
    if(N1793) begin
      r_1__31_ <= r_n_1__31_;
      r_1__30_ <= r_n_1__30_;
      r_1__29_ <= r_n_1__29_;
      r_1__28_ <= r_n_1__28_;
      r_1__27_ <= r_n_1__27_;
      r_1__26_ <= r_n_1__26_;
      r_1__25_ <= r_n_1__25_;
      r_1__24_ <= r_n_1__24_;
      r_1__23_ <= r_n_1__23_;
      r_1__22_ <= r_n_1__22_;
      r_1__21_ <= r_n_1__21_;
      r_1__20_ <= r_n_1__20_;
      r_1__19_ <= r_n_1__19_;
      r_1__18_ <= r_n_1__18_;
      r_1__17_ <= r_n_1__17_;
      r_1__16_ <= r_n_1__16_;
      r_1__15_ <= r_n_1__15_;
      r_1__14_ <= r_n_1__14_;
      r_1__13_ <= r_n_1__13_;
      r_1__12_ <= r_n_1__12_;
      r_1__11_ <= r_n_1__11_;
      r_1__10_ <= r_n_1__10_;
      r_1__9_ <= r_n_1__9_;
      r_1__8_ <= r_n_1__8_;
      r_1__7_ <= r_n_1__7_;
      r_1__6_ <= r_n_1__6_;
      r_1__5_ <= r_n_1__5_;
      r_1__4_ <= r_n_1__4_;
      r_1__3_ <= r_n_1__3_;
      r_1__2_ <= r_n_1__2_;
      r_1__1_ <= r_n_1__1_;
      r_1__0_ <= r_n_1__0_;
    end 
    if(N1794) begin
      r_2__31_ <= r_n_2__31_;
      r_2__30_ <= r_n_2__30_;
      r_2__29_ <= r_n_2__29_;
      r_2__28_ <= r_n_2__28_;
      r_2__27_ <= r_n_2__27_;
      r_2__26_ <= r_n_2__26_;
      r_2__25_ <= r_n_2__25_;
      r_2__24_ <= r_n_2__24_;
      r_2__23_ <= r_n_2__23_;
      r_2__22_ <= r_n_2__22_;
      r_2__21_ <= r_n_2__21_;
      r_2__20_ <= r_n_2__20_;
      r_2__19_ <= r_n_2__19_;
      r_2__18_ <= r_n_2__18_;
      r_2__17_ <= r_n_2__17_;
      r_2__16_ <= r_n_2__16_;
      r_2__15_ <= r_n_2__15_;
      r_2__14_ <= r_n_2__14_;
      r_2__13_ <= r_n_2__13_;
      r_2__12_ <= r_n_2__12_;
      r_2__11_ <= r_n_2__11_;
      r_2__10_ <= r_n_2__10_;
      r_2__9_ <= r_n_2__9_;
      r_2__8_ <= r_n_2__8_;
      r_2__7_ <= r_n_2__7_;
      r_2__6_ <= r_n_2__6_;
      r_2__5_ <= r_n_2__5_;
      r_2__4_ <= r_n_2__4_;
      r_2__3_ <= r_n_2__3_;
      r_2__2_ <= r_n_2__2_;
      r_2__1_ <= r_n_2__1_;
      r_2__0_ <= r_n_2__0_;
    end 
    if(N1795) begin
      r_3__31_ <= r_n_3__31_;
      r_3__30_ <= r_n_3__30_;
      r_3__29_ <= r_n_3__29_;
      r_3__28_ <= r_n_3__28_;
      r_3__27_ <= r_n_3__27_;
      r_3__26_ <= r_n_3__26_;
      r_3__25_ <= r_n_3__25_;
      r_3__24_ <= r_n_3__24_;
      r_3__23_ <= r_n_3__23_;
      r_3__22_ <= r_n_3__22_;
      r_3__21_ <= r_n_3__21_;
      r_3__20_ <= r_n_3__20_;
      r_3__19_ <= r_n_3__19_;
      r_3__18_ <= r_n_3__18_;
      r_3__17_ <= r_n_3__17_;
      r_3__16_ <= r_n_3__16_;
      r_3__15_ <= r_n_3__15_;
      r_3__14_ <= r_n_3__14_;
      r_3__13_ <= r_n_3__13_;
      r_3__12_ <= r_n_3__12_;
      r_3__11_ <= r_n_3__11_;
      r_3__10_ <= r_n_3__10_;
      r_3__9_ <= r_n_3__9_;
      r_3__8_ <= r_n_3__8_;
      r_3__7_ <= r_n_3__7_;
      r_3__6_ <= r_n_3__6_;
      r_3__5_ <= r_n_3__5_;
      r_3__4_ <= r_n_3__4_;
      r_3__3_ <= r_n_3__3_;
      r_3__2_ <= r_n_3__2_;
      r_3__1_ <= r_n_3__1_;
      r_3__0_ <= r_n_3__0_;
    end 
    if(N1796) begin
      r_4__31_ <= r_n_4__31_;
      r_4__30_ <= r_n_4__30_;
      r_4__29_ <= r_n_4__29_;
      r_4__28_ <= r_n_4__28_;
      r_4__27_ <= r_n_4__27_;
      r_4__26_ <= r_n_4__26_;
      r_4__25_ <= r_n_4__25_;
      r_4__24_ <= r_n_4__24_;
      r_4__23_ <= r_n_4__23_;
      r_4__22_ <= r_n_4__22_;
      r_4__21_ <= r_n_4__21_;
      r_4__20_ <= r_n_4__20_;
      r_4__19_ <= r_n_4__19_;
      r_4__18_ <= r_n_4__18_;
      r_4__17_ <= r_n_4__17_;
      r_4__16_ <= r_n_4__16_;
      r_4__15_ <= r_n_4__15_;
      r_4__14_ <= r_n_4__14_;
      r_4__13_ <= r_n_4__13_;
      r_4__12_ <= r_n_4__12_;
      r_4__11_ <= r_n_4__11_;
      r_4__10_ <= r_n_4__10_;
      r_4__9_ <= r_n_4__9_;
      r_4__8_ <= r_n_4__8_;
      r_4__7_ <= r_n_4__7_;
      r_4__6_ <= r_n_4__6_;
      r_4__5_ <= r_n_4__5_;
      r_4__4_ <= r_n_4__4_;
      r_4__3_ <= r_n_4__3_;
      r_4__2_ <= r_n_4__2_;
      r_4__1_ <= r_n_4__1_;
      r_4__0_ <= r_n_4__0_;
    end 
    if(N1797) begin
      r_5__31_ <= r_n_5__31_;
      r_5__30_ <= r_n_5__30_;
      r_5__29_ <= r_n_5__29_;
      r_5__28_ <= r_n_5__28_;
      r_5__27_ <= r_n_5__27_;
      r_5__26_ <= r_n_5__26_;
      r_5__25_ <= r_n_5__25_;
      r_5__24_ <= r_n_5__24_;
      r_5__23_ <= r_n_5__23_;
      r_5__22_ <= r_n_5__22_;
      r_5__21_ <= r_n_5__21_;
      r_5__20_ <= r_n_5__20_;
      r_5__19_ <= r_n_5__19_;
      r_5__18_ <= r_n_5__18_;
      r_5__17_ <= r_n_5__17_;
      r_5__16_ <= r_n_5__16_;
      r_5__15_ <= r_n_5__15_;
      r_5__14_ <= r_n_5__14_;
      r_5__13_ <= r_n_5__13_;
      r_5__12_ <= r_n_5__12_;
      r_5__11_ <= r_n_5__11_;
      r_5__10_ <= r_n_5__10_;
      r_5__9_ <= r_n_5__9_;
      r_5__8_ <= r_n_5__8_;
      r_5__7_ <= r_n_5__7_;
      r_5__6_ <= r_n_5__6_;
      r_5__5_ <= r_n_5__5_;
      r_5__4_ <= r_n_5__4_;
      r_5__3_ <= r_n_5__3_;
      r_5__2_ <= r_n_5__2_;
      r_5__1_ <= r_n_5__1_;
      r_5__0_ <= r_n_5__0_;
    end 
    if(N1798) begin
      r_6__31_ <= r_n_6__31_;
      r_6__30_ <= r_n_6__30_;
      r_6__29_ <= r_n_6__29_;
      r_6__28_ <= r_n_6__28_;
      r_6__27_ <= r_n_6__27_;
      r_6__26_ <= r_n_6__26_;
      r_6__25_ <= r_n_6__25_;
      r_6__24_ <= r_n_6__24_;
      r_6__23_ <= r_n_6__23_;
      r_6__22_ <= r_n_6__22_;
      r_6__21_ <= r_n_6__21_;
      r_6__20_ <= r_n_6__20_;
      r_6__19_ <= r_n_6__19_;
      r_6__18_ <= r_n_6__18_;
      r_6__17_ <= r_n_6__17_;
      r_6__16_ <= r_n_6__16_;
      r_6__15_ <= r_n_6__15_;
      r_6__14_ <= r_n_6__14_;
      r_6__13_ <= r_n_6__13_;
      r_6__12_ <= r_n_6__12_;
      r_6__11_ <= r_n_6__11_;
      r_6__10_ <= r_n_6__10_;
      r_6__9_ <= r_n_6__9_;
      r_6__8_ <= r_n_6__8_;
      r_6__7_ <= r_n_6__7_;
      r_6__6_ <= r_n_6__6_;
      r_6__5_ <= r_n_6__5_;
      r_6__4_ <= r_n_6__4_;
      r_6__3_ <= r_n_6__3_;
      r_6__2_ <= r_n_6__2_;
      r_6__1_ <= r_n_6__1_;
      r_6__0_ <= r_n_6__0_;
    end 
    if(N1799) begin
      r_7__31_ <= r_n_7__31_;
      r_7__30_ <= r_n_7__30_;
      r_7__29_ <= r_n_7__29_;
      r_7__28_ <= r_n_7__28_;
      r_7__27_ <= r_n_7__27_;
      r_7__26_ <= r_n_7__26_;
      r_7__25_ <= r_n_7__25_;
      r_7__24_ <= r_n_7__24_;
      r_7__23_ <= r_n_7__23_;
      r_7__22_ <= r_n_7__22_;
      r_7__21_ <= r_n_7__21_;
      r_7__20_ <= r_n_7__20_;
      r_7__19_ <= r_n_7__19_;
      r_7__18_ <= r_n_7__18_;
      r_7__17_ <= r_n_7__17_;
      r_7__16_ <= r_n_7__16_;
      r_7__15_ <= r_n_7__15_;
      r_7__14_ <= r_n_7__14_;
      r_7__13_ <= r_n_7__13_;
      r_7__12_ <= r_n_7__12_;
      r_7__11_ <= r_n_7__11_;
      r_7__10_ <= r_n_7__10_;
      r_7__9_ <= r_n_7__9_;
      r_7__8_ <= r_n_7__8_;
      r_7__7_ <= r_n_7__7_;
      r_7__6_ <= r_n_7__6_;
      r_7__5_ <= r_n_7__5_;
      r_7__4_ <= r_n_7__4_;
      r_7__3_ <= r_n_7__3_;
      r_7__2_ <= r_n_7__2_;
      r_7__1_ <= r_n_7__1_;
      r_7__0_ <= r_n_7__0_;
    end 
    if(N1800) begin
      r_8__31_ <= r_n_8__31_;
      r_8__30_ <= r_n_8__30_;
      r_8__29_ <= r_n_8__29_;
      r_8__28_ <= r_n_8__28_;
      r_8__27_ <= r_n_8__27_;
      r_8__26_ <= r_n_8__26_;
      r_8__25_ <= r_n_8__25_;
      r_8__24_ <= r_n_8__24_;
      r_8__23_ <= r_n_8__23_;
      r_8__22_ <= r_n_8__22_;
      r_8__21_ <= r_n_8__21_;
      r_8__20_ <= r_n_8__20_;
      r_8__19_ <= r_n_8__19_;
      r_8__18_ <= r_n_8__18_;
      r_8__17_ <= r_n_8__17_;
      r_8__16_ <= r_n_8__16_;
      r_8__15_ <= r_n_8__15_;
      r_8__14_ <= r_n_8__14_;
      r_8__13_ <= r_n_8__13_;
      r_8__12_ <= r_n_8__12_;
      r_8__11_ <= r_n_8__11_;
      r_8__10_ <= r_n_8__10_;
      r_8__9_ <= r_n_8__9_;
      r_8__8_ <= r_n_8__8_;
      r_8__7_ <= r_n_8__7_;
      r_8__6_ <= r_n_8__6_;
      r_8__5_ <= r_n_8__5_;
      r_8__4_ <= r_n_8__4_;
      r_8__3_ <= r_n_8__3_;
      r_8__2_ <= r_n_8__2_;
      r_8__1_ <= r_n_8__1_;
      r_8__0_ <= r_n_8__0_;
    end 
    if(N1801) begin
      r_9__31_ <= r_n_9__31_;
      r_9__30_ <= r_n_9__30_;
      r_9__29_ <= r_n_9__29_;
      r_9__28_ <= r_n_9__28_;
      r_9__27_ <= r_n_9__27_;
      r_9__26_ <= r_n_9__26_;
      r_9__25_ <= r_n_9__25_;
      r_9__24_ <= r_n_9__24_;
      r_9__23_ <= r_n_9__23_;
      r_9__22_ <= r_n_9__22_;
      r_9__21_ <= r_n_9__21_;
      r_9__20_ <= r_n_9__20_;
      r_9__19_ <= r_n_9__19_;
      r_9__18_ <= r_n_9__18_;
      r_9__17_ <= r_n_9__17_;
      r_9__16_ <= r_n_9__16_;
      r_9__15_ <= r_n_9__15_;
      r_9__14_ <= r_n_9__14_;
      r_9__13_ <= r_n_9__13_;
      r_9__12_ <= r_n_9__12_;
      r_9__11_ <= r_n_9__11_;
      r_9__10_ <= r_n_9__10_;
      r_9__9_ <= r_n_9__9_;
      r_9__8_ <= r_n_9__8_;
      r_9__7_ <= r_n_9__7_;
      r_9__6_ <= r_n_9__6_;
      r_9__5_ <= r_n_9__5_;
      r_9__4_ <= r_n_9__4_;
      r_9__3_ <= r_n_9__3_;
      r_9__2_ <= r_n_9__2_;
      r_9__1_ <= r_n_9__1_;
      r_9__0_ <= r_n_9__0_;
    end 
    if(N1802) begin
      r_10__31_ <= r_n_10__31_;
      r_10__30_ <= r_n_10__30_;
      r_10__29_ <= r_n_10__29_;
      r_10__28_ <= r_n_10__28_;
      r_10__27_ <= r_n_10__27_;
      r_10__26_ <= r_n_10__26_;
      r_10__25_ <= r_n_10__25_;
      r_10__24_ <= r_n_10__24_;
      r_10__23_ <= r_n_10__23_;
      r_10__22_ <= r_n_10__22_;
      r_10__21_ <= r_n_10__21_;
      r_10__20_ <= r_n_10__20_;
      r_10__19_ <= r_n_10__19_;
      r_10__18_ <= r_n_10__18_;
      r_10__17_ <= r_n_10__17_;
      r_10__16_ <= r_n_10__16_;
      r_10__15_ <= r_n_10__15_;
      r_10__14_ <= r_n_10__14_;
      r_10__13_ <= r_n_10__13_;
      r_10__12_ <= r_n_10__12_;
      r_10__11_ <= r_n_10__11_;
      r_10__10_ <= r_n_10__10_;
      r_10__9_ <= r_n_10__9_;
      r_10__8_ <= r_n_10__8_;
      r_10__7_ <= r_n_10__7_;
      r_10__6_ <= r_n_10__6_;
      r_10__5_ <= r_n_10__5_;
      r_10__4_ <= r_n_10__4_;
      r_10__3_ <= r_n_10__3_;
      r_10__2_ <= r_n_10__2_;
      r_10__1_ <= r_n_10__1_;
      r_10__0_ <= r_n_10__0_;
    end 
    if(N1803) begin
      r_11__31_ <= r_n_11__31_;
      r_11__30_ <= r_n_11__30_;
      r_11__29_ <= r_n_11__29_;
      r_11__28_ <= r_n_11__28_;
      r_11__27_ <= r_n_11__27_;
      r_11__26_ <= r_n_11__26_;
      r_11__25_ <= r_n_11__25_;
      r_11__24_ <= r_n_11__24_;
      r_11__23_ <= r_n_11__23_;
      r_11__22_ <= r_n_11__22_;
      r_11__21_ <= r_n_11__21_;
      r_11__20_ <= r_n_11__20_;
      r_11__19_ <= r_n_11__19_;
      r_11__18_ <= r_n_11__18_;
      r_11__17_ <= r_n_11__17_;
      r_11__16_ <= r_n_11__16_;
      r_11__15_ <= r_n_11__15_;
      r_11__14_ <= r_n_11__14_;
      r_11__13_ <= r_n_11__13_;
      r_11__12_ <= r_n_11__12_;
      r_11__11_ <= r_n_11__11_;
      r_11__10_ <= r_n_11__10_;
      r_11__9_ <= r_n_11__9_;
      r_11__8_ <= r_n_11__8_;
      r_11__7_ <= r_n_11__7_;
      r_11__6_ <= r_n_11__6_;
      r_11__5_ <= r_n_11__5_;
      r_11__4_ <= r_n_11__4_;
      r_11__3_ <= r_n_11__3_;
      r_11__2_ <= r_n_11__2_;
      r_11__1_ <= r_n_11__1_;
      r_11__0_ <= r_n_11__0_;
    end 
    if(N1804) begin
      r_12__31_ <= r_n_12__31_;
      r_12__30_ <= r_n_12__30_;
      r_12__29_ <= r_n_12__29_;
      r_12__28_ <= r_n_12__28_;
      r_12__27_ <= r_n_12__27_;
      r_12__26_ <= r_n_12__26_;
      r_12__25_ <= r_n_12__25_;
      r_12__24_ <= r_n_12__24_;
      r_12__23_ <= r_n_12__23_;
      r_12__22_ <= r_n_12__22_;
      r_12__21_ <= r_n_12__21_;
      r_12__20_ <= r_n_12__20_;
      r_12__19_ <= r_n_12__19_;
      r_12__18_ <= r_n_12__18_;
      r_12__17_ <= r_n_12__17_;
      r_12__16_ <= r_n_12__16_;
      r_12__15_ <= r_n_12__15_;
      r_12__14_ <= r_n_12__14_;
      r_12__13_ <= r_n_12__13_;
      r_12__12_ <= r_n_12__12_;
      r_12__11_ <= r_n_12__11_;
      r_12__10_ <= r_n_12__10_;
      r_12__9_ <= r_n_12__9_;
      r_12__8_ <= r_n_12__8_;
      r_12__7_ <= r_n_12__7_;
      r_12__6_ <= r_n_12__6_;
      r_12__5_ <= r_n_12__5_;
      r_12__4_ <= r_n_12__4_;
      r_12__3_ <= r_n_12__3_;
      r_12__2_ <= r_n_12__2_;
      r_12__1_ <= r_n_12__1_;
      r_12__0_ <= r_n_12__0_;
    end 
    if(N1805) begin
      r_13__31_ <= r_n_13__31_;
      r_13__30_ <= r_n_13__30_;
      r_13__29_ <= r_n_13__29_;
      r_13__28_ <= r_n_13__28_;
      r_13__27_ <= r_n_13__27_;
      r_13__26_ <= r_n_13__26_;
      r_13__25_ <= r_n_13__25_;
      r_13__24_ <= r_n_13__24_;
      r_13__23_ <= r_n_13__23_;
      r_13__22_ <= r_n_13__22_;
      r_13__21_ <= r_n_13__21_;
      r_13__20_ <= r_n_13__20_;
      r_13__19_ <= r_n_13__19_;
      r_13__18_ <= r_n_13__18_;
      r_13__17_ <= r_n_13__17_;
      r_13__16_ <= r_n_13__16_;
      r_13__15_ <= r_n_13__15_;
      r_13__14_ <= r_n_13__14_;
      r_13__13_ <= r_n_13__13_;
      r_13__12_ <= r_n_13__12_;
      r_13__11_ <= r_n_13__11_;
      r_13__10_ <= r_n_13__10_;
      r_13__9_ <= r_n_13__9_;
      r_13__8_ <= r_n_13__8_;
      r_13__7_ <= r_n_13__7_;
      r_13__6_ <= r_n_13__6_;
      r_13__5_ <= r_n_13__5_;
      r_13__4_ <= r_n_13__4_;
      r_13__3_ <= r_n_13__3_;
      r_13__2_ <= r_n_13__2_;
      r_13__1_ <= r_n_13__1_;
      r_13__0_ <= r_n_13__0_;
    end 
    if(N1806) begin
      r_14__31_ <= r_n_14__31_;
      r_14__30_ <= r_n_14__30_;
      r_14__29_ <= r_n_14__29_;
      r_14__28_ <= r_n_14__28_;
      r_14__27_ <= r_n_14__27_;
      r_14__26_ <= r_n_14__26_;
      r_14__25_ <= r_n_14__25_;
      r_14__24_ <= r_n_14__24_;
      r_14__23_ <= r_n_14__23_;
      r_14__22_ <= r_n_14__22_;
      r_14__21_ <= r_n_14__21_;
      r_14__20_ <= r_n_14__20_;
      r_14__19_ <= r_n_14__19_;
      r_14__18_ <= r_n_14__18_;
      r_14__17_ <= r_n_14__17_;
      r_14__16_ <= r_n_14__16_;
      r_14__15_ <= r_n_14__15_;
      r_14__14_ <= r_n_14__14_;
      r_14__13_ <= r_n_14__13_;
      r_14__12_ <= r_n_14__12_;
      r_14__11_ <= r_n_14__11_;
      r_14__10_ <= r_n_14__10_;
      r_14__9_ <= r_n_14__9_;
      r_14__8_ <= r_n_14__8_;
      r_14__7_ <= r_n_14__7_;
      r_14__6_ <= r_n_14__6_;
      r_14__5_ <= r_n_14__5_;
      r_14__4_ <= r_n_14__4_;
      r_14__3_ <= r_n_14__3_;
      r_14__2_ <= r_n_14__2_;
      r_14__1_ <= r_n_14__1_;
      r_14__0_ <= r_n_14__0_;
    end 
    if(N1807) begin
      r_15__31_ <= r_n_15__31_;
      r_15__30_ <= r_n_15__30_;
      r_15__29_ <= r_n_15__29_;
      r_15__28_ <= r_n_15__28_;
      r_15__27_ <= r_n_15__27_;
      r_15__26_ <= r_n_15__26_;
      r_15__25_ <= r_n_15__25_;
      r_15__24_ <= r_n_15__24_;
      r_15__23_ <= r_n_15__23_;
      r_15__22_ <= r_n_15__22_;
      r_15__21_ <= r_n_15__21_;
      r_15__20_ <= r_n_15__20_;
      r_15__19_ <= r_n_15__19_;
      r_15__18_ <= r_n_15__18_;
      r_15__17_ <= r_n_15__17_;
      r_15__16_ <= r_n_15__16_;
      r_15__15_ <= r_n_15__15_;
      r_15__14_ <= r_n_15__14_;
      r_15__13_ <= r_n_15__13_;
      r_15__12_ <= r_n_15__12_;
      r_15__11_ <= r_n_15__11_;
      r_15__10_ <= r_n_15__10_;
      r_15__9_ <= r_n_15__9_;
      r_15__8_ <= r_n_15__8_;
      r_15__7_ <= r_n_15__7_;
      r_15__6_ <= r_n_15__6_;
      r_15__5_ <= r_n_15__5_;
      r_15__4_ <= r_n_15__4_;
      r_15__3_ <= r_n_15__3_;
      r_15__2_ <= r_n_15__2_;
      r_15__1_ <= r_n_15__1_;
      r_15__0_ <= r_n_15__0_;
    end 
    if(N1808) begin
      r_16__31_ <= r_n_16__31_;
      r_16__30_ <= r_n_16__30_;
      r_16__29_ <= r_n_16__29_;
      r_16__28_ <= r_n_16__28_;
      r_16__27_ <= r_n_16__27_;
      r_16__26_ <= r_n_16__26_;
      r_16__25_ <= r_n_16__25_;
      r_16__24_ <= r_n_16__24_;
      r_16__23_ <= r_n_16__23_;
      r_16__22_ <= r_n_16__22_;
      r_16__21_ <= r_n_16__21_;
      r_16__20_ <= r_n_16__20_;
      r_16__19_ <= r_n_16__19_;
      r_16__18_ <= r_n_16__18_;
      r_16__17_ <= r_n_16__17_;
      r_16__16_ <= r_n_16__16_;
      r_16__15_ <= r_n_16__15_;
      r_16__14_ <= r_n_16__14_;
      r_16__13_ <= r_n_16__13_;
      r_16__12_ <= r_n_16__12_;
      r_16__11_ <= r_n_16__11_;
      r_16__10_ <= r_n_16__10_;
      r_16__9_ <= r_n_16__9_;
      r_16__8_ <= r_n_16__8_;
      r_16__7_ <= r_n_16__7_;
      r_16__6_ <= r_n_16__6_;
      r_16__5_ <= r_n_16__5_;
      r_16__4_ <= r_n_16__4_;
      r_16__3_ <= r_n_16__3_;
      r_16__2_ <= r_n_16__2_;
      r_16__1_ <= r_n_16__1_;
      r_16__0_ <= r_n_16__0_;
    end 
    if(N1809) begin
      r_17__31_ <= r_n_17__31_;
      r_17__30_ <= r_n_17__30_;
      r_17__29_ <= r_n_17__29_;
      r_17__28_ <= r_n_17__28_;
      r_17__27_ <= r_n_17__27_;
      r_17__26_ <= r_n_17__26_;
      r_17__25_ <= r_n_17__25_;
      r_17__24_ <= r_n_17__24_;
      r_17__23_ <= r_n_17__23_;
      r_17__22_ <= r_n_17__22_;
      r_17__21_ <= r_n_17__21_;
      r_17__20_ <= r_n_17__20_;
      r_17__19_ <= r_n_17__19_;
      r_17__18_ <= r_n_17__18_;
      r_17__17_ <= r_n_17__17_;
      r_17__16_ <= r_n_17__16_;
      r_17__15_ <= r_n_17__15_;
      r_17__14_ <= r_n_17__14_;
      r_17__13_ <= r_n_17__13_;
      r_17__12_ <= r_n_17__12_;
      r_17__11_ <= r_n_17__11_;
      r_17__10_ <= r_n_17__10_;
      r_17__9_ <= r_n_17__9_;
      r_17__8_ <= r_n_17__8_;
      r_17__7_ <= r_n_17__7_;
      r_17__6_ <= r_n_17__6_;
      r_17__5_ <= r_n_17__5_;
      r_17__4_ <= r_n_17__4_;
      r_17__3_ <= r_n_17__3_;
      r_17__2_ <= r_n_17__2_;
      r_17__1_ <= r_n_17__1_;
      r_17__0_ <= r_n_17__0_;
    end 
    if(N1810) begin
      r_18__31_ <= r_n_18__31_;
      r_18__30_ <= r_n_18__30_;
      r_18__29_ <= r_n_18__29_;
      r_18__28_ <= r_n_18__28_;
      r_18__27_ <= r_n_18__27_;
      r_18__26_ <= r_n_18__26_;
      r_18__25_ <= r_n_18__25_;
      r_18__24_ <= r_n_18__24_;
      r_18__23_ <= r_n_18__23_;
      r_18__22_ <= r_n_18__22_;
      r_18__21_ <= r_n_18__21_;
      r_18__20_ <= r_n_18__20_;
      r_18__19_ <= r_n_18__19_;
      r_18__18_ <= r_n_18__18_;
      r_18__17_ <= r_n_18__17_;
      r_18__16_ <= r_n_18__16_;
      r_18__15_ <= r_n_18__15_;
      r_18__14_ <= r_n_18__14_;
      r_18__13_ <= r_n_18__13_;
      r_18__12_ <= r_n_18__12_;
      r_18__11_ <= r_n_18__11_;
      r_18__10_ <= r_n_18__10_;
      r_18__9_ <= r_n_18__9_;
      r_18__8_ <= r_n_18__8_;
      r_18__7_ <= r_n_18__7_;
      r_18__6_ <= r_n_18__6_;
      r_18__5_ <= r_n_18__5_;
      r_18__4_ <= r_n_18__4_;
      r_18__3_ <= r_n_18__3_;
      r_18__2_ <= r_n_18__2_;
      r_18__1_ <= r_n_18__1_;
      r_18__0_ <= r_n_18__0_;
    end 
    if(N1811) begin
      r_19__31_ <= r_n_19__31_;
      r_19__30_ <= r_n_19__30_;
      r_19__29_ <= r_n_19__29_;
      r_19__28_ <= r_n_19__28_;
      r_19__27_ <= r_n_19__27_;
      r_19__26_ <= r_n_19__26_;
      r_19__25_ <= r_n_19__25_;
      r_19__24_ <= r_n_19__24_;
      r_19__23_ <= r_n_19__23_;
      r_19__22_ <= r_n_19__22_;
      r_19__21_ <= r_n_19__21_;
      r_19__20_ <= r_n_19__20_;
      r_19__19_ <= r_n_19__19_;
      r_19__18_ <= r_n_19__18_;
      r_19__17_ <= r_n_19__17_;
      r_19__16_ <= r_n_19__16_;
      r_19__15_ <= r_n_19__15_;
      r_19__14_ <= r_n_19__14_;
      r_19__13_ <= r_n_19__13_;
      r_19__12_ <= r_n_19__12_;
      r_19__11_ <= r_n_19__11_;
      r_19__10_ <= r_n_19__10_;
      r_19__9_ <= r_n_19__9_;
      r_19__8_ <= r_n_19__8_;
      r_19__7_ <= r_n_19__7_;
      r_19__6_ <= r_n_19__6_;
      r_19__5_ <= r_n_19__5_;
      r_19__4_ <= r_n_19__4_;
      r_19__3_ <= r_n_19__3_;
      r_19__2_ <= r_n_19__2_;
      r_19__1_ <= r_n_19__1_;
      r_19__0_ <= r_n_19__0_;
    end 
    if(N1812) begin
      r_20__31_ <= r_n_20__31_;
      r_20__30_ <= r_n_20__30_;
      r_20__29_ <= r_n_20__29_;
      r_20__28_ <= r_n_20__28_;
      r_20__27_ <= r_n_20__27_;
      r_20__26_ <= r_n_20__26_;
      r_20__25_ <= r_n_20__25_;
      r_20__24_ <= r_n_20__24_;
      r_20__23_ <= r_n_20__23_;
      r_20__22_ <= r_n_20__22_;
      r_20__21_ <= r_n_20__21_;
      r_20__20_ <= r_n_20__20_;
      r_20__19_ <= r_n_20__19_;
      r_20__18_ <= r_n_20__18_;
      r_20__17_ <= r_n_20__17_;
      r_20__16_ <= r_n_20__16_;
      r_20__15_ <= r_n_20__15_;
      r_20__14_ <= r_n_20__14_;
      r_20__13_ <= r_n_20__13_;
      r_20__12_ <= r_n_20__12_;
      r_20__11_ <= r_n_20__11_;
      r_20__10_ <= r_n_20__10_;
      r_20__9_ <= r_n_20__9_;
      r_20__8_ <= r_n_20__8_;
      r_20__7_ <= r_n_20__7_;
      r_20__6_ <= r_n_20__6_;
      r_20__5_ <= r_n_20__5_;
      r_20__4_ <= r_n_20__4_;
      r_20__3_ <= r_n_20__3_;
      r_20__2_ <= r_n_20__2_;
      r_20__1_ <= r_n_20__1_;
      r_20__0_ <= r_n_20__0_;
    end 
    if(N1813) begin
      r_21__31_ <= r_n_21__31_;
      r_21__30_ <= r_n_21__30_;
      r_21__29_ <= r_n_21__29_;
      r_21__28_ <= r_n_21__28_;
      r_21__27_ <= r_n_21__27_;
      r_21__26_ <= r_n_21__26_;
      r_21__25_ <= r_n_21__25_;
      r_21__24_ <= r_n_21__24_;
      r_21__23_ <= r_n_21__23_;
      r_21__22_ <= r_n_21__22_;
      r_21__21_ <= r_n_21__21_;
      r_21__20_ <= r_n_21__20_;
      r_21__19_ <= r_n_21__19_;
      r_21__18_ <= r_n_21__18_;
      r_21__17_ <= r_n_21__17_;
      r_21__16_ <= r_n_21__16_;
      r_21__15_ <= r_n_21__15_;
      r_21__14_ <= r_n_21__14_;
      r_21__13_ <= r_n_21__13_;
      r_21__12_ <= r_n_21__12_;
      r_21__11_ <= r_n_21__11_;
      r_21__10_ <= r_n_21__10_;
      r_21__9_ <= r_n_21__9_;
      r_21__8_ <= r_n_21__8_;
      r_21__7_ <= r_n_21__7_;
      r_21__6_ <= r_n_21__6_;
      r_21__5_ <= r_n_21__5_;
      r_21__4_ <= r_n_21__4_;
      r_21__3_ <= r_n_21__3_;
      r_21__2_ <= r_n_21__2_;
      r_21__1_ <= r_n_21__1_;
      r_21__0_ <= r_n_21__0_;
    end 
    if(N1814) begin
      r_22__31_ <= r_n_22__31_;
      r_22__30_ <= r_n_22__30_;
      r_22__29_ <= r_n_22__29_;
      r_22__28_ <= r_n_22__28_;
      r_22__27_ <= r_n_22__27_;
      r_22__26_ <= r_n_22__26_;
      r_22__25_ <= r_n_22__25_;
      r_22__24_ <= r_n_22__24_;
      r_22__23_ <= r_n_22__23_;
      r_22__22_ <= r_n_22__22_;
      r_22__21_ <= r_n_22__21_;
      r_22__20_ <= r_n_22__20_;
      r_22__19_ <= r_n_22__19_;
      r_22__18_ <= r_n_22__18_;
      r_22__17_ <= r_n_22__17_;
      r_22__16_ <= r_n_22__16_;
      r_22__15_ <= r_n_22__15_;
      r_22__14_ <= r_n_22__14_;
      r_22__13_ <= r_n_22__13_;
      r_22__12_ <= r_n_22__12_;
      r_22__11_ <= r_n_22__11_;
      r_22__10_ <= r_n_22__10_;
      r_22__9_ <= r_n_22__9_;
      r_22__8_ <= r_n_22__8_;
      r_22__7_ <= r_n_22__7_;
      r_22__6_ <= r_n_22__6_;
      r_22__5_ <= r_n_22__5_;
      r_22__4_ <= r_n_22__4_;
      r_22__3_ <= r_n_22__3_;
      r_22__2_ <= r_n_22__2_;
      r_22__1_ <= r_n_22__1_;
      r_22__0_ <= r_n_22__0_;
    end 
    if(N1815) begin
      r_23__31_ <= r_n_23__31_;
      r_23__30_ <= r_n_23__30_;
      r_23__29_ <= r_n_23__29_;
      r_23__28_ <= r_n_23__28_;
      r_23__27_ <= r_n_23__27_;
      r_23__26_ <= r_n_23__26_;
      r_23__25_ <= r_n_23__25_;
      r_23__24_ <= r_n_23__24_;
      r_23__23_ <= r_n_23__23_;
      r_23__22_ <= r_n_23__22_;
      r_23__21_ <= r_n_23__21_;
      r_23__20_ <= r_n_23__20_;
      r_23__19_ <= r_n_23__19_;
      r_23__18_ <= r_n_23__18_;
      r_23__17_ <= r_n_23__17_;
      r_23__16_ <= r_n_23__16_;
      r_23__15_ <= r_n_23__15_;
      r_23__14_ <= r_n_23__14_;
      r_23__13_ <= r_n_23__13_;
      r_23__12_ <= r_n_23__12_;
      r_23__11_ <= r_n_23__11_;
      r_23__10_ <= r_n_23__10_;
      r_23__9_ <= r_n_23__9_;
      r_23__8_ <= r_n_23__8_;
      r_23__7_ <= r_n_23__7_;
      r_23__6_ <= r_n_23__6_;
      r_23__5_ <= r_n_23__5_;
      r_23__4_ <= r_n_23__4_;
      r_23__3_ <= r_n_23__3_;
      r_23__2_ <= r_n_23__2_;
      r_23__1_ <= r_n_23__1_;
      r_23__0_ <= r_n_23__0_;
    end 
    if(N1816) begin
      r_24__31_ <= r_n_24__31_;
      r_24__30_ <= r_n_24__30_;
      r_24__29_ <= r_n_24__29_;
      r_24__28_ <= r_n_24__28_;
      r_24__27_ <= r_n_24__27_;
      r_24__26_ <= r_n_24__26_;
      r_24__25_ <= r_n_24__25_;
      r_24__24_ <= r_n_24__24_;
      r_24__23_ <= r_n_24__23_;
      r_24__22_ <= r_n_24__22_;
      r_24__21_ <= r_n_24__21_;
      r_24__20_ <= r_n_24__20_;
      r_24__19_ <= r_n_24__19_;
      r_24__18_ <= r_n_24__18_;
      r_24__17_ <= r_n_24__17_;
      r_24__16_ <= r_n_24__16_;
      r_24__15_ <= r_n_24__15_;
      r_24__14_ <= r_n_24__14_;
      r_24__13_ <= r_n_24__13_;
      r_24__12_ <= r_n_24__12_;
      r_24__11_ <= r_n_24__11_;
      r_24__10_ <= r_n_24__10_;
      r_24__9_ <= r_n_24__9_;
      r_24__8_ <= r_n_24__8_;
      r_24__7_ <= r_n_24__7_;
      r_24__6_ <= r_n_24__6_;
      r_24__5_ <= r_n_24__5_;
      r_24__4_ <= r_n_24__4_;
      r_24__3_ <= r_n_24__3_;
      r_24__2_ <= r_n_24__2_;
      r_24__1_ <= r_n_24__1_;
      r_24__0_ <= r_n_24__0_;
    end 
    if(N1817) begin
      r_25__31_ <= r_n_25__31_;
      r_25__30_ <= r_n_25__30_;
      r_25__29_ <= r_n_25__29_;
      r_25__28_ <= r_n_25__28_;
      r_25__27_ <= r_n_25__27_;
      r_25__26_ <= r_n_25__26_;
      r_25__25_ <= r_n_25__25_;
      r_25__24_ <= r_n_25__24_;
      r_25__23_ <= r_n_25__23_;
      r_25__22_ <= r_n_25__22_;
      r_25__21_ <= r_n_25__21_;
      r_25__20_ <= r_n_25__20_;
      r_25__19_ <= r_n_25__19_;
      r_25__18_ <= r_n_25__18_;
      r_25__17_ <= r_n_25__17_;
      r_25__16_ <= r_n_25__16_;
      r_25__15_ <= r_n_25__15_;
      r_25__14_ <= r_n_25__14_;
      r_25__13_ <= r_n_25__13_;
      r_25__12_ <= r_n_25__12_;
      r_25__11_ <= r_n_25__11_;
      r_25__10_ <= r_n_25__10_;
      r_25__9_ <= r_n_25__9_;
      r_25__8_ <= r_n_25__8_;
      r_25__7_ <= r_n_25__7_;
      r_25__6_ <= r_n_25__6_;
      r_25__5_ <= r_n_25__5_;
      r_25__4_ <= r_n_25__4_;
      r_25__3_ <= r_n_25__3_;
      r_25__2_ <= r_n_25__2_;
      r_25__1_ <= r_n_25__1_;
      r_25__0_ <= r_n_25__0_;
    end 
    if(N1818) begin
      r_26__31_ <= r_n_26__31_;
      r_26__30_ <= r_n_26__30_;
      r_26__29_ <= r_n_26__29_;
      r_26__28_ <= r_n_26__28_;
      r_26__27_ <= r_n_26__27_;
      r_26__26_ <= r_n_26__26_;
      r_26__25_ <= r_n_26__25_;
      r_26__24_ <= r_n_26__24_;
      r_26__23_ <= r_n_26__23_;
      r_26__22_ <= r_n_26__22_;
      r_26__21_ <= r_n_26__21_;
      r_26__20_ <= r_n_26__20_;
      r_26__19_ <= r_n_26__19_;
      r_26__18_ <= r_n_26__18_;
      r_26__17_ <= r_n_26__17_;
      r_26__16_ <= r_n_26__16_;
      r_26__15_ <= r_n_26__15_;
      r_26__14_ <= r_n_26__14_;
      r_26__13_ <= r_n_26__13_;
      r_26__12_ <= r_n_26__12_;
      r_26__11_ <= r_n_26__11_;
      r_26__10_ <= r_n_26__10_;
      r_26__9_ <= r_n_26__9_;
      r_26__8_ <= r_n_26__8_;
      r_26__7_ <= r_n_26__7_;
      r_26__6_ <= r_n_26__6_;
      r_26__5_ <= r_n_26__5_;
      r_26__4_ <= r_n_26__4_;
      r_26__3_ <= r_n_26__3_;
      r_26__2_ <= r_n_26__2_;
      r_26__1_ <= r_n_26__1_;
      r_26__0_ <= r_n_26__0_;
    end 
    if(N1819) begin
      r_27__31_ <= r_n_27__31_;
      r_27__30_ <= r_n_27__30_;
      r_27__29_ <= r_n_27__29_;
      r_27__28_ <= r_n_27__28_;
      r_27__27_ <= r_n_27__27_;
      r_27__26_ <= r_n_27__26_;
      r_27__25_ <= r_n_27__25_;
      r_27__24_ <= r_n_27__24_;
      r_27__23_ <= r_n_27__23_;
      r_27__22_ <= r_n_27__22_;
      r_27__21_ <= r_n_27__21_;
      r_27__20_ <= r_n_27__20_;
      r_27__19_ <= r_n_27__19_;
      r_27__18_ <= r_n_27__18_;
      r_27__17_ <= r_n_27__17_;
      r_27__16_ <= r_n_27__16_;
      r_27__15_ <= r_n_27__15_;
      r_27__14_ <= r_n_27__14_;
      r_27__13_ <= r_n_27__13_;
      r_27__12_ <= r_n_27__12_;
      r_27__11_ <= r_n_27__11_;
      r_27__10_ <= r_n_27__10_;
      r_27__9_ <= r_n_27__9_;
      r_27__8_ <= r_n_27__8_;
      r_27__7_ <= r_n_27__7_;
      r_27__6_ <= r_n_27__6_;
      r_27__5_ <= r_n_27__5_;
      r_27__4_ <= r_n_27__4_;
      r_27__3_ <= r_n_27__3_;
      r_27__2_ <= r_n_27__2_;
      r_27__1_ <= r_n_27__1_;
      r_27__0_ <= r_n_27__0_;
    end 
    if(N1820) begin
      r_28__31_ <= r_n_28__31_;
      r_28__30_ <= r_n_28__30_;
      r_28__29_ <= r_n_28__29_;
      r_28__28_ <= r_n_28__28_;
      r_28__27_ <= r_n_28__27_;
      r_28__26_ <= r_n_28__26_;
      r_28__25_ <= r_n_28__25_;
      r_28__24_ <= r_n_28__24_;
      r_28__23_ <= r_n_28__23_;
      r_28__22_ <= r_n_28__22_;
      r_28__21_ <= r_n_28__21_;
      r_28__20_ <= r_n_28__20_;
      r_28__19_ <= r_n_28__19_;
      r_28__18_ <= r_n_28__18_;
      r_28__17_ <= r_n_28__17_;
      r_28__16_ <= r_n_28__16_;
      r_28__15_ <= r_n_28__15_;
      r_28__14_ <= r_n_28__14_;
      r_28__13_ <= r_n_28__13_;
      r_28__12_ <= r_n_28__12_;
      r_28__11_ <= r_n_28__11_;
      r_28__10_ <= r_n_28__10_;
      r_28__9_ <= r_n_28__9_;
      r_28__8_ <= r_n_28__8_;
      r_28__7_ <= r_n_28__7_;
      r_28__6_ <= r_n_28__6_;
      r_28__5_ <= r_n_28__5_;
      r_28__4_ <= r_n_28__4_;
      r_28__3_ <= r_n_28__3_;
      r_28__2_ <= r_n_28__2_;
      r_28__1_ <= r_n_28__1_;
      r_28__0_ <= r_n_28__0_;
    end 
    if(N1821) begin
      r_29__31_ <= r_n_29__31_;
      r_29__30_ <= r_n_29__30_;
      r_29__29_ <= r_n_29__29_;
      r_29__28_ <= r_n_29__28_;
      r_29__27_ <= r_n_29__27_;
      r_29__26_ <= r_n_29__26_;
      r_29__25_ <= r_n_29__25_;
      r_29__24_ <= r_n_29__24_;
      r_29__23_ <= r_n_29__23_;
      r_29__22_ <= r_n_29__22_;
      r_29__21_ <= r_n_29__21_;
      r_29__20_ <= r_n_29__20_;
      r_29__19_ <= r_n_29__19_;
      r_29__18_ <= r_n_29__18_;
      r_29__17_ <= r_n_29__17_;
      r_29__16_ <= r_n_29__16_;
      r_29__15_ <= r_n_29__15_;
      r_29__14_ <= r_n_29__14_;
      r_29__13_ <= r_n_29__13_;
      r_29__12_ <= r_n_29__12_;
      r_29__11_ <= r_n_29__11_;
      r_29__10_ <= r_n_29__10_;
      r_29__9_ <= r_n_29__9_;
      r_29__8_ <= r_n_29__8_;
      r_29__7_ <= r_n_29__7_;
      r_29__6_ <= r_n_29__6_;
      r_29__5_ <= r_n_29__5_;
      r_29__4_ <= r_n_29__4_;
      r_29__3_ <= r_n_29__3_;
      r_29__2_ <= r_n_29__2_;
      r_29__1_ <= r_n_29__1_;
      r_29__0_ <= r_n_29__0_;
    end 
    if(N1822) begin
      r_30__31_ <= r_n_30__31_;
      r_30__30_ <= r_n_30__30_;
      r_30__29_ <= r_n_30__29_;
      r_30__28_ <= r_n_30__28_;
      r_30__27_ <= r_n_30__27_;
      r_30__26_ <= r_n_30__26_;
      r_30__25_ <= r_n_30__25_;
      r_30__24_ <= r_n_30__24_;
      r_30__23_ <= r_n_30__23_;
      r_30__22_ <= r_n_30__22_;
      r_30__21_ <= r_n_30__21_;
      r_30__20_ <= r_n_30__20_;
      r_30__19_ <= r_n_30__19_;
      r_30__18_ <= r_n_30__18_;
      r_30__17_ <= r_n_30__17_;
      r_30__16_ <= r_n_30__16_;
      r_30__15_ <= r_n_30__15_;
      r_30__14_ <= r_n_30__14_;
      r_30__13_ <= r_n_30__13_;
      r_30__12_ <= r_n_30__12_;
      r_30__11_ <= r_n_30__11_;
      r_30__10_ <= r_n_30__10_;
      r_30__9_ <= r_n_30__9_;
      r_30__8_ <= r_n_30__8_;
      r_30__7_ <= r_n_30__7_;
      r_30__6_ <= r_n_30__6_;
      r_30__5_ <= r_n_30__5_;
      r_30__4_ <= r_n_30__4_;
      r_30__3_ <= r_n_30__3_;
      r_30__2_ <= r_n_30__2_;
      r_30__1_ <= r_n_30__1_;
      r_30__0_ <= r_n_30__0_;
    end 
    if(N1823) begin
      r_31__31_ <= r_n_31__31_;
      r_31__30_ <= r_n_31__30_;
      r_31__29_ <= r_n_31__29_;
      r_31__28_ <= r_n_31__28_;
      r_31__27_ <= r_n_31__27_;
      r_31__26_ <= r_n_31__26_;
      r_31__25_ <= r_n_31__25_;
      r_31__24_ <= r_n_31__24_;
      r_31__23_ <= r_n_31__23_;
      r_31__22_ <= r_n_31__22_;
      r_31__21_ <= r_n_31__21_;
      r_31__20_ <= r_n_31__20_;
      r_31__19_ <= r_n_31__19_;
      r_31__18_ <= r_n_31__18_;
      r_31__17_ <= r_n_31__17_;
      r_31__16_ <= r_n_31__16_;
      r_31__15_ <= r_n_31__15_;
      r_31__14_ <= r_n_31__14_;
      r_31__13_ <= r_n_31__13_;
      r_31__12_ <= r_n_31__12_;
      r_31__11_ <= r_n_31__11_;
      r_31__10_ <= r_n_31__10_;
      r_31__9_ <= r_n_31__9_;
      r_31__8_ <= r_n_31__8_;
      r_31__7_ <= r_n_31__7_;
      r_31__6_ <= r_n_31__6_;
      r_31__5_ <= r_n_31__5_;
      r_31__4_ <= r_n_31__4_;
      r_31__3_ <= r_n_31__3_;
      r_31__2_ <= r_n_31__2_;
      r_31__1_ <= r_n_31__1_;
      r_31__0_ <= r_n_31__0_;
    end 
    if(N1824) begin
      r_32__31_ <= r_n_32__31_;
      r_32__30_ <= r_n_32__30_;
      r_32__29_ <= r_n_32__29_;
      r_32__28_ <= r_n_32__28_;
      r_32__27_ <= r_n_32__27_;
      r_32__26_ <= r_n_32__26_;
      r_32__25_ <= r_n_32__25_;
      r_32__24_ <= r_n_32__24_;
      r_32__23_ <= r_n_32__23_;
      r_32__22_ <= r_n_32__22_;
      r_32__21_ <= r_n_32__21_;
      r_32__20_ <= r_n_32__20_;
      r_32__19_ <= r_n_32__19_;
      r_32__18_ <= r_n_32__18_;
      r_32__17_ <= r_n_32__17_;
      r_32__16_ <= r_n_32__16_;
      r_32__15_ <= r_n_32__15_;
      r_32__14_ <= r_n_32__14_;
      r_32__13_ <= r_n_32__13_;
      r_32__12_ <= r_n_32__12_;
      r_32__11_ <= r_n_32__11_;
      r_32__10_ <= r_n_32__10_;
      r_32__9_ <= r_n_32__9_;
      r_32__8_ <= r_n_32__8_;
      r_32__7_ <= r_n_32__7_;
      r_32__6_ <= r_n_32__6_;
      r_32__5_ <= r_n_32__5_;
      r_32__4_ <= r_n_32__4_;
      r_32__3_ <= r_n_32__3_;
      r_32__2_ <= r_n_32__2_;
      r_32__1_ <= r_n_32__1_;
      r_32__0_ <= r_n_32__0_;
    end 
    if(N1825) begin
      r_33__31_ <= r_n_33__31_;
      r_33__30_ <= r_n_33__30_;
      r_33__29_ <= r_n_33__29_;
      r_33__28_ <= r_n_33__28_;
      r_33__27_ <= r_n_33__27_;
      r_33__26_ <= r_n_33__26_;
      r_33__25_ <= r_n_33__25_;
      r_33__24_ <= r_n_33__24_;
      r_33__23_ <= r_n_33__23_;
      r_33__22_ <= r_n_33__22_;
      r_33__21_ <= r_n_33__21_;
      r_33__20_ <= r_n_33__20_;
      r_33__19_ <= r_n_33__19_;
      r_33__18_ <= r_n_33__18_;
      r_33__17_ <= r_n_33__17_;
      r_33__16_ <= r_n_33__16_;
      r_33__15_ <= r_n_33__15_;
      r_33__14_ <= r_n_33__14_;
      r_33__13_ <= r_n_33__13_;
      r_33__12_ <= r_n_33__12_;
      r_33__11_ <= r_n_33__11_;
      r_33__10_ <= r_n_33__10_;
      r_33__9_ <= r_n_33__9_;
      r_33__8_ <= r_n_33__8_;
      r_33__7_ <= r_n_33__7_;
      r_33__6_ <= r_n_33__6_;
      r_33__5_ <= r_n_33__5_;
      r_33__4_ <= r_n_33__4_;
      r_33__3_ <= r_n_33__3_;
      r_33__2_ <= r_n_33__2_;
      r_33__1_ <= r_n_33__1_;
      r_33__0_ <= r_n_33__0_;
    end 
    if(N1826) begin
      r_34__31_ <= r_n_34__31_;
      r_34__30_ <= r_n_34__30_;
      r_34__29_ <= r_n_34__29_;
      r_34__28_ <= r_n_34__28_;
      r_34__27_ <= r_n_34__27_;
      r_34__26_ <= r_n_34__26_;
      r_34__25_ <= r_n_34__25_;
      r_34__24_ <= r_n_34__24_;
      r_34__23_ <= r_n_34__23_;
      r_34__22_ <= r_n_34__22_;
      r_34__21_ <= r_n_34__21_;
      r_34__20_ <= r_n_34__20_;
      r_34__19_ <= r_n_34__19_;
      r_34__18_ <= r_n_34__18_;
      r_34__17_ <= r_n_34__17_;
      r_34__16_ <= r_n_34__16_;
      r_34__15_ <= r_n_34__15_;
      r_34__14_ <= r_n_34__14_;
      r_34__13_ <= r_n_34__13_;
      r_34__12_ <= r_n_34__12_;
      r_34__11_ <= r_n_34__11_;
      r_34__10_ <= r_n_34__10_;
      r_34__9_ <= r_n_34__9_;
      r_34__8_ <= r_n_34__8_;
      r_34__7_ <= r_n_34__7_;
      r_34__6_ <= r_n_34__6_;
      r_34__5_ <= r_n_34__5_;
      r_34__4_ <= r_n_34__4_;
      r_34__3_ <= r_n_34__3_;
      r_34__2_ <= r_n_34__2_;
      r_34__1_ <= r_n_34__1_;
      r_34__0_ <= r_n_34__0_;
    end 
    if(N1827) begin
      r_35__31_ <= r_n_35__31_;
      r_35__30_ <= r_n_35__30_;
      r_35__29_ <= r_n_35__29_;
      r_35__28_ <= r_n_35__28_;
      r_35__27_ <= r_n_35__27_;
      r_35__26_ <= r_n_35__26_;
      r_35__25_ <= r_n_35__25_;
      r_35__24_ <= r_n_35__24_;
      r_35__23_ <= r_n_35__23_;
      r_35__22_ <= r_n_35__22_;
      r_35__21_ <= r_n_35__21_;
      r_35__20_ <= r_n_35__20_;
      r_35__19_ <= r_n_35__19_;
      r_35__18_ <= r_n_35__18_;
      r_35__17_ <= r_n_35__17_;
      r_35__16_ <= r_n_35__16_;
      r_35__15_ <= r_n_35__15_;
      r_35__14_ <= r_n_35__14_;
      r_35__13_ <= r_n_35__13_;
      r_35__12_ <= r_n_35__12_;
      r_35__11_ <= r_n_35__11_;
      r_35__10_ <= r_n_35__10_;
      r_35__9_ <= r_n_35__9_;
      r_35__8_ <= r_n_35__8_;
      r_35__7_ <= r_n_35__7_;
      r_35__6_ <= r_n_35__6_;
      r_35__5_ <= r_n_35__5_;
      r_35__4_ <= r_n_35__4_;
      r_35__3_ <= r_n_35__3_;
      r_35__2_ <= r_n_35__2_;
      r_35__1_ <= r_n_35__1_;
      r_35__0_ <= r_n_35__0_;
    end 
    if(N1828) begin
      r_36__31_ <= r_n_36__31_;
      r_36__30_ <= r_n_36__30_;
      r_36__29_ <= r_n_36__29_;
      r_36__28_ <= r_n_36__28_;
      r_36__27_ <= r_n_36__27_;
      r_36__26_ <= r_n_36__26_;
      r_36__25_ <= r_n_36__25_;
      r_36__24_ <= r_n_36__24_;
      r_36__23_ <= r_n_36__23_;
      r_36__22_ <= r_n_36__22_;
      r_36__21_ <= r_n_36__21_;
      r_36__20_ <= r_n_36__20_;
      r_36__19_ <= r_n_36__19_;
      r_36__18_ <= r_n_36__18_;
      r_36__17_ <= r_n_36__17_;
      r_36__16_ <= r_n_36__16_;
      r_36__15_ <= r_n_36__15_;
      r_36__14_ <= r_n_36__14_;
      r_36__13_ <= r_n_36__13_;
      r_36__12_ <= r_n_36__12_;
      r_36__11_ <= r_n_36__11_;
      r_36__10_ <= r_n_36__10_;
      r_36__9_ <= r_n_36__9_;
      r_36__8_ <= r_n_36__8_;
      r_36__7_ <= r_n_36__7_;
      r_36__6_ <= r_n_36__6_;
      r_36__5_ <= r_n_36__5_;
      r_36__4_ <= r_n_36__4_;
      r_36__3_ <= r_n_36__3_;
      r_36__2_ <= r_n_36__2_;
      r_36__1_ <= r_n_36__1_;
      r_36__0_ <= r_n_36__0_;
    end 
    if(N1829) begin
      r_37__31_ <= r_n_37__31_;
      r_37__30_ <= r_n_37__30_;
      r_37__29_ <= r_n_37__29_;
      r_37__28_ <= r_n_37__28_;
      r_37__27_ <= r_n_37__27_;
      r_37__26_ <= r_n_37__26_;
      r_37__25_ <= r_n_37__25_;
      r_37__24_ <= r_n_37__24_;
      r_37__23_ <= r_n_37__23_;
      r_37__22_ <= r_n_37__22_;
      r_37__21_ <= r_n_37__21_;
      r_37__20_ <= r_n_37__20_;
      r_37__19_ <= r_n_37__19_;
      r_37__18_ <= r_n_37__18_;
      r_37__17_ <= r_n_37__17_;
      r_37__16_ <= r_n_37__16_;
      r_37__15_ <= r_n_37__15_;
      r_37__14_ <= r_n_37__14_;
      r_37__13_ <= r_n_37__13_;
      r_37__12_ <= r_n_37__12_;
      r_37__11_ <= r_n_37__11_;
      r_37__10_ <= r_n_37__10_;
      r_37__9_ <= r_n_37__9_;
      r_37__8_ <= r_n_37__8_;
      r_37__7_ <= r_n_37__7_;
      r_37__6_ <= r_n_37__6_;
      r_37__5_ <= r_n_37__5_;
      r_37__4_ <= r_n_37__4_;
      r_37__3_ <= r_n_37__3_;
      r_37__2_ <= r_n_37__2_;
      r_37__1_ <= r_n_37__1_;
      r_37__0_ <= r_n_37__0_;
    end 
    if(N1830) begin
      r_38__31_ <= r_n_38__31_;
      r_38__30_ <= r_n_38__30_;
      r_38__29_ <= r_n_38__29_;
      r_38__28_ <= r_n_38__28_;
      r_38__27_ <= r_n_38__27_;
      r_38__26_ <= r_n_38__26_;
      r_38__25_ <= r_n_38__25_;
      r_38__24_ <= r_n_38__24_;
      r_38__23_ <= r_n_38__23_;
      r_38__22_ <= r_n_38__22_;
      r_38__21_ <= r_n_38__21_;
      r_38__20_ <= r_n_38__20_;
      r_38__19_ <= r_n_38__19_;
      r_38__18_ <= r_n_38__18_;
      r_38__17_ <= r_n_38__17_;
      r_38__16_ <= r_n_38__16_;
      r_38__15_ <= r_n_38__15_;
      r_38__14_ <= r_n_38__14_;
      r_38__13_ <= r_n_38__13_;
      r_38__12_ <= r_n_38__12_;
      r_38__11_ <= r_n_38__11_;
      r_38__10_ <= r_n_38__10_;
      r_38__9_ <= r_n_38__9_;
      r_38__8_ <= r_n_38__8_;
      r_38__7_ <= r_n_38__7_;
      r_38__6_ <= r_n_38__6_;
      r_38__5_ <= r_n_38__5_;
      r_38__4_ <= r_n_38__4_;
      r_38__3_ <= r_n_38__3_;
      r_38__2_ <= r_n_38__2_;
      r_38__1_ <= r_n_38__1_;
      r_38__0_ <= r_n_38__0_;
    end 
    if(N1831) begin
      r_39__31_ <= r_n_39__31_;
      r_39__30_ <= r_n_39__30_;
      r_39__29_ <= r_n_39__29_;
      r_39__28_ <= r_n_39__28_;
      r_39__27_ <= r_n_39__27_;
      r_39__26_ <= r_n_39__26_;
      r_39__25_ <= r_n_39__25_;
      r_39__24_ <= r_n_39__24_;
      r_39__23_ <= r_n_39__23_;
      r_39__22_ <= r_n_39__22_;
      r_39__21_ <= r_n_39__21_;
      r_39__20_ <= r_n_39__20_;
      r_39__19_ <= r_n_39__19_;
      r_39__18_ <= r_n_39__18_;
      r_39__17_ <= r_n_39__17_;
      r_39__16_ <= r_n_39__16_;
      r_39__15_ <= r_n_39__15_;
      r_39__14_ <= r_n_39__14_;
      r_39__13_ <= r_n_39__13_;
      r_39__12_ <= r_n_39__12_;
      r_39__11_ <= r_n_39__11_;
      r_39__10_ <= r_n_39__10_;
      r_39__9_ <= r_n_39__9_;
      r_39__8_ <= r_n_39__8_;
      r_39__7_ <= r_n_39__7_;
      r_39__6_ <= r_n_39__6_;
      r_39__5_ <= r_n_39__5_;
      r_39__4_ <= r_n_39__4_;
      r_39__3_ <= r_n_39__3_;
      r_39__2_ <= r_n_39__2_;
      r_39__1_ <= r_n_39__1_;
      r_39__0_ <= r_n_39__0_;
    end 
    if(N1832) begin
      r_40__31_ <= r_n_40__31_;
      r_40__30_ <= r_n_40__30_;
      r_40__29_ <= r_n_40__29_;
      r_40__28_ <= r_n_40__28_;
      r_40__27_ <= r_n_40__27_;
      r_40__26_ <= r_n_40__26_;
      r_40__25_ <= r_n_40__25_;
      r_40__24_ <= r_n_40__24_;
      r_40__23_ <= r_n_40__23_;
      r_40__22_ <= r_n_40__22_;
      r_40__21_ <= r_n_40__21_;
      r_40__20_ <= r_n_40__20_;
      r_40__19_ <= r_n_40__19_;
      r_40__18_ <= r_n_40__18_;
      r_40__17_ <= r_n_40__17_;
      r_40__16_ <= r_n_40__16_;
      r_40__15_ <= r_n_40__15_;
      r_40__14_ <= r_n_40__14_;
      r_40__13_ <= r_n_40__13_;
      r_40__12_ <= r_n_40__12_;
      r_40__11_ <= r_n_40__11_;
      r_40__10_ <= r_n_40__10_;
      r_40__9_ <= r_n_40__9_;
      r_40__8_ <= r_n_40__8_;
      r_40__7_ <= r_n_40__7_;
      r_40__6_ <= r_n_40__6_;
      r_40__5_ <= r_n_40__5_;
      r_40__4_ <= r_n_40__4_;
      r_40__3_ <= r_n_40__3_;
      r_40__2_ <= r_n_40__2_;
      r_40__1_ <= r_n_40__1_;
      r_40__0_ <= r_n_40__0_;
    end 
    if(N1833) begin
      r_41__31_ <= r_n_41__31_;
      r_41__30_ <= r_n_41__30_;
      r_41__29_ <= r_n_41__29_;
      r_41__28_ <= r_n_41__28_;
      r_41__27_ <= r_n_41__27_;
      r_41__26_ <= r_n_41__26_;
      r_41__25_ <= r_n_41__25_;
      r_41__24_ <= r_n_41__24_;
      r_41__23_ <= r_n_41__23_;
      r_41__22_ <= r_n_41__22_;
      r_41__21_ <= r_n_41__21_;
      r_41__20_ <= r_n_41__20_;
      r_41__19_ <= r_n_41__19_;
      r_41__18_ <= r_n_41__18_;
      r_41__17_ <= r_n_41__17_;
      r_41__16_ <= r_n_41__16_;
      r_41__15_ <= r_n_41__15_;
      r_41__14_ <= r_n_41__14_;
      r_41__13_ <= r_n_41__13_;
      r_41__12_ <= r_n_41__12_;
      r_41__11_ <= r_n_41__11_;
      r_41__10_ <= r_n_41__10_;
      r_41__9_ <= r_n_41__9_;
      r_41__8_ <= r_n_41__8_;
      r_41__7_ <= r_n_41__7_;
      r_41__6_ <= r_n_41__6_;
      r_41__5_ <= r_n_41__5_;
      r_41__4_ <= r_n_41__4_;
      r_41__3_ <= r_n_41__3_;
      r_41__2_ <= r_n_41__2_;
      r_41__1_ <= r_n_41__1_;
      r_41__0_ <= r_n_41__0_;
    end 
    if(N1834) begin
      r_42__31_ <= r_n_42__31_;
      r_42__30_ <= r_n_42__30_;
      r_42__29_ <= r_n_42__29_;
      r_42__28_ <= r_n_42__28_;
      r_42__27_ <= r_n_42__27_;
      r_42__26_ <= r_n_42__26_;
      r_42__25_ <= r_n_42__25_;
      r_42__24_ <= r_n_42__24_;
      r_42__23_ <= r_n_42__23_;
      r_42__22_ <= r_n_42__22_;
      r_42__21_ <= r_n_42__21_;
      r_42__20_ <= r_n_42__20_;
      r_42__19_ <= r_n_42__19_;
      r_42__18_ <= r_n_42__18_;
      r_42__17_ <= r_n_42__17_;
      r_42__16_ <= r_n_42__16_;
      r_42__15_ <= r_n_42__15_;
      r_42__14_ <= r_n_42__14_;
      r_42__13_ <= r_n_42__13_;
      r_42__12_ <= r_n_42__12_;
      r_42__11_ <= r_n_42__11_;
      r_42__10_ <= r_n_42__10_;
      r_42__9_ <= r_n_42__9_;
      r_42__8_ <= r_n_42__8_;
      r_42__7_ <= r_n_42__7_;
      r_42__6_ <= r_n_42__6_;
      r_42__5_ <= r_n_42__5_;
      r_42__4_ <= r_n_42__4_;
      r_42__3_ <= r_n_42__3_;
      r_42__2_ <= r_n_42__2_;
      r_42__1_ <= r_n_42__1_;
      r_42__0_ <= r_n_42__0_;
    end 
    if(N1835) begin
      r_43__31_ <= r_n_43__31_;
      r_43__30_ <= r_n_43__30_;
      r_43__29_ <= r_n_43__29_;
      r_43__28_ <= r_n_43__28_;
      r_43__27_ <= r_n_43__27_;
      r_43__26_ <= r_n_43__26_;
      r_43__25_ <= r_n_43__25_;
      r_43__24_ <= r_n_43__24_;
      r_43__23_ <= r_n_43__23_;
      r_43__22_ <= r_n_43__22_;
      r_43__21_ <= r_n_43__21_;
      r_43__20_ <= r_n_43__20_;
      r_43__19_ <= r_n_43__19_;
      r_43__18_ <= r_n_43__18_;
      r_43__17_ <= r_n_43__17_;
      r_43__16_ <= r_n_43__16_;
      r_43__15_ <= r_n_43__15_;
      r_43__14_ <= r_n_43__14_;
      r_43__13_ <= r_n_43__13_;
      r_43__12_ <= r_n_43__12_;
      r_43__11_ <= r_n_43__11_;
      r_43__10_ <= r_n_43__10_;
      r_43__9_ <= r_n_43__9_;
      r_43__8_ <= r_n_43__8_;
      r_43__7_ <= r_n_43__7_;
      r_43__6_ <= r_n_43__6_;
      r_43__5_ <= r_n_43__5_;
      r_43__4_ <= r_n_43__4_;
      r_43__3_ <= r_n_43__3_;
      r_43__2_ <= r_n_43__2_;
      r_43__1_ <= r_n_43__1_;
      r_43__0_ <= r_n_43__0_;
    end 
    if(N1836) begin
      r_44__31_ <= r_n_44__31_;
      r_44__30_ <= r_n_44__30_;
      r_44__29_ <= r_n_44__29_;
      r_44__28_ <= r_n_44__28_;
      r_44__27_ <= r_n_44__27_;
      r_44__26_ <= r_n_44__26_;
      r_44__25_ <= r_n_44__25_;
      r_44__24_ <= r_n_44__24_;
      r_44__23_ <= r_n_44__23_;
      r_44__22_ <= r_n_44__22_;
      r_44__21_ <= r_n_44__21_;
      r_44__20_ <= r_n_44__20_;
      r_44__19_ <= r_n_44__19_;
      r_44__18_ <= r_n_44__18_;
      r_44__17_ <= r_n_44__17_;
      r_44__16_ <= r_n_44__16_;
      r_44__15_ <= r_n_44__15_;
      r_44__14_ <= r_n_44__14_;
      r_44__13_ <= r_n_44__13_;
      r_44__12_ <= r_n_44__12_;
      r_44__11_ <= r_n_44__11_;
      r_44__10_ <= r_n_44__10_;
      r_44__9_ <= r_n_44__9_;
      r_44__8_ <= r_n_44__8_;
      r_44__7_ <= r_n_44__7_;
      r_44__6_ <= r_n_44__6_;
      r_44__5_ <= r_n_44__5_;
      r_44__4_ <= r_n_44__4_;
      r_44__3_ <= r_n_44__3_;
      r_44__2_ <= r_n_44__2_;
      r_44__1_ <= r_n_44__1_;
      r_44__0_ <= r_n_44__0_;
    end 
    if(N1837) begin
      r_45__31_ <= r_n_45__31_;
      r_45__30_ <= r_n_45__30_;
      r_45__29_ <= r_n_45__29_;
      r_45__28_ <= r_n_45__28_;
      r_45__27_ <= r_n_45__27_;
      r_45__26_ <= r_n_45__26_;
      r_45__25_ <= r_n_45__25_;
      r_45__24_ <= r_n_45__24_;
      r_45__23_ <= r_n_45__23_;
      r_45__22_ <= r_n_45__22_;
      r_45__21_ <= r_n_45__21_;
      r_45__20_ <= r_n_45__20_;
      r_45__19_ <= r_n_45__19_;
      r_45__18_ <= r_n_45__18_;
      r_45__17_ <= r_n_45__17_;
      r_45__16_ <= r_n_45__16_;
      r_45__15_ <= r_n_45__15_;
      r_45__14_ <= r_n_45__14_;
      r_45__13_ <= r_n_45__13_;
      r_45__12_ <= r_n_45__12_;
      r_45__11_ <= r_n_45__11_;
      r_45__10_ <= r_n_45__10_;
      r_45__9_ <= r_n_45__9_;
      r_45__8_ <= r_n_45__8_;
      r_45__7_ <= r_n_45__7_;
      r_45__6_ <= r_n_45__6_;
      r_45__5_ <= r_n_45__5_;
      r_45__4_ <= r_n_45__4_;
      r_45__3_ <= r_n_45__3_;
      r_45__2_ <= r_n_45__2_;
      r_45__1_ <= r_n_45__1_;
      r_45__0_ <= r_n_45__0_;
    end 
    if(N1838) begin
      r_46__31_ <= r_n_46__31_;
      r_46__30_ <= r_n_46__30_;
      r_46__29_ <= r_n_46__29_;
      r_46__28_ <= r_n_46__28_;
      r_46__27_ <= r_n_46__27_;
      r_46__26_ <= r_n_46__26_;
      r_46__25_ <= r_n_46__25_;
      r_46__24_ <= r_n_46__24_;
      r_46__23_ <= r_n_46__23_;
      r_46__22_ <= r_n_46__22_;
      r_46__21_ <= r_n_46__21_;
      r_46__20_ <= r_n_46__20_;
      r_46__19_ <= r_n_46__19_;
      r_46__18_ <= r_n_46__18_;
      r_46__17_ <= r_n_46__17_;
      r_46__16_ <= r_n_46__16_;
      r_46__15_ <= r_n_46__15_;
      r_46__14_ <= r_n_46__14_;
      r_46__13_ <= r_n_46__13_;
      r_46__12_ <= r_n_46__12_;
      r_46__11_ <= r_n_46__11_;
      r_46__10_ <= r_n_46__10_;
      r_46__9_ <= r_n_46__9_;
      r_46__8_ <= r_n_46__8_;
      r_46__7_ <= r_n_46__7_;
      r_46__6_ <= r_n_46__6_;
      r_46__5_ <= r_n_46__5_;
      r_46__4_ <= r_n_46__4_;
      r_46__3_ <= r_n_46__3_;
      r_46__2_ <= r_n_46__2_;
      r_46__1_ <= r_n_46__1_;
      r_46__0_ <= r_n_46__0_;
    end 
    if(N1839) begin
      r_47__31_ <= r_n_47__31_;
      r_47__30_ <= r_n_47__30_;
      r_47__29_ <= r_n_47__29_;
      r_47__28_ <= r_n_47__28_;
      r_47__27_ <= r_n_47__27_;
      r_47__26_ <= r_n_47__26_;
      r_47__25_ <= r_n_47__25_;
      r_47__24_ <= r_n_47__24_;
      r_47__23_ <= r_n_47__23_;
      r_47__22_ <= r_n_47__22_;
      r_47__21_ <= r_n_47__21_;
      r_47__20_ <= r_n_47__20_;
      r_47__19_ <= r_n_47__19_;
      r_47__18_ <= r_n_47__18_;
      r_47__17_ <= r_n_47__17_;
      r_47__16_ <= r_n_47__16_;
      r_47__15_ <= r_n_47__15_;
      r_47__14_ <= r_n_47__14_;
      r_47__13_ <= r_n_47__13_;
      r_47__12_ <= r_n_47__12_;
      r_47__11_ <= r_n_47__11_;
      r_47__10_ <= r_n_47__10_;
      r_47__9_ <= r_n_47__9_;
      r_47__8_ <= r_n_47__8_;
      r_47__7_ <= r_n_47__7_;
      r_47__6_ <= r_n_47__6_;
      r_47__5_ <= r_n_47__5_;
      r_47__4_ <= r_n_47__4_;
      r_47__3_ <= r_n_47__3_;
      r_47__2_ <= r_n_47__2_;
      r_47__1_ <= r_n_47__1_;
      r_47__0_ <= r_n_47__0_;
    end 
    if(N1840) begin
      r_48__31_ <= r_n_48__31_;
      r_48__30_ <= r_n_48__30_;
      r_48__29_ <= r_n_48__29_;
      r_48__28_ <= r_n_48__28_;
      r_48__27_ <= r_n_48__27_;
      r_48__26_ <= r_n_48__26_;
      r_48__25_ <= r_n_48__25_;
      r_48__24_ <= r_n_48__24_;
      r_48__23_ <= r_n_48__23_;
      r_48__22_ <= r_n_48__22_;
      r_48__21_ <= r_n_48__21_;
      r_48__20_ <= r_n_48__20_;
      r_48__19_ <= r_n_48__19_;
      r_48__18_ <= r_n_48__18_;
      r_48__17_ <= r_n_48__17_;
      r_48__16_ <= r_n_48__16_;
      r_48__15_ <= r_n_48__15_;
      r_48__14_ <= r_n_48__14_;
      r_48__13_ <= r_n_48__13_;
      r_48__12_ <= r_n_48__12_;
      r_48__11_ <= r_n_48__11_;
      r_48__10_ <= r_n_48__10_;
      r_48__9_ <= r_n_48__9_;
      r_48__8_ <= r_n_48__8_;
      r_48__7_ <= r_n_48__7_;
      r_48__6_ <= r_n_48__6_;
      r_48__5_ <= r_n_48__5_;
      r_48__4_ <= r_n_48__4_;
      r_48__3_ <= r_n_48__3_;
      r_48__2_ <= r_n_48__2_;
      r_48__1_ <= r_n_48__1_;
      r_48__0_ <= r_n_48__0_;
    end 
    if(N1841) begin
      r_49__31_ <= r_n_49__31_;
      r_49__30_ <= r_n_49__30_;
      r_49__29_ <= r_n_49__29_;
      r_49__28_ <= r_n_49__28_;
      r_49__27_ <= r_n_49__27_;
      r_49__26_ <= r_n_49__26_;
      r_49__25_ <= r_n_49__25_;
      r_49__24_ <= r_n_49__24_;
      r_49__23_ <= r_n_49__23_;
      r_49__22_ <= r_n_49__22_;
      r_49__21_ <= r_n_49__21_;
      r_49__20_ <= r_n_49__20_;
      r_49__19_ <= r_n_49__19_;
      r_49__18_ <= r_n_49__18_;
      r_49__17_ <= r_n_49__17_;
      r_49__16_ <= r_n_49__16_;
      r_49__15_ <= r_n_49__15_;
      r_49__14_ <= r_n_49__14_;
      r_49__13_ <= r_n_49__13_;
      r_49__12_ <= r_n_49__12_;
      r_49__11_ <= r_n_49__11_;
      r_49__10_ <= r_n_49__10_;
      r_49__9_ <= r_n_49__9_;
      r_49__8_ <= r_n_49__8_;
      r_49__7_ <= r_n_49__7_;
      r_49__6_ <= r_n_49__6_;
      r_49__5_ <= r_n_49__5_;
      r_49__4_ <= r_n_49__4_;
      r_49__3_ <= r_n_49__3_;
      r_49__2_ <= r_n_49__2_;
      r_49__1_ <= r_n_49__1_;
      r_49__0_ <= r_n_49__0_;
    end 
    if(N1842) begin
      r_50__31_ <= r_n_50__31_;
      r_50__30_ <= r_n_50__30_;
      r_50__29_ <= r_n_50__29_;
      r_50__28_ <= r_n_50__28_;
      r_50__27_ <= r_n_50__27_;
      r_50__26_ <= r_n_50__26_;
      r_50__25_ <= r_n_50__25_;
      r_50__24_ <= r_n_50__24_;
      r_50__23_ <= r_n_50__23_;
      r_50__22_ <= r_n_50__22_;
      r_50__21_ <= r_n_50__21_;
      r_50__20_ <= r_n_50__20_;
      r_50__19_ <= r_n_50__19_;
      r_50__18_ <= r_n_50__18_;
      r_50__17_ <= r_n_50__17_;
      r_50__16_ <= r_n_50__16_;
      r_50__15_ <= r_n_50__15_;
      r_50__14_ <= r_n_50__14_;
      r_50__13_ <= r_n_50__13_;
      r_50__12_ <= r_n_50__12_;
      r_50__11_ <= r_n_50__11_;
      r_50__10_ <= r_n_50__10_;
      r_50__9_ <= r_n_50__9_;
      r_50__8_ <= r_n_50__8_;
      r_50__7_ <= r_n_50__7_;
      r_50__6_ <= r_n_50__6_;
      r_50__5_ <= r_n_50__5_;
      r_50__4_ <= r_n_50__4_;
      r_50__3_ <= r_n_50__3_;
      r_50__2_ <= r_n_50__2_;
      r_50__1_ <= r_n_50__1_;
      r_50__0_ <= r_n_50__0_;
    end 
    if(N1843) begin
      r_51__31_ <= r_n_51__31_;
      r_51__30_ <= r_n_51__30_;
      r_51__29_ <= r_n_51__29_;
      r_51__28_ <= r_n_51__28_;
      r_51__27_ <= r_n_51__27_;
      r_51__26_ <= r_n_51__26_;
      r_51__25_ <= r_n_51__25_;
      r_51__24_ <= r_n_51__24_;
      r_51__23_ <= r_n_51__23_;
      r_51__22_ <= r_n_51__22_;
      r_51__21_ <= r_n_51__21_;
      r_51__20_ <= r_n_51__20_;
      r_51__19_ <= r_n_51__19_;
      r_51__18_ <= r_n_51__18_;
      r_51__17_ <= r_n_51__17_;
      r_51__16_ <= r_n_51__16_;
      r_51__15_ <= r_n_51__15_;
      r_51__14_ <= r_n_51__14_;
      r_51__13_ <= r_n_51__13_;
      r_51__12_ <= r_n_51__12_;
      r_51__11_ <= r_n_51__11_;
      r_51__10_ <= r_n_51__10_;
      r_51__9_ <= r_n_51__9_;
      r_51__8_ <= r_n_51__8_;
      r_51__7_ <= r_n_51__7_;
      r_51__6_ <= r_n_51__6_;
      r_51__5_ <= r_n_51__5_;
      r_51__4_ <= r_n_51__4_;
      r_51__3_ <= r_n_51__3_;
      r_51__2_ <= r_n_51__2_;
      r_51__1_ <= r_n_51__1_;
      r_51__0_ <= r_n_51__0_;
    end 
    if(N1844) begin
      r_52__31_ <= r_n_52__31_;
      r_52__30_ <= r_n_52__30_;
      r_52__29_ <= r_n_52__29_;
      r_52__28_ <= r_n_52__28_;
      r_52__27_ <= r_n_52__27_;
      r_52__26_ <= r_n_52__26_;
      r_52__25_ <= r_n_52__25_;
      r_52__24_ <= r_n_52__24_;
      r_52__23_ <= r_n_52__23_;
      r_52__22_ <= r_n_52__22_;
      r_52__21_ <= r_n_52__21_;
      r_52__20_ <= r_n_52__20_;
      r_52__19_ <= r_n_52__19_;
      r_52__18_ <= r_n_52__18_;
      r_52__17_ <= r_n_52__17_;
      r_52__16_ <= r_n_52__16_;
      r_52__15_ <= r_n_52__15_;
      r_52__14_ <= r_n_52__14_;
      r_52__13_ <= r_n_52__13_;
      r_52__12_ <= r_n_52__12_;
      r_52__11_ <= r_n_52__11_;
      r_52__10_ <= r_n_52__10_;
      r_52__9_ <= r_n_52__9_;
      r_52__8_ <= r_n_52__8_;
      r_52__7_ <= r_n_52__7_;
      r_52__6_ <= r_n_52__6_;
      r_52__5_ <= r_n_52__5_;
      r_52__4_ <= r_n_52__4_;
      r_52__3_ <= r_n_52__3_;
      r_52__2_ <= r_n_52__2_;
      r_52__1_ <= r_n_52__1_;
      r_52__0_ <= r_n_52__0_;
    end 
    if(N1845) begin
      r_53__31_ <= r_n_53__31_;
      r_53__30_ <= r_n_53__30_;
      r_53__29_ <= r_n_53__29_;
      r_53__28_ <= r_n_53__28_;
      r_53__27_ <= r_n_53__27_;
      r_53__26_ <= r_n_53__26_;
      r_53__25_ <= r_n_53__25_;
      r_53__24_ <= r_n_53__24_;
      r_53__23_ <= r_n_53__23_;
      r_53__22_ <= r_n_53__22_;
      r_53__21_ <= r_n_53__21_;
      r_53__20_ <= r_n_53__20_;
      r_53__19_ <= r_n_53__19_;
      r_53__18_ <= r_n_53__18_;
      r_53__17_ <= r_n_53__17_;
      r_53__16_ <= r_n_53__16_;
      r_53__15_ <= r_n_53__15_;
      r_53__14_ <= r_n_53__14_;
      r_53__13_ <= r_n_53__13_;
      r_53__12_ <= r_n_53__12_;
      r_53__11_ <= r_n_53__11_;
      r_53__10_ <= r_n_53__10_;
      r_53__9_ <= r_n_53__9_;
      r_53__8_ <= r_n_53__8_;
      r_53__7_ <= r_n_53__7_;
      r_53__6_ <= r_n_53__6_;
      r_53__5_ <= r_n_53__5_;
      r_53__4_ <= r_n_53__4_;
      r_53__3_ <= r_n_53__3_;
      r_53__2_ <= r_n_53__2_;
      r_53__1_ <= r_n_53__1_;
      r_53__0_ <= r_n_53__0_;
    end 
    if(N1846) begin
      r_54__31_ <= r_n_54__31_;
      r_54__30_ <= r_n_54__30_;
      r_54__29_ <= r_n_54__29_;
      r_54__28_ <= r_n_54__28_;
      r_54__27_ <= r_n_54__27_;
      r_54__26_ <= r_n_54__26_;
      r_54__25_ <= r_n_54__25_;
      r_54__24_ <= r_n_54__24_;
      r_54__23_ <= r_n_54__23_;
      r_54__22_ <= r_n_54__22_;
      r_54__21_ <= r_n_54__21_;
      r_54__20_ <= r_n_54__20_;
      r_54__19_ <= r_n_54__19_;
      r_54__18_ <= r_n_54__18_;
      r_54__17_ <= r_n_54__17_;
      r_54__16_ <= r_n_54__16_;
      r_54__15_ <= r_n_54__15_;
      r_54__14_ <= r_n_54__14_;
      r_54__13_ <= r_n_54__13_;
      r_54__12_ <= r_n_54__12_;
      r_54__11_ <= r_n_54__11_;
      r_54__10_ <= r_n_54__10_;
      r_54__9_ <= r_n_54__9_;
      r_54__8_ <= r_n_54__8_;
      r_54__7_ <= r_n_54__7_;
      r_54__6_ <= r_n_54__6_;
      r_54__5_ <= r_n_54__5_;
      r_54__4_ <= r_n_54__4_;
      r_54__3_ <= r_n_54__3_;
      r_54__2_ <= r_n_54__2_;
      r_54__1_ <= r_n_54__1_;
      r_54__0_ <= r_n_54__0_;
    end 
    if(N1847) begin
      r_55__31_ <= r_n_55__31_;
      r_55__30_ <= r_n_55__30_;
      r_55__29_ <= r_n_55__29_;
      r_55__28_ <= r_n_55__28_;
      r_55__27_ <= r_n_55__27_;
      r_55__26_ <= r_n_55__26_;
      r_55__25_ <= r_n_55__25_;
      r_55__24_ <= r_n_55__24_;
      r_55__23_ <= r_n_55__23_;
      r_55__22_ <= r_n_55__22_;
      r_55__21_ <= r_n_55__21_;
      r_55__20_ <= r_n_55__20_;
      r_55__19_ <= r_n_55__19_;
      r_55__18_ <= r_n_55__18_;
      r_55__17_ <= r_n_55__17_;
      r_55__16_ <= r_n_55__16_;
      r_55__15_ <= r_n_55__15_;
      r_55__14_ <= r_n_55__14_;
      r_55__13_ <= r_n_55__13_;
      r_55__12_ <= r_n_55__12_;
      r_55__11_ <= r_n_55__11_;
      r_55__10_ <= r_n_55__10_;
      r_55__9_ <= r_n_55__9_;
      r_55__8_ <= r_n_55__8_;
      r_55__7_ <= r_n_55__7_;
      r_55__6_ <= r_n_55__6_;
      r_55__5_ <= r_n_55__5_;
      r_55__4_ <= r_n_55__4_;
      r_55__3_ <= r_n_55__3_;
      r_55__2_ <= r_n_55__2_;
      r_55__1_ <= r_n_55__1_;
      r_55__0_ <= r_n_55__0_;
    end 
    if(N1848) begin
      r_56__31_ <= r_n_56__31_;
      r_56__30_ <= r_n_56__30_;
      r_56__29_ <= r_n_56__29_;
      r_56__28_ <= r_n_56__28_;
      r_56__27_ <= r_n_56__27_;
      r_56__26_ <= r_n_56__26_;
      r_56__25_ <= r_n_56__25_;
      r_56__24_ <= r_n_56__24_;
      r_56__23_ <= r_n_56__23_;
      r_56__22_ <= r_n_56__22_;
      r_56__21_ <= r_n_56__21_;
      r_56__20_ <= r_n_56__20_;
      r_56__19_ <= r_n_56__19_;
      r_56__18_ <= r_n_56__18_;
      r_56__17_ <= r_n_56__17_;
      r_56__16_ <= r_n_56__16_;
      r_56__15_ <= r_n_56__15_;
      r_56__14_ <= r_n_56__14_;
      r_56__13_ <= r_n_56__13_;
      r_56__12_ <= r_n_56__12_;
      r_56__11_ <= r_n_56__11_;
      r_56__10_ <= r_n_56__10_;
      r_56__9_ <= r_n_56__9_;
      r_56__8_ <= r_n_56__8_;
      r_56__7_ <= r_n_56__7_;
      r_56__6_ <= r_n_56__6_;
      r_56__5_ <= r_n_56__5_;
      r_56__4_ <= r_n_56__4_;
      r_56__3_ <= r_n_56__3_;
      r_56__2_ <= r_n_56__2_;
      r_56__1_ <= r_n_56__1_;
      r_56__0_ <= r_n_56__0_;
    end 
    if(N1849) begin
      r_57__31_ <= r_n_57__31_;
      r_57__30_ <= r_n_57__30_;
      r_57__29_ <= r_n_57__29_;
      r_57__28_ <= r_n_57__28_;
      r_57__27_ <= r_n_57__27_;
      r_57__26_ <= r_n_57__26_;
      r_57__25_ <= r_n_57__25_;
      r_57__24_ <= r_n_57__24_;
      r_57__23_ <= r_n_57__23_;
      r_57__22_ <= r_n_57__22_;
      r_57__21_ <= r_n_57__21_;
      r_57__20_ <= r_n_57__20_;
      r_57__19_ <= r_n_57__19_;
      r_57__18_ <= r_n_57__18_;
      r_57__17_ <= r_n_57__17_;
      r_57__16_ <= r_n_57__16_;
      r_57__15_ <= r_n_57__15_;
      r_57__14_ <= r_n_57__14_;
      r_57__13_ <= r_n_57__13_;
      r_57__12_ <= r_n_57__12_;
      r_57__11_ <= r_n_57__11_;
      r_57__10_ <= r_n_57__10_;
      r_57__9_ <= r_n_57__9_;
      r_57__8_ <= r_n_57__8_;
      r_57__7_ <= r_n_57__7_;
      r_57__6_ <= r_n_57__6_;
      r_57__5_ <= r_n_57__5_;
      r_57__4_ <= r_n_57__4_;
      r_57__3_ <= r_n_57__3_;
      r_57__2_ <= r_n_57__2_;
      r_57__1_ <= r_n_57__1_;
      r_57__0_ <= r_n_57__0_;
    end 
    if(N1850) begin
      r_58__31_ <= r_n_58__31_;
      r_58__30_ <= r_n_58__30_;
      r_58__29_ <= r_n_58__29_;
      r_58__28_ <= r_n_58__28_;
      r_58__27_ <= r_n_58__27_;
      r_58__26_ <= r_n_58__26_;
      r_58__25_ <= r_n_58__25_;
      r_58__24_ <= r_n_58__24_;
      r_58__23_ <= r_n_58__23_;
      r_58__22_ <= r_n_58__22_;
      r_58__21_ <= r_n_58__21_;
      r_58__20_ <= r_n_58__20_;
      r_58__19_ <= r_n_58__19_;
      r_58__18_ <= r_n_58__18_;
      r_58__17_ <= r_n_58__17_;
      r_58__16_ <= r_n_58__16_;
      r_58__15_ <= r_n_58__15_;
      r_58__14_ <= r_n_58__14_;
      r_58__13_ <= r_n_58__13_;
      r_58__12_ <= r_n_58__12_;
      r_58__11_ <= r_n_58__11_;
      r_58__10_ <= r_n_58__10_;
      r_58__9_ <= r_n_58__9_;
      r_58__8_ <= r_n_58__8_;
      r_58__7_ <= r_n_58__7_;
      r_58__6_ <= r_n_58__6_;
      r_58__5_ <= r_n_58__5_;
      r_58__4_ <= r_n_58__4_;
      r_58__3_ <= r_n_58__3_;
      r_58__2_ <= r_n_58__2_;
      r_58__1_ <= r_n_58__1_;
      r_58__0_ <= r_n_58__0_;
    end 
    if(N1851) begin
      r_59__31_ <= r_n_59__31_;
      r_59__30_ <= r_n_59__30_;
      r_59__29_ <= r_n_59__29_;
      r_59__28_ <= r_n_59__28_;
      r_59__27_ <= r_n_59__27_;
      r_59__26_ <= r_n_59__26_;
      r_59__25_ <= r_n_59__25_;
      r_59__24_ <= r_n_59__24_;
      r_59__23_ <= r_n_59__23_;
      r_59__22_ <= r_n_59__22_;
      r_59__21_ <= r_n_59__21_;
      r_59__20_ <= r_n_59__20_;
      r_59__19_ <= r_n_59__19_;
      r_59__18_ <= r_n_59__18_;
      r_59__17_ <= r_n_59__17_;
      r_59__16_ <= r_n_59__16_;
      r_59__15_ <= r_n_59__15_;
      r_59__14_ <= r_n_59__14_;
      r_59__13_ <= r_n_59__13_;
      r_59__12_ <= r_n_59__12_;
      r_59__11_ <= r_n_59__11_;
      r_59__10_ <= r_n_59__10_;
      r_59__9_ <= r_n_59__9_;
      r_59__8_ <= r_n_59__8_;
      r_59__7_ <= r_n_59__7_;
      r_59__6_ <= r_n_59__6_;
      r_59__5_ <= r_n_59__5_;
      r_59__4_ <= r_n_59__4_;
      r_59__3_ <= r_n_59__3_;
      r_59__2_ <= r_n_59__2_;
      r_59__1_ <= r_n_59__1_;
      r_59__0_ <= r_n_59__0_;
    end 
    if(N1852) begin
      r_60__31_ <= r_n_60__31_;
      r_60__30_ <= r_n_60__30_;
      r_60__29_ <= r_n_60__29_;
      r_60__28_ <= r_n_60__28_;
      r_60__27_ <= r_n_60__27_;
      r_60__26_ <= r_n_60__26_;
      r_60__25_ <= r_n_60__25_;
      r_60__24_ <= r_n_60__24_;
      r_60__23_ <= r_n_60__23_;
      r_60__22_ <= r_n_60__22_;
      r_60__21_ <= r_n_60__21_;
      r_60__20_ <= r_n_60__20_;
      r_60__19_ <= r_n_60__19_;
      r_60__18_ <= r_n_60__18_;
      r_60__17_ <= r_n_60__17_;
      r_60__16_ <= r_n_60__16_;
      r_60__15_ <= r_n_60__15_;
      r_60__14_ <= r_n_60__14_;
      r_60__13_ <= r_n_60__13_;
      r_60__12_ <= r_n_60__12_;
      r_60__11_ <= r_n_60__11_;
      r_60__10_ <= r_n_60__10_;
      r_60__9_ <= r_n_60__9_;
      r_60__8_ <= r_n_60__8_;
      r_60__7_ <= r_n_60__7_;
      r_60__6_ <= r_n_60__6_;
      r_60__5_ <= r_n_60__5_;
      r_60__4_ <= r_n_60__4_;
      r_60__3_ <= r_n_60__3_;
      r_60__2_ <= r_n_60__2_;
      r_60__1_ <= r_n_60__1_;
      r_60__0_ <= r_n_60__0_;
    end 
    if(N1853) begin
      r_61__31_ <= r_n_61__31_;
      r_61__30_ <= r_n_61__30_;
      r_61__29_ <= r_n_61__29_;
      r_61__28_ <= r_n_61__28_;
      r_61__27_ <= r_n_61__27_;
      r_61__26_ <= r_n_61__26_;
      r_61__25_ <= r_n_61__25_;
      r_61__24_ <= r_n_61__24_;
      r_61__23_ <= r_n_61__23_;
      r_61__22_ <= r_n_61__22_;
      r_61__21_ <= r_n_61__21_;
      r_61__20_ <= r_n_61__20_;
      r_61__19_ <= r_n_61__19_;
      r_61__18_ <= r_n_61__18_;
      r_61__17_ <= r_n_61__17_;
      r_61__16_ <= r_n_61__16_;
      r_61__15_ <= r_n_61__15_;
      r_61__14_ <= r_n_61__14_;
      r_61__13_ <= r_n_61__13_;
      r_61__12_ <= r_n_61__12_;
      r_61__11_ <= r_n_61__11_;
      r_61__10_ <= r_n_61__10_;
      r_61__9_ <= r_n_61__9_;
      r_61__8_ <= r_n_61__8_;
      r_61__7_ <= r_n_61__7_;
      r_61__6_ <= r_n_61__6_;
      r_61__5_ <= r_n_61__5_;
      r_61__4_ <= r_n_61__4_;
      r_61__3_ <= r_n_61__3_;
      r_61__2_ <= r_n_61__2_;
      r_61__1_ <= r_n_61__1_;
      r_61__0_ <= r_n_61__0_;
    end 
    if(N1854) begin
      r_62__31_ <= r_n_62__31_;
      r_62__30_ <= r_n_62__30_;
      r_62__29_ <= r_n_62__29_;
      r_62__28_ <= r_n_62__28_;
      r_62__27_ <= r_n_62__27_;
      r_62__26_ <= r_n_62__26_;
      r_62__25_ <= r_n_62__25_;
      r_62__24_ <= r_n_62__24_;
      r_62__23_ <= r_n_62__23_;
      r_62__22_ <= r_n_62__22_;
      r_62__21_ <= r_n_62__21_;
      r_62__20_ <= r_n_62__20_;
      r_62__19_ <= r_n_62__19_;
      r_62__18_ <= r_n_62__18_;
      r_62__17_ <= r_n_62__17_;
      r_62__16_ <= r_n_62__16_;
      r_62__15_ <= r_n_62__15_;
      r_62__14_ <= r_n_62__14_;
      r_62__13_ <= r_n_62__13_;
      r_62__12_ <= r_n_62__12_;
      r_62__11_ <= r_n_62__11_;
      r_62__10_ <= r_n_62__10_;
      r_62__9_ <= r_n_62__9_;
      r_62__8_ <= r_n_62__8_;
      r_62__7_ <= r_n_62__7_;
      r_62__6_ <= r_n_62__6_;
      r_62__5_ <= r_n_62__5_;
      r_62__4_ <= r_n_62__4_;
      r_62__3_ <= r_n_62__3_;
      r_62__2_ <= r_n_62__2_;
      r_62__1_ <= r_n_62__1_;
      r_62__0_ <= r_n_62__0_;
    end 
    if(N1855) begin
      r_63__31_ <= r_n_63__31_;
      r_63__30_ <= r_n_63__30_;
      r_63__29_ <= r_n_63__29_;
      r_63__28_ <= r_n_63__28_;
      r_63__27_ <= r_n_63__27_;
      r_63__26_ <= r_n_63__26_;
      r_63__25_ <= r_n_63__25_;
      r_63__24_ <= r_n_63__24_;
      r_63__23_ <= r_n_63__23_;
      r_63__22_ <= r_n_63__22_;
      r_63__21_ <= r_n_63__21_;
      r_63__20_ <= r_n_63__20_;
      r_63__19_ <= r_n_63__19_;
      r_63__18_ <= r_n_63__18_;
      r_63__17_ <= r_n_63__17_;
      r_63__16_ <= r_n_63__16_;
      r_63__15_ <= r_n_63__15_;
      r_63__14_ <= r_n_63__14_;
      r_63__13_ <= r_n_63__13_;
      r_63__12_ <= r_n_63__12_;
      r_63__11_ <= r_n_63__11_;
      r_63__10_ <= r_n_63__10_;
      r_63__9_ <= r_n_63__9_;
      r_63__8_ <= r_n_63__8_;
      r_63__7_ <= r_n_63__7_;
      r_63__6_ <= r_n_63__6_;
      r_63__5_ <= r_n_63__5_;
      r_63__4_ <= r_n_63__4_;
      r_63__3_ <= r_n_63__3_;
      r_63__2_ <= r_n_63__2_;
      r_63__1_ <= r_n_63__1_;
      r_63__0_ <= r_n_63__0_;
    end 
    if(N1856) begin
      r_64__31_ <= r_n_64__31_;
      r_64__30_ <= r_n_64__30_;
      r_64__29_ <= r_n_64__29_;
      r_64__28_ <= r_n_64__28_;
      r_64__27_ <= r_n_64__27_;
      r_64__26_ <= r_n_64__26_;
      r_64__25_ <= r_n_64__25_;
      r_64__24_ <= r_n_64__24_;
      r_64__23_ <= r_n_64__23_;
      r_64__22_ <= r_n_64__22_;
      r_64__21_ <= r_n_64__21_;
      r_64__20_ <= r_n_64__20_;
      r_64__19_ <= r_n_64__19_;
      r_64__18_ <= r_n_64__18_;
      r_64__17_ <= r_n_64__17_;
      r_64__16_ <= r_n_64__16_;
      r_64__15_ <= r_n_64__15_;
      r_64__14_ <= r_n_64__14_;
      r_64__13_ <= r_n_64__13_;
      r_64__12_ <= r_n_64__12_;
      r_64__11_ <= r_n_64__11_;
      r_64__10_ <= r_n_64__10_;
      r_64__9_ <= r_n_64__9_;
      r_64__8_ <= r_n_64__8_;
      r_64__7_ <= r_n_64__7_;
      r_64__6_ <= r_n_64__6_;
      r_64__5_ <= r_n_64__5_;
      r_64__4_ <= r_n_64__4_;
      r_64__3_ <= r_n_64__3_;
      r_64__2_ <= r_n_64__2_;
      r_64__1_ <= r_n_64__1_;
      r_64__0_ <= r_n_64__0_;
    end 
    if(N1857) begin
      r_65__31_ <= r_n_65__31_;
      r_65__30_ <= r_n_65__30_;
      r_65__29_ <= r_n_65__29_;
      r_65__28_ <= r_n_65__28_;
      r_65__27_ <= r_n_65__27_;
      r_65__26_ <= r_n_65__26_;
      r_65__25_ <= r_n_65__25_;
      r_65__24_ <= r_n_65__24_;
      r_65__23_ <= r_n_65__23_;
      r_65__22_ <= r_n_65__22_;
      r_65__21_ <= r_n_65__21_;
      r_65__20_ <= r_n_65__20_;
      r_65__19_ <= r_n_65__19_;
      r_65__18_ <= r_n_65__18_;
      r_65__17_ <= r_n_65__17_;
      r_65__16_ <= r_n_65__16_;
      r_65__15_ <= r_n_65__15_;
      r_65__14_ <= r_n_65__14_;
      r_65__13_ <= r_n_65__13_;
      r_65__12_ <= r_n_65__12_;
      r_65__11_ <= r_n_65__11_;
      r_65__10_ <= r_n_65__10_;
      r_65__9_ <= r_n_65__9_;
      r_65__8_ <= r_n_65__8_;
      r_65__7_ <= r_n_65__7_;
      r_65__6_ <= r_n_65__6_;
      r_65__5_ <= r_n_65__5_;
      r_65__4_ <= r_n_65__4_;
      r_65__3_ <= r_n_65__3_;
      r_65__2_ <= r_n_65__2_;
      r_65__1_ <= r_n_65__1_;
      r_65__0_ <= r_n_65__0_;
    end 
    if(N1858) begin
      r_66__31_ <= r_n_66__31_;
      r_66__30_ <= r_n_66__30_;
      r_66__29_ <= r_n_66__29_;
      r_66__28_ <= r_n_66__28_;
      r_66__27_ <= r_n_66__27_;
      r_66__26_ <= r_n_66__26_;
      r_66__25_ <= r_n_66__25_;
      r_66__24_ <= r_n_66__24_;
      r_66__23_ <= r_n_66__23_;
      r_66__22_ <= r_n_66__22_;
      r_66__21_ <= r_n_66__21_;
      r_66__20_ <= r_n_66__20_;
      r_66__19_ <= r_n_66__19_;
      r_66__18_ <= r_n_66__18_;
      r_66__17_ <= r_n_66__17_;
      r_66__16_ <= r_n_66__16_;
      r_66__15_ <= r_n_66__15_;
      r_66__14_ <= r_n_66__14_;
      r_66__13_ <= r_n_66__13_;
      r_66__12_ <= r_n_66__12_;
      r_66__11_ <= r_n_66__11_;
      r_66__10_ <= r_n_66__10_;
      r_66__9_ <= r_n_66__9_;
      r_66__8_ <= r_n_66__8_;
      r_66__7_ <= r_n_66__7_;
      r_66__6_ <= r_n_66__6_;
      r_66__5_ <= r_n_66__5_;
      r_66__4_ <= r_n_66__4_;
      r_66__3_ <= r_n_66__3_;
      r_66__2_ <= r_n_66__2_;
      r_66__1_ <= r_n_66__1_;
      r_66__0_ <= r_n_66__0_;
    end 
    if(N1859) begin
      r_67__31_ <= r_n_67__31_;
      r_67__30_ <= r_n_67__30_;
      r_67__29_ <= r_n_67__29_;
      r_67__28_ <= r_n_67__28_;
      r_67__27_ <= r_n_67__27_;
      r_67__26_ <= r_n_67__26_;
      r_67__25_ <= r_n_67__25_;
      r_67__24_ <= r_n_67__24_;
      r_67__23_ <= r_n_67__23_;
      r_67__22_ <= r_n_67__22_;
      r_67__21_ <= r_n_67__21_;
      r_67__20_ <= r_n_67__20_;
      r_67__19_ <= r_n_67__19_;
      r_67__18_ <= r_n_67__18_;
      r_67__17_ <= r_n_67__17_;
      r_67__16_ <= r_n_67__16_;
      r_67__15_ <= r_n_67__15_;
      r_67__14_ <= r_n_67__14_;
      r_67__13_ <= r_n_67__13_;
      r_67__12_ <= r_n_67__12_;
      r_67__11_ <= r_n_67__11_;
      r_67__10_ <= r_n_67__10_;
      r_67__9_ <= r_n_67__9_;
      r_67__8_ <= r_n_67__8_;
      r_67__7_ <= r_n_67__7_;
      r_67__6_ <= r_n_67__6_;
      r_67__5_ <= r_n_67__5_;
      r_67__4_ <= r_n_67__4_;
      r_67__3_ <= r_n_67__3_;
      r_67__2_ <= r_n_67__2_;
      r_67__1_ <= r_n_67__1_;
      r_67__0_ <= r_n_67__0_;
    end 
    if(N1860) begin
      r_68__31_ <= r_n_68__31_;
      r_68__30_ <= r_n_68__30_;
      r_68__29_ <= r_n_68__29_;
      r_68__28_ <= r_n_68__28_;
      r_68__27_ <= r_n_68__27_;
      r_68__26_ <= r_n_68__26_;
      r_68__25_ <= r_n_68__25_;
      r_68__24_ <= r_n_68__24_;
      r_68__23_ <= r_n_68__23_;
      r_68__22_ <= r_n_68__22_;
      r_68__21_ <= r_n_68__21_;
      r_68__20_ <= r_n_68__20_;
      r_68__19_ <= r_n_68__19_;
      r_68__18_ <= r_n_68__18_;
      r_68__17_ <= r_n_68__17_;
      r_68__16_ <= r_n_68__16_;
      r_68__15_ <= r_n_68__15_;
      r_68__14_ <= r_n_68__14_;
      r_68__13_ <= r_n_68__13_;
      r_68__12_ <= r_n_68__12_;
      r_68__11_ <= r_n_68__11_;
      r_68__10_ <= r_n_68__10_;
      r_68__9_ <= r_n_68__9_;
      r_68__8_ <= r_n_68__8_;
      r_68__7_ <= r_n_68__7_;
      r_68__6_ <= r_n_68__6_;
      r_68__5_ <= r_n_68__5_;
      r_68__4_ <= r_n_68__4_;
      r_68__3_ <= r_n_68__3_;
      r_68__2_ <= r_n_68__2_;
      r_68__1_ <= r_n_68__1_;
      r_68__0_ <= r_n_68__0_;
    end 
    if(N1861) begin
      r_69__31_ <= r_n_69__31_;
      r_69__30_ <= r_n_69__30_;
      r_69__29_ <= r_n_69__29_;
      r_69__28_ <= r_n_69__28_;
      r_69__27_ <= r_n_69__27_;
      r_69__26_ <= r_n_69__26_;
      r_69__25_ <= r_n_69__25_;
      r_69__24_ <= r_n_69__24_;
      r_69__23_ <= r_n_69__23_;
      r_69__22_ <= r_n_69__22_;
      r_69__21_ <= r_n_69__21_;
      r_69__20_ <= r_n_69__20_;
      r_69__19_ <= r_n_69__19_;
      r_69__18_ <= r_n_69__18_;
      r_69__17_ <= r_n_69__17_;
      r_69__16_ <= r_n_69__16_;
      r_69__15_ <= r_n_69__15_;
      r_69__14_ <= r_n_69__14_;
      r_69__13_ <= r_n_69__13_;
      r_69__12_ <= r_n_69__12_;
      r_69__11_ <= r_n_69__11_;
      r_69__10_ <= r_n_69__10_;
      r_69__9_ <= r_n_69__9_;
      r_69__8_ <= r_n_69__8_;
      r_69__7_ <= r_n_69__7_;
      r_69__6_ <= r_n_69__6_;
      r_69__5_ <= r_n_69__5_;
      r_69__4_ <= r_n_69__4_;
      r_69__3_ <= r_n_69__3_;
      r_69__2_ <= r_n_69__2_;
      r_69__1_ <= r_n_69__1_;
      r_69__0_ <= r_n_69__0_;
    end 
    if(N1862) begin
      r_70__31_ <= r_n_70__31_;
      r_70__30_ <= r_n_70__30_;
      r_70__29_ <= r_n_70__29_;
      r_70__28_ <= r_n_70__28_;
      r_70__27_ <= r_n_70__27_;
      r_70__26_ <= r_n_70__26_;
      r_70__25_ <= r_n_70__25_;
      r_70__24_ <= r_n_70__24_;
      r_70__23_ <= r_n_70__23_;
      r_70__22_ <= r_n_70__22_;
      r_70__21_ <= r_n_70__21_;
      r_70__20_ <= r_n_70__20_;
      r_70__19_ <= r_n_70__19_;
      r_70__18_ <= r_n_70__18_;
      r_70__17_ <= r_n_70__17_;
      r_70__16_ <= r_n_70__16_;
      r_70__15_ <= r_n_70__15_;
      r_70__14_ <= r_n_70__14_;
      r_70__13_ <= r_n_70__13_;
      r_70__12_ <= r_n_70__12_;
      r_70__11_ <= r_n_70__11_;
      r_70__10_ <= r_n_70__10_;
      r_70__9_ <= r_n_70__9_;
      r_70__8_ <= r_n_70__8_;
      r_70__7_ <= r_n_70__7_;
      r_70__6_ <= r_n_70__6_;
      r_70__5_ <= r_n_70__5_;
      r_70__4_ <= r_n_70__4_;
      r_70__3_ <= r_n_70__3_;
      r_70__2_ <= r_n_70__2_;
      r_70__1_ <= r_n_70__1_;
      r_70__0_ <= r_n_70__0_;
    end 
    if(N1863) begin
      r_71__31_ <= r_n_71__31_;
      r_71__30_ <= r_n_71__30_;
      r_71__29_ <= r_n_71__29_;
      r_71__28_ <= r_n_71__28_;
      r_71__27_ <= r_n_71__27_;
      r_71__26_ <= r_n_71__26_;
      r_71__25_ <= r_n_71__25_;
      r_71__24_ <= r_n_71__24_;
      r_71__23_ <= r_n_71__23_;
      r_71__22_ <= r_n_71__22_;
      r_71__21_ <= r_n_71__21_;
      r_71__20_ <= r_n_71__20_;
      r_71__19_ <= r_n_71__19_;
      r_71__18_ <= r_n_71__18_;
      r_71__17_ <= r_n_71__17_;
      r_71__16_ <= r_n_71__16_;
      r_71__15_ <= r_n_71__15_;
      r_71__14_ <= r_n_71__14_;
      r_71__13_ <= r_n_71__13_;
      r_71__12_ <= r_n_71__12_;
      r_71__11_ <= r_n_71__11_;
      r_71__10_ <= r_n_71__10_;
      r_71__9_ <= r_n_71__9_;
      r_71__8_ <= r_n_71__8_;
      r_71__7_ <= r_n_71__7_;
      r_71__6_ <= r_n_71__6_;
      r_71__5_ <= r_n_71__5_;
      r_71__4_ <= r_n_71__4_;
      r_71__3_ <= r_n_71__3_;
      r_71__2_ <= r_n_71__2_;
      r_71__1_ <= r_n_71__1_;
      r_71__0_ <= r_n_71__0_;
    end 
    if(N1864) begin
      r_72__31_ <= r_n_72__31_;
      r_72__30_ <= r_n_72__30_;
      r_72__29_ <= r_n_72__29_;
      r_72__28_ <= r_n_72__28_;
      r_72__27_ <= r_n_72__27_;
      r_72__26_ <= r_n_72__26_;
      r_72__25_ <= r_n_72__25_;
      r_72__24_ <= r_n_72__24_;
      r_72__23_ <= r_n_72__23_;
      r_72__22_ <= r_n_72__22_;
      r_72__21_ <= r_n_72__21_;
      r_72__20_ <= r_n_72__20_;
      r_72__19_ <= r_n_72__19_;
      r_72__18_ <= r_n_72__18_;
      r_72__17_ <= r_n_72__17_;
      r_72__16_ <= r_n_72__16_;
      r_72__15_ <= r_n_72__15_;
      r_72__14_ <= r_n_72__14_;
      r_72__13_ <= r_n_72__13_;
      r_72__12_ <= r_n_72__12_;
      r_72__11_ <= r_n_72__11_;
      r_72__10_ <= r_n_72__10_;
      r_72__9_ <= r_n_72__9_;
      r_72__8_ <= r_n_72__8_;
      r_72__7_ <= r_n_72__7_;
      r_72__6_ <= r_n_72__6_;
      r_72__5_ <= r_n_72__5_;
      r_72__4_ <= r_n_72__4_;
      r_72__3_ <= r_n_72__3_;
      r_72__2_ <= r_n_72__2_;
      r_72__1_ <= r_n_72__1_;
      r_72__0_ <= r_n_72__0_;
    end 
    if(N1865) begin
      r_73__31_ <= r_n_73__31_;
      r_73__30_ <= r_n_73__30_;
      r_73__29_ <= r_n_73__29_;
      r_73__28_ <= r_n_73__28_;
      r_73__27_ <= r_n_73__27_;
      r_73__26_ <= r_n_73__26_;
      r_73__25_ <= r_n_73__25_;
      r_73__24_ <= r_n_73__24_;
      r_73__23_ <= r_n_73__23_;
      r_73__22_ <= r_n_73__22_;
      r_73__21_ <= r_n_73__21_;
      r_73__20_ <= r_n_73__20_;
      r_73__19_ <= r_n_73__19_;
      r_73__18_ <= r_n_73__18_;
      r_73__17_ <= r_n_73__17_;
      r_73__16_ <= r_n_73__16_;
      r_73__15_ <= r_n_73__15_;
      r_73__14_ <= r_n_73__14_;
      r_73__13_ <= r_n_73__13_;
      r_73__12_ <= r_n_73__12_;
      r_73__11_ <= r_n_73__11_;
      r_73__10_ <= r_n_73__10_;
      r_73__9_ <= r_n_73__9_;
      r_73__8_ <= r_n_73__8_;
      r_73__7_ <= r_n_73__7_;
      r_73__6_ <= r_n_73__6_;
      r_73__5_ <= r_n_73__5_;
      r_73__4_ <= r_n_73__4_;
      r_73__3_ <= r_n_73__3_;
      r_73__2_ <= r_n_73__2_;
      r_73__1_ <= r_n_73__1_;
      r_73__0_ <= r_n_73__0_;
    end 
    if(N1866) begin
      r_74__31_ <= r_n_74__31_;
      r_74__30_ <= r_n_74__30_;
      r_74__29_ <= r_n_74__29_;
      r_74__28_ <= r_n_74__28_;
      r_74__27_ <= r_n_74__27_;
      r_74__26_ <= r_n_74__26_;
      r_74__25_ <= r_n_74__25_;
      r_74__24_ <= r_n_74__24_;
      r_74__23_ <= r_n_74__23_;
      r_74__22_ <= r_n_74__22_;
      r_74__21_ <= r_n_74__21_;
      r_74__20_ <= r_n_74__20_;
      r_74__19_ <= r_n_74__19_;
      r_74__18_ <= r_n_74__18_;
      r_74__17_ <= r_n_74__17_;
      r_74__16_ <= r_n_74__16_;
      r_74__15_ <= r_n_74__15_;
      r_74__14_ <= r_n_74__14_;
      r_74__13_ <= r_n_74__13_;
      r_74__12_ <= r_n_74__12_;
      r_74__11_ <= r_n_74__11_;
      r_74__10_ <= r_n_74__10_;
      r_74__9_ <= r_n_74__9_;
      r_74__8_ <= r_n_74__8_;
      r_74__7_ <= r_n_74__7_;
      r_74__6_ <= r_n_74__6_;
      r_74__5_ <= r_n_74__5_;
      r_74__4_ <= r_n_74__4_;
      r_74__3_ <= r_n_74__3_;
      r_74__2_ <= r_n_74__2_;
      r_74__1_ <= r_n_74__1_;
      r_74__0_ <= r_n_74__0_;
    end 
    if(N1867) begin
      r_75__31_ <= r_n_75__31_;
      r_75__30_ <= r_n_75__30_;
      r_75__29_ <= r_n_75__29_;
      r_75__28_ <= r_n_75__28_;
      r_75__27_ <= r_n_75__27_;
      r_75__26_ <= r_n_75__26_;
      r_75__25_ <= r_n_75__25_;
      r_75__24_ <= r_n_75__24_;
      r_75__23_ <= r_n_75__23_;
      r_75__22_ <= r_n_75__22_;
      r_75__21_ <= r_n_75__21_;
      r_75__20_ <= r_n_75__20_;
      r_75__19_ <= r_n_75__19_;
      r_75__18_ <= r_n_75__18_;
      r_75__17_ <= r_n_75__17_;
      r_75__16_ <= r_n_75__16_;
      r_75__15_ <= r_n_75__15_;
      r_75__14_ <= r_n_75__14_;
      r_75__13_ <= r_n_75__13_;
      r_75__12_ <= r_n_75__12_;
      r_75__11_ <= r_n_75__11_;
      r_75__10_ <= r_n_75__10_;
      r_75__9_ <= r_n_75__9_;
      r_75__8_ <= r_n_75__8_;
      r_75__7_ <= r_n_75__7_;
      r_75__6_ <= r_n_75__6_;
      r_75__5_ <= r_n_75__5_;
      r_75__4_ <= r_n_75__4_;
      r_75__3_ <= r_n_75__3_;
      r_75__2_ <= r_n_75__2_;
      r_75__1_ <= r_n_75__1_;
      r_75__0_ <= r_n_75__0_;
    end 
    if(N1868) begin
      r_76__31_ <= r_n_76__31_;
      r_76__30_ <= r_n_76__30_;
      r_76__29_ <= r_n_76__29_;
      r_76__28_ <= r_n_76__28_;
      r_76__27_ <= r_n_76__27_;
      r_76__26_ <= r_n_76__26_;
      r_76__25_ <= r_n_76__25_;
      r_76__24_ <= r_n_76__24_;
      r_76__23_ <= r_n_76__23_;
      r_76__22_ <= r_n_76__22_;
      r_76__21_ <= r_n_76__21_;
      r_76__20_ <= r_n_76__20_;
      r_76__19_ <= r_n_76__19_;
      r_76__18_ <= r_n_76__18_;
      r_76__17_ <= r_n_76__17_;
      r_76__16_ <= r_n_76__16_;
      r_76__15_ <= r_n_76__15_;
      r_76__14_ <= r_n_76__14_;
      r_76__13_ <= r_n_76__13_;
      r_76__12_ <= r_n_76__12_;
      r_76__11_ <= r_n_76__11_;
      r_76__10_ <= r_n_76__10_;
      r_76__9_ <= r_n_76__9_;
      r_76__8_ <= r_n_76__8_;
      r_76__7_ <= r_n_76__7_;
      r_76__6_ <= r_n_76__6_;
      r_76__5_ <= r_n_76__5_;
      r_76__4_ <= r_n_76__4_;
      r_76__3_ <= r_n_76__3_;
      r_76__2_ <= r_n_76__2_;
      r_76__1_ <= r_n_76__1_;
      r_76__0_ <= r_n_76__0_;
    end 
    if(N1869) begin
      r_77__31_ <= r_n_77__31_;
      r_77__30_ <= r_n_77__30_;
      r_77__29_ <= r_n_77__29_;
      r_77__28_ <= r_n_77__28_;
      r_77__27_ <= r_n_77__27_;
      r_77__26_ <= r_n_77__26_;
      r_77__25_ <= r_n_77__25_;
      r_77__24_ <= r_n_77__24_;
      r_77__23_ <= r_n_77__23_;
      r_77__22_ <= r_n_77__22_;
      r_77__21_ <= r_n_77__21_;
      r_77__20_ <= r_n_77__20_;
      r_77__19_ <= r_n_77__19_;
      r_77__18_ <= r_n_77__18_;
      r_77__17_ <= r_n_77__17_;
      r_77__16_ <= r_n_77__16_;
      r_77__15_ <= r_n_77__15_;
      r_77__14_ <= r_n_77__14_;
      r_77__13_ <= r_n_77__13_;
      r_77__12_ <= r_n_77__12_;
      r_77__11_ <= r_n_77__11_;
      r_77__10_ <= r_n_77__10_;
      r_77__9_ <= r_n_77__9_;
      r_77__8_ <= r_n_77__8_;
      r_77__7_ <= r_n_77__7_;
      r_77__6_ <= r_n_77__6_;
      r_77__5_ <= r_n_77__5_;
      r_77__4_ <= r_n_77__4_;
      r_77__3_ <= r_n_77__3_;
      r_77__2_ <= r_n_77__2_;
      r_77__1_ <= r_n_77__1_;
      r_77__0_ <= r_n_77__0_;
    end 
    if(N1870) begin
      r_78__31_ <= r_n_78__31_;
      r_78__30_ <= r_n_78__30_;
      r_78__29_ <= r_n_78__29_;
      r_78__28_ <= r_n_78__28_;
      r_78__27_ <= r_n_78__27_;
      r_78__26_ <= r_n_78__26_;
      r_78__25_ <= r_n_78__25_;
      r_78__24_ <= r_n_78__24_;
      r_78__23_ <= r_n_78__23_;
      r_78__22_ <= r_n_78__22_;
      r_78__21_ <= r_n_78__21_;
      r_78__20_ <= r_n_78__20_;
      r_78__19_ <= r_n_78__19_;
      r_78__18_ <= r_n_78__18_;
      r_78__17_ <= r_n_78__17_;
      r_78__16_ <= r_n_78__16_;
      r_78__15_ <= r_n_78__15_;
      r_78__14_ <= r_n_78__14_;
      r_78__13_ <= r_n_78__13_;
      r_78__12_ <= r_n_78__12_;
      r_78__11_ <= r_n_78__11_;
      r_78__10_ <= r_n_78__10_;
      r_78__9_ <= r_n_78__9_;
      r_78__8_ <= r_n_78__8_;
      r_78__7_ <= r_n_78__7_;
      r_78__6_ <= r_n_78__6_;
      r_78__5_ <= r_n_78__5_;
      r_78__4_ <= r_n_78__4_;
      r_78__3_ <= r_n_78__3_;
      r_78__2_ <= r_n_78__2_;
      r_78__1_ <= r_n_78__1_;
      r_78__0_ <= r_n_78__0_;
    end 
    if(N1871) begin
      r_79__31_ <= r_n_79__31_;
      r_79__30_ <= r_n_79__30_;
      r_79__29_ <= r_n_79__29_;
      r_79__28_ <= r_n_79__28_;
      r_79__27_ <= r_n_79__27_;
      r_79__26_ <= r_n_79__26_;
      r_79__25_ <= r_n_79__25_;
      r_79__24_ <= r_n_79__24_;
      r_79__23_ <= r_n_79__23_;
      r_79__22_ <= r_n_79__22_;
      r_79__21_ <= r_n_79__21_;
      r_79__20_ <= r_n_79__20_;
      r_79__19_ <= r_n_79__19_;
      r_79__18_ <= r_n_79__18_;
      r_79__17_ <= r_n_79__17_;
      r_79__16_ <= r_n_79__16_;
      r_79__15_ <= r_n_79__15_;
      r_79__14_ <= r_n_79__14_;
      r_79__13_ <= r_n_79__13_;
      r_79__12_ <= r_n_79__12_;
      r_79__11_ <= r_n_79__11_;
      r_79__10_ <= r_n_79__10_;
      r_79__9_ <= r_n_79__9_;
      r_79__8_ <= r_n_79__8_;
      r_79__7_ <= r_n_79__7_;
      r_79__6_ <= r_n_79__6_;
      r_79__5_ <= r_n_79__5_;
      r_79__4_ <= r_n_79__4_;
      r_79__3_ <= r_n_79__3_;
      r_79__2_ <= r_n_79__2_;
      r_79__1_ <= r_n_79__1_;
      r_79__0_ <= r_n_79__0_;
    end 
    if(N1872) begin
      r_80__31_ <= r_n_80__31_;
      r_80__30_ <= r_n_80__30_;
      r_80__29_ <= r_n_80__29_;
      r_80__28_ <= r_n_80__28_;
      r_80__27_ <= r_n_80__27_;
      r_80__26_ <= r_n_80__26_;
      r_80__25_ <= r_n_80__25_;
      r_80__24_ <= r_n_80__24_;
      r_80__23_ <= r_n_80__23_;
      r_80__22_ <= r_n_80__22_;
      r_80__21_ <= r_n_80__21_;
      r_80__20_ <= r_n_80__20_;
      r_80__19_ <= r_n_80__19_;
      r_80__18_ <= r_n_80__18_;
      r_80__17_ <= r_n_80__17_;
      r_80__16_ <= r_n_80__16_;
      r_80__15_ <= r_n_80__15_;
      r_80__14_ <= r_n_80__14_;
      r_80__13_ <= r_n_80__13_;
      r_80__12_ <= r_n_80__12_;
      r_80__11_ <= r_n_80__11_;
      r_80__10_ <= r_n_80__10_;
      r_80__9_ <= r_n_80__9_;
      r_80__8_ <= r_n_80__8_;
      r_80__7_ <= r_n_80__7_;
      r_80__6_ <= r_n_80__6_;
      r_80__5_ <= r_n_80__5_;
      r_80__4_ <= r_n_80__4_;
      r_80__3_ <= r_n_80__3_;
      r_80__2_ <= r_n_80__2_;
      r_80__1_ <= r_n_80__1_;
      r_80__0_ <= r_n_80__0_;
    end 
    if(N1873) begin
      r_81__31_ <= r_n_81__31_;
      r_81__30_ <= r_n_81__30_;
      r_81__29_ <= r_n_81__29_;
      r_81__28_ <= r_n_81__28_;
      r_81__27_ <= r_n_81__27_;
      r_81__26_ <= r_n_81__26_;
      r_81__25_ <= r_n_81__25_;
      r_81__24_ <= r_n_81__24_;
      r_81__23_ <= r_n_81__23_;
      r_81__22_ <= r_n_81__22_;
      r_81__21_ <= r_n_81__21_;
      r_81__20_ <= r_n_81__20_;
      r_81__19_ <= r_n_81__19_;
      r_81__18_ <= r_n_81__18_;
      r_81__17_ <= r_n_81__17_;
      r_81__16_ <= r_n_81__16_;
      r_81__15_ <= r_n_81__15_;
      r_81__14_ <= r_n_81__14_;
      r_81__13_ <= r_n_81__13_;
      r_81__12_ <= r_n_81__12_;
      r_81__11_ <= r_n_81__11_;
      r_81__10_ <= r_n_81__10_;
      r_81__9_ <= r_n_81__9_;
      r_81__8_ <= r_n_81__8_;
      r_81__7_ <= r_n_81__7_;
      r_81__6_ <= r_n_81__6_;
      r_81__5_ <= r_n_81__5_;
      r_81__4_ <= r_n_81__4_;
      r_81__3_ <= r_n_81__3_;
      r_81__2_ <= r_n_81__2_;
      r_81__1_ <= r_n_81__1_;
      r_81__0_ <= r_n_81__0_;
    end 
    if(N1874) begin
      r_82__31_ <= r_n_82__31_;
      r_82__30_ <= r_n_82__30_;
      r_82__29_ <= r_n_82__29_;
      r_82__28_ <= r_n_82__28_;
      r_82__27_ <= r_n_82__27_;
      r_82__26_ <= r_n_82__26_;
      r_82__25_ <= r_n_82__25_;
      r_82__24_ <= r_n_82__24_;
      r_82__23_ <= r_n_82__23_;
      r_82__22_ <= r_n_82__22_;
      r_82__21_ <= r_n_82__21_;
      r_82__20_ <= r_n_82__20_;
      r_82__19_ <= r_n_82__19_;
      r_82__18_ <= r_n_82__18_;
      r_82__17_ <= r_n_82__17_;
      r_82__16_ <= r_n_82__16_;
      r_82__15_ <= r_n_82__15_;
      r_82__14_ <= r_n_82__14_;
      r_82__13_ <= r_n_82__13_;
      r_82__12_ <= r_n_82__12_;
      r_82__11_ <= r_n_82__11_;
      r_82__10_ <= r_n_82__10_;
      r_82__9_ <= r_n_82__9_;
      r_82__8_ <= r_n_82__8_;
      r_82__7_ <= r_n_82__7_;
      r_82__6_ <= r_n_82__6_;
      r_82__5_ <= r_n_82__5_;
      r_82__4_ <= r_n_82__4_;
      r_82__3_ <= r_n_82__3_;
      r_82__2_ <= r_n_82__2_;
      r_82__1_ <= r_n_82__1_;
      r_82__0_ <= r_n_82__0_;
    end 
    if(N1875) begin
      r_83__31_ <= r_n_83__31_;
      r_83__30_ <= r_n_83__30_;
      r_83__29_ <= r_n_83__29_;
      r_83__28_ <= r_n_83__28_;
      r_83__27_ <= r_n_83__27_;
      r_83__26_ <= r_n_83__26_;
      r_83__25_ <= r_n_83__25_;
      r_83__24_ <= r_n_83__24_;
      r_83__23_ <= r_n_83__23_;
      r_83__22_ <= r_n_83__22_;
      r_83__21_ <= r_n_83__21_;
      r_83__20_ <= r_n_83__20_;
      r_83__19_ <= r_n_83__19_;
      r_83__18_ <= r_n_83__18_;
      r_83__17_ <= r_n_83__17_;
      r_83__16_ <= r_n_83__16_;
      r_83__15_ <= r_n_83__15_;
      r_83__14_ <= r_n_83__14_;
      r_83__13_ <= r_n_83__13_;
      r_83__12_ <= r_n_83__12_;
      r_83__11_ <= r_n_83__11_;
      r_83__10_ <= r_n_83__10_;
      r_83__9_ <= r_n_83__9_;
      r_83__8_ <= r_n_83__8_;
      r_83__7_ <= r_n_83__7_;
      r_83__6_ <= r_n_83__6_;
      r_83__5_ <= r_n_83__5_;
      r_83__4_ <= r_n_83__4_;
      r_83__3_ <= r_n_83__3_;
      r_83__2_ <= r_n_83__2_;
      r_83__1_ <= r_n_83__1_;
      r_83__0_ <= r_n_83__0_;
    end 
    if(N1876) begin
      r_84__31_ <= r_n_84__31_;
      r_84__30_ <= r_n_84__30_;
      r_84__29_ <= r_n_84__29_;
      r_84__28_ <= r_n_84__28_;
      r_84__27_ <= r_n_84__27_;
      r_84__26_ <= r_n_84__26_;
      r_84__25_ <= r_n_84__25_;
      r_84__24_ <= r_n_84__24_;
      r_84__23_ <= r_n_84__23_;
      r_84__22_ <= r_n_84__22_;
      r_84__21_ <= r_n_84__21_;
      r_84__20_ <= r_n_84__20_;
      r_84__19_ <= r_n_84__19_;
      r_84__18_ <= r_n_84__18_;
      r_84__17_ <= r_n_84__17_;
      r_84__16_ <= r_n_84__16_;
      r_84__15_ <= r_n_84__15_;
      r_84__14_ <= r_n_84__14_;
      r_84__13_ <= r_n_84__13_;
      r_84__12_ <= r_n_84__12_;
      r_84__11_ <= r_n_84__11_;
      r_84__10_ <= r_n_84__10_;
      r_84__9_ <= r_n_84__9_;
      r_84__8_ <= r_n_84__8_;
      r_84__7_ <= r_n_84__7_;
      r_84__6_ <= r_n_84__6_;
      r_84__5_ <= r_n_84__5_;
      r_84__4_ <= r_n_84__4_;
      r_84__3_ <= r_n_84__3_;
      r_84__2_ <= r_n_84__2_;
      r_84__1_ <= r_n_84__1_;
      r_84__0_ <= r_n_84__0_;
    end 
    if(N1877) begin
      r_85__31_ <= r_n_85__31_;
      r_85__30_ <= r_n_85__30_;
      r_85__29_ <= r_n_85__29_;
      r_85__28_ <= r_n_85__28_;
      r_85__27_ <= r_n_85__27_;
      r_85__26_ <= r_n_85__26_;
      r_85__25_ <= r_n_85__25_;
      r_85__24_ <= r_n_85__24_;
      r_85__23_ <= r_n_85__23_;
      r_85__22_ <= r_n_85__22_;
      r_85__21_ <= r_n_85__21_;
      r_85__20_ <= r_n_85__20_;
      r_85__19_ <= r_n_85__19_;
      r_85__18_ <= r_n_85__18_;
      r_85__17_ <= r_n_85__17_;
      r_85__16_ <= r_n_85__16_;
      r_85__15_ <= r_n_85__15_;
      r_85__14_ <= r_n_85__14_;
      r_85__13_ <= r_n_85__13_;
      r_85__12_ <= r_n_85__12_;
      r_85__11_ <= r_n_85__11_;
      r_85__10_ <= r_n_85__10_;
      r_85__9_ <= r_n_85__9_;
      r_85__8_ <= r_n_85__8_;
      r_85__7_ <= r_n_85__7_;
      r_85__6_ <= r_n_85__6_;
      r_85__5_ <= r_n_85__5_;
      r_85__4_ <= r_n_85__4_;
      r_85__3_ <= r_n_85__3_;
      r_85__2_ <= r_n_85__2_;
      r_85__1_ <= r_n_85__1_;
      r_85__0_ <= r_n_85__0_;
    end 
    if(N1878) begin
      r_86__31_ <= r_n_86__31_;
      r_86__30_ <= r_n_86__30_;
      r_86__29_ <= r_n_86__29_;
      r_86__28_ <= r_n_86__28_;
      r_86__27_ <= r_n_86__27_;
      r_86__26_ <= r_n_86__26_;
      r_86__25_ <= r_n_86__25_;
      r_86__24_ <= r_n_86__24_;
      r_86__23_ <= r_n_86__23_;
      r_86__22_ <= r_n_86__22_;
      r_86__21_ <= r_n_86__21_;
      r_86__20_ <= r_n_86__20_;
      r_86__19_ <= r_n_86__19_;
      r_86__18_ <= r_n_86__18_;
      r_86__17_ <= r_n_86__17_;
      r_86__16_ <= r_n_86__16_;
      r_86__15_ <= r_n_86__15_;
      r_86__14_ <= r_n_86__14_;
      r_86__13_ <= r_n_86__13_;
      r_86__12_ <= r_n_86__12_;
      r_86__11_ <= r_n_86__11_;
      r_86__10_ <= r_n_86__10_;
      r_86__9_ <= r_n_86__9_;
      r_86__8_ <= r_n_86__8_;
      r_86__7_ <= r_n_86__7_;
      r_86__6_ <= r_n_86__6_;
      r_86__5_ <= r_n_86__5_;
      r_86__4_ <= r_n_86__4_;
      r_86__3_ <= r_n_86__3_;
      r_86__2_ <= r_n_86__2_;
      r_86__1_ <= r_n_86__1_;
      r_86__0_ <= r_n_86__0_;
    end 
    if(N1879) begin
      r_87__31_ <= r_n_87__31_;
      r_87__30_ <= r_n_87__30_;
      r_87__29_ <= r_n_87__29_;
      r_87__28_ <= r_n_87__28_;
      r_87__27_ <= r_n_87__27_;
      r_87__26_ <= r_n_87__26_;
      r_87__25_ <= r_n_87__25_;
      r_87__24_ <= r_n_87__24_;
      r_87__23_ <= r_n_87__23_;
      r_87__22_ <= r_n_87__22_;
      r_87__21_ <= r_n_87__21_;
      r_87__20_ <= r_n_87__20_;
      r_87__19_ <= r_n_87__19_;
      r_87__18_ <= r_n_87__18_;
      r_87__17_ <= r_n_87__17_;
      r_87__16_ <= r_n_87__16_;
      r_87__15_ <= r_n_87__15_;
      r_87__14_ <= r_n_87__14_;
      r_87__13_ <= r_n_87__13_;
      r_87__12_ <= r_n_87__12_;
      r_87__11_ <= r_n_87__11_;
      r_87__10_ <= r_n_87__10_;
      r_87__9_ <= r_n_87__9_;
      r_87__8_ <= r_n_87__8_;
      r_87__7_ <= r_n_87__7_;
      r_87__6_ <= r_n_87__6_;
      r_87__5_ <= r_n_87__5_;
      r_87__4_ <= r_n_87__4_;
      r_87__3_ <= r_n_87__3_;
      r_87__2_ <= r_n_87__2_;
      r_87__1_ <= r_n_87__1_;
      r_87__0_ <= r_n_87__0_;
    end 
    if(N1880) begin
      r_88__31_ <= r_n_88__31_;
      r_88__30_ <= r_n_88__30_;
      r_88__29_ <= r_n_88__29_;
      r_88__28_ <= r_n_88__28_;
      r_88__27_ <= r_n_88__27_;
      r_88__26_ <= r_n_88__26_;
      r_88__25_ <= r_n_88__25_;
      r_88__24_ <= r_n_88__24_;
      r_88__23_ <= r_n_88__23_;
      r_88__22_ <= r_n_88__22_;
      r_88__21_ <= r_n_88__21_;
      r_88__20_ <= r_n_88__20_;
      r_88__19_ <= r_n_88__19_;
      r_88__18_ <= r_n_88__18_;
      r_88__17_ <= r_n_88__17_;
      r_88__16_ <= r_n_88__16_;
      r_88__15_ <= r_n_88__15_;
      r_88__14_ <= r_n_88__14_;
      r_88__13_ <= r_n_88__13_;
      r_88__12_ <= r_n_88__12_;
      r_88__11_ <= r_n_88__11_;
      r_88__10_ <= r_n_88__10_;
      r_88__9_ <= r_n_88__9_;
      r_88__8_ <= r_n_88__8_;
      r_88__7_ <= r_n_88__7_;
      r_88__6_ <= r_n_88__6_;
      r_88__5_ <= r_n_88__5_;
      r_88__4_ <= r_n_88__4_;
      r_88__3_ <= r_n_88__3_;
      r_88__2_ <= r_n_88__2_;
      r_88__1_ <= r_n_88__1_;
      r_88__0_ <= r_n_88__0_;
    end 
    if(N1881) begin
      r_89__31_ <= r_n_89__31_;
      r_89__30_ <= r_n_89__30_;
      r_89__29_ <= r_n_89__29_;
      r_89__28_ <= r_n_89__28_;
      r_89__27_ <= r_n_89__27_;
      r_89__26_ <= r_n_89__26_;
      r_89__25_ <= r_n_89__25_;
      r_89__24_ <= r_n_89__24_;
      r_89__23_ <= r_n_89__23_;
      r_89__22_ <= r_n_89__22_;
      r_89__21_ <= r_n_89__21_;
      r_89__20_ <= r_n_89__20_;
      r_89__19_ <= r_n_89__19_;
      r_89__18_ <= r_n_89__18_;
      r_89__17_ <= r_n_89__17_;
      r_89__16_ <= r_n_89__16_;
      r_89__15_ <= r_n_89__15_;
      r_89__14_ <= r_n_89__14_;
      r_89__13_ <= r_n_89__13_;
      r_89__12_ <= r_n_89__12_;
      r_89__11_ <= r_n_89__11_;
      r_89__10_ <= r_n_89__10_;
      r_89__9_ <= r_n_89__9_;
      r_89__8_ <= r_n_89__8_;
      r_89__7_ <= r_n_89__7_;
      r_89__6_ <= r_n_89__6_;
      r_89__5_ <= r_n_89__5_;
      r_89__4_ <= r_n_89__4_;
      r_89__3_ <= r_n_89__3_;
      r_89__2_ <= r_n_89__2_;
      r_89__1_ <= r_n_89__1_;
      r_89__0_ <= r_n_89__0_;
    end 
    if(N1882) begin
      r_90__31_ <= r_n_90__31_;
      r_90__30_ <= r_n_90__30_;
      r_90__29_ <= r_n_90__29_;
      r_90__28_ <= r_n_90__28_;
      r_90__27_ <= r_n_90__27_;
      r_90__26_ <= r_n_90__26_;
      r_90__25_ <= r_n_90__25_;
      r_90__24_ <= r_n_90__24_;
      r_90__23_ <= r_n_90__23_;
      r_90__22_ <= r_n_90__22_;
      r_90__21_ <= r_n_90__21_;
      r_90__20_ <= r_n_90__20_;
      r_90__19_ <= r_n_90__19_;
      r_90__18_ <= r_n_90__18_;
      r_90__17_ <= r_n_90__17_;
      r_90__16_ <= r_n_90__16_;
      r_90__15_ <= r_n_90__15_;
      r_90__14_ <= r_n_90__14_;
      r_90__13_ <= r_n_90__13_;
      r_90__12_ <= r_n_90__12_;
      r_90__11_ <= r_n_90__11_;
      r_90__10_ <= r_n_90__10_;
      r_90__9_ <= r_n_90__9_;
      r_90__8_ <= r_n_90__8_;
      r_90__7_ <= r_n_90__7_;
      r_90__6_ <= r_n_90__6_;
      r_90__5_ <= r_n_90__5_;
      r_90__4_ <= r_n_90__4_;
      r_90__3_ <= r_n_90__3_;
      r_90__2_ <= r_n_90__2_;
      r_90__1_ <= r_n_90__1_;
      r_90__0_ <= r_n_90__0_;
    end 
    if(N1883) begin
      r_91__31_ <= r_n_91__31_;
      r_91__30_ <= r_n_91__30_;
      r_91__29_ <= r_n_91__29_;
      r_91__28_ <= r_n_91__28_;
      r_91__27_ <= r_n_91__27_;
      r_91__26_ <= r_n_91__26_;
      r_91__25_ <= r_n_91__25_;
      r_91__24_ <= r_n_91__24_;
      r_91__23_ <= r_n_91__23_;
      r_91__22_ <= r_n_91__22_;
      r_91__21_ <= r_n_91__21_;
      r_91__20_ <= r_n_91__20_;
      r_91__19_ <= r_n_91__19_;
      r_91__18_ <= r_n_91__18_;
      r_91__17_ <= r_n_91__17_;
      r_91__16_ <= r_n_91__16_;
      r_91__15_ <= r_n_91__15_;
      r_91__14_ <= r_n_91__14_;
      r_91__13_ <= r_n_91__13_;
      r_91__12_ <= r_n_91__12_;
      r_91__11_ <= r_n_91__11_;
      r_91__10_ <= r_n_91__10_;
      r_91__9_ <= r_n_91__9_;
      r_91__8_ <= r_n_91__8_;
      r_91__7_ <= r_n_91__7_;
      r_91__6_ <= r_n_91__6_;
      r_91__5_ <= r_n_91__5_;
      r_91__4_ <= r_n_91__4_;
      r_91__3_ <= r_n_91__3_;
      r_91__2_ <= r_n_91__2_;
      r_91__1_ <= r_n_91__1_;
      r_91__0_ <= r_n_91__0_;
    end 
    if(N1884) begin
      r_92__31_ <= r_n_92__31_;
      r_92__30_ <= r_n_92__30_;
      r_92__29_ <= r_n_92__29_;
      r_92__28_ <= r_n_92__28_;
      r_92__27_ <= r_n_92__27_;
      r_92__26_ <= r_n_92__26_;
      r_92__25_ <= r_n_92__25_;
      r_92__24_ <= r_n_92__24_;
      r_92__23_ <= r_n_92__23_;
      r_92__22_ <= r_n_92__22_;
      r_92__21_ <= r_n_92__21_;
      r_92__20_ <= r_n_92__20_;
      r_92__19_ <= r_n_92__19_;
      r_92__18_ <= r_n_92__18_;
      r_92__17_ <= r_n_92__17_;
      r_92__16_ <= r_n_92__16_;
      r_92__15_ <= r_n_92__15_;
      r_92__14_ <= r_n_92__14_;
      r_92__13_ <= r_n_92__13_;
      r_92__12_ <= r_n_92__12_;
      r_92__11_ <= r_n_92__11_;
      r_92__10_ <= r_n_92__10_;
      r_92__9_ <= r_n_92__9_;
      r_92__8_ <= r_n_92__8_;
      r_92__7_ <= r_n_92__7_;
      r_92__6_ <= r_n_92__6_;
      r_92__5_ <= r_n_92__5_;
      r_92__4_ <= r_n_92__4_;
      r_92__3_ <= r_n_92__3_;
      r_92__2_ <= r_n_92__2_;
      r_92__1_ <= r_n_92__1_;
      r_92__0_ <= r_n_92__0_;
    end 
    if(N1885) begin
      r_93__31_ <= r_n_93__31_;
      r_93__30_ <= r_n_93__30_;
      r_93__29_ <= r_n_93__29_;
      r_93__28_ <= r_n_93__28_;
      r_93__27_ <= r_n_93__27_;
      r_93__26_ <= r_n_93__26_;
      r_93__25_ <= r_n_93__25_;
      r_93__24_ <= r_n_93__24_;
      r_93__23_ <= r_n_93__23_;
      r_93__22_ <= r_n_93__22_;
      r_93__21_ <= r_n_93__21_;
      r_93__20_ <= r_n_93__20_;
      r_93__19_ <= r_n_93__19_;
      r_93__18_ <= r_n_93__18_;
      r_93__17_ <= r_n_93__17_;
      r_93__16_ <= r_n_93__16_;
      r_93__15_ <= r_n_93__15_;
      r_93__14_ <= r_n_93__14_;
      r_93__13_ <= r_n_93__13_;
      r_93__12_ <= r_n_93__12_;
      r_93__11_ <= r_n_93__11_;
      r_93__10_ <= r_n_93__10_;
      r_93__9_ <= r_n_93__9_;
      r_93__8_ <= r_n_93__8_;
      r_93__7_ <= r_n_93__7_;
      r_93__6_ <= r_n_93__6_;
      r_93__5_ <= r_n_93__5_;
      r_93__4_ <= r_n_93__4_;
      r_93__3_ <= r_n_93__3_;
      r_93__2_ <= r_n_93__2_;
      r_93__1_ <= r_n_93__1_;
      r_93__0_ <= r_n_93__0_;
    end 
    if(N1886) begin
      r_94__31_ <= r_n_94__31_;
      r_94__30_ <= r_n_94__30_;
      r_94__29_ <= r_n_94__29_;
      r_94__28_ <= r_n_94__28_;
      r_94__27_ <= r_n_94__27_;
      r_94__26_ <= r_n_94__26_;
      r_94__25_ <= r_n_94__25_;
      r_94__24_ <= r_n_94__24_;
      r_94__23_ <= r_n_94__23_;
      r_94__22_ <= r_n_94__22_;
      r_94__21_ <= r_n_94__21_;
      r_94__20_ <= r_n_94__20_;
      r_94__19_ <= r_n_94__19_;
      r_94__18_ <= r_n_94__18_;
      r_94__17_ <= r_n_94__17_;
      r_94__16_ <= r_n_94__16_;
      r_94__15_ <= r_n_94__15_;
      r_94__14_ <= r_n_94__14_;
      r_94__13_ <= r_n_94__13_;
      r_94__12_ <= r_n_94__12_;
      r_94__11_ <= r_n_94__11_;
      r_94__10_ <= r_n_94__10_;
      r_94__9_ <= r_n_94__9_;
      r_94__8_ <= r_n_94__8_;
      r_94__7_ <= r_n_94__7_;
      r_94__6_ <= r_n_94__6_;
      r_94__5_ <= r_n_94__5_;
      r_94__4_ <= r_n_94__4_;
      r_94__3_ <= r_n_94__3_;
      r_94__2_ <= r_n_94__2_;
      r_94__1_ <= r_n_94__1_;
      r_94__0_ <= r_n_94__0_;
    end 
    if(N1887) begin
      r_95__31_ <= r_n_95__31_;
      r_95__30_ <= r_n_95__30_;
      r_95__29_ <= r_n_95__29_;
      r_95__28_ <= r_n_95__28_;
      r_95__27_ <= r_n_95__27_;
      r_95__26_ <= r_n_95__26_;
      r_95__25_ <= r_n_95__25_;
      r_95__24_ <= r_n_95__24_;
      r_95__23_ <= r_n_95__23_;
      r_95__22_ <= r_n_95__22_;
      r_95__21_ <= r_n_95__21_;
      r_95__20_ <= r_n_95__20_;
      r_95__19_ <= r_n_95__19_;
      r_95__18_ <= r_n_95__18_;
      r_95__17_ <= r_n_95__17_;
      r_95__16_ <= r_n_95__16_;
      r_95__15_ <= r_n_95__15_;
      r_95__14_ <= r_n_95__14_;
      r_95__13_ <= r_n_95__13_;
      r_95__12_ <= r_n_95__12_;
      r_95__11_ <= r_n_95__11_;
      r_95__10_ <= r_n_95__10_;
      r_95__9_ <= r_n_95__9_;
      r_95__8_ <= r_n_95__8_;
      r_95__7_ <= r_n_95__7_;
      r_95__6_ <= r_n_95__6_;
      r_95__5_ <= r_n_95__5_;
      r_95__4_ <= r_n_95__4_;
      r_95__3_ <= r_n_95__3_;
      r_95__2_ <= r_n_95__2_;
      r_95__1_ <= r_n_95__1_;
      r_95__0_ <= r_n_95__0_;
    end 
    if(N1888) begin
      r_96__31_ <= r_n_96__31_;
      r_96__30_ <= r_n_96__30_;
      r_96__29_ <= r_n_96__29_;
      r_96__28_ <= r_n_96__28_;
      r_96__27_ <= r_n_96__27_;
      r_96__26_ <= r_n_96__26_;
      r_96__25_ <= r_n_96__25_;
      r_96__24_ <= r_n_96__24_;
      r_96__23_ <= r_n_96__23_;
      r_96__22_ <= r_n_96__22_;
      r_96__21_ <= r_n_96__21_;
      r_96__20_ <= r_n_96__20_;
      r_96__19_ <= r_n_96__19_;
      r_96__18_ <= r_n_96__18_;
      r_96__17_ <= r_n_96__17_;
      r_96__16_ <= r_n_96__16_;
      r_96__15_ <= r_n_96__15_;
      r_96__14_ <= r_n_96__14_;
      r_96__13_ <= r_n_96__13_;
      r_96__12_ <= r_n_96__12_;
      r_96__11_ <= r_n_96__11_;
      r_96__10_ <= r_n_96__10_;
      r_96__9_ <= r_n_96__9_;
      r_96__8_ <= r_n_96__8_;
      r_96__7_ <= r_n_96__7_;
      r_96__6_ <= r_n_96__6_;
      r_96__5_ <= r_n_96__5_;
      r_96__4_ <= r_n_96__4_;
      r_96__3_ <= r_n_96__3_;
      r_96__2_ <= r_n_96__2_;
      r_96__1_ <= r_n_96__1_;
      r_96__0_ <= r_n_96__0_;
    end 
    if(N1889) begin
      r_97__31_ <= r_n_97__31_;
      r_97__30_ <= r_n_97__30_;
      r_97__29_ <= r_n_97__29_;
      r_97__28_ <= r_n_97__28_;
      r_97__27_ <= r_n_97__27_;
      r_97__26_ <= r_n_97__26_;
      r_97__25_ <= r_n_97__25_;
      r_97__24_ <= r_n_97__24_;
      r_97__23_ <= r_n_97__23_;
      r_97__22_ <= r_n_97__22_;
      r_97__21_ <= r_n_97__21_;
      r_97__20_ <= r_n_97__20_;
      r_97__19_ <= r_n_97__19_;
      r_97__18_ <= r_n_97__18_;
      r_97__17_ <= r_n_97__17_;
      r_97__16_ <= r_n_97__16_;
      r_97__15_ <= r_n_97__15_;
      r_97__14_ <= r_n_97__14_;
      r_97__13_ <= r_n_97__13_;
      r_97__12_ <= r_n_97__12_;
      r_97__11_ <= r_n_97__11_;
      r_97__10_ <= r_n_97__10_;
      r_97__9_ <= r_n_97__9_;
      r_97__8_ <= r_n_97__8_;
      r_97__7_ <= r_n_97__7_;
      r_97__6_ <= r_n_97__6_;
      r_97__5_ <= r_n_97__5_;
      r_97__4_ <= r_n_97__4_;
      r_97__3_ <= r_n_97__3_;
      r_97__2_ <= r_n_97__2_;
      r_97__1_ <= r_n_97__1_;
      r_97__0_ <= r_n_97__0_;
    end 
    if(N1890) begin
      r_98__31_ <= r_n_98__31_;
      r_98__30_ <= r_n_98__30_;
      r_98__29_ <= r_n_98__29_;
      r_98__28_ <= r_n_98__28_;
      r_98__27_ <= r_n_98__27_;
      r_98__26_ <= r_n_98__26_;
      r_98__25_ <= r_n_98__25_;
      r_98__24_ <= r_n_98__24_;
      r_98__23_ <= r_n_98__23_;
      r_98__22_ <= r_n_98__22_;
      r_98__21_ <= r_n_98__21_;
      r_98__20_ <= r_n_98__20_;
      r_98__19_ <= r_n_98__19_;
      r_98__18_ <= r_n_98__18_;
      r_98__17_ <= r_n_98__17_;
      r_98__16_ <= r_n_98__16_;
      r_98__15_ <= r_n_98__15_;
      r_98__14_ <= r_n_98__14_;
      r_98__13_ <= r_n_98__13_;
      r_98__12_ <= r_n_98__12_;
      r_98__11_ <= r_n_98__11_;
      r_98__10_ <= r_n_98__10_;
      r_98__9_ <= r_n_98__9_;
      r_98__8_ <= r_n_98__8_;
      r_98__7_ <= r_n_98__7_;
      r_98__6_ <= r_n_98__6_;
      r_98__5_ <= r_n_98__5_;
      r_98__4_ <= r_n_98__4_;
      r_98__3_ <= r_n_98__3_;
      r_98__2_ <= r_n_98__2_;
      r_98__1_ <= r_n_98__1_;
      r_98__0_ <= r_n_98__0_;
    end 
    if(N1891) begin
      r_99__31_ <= r_n_99__31_;
      r_99__30_ <= r_n_99__30_;
      r_99__29_ <= r_n_99__29_;
      r_99__28_ <= r_n_99__28_;
      r_99__27_ <= r_n_99__27_;
      r_99__26_ <= r_n_99__26_;
      r_99__25_ <= r_n_99__25_;
      r_99__24_ <= r_n_99__24_;
      r_99__23_ <= r_n_99__23_;
      r_99__22_ <= r_n_99__22_;
      r_99__21_ <= r_n_99__21_;
      r_99__20_ <= r_n_99__20_;
      r_99__19_ <= r_n_99__19_;
      r_99__18_ <= r_n_99__18_;
      r_99__17_ <= r_n_99__17_;
      r_99__16_ <= r_n_99__16_;
      r_99__15_ <= r_n_99__15_;
      r_99__14_ <= r_n_99__14_;
      r_99__13_ <= r_n_99__13_;
      r_99__12_ <= r_n_99__12_;
      r_99__11_ <= r_n_99__11_;
      r_99__10_ <= r_n_99__10_;
      r_99__9_ <= r_n_99__9_;
      r_99__8_ <= r_n_99__8_;
      r_99__7_ <= r_n_99__7_;
      r_99__6_ <= r_n_99__6_;
      r_99__5_ <= r_n_99__5_;
      r_99__4_ <= r_n_99__4_;
      r_99__3_ <= r_n_99__3_;
      r_99__2_ <= r_n_99__2_;
      r_99__1_ <= r_n_99__1_;
      r_99__0_ <= r_n_99__0_;
    end 
    if(N1892) begin
      r_100__31_ <= r_n_100__31_;
      r_100__30_ <= r_n_100__30_;
      r_100__29_ <= r_n_100__29_;
      r_100__28_ <= r_n_100__28_;
      r_100__27_ <= r_n_100__27_;
      r_100__26_ <= r_n_100__26_;
      r_100__25_ <= r_n_100__25_;
      r_100__24_ <= r_n_100__24_;
      r_100__23_ <= r_n_100__23_;
      r_100__22_ <= r_n_100__22_;
      r_100__21_ <= r_n_100__21_;
      r_100__20_ <= r_n_100__20_;
      r_100__19_ <= r_n_100__19_;
      r_100__18_ <= r_n_100__18_;
      r_100__17_ <= r_n_100__17_;
      r_100__16_ <= r_n_100__16_;
      r_100__15_ <= r_n_100__15_;
      r_100__14_ <= r_n_100__14_;
      r_100__13_ <= r_n_100__13_;
      r_100__12_ <= r_n_100__12_;
      r_100__11_ <= r_n_100__11_;
      r_100__10_ <= r_n_100__10_;
      r_100__9_ <= r_n_100__9_;
      r_100__8_ <= r_n_100__8_;
      r_100__7_ <= r_n_100__7_;
      r_100__6_ <= r_n_100__6_;
      r_100__5_ <= r_n_100__5_;
      r_100__4_ <= r_n_100__4_;
      r_100__3_ <= r_n_100__3_;
      r_100__2_ <= r_n_100__2_;
      r_100__1_ <= r_n_100__1_;
      r_100__0_ <= r_n_100__0_;
    end 
    if(N1893) begin
      r_101__31_ <= r_n_101__31_;
      r_101__30_ <= r_n_101__30_;
      r_101__29_ <= r_n_101__29_;
      r_101__28_ <= r_n_101__28_;
      r_101__27_ <= r_n_101__27_;
      r_101__26_ <= r_n_101__26_;
      r_101__25_ <= r_n_101__25_;
      r_101__24_ <= r_n_101__24_;
      r_101__23_ <= r_n_101__23_;
      r_101__22_ <= r_n_101__22_;
      r_101__21_ <= r_n_101__21_;
      r_101__20_ <= r_n_101__20_;
      r_101__19_ <= r_n_101__19_;
      r_101__18_ <= r_n_101__18_;
      r_101__17_ <= r_n_101__17_;
      r_101__16_ <= r_n_101__16_;
      r_101__15_ <= r_n_101__15_;
      r_101__14_ <= r_n_101__14_;
      r_101__13_ <= r_n_101__13_;
      r_101__12_ <= r_n_101__12_;
      r_101__11_ <= r_n_101__11_;
      r_101__10_ <= r_n_101__10_;
      r_101__9_ <= r_n_101__9_;
      r_101__8_ <= r_n_101__8_;
      r_101__7_ <= r_n_101__7_;
      r_101__6_ <= r_n_101__6_;
      r_101__5_ <= r_n_101__5_;
      r_101__4_ <= r_n_101__4_;
      r_101__3_ <= r_n_101__3_;
      r_101__2_ <= r_n_101__2_;
      r_101__1_ <= r_n_101__1_;
      r_101__0_ <= r_n_101__0_;
    end 
    if(N1894) begin
      r_102__31_ <= r_n_102__31_;
      r_102__30_ <= r_n_102__30_;
      r_102__29_ <= r_n_102__29_;
      r_102__28_ <= r_n_102__28_;
      r_102__27_ <= r_n_102__27_;
      r_102__26_ <= r_n_102__26_;
      r_102__25_ <= r_n_102__25_;
      r_102__24_ <= r_n_102__24_;
      r_102__23_ <= r_n_102__23_;
      r_102__22_ <= r_n_102__22_;
      r_102__21_ <= r_n_102__21_;
      r_102__20_ <= r_n_102__20_;
      r_102__19_ <= r_n_102__19_;
      r_102__18_ <= r_n_102__18_;
      r_102__17_ <= r_n_102__17_;
      r_102__16_ <= r_n_102__16_;
      r_102__15_ <= r_n_102__15_;
      r_102__14_ <= r_n_102__14_;
      r_102__13_ <= r_n_102__13_;
      r_102__12_ <= r_n_102__12_;
      r_102__11_ <= r_n_102__11_;
      r_102__10_ <= r_n_102__10_;
      r_102__9_ <= r_n_102__9_;
      r_102__8_ <= r_n_102__8_;
      r_102__7_ <= r_n_102__7_;
      r_102__6_ <= r_n_102__6_;
      r_102__5_ <= r_n_102__5_;
      r_102__4_ <= r_n_102__4_;
      r_102__3_ <= r_n_102__3_;
      r_102__2_ <= r_n_102__2_;
      r_102__1_ <= r_n_102__1_;
      r_102__0_ <= r_n_102__0_;
    end 
    if(N1895) begin
      r_103__31_ <= r_n_103__31_;
      r_103__30_ <= r_n_103__30_;
      r_103__29_ <= r_n_103__29_;
      r_103__28_ <= r_n_103__28_;
      r_103__27_ <= r_n_103__27_;
      r_103__26_ <= r_n_103__26_;
      r_103__25_ <= r_n_103__25_;
      r_103__24_ <= r_n_103__24_;
      r_103__23_ <= r_n_103__23_;
      r_103__22_ <= r_n_103__22_;
      r_103__21_ <= r_n_103__21_;
      r_103__20_ <= r_n_103__20_;
      r_103__19_ <= r_n_103__19_;
      r_103__18_ <= r_n_103__18_;
      r_103__17_ <= r_n_103__17_;
      r_103__16_ <= r_n_103__16_;
      r_103__15_ <= r_n_103__15_;
      r_103__14_ <= r_n_103__14_;
      r_103__13_ <= r_n_103__13_;
      r_103__12_ <= r_n_103__12_;
      r_103__11_ <= r_n_103__11_;
      r_103__10_ <= r_n_103__10_;
      r_103__9_ <= r_n_103__9_;
      r_103__8_ <= r_n_103__8_;
      r_103__7_ <= r_n_103__7_;
      r_103__6_ <= r_n_103__6_;
      r_103__5_ <= r_n_103__5_;
      r_103__4_ <= r_n_103__4_;
      r_103__3_ <= r_n_103__3_;
      r_103__2_ <= r_n_103__2_;
      r_103__1_ <= r_n_103__1_;
      r_103__0_ <= r_n_103__0_;
    end 
    if(N1896) begin
      r_104__31_ <= r_n_104__31_;
      r_104__30_ <= r_n_104__30_;
      r_104__29_ <= r_n_104__29_;
      r_104__28_ <= r_n_104__28_;
      r_104__27_ <= r_n_104__27_;
      r_104__26_ <= r_n_104__26_;
      r_104__25_ <= r_n_104__25_;
      r_104__24_ <= r_n_104__24_;
      r_104__23_ <= r_n_104__23_;
      r_104__22_ <= r_n_104__22_;
      r_104__21_ <= r_n_104__21_;
      r_104__20_ <= r_n_104__20_;
      r_104__19_ <= r_n_104__19_;
      r_104__18_ <= r_n_104__18_;
      r_104__17_ <= r_n_104__17_;
      r_104__16_ <= r_n_104__16_;
      r_104__15_ <= r_n_104__15_;
      r_104__14_ <= r_n_104__14_;
      r_104__13_ <= r_n_104__13_;
      r_104__12_ <= r_n_104__12_;
      r_104__11_ <= r_n_104__11_;
      r_104__10_ <= r_n_104__10_;
      r_104__9_ <= r_n_104__9_;
      r_104__8_ <= r_n_104__8_;
      r_104__7_ <= r_n_104__7_;
      r_104__6_ <= r_n_104__6_;
      r_104__5_ <= r_n_104__5_;
      r_104__4_ <= r_n_104__4_;
      r_104__3_ <= r_n_104__3_;
      r_104__2_ <= r_n_104__2_;
      r_104__1_ <= r_n_104__1_;
      r_104__0_ <= r_n_104__0_;
    end 
    if(N1897) begin
      r_105__31_ <= r_n_105__31_;
      r_105__30_ <= r_n_105__30_;
      r_105__29_ <= r_n_105__29_;
      r_105__28_ <= r_n_105__28_;
      r_105__27_ <= r_n_105__27_;
      r_105__26_ <= r_n_105__26_;
      r_105__25_ <= r_n_105__25_;
      r_105__24_ <= r_n_105__24_;
      r_105__23_ <= r_n_105__23_;
      r_105__22_ <= r_n_105__22_;
      r_105__21_ <= r_n_105__21_;
      r_105__20_ <= r_n_105__20_;
      r_105__19_ <= r_n_105__19_;
      r_105__18_ <= r_n_105__18_;
      r_105__17_ <= r_n_105__17_;
      r_105__16_ <= r_n_105__16_;
      r_105__15_ <= r_n_105__15_;
      r_105__14_ <= r_n_105__14_;
      r_105__13_ <= r_n_105__13_;
      r_105__12_ <= r_n_105__12_;
      r_105__11_ <= r_n_105__11_;
      r_105__10_ <= r_n_105__10_;
      r_105__9_ <= r_n_105__9_;
      r_105__8_ <= r_n_105__8_;
      r_105__7_ <= r_n_105__7_;
      r_105__6_ <= r_n_105__6_;
      r_105__5_ <= r_n_105__5_;
      r_105__4_ <= r_n_105__4_;
      r_105__3_ <= r_n_105__3_;
      r_105__2_ <= r_n_105__2_;
      r_105__1_ <= r_n_105__1_;
      r_105__0_ <= r_n_105__0_;
    end 
    if(N1898) begin
      r_106__31_ <= r_n_106__31_;
      r_106__30_ <= r_n_106__30_;
      r_106__29_ <= r_n_106__29_;
      r_106__28_ <= r_n_106__28_;
      r_106__27_ <= r_n_106__27_;
      r_106__26_ <= r_n_106__26_;
      r_106__25_ <= r_n_106__25_;
      r_106__24_ <= r_n_106__24_;
      r_106__23_ <= r_n_106__23_;
      r_106__22_ <= r_n_106__22_;
      r_106__21_ <= r_n_106__21_;
      r_106__20_ <= r_n_106__20_;
      r_106__19_ <= r_n_106__19_;
      r_106__18_ <= r_n_106__18_;
      r_106__17_ <= r_n_106__17_;
      r_106__16_ <= r_n_106__16_;
      r_106__15_ <= r_n_106__15_;
      r_106__14_ <= r_n_106__14_;
      r_106__13_ <= r_n_106__13_;
      r_106__12_ <= r_n_106__12_;
      r_106__11_ <= r_n_106__11_;
      r_106__10_ <= r_n_106__10_;
      r_106__9_ <= r_n_106__9_;
      r_106__8_ <= r_n_106__8_;
      r_106__7_ <= r_n_106__7_;
      r_106__6_ <= r_n_106__6_;
      r_106__5_ <= r_n_106__5_;
      r_106__4_ <= r_n_106__4_;
      r_106__3_ <= r_n_106__3_;
      r_106__2_ <= r_n_106__2_;
      r_106__1_ <= r_n_106__1_;
      r_106__0_ <= r_n_106__0_;
    end 
    if(N1899) begin
      r_107__31_ <= r_n_107__31_;
      r_107__30_ <= r_n_107__30_;
      r_107__29_ <= r_n_107__29_;
      r_107__28_ <= r_n_107__28_;
      r_107__27_ <= r_n_107__27_;
      r_107__26_ <= r_n_107__26_;
      r_107__25_ <= r_n_107__25_;
      r_107__24_ <= r_n_107__24_;
      r_107__23_ <= r_n_107__23_;
      r_107__22_ <= r_n_107__22_;
      r_107__21_ <= r_n_107__21_;
      r_107__20_ <= r_n_107__20_;
      r_107__19_ <= r_n_107__19_;
      r_107__18_ <= r_n_107__18_;
      r_107__17_ <= r_n_107__17_;
      r_107__16_ <= r_n_107__16_;
      r_107__15_ <= r_n_107__15_;
      r_107__14_ <= r_n_107__14_;
      r_107__13_ <= r_n_107__13_;
      r_107__12_ <= r_n_107__12_;
      r_107__11_ <= r_n_107__11_;
      r_107__10_ <= r_n_107__10_;
      r_107__9_ <= r_n_107__9_;
      r_107__8_ <= r_n_107__8_;
      r_107__7_ <= r_n_107__7_;
      r_107__6_ <= r_n_107__6_;
      r_107__5_ <= r_n_107__5_;
      r_107__4_ <= r_n_107__4_;
      r_107__3_ <= r_n_107__3_;
      r_107__2_ <= r_n_107__2_;
      r_107__1_ <= r_n_107__1_;
      r_107__0_ <= r_n_107__0_;
    end 
    if(N1900) begin
      r_108__31_ <= r_n_108__31_;
      r_108__30_ <= r_n_108__30_;
      r_108__29_ <= r_n_108__29_;
      r_108__28_ <= r_n_108__28_;
      r_108__27_ <= r_n_108__27_;
      r_108__26_ <= r_n_108__26_;
      r_108__25_ <= r_n_108__25_;
      r_108__24_ <= r_n_108__24_;
      r_108__23_ <= r_n_108__23_;
      r_108__22_ <= r_n_108__22_;
      r_108__21_ <= r_n_108__21_;
      r_108__20_ <= r_n_108__20_;
      r_108__19_ <= r_n_108__19_;
      r_108__18_ <= r_n_108__18_;
      r_108__17_ <= r_n_108__17_;
      r_108__16_ <= r_n_108__16_;
      r_108__15_ <= r_n_108__15_;
      r_108__14_ <= r_n_108__14_;
      r_108__13_ <= r_n_108__13_;
      r_108__12_ <= r_n_108__12_;
      r_108__11_ <= r_n_108__11_;
      r_108__10_ <= r_n_108__10_;
      r_108__9_ <= r_n_108__9_;
      r_108__8_ <= r_n_108__8_;
      r_108__7_ <= r_n_108__7_;
      r_108__6_ <= r_n_108__6_;
      r_108__5_ <= r_n_108__5_;
      r_108__4_ <= r_n_108__4_;
      r_108__3_ <= r_n_108__3_;
      r_108__2_ <= r_n_108__2_;
      r_108__1_ <= r_n_108__1_;
      r_108__0_ <= r_n_108__0_;
    end 
    if(N1901) begin
      r_109__31_ <= r_n_109__31_;
      r_109__30_ <= r_n_109__30_;
      r_109__29_ <= r_n_109__29_;
      r_109__28_ <= r_n_109__28_;
      r_109__27_ <= r_n_109__27_;
      r_109__26_ <= r_n_109__26_;
      r_109__25_ <= r_n_109__25_;
      r_109__24_ <= r_n_109__24_;
      r_109__23_ <= r_n_109__23_;
      r_109__22_ <= r_n_109__22_;
      r_109__21_ <= r_n_109__21_;
      r_109__20_ <= r_n_109__20_;
      r_109__19_ <= r_n_109__19_;
      r_109__18_ <= r_n_109__18_;
      r_109__17_ <= r_n_109__17_;
      r_109__16_ <= r_n_109__16_;
      r_109__15_ <= r_n_109__15_;
      r_109__14_ <= r_n_109__14_;
      r_109__13_ <= r_n_109__13_;
      r_109__12_ <= r_n_109__12_;
      r_109__11_ <= r_n_109__11_;
      r_109__10_ <= r_n_109__10_;
      r_109__9_ <= r_n_109__9_;
      r_109__8_ <= r_n_109__8_;
      r_109__7_ <= r_n_109__7_;
      r_109__6_ <= r_n_109__6_;
      r_109__5_ <= r_n_109__5_;
      r_109__4_ <= r_n_109__4_;
      r_109__3_ <= r_n_109__3_;
      r_109__2_ <= r_n_109__2_;
      r_109__1_ <= r_n_109__1_;
      r_109__0_ <= r_n_109__0_;
    end 
    if(N1902) begin
      r_110__31_ <= r_n_110__31_;
      r_110__30_ <= r_n_110__30_;
      r_110__29_ <= r_n_110__29_;
      r_110__28_ <= r_n_110__28_;
      r_110__27_ <= r_n_110__27_;
      r_110__26_ <= r_n_110__26_;
      r_110__25_ <= r_n_110__25_;
      r_110__24_ <= r_n_110__24_;
      r_110__23_ <= r_n_110__23_;
      r_110__22_ <= r_n_110__22_;
      r_110__21_ <= r_n_110__21_;
      r_110__20_ <= r_n_110__20_;
      r_110__19_ <= r_n_110__19_;
      r_110__18_ <= r_n_110__18_;
      r_110__17_ <= r_n_110__17_;
      r_110__16_ <= r_n_110__16_;
      r_110__15_ <= r_n_110__15_;
      r_110__14_ <= r_n_110__14_;
      r_110__13_ <= r_n_110__13_;
      r_110__12_ <= r_n_110__12_;
      r_110__11_ <= r_n_110__11_;
      r_110__10_ <= r_n_110__10_;
      r_110__9_ <= r_n_110__9_;
      r_110__8_ <= r_n_110__8_;
      r_110__7_ <= r_n_110__7_;
      r_110__6_ <= r_n_110__6_;
      r_110__5_ <= r_n_110__5_;
      r_110__4_ <= r_n_110__4_;
      r_110__3_ <= r_n_110__3_;
      r_110__2_ <= r_n_110__2_;
      r_110__1_ <= r_n_110__1_;
      r_110__0_ <= r_n_110__0_;
    end 
    if(N1903) begin
      r_111__31_ <= r_n_111__31_;
      r_111__30_ <= r_n_111__30_;
      r_111__29_ <= r_n_111__29_;
      r_111__28_ <= r_n_111__28_;
      r_111__27_ <= r_n_111__27_;
      r_111__26_ <= r_n_111__26_;
      r_111__25_ <= r_n_111__25_;
      r_111__24_ <= r_n_111__24_;
      r_111__23_ <= r_n_111__23_;
      r_111__22_ <= r_n_111__22_;
      r_111__21_ <= r_n_111__21_;
      r_111__20_ <= r_n_111__20_;
      r_111__19_ <= r_n_111__19_;
      r_111__18_ <= r_n_111__18_;
      r_111__17_ <= r_n_111__17_;
      r_111__16_ <= r_n_111__16_;
      r_111__15_ <= r_n_111__15_;
      r_111__14_ <= r_n_111__14_;
      r_111__13_ <= r_n_111__13_;
      r_111__12_ <= r_n_111__12_;
      r_111__11_ <= r_n_111__11_;
      r_111__10_ <= r_n_111__10_;
      r_111__9_ <= r_n_111__9_;
      r_111__8_ <= r_n_111__8_;
      r_111__7_ <= r_n_111__7_;
      r_111__6_ <= r_n_111__6_;
      r_111__5_ <= r_n_111__5_;
      r_111__4_ <= r_n_111__4_;
      r_111__3_ <= r_n_111__3_;
      r_111__2_ <= r_n_111__2_;
      r_111__1_ <= r_n_111__1_;
      r_111__0_ <= r_n_111__0_;
    end 
    if(N1904) begin
      r_112__31_ <= r_n_112__31_;
      r_112__30_ <= r_n_112__30_;
      r_112__29_ <= r_n_112__29_;
      r_112__28_ <= r_n_112__28_;
      r_112__27_ <= r_n_112__27_;
      r_112__26_ <= r_n_112__26_;
      r_112__25_ <= r_n_112__25_;
      r_112__24_ <= r_n_112__24_;
      r_112__23_ <= r_n_112__23_;
      r_112__22_ <= r_n_112__22_;
      r_112__21_ <= r_n_112__21_;
      r_112__20_ <= r_n_112__20_;
      r_112__19_ <= r_n_112__19_;
      r_112__18_ <= r_n_112__18_;
      r_112__17_ <= r_n_112__17_;
      r_112__16_ <= r_n_112__16_;
      r_112__15_ <= r_n_112__15_;
      r_112__14_ <= r_n_112__14_;
      r_112__13_ <= r_n_112__13_;
      r_112__12_ <= r_n_112__12_;
      r_112__11_ <= r_n_112__11_;
      r_112__10_ <= r_n_112__10_;
      r_112__9_ <= r_n_112__9_;
      r_112__8_ <= r_n_112__8_;
      r_112__7_ <= r_n_112__7_;
      r_112__6_ <= r_n_112__6_;
      r_112__5_ <= r_n_112__5_;
      r_112__4_ <= r_n_112__4_;
      r_112__3_ <= r_n_112__3_;
      r_112__2_ <= r_n_112__2_;
      r_112__1_ <= r_n_112__1_;
      r_112__0_ <= r_n_112__0_;
    end 
    if(N1905) begin
      r_113__31_ <= r_n_113__31_;
      r_113__30_ <= r_n_113__30_;
      r_113__29_ <= r_n_113__29_;
      r_113__28_ <= r_n_113__28_;
      r_113__27_ <= r_n_113__27_;
      r_113__26_ <= r_n_113__26_;
      r_113__25_ <= r_n_113__25_;
      r_113__24_ <= r_n_113__24_;
      r_113__23_ <= r_n_113__23_;
      r_113__22_ <= r_n_113__22_;
      r_113__21_ <= r_n_113__21_;
      r_113__20_ <= r_n_113__20_;
      r_113__19_ <= r_n_113__19_;
      r_113__18_ <= r_n_113__18_;
      r_113__17_ <= r_n_113__17_;
      r_113__16_ <= r_n_113__16_;
      r_113__15_ <= r_n_113__15_;
      r_113__14_ <= r_n_113__14_;
      r_113__13_ <= r_n_113__13_;
      r_113__12_ <= r_n_113__12_;
      r_113__11_ <= r_n_113__11_;
      r_113__10_ <= r_n_113__10_;
      r_113__9_ <= r_n_113__9_;
      r_113__8_ <= r_n_113__8_;
      r_113__7_ <= r_n_113__7_;
      r_113__6_ <= r_n_113__6_;
      r_113__5_ <= r_n_113__5_;
      r_113__4_ <= r_n_113__4_;
      r_113__3_ <= r_n_113__3_;
      r_113__2_ <= r_n_113__2_;
      r_113__1_ <= r_n_113__1_;
      r_113__0_ <= r_n_113__0_;
    end 
    if(N1906) begin
      r_114__31_ <= r_n_114__31_;
      r_114__30_ <= r_n_114__30_;
      r_114__29_ <= r_n_114__29_;
      r_114__28_ <= r_n_114__28_;
      r_114__27_ <= r_n_114__27_;
      r_114__26_ <= r_n_114__26_;
      r_114__25_ <= r_n_114__25_;
      r_114__24_ <= r_n_114__24_;
      r_114__23_ <= r_n_114__23_;
      r_114__22_ <= r_n_114__22_;
      r_114__21_ <= r_n_114__21_;
      r_114__20_ <= r_n_114__20_;
      r_114__19_ <= r_n_114__19_;
      r_114__18_ <= r_n_114__18_;
      r_114__17_ <= r_n_114__17_;
      r_114__16_ <= r_n_114__16_;
      r_114__15_ <= r_n_114__15_;
      r_114__14_ <= r_n_114__14_;
      r_114__13_ <= r_n_114__13_;
      r_114__12_ <= r_n_114__12_;
      r_114__11_ <= r_n_114__11_;
      r_114__10_ <= r_n_114__10_;
      r_114__9_ <= r_n_114__9_;
      r_114__8_ <= r_n_114__8_;
      r_114__7_ <= r_n_114__7_;
      r_114__6_ <= r_n_114__6_;
      r_114__5_ <= r_n_114__5_;
      r_114__4_ <= r_n_114__4_;
      r_114__3_ <= r_n_114__3_;
      r_114__2_ <= r_n_114__2_;
      r_114__1_ <= r_n_114__1_;
      r_114__0_ <= r_n_114__0_;
    end 
    if(N1907) begin
      r_115__31_ <= r_n_115__31_;
      r_115__30_ <= r_n_115__30_;
      r_115__29_ <= r_n_115__29_;
      r_115__28_ <= r_n_115__28_;
      r_115__27_ <= r_n_115__27_;
      r_115__26_ <= r_n_115__26_;
      r_115__25_ <= r_n_115__25_;
      r_115__24_ <= r_n_115__24_;
      r_115__23_ <= r_n_115__23_;
      r_115__22_ <= r_n_115__22_;
      r_115__21_ <= r_n_115__21_;
      r_115__20_ <= r_n_115__20_;
      r_115__19_ <= r_n_115__19_;
      r_115__18_ <= r_n_115__18_;
      r_115__17_ <= r_n_115__17_;
      r_115__16_ <= r_n_115__16_;
      r_115__15_ <= r_n_115__15_;
      r_115__14_ <= r_n_115__14_;
      r_115__13_ <= r_n_115__13_;
      r_115__12_ <= r_n_115__12_;
      r_115__11_ <= r_n_115__11_;
      r_115__10_ <= r_n_115__10_;
      r_115__9_ <= r_n_115__9_;
      r_115__8_ <= r_n_115__8_;
      r_115__7_ <= r_n_115__7_;
      r_115__6_ <= r_n_115__6_;
      r_115__5_ <= r_n_115__5_;
      r_115__4_ <= r_n_115__4_;
      r_115__3_ <= r_n_115__3_;
      r_115__2_ <= r_n_115__2_;
      r_115__1_ <= r_n_115__1_;
      r_115__0_ <= r_n_115__0_;
    end 
    if(N1908) begin
      r_116__31_ <= r_n_116__31_;
      r_116__30_ <= r_n_116__30_;
      r_116__29_ <= r_n_116__29_;
      r_116__28_ <= r_n_116__28_;
      r_116__27_ <= r_n_116__27_;
      r_116__26_ <= r_n_116__26_;
      r_116__25_ <= r_n_116__25_;
      r_116__24_ <= r_n_116__24_;
      r_116__23_ <= r_n_116__23_;
      r_116__22_ <= r_n_116__22_;
      r_116__21_ <= r_n_116__21_;
      r_116__20_ <= r_n_116__20_;
      r_116__19_ <= r_n_116__19_;
      r_116__18_ <= r_n_116__18_;
      r_116__17_ <= r_n_116__17_;
      r_116__16_ <= r_n_116__16_;
      r_116__15_ <= r_n_116__15_;
      r_116__14_ <= r_n_116__14_;
      r_116__13_ <= r_n_116__13_;
      r_116__12_ <= r_n_116__12_;
      r_116__11_ <= r_n_116__11_;
      r_116__10_ <= r_n_116__10_;
      r_116__9_ <= r_n_116__9_;
      r_116__8_ <= r_n_116__8_;
      r_116__7_ <= r_n_116__7_;
      r_116__6_ <= r_n_116__6_;
      r_116__5_ <= r_n_116__5_;
      r_116__4_ <= r_n_116__4_;
      r_116__3_ <= r_n_116__3_;
      r_116__2_ <= r_n_116__2_;
      r_116__1_ <= r_n_116__1_;
      r_116__0_ <= r_n_116__0_;
    end 
    if(N1909) begin
      r_117__31_ <= r_n_117__31_;
      r_117__30_ <= r_n_117__30_;
      r_117__29_ <= r_n_117__29_;
      r_117__28_ <= r_n_117__28_;
      r_117__27_ <= r_n_117__27_;
      r_117__26_ <= r_n_117__26_;
      r_117__25_ <= r_n_117__25_;
      r_117__24_ <= r_n_117__24_;
      r_117__23_ <= r_n_117__23_;
      r_117__22_ <= r_n_117__22_;
      r_117__21_ <= r_n_117__21_;
      r_117__20_ <= r_n_117__20_;
      r_117__19_ <= r_n_117__19_;
      r_117__18_ <= r_n_117__18_;
      r_117__17_ <= r_n_117__17_;
      r_117__16_ <= r_n_117__16_;
      r_117__15_ <= r_n_117__15_;
      r_117__14_ <= r_n_117__14_;
      r_117__13_ <= r_n_117__13_;
      r_117__12_ <= r_n_117__12_;
      r_117__11_ <= r_n_117__11_;
      r_117__10_ <= r_n_117__10_;
      r_117__9_ <= r_n_117__9_;
      r_117__8_ <= r_n_117__8_;
      r_117__7_ <= r_n_117__7_;
      r_117__6_ <= r_n_117__6_;
      r_117__5_ <= r_n_117__5_;
      r_117__4_ <= r_n_117__4_;
      r_117__3_ <= r_n_117__3_;
      r_117__2_ <= r_n_117__2_;
      r_117__1_ <= r_n_117__1_;
      r_117__0_ <= r_n_117__0_;
    end 
    if(N1910) begin
      r_118__31_ <= r_n_118__31_;
      r_118__30_ <= r_n_118__30_;
      r_118__29_ <= r_n_118__29_;
      r_118__28_ <= r_n_118__28_;
      r_118__27_ <= r_n_118__27_;
      r_118__26_ <= r_n_118__26_;
      r_118__25_ <= r_n_118__25_;
      r_118__24_ <= r_n_118__24_;
      r_118__23_ <= r_n_118__23_;
      r_118__22_ <= r_n_118__22_;
      r_118__21_ <= r_n_118__21_;
      r_118__20_ <= r_n_118__20_;
      r_118__19_ <= r_n_118__19_;
      r_118__18_ <= r_n_118__18_;
      r_118__17_ <= r_n_118__17_;
      r_118__16_ <= r_n_118__16_;
      r_118__15_ <= r_n_118__15_;
      r_118__14_ <= r_n_118__14_;
      r_118__13_ <= r_n_118__13_;
      r_118__12_ <= r_n_118__12_;
      r_118__11_ <= r_n_118__11_;
      r_118__10_ <= r_n_118__10_;
      r_118__9_ <= r_n_118__9_;
      r_118__8_ <= r_n_118__8_;
      r_118__7_ <= r_n_118__7_;
      r_118__6_ <= r_n_118__6_;
      r_118__5_ <= r_n_118__5_;
      r_118__4_ <= r_n_118__4_;
      r_118__3_ <= r_n_118__3_;
      r_118__2_ <= r_n_118__2_;
      r_118__1_ <= r_n_118__1_;
      r_118__0_ <= r_n_118__0_;
    end 
    if(N1911) begin
      r_119__31_ <= r_n_119__31_;
      r_119__30_ <= r_n_119__30_;
      r_119__29_ <= r_n_119__29_;
      r_119__28_ <= r_n_119__28_;
      r_119__27_ <= r_n_119__27_;
      r_119__26_ <= r_n_119__26_;
      r_119__25_ <= r_n_119__25_;
      r_119__24_ <= r_n_119__24_;
      r_119__23_ <= r_n_119__23_;
      r_119__22_ <= r_n_119__22_;
      r_119__21_ <= r_n_119__21_;
      r_119__20_ <= r_n_119__20_;
      r_119__19_ <= r_n_119__19_;
      r_119__18_ <= r_n_119__18_;
      r_119__17_ <= r_n_119__17_;
      r_119__16_ <= r_n_119__16_;
      r_119__15_ <= r_n_119__15_;
      r_119__14_ <= r_n_119__14_;
      r_119__13_ <= r_n_119__13_;
      r_119__12_ <= r_n_119__12_;
      r_119__11_ <= r_n_119__11_;
      r_119__10_ <= r_n_119__10_;
      r_119__9_ <= r_n_119__9_;
      r_119__8_ <= r_n_119__8_;
      r_119__7_ <= r_n_119__7_;
      r_119__6_ <= r_n_119__6_;
      r_119__5_ <= r_n_119__5_;
      r_119__4_ <= r_n_119__4_;
      r_119__3_ <= r_n_119__3_;
      r_119__2_ <= r_n_119__2_;
      r_119__1_ <= r_n_119__1_;
      r_119__0_ <= r_n_119__0_;
    end 
    if(N1912) begin
      r_120__31_ <= r_n_120__31_;
      r_120__30_ <= r_n_120__30_;
      r_120__29_ <= r_n_120__29_;
      r_120__28_ <= r_n_120__28_;
      r_120__27_ <= r_n_120__27_;
      r_120__26_ <= r_n_120__26_;
      r_120__25_ <= r_n_120__25_;
      r_120__24_ <= r_n_120__24_;
      r_120__23_ <= r_n_120__23_;
      r_120__22_ <= r_n_120__22_;
      r_120__21_ <= r_n_120__21_;
      r_120__20_ <= r_n_120__20_;
      r_120__19_ <= r_n_120__19_;
      r_120__18_ <= r_n_120__18_;
      r_120__17_ <= r_n_120__17_;
      r_120__16_ <= r_n_120__16_;
      r_120__15_ <= r_n_120__15_;
      r_120__14_ <= r_n_120__14_;
      r_120__13_ <= r_n_120__13_;
      r_120__12_ <= r_n_120__12_;
      r_120__11_ <= r_n_120__11_;
      r_120__10_ <= r_n_120__10_;
      r_120__9_ <= r_n_120__9_;
      r_120__8_ <= r_n_120__8_;
      r_120__7_ <= r_n_120__7_;
      r_120__6_ <= r_n_120__6_;
      r_120__5_ <= r_n_120__5_;
      r_120__4_ <= r_n_120__4_;
      r_120__3_ <= r_n_120__3_;
      r_120__2_ <= r_n_120__2_;
      r_120__1_ <= r_n_120__1_;
      r_120__0_ <= r_n_120__0_;
    end 
    if(N1913) begin
      r_121__31_ <= r_n_121__31_;
      r_121__30_ <= r_n_121__30_;
      r_121__29_ <= r_n_121__29_;
      r_121__28_ <= r_n_121__28_;
      r_121__27_ <= r_n_121__27_;
      r_121__26_ <= r_n_121__26_;
      r_121__25_ <= r_n_121__25_;
      r_121__24_ <= r_n_121__24_;
      r_121__23_ <= r_n_121__23_;
      r_121__22_ <= r_n_121__22_;
      r_121__21_ <= r_n_121__21_;
      r_121__20_ <= r_n_121__20_;
      r_121__19_ <= r_n_121__19_;
      r_121__18_ <= r_n_121__18_;
      r_121__17_ <= r_n_121__17_;
      r_121__16_ <= r_n_121__16_;
      r_121__15_ <= r_n_121__15_;
      r_121__14_ <= r_n_121__14_;
      r_121__13_ <= r_n_121__13_;
      r_121__12_ <= r_n_121__12_;
      r_121__11_ <= r_n_121__11_;
      r_121__10_ <= r_n_121__10_;
      r_121__9_ <= r_n_121__9_;
      r_121__8_ <= r_n_121__8_;
      r_121__7_ <= r_n_121__7_;
      r_121__6_ <= r_n_121__6_;
      r_121__5_ <= r_n_121__5_;
      r_121__4_ <= r_n_121__4_;
      r_121__3_ <= r_n_121__3_;
      r_121__2_ <= r_n_121__2_;
      r_121__1_ <= r_n_121__1_;
      r_121__0_ <= r_n_121__0_;
    end 
    if(N1914) begin
      r_122__31_ <= r_n_122__31_;
      r_122__30_ <= r_n_122__30_;
      r_122__29_ <= r_n_122__29_;
      r_122__28_ <= r_n_122__28_;
      r_122__27_ <= r_n_122__27_;
      r_122__26_ <= r_n_122__26_;
      r_122__25_ <= r_n_122__25_;
      r_122__24_ <= r_n_122__24_;
      r_122__23_ <= r_n_122__23_;
      r_122__22_ <= r_n_122__22_;
      r_122__21_ <= r_n_122__21_;
      r_122__20_ <= r_n_122__20_;
      r_122__19_ <= r_n_122__19_;
      r_122__18_ <= r_n_122__18_;
      r_122__17_ <= r_n_122__17_;
      r_122__16_ <= r_n_122__16_;
      r_122__15_ <= r_n_122__15_;
      r_122__14_ <= r_n_122__14_;
      r_122__13_ <= r_n_122__13_;
      r_122__12_ <= r_n_122__12_;
      r_122__11_ <= r_n_122__11_;
      r_122__10_ <= r_n_122__10_;
      r_122__9_ <= r_n_122__9_;
      r_122__8_ <= r_n_122__8_;
      r_122__7_ <= r_n_122__7_;
      r_122__6_ <= r_n_122__6_;
      r_122__5_ <= r_n_122__5_;
      r_122__4_ <= r_n_122__4_;
      r_122__3_ <= r_n_122__3_;
      r_122__2_ <= r_n_122__2_;
      r_122__1_ <= r_n_122__1_;
      r_122__0_ <= r_n_122__0_;
    end 
    if(N1915) begin
      r_123__31_ <= r_n_123__31_;
      r_123__30_ <= r_n_123__30_;
      r_123__29_ <= r_n_123__29_;
      r_123__28_ <= r_n_123__28_;
      r_123__27_ <= r_n_123__27_;
      r_123__26_ <= r_n_123__26_;
      r_123__25_ <= r_n_123__25_;
      r_123__24_ <= r_n_123__24_;
      r_123__23_ <= r_n_123__23_;
      r_123__22_ <= r_n_123__22_;
      r_123__21_ <= r_n_123__21_;
      r_123__20_ <= r_n_123__20_;
      r_123__19_ <= r_n_123__19_;
      r_123__18_ <= r_n_123__18_;
      r_123__17_ <= r_n_123__17_;
      r_123__16_ <= r_n_123__16_;
      r_123__15_ <= r_n_123__15_;
      r_123__14_ <= r_n_123__14_;
      r_123__13_ <= r_n_123__13_;
      r_123__12_ <= r_n_123__12_;
      r_123__11_ <= r_n_123__11_;
      r_123__10_ <= r_n_123__10_;
      r_123__9_ <= r_n_123__9_;
      r_123__8_ <= r_n_123__8_;
      r_123__7_ <= r_n_123__7_;
      r_123__6_ <= r_n_123__6_;
      r_123__5_ <= r_n_123__5_;
      r_123__4_ <= r_n_123__4_;
      r_123__3_ <= r_n_123__3_;
      r_123__2_ <= r_n_123__2_;
      r_123__1_ <= r_n_123__1_;
      r_123__0_ <= r_n_123__0_;
    end 
    if(N1916) begin
      r_124__31_ <= r_n_124__31_;
      r_124__30_ <= r_n_124__30_;
      r_124__29_ <= r_n_124__29_;
      r_124__28_ <= r_n_124__28_;
      r_124__27_ <= r_n_124__27_;
      r_124__26_ <= r_n_124__26_;
      r_124__25_ <= r_n_124__25_;
      r_124__24_ <= r_n_124__24_;
      r_124__23_ <= r_n_124__23_;
      r_124__22_ <= r_n_124__22_;
      r_124__21_ <= r_n_124__21_;
      r_124__20_ <= r_n_124__20_;
      r_124__19_ <= r_n_124__19_;
      r_124__18_ <= r_n_124__18_;
      r_124__17_ <= r_n_124__17_;
      r_124__16_ <= r_n_124__16_;
      r_124__15_ <= r_n_124__15_;
      r_124__14_ <= r_n_124__14_;
      r_124__13_ <= r_n_124__13_;
      r_124__12_ <= r_n_124__12_;
      r_124__11_ <= r_n_124__11_;
      r_124__10_ <= r_n_124__10_;
      r_124__9_ <= r_n_124__9_;
      r_124__8_ <= r_n_124__8_;
      r_124__7_ <= r_n_124__7_;
      r_124__6_ <= r_n_124__6_;
      r_124__5_ <= r_n_124__5_;
      r_124__4_ <= r_n_124__4_;
      r_124__3_ <= r_n_124__3_;
      r_124__2_ <= r_n_124__2_;
      r_124__1_ <= r_n_124__1_;
      r_124__0_ <= r_n_124__0_;
    end 
    if(N1917) begin
      r_125__31_ <= r_n_125__31_;
      r_125__30_ <= r_n_125__30_;
      r_125__29_ <= r_n_125__29_;
      r_125__28_ <= r_n_125__28_;
      r_125__27_ <= r_n_125__27_;
      r_125__26_ <= r_n_125__26_;
      r_125__25_ <= r_n_125__25_;
      r_125__24_ <= r_n_125__24_;
      r_125__23_ <= r_n_125__23_;
      r_125__22_ <= r_n_125__22_;
      r_125__21_ <= r_n_125__21_;
      r_125__20_ <= r_n_125__20_;
      r_125__19_ <= r_n_125__19_;
      r_125__18_ <= r_n_125__18_;
      r_125__17_ <= r_n_125__17_;
      r_125__16_ <= r_n_125__16_;
      r_125__15_ <= r_n_125__15_;
      r_125__14_ <= r_n_125__14_;
      r_125__13_ <= r_n_125__13_;
      r_125__12_ <= r_n_125__12_;
      r_125__11_ <= r_n_125__11_;
      r_125__10_ <= r_n_125__10_;
      r_125__9_ <= r_n_125__9_;
      r_125__8_ <= r_n_125__8_;
      r_125__7_ <= r_n_125__7_;
      r_125__6_ <= r_n_125__6_;
      r_125__5_ <= r_n_125__5_;
      r_125__4_ <= r_n_125__4_;
      r_125__3_ <= r_n_125__3_;
      r_125__2_ <= r_n_125__2_;
      r_125__1_ <= r_n_125__1_;
      r_125__0_ <= r_n_125__0_;
    end 
    if(N1918) begin
      r_126__31_ <= r_n_126__31_;
      r_126__30_ <= r_n_126__30_;
      r_126__29_ <= r_n_126__29_;
      r_126__28_ <= r_n_126__28_;
      r_126__27_ <= r_n_126__27_;
      r_126__26_ <= r_n_126__26_;
      r_126__25_ <= r_n_126__25_;
      r_126__24_ <= r_n_126__24_;
      r_126__23_ <= r_n_126__23_;
      r_126__22_ <= r_n_126__22_;
      r_126__21_ <= r_n_126__21_;
      r_126__20_ <= r_n_126__20_;
      r_126__19_ <= r_n_126__19_;
      r_126__18_ <= r_n_126__18_;
      r_126__17_ <= r_n_126__17_;
      r_126__16_ <= r_n_126__16_;
      r_126__15_ <= r_n_126__15_;
      r_126__14_ <= r_n_126__14_;
      r_126__13_ <= r_n_126__13_;
      r_126__12_ <= r_n_126__12_;
      r_126__11_ <= r_n_126__11_;
      r_126__10_ <= r_n_126__10_;
      r_126__9_ <= r_n_126__9_;
      r_126__8_ <= r_n_126__8_;
      r_126__7_ <= r_n_126__7_;
      r_126__6_ <= r_n_126__6_;
      r_126__5_ <= r_n_126__5_;
      r_126__4_ <= r_n_126__4_;
      r_126__3_ <= r_n_126__3_;
      r_126__2_ <= r_n_126__2_;
      r_126__1_ <= r_n_126__1_;
      r_126__0_ <= r_n_126__0_;
    end 
    if(N1919) begin
      r_127__31_ <= r_n_127__31_;
      r_127__30_ <= r_n_127__30_;
      r_127__29_ <= r_n_127__29_;
      r_127__28_ <= r_n_127__28_;
      r_127__27_ <= r_n_127__27_;
      r_127__26_ <= r_n_127__26_;
      r_127__25_ <= r_n_127__25_;
      r_127__24_ <= r_n_127__24_;
      r_127__23_ <= r_n_127__23_;
      r_127__22_ <= r_n_127__22_;
      r_127__21_ <= r_n_127__21_;
      r_127__20_ <= r_n_127__20_;
      r_127__19_ <= r_n_127__19_;
      r_127__18_ <= r_n_127__18_;
      r_127__17_ <= r_n_127__17_;
      r_127__16_ <= r_n_127__16_;
      r_127__15_ <= r_n_127__15_;
      r_127__14_ <= r_n_127__14_;
      r_127__13_ <= r_n_127__13_;
      r_127__12_ <= r_n_127__12_;
      r_127__11_ <= r_n_127__11_;
      r_127__10_ <= r_n_127__10_;
      r_127__9_ <= r_n_127__9_;
      r_127__8_ <= r_n_127__8_;
      r_127__7_ <= r_n_127__7_;
      r_127__6_ <= r_n_127__6_;
      r_127__5_ <= r_n_127__5_;
      r_127__4_ <= r_n_127__4_;
      r_127__3_ <= r_n_127__3_;
      r_127__2_ <= r_n_127__2_;
      r_127__1_ <= r_n_127__1_;
      r_127__0_ <= r_n_127__0_;
    end 
    if(N1920) begin
      r_128__31_ <= r_n_128__31_;
      r_128__30_ <= r_n_128__30_;
      r_128__29_ <= r_n_128__29_;
      r_128__28_ <= r_n_128__28_;
      r_128__27_ <= r_n_128__27_;
      r_128__26_ <= r_n_128__26_;
      r_128__25_ <= r_n_128__25_;
      r_128__24_ <= r_n_128__24_;
      r_128__23_ <= r_n_128__23_;
      r_128__22_ <= r_n_128__22_;
      r_128__21_ <= r_n_128__21_;
      r_128__20_ <= r_n_128__20_;
      r_128__19_ <= r_n_128__19_;
      r_128__18_ <= r_n_128__18_;
      r_128__17_ <= r_n_128__17_;
      r_128__16_ <= r_n_128__16_;
      r_128__15_ <= r_n_128__15_;
      r_128__14_ <= r_n_128__14_;
      r_128__13_ <= r_n_128__13_;
      r_128__12_ <= r_n_128__12_;
      r_128__11_ <= r_n_128__11_;
      r_128__10_ <= r_n_128__10_;
      r_128__9_ <= r_n_128__9_;
      r_128__8_ <= r_n_128__8_;
      r_128__7_ <= r_n_128__7_;
      r_128__6_ <= r_n_128__6_;
      r_128__5_ <= r_n_128__5_;
      r_128__4_ <= r_n_128__4_;
      r_128__3_ <= r_n_128__3_;
      r_128__2_ <= r_n_128__2_;
      r_128__1_ <= r_n_128__1_;
      r_128__0_ <= r_n_128__0_;
    end 
    if(N1921) begin
      r_129__31_ <= r_n_129__31_;
      r_129__30_ <= r_n_129__30_;
      r_129__29_ <= r_n_129__29_;
      r_129__28_ <= r_n_129__28_;
      r_129__27_ <= r_n_129__27_;
      r_129__26_ <= r_n_129__26_;
      r_129__25_ <= r_n_129__25_;
      r_129__24_ <= r_n_129__24_;
      r_129__23_ <= r_n_129__23_;
      r_129__22_ <= r_n_129__22_;
      r_129__21_ <= r_n_129__21_;
      r_129__20_ <= r_n_129__20_;
      r_129__19_ <= r_n_129__19_;
      r_129__18_ <= r_n_129__18_;
      r_129__17_ <= r_n_129__17_;
      r_129__16_ <= r_n_129__16_;
      r_129__15_ <= r_n_129__15_;
      r_129__14_ <= r_n_129__14_;
      r_129__13_ <= r_n_129__13_;
      r_129__12_ <= r_n_129__12_;
      r_129__11_ <= r_n_129__11_;
      r_129__10_ <= r_n_129__10_;
      r_129__9_ <= r_n_129__9_;
      r_129__8_ <= r_n_129__8_;
      r_129__7_ <= r_n_129__7_;
      r_129__6_ <= r_n_129__6_;
      r_129__5_ <= r_n_129__5_;
      r_129__4_ <= r_n_129__4_;
      r_129__3_ <= r_n_129__3_;
      r_129__2_ <= r_n_129__2_;
      r_129__1_ <= r_n_129__1_;
      r_129__0_ <= r_n_129__0_;
    end 
    if(N1922) begin
      r_130__31_ <= r_n_130__31_;
      r_130__30_ <= r_n_130__30_;
      r_130__29_ <= r_n_130__29_;
      r_130__28_ <= r_n_130__28_;
      r_130__27_ <= r_n_130__27_;
      r_130__26_ <= r_n_130__26_;
      r_130__25_ <= r_n_130__25_;
      r_130__24_ <= r_n_130__24_;
      r_130__23_ <= r_n_130__23_;
      r_130__22_ <= r_n_130__22_;
      r_130__21_ <= r_n_130__21_;
      r_130__20_ <= r_n_130__20_;
      r_130__19_ <= r_n_130__19_;
      r_130__18_ <= r_n_130__18_;
      r_130__17_ <= r_n_130__17_;
      r_130__16_ <= r_n_130__16_;
      r_130__15_ <= r_n_130__15_;
      r_130__14_ <= r_n_130__14_;
      r_130__13_ <= r_n_130__13_;
      r_130__12_ <= r_n_130__12_;
      r_130__11_ <= r_n_130__11_;
      r_130__10_ <= r_n_130__10_;
      r_130__9_ <= r_n_130__9_;
      r_130__8_ <= r_n_130__8_;
      r_130__7_ <= r_n_130__7_;
      r_130__6_ <= r_n_130__6_;
      r_130__5_ <= r_n_130__5_;
      r_130__4_ <= r_n_130__4_;
      r_130__3_ <= r_n_130__3_;
      r_130__2_ <= r_n_130__2_;
      r_130__1_ <= r_n_130__1_;
      r_130__0_ <= r_n_130__0_;
    end 
    if(N1923) begin
      r_131__31_ <= r_n_131__31_;
      r_131__30_ <= r_n_131__30_;
      r_131__29_ <= r_n_131__29_;
      r_131__28_ <= r_n_131__28_;
      r_131__27_ <= r_n_131__27_;
      r_131__26_ <= r_n_131__26_;
      r_131__25_ <= r_n_131__25_;
      r_131__24_ <= r_n_131__24_;
      r_131__23_ <= r_n_131__23_;
      r_131__22_ <= r_n_131__22_;
      r_131__21_ <= r_n_131__21_;
      r_131__20_ <= r_n_131__20_;
      r_131__19_ <= r_n_131__19_;
      r_131__18_ <= r_n_131__18_;
      r_131__17_ <= r_n_131__17_;
      r_131__16_ <= r_n_131__16_;
      r_131__15_ <= r_n_131__15_;
      r_131__14_ <= r_n_131__14_;
      r_131__13_ <= r_n_131__13_;
      r_131__12_ <= r_n_131__12_;
      r_131__11_ <= r_n_131__11_;
      r_131__10_ <= r_n_131__10_;
      r_131__9_ <= r_n_131__9_;
      r_131__8_ <= r_n_131__8_;
      r_131__7_ <= r_n_131__7_;
      r_131__6_ <= r_n_131__6_;
      r_131__5_ <= r_n_131__5_;
      r_131__4_ <= r_n_131__4_;
      r_131__3_ <= r_n_131__3_;
      r_131__2_ <= r_n_131__2_;
      r_131__1_ <= r_n_131__1_;
      r_131__0_ <= r_n_131__0_;
    end 
    if(N1924) begin
      r_132__31_ <= r_n_132__31_;
      r_132__30_ <= r_n_132__30_;
      r_132__29_ <= r_n_132__29_;
      r_132__28_ <= r_n_132__28_;
      r_132__27_ <= r_n_132__27_;
      r_132__26_ <= r_n_132__26_;
      r_132__25_ <= r_n_132__25_;
      r_132__24_ <= r_n_132__24_;
      r_132__23_ <= r_n_132__23_;
      r_132__22_ <= r_n_132__22_;
      r_132__21_ <= r_n_132__21_;
      r_132__20_ <= r_n_132__20_;
      r_132__19_ <= r_n_132__19_;
      r_132__18_ <= r_n_132__18_;
      r_132__17_ <= r_n_132__17_;
      r_132__16_ <= r_n_132__16_;
      r_132__15_ <= r_n_132__15_;
      r_132__14_ <= r_n_132__14_;
      r_132__13_ <= r_n_132__13_;
      r_132__12_ <= r_n_132__12_;
      r_132__11_ <= r_n_132__11_;
      r_132__10_ <= r_n_132__10_;
      r_132__9_ <= r_n_132__9_;
      r_132__8_ <= r_n_132__8_;
      r_132__7_ <= r_n_132__7_;
      r_132__6_ <= r_n_132__6_;
      r_132__5_ <= r_n_132__5_;
      r_132__4_ <= r_n_132__4_;
      r_132__3_ <= r_n_132__3_;
      r_132__2_ <= r_n_132__2_;
      r_132__1_ <= r_n_132__1_;
      r_132__0_ <= r_n_132__0_;
    end 
    if(N1925) begin
      r_133__31_ <= r_n_133__31_;
      r_133__30_ <= r_n_133__30_;
      r_133__29_ <= r_n_133__29_;
      r_133__28_ <= r_n_133__28_;
      r_133__27_ <= r_n_133__27_;
      r_133__26_ <= r_n_133__26_;
      r_133__25_ <= r_n_133__25_;
      r_133__24_ <= r_n_133__24_;
      r_133__23_ <= r_n_133__23_;
      r_133__22_ <= r_n_133__22_;
      r_133__21_ <= r_n_133__21_;
      r_133__20_ <= r_n_133__20_;
      r_133__19_ <= r_n_133__19_;
      r_133__18_ <= r_n_133__18_;
      r_133__17_ <= r_n_133__17_;
      r_133__16_ <= r_n_133__16_;
      r_133__15_ <= r_n_133__15_;
      r_133__14_ <= r_n_133__14_;
      r_133__13_ <= r_n_133__13_;
      r_133__12_ <= r_n_133__12_;
      r_133__11_ <= r_n_133__11_;
      r_133__10_ <= r_n_133__10_;
      r_133__9_ <= r_n_133__9_;
      r_133__8_ <= r_n_133__8_;
      r_133__7_ <= r_n_133__7_;
      r_133__6_ <= r_n_133__6_;
      r_133__5_ <= r_n_133__5_;
      r_133__4_ <= r_n_133__4_;
      r_133__3_ <= r_n_133__3_;
      r_133__2_ <= r_n_133__2_;
      r_133__1_ <= r_n_133__1_;
      r_133__0_ <= r_n_133__0_;
    end 
    if(N1926) begin
      r_134__31_ <= r_n_134__31_;
      r_134__30_ <= r_n_134__30_;
      r_134__29_ <= r_n_134__29_;
      r_134__28_ <= r_n_134__28_;
      r_134__27_ <= r_n_134__27_;
      r_134__26_ <= r_n_134__26_;
      r_134__25_ <= r_n_134__25_;
      r_134__24_ <= r_n_134__24_;
      r_134__23_ <= r_n_134__23_;
      r_134__22_ <= r_n_134__22_;
      r_134__21_ <= r_n_134__21_;
      r_134__20_ <= r_n_134__20_;
      r_134__19_ <= r_n_134__19_;
      r_134__18_ <= r_n_134__18_;
      r_134__17_ <= r_n_134__17_;
      r_134__16_ <= r_n_134__16_;
      r_134__15_ <= r_n_134__15_;
      r_134__14_ <= r_n_134__14_;
      r_134__13_ <= r_n_134__13_;
      r_134__12_ <= r_n_134__12_;
      r_134__11_ <= r_n_134__11_;
      r_134__10_ <= r_n_134__10_;
      r_134__9_ <= r_n_134__9_;
      r_134__8_ <= r_n_134__8_;
      r_134__7_ <= r_n_134__7_;
      r_134__6_ <= r_n_134__6_;
      r_134__5_ <= r_n_134__5_;
      r_134__4_ <= r_n_134__4_;
      r_134__3_ <= r_n_134__3_;
      r_134__2_ <= r_n_134__2_;
      r_134__1_ <= r_n_134__1_;
      r_134__0_ <= r_n_134__0_;
    end 
    if(N1927) begin
      r_135__31_ <= r_n_135__31_;
      r_135__30_ <= r_n_135__30_;
      r_135__29_ <= r_n_135__29_;
      r_135__28_ <= r_n_135__28_;
      r_135__27_ <= r_n_135__27_;
      r_135__26_ <= r_n_135__26_;
      r_135__25_ <= r_n_135__25_;
      r_135__24_ <= r_n_135__24_;
      r_135__23_ <= r_n_135__23_;
      r_135__22_ <= r_n_135__22_;
      r_135__21_ <= r_n_135__21_;
      r_135__20_ <= r_n_135__20_;
      r_135__19_ <= r_n_135__19_;
      r_135__18_ <= r_n_135__18_;
      r_135__17_ <= r_n_135__17_;
      r_135__16_ <= r_n_135__16_;
      r_135__15_ <= r_n_135__15_;
      r_135__14_ <= r_n_135__14_;
      r_135__13_ <= r_n_135__13_;
      r_135__12_ <= r_n_135__12_;
      r_135__11_ <= r_n_135__11_;
      r_135__10_ <= r_n_135__10_;
      r_135__9_ <= r_n_135__9_;
      r_135__8_ <= r_n_135__8_;
      r_135__7_ <= r_n_135__7_;
      r_135__6_ <= r_n_135__6_;
      r_135__5_ <= r_n_135__5_;
      r_135__4_ <= r_n_135__4_;
      r_135__3_ <= r_n_135__3_;
      r_135__2_ <= r_n_135__2_;
      r_135__1_ <= r_n_135__1_;
      r_135__0_ <= r_n_135__0_;
    end 
    if(N1928) begin
      r_136__31_ <= r_n_136__31_;
      r_136__30_ <= r_n_136__30_;
      r_136__29_ <= r_n_136__29_;
      r_136__28_ <= r_n_136__28_;
      r_136__27_ <= r_n_136__27_;
      r_136__26_ <= r_n_136__26_;
      r_136__25_ <= r_n_136__25_;
      r_136__24_ <= r_n_136__24_;
      r_136__23_ <= r_n_136__23_;
      r_136__22_ <= r_n_136__22_;
      r_136__21_ <= r_n_136__21_;
      r_136__20_ <= r_n_136__20_;
      r_136__19_ <= r_n_136__19_;
      r_136__18_ <= r_n_136__18_;
      r_136__17_ <= r_n_136__17_;
      r_136__16_ <= r_n_136__16_;
      r_136__15_ <= r_n_136__15_;
      r_136__14_ <= r_n_136__14_;
      r_136__13_ <= r_n_136__13_;
      r_136__12_ <= r_n_136__12_;
      r_136__11_ <= r_n_136__11_;
      r_136__10_ <= r_n_136__10_;
      r_136__9_ <= r_n_136__9_;
      r_136__8_ <= r_n_136__8_;
      r_136__7_ <= r_n_136__7_;
      r_136__6_ <= r_n_136__6_;
      r_136__5_ <= r_n_136__5_;
      r_136__4_ <= r_n_136__4_;
      r_136__3_ <= r_n_136__3_;
      r_136__2_ <= r_n_136__2_;
      r_136__1_ <= r_n_136__1_;
      r_136__0_ <= r_n_136__0_;
    end 
    if(N1929) begin
      r_137__31_ <= r_n_137__31_;
      r_137__30_ <= r_n_137__30_;
      r_137__29_ <= r_n_137__29_;
      r_137__28_ <= r_n_137__28_;
      r_137__27_ <= r_n_137__27_;
      r_137__26_ <= r_n_137__26_;
      r_137__25_ <= r_n_137__25_;
      r_137__24_ <= r_n_137__24_;
      r_137__23_ <= r_n_137__23_;
      r_137__22_ <= r_n_137__22_;
      r_137__21_ <= r_n_137__21_;
      r_137__20_ <= r_n_137__20_;
      r_137__19_ <= r_n_137__19_;
      r_137__18_ <= r_n_137__18_;
      r_137__17_ <= r_n_137__17_;
      r_137__16_ <= r_n_137__16_;
      r_137__15_ <= r_n_137__15_;
      r_137__14_ <= r_n_137__14_;
      r_137__13_ <= r_n_137__13_;
      r_137__12_ <= r_n_137__12_;
      r_137__11_ <= r_n_137__11_;
      r_137__10_ <= r_n_137__10_;
      r_137__9_ <= r_n_137__9_;
      r_137__8_ <= r_n_137__8_;
      r_137__7_ <= r_n_137__7_;
      r_137__6_ <= r_n_137__6_;
      r_137__5_ <= r_n_137__5_;
      r_137__4_ <= r_n_137__4_;
      r_137__3_ <= r_n_137__3_;
      r_137__2_ <= r_n_137__2_;
      r_137__1_ <= r_n_137__1_;
      r_137__0_ <= r_n_137__0_;
    end 
    if(N1930) begin
      r_138__31_ <= r_n_138__31_;
      r_138__30_ <= r_n_138__30_;
      r_138__29_ <= r_n_138__29_;
      r_138__28_ <= r_n_138__28_;
      r_138__27_ <= r_n_138__27_;
      r_138__26_ <= r_n_138__26_;
      r_138__25_ <= r_n_138__25_;
      r_138__24_ <= r_n_138__24_;
      r_138__23_ <= r_n_138__23_;
      r_138__22_ <= r_n_138__22_;
      r_138__21_ <= r_n_138__21_;
      r_138__20_ <= r_n_138__20_;
      r_138__19_ <= r_n_138__19_;
      r_138__18_ <= r_n_138__18_;
      r_138__17_ <= r_n_138__17_;
      r_138__16_ <= r_n_138__16_;
      r_138__15_ <= r_n_138__15_;
      r_138__14_ <= r_n_138__14_;
      r_138__13_ <= r_n_138__13_;
      r_138__12_ <= r_n_138__12_;
      r_138__11_ <= r_n_138__11_;
      r_138__10_ <= r_n_138__10_;
      r_138__9_ <= r_n_138__9_;
      r_138__8_ <= r_n_138__8_;
      r_138__7_ <= r_n_138__7_;
      r_138__6_ <= r_n_138__6_;
      r_138__5_ <= r_n_138__5_;
      r_138__4_ <= r_n_138__4_;
      r_138__3_ <= r_n_138__3_;
      r_138__2_ <= r_n_138__2_;
      r_138__1_ <= r_n_138__1_;
      r_138__0_ <= r_n_138__0_;
    end 
    if(N1931) begin
      r_139__31_ <= r_n_139__31_;
      r_139__30_ <= r_n_139__30_;
      r_139__29_ <= r_n_139__29_;
      r_139__28_ <= r_n_139__28_;
      r_139__27_ <= r_n_139__27_;
      r_139__26_ <= r_n_139__26_;
      r_139__25_ <= r_n_139__25_;
      r_139__24_ <= r_n_139__24_;
      r_139__23_ <= r_n_139__23_;
      r_139__22_ <= r_n_139__22_;
      r_139__21_ <= r_n_139__21_;
      r_139__20_ <= r_n_139__20_;
      r_139__19_ <= r_n_139__19_;
      r_139__18_ <= r_n_139__18_;
      r_139__17_ <= r_n_139__17_;
      r_139__16_ <= r_n_139__16_;
      r_139__15_ <= r_n_139__15_;
      r_139__14_ <= r_n_139__14_;
      r_139__13_ <= r_n_139__13_;
      r_139__12_ <= r_n_139__12_;
      r_139__11_ <= r_n_139__11_;
      r_139__10_ <= r_n_139__10_;
      r_139__9_ <= r_n_139__9_;
      r_139__8_ <= r_n_139__8_;
      r_139__7_ <= r_n_139__7_;
      r_139__6_ <= r_n_139__6_;
      r_139__5_ <= r_n_139__5_;
      r_139__4_ <= r_n_139__4_;
      r_139__3_ <= r_n_139__3_;
      r_139__2_ <= r_n_139__2_;
      r_139__1_ <= r_n_139__1_;
      r_139__0_ <= r_n_139__0_;
    end 
    if(N1932) begin
      r_140__31_ <= r_n_140__31_;
      r_140__30_ <= r_n_140__30_;
      r_140__29_ <= r_n_140__29_;
      r_140__28_ <= r_n_140__28_;
      r_140__27_ <= r_n_140__27_;
      r_140__26_ <= r_n_140__26_;
      r_140__25_ <= r_n_140__25_;
      r_140__24_ <= r_n_140__24_;
      r_140__23_ <= r_n_140__23_;
      r_140__22_ <= r_n_140__22_;
      r_140__21_ <= r_n_140__21_;
      r_140__20_ <= r_n_140__20_;
      r_140__19_ <= r_n_140__19_;
      r_140__18_ <= r_n_140__18_;
      r_140__17_ <= r_n_140__17_;
      r_140__16_ <= r_n_140__16_;
      r_140__15_ <= r_n_140__15_;
      r_140__14_ <= r_n_140__14_;
      r_140__13_ <= r_n_140__13_;
      r_140__12_ <= r_n_140__12_;
      r_140__11_ <= r_n_140__11_;
      r_140__10_ <= r_n_140__10_;
      r_140__9_ <= r_n_140__9_;
      r_140__8_ <= r_n_140__8_;
      r_140__7_ <= r_n_140__7_;
      r_140__6_ <= r_n_140__6_;
      r_140__5_ <= r_n_140__5_;
      r_140__4_ <= r_n_140__4_;
      r_140__3_ <= r_n_140__3_;
      r_140__2_ <= r_n_140__2_;
      r_140__1_ <= r_n_140__1_;
      r_140__0_ <= r_n_140__0_;
    end 
    if(N1933) begin
      r_141__31_ <= r_n_141__31_;
      r_141__30_ <= r_n_141__30_;
      r_141__29_ <= r_n_141__29_;
      r_141__28_ <= r_n_141__28_;
      r_141__27_ <= r_n_141__27_;
      r_141__26_ <= r_n_141__26_;
      r_141__25_ <= r_n_141__25_;
      r_141__24_ <= r_n_141__24_;
      r_141__23_ <= r_n_141__23_;
      r_141__22_ <= r_n_141__22_;
      r_141__21_ <= r_n_141__21_;
      r_141__20_ <= r_n_141__20_;
      r_141__19_ <= r_n_141__19_;
      r_141__18_ <= r_n_141__18_;
      r_141__17_ <= r_n_141__17_;
      r_141__16_ <= r_n_141__16_;
      r_141__15_ <= r_n_141__15_;
      r_141__14_ <= r_n_141__14_;
      r_141__13_ <= r_n_141__13_;
      r_141__12_ <= r_n_141__12_;
      r_141__11_ <= r_n_141__11_;
      r_141__10_ <= r_n_141__10_;
      r_141__9_ <= r_n_141__9_;
      r_141__8_ <= r_n_141__8_;
      r_141__7_ <= r_n_141__7_;
      r_141__6_ <= r_n_141__6_;
      r_141__5_ <= r_n_141__5_;
      r_141__4_ <= r_n_141__4_;
      r_141__3_ <= r_n_141__3_;
      r_141__2_ <= r_n_141__2_;
      r_141__1_ <= r_n_141__1_;
      r_141__0_ <= r_n_141__0_;
    end 
    if(N1934) begin
      r_142__31_ <= r_n_142__31_;
      r_142__30_ <= r_n_142__30_;
      r_142__29_ <= r_n_142__29_;
      r_142__28_ <= r_n_142__28_;
      r_142__27_ <= r_n_142__27_;
      r_142__26_ <= r_n_142__26_;
      r_142__25_ <= r_n_142__25_;
      r_142__24_ <= r_n_142__24_;
      r_142__23_ <= r_n_142__23_;
      r_142__22_ <= r_n_142__22_;
      r_142__21_ <= r_n_142__21_;
      r_142__20_ <= r_n_142__20_;
      r_142__19_ <= r_n_142__19_;
      r_142__18_ <= r_n_142__18_;
      r_142__17_ <= r_n_142__17_;
      r_142__16_ <= r_n_142__16_;
      r_142__15_ <= r_n_142__15_;
      r_142__14_ <= r_n_142__14_;
      r_142__13_ <= r_n_142__13_;
      r_142__12_ <= r_n_142__12_;
      r_142__11_ <= r_n_142__11_;
      r_142__10_ <= r_n_142__10_;
      r_142__9_ <= r_n_142__9_;
      r_142__8_ <= r_n_142__8_;
      r_142__7_ <= r_n_142__7_;
      r_142__6_ <= r_n_142__6_;
      r_142__5_ <= r_n_142__5_;
      r_142__4_ <= r_n_142__4_;
      r_142__3_ <= r_n_142__3_;
      r_142__2_ <= r_n_142__2_;
      r_142__1_ <= r_n_142__1_;
      r_142__0_ <= r_n_142__0_;
    end 
    if(N1935) begin
      r_143__31_ <= r_n_143__31_;
      r_143__30_ <= r_n_143__30_;
      r_143__29_ <= r_n_143__29_;
      r_143__28_ <= r_n_143__28_;
      r_143__27_ <= r_n_143__27_;
      r_143__26_ <= r_n_143__26_;
      r_143__25_ <= r_n_143__25_;
      r_143__24_ <= r_n_143__24_;
      r_143__23_ <= r_n_143__23_;
      r_143__22_ <= r_n_143__22_;
      r_143__21_ <= r_n_143__21_;
      r_143__20_ <= r_n_143__20_;
      r_143__19_ <= r_n_143__19_;
      r_143__18_ <= r_n_143__18_;
      r_143__17_ <= r_n_143__17_;
      r_143__16_ <= r_n_143__16_;
      r_143__15_ <= r_n_143__15_;
      r_143__14_ <= r_n_143__14_;
      r_143__13_ <= r_n_143__13_;
      r_143__12_ <= r_n_143__12_;
      r_143__11_ <= r_n_143__11_;
      r_143__10_ <= r_n_143__10_;
      r_143__9_ <= r_n_143__9_;
      r_143__8_ <= r_n_143__8_;
      r_143__7_ <= r_n_143__7_;
      r_143__6_ <= r_n_143__6_;
      r_143__5_ <= r_n_143__5_;
      r_143__4_ <= r_n_143__4_;
      r_143__3_ <= r_n_143__3_;
      r_143__2_ <= r_n_143__2_;
      r_143__1_ <= r_n_143__1_;
      r_143__0_ <= r_n_143__0_;
    end 
    if(N1936) begin
      r_144__31_ <= r_n_144__31_;
      r_144__30_ <= r_n_144__30_;
      r_144__29_ <= r_n_144__29_;
      r_144__28_ <= r_n_144__28_;
      r_144__27_ <= r_n_144__27_;
      r_144__26_ <= r_n_144__26_;
      r_144__25_ <= r_n_144__25_;
      r_144__24_ <= r_n_144__24_;
      r_144__23_ <= r_n_144__23_;
      r_144__22_ <= r_n_144__22_;
      r_144__21_ <= r_n_144__21_;
      r_144__20_ <= r_n_144__20_;
      r_144__19_ <= r_n_144__19_;
      r_144__18_ <= r_n_144__18_;
      r_144__17_ <= r_n_144__17_;
      r_144__16_ <= r_n_144__16_;
      r_144__15_ <= r_n_144__15_;
      r_144__14_ <= r_n_144__14_;
      r_144__13_ <= r_n_144__13_;
      r_144__12_ <= r_n_144__12_;
      r_144__11_ <= r_n_144__11_;
      r_144__10_ <= r_n_144__10_;
      r_144__9_ <= r_n_144__9_;
      r_144__8_ <= r_n_144__8_;
      r_144__7_ <= r_n_144__7_;
      r_144__6_ <= r_n_144__6_;
      r_144__5_ <= r_n_144__5_;
      r_144__4_ <= r_n_144__4_;
      r_144__3_ <= r_n_144__3_;
      r_144__2_ <= r_n_144__2_;
      r_144__1_ <= r_n_144__1_;
      r_144__0_ <= r_n_144__0_;
    end 
    if(N1937) begin
      r_145__31_ <= r_n_145__31_;
      r_145__30_ <= r_n_145__30_;
      r_145__29_ <= r_n_145__29_;
      r_145__28_ <= r_n_145__28_;
      r_145__27_ <= r_n_145__27_;
      r_145__26_ <= r_n_145__26_;
      r_145__25_ <= r_n_145__25_;
      r_145__24_ <= r_n_145__24_;
      r_145__23_ <= r_n_145__23_;
      r_145__22_ <= r_n_145__22_;
      r_145__21_ <= r_n_145__21_;
      r_145__20_ <= r_n_145__20_;
      r_145__19_ <= r_n_145__19_;
      r_145__18_ <= r_n_145__18_;
      r_145__17_ <= r_n_145__17_;
      r_145__16_ <= r_n_145__16_;
      r_145__15_ <= r_n_145__15_;
      r_145__14_ <= r_n_145__14_;
      r_145__13_ <= r_n_145__13_;
      r_145__12_ <= r_n_145__12_;
      r_145__11_ <= r_n_145__11_;
      r_145__10_ <= r_n_145__10_;
      r_145__9_ <= r_n_145__9_;
      r_145__8_ <= r_n_145__8_;
      r_145__7_ <= r_n_145__7_;
      r_145__6_ <= r_n_145__6_;
      r_145__5_ <= r_n_145__5_;
      r_145__4_ <= r_n_145__4_;
      r_145__3_ <= r_n_145__3_;
      r_145__2_ <= r_n_145__2_;
      r_145__1_ <= r_n_145__1_;
      r_145__0_ <= r_n_145__0_;
    end 
    if(N1938) begin
      r_146__31_ <= r_n_146__31_;
      r_146__30_ <= r_n_146__30_;
      r_146__29_ <= r_n_146__29_;
      r_146__28_ <= r_n_146__28_;
      r_146__27_ <= r_n_146__27_;
      r_146__26_ <= r_n_146__26_;
      r_146__25_ <= r_n_146__25_;
      r_146__24_ <= r_n_146__24_;
      r_146__23_ <= r_n_146__23_;
      r_146__22_ <= r_n_146__22_;
      r_146__21_ <= r_n_146__21_;
      r_146__20_ <= r_n_146__20_;
      r_146__19_ <= r_n_146__19_;
      r_146__18_ <= r_n_146__18_;
      r_146__17_ <= r_n_146__17_;
      r_146__16_ <= r_n_146__16_;
      r_146__15_ <= r_n_146__15_;
      r_146__14_ <= r_n_146__14_;
      r_146__13_ <= r_n_146__13_;
      r_146__12_ <= r_n_146__12_;
      r_146__11_ <= r_n_146__11_;
      r_146__10_ <= r_n_146__10_;
      r_146__9_ <= r_n_146__9_;
      r_146__8_ <= r_n_146__8_;
      r_146__7_ <= r_n_146__7_;
      r_146__6_ <= r_n_146__6_;
      r_146__5_ <= r_n_146__5_;
      r_146__4_ <= r_n_146__4_;
      r_146__3_ <= r_n_146__3_;
      r_146__2_ <= r_n_146__2_;
      r_146__1_ <= r_n_146__1_;
      r_146__0_ <= r_n_146__0_;
    end 
    if(N1939) begin
      r_147__31_ <= r_n_147__31_;
      r_147__30_ <= r_n_147__30_;
      r_147__29_ <= r_n_147__29_;
      r_147__28_ <= r_n_147__28_;
      r_147__27_ <= r_n_147__27_;
      r_147__26_ <= r_n_147__26_;
      r_147__25_ <= r_n_147__25_;
      r_147__24_ <= r_n_147__24_;
      r_147__23_ <= r_n_147__23_;
      r_147__22_ <= r_n_147__22_;
      r_147__21_ <= r_n_147__21_;
      r_147__20_ <= r_n_147__20_;
      r_147__19_ <= r_n_147__19_;
      r_147__18_ <= r_n_147__18_;
      r_147__17_ <= r_n_147__17_;
      r_147__16_ <= r_n_147__16_;
      r_147__15_ <= r_n_147__15_;
      r_147__14_ <= r_n_147__14_;
      r_147__13_ <= r_n_147__13_;
      r_147__12_ <= r_n_147__12_;
      r_147__11_ <= r_n_147__11_;
      r_147__10_ <= r_n_147__10_;
      r_147__9_ <= r_n_147__9_;
      r_147__8_ <= r_n_147__8_;
      r_147__7_ <= r_n_147__7_;
      r_147__6_ <= r_n_147__6_;
      r_147__5_ <= r_n_147__5_;
      r_147__4_ <= r_n_147__4_;
      r_147__3_ <= r_n_147__3_;
      r_147__2_ <= r_n_147__2_;
      r_147__1_ <= r_n_147__1_;
      r_147__0_ <= r_n_147__0_;
    end 
    if(N1940) begin
      r_148__31_ <= r_n_148__31_;
      r_148__30_ <= r_n_148__30_;
      r_148__29_ <= r_n_148__29_;
      r_148__28_ <= r_n_148__28_;
      r_148__27_ <= r_n_148__27_;
      r_148__26_ <= r_n_148__26_;
      r_148__25_ <= r_n_148__25_;
      r_148__24_ <= r_n_148__24_;
      r_148__23_ <= r_n_148__23_;
      r_148__22_ <= r_n_148__22_;
      r_148__21_ <= r_n_148__21_;
      r_148__20_ <= r_n_148__20_;
      r_148__19_ <= r_n_148__19_;
      r_148__18_ <= r_n_148__18_;
      r_148__17_ <= r_n_148__17_;
      r_148__16_ <= r_n_148__16_;
      r_148__15_ <= r_n_148__15_;
      r_148__14_ <= r_n_148__14_;
      r_148__13_ <= r_n_148__13_;
      r_148__12_ <= r_n_148__12_;
      r_148__11_ <= r_n_148__11_;
      r_148__10_ <= r_n_148__10_;
      r_148__9_ <= r_n_148__9_;
      r_148__8_ <= r_n_148__8_;
      r_148__7_ <= r_n_148__7_;
      r_148__6_ <= r_n_148__6_;
      r_148__5_ <= r_n_148__5_;
      r_148__4_ <= r_n_148__4_;
      r_148__3_ <= r_n_148__3_;
      r_148__2_ <= r_n_148__2_;
      r_148__1_ <= r_n_148__1_;
      r_148__0_ <= r_n_148__0_;
    end 
    if(N1941) begin
      r_149__31_ <= r_n_149__31_;
      r_149__30_ <= r_n_149__30_;
      r_149__29_ <= r_n_149__29_;
      r_149__28_ <= r_n_149__28_;
      r_149__27_ <= r_n_149__27_;
      r_149__26_ <= r_n_149__26_;
      r_149__25_ <= r_n_149__25_;
      r_149__24_ <= r_n_149__24_;
      r_149__23_ <= r_n_149__23_;
      r_149__22_ <= r_n_149__22_;
      r_149__21_ <= r_n_149__21_;
      r_149__20_ <= r_n_149__20_;
      r_149__19_ <= r_n_149__19_;
      r_149__18_ <= r_n_149__18_;
      r_149__17_ <= r_n_149__17_;
      r_149__16_ <= r_n_149__16_;
      r_149__15_ <= r_n_149__15_;
      r_149__14_ <= r_n_149__14_;
      r_149__13_ <= r_n_149__13_;
      r_149__12_ <= r_n_149__12_;
      r_149__11_ <= r_n_149__11_;
      r_149__10_ <= r_n_149__10_;
      r_149__9_ <= r_n_149__9_;
      r_149__8_ <= r_n_149__8_;
      r_149__7_ <= r_n_149__7_;
      r_149__6_ <= r_n_149__6_;
      r_149__5_ <= r_n_149__5_;
      r_149__4_ <= r_n_149__4_;
      r_149__3_ <= r_n_149__3_;
      r_149__2_ <= r_n_149__2_;
      r_149__1_ <= r_n_149__1_;
      r_149__0_ <= r_n_149__0_;
    end 
    if(N1942) begin
      r_150__31_ <= r_n_150__31_;
      r_150__30_ <= r_n_150__30_;
      r_150__29_ <= r_n_150__29_;
      r_150__28_ <= r_n_150__28_;
      r_150__27_ <= r_n_150__27_;
      r_150__26_ <= r_n_150__26_;
      r_150__25_ <= r_n_150__25_;
      r_150__24_ <= r_n_150__24_;
      r_150__23_ <= r_n_150__23_;
      r_150__22_ <= r_n_150__22_;
      r_150__21_ <= r_n_150__21_;
      r_150__20_ <= r_n_150__20_;
      r_150__19_ <= r_n_150__19_;
      r_150__18_ <= r_n_150__18_;
      r_150__17_ <= r_n_150__17_;
      r_150__16_ <= r_n_150__16_;
      r_150__15_ <= r_n_150__15_;
      r_150__14_ <= r_n_150__14_;
      r_150__13_ <= r_n_150__13_;
      r_150__12_ <= r_n_150__12_;
      r_150__11_ <= r_n_150__11_;
      r_150__10_ <= r_n_150__10_;
      r_150__9_ <= r_n_150__9_;
      r_150__8_ <= r_n_150__8_;
      r_150__7_ <= r_n_150__7_;
      r_150__6_ <= r_n_150__6_;
      r_150__5_ <= r_n_150__5_;
      r_150__4_ <= r_n_150__4_;
      r_150__3_ <= r_n_150__3_;
      r_150__2_ <= r_n_150__2_;
      r_150__1_ <= r_n_150__1_;
      r_150__0_ <= r_n_150__0_;
    end 
    if(N1943) begin
      r_151__31_ <= r_n_151__31_;
      r_151__30_ <= r_n_151__30_;
      r_151__29_ <= r_n_151__29_;
      r_151__28_ <= r_n_151__28_;
      r_151__27_ <= r_n_151__27_;
      r_151__26_ <= r_n_151__26_;
      r_151__25_ <= r_n_151__25_;
      r_151__24_ <= r_n_151__24_;
      r_151__23_ <= r_n_151__23_;
      r_151__22_ <= r_n_151__22_;
      r_151__21_ <= r_n_151__21_;
      r_151__20_ <= r_n_151__20_;
      r_151__19_ <= r_n_151__19_;
      r_151__18_ <= r_n_151__18_;
      r_151__17_ <= r_n_151__17_;
      r_151__16_ <= r_n_151__16_;
      r_151__15_ <= r_n_151__15_;
      r_151__14_ <= r_n_151__14_;
      r_151__13_ <= r_n_151__13_;
      r_151__12_ <= r_n_151__12_;
      r_151__11_ <= r_n_151__11_;
      r_151__10_ <= r_n_151__10_;
      r_151__9_ <= r_n_151__9_;
      r_151__8_ <= r_n_151__8_;
      r_151__7_ <= r_n_151__7_;
      r_151__6_ <= r_n_151__6_;
      r_151__5_ <= r_n_151__5_;
      r_151__4_ <= r_n_151__4_;
      r_151__3_ <= r_n_151__3_;
      r_151__2_ <= r_n_151__2_;
      r_151__1_ <= r_n_151__1_;
      r_151__0_ <= r_n_151__0_;
    end 
    if(N1944) begin
      r_152__31_ <= r_n_152__31_;
      r_152__30_ <= r_n_152__30_;
      r_152__29_ <= r_n_152__29_;
      r_152__28_ <= r_n_152__28_;
      r_152__27_ <= r_n_152__27_;
      r_152__26_ <= r_n_152__26_;
      r_152__25_ <= r_n_152__25_;
      r_152__24_ <= r_n_152__24_;
      r_152__23_ <= r_n_152__23_;
      r_152__22_ <= r_n_152__22_;
      r_152__21_ <= r_n_152__21_;
      r_152__20_ <= r_n_152__20_;
      r_152__19_ <= r_n_152__19_;
      r_152__18_ <= r_n_152__18_;
      r_152__17_ <= r_n_152__17_;
      r_152__16_ <= r_n_152__16_;
      r_152__15_ <= r_n_152__15_;
      r_152__14_ <= r_n_152__14_;
      r_152__13_ <= r_n_152__13_;
      r_152__12_ <= r_n_152__12_;
      r_152__11_ <= r_n_152__11_;
      r_152__10_ <= r_n_152__10_;
      r_152__9_ <= r_n_152__9_;
      r_152__8_ <= r_n_152__8_;
      r_152__7_ <= r_n_152__7_;
      r_152__6_ <= r_n_152__6_;
      r_152__5_ <= r_n_152__5_;
      r_152__4_ <= r_n_152__4_;
      r_152__3_ <= r_n_152__3_;
      r_152__2_ <= r_n_152__2_;
      r_152__1_ <= r_n_152__1_;
      r_152__0_ <= r_n_152__0_;
    end 
    if(N1945) begin
      r_153__31_ <= r_n_153__31_;
      r_153__30_ <= r_n_153__30_;
      r_153__29_ <= r_n_153__29_;
      r_153__28_ <= r_n_153__28_;
      r_153__27_ <= r_n_153__27_;
      r_153__26_ <= r_n_153__26_;
      r_153__25_ <= r_n_153__25_;
      r_153__24_ <= r_n_153__24_;
      r_153__23_ <= r_n_153__23_;
      r_153__22_ <= r_n_153__22_;
      r_153__21_ <= r_n_153__21_;
      r_153__20_ <= r_n_153__20_;
      r_153__19_ <= r_n_153__19_;
      r_153__18_ <= r_n_153__18_;
      r_153__17_ <= r_n_153__17_;
      r_153__16_ <= r_n_153__16_;
      r_153__15_ <= r_n_153__15_;
      r_153__14_ <= r_n_153__14_;
      r_153__13_ <= r_n_153__13_;
      r_153__12_ <= r_n_153__12_;
      r_153__11_ <= r_n_153__11_;
      r_153__10_ <= r_n_153__10_;
      r_153__9_ <= r_n_153__9_;
      r_153__8_ <= r_n_153__8_;
      r_153__7_ <= r_n_153__7_;
      r_153__6_ <= r_n_153__6_;
      r_153__5_ <= r_n_153__5_;
      r_153__4_ <= r_n_153__4_;
      r_153__3_ <= r_n_153__3_;
      r_153__2_ <= r_n_153__2_;
      r_153__1_ <= r_n_153__1_;
      r_153__0_ <= r_n_153__0_;
    end 
    if(N1946) begin
      r_154__31_ <= r_n_154__31_;
      r_154__30_ <= r_n_154__30_;
      r_154__29_ <= r_n_154__29_;
      r_154__28_ <= r_n_154__28_;
      r_154__27_ <= r_n_154__27_;
      r_154__26_ <= r_n_154__26_;
      r_154__25_ <= r_n_154__25_;
      r_154__24_ <= r_n_154__24_;
      r_154__23_ <= r_n_154__23_;
      r_154__22_ <= r_n_154__22_;
      r_154__21_ <= r_n_154__21_;
      r_154__20_ <= r_n_154__20_;
      r_154__19_ <= r_n_154__19_;
      r_154__18_ <= r_n_154__18_;
      r_154__17_ <= r_n_154__17_;
      r_154__16_ <= r_n_154__16_;
      r_154__15_ <= r_n_154__15_;
      r_154__14_ <= r_n_154__14_;
      r_154__13_ <= r_n_154__13_;
      r_154__12_ <= r_n_154__12_;
      r_154__11_ <= r_n_154__11_;
      r_154__10_ <= r_n_154__10_;
      r_154__9_ <= r_n_154__9_;
      r_154__8_ <= r_n_154__8_;
      r_154__7_ <= r_n_154__7_;
      r_154__6_ <= r_n_154__6_;
      r_154__5_ <= r_n_154__5_;
      r_154__4_ <= r_n_154__4_;
      r_154__3_ <= r_n_154__3_;
      r_154__2_ <= r_n_154__2_;
      r_154__1_ <= r_n_154__1_;
      r_154__0_ <= r_n_154__0_;
    end 
    if(N1947) begin
      r_155__31_ <= r_n_155__31_;
      r_155__30_ <= r_n_155__30_;
      r_155__29_ <= r_n_155__29_;
      r_155__28_ <= r_n_155__28_;
      r_155__27_ <= r_n_155__27_;
      r_155__26_ <= r_n_155__26_;
      r_155__25_ <= r_n_155__25_;
      r_155__24_ <= r_n_155__24_;
      r_155__23_ <= r_n_155__23_;
      r_155__22_ <= r_n_155__22_;
      r_155__21_ <= r_n_155__21_;
      r_155__20_ <= r_n_155__20_;
      r_155__19_ <= r_n_155__19_;
      r_155__18_ <= r_n_155__18_;
      r_155__17_ <= r_n_155__17_;
      r_155__16_ <= r_n_155__16_;
      r_155__15_ <= r_n_155__15_;
      r_155__14_ <= r_n_155__14_;
      r_155__13_ <= r_n_155__13_;
      r_155__12_ <= r_n_155__12_;
      r_155__11_ <= r_n_155__11_;
      r_155__10_ <= r_n_155__10_;
      r_155__9_ <= r_n_155__9_;
      r_155__8_ <= r_n_155__8_;
      r_155__7_ <= r_n_155__7_;
      r_155__6_ <= r_n_155__6_;
      r_155__5_ <= r_n_155__5_;
      r_155__4_ <= r_n_155__4_;
      r_155__3_ <= r_n_155__3_;
      r_155__2_ <= r_n_155__2_;
      r_155__1_ <= r_n_155__1_;
      r_155__0_ <= r_n_155__0_;
    end 
    if(N1948) begin
      r_156__31_ <= r_n_156__31_;
      r_156__30_ <= r_n_156__30_;
      r_156__29_ <= r_n_156__29_;
      r_156__28_ <= r_n_156__28_;
      r_156__27_ <= r_n_156__27_;
      r_156__26_ <= r_n_156__26_;
      r_156__25_ <= r_n_156__25_;
      r_156__24_ <= r_n_156__24_;
      r_156__23_ <= r_n_156__23_;
      r_156__22_ <= r_n_156__22_;
      r_156__21_ <= r_n_156__21_;
      r_156__20_ <= r_n_156__20_;
      r_156__19_ <= r_n_156__19_;
      r_156__18_ <= r_n_156__18_;
      r_156__17_ <= r_n_156__17_;
      r_156__16_ <= r_n_156__16_;
      r_156__15_ <= r_n_156__15_;
      r_156__14_ <= r_n_156__14_;
      r_156__13_ <= r_n_156__13_;
      r_156__12_ <= r_n_156__12_;
      r_156__11_ <= r_n_156__11_;
      r_156__10_ <= r_n_156__10_;
      r_156__9_ <= r_n_156__9_;
      r_156__8_ <= r_n_156__8_;
      r_156__7_ <= r_n_156__7_;
      r_156__6_ <= r_n_156__6_;
      r_156__5_ <= r_n_156__5_;
      r_156__4_ <= r_n_156__4_;
      r_156__3_ <= r_n_156__3_;
      r_156__2_ <= r_n_156__2_;
      r_156__1_ <= r_n_156__1_;
      r_156__0_ <= r_n_156__0_;
    end 
    if(N1949) begin
      r_157__31_ <= r_n_157__31_;
      r_157__30_ <= r_n_157__30_;
      r_157__29_ <= r_n_157__29_;
      r_157__28_ <= r_n_157__28_;
      r_157__27_ <= r_n_157__27_;
      r_157__26_ <= r_n_157__26_;
      r_157__25_ <= r_n_157__25_;
      r_157__24_ <= r_n_157__24_;
      r_157__23_ <= r_n_157__23_;
      r_157__22_ <= r_n_157__22_;
      r_157__21_ <= r_n_157__21_;
      r_157__20_ <= r_n_157__20_;
      r_157__19_ <= r_n_157__19_;
      r_157__18_ <= r_n_157__18_;
      r_157__17_ <= r_n_157__17_;
      r_157__16_ <= r_n_157__16_;
      r_157__15_ <= r_n_157__15_;
      r_157__14_ <= r_n_157__14_;
      r_157__13_ <= r_n_157__13_;
      r_157__12_ <= r_n_157__12_;
      r_157__11_ <= r_n_157__11_;
      r_157__10_ <= r_n_157__10_;
      r_157__9_ <= r_n_157__9_;
      r_157__8_ <= r_n_157__8_;
      r_157__7_ <= r_n_157__7_;
      r_157__6_ <= r_n_157__6_;
      r_157__5_ <= r_n_157__5_;
      r_157__4_ <= r_n_157__4_;
      r_157__3_ <= r_n_157__3_;
      r_157__2_ <= r_n_157__2_;
      r_157__1_ <= r_n_157__1_;
      r_157__0_ <= r_n_157__0_;
    end 
    if(N1950) begin
      r_158__31_ <= r_n_158__31_;
      r_158__30_ <= r_n_158__30_;
      r_158__29_ <= r_n_158__29_;
      r_158__28_ <= r_n_158__28_;
      r_158__27_ <= r_n_158__27_;
      r_158__26_ <= r_n_158__26_;
      r_158__25_ <= r_n_158__25_;
      r_158__24_ <= r_n_158__24_;
      r_158__23_ <= r_n_158__23_;
      r_158__22_ <= r_n_158__22_;
      r_158__21_ <= r_n_158__21_;
      r_158__20_ <= r_n_158__20_;
      r_158__19_ <= r_n_158__19_;
      r_158__18_ <= r_n_158__18_;
      r_158__17_ <= r_n_158__17_;
      r_158__16_ <= r_n_158__16_;
      r_158__15_ <= r_n_158__15_;
      r_158__14_ <= r_n_158__14_;
      r_158__13_ <= r_n_158__13_;
      r_158__12_ <= r_n_158__12_;
      r_158__11_ <= r_n_158__11_;
      r_158__10_ <= r_n_158__10_;
      r_158__9_ <= r_n_158__9_;
      r_158__8_ <= r_n_158__8_;
      r_158__7_ <= r_n_158__7_;
      r_158__6_ <= r_n_158__6_;
      r_158__5_ <= r_n_158__5_;
      r_158__4_ <= r_n_158__4_;
      r_158__3_ <= r_n_158__3_;
      r_158__2_ <= r_n_158__2_;
      r_158__1_ <= r_n_158__1_;
      r_158__0_ <= r_n_158__0_;
    end 
    if(N1951) begin
      r_159__31_ <= r_n_159__31_;
      r_159__30_ <= r_n_159__30_;
      r_159__29_ <= r_n_159__29_;
      r_159__28_ <= r_n_159__28_;
      r_159__27_ <= r_n_159__27_;
      r_159__26_ <= r_n_159__26_;
      r_159__25_ <= r_n_159__25_;
      r_159__24_ <= r_n_159__24_;
      r_159__23_ <= r_n_159__23_;
      r_159__22_ <= r_n_159__22_;
      r_159__21_ <= r_n_159__21_;
      r_159__20_ <= r_n_159__20_;
      r_159__19_ <= r_n_159__19_;
      r_159__18_ <= r_n_159__18_;
      r_159__17_ <= r_n_159__17_;
      r_159__16_ <= r_n_159__16_;
      r_159__15_ <= r_n_159__15_;
      r_159__14_ <= r_n_159__14_;
      r_159__13_ <= r_n_159__13_;
      r_159__12_ <= r_n_159__12_;
      r_159__11_ <= r_n_159__11_;
      r_159__10_ <= r_n_159__10_;
      r_159__9_ <= r_n_159__9_;
      r_159__8_ <= r_n_159__8_;
      r_159__7_ <= r_n_159__7_;
      r_159__6_ <= r_n_159__6_;
      r_159__5_ <= r_n_159__5_;
      r_159__4_ <= r_n_159__4_;
      r_159__3_ <= r_n_159__3_;
      r_159__2_ <= r_n_159__2_;
      r_159__1_ <= r_n_159__1_;
      r_159__0_ <= r_n_159__0_;
    end 
    if(N1952) begin
      r_160__31_ <= r_n_160__31_;
      r_160__30_ <= r_n_160__30_;
      r_160__29_ <= r_n_160__29_;
      r_160__28_ <= r_n_160__28_;
      r_160__27_ <= r_n_160__27_;
      r_160__26_ <= r_n_160__26_;
      r_160__25_ <= r_n_160__25_;
      r_160__24_ <= r_n_160__24_;
      r_160__23_ <= r_n_160__23_;
      r_160__22_ <= r_n_160__22_;
      r_160__21_ <= r_n_160__21_;
      r_160__20_ <= r_n_160__20_;
      r_160__19_ <= r_n_160__19_;
      r_160__18_ <= r_n_160__18_;
      r_160__17_ <= r_n_160__17_;
      r_160__16_ <= r_n_160__16_;
      r_160__15_ <= r_n_160__15_;
      r_160__14_ <= r_n_160__14_;
      r_160__13_ <= r_n_160__13_;
      r_160__12_ <= r_n_160__12_;
      r_160__11_ <= r_n_160__11_;
      r_160__10_ <= r_n_160__10_;
      r_160__9_ <= r_n_160__9_;
      r_160__8_ <= r_n_160__8_;
      r_160__7_ <= r_n_160__7_;
      r_160__6_ <= r_n_160__6_;
      r_160__5_ <= r_n_160__5_;
      r_160__4_ <= r_n_160__4_;
      r_160__3_ <= r_n_160__3_;
      r_160__2_ <= r_n_160__2_;
      r_160__1_ <= r_n_160__1_;
      r_160__0_ <= r_n_160__0_;
    end 
    if(N1953) begin
      r_161__31_ <= r_n_161__31_;
      r_161__30_ <= r_n_161__30_;
      r_161__29_ <= r_n_161__29_;
      r_161__28_ <= r_n_161__28_;
      r_161__27_ <= r_n_161__27_;
      r_161__26_ <= r_n_161__26_;
      r_161__25_ <= r_n_161__25_;
      r_161__24_ <= r_n_161__24_;
      r_161__23_ <= r_n_161__23_;
      r_161__22_ <= r_n_161__22_;
      r_161__21_ <= r_n_161__21_;
      r_161__20_ <= r_n_161__20_;
      r_161__19_ <= r_n_161__19_;
      r_161__18_ <= r_n_161__18_;
      r_161__17_ <= r_n_161__17_;
      r_161__16_ <= r_n_161__16_;
      r_161__15_ <= r_n_161__15_;
      r_161__14_ <= r_n_161__14_;
      r_161__13_ <= r_n_161__13_;
      r_161__12_ <= r_n_161__12_;
      r_161__11_ <= r_n_161__11_;
      r_161__10_ <= r_n_161__10_;
      r_161__9_ <= r_n_161__9_;
      r_161__8_ <= r_n_161__8_;
      r_161__7_ <= r_n_161__7_;
      r_161__6_ <= r_n_161__6_;
      r_161__5_ <= r_n_161__5_;
      r_161__4_ <= r_n_161__4_;
      r_161__3_ <= r_n_161__3_;
      r_161__2_ <= r_n_161__2_;
      r_161__1_ <= r_n_161__1_;
      r_161__0_ <= r_n_161__0_;
    end 
    if(N1954) begin
      r_162__31_ <= r_n_162__31_;
      r_162__30_ <= r_n_162__30_;
      r_162__29_ <= r_n_162__29_;
      r_162__28_ <= r_n_162__28_;
      r_162__27_ <= r_n_162__27_;
      r_162__26_ <= r_n_162__26_;
      r_162__25_ <= r_n_162__25_;
      r_162__24_ <= r_n_162__24_;
      r_162__23_ <= r_n_162__23_;
      r_162__22_ <= r_n_162__22_;
      r_162__21_ <= r_n_162__21_;
      r_162__20_ <= r_n_162__20_;
      r_162__19_ <= r_n_162__19_;
      r_162__18_ <= r_n_162__18_;
      r_162__17_ <= r_n_162__17_;
      r_162__16_ <= r_n_162__16_;
      r_162__15_ <= r_n_162__15_;
      r_162__14_ <= r_n_162__14_;
      r_162__13_ <= r_n_162__13_;
      r_162__12_ <= r_n_162__12_;
      r_162__11_ <= r_n_162__11_;
      r_162__10_ <= r_n_162__10_;
      r_162__9_ <= r_n_162__9_;
      r_162__8_ <= r_n_162__8_;
      r_162__7_ <= r_n_162__7_;
      r_162__6_ <= r_n_162__6_;
      r_162__5_ <= r_n_162__5_;
      r_162__4_ <= r_n_162__4_;
      r_162__3_ <= r_n_162__3_;
      r_162__2_ <= r_n_162__2_;
      r_162__1_ <= r_n_162__1_;
      r_162__0_ <= r_n_162__0_;
    end 
    if(N1955) begin
      r_163__31_ <= r_n_163__31_;
      r_163__30_ <= r_n_163__30_;
      r_163__29_ <= r_n_163__29_;
      r_163__28_ <= r_n_163__28_;
      r_163__27_ <= r_n_163__27_;
      r_163__26_ <= r_n_163__26_;
      r_163__25_ <= r_n_163__25_;
      r_163__24_ <= r_n_163__24_;
      r_163__23_ <= r_n_163__23_;
      r_163__22_ <= r_n_163__22_;
      r_163__21_ <= r_n_163__21_;
      r_163__20_ <= r_n_163__20_;
      r_163__19_ <= r_n_163__19_;
      r_163__18_ <= r_n_163__18_;
      r_163__17_ <= r_n_163__17_;
      r_163__16_ <= r_n_163__16_;
      r_163__15_ <= r_n_163__15_;
      r_163__14_ <= r_n_163__14_;
      r_163__13_ <= r_n_163__13_;
      r_163__12_ <= r_n_163__12_;
      r_163__11_ <= r_n_163__11_;
      r_163__10_ <= r_n_163__10_;
      r_163__9_ <= r_n_163__9_;
      r_163__8_ <= r_n_163__8_;
      r_163__7_ <= r_n_163__7_;
      r_163__6_ <= r_n_163__6_;
      r_163__5_ <= r_n_163__5_;
      r_163__4_ <= r_n_163__4_;
      r_163__3_ <= r_n_163__3_;
      r_163__2_ <= r_n_163__2_;
      r_163__1_ <= r_n_163__1_;
      r_163__0_ <= r_n_163__0_;
    end 
    if(N1956) begin
      r_164__31_ <= r_n_164__31_;
      r_164__30_ <= r_n_164__30_;
      r_164__29_ <= r_n_164__29_;
      r_164__28_ <= r_n_164__28_;
      r_164__27_ <= r_n_164__27_;
      r_164__26_ <= r_n_164__26_;
      r_164__25_ <= r_n_164__25_;
      r_164__24_ <= r_n_164__24_;
      r_164__23_ <= r_n_164__23_;
      r_164__22_ <= r_n_164__22_;
      r_164__21_ <= r_n_164__21_;
      r_164__20_ <= r_n_164__20_;
      r_164__19_ <= r_n_164__19_;
      r_164__18_ <= r_n_164__18_;
      r_164__17_ <= r_n_164__17_;
      r_164__16_ <= r_n_164__16_;
      r_164__15_ <= r_n_164__15_;
      r_164__14_ <= r_n_164__14_;
      r_164__13_ <= r_n_164__13_;
      r_164__12_ <= r_n_164__12_;
      r_164__11_ <= r_n_164__11_;
      r_164__10_ <= r_n_164__10_;
      r_164__9_ <= r_n_164__9_;
      r_164__8_ <= r_n_164__8_;
      r_164__7_ <= r_n_164__7_;
      r_164__6_ <= r_n_164__6_;
      r_164__5_ <= r_n_164__5_;
      r_164__4_ <= r_n_164__4_;
      r_164__3_ <= r_n_164__3_;
      r_164__2_ <= r_n_164__2_;
      r_164__1_ <= r_n_164__1_;
      r_164__0_ <= r_n_164__0_;
    end 
    if(N1957) begin
      r_165__31_ <= r_n_165__31_;
      r_165__30_ <= r_n_165__30_;
      r_165__29_ <= r_n_165__29_;
      r_165__28_ <= r_n_165__28_;
      r_165__27_ <= r_n_165__27_;
      r_165__26_ <= r_n_165__26_;
      r_165__25_ <= r_n_165__25_;
      r_165__24_ <= r_n_165__24_;
      r_165__23_ <= r_n_165__23_;
      r_165__22_ <= r_n_165__22_;
      r_165__21_ <= r_n_165__21_;
      r_165__20_ <= r_n_165__20_;
      r_165__19_ <= r_n_165__19_;
      r_165__18_ <= r_n_165__18_;
      r_165__17_ <= r_n_165__17_;
      r_165__16_ <= r_n_165__16_;
      r_165__15_ <= r_n_165__15_;
      r_165__14_ <= r_n_165__14_;
      r_165__13_ <= r_n_165__13_;
      r_165__12_ <= r_n_165__12_;
      r_165__11_ <= r_n_165__11_;
      r_165__10_ <= r_n_165__10_;
      r_165__9_ <= r_n_165__9_;
      r_165__8_ <= r_n_165__8_;
      r_165__7_ <= r_n_165__7_;
      r_165__6_ <= r_n_165__6_;
      r_165__5_ <= r_n_165__5_;
      r_165__4_ <= r_n_165__4_;
      r_165__3_ <= r_n_165__3_;
      r_165__2_ <= r_n_165__2_;
      r_165__1_ <= r_n_165__1_;
      r_165__0_ <= r_n_165__0_;
    end 
    if(N1958) begin
      r_166__31_ <= r_n_166__31_;
      r_166__30_ <= r_n_166__30_;
      r_166__29_ <= r_n_166__29_;
      r_166__28_ <= r_n_166__28_;
      r_166__27_ <= r_n_166__27_;
      r_166__26_ <= r_n_166__26_;
      r_166__25_ <= r_n_166__25_;
      r_166__24_ <= r_n_166__24_;
      r_166__23_ <= r_n_166__23_;
      r_166__22_ <= r_n_166__22_;
      r_166__21_ <= r_n_166__21_;
      r_166__20_ <= r_n_166__20_;
      r_166__19_ <= r_n_166__19_;
      r_166__18_ <= r_n_166__18_;
      r_166__17_ <= r_n_166__17_;
      r_166__16_ <= r_n_166__16_;
      r_166__15_ <= r_n_166__15_;
      r_166__14_ <= r_n_166__14_;
      r_166__13_ <= r_n_166__13_;
      r_166__12_ <= r_n_166__12_;
      r_166__11_ <= r_n_166__11_;
      r_166__10_ <= r_n_166__10_;
      r_166__9_ <= r_n_166__9_;
      r_166__8_ <= r_n_166__8_;
      r_166__7_ <= r_n_166__7_;
      r_166__6_ <= r_n_166__6_;
      r_166__5_ <= r_n_166__5_;
      r_166__4_ <= r_n_166__4_;
      r_166__3_ <= r_n_166__3_;
      r_166__2_ <= r_n_166__2_;
      r_166__1_ <= r_n_166__1_;
      r_166__0_ <= r_n_166__0_;
    end 
    if(N1959) begin
      r_167__31_ <= r_n_167__31_;
      r_167__30_ <= r_n_167__30_;
      r_167__29_ <= r_n_167__29_;
      r_167__28_ <= r_n_167__28_;
      r_167__27_ <= r_n_167__27_;
      r_167__26_ <= r_n_167__26_;
      r_167__25_ <= r_n_167__25_;
      r_167__24_ <= r_n_167__24_;
      r_167__23_ <= r_n_167__23_;
      r_167__22_ <= r_n_167__22_;
      r_167__21_ <= r_n_167__21_;
      r_167__20_ <= r_n_167__20_;
      r_167__19_ <= r_n_167__19_;
      r_167__18_ <= r_n_167__18_;
      r_167__17_ <= r_n_167__17_;
      r_167__16_ <= r_n_167__16_;
      r_167__15_ <= r_n_167__15_;
      r_167__14_ <= r_n_167__14_;
      r_167__13_ <= r_n_167__13_;
      r_167__12_ <= r_n_167__12_;
      r_167__11_ <= r_n_167__11_;
      r_167__10_ <= r_n_167__10_;
      r_167__9_ <= r_n_167__9_;
      r_167__8_ <= r_n_167__8_;
      r_167__7_ <= r_n_167__7_;
      r_167__6_ <= r_n_167__6_;
      r_167__5_ <= r_n_167__5_;
      r_167__4_ <= r_n_167__4_;
      r_167__3_ <= r_n_167__3_;
      r_167__2_ <= r_n_167__2_;
      r_167__1_ <= r_n_167__1_;
      r_167__0_ <= r_n_167__0_;
    end 
    if(N1960) begin
      r_168__31_ <= r_n_168__31_;
      r_168__30_ <= r_n_168__30_;
      r_168__29_ <= r_n_168__29_;
      r_168__28_ <= r_n_168__28_;
      r_168__27_ <= r_n_168__27_;
      r_168__26_ <= r_n_168__26_;
      r_168__25_ <= r_n_168__25_;
      r_168__24_ <= r_n_168__24_;
      r_168__23_ <= r_n_168__23_;
      r_168__22_ <= r_n_168__22_;
      r_168__21_ <= r_n_168__21_;
      r_168__20_ <= r_n_168__20_;
      r_168__19_ <= r_n_168__19_;
      r_168__18_ <= r_n_168__18_;
      r_168__17_ <= r_n_168__17_;
      r_168__16_ <= r_n_168__16_;
      r_168__15_ <= r_n_168__15_;
      r_168__14_ <= r_n_168__14_;
      r_168__13_ <= r_n_168__13_;
      r_168__12_ <= r_n_168__12_;
      r_168__11_ <= r_n_168__11_;
      r_168__10_ <= r_n_168__10_;
      r_168__9_ <= r_n_168__9_;
      r_168__8_ <= r_n_168__8_;
      r_168__7_ <= r_n_168__7_;
      r_168__6_ <= r_n_168__6_;
      r_168__5_ <= r_n_168__5_;
      r_168__4_ <= r_n_168__4_;
      r_168__3_ <= r_n_168__3_;
      r_168__2_ <= r_n_168__2_;
      r_168__1_ <= r_n_168__1_;
      r_168__0_ <= r_n_168__0_;
    end 
    if(N1961) begin
      r_169__31_ <= r_n_169__31_;
      r_169__30_ <= r_n_169__30_;
      r_169__29_ <= r_n_169__29_;
      r_169__28_ <= r_n_169__28_;
      r_169__27_ <= r_n_169__27_;
      r_169__26_ <= r_n_169__26_;
      r_169__25_ <= r_n_169__25_;
      r_169__24_ <= r_n_169__24_;
      r_169__23_ <= r_n_169__23_;
      r_169__22_ <= r_n_169__22_;
      r_169__21_ <= r_n_169__21_;
      r_169__20_ <= r_n_169__20_;
      r_169__19_ <= r_n_169__19_;
      r_169__18_ <= r_n_169__18_;
      r_169__17_ <= r_n_169__17_;
      r_169__16_ <= r_n_169__16_;
      r_169__15_ <= r_n_169__15_;
      r_169__14_ <= r_n_169__14_;
      r_169__13_ <= r_n_169__13_;
      r_169__12_ <= r_n_169__12_;
      r_169__11_ <= r_n_169__11_;
      r_169__10_ <= r_n_169__10_;
      r_169__9_ <= r_n_169__9_;
      r_169__8_ <= r_n_169__8_;
      r_169__7_ <= r_n_169__7_;
      r_169__6_ <= r_n_169__6_;
      r_169__5_ <= r_n_169__5_;
      r_169__4_ <= r_n_169__4_;
      r_169__3_ <= r_n_169__3_;
      r_169__2_ <= r_n_169__2_;
      r_169__1_ <= r_n_169__1_;
      r_169__0_ <= r_n_169__0_;
    end 
    if(N1962) begin
      r_170__31_ <= r_n_170__31_;
      r_170__30_ <= r_n_170__30_;
      r_170__29_ <= r_n_170__29_;
      r_170__28_ <= r_n_170__28_;
      r_170__27_ <= r_n_170__27_;
      r_170__26_ <= r_n_170__26_;
      r_170__25_ <= r_n_170__25_;
      r_170__24_ <= r_n_170__24_;
      r_170__23_ <= r_n_170__23_;
      r_170__22_ <= r_n_170__22_;
      r_170__21_ <= r_n_170__21_;
      r_170__20_ <= r_n_170__20_;
      r_170__19_ <= r_n_170__19_;
      r_170__18_ <= r_n_170__18_;
      r_170__17_ <= r_n_170__17_;
      r_170__16_ <= r_n_170__16_;
      r_170__15_ <= r_n_170__15_;
      r_170__14_ <= r_n_170__14_;
      r_170__13_ <= r_n_170__13_;
      r_170__12_ <= r_n_170__12_;
      r_170__11_ <= r_n_170__11_;
      r_170__10_ <= r_n_170__10_;
      r_170__9_ <= r_n_170__9_;
      r_170__8_ <= r_n_170__8_;
      r_170__7_ <= r_n_170__7_;
      r_170__6_ <= r_n_170__6_;
      r_170__5_ <= r_n_170__5_;
      r_170__4_ <= r_n_170__4_;
      r_170__3_ <= r_n_170__3_;
      r_170__2_ <= r_n_170__2_;
      r_170__1_ <= r_n_170__1_;
      r_170__0_ <= r_n_170__0_;
    end 
    if(N1963) begin
      r_171__31_ <= r_n_171__31_;
      r_171__30_ <= r_n_171__30_;
      r_171__29_ <= r_n_171__29_;
      r_171__28_ <= r_n_171__28_;
      r_171__27_ <= r_n_171__27_;
      r_171__26_ <= r_n_171__26_;
      r_171__25_ <= r_n_171__25_;
      r_171__24_ <= r_n_171__24_;
      r_171__23_ <= r_n_171__23_;
      r_171__22_ <= r_n_171__22_;
      r_171__21_ <= r_n_171__21_;
      r_171__20_ <= r_n_171__20_;
      r_171__19_ <= r_n_171__19_;
      r_171__18_ <= r_n_171__18_;
      r_171__17_ <= r_n_171__17_;
      r_171__16_ <= r_n_171__16_;
      r_171__15_ <= r_n_171__15_;
      r_171__14_ <= r_n_171__14_;
      r_171__13_ <= r_n_171__13_;
      r_171__12_ <= r_n_171__12_;
      r_171__11_ <= r_n_171__11_;
      r_171__10_ <= r_n_171__10_;
      r_171__9_ <= r_n_171__9_;
      r_171__8_ <= r_n_171__8_;
      r_171__7_ <= r_n_171__7_;
      r_171__6_ <= r_n_171__6_;
      r_171__5_ <= r_n_171__5_;
      r_171__4_ <= r_n_171__4_;
      r_171__3_ <= r_n_171__3_;
      r_171__2_ <= r_n_171__2_;
      r_171__1_ <= r_n_171__1_;
      r_171__0_ <= r_n_171__0_;
    end 
    if(N1964) begin
      r_172__31_ <= r_n_172__31_;
      r_172__30_ <= r_n_172__30_;
      r_172__29_ <= r_n_172__29_;
      r_172__28_ <= r_n_172__28_;
      r_172__27_ <= r_n_172__27_;
      r_172__26_ <= r_n_172__26_;
      r_172__25_ <= r_n_172__25_;
      r_172__24_ <= r_n_172__24_;
      r_172__23_ <= r_n_172__23_;
      r_172__22_ <= r_n_172__22_;
      r_172__21_ <= r_n_172__21_;
      r_172__20_ <= r_n_172__20_;
      r_172__19_ <= r_n_172__19_;
      r_172__18_ <= r_n_172__18_;
      r_172__17_ <= r_n_172__17_;
      r_172__16_ <= r_n_172__16_;
      r_172__15_ <= r_n_172__15_;
      r_172__14_ <= r_n_172__14_;
      r_172__13_ <= r_n_172__13_;
      r_172__12_ <= r_n_172__12_;
      r_172__11_ <= r_n_172__11_;
      r_172__10_ <= r_n_172__10_;
      r_172__9_ <= r_n_172__9_;
      r_172__8_ <= r_n_172__8_;
      r_172__7_ <= r_n_172__7_;
      r_172__6_ <= r_n_172__6_;
      r_172__5_ <= r_n_172__5_;
      r_172__4_ <= r_n_172__4_;
      r_172__3_ <= r_n_172__3_;
      r_172__2_ <= r_n_172__2_;
      r_172__1_ <= r_n_172__1_;
      r_172__0_ <= r_n_172__0_;
    end 
    if(N1965) begin
      r_173__31_ <= r_n_173__31_;
      r_173__30_ <= r_n_173__30_;
      r_173__29_ <= r_n_173__29_;
      r_173__28_ <= r_n_173__28_;
      r_173__27_ <= r_n_173__27_;
      r_173__26_ <= r_n_173__26_;
      r_173__25_ <= r_n_173__25_;
      r_173__24_ <= r_n_173__24_;
      r_173__23_ <= r_n_173__23_;
      r_173__22_ <= r_n_173__22_;
      r_173__21_ <= r_n_173__21_;
      r_173__20_ <= r_n_173__20_;
      r_173__19_ <= r_n_173__19_;
      r_173__18_ <= r_n_173__18_;
      r_173__17_ <= r_n_173__17_;
      r_173__16_ <= r_n_173__16_;
      r_173__15_ <= r_n_173__15_;
      r_173__14_ <= r_n_173__14_;
      r_173__13_ <= r_n_173__13_;
      r_173__12_ <= r_n_173__12_;
      r_173__11_ <= r_n_173__11_;
      r_173__10_ <= r_n_173__10_;
      r_173__9_ <= r_n_173__9_;
      r_173__8_ <= r_n_173__8_;
      r_173__7_ <= r_n_173__7_;
      r_173__6_ <= r_n_173__6_;
      r_173__5_ <= r_n_173__5_;
      r_173__4_ <= r_n_173__4_;
      r_173__3_ <= r_n_173__3_;
      r_173__2_ <= r_n_173__2_;
      r_173__1_ <= r_n_173__1_;
      r_173__0_ <= r_n_173__0_;
    end 
    if(N1966) begin
      r_174__31_ <= r_n_174__31_;
      r_174__30_ <= r_n_174__30_;
      r_174__29_ <= r_n_174__29_;
      r_174__28_ <= r_n_174__28_;
      r_174__27_ <= r_n_174__27_;
      r_174__26_ <= r_n_174__26_;
      r_174__25_ <= r_n_174__25_;
      r_174__24_ <= r_n_174__24_;
      r_174__23_ <= r_n_174__23_;
      r_174__22_ <= r_n_174__22_;
      r_174__21_ <= r_n_174__21_;
      r_174__20_ <= r_n_174__20_;
      r_174__19_ <= r_n_174__19_;
      r_174__18_ <= r_n_174__18_;
      r_174__17_ <= r_n_174__17_;
      r_174__16_ <= r_n_174__16_;
      r_174__15_ <= r_n_174__15_;
      r_174__14_ <= r_n_174__14_;
      r_174__13_ <= r_n_174__13_;
      r_174__12_ <= r_n_174__12_;
      r_174__11_ <= r_n_174__11_;
      r_174__10_ <= r_n_174__10_;
      r_174__9_ <= r_n_174__9_;
      r_174__8_ <= r_n_174__8_;
      r_174__7_ <= r_n_174__7_;
      r_174__6_ <= r_n_174__6_;
      r_174__5_ <= r_n_174__5_;
      r_174__4_ <= r_n_174__4_;
      r_174__3_ <= r_n_174__3_;
      r_174__2_ <= r_n_174__2_;
      r_174__1_ <= r_n_174__1_;
      r_174__0_ <= r_n_174__0_;
    end 
    if(N1967) begin
      r_175__31_ <= r_n_175__31_;
      r_175__30_ <= r_n_175__30_;
      r_175__29_ <= r_n_175__29_;
      r_175__28_ <= r_n_175__28_;
      r_175__27_ <= r_n_175__27_;
      r_175__26_ <= r_n_175__26_;
      r_175__25_ <= r_n_175__25_;
      r_175__24_ <= r_n_175__24_;
      r_175__23_ <= r_n_175__23_;
      r_175__22_ <= r_n_175__22_;
      r_175__21_ <= r_n_175__21_;
      r_175__20_ <= r_n_175__20_;
      r_175__19_ <= r_n_175__19_;
      r_175__18_ <= r_n_175__18_;
      r_175__17_ <= r_n_175__17_;
      r_175__16_ <= r_n_175__16_;
      r_175__15_ <= r_n_175__15_;
      r_175__14_ <= r_n_175__14_;
      r_175__13_ <= r_n_175__13_;
      r_175__12_ <= r_n_175__12_;
      r_175__11_ <= r_n_175__11_;
      r_175__10_ <= r_n_175__10_;
      r_175__9_ <= r_n_175__9_;
      r_175__8_ <= r_n_175__8_;
      r_175__7_ <= r_n_175__7_;
      r_175__6_ <= r_n_175__6_;
      r_175__5_ <= r_n_175__5_;
      r_175__4_ <= r_n_175__4_;
      r_175__3_ <= r_n_175__3_;
      r_175__2_ <= r_n_175__2_;
      r_175__1_ <= r_n_175__1_;
      r_175__0_ <= r_n_175__0_;
    end 
    if(N1968) begin
      r_176__31_ <= r_n_176__31_;
      r_176__30_ <= r_n_176__30_;
      r_176__29_ <= r_n_176__29_;
      r_176__28_ <= r_n_176__28_;
      r_176__27_ <= r_n_176__27_;
      r_176__26_ <= r_n_176__26_;
      r_176__25_ <= r_n_176__25_;
      r_176__24_ <= r_n_176__24_;
      r_176__23_ <= r_n_176__23_;
      r_176__22_ <= r_n_176__22_;
      r_176__21_ <= r_n_176__21_;
      r_176__20_ <= r_n_176__20_;
      r_176__19_ <= r_n_176__19_;
      r_176__18_ <= r_n_176__18_;
      r_176__17_ <= r_n_176__17_;
      r_176__16_ <= r_n_176__16_;
      r_176__15_ <= r_n_176__15_;
      r_176__14_ <= r_n_176__14_;
      r_176__13_ <= r_n_176__13_;
      r_176__12_ <= r_n_176__12_;
      r_176__11_ <= r_n_176__11_;
      r_176__10_ <= r_n_176__10_;
      r_176__9_ <= r_n_176__9_;
      r_176__8_ <= r_n_176__8_;
      r_176__7_ <= r_n_176__7_;
      r_176__6_ <= r_n_176__6_;
      r_176__5_ <= r_n_176__5_;
      r_176__4_ <= r_n_176__4_;
      r_176__3_ <= r_n_176__3_;
      r_176__2_ <= r_n_176__2_;
      r_176__1_ <= r_n_176__1_;
      r_176__0_ <= r_n_176__0_;
    end 
    if(N1969) begin
      r_177__31_ <= r_n_177__31_;
      r_177__30_ <= r_n_177__30_;
      r_177__29_ <= r_n_177__29_;
      r_177__28_ <= r_n_177__28_;
      r_177__27_ <= r_n_177__27_;
      r_177__26_ <= r_n_177__26_;
      r_177__25_ <= r_n_177__25_;
      r_177__24_ <= r_n_177__24_;
      r_177__23_ <= r_n_177__23_;
      r_177__22_ <= r_n_177__22_;
      r_177__21_ <= r_n_177__21_;
      r_177__20_ <= r_n_177__20_;
      r_177__19_ <= r_n_177__19_;
      r_177__18_ <= r_n_177__18_;
      r_177__17_ <= r_n_177__17_;
      r_177__16_ <= r_n_177__16_;
      r_177__15_ <= r_n_177__15_;
      r_177__14_ <= r_n_177__14_;
      r_177__13_ <= r_n_177__13_;
      r_177__12_ <= r_n_177__12_;
      r_177__11_ <= r_n_177__11_;
      r_177__10_ <= r_n_177__10_;
      r_177__9_ <= r_n_177__9_;
      r_177__8_ <= r_n_177__8_;
      r_177__7_ <= r_n_177__7_;
      r_177__6_ <= r_n_177__6_;
      r_177__5_ <= r_n_177__5_;
      r_177__4_ <= r_n_177__4_;
      r_177__3_ <= r_n_177__3_;
      r_177__2_ <= r_n_177__2_;
      r_177__1_ <= r_n_177__1_;
      r_177__0_ <= r_n_177__0_;
    end 
    if(N1970) begin
      r_178__31_ <= r_n_178__31_;
      r_178__30_ <= r_n_178__30_;
      r_178__29_ <= r_n_178__29_;
      r_178__28_ <= r_n_178__28_;
      r_178__27_ <= r_n_178__27_;
      r_178__26_ <= r_n_178__26_;
      r_178__25_ <= r_n_178__25_;
      r_178__24_ <= r_n_178__24_;
      r_178__23_ <= r_n_178__23_;
      r_178__22_ <= r_n_178__22_;
      r_178__21_ <= r_n_178__21_;
      r_178__20_ <= r_n_178__20_;
      r_178__19_ <= r_n_178__19_;
      r_178__18_ <= r_n_178__18_;
      r_178__17_ <= r_n_178__17_;
      r_178__16_ <= r_n_178__16_;
      r_178__15_ <= r_n_178__15_;
      r_178__14_ <= r_n_178__14_;
      r_178__13_ <= r_n_178__13_;
      r_178__12_ <= r_n_178__12_;
      r_178__11_ <= r_n_178__11_;
      r_178__10_ <= r_n_178__10_;
      r_178__9_ <= r_n_178__9_;
      r_178__8_ <= r_n_178__8_;
      r_178__7_ <= r_n_178__7_;
      r_178__6_ <= r_n_178__6_;
      r_178__5_ <= r_n_178__5_;
      r_178__4_ <= r_n_178__4_;
      r_178__3_ <= r_n_178__3_;
      r_178__2_ <= r_n_178__2_;
      r_178__1_ <= r_n_178__1_;
      r_178__0_ <= r_n_178__0_;
    end 
    if(N1971) begin
      r_179__31_ <= r_n_179__31_;
      r_179__30_ <= r_n_179__30_;
      r_179__29_ <= r_n_179__29_;
      r_179__28_ <= r_n_179__28_;
      r_179__27_ <= r_n_179__27_;
      r_179__26_ <= r_n_179__26_;
      r_179__25_ <= r_n_179__25_;
      r_179__24_ <= r_n_179__24_;
      r_179__23_ <= r_n_179__23_;
      r_179__22_ <= r_n_179__22_;
      r_179__21_ <= r_n_179__21_;
      r_179__20_ <= r_n_179__20_;
      r_179__19_ <= r_n_179__19_;
      r_179__18_ <= r_n_179__18_;
      r_179__17_ <= r_n_179__17_;
      r_179__16_ <= r_n_179__16_;
      r_179__15_ <= r_n_179__15_;
      r_179__14_ <= r_n_179__14_;
      r_179__13_ <= r_n_179__13_;
      r_179__12_ <= r_n_179__12_;
      r_179__11_ <= r_n_179__11_;
      r_179__10_ <= r_n_179__10_;
      r_179__9_ <= r_n_179__9_;
      r_179__8_ <= r_n_179__8_;
      r_179__7_ <= r_n_179__7_;
      r_179__6_ <= r_n_179__6_;
      r_179__5_ <= r_n_179__5_;
      r_179__4_ <= r_n_179__4_;
      r_179__3_ <= r_n_179__3_;
      r_179__2_ <= r_n_179__2_;
      r_179__1_ <= r_n_179__1_;
      r_179__0_ <= r_n_179__0_;
    end 
    if(N1972) begin
      r_180__31_ <= r_n_180__31_;
      r_180__30_ <= r_n_180__30_;
      r_180__29_ <= r_n_180__29_;
      r_180__28_ <= r_n_180__28_;
      r_180__27_ <= r_n_180__27_;
      r_180__26_ <= r_n_180__26_;
      r_180__25_ <= r_n_180__25_;
      r_180__24_ <= r_n_180__24_;
      r_180__23_ <= r_n_180__23_;
      r_180__22_ <= r_n_180__22_;
      r_180__21_ <= r_n_180__21_;
      r_180__20_ <= r_n_180__20_;
      r_180__19_ <= r_n_180__19_;
      r_180__18_ <= r_n_180__18_;
      r_180__17_ <= r_n_180__17_;
      r_180__16_ <= r_n_180__16_;
      r_180__15_ <= r_n_180__15_;
      r_180__14_ <= r_n_180__14_;
      r_180__13_ <= r_n_180__13_;
      r_180__12_ <= r_n_180__12_;
      r_180__11_ <= r_n_180__11_;
      r_180__10_ <= r_n_180__10_;
      r_180__9_ <= r_n_180__9_;
      r_180__8_ <= r_n_180__8_;
      r_180__7_ <= r_n_180__7_;
      r_180__6_ <= r_n_180__6_;
      r_180__5_ <= r_n_180__5_;
      r_180__4_ <= r_n_180__4_;
      r_180__3_ <= r_n_180__3_;
      r_180__2_ <= r_n_180__2_;
      r_180__1_ <= r_n_180__1_;
      r_180__0_ <= r_n_180__0_;
    end 
    if(N1973) begin
      r_181__31_ <= r_n_181__31_;
      r_181__30_ <= r_n_181__30_;
      r_181__29_ <= r_n_181__29_;
      r_181__28_ <= r_n_181__28_;
      r_181__27_ <= r_n_181__27_;
      r_181__26_ <= r_n_181__26_;
      r_181__25_ <= r_n_181__25_;
      r_181__24_ <= r_n_181__24_;
      r_181__23_ <= r_n_181__23_;
      r_181__22_ <= r_n_181__22_;
      r_181__21_ <= r_n_181__21_;
      r_181__20_ <= r_n_181__20_;
      r_181__19_ <= r_n_181__19_;
      r_181__18_ <= r_n_181__18_;
      r_181__17_ <= r_n_181__17_;
      r_181__16_ <= r_n_181__16_;
      r_181__15_ <= r_n_181__15_;
      r_181__14_ <= r_n_181__14_;
      r_181__13_ <= r_n_181__13_;
      r_181__12_ <= r_n_181__12_;
      r_181__11_ <= r_n_181__11_;
      r_181__10_ <= r_n_181__10_;
      r_181__9_ <= r_n_181__9_;
      r_181__8_ <= r_n_181__8_;
      r_181__7_ <= r_n_181__7_;
      r_181__6_ <= r_n_181__6_;
      r_181__5_ <= r_n_181__5_;
      r_181__4_ <= r_n_181__4_;
      r_181__3_ <= r_n_181__3_;
      r_181__2_ <= r_n_181__2_;
      r_181__1_ <= r_n_181__1_;
      r_181__0_ <= r_n_181__0_;
    end 
    if(N1974) begin
      r_182__31_ <= r_n_182__31_;
      r_182__30_ <= r_n_182__30_;
      r_182__29_ <= r_n_182__29_;
      r_182__28_ <= r_n_182__28_;
      r_182__27_ <= r_n_182__27_;
      r_182__26_ <= r_n_182__26_;
      r_182__25_ <= r_n_182__25_;
      r_182__24_ <= r_n_182__24_;
      r_182__23_ <= r_n_182__23_;
      r_182__22_ <= r_n_182__22_;
      r_182__21_ <= r_n_182__21_;
      r_182__20_ <= r_n_182__20_;
      r_182__19_ <= r_n_182__19_;
      r_182__18_ <= r_n_182__18_;
      r_182__17_ <= r_n_182__17_;
      r_182__16_ <= r_n_182__16_;
      r_182__15_ <= r_n_182__15_;
      r_182__14_ <= r_n_182__14_;
      r_182__13_ <= r_n_182__13_;
      r_182__12_ <= r_n_182__12_;
      r_182__11_ <= r_n_182__11_;
      r_182__10_ <= r_n_182__10_;
      r_182__9_ <= r_n_182__9_;
      r_182__8_ <= r_n_182__8_;
      r_182__7_ <= r_n_182__7_;
      r_182__6_ <= r_n_182__6_;
      r_182__5_ <= r_n_182__5_;
      r_182__4_ <= r_n_182__4_;
      r_182__3_ <= r_n_182__3_;
      r_182__2_ <= r_n_182__2_;
      r_182__1_ <= r_n_182__1_;
      r_182__0_ <= r_n_182__0_;
    end 
    if(N1975) begin
      r_183__31_ <= r_n_183__31_;
      r_183__30_ <= r_n_183__30_;
      r_183__29_ <= r_n_183__29_;
      r_183__28_ <= r_n_183__28_;
      r_183__27_ <= r_n_183__27_;
      r_183__26_ <= r_n_183__26_;
      r_183__25_ <= r_n_183__25_;
      r_183__24_ <= r_n_183__24_;
      r_183__23_ <= r_n_183__23_;
      r_183__22_ <= r_n_183__22_;
      r_183__21_ <= r_n_183__21_;
      r_183__20_ <= r_n_183__20_;
      r_183__19_ <= r_n_183__19_;
      r_183__18_ <= r_n_183__18_;
      r_183__17_ <= r_n_183__17_;
      r_183__16_ <= r_n_183__16_;
      r_183__15_ <= r_n_183__15_;
      r_183__14_ <= r_n_183__14_;
      r_183__13_ <= r_n_183__13_;
      r_183__12_ <= r_n_183__12_;
      r_183__11_ <= r_n_183__11_;
      r_183__10_ <= r_n_183__10_;
      r_183__9_ <= r_n_183__9_;
      r_183__8_ <= r_n_183__8_;
      r_183__7_ <= r_n_183__7_;
      r_183__6_ <= r_n_183__6_;
      r_183__5_ <= r_n_183__5_;
      r_183__4_ <= r_n_183__4_;
      r_183__3_ <= r_n_183__3_;
      r_183__2_ <= r_n_183__2_;
      r_183__1_ <= r_n_183__1_;
      r_183__0_ <= r_n_183__0_;
    end 
    if(N1976) begin
      r_184__31_ <= r_n_184__31_;
      r_184__30_ <= r_n_184__30_;
      r_184__29_ <= r_n_184__29_;
      r_184__28_ <= r_n_184__28_;
      r_184__27_ <= r_n_184__27_;
      r_184__26_ <= r_n_184__26_;
      r_184__25_ <= r_n_184__25_;
      r_184__24_ <= r_n_184__24_;
      r_184__23_ <= r_n_184__23_;
      r_184__22_ <= r_n_184__22_;
      r_184__21_ <= r_n_184__21_;
      r_184__20_ <= r_n_184__20_;
      r_184__19_ <= r_n_184__19_;
      r_184__18_ <= r_n_184__18_;
      r_184__17_ <= r_n_184__17_;
      r_184__16_ <= r_n_184__16_;
      r_184__15_ <= r_n_184__15_;
      r_184__14_ <= r_n_184__14_;
      r_184__13_ <= r_n_184__13_;
      r_184__12_ <= r_n_184__12_;
      r_184__11_ <= r_n_184__11_;
      r_184__10_ <= r_n_184__10_;
      r_184__9_ <= r_n_184__9_;
      r_184__8_ <= r_n_184__8_;
      r_184__7_ <= r_n_184__7_;
      r_184__6_ <= r_n_184__6_;
      r_184__5_ <= r_n_184__5_;
      r_184__4_ <= r_n_184__4_;
      r_184__3_ <= r_n_184__3_;
      r_184__2_ <= r_n_184__2_;
      r_184__1_ <= r_n_184__1_;
      r_184__0_ <= r_n_184__0_;
    end 
    if(N1977) begin
      r_185__31_ <= r_n_185__31_;
      r_185__30_ <= r_n_185__30_;
      r_185__29_ <= r_n_185__29_;
      r_185__28_ <= r_n_185__28_;
      r_185__27_ <= r_n_185__27_;
      r_185__26_ <= r_n_185__26_;
      r_185__25_ <= r_n_185__25_;
      r_185__24_ <= r_n_185__24_;
      r_185__23_ <= r_n_185__23_;
      r_185__22_ <= r_n_185__22_;
      r_185__21_ <= r_n_185__21_;
      r_185__20_ <= r_n_185__20_;
      r_185__19_ <= r_n_185__19_;
      r_185__18_ <= r_n_185__18_;
      r_185__17_ <= r_n_185__17_;
      r_185__16_ <= r_n_185__16_;
      r_185__15_ <= r_n_185__15_;
      r_185__14_ <= r_n_185__14_;
      r_185__13_ <= r_n_185__13_;
      r_185__12_ <= r_n_185__12_;
      r_185__11_ <= r_n_185__11_;
      r_185__10_ <= r_n_185__10_;
      r_185__9_ <= r_n_185__9_;
      r_185__8_ <= r_n_185__8_;
      r_185__7_ <= r_n_185__7_;
      r_185__6_ <= r_n_185__6_;
      r_185__5_ <= r_n_185__5_;
      r_185__4_ <= r_n_185__4_;
      r_185__3_ <= r_n_185__3_;
      r_185__2_ <= r_n_185__2_;
      r_185__1_ <= r_n_185__1_;
      r_185__0_ <= r_n_185__0_;
    end 
    if(N1978) begin
      r_186__31_ <= r_n_186__31_;
      r_186__30_ <= r_n_186__30_;
      r_186__29_ <= r_n_186__29_;
      r_186__28_ <= r_n_186__28_;
      r_186__27_ <= r_n_186__27_;
      r_186__26_ <= r_n_186__26_;
      r_186__25_ <= r_n_186__25_;
      r_186__24_ <= r_n_186__24_;
      r_186__23_ <= r_n_186__23_;
      r_186__22_ <= r_n_186__22_;
      r_186__21_ <= r_n_186__21_;
      r_186__20_ <= r_n_186__20_;
      r_186__19_ <= r_n_186__19_;
      r_186__18_ <= r_n_186__18_;
      r_186__17_ <= r_n_186__17_;
      r_186__16_ <= r_n_186__16_;
      r_186__15_ <= r_n_186__15_;
      r_186__14_ <= r_n_186__14_;
      r_186__13_ <= r_n_186__13_;
      r_186__12_ <= r_n_186__12_;
      r_186__11_ <= r_n_186__11_;
      r_186__10_ <= r_n_186__10_;
      r_186__9_ <= r_n_186__9_;
      r_186__8_ <= r_n_186__8_;
      r_186__7_ <= r_n_186__7_;
      r_186__6_ <= r_n_186__6_;
      r_186__5_ <= r_n_186__5_;
      r_186__4_ <= r_n_186__4_;
      r_186__3_ <= r_n_186__3_;
      r_186__2_ <= r_n_186__2_;
      r_186__1_ <= r_n_186__1_;
      r_186__0_ <= r_n_186__0_;
    end 
    if(N1979) begin
      r_187__31_ <= r_n_187__31_;
      r_187__30_ <= r_n_187__30_;
      r_187__29_ <= r_n_187__29_;
      r_187__28_ <= r_n_187__28_;
      r_187__27_ <= r_n_187__27_;
      r_187__26_ <= r_n_187__26_;
      r_187__25_ <= r_n_187__25_;
      r_187__24_ <= r_n_187__24_;
      r_187__23_ <= r_n_187__23_;
      r_187__22_ <= r_n_187__22_;
      r_187__21_ <= r_n_187__21_;
      r_187__20_ <= r_n_187__20_;
      r_187__19_ <= r_n_187__19_;
      r_187__18_ <= r_n_187__18_;
      r_187__17_ <= r_n_187__17_;
      r_187__16_ <= r_n_187__16_;
      r_187__15_ <= r_n_187__15_;
      r_187__14_ <= r_n_187__14_;
      r_187__13_ <= r_n_187__13_;
      r_187__12_ <= r_n_187__12_;
      r_187__11_ <= r_n_187__11_;
      r_187__10_ <= r_n_187__10_;
      r_187__9_ <= r_n_187__9_;
      r_187__8_ <= r_n_187__8_;
      r_187__7_ <= r_n_187__7_;
      r_187__6_ <= r_n_187__6_;
      r_187__5_ <= r_n_187__5_;
      r_187__4_ <= r_n_187__4_;
      r_187__3_ <= r_n_187__3_;
      r_187__2_ <= r_n_187__2_;
      r_187__1_ <= r_n_187__1_;
      r_187__0_ <= r_n_187__0_;
    end 
    if(N1980) begin
      r_188__31_ <= r_n_188__31_;
      r_188__30_ <= r_n_188__30_;
      r_188__29_ <= r_n_188__29_;
      r_188__28_ <= r_n_188__28_;
      r_188__27_ <= r_n_188__27_;
      r_188__26_ <= r_n_188__26_;
      r_188__25_ <= r_n_188__25_;
      r_188__24_ <= r_n_188__24_;
      r_188__23_ <= r_n_188__23_;
      r_188__22_ <= r_n_188__22_;
      r_188__21_ <= r_n_188__21_;
      r_188__20_ <= r_n_188__20_;
      r_188__19_ <= r_n_188__19_;
      r_188__18_ <= r_n_188__18_;
      r_188__17_ <= r_n_188__17_;
      r_188__16_ <= r_n_188__16_;
      r_188__15_ <= r_n_188__15_;
      r_188__14_ <= r_n_188__14_;
      r_188__13_ <= r_n_188__13_;
      r_188__12_ <= r_n_188__12_;
      r_188__11_ <= r_n_188__11_;
      r_188__10_ <= r_n_188__10_;
      r_188__9_ <= r_n_188__9_;
      r_188__8_ <= r_n_188__8_;
      r_188__7_ <= r_n_188__7_;
      r_188__6_ <= r_n_188__6_;
      r_188__5_ <= r_n_188__5_;
      r_188__4_ <= r_n_188__4_;
      r_188__3_ <= r_n_188__3_;
      r_188__2_ <= r_n_188__2_;
      r_188__1_ <= r_n_188__1_;
      r_188__0_ <= r_n_188__0_;
    end 
    if(N1981) begin
      r_189__31_ <= r_n_189__31_;
      r_189__30_ <= r_n_189__30_;
      r_189__29_ <= r_n_189__29_;
      r_189__28_ <= r_n_189__28_;
      r_189__27_ <= r_n_189__27_;
      r_189__26_ <= r_n_189__26_;
      r_189__25_ <= r_n_189__25_;
      r_189__24_ <= r_n_189__24_;
      r_189__23_ <= r_n_189__23_;
      r_189__22_ <= r_n_189__22_;
      r_189__21_ <= r_n_189__21_;
      r_189__20_ <= r_n_189__20_;
      r_189__19_ <= r_n_189__19_;
      r_189__18_ <= r_n_189__18_;
      r_189__17_ <= r_n_189__17_;
      r_189__16_ <= r_n_189__16_;
      r_189__15_ <= r_n_189__15_;
      r_189__14_ <= r_n_189__14_;
      r_189__13_ <= r_n_189__13_;
      r_189__12_ <= r_n_189__12_;
      r_189__11_ <= r_n_189__11_;
      r_189__10_ <= r_n_189__10_;
      r_189__9_ <= r_n_189__9_;
      r_189__8_ <= r_n_189__8_;
      r_189__7_ <= r_n_189__7_;
      r_189__6_ <= r_n_189__6_;
      r_189__5_ <= r_n_189__5_;
      r_189__4_ <= r_n_189__4_;
      r_189__3_ <= r_n_189__3_;
      r_189__2_ <= r_n_189__2_;
      r_189__1_ <= r_n_189__1_;
      r_189__0_ <= r_n_189__0_;
    end 
    if(N1982) begin
      r_190__31_ <= r_n_190__31_;
      r_190__30_ <= r_n_190__30_;
      r_190__29_ <= r_n_190__29_;
      r_190__28_ <= r_n_190__28_;
      r_190__27_ <= r_n_190__27_;
      r_190__26_ <= r_n_190__26_;
      r_190__25_ <= r_n_190__25_;
      r_190__24_ <= r_n_190__24_;
      r_190__23_ <= r_n_190__23_;
      r_190__22_ <= r_n_190__22_;
      r_190__21_ <= r_n_190__21_;
      r_190__20_ <= r_n_190__20_;
      r_190__19_ <= r_n_190__19_;
      r_190__18_ <= r_n_190__18_;
      r_190__17_ <= r_n_190__17_;
      r_190__16_ <= r_n_190__16_;
      r_190__15_ <= r_n_190__15_;
      r_190__14_ <= r_n_190__14_;
      r_190__13_ <= r_n_190__13_;
      r_190__12_ <= r_n_190__12_;
      r_190__11_ <= r_n_190__11_;
      r_190__10_ <= r_n_190__10_;
      r_190__9_ <= r_n_190__9_;
      r_190__8_ <= r_n_190__8_;
      r_190__7_ <= r_n_190__7_;
      r_190__6_ <= r_n_190__6_;
      r_190__5_ <= r_n_190__5_;
      r_190__4_ <= r_n_190__4_;
      r_190__3_ <= r_n_190__3_;
      r_190__2_ <= r_n_190__2_;
      r_190__1_ <= r_n_190__1_;
      r_190__0_ <= r_n_190__0_;
    end 
    if(N1983) begin
      r_191__31_ <= r_n_191__31_;
      r_191__30_ <= r_n_191__30_;
      r_191__29_ <= r_n_191__29_;
      r_191__28_ <= r_n_191__28_;
      r_191__27_ <= r_n_191__27_;
      r_191__26_ <= r_n_191__26_;
      r_191__25_ <= r_n_191__25_;
      r_191__24_ <= r_n_191__24_;
      r_191__23_ <= r_n_191__23_;
      r_191__22_ <= r_n_191__22_;
      r_191__21_ <= r_n_191__21_;
      r_191__20_ <= r_n_191__20_;
      r_191__19_ <= r_n_191__19_;
      r_191__18_ <= r_n_191__18_;
      r_191__17_ <= r_n_191__17_;
      r_191__16_ <= r_n_191__16_;
      r_191__15_ <= r_n_191__15_;
      r_191__14_ <= r_n_191__14_;
      r_191__13_ <= r_n_191__13_;
      r_191__12_ <= r_n_191__12_;
      r_191__11_ <= r_n_191__11_;
      r_191__10_ <= r_n_191__10_;
      r_191__9_ <= r_n_191__9_;
      r_191__8_ <= r_n_191__8_;
      r_191__7_ <= r_n_191__7_;
      r_191__6_ <= r_n_191__6_;
      r_191__5_ <= r_n_191__5_;
      r_191__4_ <= r_n_191__4_;
      r_191__3_ <= r_n_191__3_;
      r_191__2_ <= r_n_191__2_;
      r_191__1_ <= r_n_191__1_;
      r_191__0_ <= r_n_191__0_;
    end 
    if(N1984) begin
      r_192__31_ <= r_n_192__31_;
      r_192__30_ <= r_n_192__30_;
      r_192__29_ <= r_n_192__29_;
      r_192__28_ <= r_n_192__28_;
      r_192__27_ <= r_n_192__27_;
      r_192__26_ <= r_n_192__26_;
      r_192__25_ <= r_n_192__25_;
      r_192__24_ <= r_n_192__24_;
      r_192__23_ <= r_n_192__23_;
      r_192__22_ <= r_n_192__22_;
      r_192__21_ <= r_n_192__21_;
      r_192__20_ <= r_n_192__20_;
      r_192__19_ <= r_n_192__19_;
      r_192__18_ <= r_n_192__18_;
      r_192__17_ <= r_n_192__17_;
      r_192__16_ <= r_n_192__16_;
      r_192__15_ <= r_n_192__15_;
      r_192__14_ <= r_n_192__14_;
      r_192__13_ <= r_n_192__13_;
      r_192__12_ <= r_n_192__12_;
      r_192__11_ <= r_n_192__11_;
      r_192__10_ <= r_n_192__10_;
      r_192__9_ <= r_n_192__9_;
      r_192__8_ <= r_n_192__8_;
      r_192__7_ <= r_n_192__7_;
      r_192__6_ <= r_n_192__6_;
      r_192__5_ <= r_n_192__5_;
      r_192__4_ <= r_n_192__4_;
      r_192__3_ <= r_n_192__3_;
      r_192__2_ <= r_n_192__2_;
      r_192__1_ <= r_n_192__1_;
      r_192__0_ <= r_n_192__0_;
    end 
    if(N1985) begin
      r_193__31_ <= r_n_193__31_;
      r_193__30_ <= r_n_193__30_;
      r_193__29_ <= r_n_193__29_;
      r_193__28_ <= r_n_193__28_;
      r_193__27_ <= r_n_193__27_;
      r_193__26_ <= r_n_193__26_;
      r_193__25_ <= r_n_193__25_;
      r_193__24_ <= r_n_193__24_;
      r_193__23_ <= r_n_193__23_;
      r_193__22_ <= r_n_193__22_;
      r_193__21_ <= r_n_193__21_;
      r_193__20_ <= r_n_193__20_;
      r_193__19_ <= r_n_193__19_;
      r_193__18_ <= r_n_193__18_;
      r_193__17_ <= r_n_193__17_;
      r_193__16_ <= r_n_193__16_;
      r_193__15_ <= r_n_193__15_;
      r_193__14_ <= r_n_193__14_;
      r_193__13_ <= r_n_193__13_;
      r_193__12_ <= r_n_193__12_;
      r_193__11_ <= r_n_193__11_;
      r_193__10_ <= r_n_193__10_;
      r_193__9_ <= r_n_193__9_;
      r_193__8_ <= r_n_193__8_;
      r_193__7_ <= r_n_193__7_;
      r_193__6_ <= r_n_193__6_;
      r_193__5_ <= r_n_193__5_;
      r_193__4_ <= r_n_193__4_;
      r_193__3_ <= r_n_193__3_;
      r_193__2_ <= r_n_193__2_;
      r_193__1_ <= r_n_193__1_;
      r_193__0_ <= r_n_193__0_;
    end 
    if(N1986) begin
      r_194__31_ <= r_n_194__31_;
      r_194__30_ <= r_n_194__30_;
      r_194__29_ <= r_n_194__29_;
      r_194__28_ <= r_n_194__28_;
      r_194__27_ <= r_n_194__27_;
      r_194__26_ <= r_n_194__26_;
      r_194__25_ <= r_n_194__25_;
      r_194__24_ <= r_n_194__24_;
      r_194__23_ <= r_n_194__23_;
      r_194__22_ <= r_n_194__22_;
      r_194__21_ <= r_n_194__21_;
      r_194__20_ <= r_n_194__20_;
      r_194__19_ <= r_n_194__19_;
      r_194__18_ <= r_n_194__18_;
      r_194__17_ <= r_n_194__17_;
      r_194__16_ <= r_n_194__16_;
      r_194__15_ <= r_n_194__15_;
      r_194__14_ <= r_n_194__14_;
      r_194__13_ <= r_n_194__13_;
      r_194__12_ <= r_n_194__12_;
      r_194__11_ <= r_n_194__11_;
      r_194__10_ <= r_n_194__10_;
      r_194__9_ <= r_n_194__9_;
      r_194__8_ <= r_n_194__8_;
      r_194__7_ <= r_n_194__7_;
      r_194__6_ <= r_n_194__6_;
      r_194__5_ <= r_n_194__5_;
      r_194__4_ <= r_n_194__4_;
      r_194__3_ <= r_n_194__3_;
      r_194__2_ <= r_n_194__2_;
      r_194__1_ <= r_n_194__1_;
      r_194__0_ <= r_n_194__0_;
    end 
    if(N1987) begin
      r_195__31_ <= r_n_195__31_;
      r_195__30_ <= r_n_195__30_;
      r_195__29_ <= r_n_195__29_;
      r_195__28_ <= r_n_195__28_;
      r_195__27_ <= r_n_195__27_;
      r_195__26_ <= r_n_195__26_;
      r_195__25_ <= r_n_195__25_;
      r_195__24_ <= r_n_195__24_;
      r_195__23_ <= r_n_195__23_;
      r_195__22_ <= r_n_195__22_;
      r_195__21_ <= r_n_195__21_;
      r_195__20_ <= r_n_195__20_;
      r_195__19_ <= r_n_195__19_;
      r_195__18_ <= r_n_195__18_;
      r_195__17_ <= r_n_195__17_;
      r_195__16_ <= r_n_195__16_;
      r_195__15_ <= r_n_195__15_;
      r_195__14_ <= r_n_195__14_;
      r_195__13_ <= r_n_195__13_;
      r_195__12_ <= r_n_195__12_;
      r_195__11_ <= r_n_195__11_;
      r_195__10_ <= r_n_195__10_;
      r_195__9_ <= r_n_195__9_;
      r_195__8_ <= r_n_195__8_;
      r_195__7_ <= r_n_195__7_;
      r_195__6_ <= r_n_195__6_;
      r_195__5_ <= r_n_195__5_;
      r_195__4_ <= r_n_195__4_;
      r_195__3_ <= r_n_195__3_;
      r_195__2_ <= r_n_195__2_;
      r_195__1_ <= r_n_195__1_;
      r_195__0_ <= r_n_195__0_;
    end 
    if(N1988) begin
      r_196__31_ <= r_n_196__31_;
      r_196__30_ <= r_n_196__30_;
      r_196__29_ <= r_n_196__29_;
      r_196__28_ <= r_n_196__28_;
      r_196__27_ <= r_n_196__27_;
      r_196__26_ <= r_n_196__26_;
      r_196__25_ <= r_n_196__25_;
      r_196__24_ <= r_n_196__24_;
      r_196__23_ <= r_n_196__23_;
      r_196__22_ <= r_n_196__22_;
      r_196__21_ <= r_n_196__21_;
      r_196__20_ <= r_n_196__20_;
      r_196__19_ <= r_n_196__19_;
      r_196__18_ <= r_n_196__18_;
      r_196__17_ <= r_n_196__17_;
      r_196__16_ <= r_n_196__16_;
      r_196__15_ <= r_n_196__15_;
      r_196__14_ <= r_n_196__14_;
      r_196__13_ <= r_n_196__13_;
      r_196__12_ <= r_n_196__12_;
      r_196__11_ <= r_n_196__11_;
      r_196__10_ <= r_n_196__10_;
      r_196__9_ <= r_n_196__9_;
      r_196__8_ <= r_n_196__8_;
      r_196__7_ <= r_n_196__7_;
      r_196__6_ <= r_n_196__6_;
      r_196__5_ <= r_n_196__5_;
      r_196__4_ <= r_n_196__4_;
      r_196__3_ <= r_n_196__3_;
      r_196__2_ <= r_n_196__2_;
      r_196__1_ <= r_n_196__1_;
      r_196__0_ <= r_n_196__0_;
    end 
    if(N1989) begin
      r_197__31_ <= r_n_197__31_;
      r_197__30_ <= r_n_197__30_;
      r_197__29_ <= r_n_197__29_;
      r_197__28_ <= r_n_197__28_;
      r_197__27_ <= r_n_197__27_;
      r_197__26_ <= r_n_197__26_;
      r_197__25_ <= r_n_197__25_;
      r_197__24_ <= r_n_197__24_;
      r_197__23_ <= r_n_197__23_;
      r_197__22_ <= r_n_197__22_;
      r_197__21_ <= r_n_197__21_;
      r_197__20_ <= r_n_197__20_;
      r_197__19_ <= r_n_197__19_;
      r_197__18_ <= r_n_197__18_;
      r_197__17_ <= r_n_197__17_;
      r_197__16_ <= r_n_197__16_;
      r_197__15_ <= r_n_197__15_;
      r_197__14_ <= r_n_197__14_;
      r_197__13_ <= r_n_197__13_;
      r_197__12_ <= r_n_197__12_;
      r_197__11_ <= r_n_197__11_;
      r_197__10_ <= r_n_197__10_;
      r_197__9_ <= r_n_197__9_;
      r_197__8_ <= r_n_197__8_;
      r_197__7_ <= r_n_197__7_;
      r_197__6_ <= r_n_197__6_;
      r_197__5_ <= r_n_197__5_;
      r_197__4_ <= r_n_197__4_;
      r_197__3_ <= r_n_197__3_;
      r_197__2_ <= r_n_197__2_;
      r_197__1_ <= r_n_197__1_;
      r_197__0_ <= r_n_197__0_;
    end 
    if(N1990) begin
      r_198__31_ <= r_n_198__31_;
      r_198__30_ <= r_n_198__30_;
      r_198__29_ <= r_n_198__29_;
      r_198__28_ <= r_n_198__28_;
      r_198__27_ <= r_n_198__27_;
      r_198__26_ <= r_n_198__26_;
      r_198__25_ <= r_n_198__25_;
      r_198__24_ <= r_n_198__24_;
      r_198__23_ <= r_n_198__23_;
      r_198__22_ <= r_n_198__22_;
      r_198__21_ <= r_n_198__21_;
      r_198__20_ <= r_n_198__20_;
      r_198__19_ <= r_n_198__19_;
      r_198__18_ <= r_n_198__18_;
      r_198__17_ <= r_n_198__17_;
      r_198__16_ <= r_n_198__16_;
      r_198__15_ <= r_n_198__15_;
      r_198__14_ <= r_n_198__14_;
      r_198__13_ <= r_n_198__13_;
      r_198__12_ <= r_n_198__12_;
      r_198__11_ <= r_n_198__11_;
      r_198__10_ <= r_n_198__10_;
      r_198__9_ <= r_n_198__9_;
      r_198__8_ <= r_n_198__8_;
      r_198__7_ <= r_n_198__7_;
      r_198__6_ <= r_n_198__6_;
      r_198__5_ <= r_n_198__5_;
      r_198__4_ <= r_n_198__4_;
      r_198__3_ <= r_n_198__3_;
      r_198__2_ <= r_n_198__2_;
      r_198__1_ <= r_n_198__1_;
      r_198__0_ <= r_n_198__0_;
    end 
    if(N1991) begin
      r_199__31_ <= r_n_199__31_;
      r_199__30_ <= r_n_199__30_;
      r_199__29_ <= r_n_199__29_;
      r_199__28_ <= r_n_199__28_;
      r_199__27_ <= r_n_199__27_;
      r_199__26_ <= r_n_199__26_;
      r_199__25_ <= r_n_199__25_;
      r_199__24_ <= r_n_199__24_;
      r_199__23_ <= r_n_199__23_;
      r_199__22_ <= r_n_199__22_;
      r_199__21_ <= r_n_199__21_;
      r_199__20_ <= r_n_199__20_;
      r_199__19_ <= r_n_199__19_;
      r_199__18_ <= r_n_199__18_;
      r_199__17_ <= r_n_199__17_;
      r_199__16_ <= r_n_199__16_;
      r_199__15_ <= r_n_199__15_;
      r_199__14_ <= r_n_199__14_;
      r_199__13_ <= r_n_199__13_;
      r_199__12_ <= r_n_199__12_;
      r_199__11_ <= r_n_199__11_;
      r_199__10_ <= r_n_199__10_;
      r_199__9_ <= r_n_199__9_;
      r_199__8_ <= r_n_199__8_;
      r_199__7_ <= r_n_199__7_;
      r_199__6_ <= r_n_199__6_;
      r_199__5_ <= r_n_199__5_;
      r_199__4_ <= r_n_199__4_;
      r_199__3_ <= r_n_199__3_;
      r_199__2_ <= r_n_199__2_;
      r_199__1_ <= r_n_199__1_;
      r_199__0_ <= r_n_199__0_;
    end 
    if(N1992) begin
      r_200__31_ <= r_n_200__31_;
      r_200__30_ <= r_n_200__30_;
      r_200__29_ <= r_n_200__29_;
      r_200__28_ <= r_n_200__28_;
      r_200__27_ <= r_n_200__27_;
      r_200__26_ <= r_n_200__26_;
      r_200__25_ <= r_n_200__25_;
      r_200__24_ <= r_n_200__24_;
      r_200__23_ <= r_n_200__23_;
      r_200__22_ <= r_n_200__22_;
      r_200__21_ <= r_n_200__21_;
      r_200__20_ <= r_n_200__20_;
      r_200__19_ <= r_n_200__19_;
      r_200__18_ <= r_n_200__18_;
      r_200__17_ <= r_n_200__17_;
      r_200__16_ <= r_n_200__16_;
      r_200__15_ <= r_n_200__15_;
      r_200__14_ <= r_n_200__14_;
      r_200__13_ <= r_n_200__13_;
      r_200__12_ <= r_n_200__12_;
      r_200__11_ <= r_n_200__11_;
      r_200__10_ <= r_n_200__10_;
      r_200__9_ <= r_n_200__9_;
      r_200__8_ <= r_n_200__8_;
      r_200__7_ <= r_n_200__7_;
      r_200__6_ <= r_n_200__6_;
      r_200__5_ <= r_n_200__5_;
      r_200__4_ <= r_n_200__4_;
      r_200__3_ <= r_n_200__3_;
      r_200__2_ <= r_n_200__2_;
      r_200__1_ <= r_n_200__1_;
      r_200__0_ <= r_n_200__0_;
    end 
    if(N1993) begin
      r_201__31_ <= r_n_201__31_;
      r_201__30_ <= r_n_201__30_;
      r_201__29_ <= r_n_201__29_;
      r_201__28_ <= r_n_201__28_;
      r_201__27_ <= r_n_201__27_;
      r_201__26_ <= r_n_201__26_;
      r_201__25_ <= r_n_201__25_;
      r_201__24_ <= r_n_201__24_;
      r_201__23_ <= r_n_201__23_;
      r_201__22_ <= r_n_201__22_;
      r_201__21_ <= r_n_201__21_;
      r_201__20_ <= r_n_201__20_;
      r_201__19_ <= r_n_201__19_;
      r_201__18_ <= r_n_201__18_;
      r_201__17_ <= r_n_201__17_;
      r_201__16_ <= r_n_201__16_;
      r_201__15_ <= r_n_201__15_;
      r_201__14_ <= r_n_201__14_;
      r_201__13_ <= r_n_201__13_;
      r_201__12_ <= r_n_201__12_;
      r_201__11_ <= r_n_201__11_;
      r_201__10_ <= r_n_201__10_;
      r_201__9_ <= r_n_201__9_;
      r_201__8_ <= r_n_201__8_;
      r_201__7_ <= r_n_201__7_;
      r_201__6_ <= r_n_201__6_;
      r_201__5_ <= r_n_201__5_;
      r_201__4_ <= r_n_201__4_;
      r_201__3_ <= r_n_201__3_;
      r_201__2_ <= r_n_201__2_;
      r_201__1_ <= r_n_201__1_;
      r_201__0_ <= r_n_201__0_;
    end 
    if(N1994) begin
      r_202__31_ <= r_n_202__31_;
      r_202__30_ <= r_n_202__30_;
      r_202__29_ <= r_n_202__29_;
      r_202__28_ <= r_n_202__28_;
      r_202__27_ <= r_n_202__27_;
      r_202__26_ <= r_n_202__26_;
      r_202__25_ <= r_n_202__25_;
      r_202__24_ <= r_n_202__24_;
      r_202__23_ <= r_n_202__23_;
      r_202__22_ <= r_n_202__22_;
      r_202__21_ <= r_n_202__21_;
      r_202__20_ <= r_n_202__20_;
      r_202__19_ <= r_n_202__19_;
      r_202__18_ <= r_n_202__18_;
      r_202__17_ <= r_n_202__17_;
      r_202__16_ <= r_n_202__16_;
      r_202__15_ <= r_n_202__15_;
      r_202__14_ <= r_n_202__14_;
      r_202__13_ <= r_n_202__13_;
      r_202__12_ <= r_n_202__12_;
      r_202__11_ <= r_n_202__11_;
      r_202__10_ <= r_n_202__10_;
      r_202__9_ <= r_n_202__9_;
      r_202__8_ <= r_n_202__8_;
      r_202__7_ <= r_n_202__7_;
      r_202__6_ <= r_n_202__6_;
      r_202__5_ <= r_n_202__5_;
      r_202__4_ <= r_n_202__4_;
      r_202__3_ <= r_n_202__3_;
      r_202__2_ <= r_n_202__2_;
      r_202__1_ <= r_n_202__1_;
      r_202__0_ <= r_n_202__0_;
    end 
    if(N1995) begin
      r_203__31_ <= r_n_203__31_;
      r_203__30_ <= r_n_203__30_;
      r_203__29_ <= r_n_203__29_;
      r_203__28_ <= r_n_203__28_;
      r_203__27_ <= r_n_203__27_;
      r_203__26_ <= r_n_203__26_;
      r_203__25_ <= r_n_203__25_;
      r_203__24_ <= r_n_203__24_;
      r_203__23_ <= r_n_203__23_;
      r_203__22_ <= r_n_203__22_;
      r_203__21_ <= r_n_203__21_;
      r_203__20_ <= r_n_203__20_;
      r_203__19_ <= r_n_203__19_;
      r_203__18_ <= r_n_203__18_;
      r_203__17_ <= r_n_203__17_;
      r_203__16_ <= r_n_203__16_;
      r_203__15_ <= r_n_203__15_;
      r_203__14_ <= r_n_203__14_;
      r_203__13_ <= r_n_203__13_;
      r_203__12_ <= r_n_203__12_;
      r_203__11_ <= r_n_203__11_;
      r_203__10_ <= r_n_203__10_;
      r_203__9_ <= r_n_203__9_;
      r_203__8_ <= r_n_203__8_;
      r_203__7_ <= r_n_203__7_;
      r_203__6_ <= r_n_203__6_;
      r_203__5_ <= r_n_203__5_;
      r_203__4_ <= r_n_203__4_;
      r_203__3_ <= r_n_203__3_;
      r_203__2_ <= r_n_203__2_;
      r_203__1_ <= r_n_203__1_;
      r_203__0_ <= r_n_203__0_;
    end 
    if(N1996) begin
      r_204__31_ <= r_n_204__31_;
      r_204__30_ <= r_n_204__30_;
      r_204__29_ <= r_n_204__29_;
      r_204__28_ <= r_n_204__28_;
      r_204__27_ <= r_n_204__27_;
      r_204__26_ <= r_n_204__26_;
      r_204__25_ <= r_n_204__25_;
      r_204__24_ <= r_n_204__24_;
      r_204__23_ <= r_n_204__23_;
      r_204__22_ <= r_n_204__22_;
      r_204__21_ <= r_n_204__21_;
      r_204__20_ <= r_n_204__20_;
      r_204__19_ <= r_n_204__19_;
      r_204__18_ <= r_n_204__18_;
      r_204__17_ <= r_n_204__17_;
      r_204__16_ <= r_n_204__16_;
      r_204__15_ <= r_n_204__15_;
      r_204__14_ <= r_n_204__14_;
      r_204__13_ <= r_n_204__13_;
      r_204__12_ <= r_n_204__12_;
      r_204__11_ <= r_n_204__11_;
      r_204__10_ <= r_n_204__10_;
      r_204__9_ <= r_n_204__9_;
      r_204__8_ <= r_n_204__8_;
      r_204__7_ <= r_n_204__7_;
      r_204__6_ <= r_n_204__6_;
      r_204__5_ <= r_n_204__5_;
      r_204__4_ <= r_n_204__4_;
      r_204__3_ <= r_n_204__3_;
      r_204__2_ <= r_n_204__2_;
      r_204__1_ <= r_n_204__1_;
      r_204__0_ <= r_n_204__0_;
    end 
    if(N1997) begin
      r_205__31_ <= r_n_205__31_;
      r_205__30_ <= r_n_205__30_;
      r_205__29_ <= r_n_205__29_;
      r_205__28_ <= r_n_205__28_;
      r_205__27_ <= r_n_205__27_;
      r_205__26_ <= r_n_205__26_;
      r_205__25_ <= r_n_205__25_;
      r_205__24_ <= r_n_205__24_;
      r_205__23_ <= r_n_205__23_;
      r_205__22_ <= r_n_205__22_;
      r_205__21_ <= r_n_205__21_;
      r_205__20_ <= r_n_205__20_;
      r_205__19_ <= r_n_205__19_;
      r_205__18_ <= r_n_205__18_;
      r_205__17_ <= r_n_205__17_;
      r_205__16_ <= r_n_205__16_;
      r_205__15_ <= r_n_205__15_;
      r_205__14_ <= r_n_205__14_;
      r_205__13_ <= r_n_205__13_;
      r_205__12_ <= r_n_205__12_;
      r_205__11_ <= r_n_205__11_;
      r_205__10_ <= r_n_205__10_;
      r_205__9_ <= r_n_205__9_;
      r_205__8_ <= r_n_205__8_;
      r_205__7_ <= r_n_205__7_;
      r_205__6_ <= r_n_205__6_;
      r_205__5_ <= r_n_205__5_;
      r_205__4_ <= r_n_205__4_;
      r_205__3_ <= r_n_205__3_;
      r_205__2_ <= r_n_205__2_;
      r_205__1_ <= r_n_205__1_;
      r_205__0_ <= r_n_205__0_;
    end 
    if(N1998) begin
      r_206__31_ <= r_n_206__31_;
      r_206__30_ <= r_n_206__30_;
      r_206__29_ <= r_n_206__29_;
      r_206__28_ <= r_n_206__28_;
      r_206__27_ <= r_n_206__27_;
      r_206__26_ <= r_n_206__26_;
      r_206__25_ <= r_n_206__25_;
      r_206__24_ <= r_n_206__24_;
      r_206__23_ <= r_n_206__23_;
      r_206__22_ <= r_n_206__22_;
      r_206__21_ <= r_n_206__21_;
      r_206__20_ <= r_n_206__20_;
      r_206__19_ <= r_n_206__19_;
      r_206__18_ <= r_n_206__18_;
      r_206__17_ <= r_n_206__17_;
      r_206__16_ <= r_n_206__16_;
      r_206__15_ <= r_n_206__15_;
      r_206__14_ <= r_n_206__14_;
      r_206__13_ <= r_n_206__13_;
      r_206__12_ <= r_n_206__12_;
      r_206__11_ <= r_n_206__11_;
      r_206__10_ <= r_n_206__10_;
      r_206__9_ <= r_n_206__9_;
      r_206__8_ <= r_n_206__8_;
      r_206__7_ <= r_n_206__7_;
      r_206__6_ <= r_n_206__6_;
      r_206__5_ <= r_n_206__5_;
      r_206__4_ <= r_n_206__4_;
      r_206__3_ <= r_n_206__3_;
      r_206__2_ <= r_n_206__2_;
      r_206__1_ <= r_n_206__1_;
      r_206__0_ <= r_n_206__0_;
    end 
    if(N1999) begin
      r_207__31_ <= r_n_207__31_;
      r_207__30_ <= r_n_207__30_;
      r_207__29_ <= r_n_207__29_;
      r_207__28_ <= r_n_207__28_;
      r_207__27_ <= r_n_207__27_;
      r_207__26_ <= r_n_207__26_;
      r_207__25_ <= r_n_207__25_;
      r_207__24_ <= r_n_207__24_;
      r_207__23_ <= r_n_207__23_;
      r_207__22_ <= r_n_207__22_;
      r_207__21_ <= r_n_207__21_;
      r_207__20_ <= r_n_207__20_;
      r_207__19_ <= r_n_207__19_;
      r_207__18_ <= r_n_207__18_;
      r_207__17_ <= r_n_207__17_;
      r_207__16_ <= r_n_207__16_;
      r_207__15_ <= r_n_207__15_;
      r_207__14_ <= r_n_207__14_;
      r_207__13_ <= r_n_207__13_;
      r_207__12_ <= r_n_207__12_;
      r_207__11_ <= r_n_207__11_;
      r_207__10_ <= r_n_207__10_;
      r_207__9_ <= r_n_207__9_;
      r_207__8_ <= r_n_207__8_;
      r_207__7_ <= r_n_207__7_;
      r_207__6_ <= r_n_207__6_;
      r_207__5_ <= r_n_207__5_;
      r_207__4_ <= r_n_207__4_;
      r_207__3_ <= r_n_207__3_;
      r_207__2_ <= r_n_207__2_;
      r_207__1_ <= r_n_207__1_;
      r_207__0_ <= r_n_207__0_;
    end 
    if(N2000) begin
      r_208__31_ <= r_n_208__31_;
      r_208__30_ <= r_n_208__30_;
      r_208__29_ <= r_n_208__29_;
      r_208__28_ <= r_n_208__28_;
      r_208__27_ <= r_n_208__27_;
      r_208__26_ <= r_n_208__26_;
      r_208__25_ <= r_n_208__25_;
      r_208__24_ <= r_n_208__24_;
      r_208__23_ <= r_n_208__23_;
      r_208__22_ <= r_n_208__22_;
      r_208__21_ <= r_n_208__21_;
      r_208__20_ <= r_n_208__20_;
      r_208__19_ <= r_n_208__19_;
      r_208__18_ <= r_n_208__18_;
      r_208__17_ <= r_n_208__17_;
      r_208__16_ <= r_n_208__16_;
      r_208__15_ <= r_n_208__15_;
      r_208__14_ <= r_n_208__14_;
      r_208__13_ <= r_n_208__13_;
      r_208__12_ <= r_n_208__12_;
      r_208__11_ <= r_n_208__11_;
      r_208__10_ <= r_n_208__10_;
      r_208__9_ <= r_n_208__9_;
      r_208__8_ <= r_n_208__8_;
      r_208__7_ <= r_n_208__7_;
      r_208__6_ <= r_n_208__6_;
      r_208__5_ <= r_n_208__5_;
      r_208__4_ <= r_n_208__4_;
      r_208__3_ <= r_n_208__3_;
      r_208__2_ <= r_n_208__2_;
      r_208__1_ <= r_n_208__1_;
      r_208__0_ <= r_n_208__0_;
    end 
    if(N2001) begin
      r_209__31_ <= r_n_209__31_;
      r_209__30_ <= r_n_209__30_;
      r_209__29_ <= r_n_209__29_;
      r_209__28_ <= r_n_209__28_;
      r_209__27_ <= r_n_209__27_;
      r_209__26_ <= r_n_209__26_;
      r_209__25_ <= r_n_209__25_;
      r_209__24_ <= r_n_209__24_;
      r_209__23_ <= r_n_209__23_;
      r_209__22_ <= r_n_209__22_;
      r_209__21_ <= r_n_209__21_;
      r_209__20_ <= r_n_209__20_;
      r_209__19_ <= r_n_209__19_;
      r_209__18_ <= r_n_209__18_;
      r_209__17_ <= r_n_209__17_;
      r_209__16_ <= r_n_209__16_;
      r_209__15_ <= r_n_209__15_;
      r_209__14_ <= r_n_209__14_;
      r_209__13_ <= r_n_209__13_;
      r_209__12_ <= r_n_209__12_;
      r_209__11_ <= r_n_209__11_;
      r_209__10_ <= r_n_209__10_;
      r_209__9_ <= r_n_209__9_;
      r_209__8_ <= r_n_209__8_;
      r_209__7_ <= r_n_209__7_;
      r_209__6_ <= r_n_209__6_;
      r_209__5_ <= r_n_209__5_;
      r_209__4_ <= r_n_209__4_;
      r_209__3_ <= r_n_209__3_;
      r_209__2_ <= r_n_209__2_;
      r_209__1_ <= r_n_209__1_;
      r_209__0_ <= r_n_209__0_;
    end 
    if(N2002) begin
      r_210__31_ <= r_n_210__31_;
      r_210__30_ <= r_n_210__30_;
      r_210__29_ <= r_n_210__29_;
      r_210__28_ <= r_n_210__28_;
      r_210__27_ <= r_n_210__27_;
      r_210__26_ <= r_n_210__26_;
      r_210__25_ <= r_n_210__25_;
      r_210__24_ <= r_n_210__24_;
      r_210__23_ <= r_n_210__23_;
      r_210__22_ <= r_n_210__22_;
      r_210__21_ <= r_n_210__21_;
      r_210__20_ <= r_n_210__20_;
      r_210__19_ <= r_n_210__19_;
      r_210__18_ <= r_n_210__18_;
      r_210__17_ <= r_n_210__17_;
      r_210__16_ <= r_n_210__16_;
      r_210__15_ <= r_n_210__15_;
      r_210__14_ <= r_n_210__14_;
      r_210__13_ <= r_n_210__13_;
      r_210__12_ <= r_n_210__12_;
      r_210__11_ <= r_n_210__11_;
      r_210__10_ <= r_n_210__10_;
      r_210__9_ <= r_n_210__9_;
      r_210__8_ <= r_n_210__8_;
      r_210__7_ <= r_n_210__7_;
      r_210__6_ <= r_n_210__6_;
      r_210__5_ <= r_n_210__5_;
      r_210__4_ <= r_n_210__4_;
      r_210__3_ <= r_n_210__3_;
      r_210__2_ <= r_n_210__2_;
      r_210__1_ <= r_n_210__1_;
      r_210__0_ <= r_n_210__0_;
    end 
    if(N2003) begin
      r_211__31_ <= r_n_211__31_;
      r_211__30_ <= r_n_211__30_;
      r_211__29_ <= r_n_211__29_;
      r_211__28_ <= r_n_211__28_;
      r_211__27_ <= r_n_211__27_;
      r_211__26_ <= r_n_211__26_;
      r_211__25_ <= r_n_211__25_;
      r_211__24_ <= r_n_211__24_;
      r_211__23_ <= r_n_211__23_;
      r_211__22_ <= r_n_211__22_;
      r_211__21_ <= r_n_211__21_;
      r_211__20_ <= r_n_211__20_;
      r_211__19_ <= r_n_211__19_;
      r_211__18_ <= r_n_211__18_;
      r_211__17_ <= r_n_211__17_;
      r_211__16_ <= r_n_211__16_;
      r_211__15_ <= r_n_211__15_;
      r_211__14_ <= r_n_211__14_;
      r_211__13_ <= r_n_211__13_;
      r_211__12_ <= r_n_211__12_;
      r_211__11_ <= r_n_211__11_;
      r_211__10_ <= r_n_211__10_;
      r_211__9_ <= r_n_211__9_;
      r_211__8_ <= r_n_211__8_;
      r_211__7_ <= r_n_211__7_;
      r_211__6_ <= r_n_211__6_;
      r_211__5_ <= r_n_211__5_;
      r_211__4_ <= r_n_211__4_;
      r_211__3_ <= r_n_211__3_;
      r_211__2_ <= r_n_211__2_;
      r_211__1_ <= r_n_211__1_;
      r_211__0_ <= r_n_211__0_;
    end 
    if(N2004) begin
      r_212__31_ <= r_n_212__31_;
      r_212__30_ <= r_n_212__30_;
      r_212__29_ <= r_n_212__29_;
      r_212__28_ <= r_n_212__28_;
      r_212__27_ <= r_n_212__27_;
      r_212__26_ <= r_n_212__26_;
      r_212__25_ <= r_n_212__25_;
      r_212__24_ <= r_n_212__24_;
      r_212__23_ <= r_n_212__23_;
      r_212__22_ <= r_n_212__22_;
      r_212__21_ <= r_n_212__21_;
      r_212__20_ <= r_n_212__20_;
      r_212__19_ <= r_n_212__19_;
      r_212__18_ <= r_n_212__18_;
      r_212__17_ <= r_n_212__17_;
      r_212__16_ <= r_n_212__16_;
      r_212__15_ <= r_n_212__15_;
      r_212__14_ <= r_n_212__14_;
      r_212__13_ <= r_n_212__13_;
      r_212__12_ <= r_n_212__12_;
      r_212__11_ <= r_n_212__11_;
      r_212__10_ <= r_n_212__10_;
      r_212__9_ <= r_n_212__9_;
      r_212__8_ <= r_n_212__8_;
      r_212__7_ <= r_n_212__7_;
      r_212__6_ <= r_n_212__6_;
      r_212__5_ <= r_n_212__5_;
      r_212__4_ <= r_n_212__4_;
      r_212__3_ <= r_n_212__3_;
      r_212__2_ <= r_n_212__2_;
      r_212__1_ <= r_n_212__1_;
      r_212__0_ <= r_n_212__0_;
    end 
    if(N2005) begin
      r_213__31_ <= r_n_213__31_;
      r_213__30_ <= r_n_213__30_;
      r_213__29_ <= r_n_213__29_;
      r_213__28_ <= r_n_213__28_;
      r_213__27_ <= r_n_213__27_;
      r_213__26_ <= r_n_213__26_;
      r_213__25_ <= r_n_213__25_;
      r_213__24_ <= r_n_213__24_;
      r_213__23_ <= r_n_213__23_;
      r_213__22_ <= r_n_213__22_;
      r_213__21_ <= r_n_213__21_;
      r_213__20_ <= r_n_213__20_;
      r_213__19_ <= r_n_213__19_;
      r_213__18_ <= r_n_213__18_;
      r_213__17_ <= r_n_213__17_;
      r_213__16_ <= r_n_213__16_;
      r_213__15_ <= r_n_213__15_;
      r_213__14_ <= r_n_213__14_;
      r_213__13_ <= r_n_213__13_;
      r_213__12_ <= r_n_213__12_;
      r_213__11_ <= r_n_213__11_;
      r_213__10_ <= r_n_213__10_;
      r_213__9_ <= r_n_213__9_;
      r_213__8_ <= r_n_213__8_;
      r_213__7_ <= r_n_213__7_;
      r_213__6_ <= r_n_213__6_;
      r_213__5_ <= r_n_213__5_;
      r_213__4_ <= r_n_213__4_;
      r_213__3_ <= r_n_213__3_;
      r_213__2_ <= r_n_213__2_;
      r_213__1_ <= r_n_213__1_;
      r_213__0_ <= r_n_213__0_;
    end 
    if(N2006) begin
      r_214__31_ <= r_n_214__31_;
      r_214__30_ <= r_n_214__30_;
      r_214__29_ <= r_n_214__29_;
      r_214__28_ <= r_n_214__28_;
      r_214__27_ <= r_n_214__27_;
      r_214__26_ <= r_n_214__26_;
      r_214__25_ <= r_n_214__25_;
      r_214__24_ <= r_n_214__24_;
      r_214__23_ <= r_n_214__23_;
      r_214__22_ <= r_n_214__22_;
      r_214__21_ <= r_n_214__21_;
      r_214__20_ <= r_n_214__20_;
      r_214__19_ <= r_n_214__19_;
      r_214__18_ <= r_n_214__18_;
      r_214__17_ <= r_n_214__17_;
      r_214__16_ <= r_n_214__16_;
      r_214__15_ <= r_n_214__15_;
      r_214__14_ <= r_n_214__14_;
      r_214__13_ <= r_n_214__13_;
      r_214__12_ <= r_n_214__12_;
      r_214__11_ <= r_n_214__11_;
      r_214__10_ <= r_n_214__10_;
      r_214__9_ <= r_n_214__9_;
      r_214__8_ <= r_n_214__8_;
      r_214__7_ <= r_n_214__7_;
      r_214__6_ <= r_n_214__6_;
      r_214__5_ <= r_n_214__5_;
      r_214__4_ <= r_n_214__4_;
      r_214__3_ <= r_n_214__3_;
      r_214__2_ <= r_n_214__2_;
      r_214__1_ <= r_n_214__1_;
      r_214__0_ <= r_n_214__0_;
    end 
    if(N2007) begin
      r_215__31_ <= r_n_215__31_;
      r_215__30_ <= r_n_215__30_;
      r_215__29_ <= r_n_215__29_;
      r_215__28_ <= r_n_215__28_;
      r_215__27_ <= r_n_215__27_;
      r_215__26_ <= r_n_215__26_;
      r_215__25_ <= r_n_215__25_;
      r_215__24_ <= r_n_215__24_;
      r_215__23_ <= r_n_215__23_;
      r_215__22_ <= r_n_215__22_;
      r_215__21_ <= r_n_215__21_;
      r_215__20_ <= r_n_215__20_;
      r_215__19_ <= r_n_215__19_;
      r_215__18_ <= r_n_215__18_;
      r_215__17_ <= r_n_215__17_;
      r_215__16_ <= r_n_215__16_;
      r_215__15_ <= r_n_215__15_;
      r_215__14_ <= r_n_215__14_;
      r_215__13_ <= r_n_215__13_;
      r_215__12_ <= r_n_215__12_;
      r_215__11_ <= r_n_215__11_;
      r_215__10_ <= r_n_215__10_;
      r_215__9_ <= r_n_215__9_;
      r_215__8_ <= r_n_215__8_;
      r_215__7_ <= r_n_215__7_;
      r_215__6_ <= r_n_215__6_;
      r_215__5_ <= r_n_215__5_;
      r_215__4_ <= r_n_215__4_;
      r_215__3_ <= r_n_215__3_;
      r_215__2_ <= r_n_215__2_;
      r_215__1_ <= r_n_215__1_;
      r_215__0_ <= r_n_215__0_;
    end 
    if(N2008) begin
      r_216__31_ <= r_n_216__31_;
      r_216__30_ <= r_n_216__30_;
      r_216__29_ <= r_n_216__29_;
      r_216__28_ <= r_n_216__28_;
      r_216__27_ <= r_n_216__27_;
      r_216__26_ <= r_n_216__26_;
      r_216__25_ <= r_n_216__25_;
      r_216__24_ <= r_n_216__24_;
      r_216__23_ <= r_n_216__23_;
      r_216__22_ <= r_n_216__22_;
      r_216__21_ <= r_n_216__21_;
      r_216__20_ <= r_n_216__20_;
      r_216__19_ <= r_n_216__19_;
      r_216__18_ <= r_n_216__18_;
      r_216__17_ <= r_n_216__17_;
      r_216__16_ <= r_n_216__16_;
      r_216__15_ <= r_n_216__15_;
      r_216__14_ <= r_n_216__14_;
      r_216__13_ <= r_n_216__13_;
      r_216__12_ <= r_n_216__12_;
      r_216__11_ <= r_n_216__11_;
      r_216__10_ <= r_n_216__10_;
      r_216__9_ <= r_n_216__9_;
      r_216__8_ <= r_n_216__8_;
      r_216__7_ <= r_n_216__7_;
      r_216__6_ <= r_n_216__6_;
      r_216__5_ <= r_n_216__5_;
      r_216__4_ <= r_n_216__4_;
      r_216__3_ <= r_n_216__3_;
      r_216__2_ <= r_n_216__2_;
      r_216__1_ <= r_n_216__1_;
      r_216__0_ <= r_n_216__0_;
    end 
    if(N2009) begin
      r_217__31_ <= r_n_217__31_;
      r_217__30_ <= r_n_217__30_;
      r_217__29_ <= r_n_217__29_;
      r_217__28_ <= r_n_217__28_;
      r_217__27_ <= r_n_217__27_;
      r_217__26_ <= r_n_217__26_;
      r_217__25_ <= r_n_217__25_;
      r_217__24_ <= r_n_217__24_;
      r_217__23_ <= r_n_217__23_;
      r_217__22_ <= r_n_217__22_;
      r_217__21_ <= r_n_217__21_;
      r_217__20_ <= r_n_217__20_;
      r_217__19_ <= r_n_217__19_;
      r_217__18_ <= r_n_217__18_;
      r_217__17_ <= r_n_217__17_;
      r_217__16_ <= r_n_217__16_;
      r_217__15_ <= r_n_217__15_;
      r_217__14_ <= r_n_217__14_;
      r_217__13_ <= r_n_217__13_;
      r_217__12_ <= r_n_217__12_;
      r_217__11_ <= r_n_217__11_;
      r_217__10_ <= r_n_217__10_;
      r_217__9_ <= r_n_217__9_;
      r_217__8_ <= r_n_217__8_;
      r_217__7_ <= r_n_217__7_;
      r_217__6_ <= r_n_217__6_;
      r_217__5_ <= r_n_217__5_;
      r_217__4_ <= r_n_217__4_;
      r_217__3_ <= r_n_217__3_;
      r_217__2_ <= r_n_217__2_;
      r_217__1_ <= r_n_217__1_;
      r_217__0_ <= r_n_217__0_;
    end 
    if(N2010) begin
      r_218__31_ <= r_n_218__31_;
      r_218__30_ <= r_n_218__30_;
      r_218__29_ <= r_n_218__29_;
      r_218__28_ <= r_n_218__28_;
      r_218__27_ <= r_n_218__27_;
      r_218__26_ <= r_n_218__26_;
      r_218__25_ <= r_n_218__25_;
      r_218__24_ <= r_n_218__24_;
      r_218__23_ <= r_n_218__23_;
      r_218__22_ <= r_n_218__22_;
      r_218__21_ <= r_n_218__21_;
      r_218__20_ <= r_n_218__20_;
      r_218__19_ <= r_n_218__19_;
      r_218__18_ <= r_n_218__18_;
      r_218__17_ <= r_n_218__17_;
      r_218__16_ <= r_n_218__16_;
      r_218__15_ <= r_n_218__15_;
      r_218__14_ <= r_n_218__14_;
      r_218__13_ <= r_n_218__13_;
      r_218__12_ <= r_n_218__12_;
      r_218__11_ <= r_n_218__11_;
      r_218__10_ <= r_n_218__10_;
      r_218__9_ <= r_n_218__9_;
      r_218__8_ <= r_n_218__8_;
      r_218__7_ <= r_n_218__7_;
      r_218__6_ <= r_n_218__6_;
      r_218__5_ <= r_n_218__5_;
      r_218__4_ <= r_n_218__4_;
      r_218__3_ <= r_n_218__3_;
      r_218__2_ <= r_n_218__2_;
      r_218__1_ <= r_n_218__1_;
      r_218__0_ <= r_n_218__0_;
    end 
    if(N2011) begin
      r_219__31_ <= r_n_219__31_;
      r_219__30_ <= r_n_219__30_;
      r_219__29_ <= r_n_219__29_;
      r_219__28_ <= r_n_219__28_;
      r_219__27_ <= r_n_219__27_;
      r_219__26_ <= r_n_219__26_;
      r_219__25_ <= r_n_219__25_;
      r_219__24_ <= r_n_219__24_;
      r_219__23_ <= r_n_219__23_;
      r_219__22_ <= r_n_219__22_;
      r_219__21_ <= r_n_219__21_;
      r_219__20_ <= r_n_219__20_;
      r_219__19_ <= r_n_219__19_;
      r_219__18_ <= r_n_219__18_;
      r_219__17_ <= r_n_219__17_;
      r_219__16_ <= r_n_219__16_;
      r_219__15_ <= r_n_219__15_;
      r_219__14_ <= r_n_219__14_;
      r_219__13_ <= r_n_219__13_;
      r_219__12_ <= r_n_219__12_;
      r_219__11_ <= r_n_219__11_;
      r_219__10_ <= r_n_219__10_;
      r_219__9_ <= r_n_219__9_;
      r_219__8_ <= r_n_219__8_;
      r_219__7_ <= r_n_219__7_;
      r_219__6_ <= r_n_219__6_;
      r_219__5_ <= r_n_219__5_;
      r_219__4_ <= r_n_219__4_;
      r_219__3_ <= r_n_219__3_;
      r_219__2_ <= r_n_219__2_;
      r_219__1_ <= r_n_219__1_;
      r_219__0_ <= r_n_219__0_;
    end 
    if(N2012) begin
      r_220__31_ <= r_n_220__31_;
      r_220__30_ <= r_n_220__30_;
      r_220__29_ <= r_n_220__29_;
      r_220__28_ <= r_n_220__28_;
      r_220__27_ <= r_n_220__27_;
      r_220__26_ <= r_n_220__26_;
      r_220__25_ <= r_n_220__25_;
      r_220__24_ <= r_n_220__24_;
      r_220__23_ <= r_n_220__23_;
      r_220__22_ <= r_n_220__22_;
      r_220__21_ <= r_n_220__21_;
      r_220__20_ <= r_n_220__20_;
      r_220__19_ <= r_n_220__19_;
      r_220__18_ <= r_n_220__18_;
      r_220__17_ <= r_n_220__17_;
      r_220__16_ <= r_n_220__16_;
      r_220__15_ <= r_n_220__15_;
      r_220__14_ <= r_n_220__14_;
      r_220__13_ <= r_n_220__13_;
      r_220__12_ <= r_n_220__12_;
      r_220__11_ <= r_n_220__11_;
      r_220__10_ <= r_n_220__10_;
      r_220__9_ <= r_n_220__9_;
      r_220__8_ <= r_n_220__8_;
      r_220__7_ <= r_n_220__7_;
      r_220__6_ <= r_n_220__6_;
      r_220__5_ <= r_n_220__5_;
      r_220__4_ <= r_n_220__4_;
      r_220__3_ <= r_n_220__3_;
      r_220__2_ <= r_n_220__2_;
      r_220__1_ <= r_n_220__1_;
      r_220__0_ <= r_n_220__0_;
    end 
    if(N2013) begin
      r_221__31_ <= r_n_221__31_;
      r_221__30_ <= r_n_221__30_;
      r_221__29_ <= r_n_221__29_;
      r_221__28_ <= r_n_221__28_;
      r_221__27_ <= r_n_221__27_;
      r_221__26_ <= r_n_221__26_;
      r_221__25_ <= r_n_221__25_;
      r_221__24_ <= r_n_221__24_;
      r_221__23_ <= r_n_221__23_;
      r_221__22_ <= r_n_221__22_;
      r_221__21_ <= r_n_221__21_;
      r_221__20_ <= r_n_221__20_;
      r_221__19_ <= r_n_221__19_;
      r_221__18_ <= r_n_221__18_;
      r_221__17_ <= r_n_221__17_;
      r_221__16_ <= r_n_221__16_;
      r_221__15_ <= r_n_221__15_;
      r_221__14_ <= r_n_221__14_;
      r_221__13_ <= r_n_221__13_;
      r_221__12_ <= r_n_221__12_;
      r_221__11_ <= r_n_221__11_;
      r_221__10_ <= r_n_221__10_;
      r_221__9_ <= r_n_221__9_;
      r_221__8_ <= r_n_221__8_;
      r_221__7_ <= r_n_221__7_;
      r_221__6_ <= r_n_221__6_;
      r_221__5_ <= r_n_221__5_;
      r_221__4_ <= r_n_221__4_;
      r_221__3_ <= r_n_221__3_;
      r_221__2_ <= r_n_221__2_;
      r_221__1_ <= r_n_221__1_;
      r_221__0_ <= r_n_221__0_;
    end 
    if(N2014) begin
      r_222__31_ <= r_n_222__31_;
      r_222__30_ <= r_n_222__30_;
      r_222__29_ <= r_n_222__29_;
      r_222__28_ <= r_n_222__28_;
      r_222__27_ <= r_n_222__27_;
      r_222__26_ <= r_n_222__26_;
      r_222__25_ <= r_n_222__25_;
      r_222__24_ <= r_n_222__24_;
      r_222__23_ <= r_n_222__23_;
      r_222__22_ <= r_n_222__22_;
      r_222__21_ <= r_n_222__21_;
      r_222__20_ <= r_n_222__20_;
      r_222__19_ <= r_n_222__19_;
      r_222__18_ <= r_n_222__18_;
      r_222__17_ <= r_n_222__17_;
      r_222__16_ <= r_n_222__16_;
      r_222__15_ <= r_n_222__15_;
      r_222__14_ <= r_n_222__14_;
      r_222__13_ <= r_n_222__13_;
      r_222__12_ <= r_n_222__12_;
      r_222__11_ <= r_n_222__11_;
      r_222__10_ <= r_n_222__10_;
      r_222__9_ <= r_n_222__9_;
      r_222__8_ <= r_n_222__8_;
      r_222__7_ <= r_n_222__7_;
      r_222__6_ <= r_n_222__6_;
      r_222__5_ <= r_n_222__5_;
      r_222__4_ <= r_n_222__4_;
      r_222__3_ <= r_n_222__3_;
      r_222__2_ <= r_n_222__2_;
      r_222__1_ <= r_n_222__1_;
      r_222__0_ <= r_n_222__0_;
    end 
    if(N2015) begin
      r_223__31_ <= r_n_223__31_;
      r_223__30_ <= r_n_223__30_;
      r_223__29_ <= r_n_223__29_;
      r_223__28_ <= r_n_223__28_;
      r_223__27_ <= r_n_223__27_;
      r_223__26_ <= r_n_223__26_;
      r_223__25_ <= r_n_223__25_;
      r_223__24_ <= r_n_223__24_;
      r_223__23_ <= r_n_223__23_;
      r_223__22_ <= r_n_223__22_;
      r_223__21_ <= r_n_223__21_;
      r_223__20_ <= r_n_223__20_;
      r_223__19_ <= r_n_223__19_;
      r_223__18_ <= r_n_223__18_;
      r_223__17_ <= r_n_223__17_;
      r_223__16_ <= r_n_223__16_;
      r_223__15_ <= r_n_223__15_;
      r_223__14_ <= r_n_223__14_;
      r_223__13_ <= r_n_223__13_;
      r_223__12_ <= r_n_223__12_;
      r_223__11_ <= r_n_223__11_;
      r_223__10_ <= r_n_223__10_;
      r_223__9_ <= r_n_223__9_;
      r_223__8_ <= r_n_223__8_;
      r_223__7_ <= r_n_223__7_;
      r_223__6_ <= r_n_223__6_;
      r_223__5_ <= r_n_223__5_;
      r_223__4_ <= r_n_223__4_;
      r_223__3_ <= r_n_223__3_;
      r_223__2_ <= r_n_223__2_;
      r_223__1_ <= r_n_223__1_;
      r_223__0_ <= r_n_223__0_;
    end 
    if(N2016) begin
      r_224__31_ <= r_n_224__31_;
      r_224__30_ <= r_n_224__30_;
      r_224__29_ <= r_n_224__29_;
      r_224__28_ <= r_n_224__28_;
      r_224__27_ <= r_n_224__27_;
      r_224__26_ <= r_n_224__26_;
      r_224__25_ <= r_n_224__25_;
      r_224__24_ <= r_n_224__24_;
      r_224__23_ <= r_n_224__23_;
      r_224__22_ <= r_n_224__22_;
      r_224__21_ <= r_n_224__21_;
      r_224__20_ <= r_n_224__20_;
      r_224__19_ <= r_n_224__19_;
      r_224__18_ <= r_n_224__18_;
      r_224__17_ <= r_n_224__17_;
      r_224__16_ <= r_n_224__16_;
      r_224__15_ <= r_n_224__15_;
      r_224__14_ <= r_n_224__14_;
      r_224__13_ <= r_n_224__13_;
      r_224__12_ <= r_n_224__12_;
      r_224__11_ <= r_n_224__11_;
      r_224__10_ <= r_n_224__10_;
      r_224__9_ <= r_n_224__9_;
      r_224__8_ <= r_n_224__8_;
      r_224__7_ <= r_n_224__7_;
      r_224__6_ <= r_n_224__6_;
      r_224__5_ <= r_n_224__5_;
      r_224__4_ <= r_n_224__4_;
      r_224__3_ <= r_n_224__3_;
      r_224__2_ <= r_n_224__2_;
      r_224__1_ <= r_n_224__1_;
      r_224__0_ <= r_n_224__0_;
    end 
    if(N2017) begin
      r_225__31_ <= r_n_225__31_;
      r_225__30_ <= r_n_225__30_;
      r_225__29_ <= r_n_225__29_;
      r_225__28_ <= r_n_225__28_;
      r_225__27_ <= r_n_225__27_;
      r_225__26_ <= r_n_225__26_;
      r_225__25_ <= r_n_225__25_;
      r_225__24_ <= r_n_225__24_;
      r_225__23_ <= r_n_225__23_;
      r_225__22_ <= r_n_225__22_;
      r_225__21_ <= r_n_225__21_;
      r_225__20_ <= r_n_225__20_;
      r_225__19_ <= r_n_225__19_;
      r_225__18_ <= r_n_225__18_;
      r_225__17_ <= r_n_225__17_;
      r_225__16_ <= r_n_225__16_;
      r_225__15_ <= r_n_225__15_;
      r_225__14_ <= r_n_225__14_;
      r_225__13_ <= r_n_225__13_;
      r_225__12_ <= r_n_225__12_;
      r_225__11_ <= r_n_225__11_;
      r_225__10_ <= r_n_225__10_;
      r_225__9_ <= r_n_225__9_;
      r_225__8_ <= r_n_225__8_;
      r_225__7_ <= r_n_225__7_;
      r_225__6_ <= r_n_225__6_;
      r_225__5_ <= r_n_225__5_;
      r_225__4_ <= r_n_225__4_;
      r_225__3_ <= r_n_225__3_;
      r_225__2_ <= r_n_225__2_;
      r_225__1_ <= r_n_225__1_;
      r_225__0_ <= r_n_225__0_;
    end 
    if(N2018) begin
      r_226__31_ <= r_n_226__31_;
      r_226__30_ <= r_n_226__30_;
      r_226__29_ <= r_n_226__29_;
      r_226__28_ <= r_n_226__28_;
      r_226__27_ <= r_n_226__27_;
      r_226__26_ <= r_n_226__26_;
      r_226__25_ <= r_n_226__25_;
      r_226__24_ <= r_n_226__24_;
      r_226__23_ <= r_n_226__23_;
      r_226__22_ <= r_n_226__22_;
      r_226__21_ <= r_n_226__21_;
      r_226__20_ <= r_n_226__20_;
      r_226__19_ <= r_n_226__19_;
      r_226__18_ <= r_n_226__18_;
      r_226__17_ <= r_n_226__17_;
      r_226__16_ <= r_n_226__16_;
      r_226__15_ <= r_n_226__15_;
      r_226__14_ <= r_n_226__14_;
      r_226__13_ <= r_n_226__13_;
      r_226__12_ <= r_n_226__12_;
      r_226__11_ <= r_n_226__11_;
      r_226__10_ <= r_n_226__10_;
      r_226__9_ <= r_n_226__9_;
      r_226__8_ <= r_n_226__8_;
      r_226__7_ <= r_n_226__7_;
      r_226__6_ <= r_n_226__6_;
      r_226__5_ <= r_n_226__5_;
      r_226__4_ <= r_n_226__4_;
      r_226__3_ <= r_n_226__3_;
      r_226__2_ <= r_n_226__2_;
      r_226__1_ <= r_n_226__1_;
      r_226__0_ <= r_n_226__0_;
    end 
    if(N2019) begin
      r_227__31_ <= r_n_227__31_;
      r_227__30_ <= r_n_227__30_;
      r_227__29_ <= r_n_227__29_;
      r_227__28_ <= r_n_227__28_;
      r_227__27_ <= r_n_227__27_;
      r_227__26_ <= r_n_227__26_;
      r_227__25_ <= r_n_227__25_;
      r_227__24_ <= r_n_227__24_;
      r_227__23_ <= r_n_227__23_;
      r_227__22_ <= r_n_227__22_;
      r_227__21_ <= r_n_227__21_;
      r_227__20_ <= r_n_227__20_;
      r_227__19_ <= r_n_227__19_;
      r_227__18_ <= r_n_227__18_;
      r_227__17_ <= r_n_227__17_;
      r_227__16_ <= r_n_227__16_;
      r_227__15_ <= r_n_227__15_;
      r_227__14_ <= r_n_227__14_;
      r_227__13_ <= r_n_227__13_;
      r_227__12_ <= r_n_227__12_;
      r_227__11_ <= r_n_227__11_;
      r_227__10_ <= r_n_227__10_;
      r_227__9_ <= r_n_227__9_;
      r_227__8_ <= r_n_227__8_;
      r_227__7_ <= r_n_227__7_;
      r_227__6_ <= r_n_227__6_;
      r_227__5_ <= r_n_227__5_;
      r_227__4_ <= r_n_227__4_;
      r_227__3_ <= r_n_227__3_;
      r_227__2_ <= r_n_227__2_;
      r_227__1_ <= r_n_227__1_;
      r_227__0_ <= r_n_227__0_;
    end 
    if(N2020) begin
      r_228__31_ <= r_n_228__31_;
      r_228__30_ <= r_n_228__30_;
      r_228__29_ <= r_n_228__29_;
      r_228__28_ <= r_n_228__28_;
      r_228__27_ <= r_n_228__27_;
      r_228__26_ <= r_n_228__26_;
      r_228__25_ <= r_n_228__25_;
      r_228__24_ <= r_n_228__24_;
      r_228__23_ <= r_n_228__23_;
      r_228__22_ <= r_n_228__22_;
      r_228__21_ <= r_n_228__21_;
      r_228__20_ <= r_n_228__20_;
      r_228__19_ <= r_n_228__19_;
      r_228__18_ <= r_n_228__18_;
      r_228__17_ <= r_n_228__17_;
      r_228__16_ <= r_n_228__16_;
      r_228__15_ <= r_n_228__15_;
      r_228__14_ <= r_n_228__14_;
      r_228__13_ <= r_n_228__13_;
      r_228__12_ <= r_n_228__12_;
      r_228__11_ <= r_n_228__11_;
      r_228__10_ <= r_n_228__10_;
      r_228__9_ <= r_n_228__9_;
      r_228__8_ <= r_n_228__8_;
      r_228__7_ <= r_n_228__7_;
      r_228__6_ <= r_n_228__6_;
      r_228__5_ <= r_n_228__5_;
      r_228__4_ <= r_n_228__4_;
      r_228__3_ <= r_n_228__3_;
      r_228__2_ <= r_n_228__2_;
      r_228__1_ <= r_n_228__1_;
      r_228__0_ <= r_n_228__0_;
    end 
    if(N2021) begin
      r_229__31_ <= r_n_229__31_;
      r_229__30_ <= r_n_229__30_;
      r_229__29_ <= r_n_229__29_;
      r_229__28_ <= r_n_229__28_;
      r_229__27_ <= r_n_229__27_;
      r_229__26_ <= r_n_229__26_;
      r_229__25_ <= r_n_229__25_;
      r_229__24_ <= r_n_229__24_;
      r_229__23_ <= r_n_229__23_;
      r_229__22_ <= r_n_229__22_;
      r_229__21_ <= r_n_229__21_;
      r_229__20_ <= r_n_229__20_;
      r_229__19_ <= r_n_229__19_;
      r_229__18_ <= r_n_229__18_;
      r_229__17_ <= r_n_229__17_;
      r_229__16_ <= r_n_229__16_;
      r_229__15_ <= r_n_229__15_;
      r_229__14_ <= r_n_229__14_;
      r_229__13_ <= r_n_229__13_;
      r_229__12_ <= r_n_229__12_;
      r_229__11_ <= r_n_229__11_;
      r_229__10_ <= r_n_229__10_;
      r_229__9_ <= r_n_229__9_;
      r_229__8_ <= r_n_229__8_;
      r_229__7_ <= r_n_229__7_;
      r_229__6_ <= r_n_229__6_;
      r_229__5_ <= r_n_229__5_;
      r_229__4_ <= r_n_229__4_;
      r_229__3_ <= r_n_229__3_;
      r_229__2_ <= r_n_229__2_;
      r_229__1_ <= r_n_229__1_;
      r_229__0_ <= r_n_229__0_;
    end 
    if(N2022) begin
      r_230__31_ <= r_n_230__31_;
      r_230__30_ <= r_n_230__30_;
      r_230__29_ <= r_n_230__29_;
      r_230__28_ <= r_n_230__28_;
      r_230__27_ <= r_n_230__27_;
      r_230__26_ <= r_n_230__26_;
      r_230__25_ <= r_n_230__25_;
      r_230__24_ <= r_n_230__24_;
      r_230__23_ <= r_n_230__23_;
      r_230__22_ <= r_n_230__22_;
      r_230__21_ <= r_n_230__21_;
      r_230__20_ <= r_n_230__20_;
      r_230__19_ <= r_n_230__19_;
      r_230__18_ <= r_n_230__18_;
      r_230__17_ <= r_n_230__17_;
      r_230__16_ <= r_n_230__16_;
      r_230__15_ <= r_n_230__15_;
      r_230__14_ <= r_n_230__14_;
      r_230__13_ <= r_n_230__13_;
      r_230__12_ <= r_n_230__12_;
      r_230__11_ <= r_n_230__11_;
      r_230__10_ <= r_n_230__10_;
      r_230__9_ <= r_n_230__9_;
      r_230__8_ <= r_n_230__8_;
      r_230__7_ <= r_n_230__7_;
      r_230__6_ <= r_n_230__6_;
      r_230__5_ <= r_n_230__5_;
      r_230__4_ <= r_n_230__4_;
      r_230__3_ <= r_n_230__3_;
      r_230__2_ <= r_n_230__2_;
      r_230__1_ <= r_n_230__1_;
      r_230__0_ <= r_n_230__0_;
    end 
    if(N2023) begin
      r_231__31_ <= r_n_231__31_;
      r_231__30_ <= r_n_231__30_;
      r_231__29_ <= r_n_231__29_;
      r_231__28_ <= r_n_231__28_;
      r_231__27_ <= r_n_231__27_;
      r_231__26_ <= r_n_231__26_;
      r_231__25_ <= r_n_231__25_;
      r_231__24_ <= r_n_231__24_;
      r_231__23_ <= r_n_231__23_;
      r_231__22_ <= r_n_231__22_;
      r_231__21_ <= r_n_231__21_;
      r_231__20_ <= r_n_231__20_;
      r_231__19_ <= r_n_231__19_;
      r_231__18_ <= r_n_231__18_;
      r_231__17_ <= r_n_231__17_;
      r_231__16_ <= r_n_231__16_;
      r_231__15_ <= r_n_231__15_;
      r_231__14_ <= r_n_231__14_;
      r_231__13_ <= r_n_231__13_;
      r_231__12_ <= r_n_231__12_;
      r_231__11_ <= r_n_231__11_;
      r_231__10_ <= r_n_231__10_;
      r_231__9_ <= r_n_231__9_;
      r_231__8_ <= r_n_231__8_;
      r_231__7_ <= r_n_231__7_;
      r_231__6_ <= r_n_231__6_;
      r_231__5_ <= r_n_231__5_;
      r_231__4_ <= r_n_231__4_;
      r_231__3_ <= r_n_231__3_;
      r_231__2_ <= r_n_231__2_;
      r_231__1_ <= r_n_231__1_;
      r_231__0_ <= r_n_231__0_;
    end 
    if(N2024) begin
      r_232__31_ <= r_n_232__31_;
      r_232__30_ <= r_n_232__30_;
      r_232__29_ <= r_n_232__29_;
      r_232__28_ <= r_n_232__28_;
      r_232__27_ <= r_n_232__27_;
      r_232__26_ <= r_n_232__26_;
      r_232__25_ <= r_n_232__25_;
      r_232__24_ <= r_n_232__24_;
      r_232__23_ <= r_n_232__23_;
      r_232__22_ <= r_n_232__22_;
      r_232__21_ <= r_n_232__21_;
      r_232__20_ <= r_n_232__20_;
      r_232__19_ <= r_n_232__19_;
      r_232__18_ <= r_n_232__18_;
      r_232__17_ <= r_n_232__17_;
      r_232__16_ <= r_n_232__16_;
      r_232__15_ <= r_n_232__15_;
      r_232__14_ <= r_n_232__14_;
      r_232__13_ <= r_n_232__13_;
      r_232__12_ <= r_n_232__12_;
      r_232__11_ <= r_n_232__11_;
      r_232__10_ <= r_n_232__10_;
      r_232__9_ <= r_n_232__9_;
      r_232__8_ <= r_n_232__8_;
      r_232__7_ <= r_n_232__7_;
      r_232__6_ <= r_n_232__6_;
      r_232__5_ <= r_n_232__5_;
      r_232__4_ <= r_n_232__4_;
      r_232__3_ <= r_n_232__3_;
      r_232__2_ <= r_n_232__2_;
      r_232__1_ <= r_n_232__1_;
      r_232__0_ <= r_n_232__0_;
    end 
    if(N2025) begin
      r_233__31_ <= r_n_233__31_;
      r_233__30_ <= r_n_233__30_;
      r_233__29_ <= r_n_233__29_;
      r_233__28_ <= r_n_233__28_;
      r_233__27_ <= r_n_233__27_;
      r_233__26_ <= r_n_233__26_;
      r_233__25_ <= r_n_233__25_;
      r_233__24_ <= r_n_233__24_;
      r_233__23_ <= r_n_233__23_;
      r_233__22_ <= r_n_233__22_;
      r_233__21_ <= r_n_233__21_;
      r_233__20_ <= r_n_233__20_;
      r_233__19_ <= r_n_233__19_;
      r_233__18_ <= r_n_233__18_;
      r_233__17_ <= r_n_233__17_;
      r_233__16_ <= r_n_233__16_;
      r_233__15_ <= r_n_233__15_;
      r_233__14_ <= r_n_233__14_;
      r_233__13_ <= r_n_233__13_;
      r_233__12_ <= r_n_233__12_;
      r_233__11_ <= r_n_233__11_;
      r_233__10_ <= r_n_233__10_;
      r_233__9_ <= r_n_233__9_;
      r_233__8_ <= r_n_233__8_;
      r_233__7_ <= r_n_233__7_;
      r_233__6_ <= r_n_233__6_;
      r_233__5_ <= r_n_233__5_;
      r_233__4_ <= r_n_233__4_;
      r_233__3_ <= r_n_233__3_;
      r_233__2_ <= r_n_233__2_;
      r_233__1_ <= r_n_233__1_;
      r_233__0_ <= r_n_233__0_;
    end 
    if(N2026) begin
      r_234__31_ <= r_n_234__31_;
      r_234__30_ <= r_n_234__30_;
      r_234__29_ <= r_n_234__29_;
      r_234__28_ <= r_n_234__28_;
      r_234__27_ <= r_n_234__27_;
      r_234__26_ <= r_n_234__26_;
      r_234__25_ <= r_n_234__25_;
      r_234__24_ <= r_n_234__24_;
      r_234__23_ <= r_n_234__23_;
      r_234__22_ <= r_n_234__22_;
      r_234__21_ <= r_n_234__21_;
      r_234__20_ <= r_n_234__20_;
      r_234__19_ <= r_n_234__19_;
      r_234__18_ <= r_n_234__18_;
      r_234__17_ <= r_n_234__17_;
      r_234__16_ <= r_n_234__16_;
      r_234__15_ <= r_n_234__15_;
      r_234__14_ <= r_n_234__14_;
      r_234__13_ <= r_n_234__13_;
      r_234__12_ <= r_n_234__12_;
      r_234__11_ <= r_n_234__11_;
      r_234__10_ <= r_n_234__10_;
      r_234__9_ <= r_n_234__9_;
      r_234__8_ <= r_n_234__8_;
      r_234__7_ <= r_n_234__7_;
      r_234__6_ <= r_n_234__6_;
      r_234__5_ <= r_n_234__5_;
      r_234__4_ <= r_n_234__4_;
      r_234__3_ <= r_n_234__3_;
      r_234__2_ <= r_n_234__2_;
      r_234__1_ <= r_n_234__1_;
      r_234__0_ <= r_n_234__0_;
    end 
    if(N2027) begin
      r_235__31_ <= r_n_235__31_;
      r_235__30_ <= r_n_235__30_;
      r_235__29_ <= r_n_235__29_;
      r_235__28_ <= r_n_235__28_;
      r_235__27_ <= r_n_235__27_;
      r_235__26_ <= r_n_235__26_;
      r_235__25_ <= r_n_235__25_;
      r_235__24_ <= r_n_235__24_;
      r_235__23_ <= r_n_235__23_;
      r_235__22_ <= r_n_235__22_;
      r_235__21_ <= r_n_235__21_;
      r_235__20_ <= r_n_235__20_;
      r_235__19_ <= r_n_235__19_;
      r_235__18_ <= r_n_235__18_;
      r_235__17_ <= r_n_235__17_;
      r_235__16_ <= r_n_235__16_;
      r_235__15_ <= r_n_235__15_;
      r_235__14_ <= r_n_235__14_;
      r_235__13_ <= r_n_235__13_;
      r_235__12_ <= r_n_235__12_;
      r_235__11_ <= r_n_235__11_;
      r_235__10_ <= r_n_235__10_;
      r_235__9_ <= r_n_235__9_;
      r_235__8_ <= r_n_235__8_;
      r_235__7_ <= r_n_235__7_;
      r_235__6_ <= r_n_235__6_;
      r_235__5_ <= r_n_235__5_;
      r_235__4_ <= r_n_235__4_;
      r_235__3_ <= r_n_235__3_;
      r_235__2_ <= r_n_235__2_;
      r_235__1_ <= r_n_235__1_;
      r_235__0_ <= r_n_235__0_;
    end 
    if(N2028) begin
      r_236__31_ <= r_n_236__31_;
      r_236__30_ <= r_n_236__30_;
      r_236__29_ <= r_n_236__29_;
      r_236__28_ <= r_n_236__28_;
      r_236__27_ <= r_n_236__27_;
      r_236__26_ <= r_n_236__26_;
      r_236__25_ <= r_n_236__25_;
      r_236__24_ <= r_n_236__24_;
      r_236__23_ <= r_n_236__23_;
      r_236__22_ <= r_n_236__22_;
      r_236__21_ <= r_n_236__21_;
      r_236__20_ <= r_n_236__20_;
      r_236__19_ <= r_n_236__19_;
      r_236__18_ <= r_n_236__18_;
      r_236__17_ <= r_n_236__17_;
      r_236__16_ <= r_n_236__16_;
      r_236__15_ <= r_n_236__15_;
      r_236__14_ <= r_n_236__14_;
      r_236__13_ <= r_n_236__13_;
      r_236__12_ <= r_n_236__12_;
      r_236__11_ <= r_n_236__11_;
      r_236__10_ <= r_n_236__10_;
      r_236__9_ <= r_n_236__9_;
      r_236__8_ <= r_n_236__8_;
      r_236__7_ <= r_n_236__7_;
      r_236__6_ <= r_n_236__6_;
      r_236__5_ <= r_n_236__5_;
      r_236__4_ <= r_n_236__4_;
      r_236__3_ <= r_n_236__3_;
      r_236__2_ <= r_n_236__2_;
      r_236__1_ <= r_n_236__1_;
      r_236__0_ <= r_n_236__0_;
    end 
    if(N2029) begin
      r_237__31_ <= r_n_237__31_;
      r_237__30_ <= r_n_237__30_;
      r_237__29_ <= r_n_237__29_;
      r_237__28_ <= r_n_237__28_;
      r_237__27_ <= r_n_237__27_;
      r_237__26_ <= r_n_237__26_;
      r_237__25_ <= r_n_237__25_;
      r_237__24_ <= r_n_237__24_;
      r_237__23_ <= r_n_237__23_;
      r_237__22_ <= r_n_237__22_;
      r_237__21_ <= r_n_237__21_;
      r_237__20_ <= r_n_237__20_;
      r_237__19_ <= r_n_237__19_;
      r_237__18_ <= r_n_237__18_;
      r_237__17_ <= r_n_237__17_;
      r_237__16_ <= r_n_237__16_;
      r_237__15_ <= r_n_237__15_;
      r_237__14_ <= r_n_237__14_;
      r_237__13_ <= r_n_237__13_;
      r_237__12_ <= r_n_237__12_;
      r_237__11_ <= r_n_237__11_;
      r_237__10_ <= r_n_237__10_;
      r_237__9_ <= r_n_237__9_;
      r_237__8_ <= r_n_237__8_;
      r_237__7_ <= r_n_237__7_;
      r_237__6_ <= r_n_237__6_;
      r_237__5_ <= r_n_237__5_;
      r_237__4_ <= r_n_237__4_;
      r_237__3_ <= r_n_237__3_;
      r_237__2_ <= r_n_237__2_;
      r_237__1_ <= r_n_237__1_;
      r_237__0_ <= r_n_237__0_;
    end 
    if(N2030) begin
      r_238__31_ <= r_n_238__31_;
      r_238__30_ <= r_n_238__30_;
      r_238__29_ <= r_n_238__29_;
      r_238__28_ <= r_n_238__28_;
      r_238__27_ <= r_n_238__27_;
      r_238__26_ <= r_n_238__26_;
      r_238__25_ <= r_n_238__25_;
      r_238__24_ <= r_n_238__24_;
      r_238__23_ <= r_n_238__23_;
      r_238__22_ <= r_n_238__22_;
      r_238__21_ <= r_n_238__21_;
      r_238__20_ <= r_n_238__20_;
      r_238__19_ <= r_n_238__19_;
      r_238__18_ <= r_n_238__18_;
      r_238__17_ <= r_n_238__17_;
      r_238__16_ <= r_n_238__16_;
      r_238__15_ <= r_n_238__15_;
      r_238__14_ <= r_n_238__14_;
      r_238__13_ <= r_n_238__13_;
      r_238__12_ <= r_n_238__12_;
      r_238__11_ <= r_n_238__11_;
      r_238__10_ <= r_n_238__10_;
      r_238__9_ <= r_n_238__9_;
      r_238__8_ <= r_n_238__8_;
      r_238__7_ <= r_n_238__7_;
      r_238__6_ <= r_n_238__6_;
      r_238__5_ <= r_n_238__5_;
      r_238__4_ <= r_n_238__4_;
      r_238__3_ <= r_n_238__3_;
      r_238__2_ <= r_n_238__2_;
      r_238__1_ <= r_n_238__1_;
      r_238__0_ <= r_n_238__0_;
    end 
    if(N2031) begin
      r_239__31_ <= r_n_239__31_;
      r_239__30_ <= r_n_239__30_;
      r_239__29_ <= r_n_239__29_;
      r_239__28_ <= r_n_239__28_;
      r_239__27_ <= r_n_239__27_;
      r_239__26_ <= r_n_239__26_;
      r_239__25_ <= r_n_239__25_;
      r_239__24_ <= r_n_239__24_;
      r_239__23_ <= r_n_239__23_;
      r_239__22_ <= r_n_239__22_;
      r_239__21_ <= r_n_239__21_;
      r_239__20_ <= r_n_239__20_;
      r_239__19_ <= r_n_239__19_;
      r_239__18_ <= r_n_239__18_;
      r_239__17_ <= r_n_239__17_;
      r_239__16_ <= r_n_239__16_;
      r_239__15_ <= r_n_239__15_;
      r_239__14_ <= r_n_239__14_;
      r_239__13_ <= r_n_239__13_;
      r_239__12_ <= r_n_239__12_;
      r_239__11_ <= r_n_239__11_;
      r_239__10_ <= r_n_239__10_;
      r_239__9_ <= r_n_239__9_;
      r_239__8_ <= r_n_239__8_;
      r_239__7_ <= r_n_239__7_;
      r_239__6_ <= r_n_239__6_;
      r_239__5_ <= r_n_239__5_;
      r_239__4_ <= r_n_239__4_;
      r_239__3_ <= r_n_239__3_;
      r_239__2_ <= r_n_239__2_;
      r_239__1_ <= r_n_239__1_;
      r_239__0_ <= r_n_239__0_;
    end 
    if(N2032) begin
      r_240__31_ <= r_n_240__31_;
      r_240__30_ <= r_n_240__30_;
      r_240__29_ <= r_n_240__29_;
      r_240__28_ <= r_n_240__28_;
      r_240__27_ <= r_n_240__27_;
      r_240__26_ <= r_n_240__26_;
      r_240__25_ <= r_n_240__25_;
      r_240__24_ <= r_n_240__24_;
      r_240__23_ <= r_n_240__23_;
      r_240__22_ <= r_n_240__22_;
      r_240__21_ <= r_n_240__21_;
      r_240__20_ <= r_n_240__20_;
      r_240__19_ <= r_n_240__19_;
      r_240__18_ <= r_n_240__18_;
      r_240__17_ <= r_n_240__17_;
      r_240__16_ <= r_n_240__16_;
      r_240__15_ <= r_n_240__15_;
      r_240__14_ <= r_n_240__14_;
      r_240__13_ <= r_n_240__13_;
      r_240__12_ <= r_n_240__12_;
      r_240__11_ <= r_n_240__11_;
      r_240__10_ <= r_n_240__10_;
      r_240__9_ <= r_n_240__9_;
      r_240__8_ <= r_n_240__8_;
      r_240__7_ <= r_n_240__7_;
      r_240__6_ <= r_n_240__6_;
      r_240__5_ <= r_n_240__5_;
      r_240__4_ <= r_n_240__4_;
      r_240__3_ <= r_n_240__3_;
      r_240__2_ <= r_n_240__2_;
      r_240__1_ <= r_n_240__1_;
      r_240__0_ <= r_n_240__0_;
    end 
    if(N2033) begin
      r_241__31_ <= r_n_241__31_;
      r_241__30_ <= r_n_241__30_;
      r_241__29_ <= r_n_241__29_;
      r_241__28_ <= r_n_241__28_;
      r_241__27_ <= r_n_241__27_;
      r_241__26_ <= r_n_241__26_;
      r_241__25_ <= r_n_241__25_;
      r_241__24_ <= r_n_241__24_;
      r_241__23_ <= r_n_241__23_;
      r_241__22_ <= r_n_241__22_;
      r_241__21_ <= r_n_241__21_;
      r_241__20_ <= r_n_241__20_;
      r_241__19_ <= r_n_241__19_;
      r_241__18_ <= r_n_241__18_;
      r_241__17_ <= r_n_241__17_;
      r_241__16_ <= r_n_241__16_;
      r_241__15_ <= r_n_241__15_;
      r_241__14_ <= r_n_241__14_;
      r_241__13_ <= r_n_241__13_;
      r_241__12_ <= r_n_241__12_;
      r_241__11_ <= r_n_241__11_;
      r_241__10_ <= r_n_241__10_;
      r_241__9_ <= r_n_241__9_;
      r_241__8_ <= r_n_241__8_;
      r_241__7_ <= r_n_241__7_;
      r_241__6_ <= r_n_241__6_;
      r_241__5_ <= r_n_241__5_;
      r_241__4_ <= r_n_241__4_;
      r_241__3_ <= r_n_241__3_;
      r_241__2_ <= r_n_241__2_;
      r_241__1_ <= r_n_241__1_;
      r_241__0_ <= r_n_241__0_;
    end 
    if(N2034) begin
      r_242__31_ <= r_n_242__31_;
      r_242__30_ <= r_n_242__30_;
      r_242__29_ <= r_n_242__29_;
      r_242__28_ <= r_n_242__28_;
      r_242__27_ <= r_n_242__27_;
      r_242__26_ <= r_n_242__26_;
      r_242__25_ <= r_n_242__25_;
      r_242__24_ <= r_n_242__24_;
      r_242__23_ <= r_n_242__23_;
      r_242__22_ <= r_n_242__22_;
      r_242__21_ <= r_n_242__21_;
      r_242__20_ <= r_n_242__20_;
      r_242__19_ <= r_n_242__19_;
      r_242__18_ <= r_n_242__18_;
      r_242__17_ <= r_n_242__17_;
      r_242__16_ <= r_n_242__16_;
      r_242__15_ <= r_n_242__15_;
      r_242__14_ <= r_n_242__14_;
      r_242__13_ <= r_n_242__13_;
      r_242__12_ <= r_n_242__12_;
      r_242__11_ <= r_n_242__11_;
      r_242__10_ <= r_n_242__10_;
      r_242__9_ <= r_n_242__9_;
      r_242__8_ <= r_n_242__8_;
      r_242__7_ <= r_n_242__7_;
      r_242__6_ <= r_n_242__6_;
      r_242__5_ <= r_n_242__5_;
      r_242__4_ <= r_n_242__4_;
      r_242__3_ <= r_n_242__3_;
      r_242__2_ <= r_n_242__2_;
      r_242__1_ <= r_n_242__1_;
      r_242__0_ <= r_n_242__0_;
    end 
    if(N2035) begin
      r_243__31_ <= r_n_243__31_;
      r_243__30_ <= r_n_243__30_;
      r_243__29_ <= r_n_243__29_;
      r_243__28_ <= r_n_243__28_;
      r_243__27_ <= r_n_243__27_;
      r_243__26_ <= r_n_243__26_;
      r_243__25_ <= r_n_243__25_;
      r_243__24_ <= r_n_243__24_;
      r_243__23_ <= r_n_243__23_;
      r_243__22_ <= r_n_243__22_;
      r_243__21_ <= r_n_243__21_;
      r_243__20_ <= r_n_243__20_;
      r_243__19_ <= r_n_243__19_;
      r_243__18_ <= r_n_243__18_;
      r_243__17_ <= r_n_243__17_;
      r_243__16_ <= r_n_243__16_;
      r_243__15_ <= r_n_243__15_;
      r_243__14_ <= r_n_243__14_;
      r_243__13_ <= r_n_243__13_;
      r_243__12_ <= r_n_243__12_;
      r_243__11_ <= r_n_243__11_;
      r_243__10_ <= r_n_243__10_;
      r_243__9_ <= r_n_243__9_;
      r_243__8_ <= r_n_243__8_;
      r_243__7_ <= r_n_243__7_;
      r_243__6_ <= r_n_243__6_;
      r_243__5_ <= r_n_243__5_;
      r_243__4_ <= r_n_243__4_;
      r_243__3_ <= r_n_243__3_;
      r_243__2_ <= r_n_243__2_;
      r_243__1_ <= r_n_243__1_;
      r_243__0_ <= r_n_243__0_;
    end 
    if(N2036) begin
      r_244__31_ <= r_n_244__31_;
      r_244__30_ <= r_n_244__30_;
      r_244__29_ <= r_n_244__29_;
      r_244__28_ <= r_n_244__28_;
      r_244__27_ <= r_n_244__27_;
      r_244__26_ <= r_n_244__26_;
      r_244__25_ <= r_n_244__25_;
      r_244__24_ <= r_n_244__24_;
      r_244__23_ <= r_n_244__23_;
      r_244__22_ <= r_n_244__22_;
      r_244__21_ <= r_n_244__21_;
      r_244__20_ <= r_n_244__20_;
      r_244__19_ <= r_n_244__19_;
      r_244__18_ <= r_n_244__18_;
      r_244__17_ <= r_n_244__17_;
      r_244__16_ <= r_n_244__16_;
      r_244__15_ <= r_n_244__15_;
      r_244__14_ <= r_n_244__14_;
      r_244__13_ <= r_n_244__13_;
      r_244__12_ <= r_n_244__12_;
      r_244__11_ <= r_n_244__11_;
      r_244__10_ <= r_n_244__10_;
      r_244__9_ <= r_n_244__9_;
      r_244__8_ <= r_n_244__8_;
      r_244__7_ <= r_n_244__7_;
      r_244__6_ <= r_n_244__6_;
      r_244__5_ <= r_n_244__5_;
      r_244__4_ <= r_n_244__4_;
      r_244__3_ <= r_n_244__3_;
      r_244__2_ <= r_n_244__2_;
      r_244__1_ <= r_n_244__1_;
      r_244__0_ <= r_n_244__0_;
    end 
    if(N2037) begin
      r_245__31_ <= r_n_245__31_;
      r_245__30_ <= r_n_245__30_;
      r_245__29_ <= r_n_245__29_;
      r_245__28_ <= r_n_245__28_;
      r_245__27_ <= r_n_245__27_;
      r_245__26_ <= r_n_245__26_;
      r_245__25_ <= r_n_245__25_;
      r_245__24_ <= r_n_245__24_;
      r_245__23_ <= r_n_245__23_;
      r_245__22_ <= r_n_245__22_;
      r_245__21_ <= r_n_245__21_;
      r_245__20_ <= r_n_245__20_;
      r_245__19_ <= r_n_245__19_;
      r_245__18_ <= r_n_245__18_;
      r_245__17_ <= r_n_245__17_;
      r_245__16_ <= r_n_245__16_;
      r_245__15_ <= r_n_245__15_;
      r_245__14_ <= r_n_245__14_;
      r_245__13_ <= r_n_245__13_;
      r_245__12_ <= r_n_245__12_;
      r_245__11_ <= r_n_245__11_;
      r_245__10_ <= r_n_245__10_;
      r_245__9_ <= r_n_245__9_;
      r_245__8_ <= r_n_245__8_;
      r_245__7_ <= r_n_245__7_;
      r_245__6_ <= r_n_245__6_;
      r_245__5_ <= r_n_245__5_;
      r_245__4_ <= r_n_245__4_;
      r_245__3_ <= r_n_245__3_;
      r_245__2_ <= r_n_245__2_;
      r_245__1_ <= r_n_245__1_;
      r_245__0_ <= r_n_245__0_;
    end 
    if(N2038) begin
      r_246__31_ <= r_n_246__31_;
      r_246__30_ <= r_n_246__30_;
      r_246__29_ <= r_n_246__29_;
      r_246__28_ <= r_n_246__28_;
      r_246__27_ <= r_n_246__27_;
      r_246__26_ <= r_n_246__26_;
      r_246__25_ <= r_n_246__25_;
      r_246__24_ <= r_n_246__24_;
      r_246__23_ <= r_n_246__23_;
      r_246__22_ <= r_n_246__22_;
      r_246__21_ <= r_n_246__21_;
      r_246__20_ <= r_n_246__20_;
      r_246__19_ <= r_n_246__19_;
      r_246__18_ <= r_n_246__18_;
      r_246__17_ <= r_n_246__17_;
      r_246__16_ <= r_n_246__16_;
      r_246__15_ <= r_n_246__15_;
      r_246__14_ <= r_n_246__14_;
      r_246__13_ <= r_n_246__13_;
      r_246__12_ <= r_n_246__12_;
      r_246__11_ <= r_n_246__11_;
      r_246__10_ <= r_n_246__10_;
      r_246__9_ <= r_n_246__9_;
      r_246__8_ <= r_n_246__8_;
      r_246__7_ <= r_n_246__7_;
      r_246__6_ <= r_n_246__6_;
      r_246__5_ <= r_n_246__5_;
      r_246__4_ <= r_n_246__4_;
      r_246__3_ <= r_n_246__3_;
      r_246__2_ <= r_n_246__2_;
      r_246__1_ <= r_n_246__1_;
      r_246__0_ <= r_n_246__0_;
    end 
    if(N2039) begin
      r_247__31_ <= r_n_247__31_;
      r_247__30_ <= r_n_247__30_;
      r_247__29_ <= r_n_247__29_;
      r_247__28_ <= r_n_247__28_;
      r_247__27_ <= r_n_247__27_;
      r_247__26_ <= r_n_247__26_;
      r_247__25_ <= r_n_247__25_;
      r_247__24_ <= r_n_247__24_;
      r_247__23_ <= r_n_247__23_;
      r_247__22_ <= r_n_247__22_;
      r_247__21_ <= r_n_247__21_;
      r_247__20_ <= r_n_247__20_;
      r_247__19_ <= r_n_247__19_;
      r_247__18_ <= r_n_247__18_;
      r_247__17_ <= r_n_247__17_;
      r_247__16_ <= r_n_247__16_;
      r_247__15_ <= r_n_247__15_;
      r_247__14_ <= r_n_247__14_;
      r_247__13_ <= r_n_247__13_;
      r_247__12_ <= r_n_247__12_;
      r_247__11_ <= r_n_247__11_;
      r_247__10_ <= r_n_247__10_;
      r_247__9_ <= r_n_247__9_;
      r_247__8_ <= r_n_247__8_;
      r_247__7_ <= r_n_247__7_;
      r_247__6_ <= r_n_247__6_;
      r_247__5_ <= r_n_247__5_;
      r_247__4_ <= r_n_247__4_;
      r_247__3_ <= r_n_247__3_;
      r_247__2_ <= r_n_247__2_;
      r_247__1_ <= r_n_247__1_;
      r_247__0_ <= r_n_247__0_;
    end 
    if(N2040) begin
      r_248__31_ <= r_n_248__31_;
      r_248__30_ <= r_n_248__30_;
      r_248__29_ <= r_n_248__29_;
      r_248__28_ <= r_n_248__28_;
      r_248__27_ <= r_n_248__27_;
      r_248__26_ <= r_n_248__26_;
      r_248__25_ <= r_n_248__25_;
      r_248__24_ <= r_n_248__24_;
      r_248__23_ <= r_n_248__23_;
      r_248__22_ <= r_n_248__22_;
      r_248__21_ <= r_n_248__21_;
      r_248__20_ <= r_n_248__20_;
      r_248__19_ <= r_n_248__19_;
      r_248__18_ <= r_n_248__18_;
      r_248__17_ <= r_n_248__17_;
      r_248__16_ <= r_n_248__16_;
      r_248__15_ <= r_n_248__15_;
      r_248__14_ <= r_n_248__14_;
      r_248__13_ <= r_n_248__13_;
      r_248__12_ <= r_n_248__12_;
      r_248__11_ <= r_n_248__11_;
      r_248__10_ <= r_n_248__10_;
      r_248__9_ <= r_n_248__9_;
      r_248__8_ <= r_n_248__8_;
      r_248__7_ <= r_n_248__7_;
      r_248__6_ <= r_n_248__6_;
      r_248__5_ <= r_n_248__5_;
      r_248__4_ <= r_n_248__4_;
      r_248__3_ <= r_n_248__3_;
      r_248__2_ <= r_n_248__2_;
      r_248__1_ <= r_n_248__1_;
      r_248__0_ <= r_n_248__0_;
    end 
    if(N2041) begin
      r_249__31_ <= r_n_249__31_;
      r_249__30_ <= r_n_249__30_;
      r_249__29_ <= r_n_249__29_;
      r_249__28_ <= r_n_249__28_;
      r_249__27_ <= r_n_249__27_;
      r_249__26_ <= r_n_249__26_;
      r_249__25_ <= r_n_249__25_;
      r_249__24_ <= r_n_249__24_;
      r_249__23_ <= r_n_249__23_;
      r_249__22_ <= r_n_249__22_;
      r_249__21_ <= r_n_249__21_;
      r_249__20_ <= r_n_249__20_;
      r_249__19_ <= r_n_249__19_;
      r_249__18_ <= r_n_249__18_;
      r_249__17_ <= r_n_249__17_;
      r_249__16_ <= r_n_249__16_;
      r_249__15_ <= r_n_249__15_;
      r_249__14_ <= r_n_249__14_;
      r_249__13_ <= r_n_249__13_;
      r_249__12_ <= r_n_249__12_;
      r_249__11_ <= r_n_249__11_;
      r_249__10_ <= r_n_249__10_;
      r_249__9_ <= r_n_249__9_;
      r_249__8_ <= r_n_249__8_;
      r_249__7_ <= r_n_249__7_;
      r_249__6_ <= r_n_249__6_;
      r_249__5_ <= r_n_249__5_;
      r_249__4_ <= r_n_249__4_;
      r_249__3_ <= r_n_249__3_;
      r_249__2_ <= r_n_249__2_;
      r_249__1_ <= r_n_249__1_;
      r_249__0_ <= r_n_249__0_;
    end 
    if(N2042) begin
      r_250__31_ <= r_n_250__31_;
      r_250__30_ <= r_n_250__30_;
      r_250__29_ <= r_n_250__29_;
      r_250__28_ <= r_n_250__28_;
      r_250__27_ <= r_n_250__27_;
      r_250__26_ <= r_n_250__26_;
      r_250__25_ <= r_n_250__25_;
      r_250__24_ <= r_n_250__24_;
      r_250__23_ <= r_n_250__23_;
      r_250__22_ <= r_n_250__22_;
      r_250__21_ <= r_n_250__21_;
      r_250__20_ <= r_n_250__20_;
      r_250__19_ <= r_n_250__19_;
      r_250__18_ <= r_n_250__18_;
      r_250__17_ <= r_n_250__17_;
      r_250__16_ <= r_n_250__16_;
      r_250__15_ <= r_n_250__15_;
      r_250__14_ <= r_n_250__14_;
      r_250__13_ <= r_n_250__13_;
      r_250__12_ <= r_n_250__12_;
      r_250__11_ <= r_n_250__11_;
      r_250__10_ <= r_n_250__10_;
      r_250__9_ <= r_n_250__9_;
      r_250__8_ <= r_n_250__8_;
      r_250__7_ <= r_n_250__7_;
      r_250__6_ <= r_n_250__6_;
      r_250__5_ <= r_n_250__5_;
      r_250__4_ <= r_n_250__4_;
      r_250__3_ <= r_n_250__3_;
      r_250__2_ <= r_n_250__2_;
      r_250__1_ <= r_n_250__1_;
      r_250__0_ <= r_n_250__0_;
    end 
    if(N2043) begin
      r_251__31_ <= r_n_251__31_;
      r_251__30_ <= r_n_251__30_;
      r_251__29_ <= r_n_251__29_;
      r_251__28_ <= r_n_251__28_;
      r_251__27_ <= r_n_251__27_;
      r_251__26_ <= r_n_251__26_;
      r_251__25_ <= r_n_251__25_;
      r_251__24_ <= r_n_251__24_;
      r_251__23_ <= r_n_251__23_;
      r_251__22_ <= r_n_251__22_;
      r_251__21_ <= r_n_251__21_;
      r_251__20_ <= r_n_251__20_;
      r_251__19_ <= r_n_251__19_;
      r_251__18_ <= r_n_251__18_;
      r_251__17_ <= r_n_251__17_;
      r_251__16_ <= r_n_251__16_;
      r_251__15_ <= r_n_251__15_;
      r_251__14_ <= r_n_251__14_;
      r_251__13_ <= r_n_251__13_;
      r_251__12_ <= r_n_251__12_;
      r_251__11_ <= r_n_251__11_;
      r_251__10_ <= r_n_251__10_;
      r_251__9_ <= r_n_251__9_;
      r_251__8_ <= r_n_251__8_;
      r_251__7_ <= r_n_251__7_;
      r_251__6_ <= r_n_251__6_;
      r_251__5_ <= r_n_251__5_;
      r_251__4_ <= r_n_251__4_;
      r_251__3_ <= r_n_251__3_;
      r_251__2_ <= r_n_251__2_;
      r_251__1_ <= r_n_251__1_;
      r_251__0_ <= r_n_251__0_;
    end 
    if(N2044) begin
      r_252__31_ <= r_n_252__31_;
      r_252__30_ <= r_n_252__30_;
      r_252__29_ <= r_n_252__29_;
      r_252__28_ <= r_n_252__28_;
      r_252__27_ <= r_n_252__27_;
      r_252__26_ <= r_n_252__26_;
      r_252__25_ <= r_n_252__25_;
      r_252__24_ <= r_n_252__24_;
      r_252__23_ <= r_n_252__23_;
      r_252__22_ <= r_n_252__22_;
      r_252__21_ <= r_n_252__21_;
      r_252__20_ <= r_n_252__20_;
      r_252__19_ <= r_n_252__19_;
      r_252__18_ <= r_n_252__18_;
      r_252__17_ <= r_n_252__17_;
      r_252__16_ <= r_n_252__16_;
      r_252__15_ <= r_n_252__15_;
      r_252__14_ <= r_n_252__14_;
      r_252__13_ <= r_n_252__13_;
      r_252__12_ <= r_n_252__12_;
      r_252__11_ <= r_n_252__11_;
      r_252__10_ <= r_n_252__10_;
      r_252__9_ <= r_n_252__9_;
      r_252__8_ <= r_n_252__8_;
      r_252__7_ <= r_n_252__7_;
      r_252__6_ <= r_n_252__6_;
      r_252__5_ <= r_n_252__5_;
      r_252__4_ <= r_n_252__4_;
      r_252__3_ <= r_n_252__3_;
      r_252__2_ <= r_n_252__2_;
      r_252__1_ <= r_n_252__1_;
      r_252__0_ <= r_n_252__0_;
    end 
    if(N2045) begin
      r_253__31_ <= r_n_253__31_;
      r_253__30_ <= r_n_253__30_;
      r_253__29_ <= r_n_253__29_;
      r_253__28_ <= r_n_253__28_;
      r_253__27_ <= r_n_253__27_;
      r_253__26_ <= r_n_253__26_;
      r_253__25_ <= r_n_253__25_;
      r_253__24_ <= r_n_253__24_;
      r_253__23_ <= r_n_253__23_;
      r_253__22_ <= r_n_253__22_;
      r_253__21_ <= r_n_253__21_;
      r_253__20_ <= r_n_253__20_;
      r_253__19_ <= r_n_253__19_;
      r_253__18_ <= r_n_253__18_;
      r_253__17_ <= r_n_253__17_;
      r_253__16_ <= r_n_253__16_;
      r_253__15_ <= r_n_253__15_;
      r_253__14_ <= r_n_253__14_;
      r_253__13_ <= r_n_253__13_;
      r_253__12_ <= r_n_253__12_;
      r_253__11_ <= r_n_253__11_;
      r_253__10_ <= r_n_253__10_;
      r_253__9_ <= r_n_253__9_;
      r_253__8_ <= r_n_253__8_;
      r_253__7_ <= r_n_253__7_;
      r_253__6_ <= r_n_253__6_;
      r_253__5_ <= r_n_253__5_;
      r_253__4_ <= r_n_253__4_;
      r_253__3_ <= r_n_253__3_;
      r_253__2_ <= r_n_253__2_;
      r_253__1_ <= r_n_253__1_;
      r_253__0_ <= r_n_253__0_;
    end 
    if(N2046) begin
      r_254__31_ <= r_n_254__31_;
      r_254__30_ <= r_n_254__30_;
      r_254__29_ <= r_n_254__29_;
      r_254__28_ <= r_n_254__28_;
      r_254__27_ <= r_n_254__27_;
      r_254__26_ <= r_n_254__26_;
      r_254__25_ <= r_n_254__25_;
      r_254__24_ <= r_n_254__24_;
      r_254__23_ <= r_n_254__23_;
      r_254__22_ <= r_n_254__22_;
      r_254__21_ <= r_n_254__21_;
      r_254__20_ <= r_n_254__20_;
      r_254__19_ <= r_n_254__19_;
      r_254__18_ <= r_n_254__18_;
      r_254__17_ <= r_n_254__17_;
      r_254__16_ <= r_n_254__16_;
      r_254__15_ <= r_n_254__15_;
      r_254__14_ <= r_n_254__14_;
      r_254__13_ <= r_n_254__13_;
      r_254__12_ <= r_n_254__12_;
      r_254__11_ <= r_n_254__11_;
      r_254__10_ <= r_n_254__10_;
      r_254__9_ <= r_n_254__9_;
      r_254__8_ <= r_n_254__8_;
      r_254__7_ <= r_n_254__7_;
      r_254__6_ <= r_n_254__6_;
      r_254__5_ <= r_n_254__5_;
      r_254__4_ <= r_n_254__4_;
      r_254__3_ <= r_n_254__3_;
      r_254__2_ <= r_n_254__2_;
      r_254__1_ <= r_n_254__1_;
      r_254__0_ <= r_n_254__0_;
    end 
    if(N2047) begin
      r_255__31_ <= r_n_255__31_;
      r_255__30_ <= r_n_255__30_;
      r_255__29_ <= r_n_255__29_;
      r_255__28_ <= r_n_255__28_;
      r_255__27_ <= r_n_255__27_;
      r_255__26_ <= r_n_255__26_;
      r_255__25_ <= r_n_255__25_;
      r_255__24_ <= r_n_255__24_;
      r_255__23_ <= r_n_255__23_;
      r_255__22_ <= r_n_255__22_;
      r_255__21_ <= r_n_255__21_;
      r_255__20_ <= r_n_255__20_;
      r_255__19_ <= r_n_255__19_;
      r_255__18_ <= r_n_255__18_;
      r_255__17_ <= r_n_255__17_;
      r_255__16_ <= r_n_255__16_;
      r_255__15_ <= r_n_255__15_;
      r_255__14_ <= r_n_255__14_;
      r_255__13_ <= r_n_255__13_;
      r_255__12_ <= r_n_255__12_;
      r_255__11_ <= r_n_255__11_;
      r_255__10_ <= r_n_255__10_;
      r_255__9_ <= r_n_255__9_;
      r_255__8_ <= r_n_255__8_;
      r_255__7_ <= r_n_255__7_;
      r_255__6_ <= r_n_255__6_;
      r_255__5_ <= r_n_255__5_;
      r_255__4_ <= r_n_255__4_;
      r_255__3_ <= r_n_255__3_;
      r_255__2_ <= r_n_255__2_;
      r_255__1_ <= r_n_255__1_;
      r_255__0_ <= r_n_255__0_;
    end 
  end


endmodule

