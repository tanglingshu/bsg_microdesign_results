

module top
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [8191:0] data_i;
  input [63:0] sel_one_hot_i;
  output [127:0] data_o;

  bsg_mux_one_hot
  wrapper
  (
    .data_i(data_i),
    .sel_one_hot_i(sel_one_hot_i),
    .data_o(data_o)
  );


endmodule



module bsg_mux_one_hot
(
  data_i,
  sel_one_hot_i,
  data_o
);

  input [8191:0] data_i;
  input [63:0] sel_one_hot_i;
  output [127:0] data_o;
  wire [127:0] data_o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022,N1023,N1024,
  N1025,N1026,N1027,N1028,N1029,N1030,N1031,N1032,N1033,N1034,N1035,N1036,N1037,
  N1038,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046,N1047,N1048,N1049,N1050,
  N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062,N1063,N1064,
  N1065,N1066,N1067,N1068,N1069,N1070,N1071,N1072,N1073,N1074,N1075,N1076,N1077,
  N1078,N1079,N1080,N1081,N1082,N1083,N1084,N1085,N1086,N1087,N1088,N1089,N1090,
  N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,N1099,N1100,N1101,N1102,N1103,N1104,
  N1105,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113,N1114,N1115,N1116,N1117,
  N1118,N1119,N1120,N1121,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129,N1130,
  N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,N1139,N1140,N1141,N1142,N1143,N1144,
  N1145,N1146,N1147,N1148,N1149,N1150,N1151,N1152,N1153,N1154,N1155,N1156,N1157,
  N1158,N1159,N1160,N1161,N1162,N1163,N1164,N1165,N1166,N1167,N1168,N1169,N1170,
  N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,N1179,N1180,N1181,N1182,N1183,N1184,
  N1185,N1186,N1187,N1188,N1189,N1190,N1191,N1192,N1193,N1194,N1195,N1196,N1197,
  N1198,N1199,N1200,N1201,N1202,N1203,N1204,N1205,N1206,N1207,N1208,N1209,N1210,
  N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224,
  N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232,N1233,N1234,N1235,N1236,N1237,
  N1238,N1239,N1240,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248,N1249,N1250,
  N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
  N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272,N1273,N1274,N1275,N1276,N1277,
  N1278,N1279,N1280,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288,N1289,N1290,
  N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304,
  N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312,N1313,N1314,N1315,N1316,N1317,
  N1318,N1319,N1320,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328,N1329,N1330,
  N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344,
  N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354,N1355,N1356,N1357,
  N1358,N1359,N1360,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368,N1369,N1370,
  N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384,
  N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392,N1393,N1394,N1395,N1396,N1397,
  N1398,N1399,N1400,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408,N1409,N1410,
  N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424,
  N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434,N1435,N1436,N1437,
  N1438,N1439,N1440,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1450,
  N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,N1463,N1464,
  N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474,N1475,N1476,N1477,
  N1478,N1479,N1480,N1481,N1482,N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,
  N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504,
  N1505,N1506,N1507,N1508,N1509,N1510,N1511,N1512,N1513,N1514,N1515,N1516,N1517,
  N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530,
  N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542,N1543,N1544,
  N1545,N1546,N1547,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557,
  N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568,N1569,N1570,
  N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581,N1582,N1583,N1584,
  N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597,
  N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610,
  N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622,N1623,N1624,
  N1625,N1626,N1627,N1628,N1629,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637,
  N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646,N1647,N1648,N1649,N1650,
  N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1664,
  N1665,N1666,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677,
  N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686,N1687,N1688,N1689,N1690,
  N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702,N1703,N1704,
  N1705,N1706,N1707,N1708,N1709,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717,
  N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728,N1729,N1730,
  N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744,
  N1745,N1746,N1747,N1748,N1749,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757,
  N1758,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1766,N1767,N1768,N1769,N1770,
  N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783,N1784,
  N1785,N1786,N1787,N1788,N1789,N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,
  N1798,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806,N1807,N1808,N1809,N1810,
  N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822,N1823,N1824,
  N1825,N1826,N1827,N1828,N1829,N1830,N1831,N1832,N1833,N1834,N1835,N1836,N1837,
  N1838,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,N1850,
  N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862,N1863,N1864,
  N1865,N1866,N1867,N1868,N1869,N1870,N1871,N1872,N1873,N1874,N1875,N1876,N1877,
  N1878,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886,N1887,N1888,N1889,N1890,
  N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902,N1903,N1904,
  N1905,N1906,N1907,N1908,N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,
  N1918,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926,N1927,N1928,N1929,N1930,
  N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942,N1943,N1944,
  N1945,N1946,N1947,N1948,N1949,N1950,N1951,N1952,N1953,N1954,N1955,N1956,N1957,
  N1958,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966,N1967,N1968,N1969,N1970,
  N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982,N1983,N1984,
  N1985,N1986,N1987,N1988,N1989,N1990,N1991,N1992,N1993,N1994,N1995,N1996,N1997,
  N1998,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006,N2007,N2008,N2009,N2010,
  N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022,N2023,N2024,
  N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2035,N2036,N2037,
  N2038,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046,N2047,N2048,N2049,N2050,
  N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062,N2063,N2064,
  N2065,N2066,N2067,N2068,N2069,N2070,N2071,N2072,N2073,N2074,N2075,N2076,N2077,
  N2078,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086,N2087,N2088,N2089,N2090,
  N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102,N2103,N2104,
  N2105,N2106,N2107,N2108,N2109,N2110,N2111,N2112,N2113,N2114,N2115,N2116,N2117,
  N2118,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126,N2127,N2128,N2129,N2130,
  N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142,N2143,N2144,
  N2145,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,
  N2158,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166,N2167,N2168,N2169,N2170,
  N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184,
  N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196,N2197,
  N2198,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209,N2210,
  N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223,N2224,
  N2225,N2226,N2227,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235,N2236,N2237,
  N2238,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246,N2247,N2248,N2249,N2250,
  N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262,N2263,N2264,
  N2265,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273,N2274,N2275,N2276,N2277,
  N2278,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290,
  N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302,N2303,N2304,
  N2305,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,
  N2318,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,N2329,N2330,
  N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342,N2343,N2344,
  N2345,N2346,N2347,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355,N2356,N2357,
  N2358,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366,N2367,N2368,N2369,N2370,
  N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384,
  N2385,N2386,N2387,N2388,N2389,N2390,N2391,N2392,N2393,N2394,N2395,N2396,N2397,
  N2398,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410,
  N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422,N2423,N2424,
  N2425,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433,N2434,N2435,N2436,N2437,
  N2438,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446,N2447,N2448,N2449,N2450,
  N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462,N2463,N2464,
  N2465,N2466,N2467,N2468,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476,N2477,
  N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487,N2488,N2489,N2490,
  N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504,
  N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512,N2513,N2514,N2515,N2516,N2517,
  N2518,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526,N2527,N2528,N2529,N2530,
  N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542,N2543,N2544,
  N2545,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556,N2557,
  N2558,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566,N2567,N2568,N2569,N2570,
  N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582,N2583,N2584,
  N2585,N2586,N2587,N2588,N2589,N2590,N2591,N2592,N2593,N2594,N2595,N2596,N2597,
  N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606,N2607,N2608,N2609,N2610,
  N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624,
  N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2637,
  N2638,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,N2649,N2650,
  N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662,N2663,N2664,
  N2665,N2666,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,
  N2678,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686,N2687,N2688,N2689,N2690,
  N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2704,
  N2705,N2706,N2707,N2708,N2709,N2710,N2711,N2712,N2713,N2714,N2715,N2716,N2717,
  N2718,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726,N2727,N2728,N2729,N2730,
  N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744,
  N2745,N2746,N2747,N2748,N2749,N2750,N2751,N2752,N2753,N2754,N2755,N2756,N2757,
  N2758,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769,N2770,
  N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783,N2784,
  N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793,N2794,N2795,N2796,N2797,
  N2798,N2799,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2810,
  N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,N2819,N2820,N2821,N2822,N2823,N2824,
  N2825,N2826,N2827,N2828,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836,N2837,
  N2838,N2839,N2840,N2841,N2842,N2843,N2844,N2845,N2846,N2847,N2848,N2849,N2850,
  N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862,N2863,N2864,
  N2865,N2866,N2867,N2868,N2869,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877,
  N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887,N2888,N2889,N2890,
  N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904,
  N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912,N2913,N2914,N2915,N2916,N2917,
  N2918,N2919,N2920,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928,N2929,N2930,
  N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,N2939,N2940,N2941,N2942,N2943,N2944,
  N2945,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954,N2955,N2956,N2957,
  N2958,N2959,N2960,N2961,N2962,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970,
  N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980,N2981,N2982,N2983,N2984,
  N2985,N2986,N2987,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996,N2997,
  N2998,N2999,N3000,N3001,N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,
  N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,N3022,N3023,N3024,
  N3025,N3026,N3027,N3028,N3029,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037,
  N3038,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,
  N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3062,N3063,N3064,
  N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077,
  N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,
  N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,N3102,N3103,N3104,
  N3105,N3106,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114,N3115,N3116,N3117,
  N3118,N3119,N3120,N3121,N3122,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130,
  N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139,N3140,N3141,N3142,N3143,N3144,
  N3145,N3146,N3147,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155,N3156,N3157,
  N3158,N3159,N3160,N3161,N3162,N3163,N3164,N3165,N3166,N3167,N3168,N3169,N3170,
  N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182,N3183,N3184,
  N3185,N3186,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,N3195,N3196,N3197,
  N3198,N3199,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207,N3208,N3209,N3210,
  N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223,N3224,
  N3225,N3226,N3227,N3228,N3229,N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,
  N3238,N3239,N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,N3250,
  N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,N3260,N3261,N3262,N3263,N3264,
  N3265,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,
  N3278,N3279,N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290,
  N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,N3300,N3301,N3302,N3303,N3304,
  N3305,N3306,N3307,N3308,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,
  N3318,N3319,N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,N3330,
  N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341,N3342,N3343,N3344,
  N3345,N3346,N3347,N3348,N3349,N3350,N3351,N3352,N3353,N3354,N3355,N3356,N3357,
  N3358,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367,N3368,N3369,N3370,
  N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383,N3384,
  N3385,N3386,N3387,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,
  N3398,N3399,N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3408,N3409,N3410,
  N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420,N3421,N3422,N3423,N3424,
  N3425,N3426,N3427,N3428,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436,N3437,
  N3438,N3439,N3440,N3441,N3442,N3443,N3444,N3445,N3446,N3447,N3448,N3449,N3450,
  N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460,N3461,N3462,N3463,N3464,
  N3465,N3466,N3467,N3468,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476,N3477,
  N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,N3487,N3488,N3489,N3490,
  N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501,N3502,N3503,N3504,
  N3505,N3506,N3507,N3508,N3509,N3510,N3511,N3512,N3513,N3514,N3515,N3516,N3517,
  N3518,N3519,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527,N3528,N3529,N3530,
  N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543,N3544,
  N3545,N3546,N3547,N3548,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556,N3557,
  N3558,N3559,N3560,N3561,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569,N3570,
  N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,N3579,N3580,N3581,N3582,N3583,N3584,
  N3585,N3586,N3587,N3588,N3589,N3590,N3591,N3592,N3593,N3594,N3595,N3596,N3597,
  N3598,N3599,N3600,N3601,N3602,N3603,N3604,N3605,N3606,N3607,N3608,N3609,N3610,
  N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3620,N3621,N3622,N3623,N3624,
  N3625,N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3636,N3637,
  N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,N3646,N3647,N3648,N3649,N3650,
  N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,N3659,N3660,N3661,N3662,N3663,N3664,
  N3665,N3666,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674,N3675,N3676,N3677,
  N3678,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686,N3687,N3688,N3689,N3690,
  N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699,N3700,N3701,N3702,N3703,N3704,
  N3705,N3706,N3707,N3708,N3709,N3710,N3711,N3712,N3713,N3714,N3715,N3716,N3717,
  N3718,N3719,N3720,N3721,N3722,N3723,N3724,N3725,N3726,N3727,N3728,N3729,N3730,
  N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742,N3743,N3744,
  N3745,N3746,N3747,N3748,N3749,N3750,N3751,N3752,N3753,N3754,N3755,N3756,N3757,
  N3758,N3759,N3760,N3761,N3762,N3763,N3764,N3765,N3766,N3767,N3768,N3769,N3770,
  N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3781,N3782,N3783,N3784,
  N3785,N3786,N3787,N3788,N3789,N3790,N3791,N3792,N3793,N3794,N3795,N3796,N3797,
  N3798,N3799,N3800,N3801,N3802,N3803,N3804,N3805,N3806,N3807,N3808,N3809,N3810,
  N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,N3824,
  N3825,N3826,N3827,N3828,N3829,N3830,N3831,N3832,N3833,N3834,N3835,N3836,N3837,
  N3838,N3839,N3840,N3841,N3842,N3843,N3844,N3845,N3846,N3847,N3848,N3849,N3850,
  N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,N3859,N3860,N3861,N3862,N3863,N3864,
  N3865,N3866,N3867,N3868,N3869,N3870,N3871,N3872,N3873,N3874,N3875,N3876,N3877,
  N3878,N3879,N3880,N3881,N3882,N3883,N3884,N3885,N3886,N3887,N3888,N3889,N3890,
  N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,N3899,N3900,N3901,N3902,N3903,N3904,
  N3905,N3906,N3907,N3908,N3909,N3910,N3911,N3912,N3913,N3914,N3915,N3916,N3917,
  N3918,N3919,N3920,N3921,N3922,N3923,N3924,N3925,N3926,N3927,N3928,N3929,N3930,
  N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,N3939,N3940,N3941,N3942,N3943,N3944,
  N3945,N3946,N3947,N3948,N3949,N3950,N3951,N3952,N3953,N3954,N3955,N3956,N3957,
  N3958,N3959,N3960,N3961,N3962,N3963,N3964,N3965,N3966,N3967,N3968,N3969,N3970,
  N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,N3979,N3980,N3981,N3982,N3983,N3984,
  N3985,N3986,N3987,N3988,N3989,N3990,N3991,N3992,N3993,N3994,N3995,N3996,N3997,
  N3998,N3999,N4000,N4001,N4002,N4003,N4004,N4005,N4006,N4007,N4008,N4009,N4010,
  N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,N4019,N4020,N4021,N4022,N4023,N4024,
  N4025,N4026,N4027,N4028,N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4036,N4037,
  N4038,N4039,N4040,N4041,N4042,N4043,N4044,N4045,N4046,N4047,N4048,N4049,N4050,
  N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,N4059,N4060,N4061,N4062,N4063,N4064,
  N4065,N4066,N4067,N4068,N4069,N4070,N4071,N4072,N4073,N4074,N4075,N4076,N4077,
  N4078,N4079,N4080,N4081,N4082,N4083,N4084,N4085,N4086,N4087,N4088,N4089,N4090,
  N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,N4099,N4100,N4101,N4102,N4103,N4104,
  N4105,N4106,N4107,N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4117,
  N4118,N4119,N4120,N4121,N4122,N4123,N4124,N4125,N4126,N4127,N4128,N4129,N4130,
  N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,N4139,N4140,N4141,N4142,N4143,N4144,
  N4145,N4146,N4147,N4148,N4149,N4150,N4151,N4152,N4153,N4154,N4155,N4156,N4157,
  N4158,N4159,N4160,N4161,N4162,N4163,N4164,N4165,N4166,N4167,N4168,N4169,N4170,
  N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,N4179,N4180,N4181,N4182,N4183,N4184,
  N4185,N4186,N4187,N4188,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,
  N4198,N4199,N4200,N4201,N4202,N4203,N4204,N4205,N4206,N4207,N4208,N4209,N4210,
  N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,N4219,N4220,N4221,N4222,N4223,N4224,
  N4225,N4226,N4227,N4228,N4229,N4230,N4231,N4232,N4233,N4234,N4235,N4236,N4237,
  N4238,N4239,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247,N4248,N4249,N4250,
  N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4259,N4260,N4261,N4262,N4263,N4264,
  N4265,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4273,N4274,N4275,N4276,N4277,
  N4278,N4279,N4280,N4281,N4282,N4283,N4284,N4285,N4286,N4287,N4288,N4289,N4290,
  N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,N4299,N4300,N4301,N4302,N4303,N4304,
  N4305,N4306,N4307,N4308,N4309,N4310,N4311,N4312,N4313,N4314,N4315,N4316,N4317,
  N4318,N4319,N4320,N4321,N4322,N4323,N4324,N4325,N4326,N4327,N4328,N4329,N4330,
  N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,N4339,N4340,N4341,N4342,N4343,N4344,
  N4345,N4346,N4347,N4348,N4349,N4350,N4351,N4352,N4353,N4354,N4355,N4356,N4357,
  N4358,N4359,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367,N4368,N4369,N4370,
  N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,N4379,N4380,N4381,N4382,N4383,N4384,
  N4385,N4386,N4387,N4388,N4389,N4390,N4391,N4392,N4393,N4394,N4395,N4396,N4397,
  N4398,N4399,N4400,N4401,N4402,N4403,N4404,N4405,N4406,N4407,N4408,N4409,N4410,
  N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,N4419,N4420,N4421,N4422,N4423,N4424,
  N4425,N4426,N4427,N4428,N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436,N4437,
  N4438,N4439,N4440,N4441,N4442,N4443,N4444,N4445,N4446,N4447,N4448,N4449,N4450,
  N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,N4459,N4460,N4461,N4462,N4463,N4464,
  N4465,N4466,N4467,N4468,N4469,N4470,N4471,N4472,N4473,N4474,N4475,N4476,N4477,
  N4478,N4479,N4480,N4481,N4482,N4483,N4484,N4485,N4486,N4487,N4488,N4489,N4490,
  N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502,N4503,N4504,
  N4505,N4506,N4507,N4508,N4509,N4510,N4511,N4512,N4513,N4514,N4515,N4516,N4517,
  N4518,N4519,N4520,N4521,N4522,N4523,N4524,N4525,N4526,N4527,N4528,N4529,N4530,
  N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540,N4541,N4542,N4543,N4544,
  N4545,N4546,N4547,N4548,N4549,N4550,N4551,N4552,N4553,N4554,N4555,N4556,N4557,
  N4558,N4559,N4560,N4561,N4562,N4563,N4564,N4565,N4566,N4567,N4568,N4569,N4570,
  N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,N4579,N4580,N4581,N4582,N4583,N4584,
  N4585,N4586,N4587,N4588,N4589,N4590,N4591,N4592,N4593,N4594,N4595,N4596,N4597,
  N4598,N4599,N4600,N4601,N4602,N4603,N4604,N4605,N4606,N4607,N4608,N4609,N4610,
  N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,N4619,N4620,N4621,N4622,N4623,N4624,
  N4625,N4626,N4627,N4628,N4629,N4630,N4631,N4632,N4633,N4634,N4635,N4636,N4637,
  N4638,N4639,N4640,N4641,N4642,N4643,N4644,N4645,N4646,N4647,N4648,N4649,N4650,
  N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,N4659,N4660,N4661,N4662,N4663,N4664,
  N4665,N4666,N4667,N4668,N4669,N4670,N4671,N4672,N4673,N4674,N4675,N4676,N4677,
  N4678,N4679,N4680,N4681,N4682,N4683,N4684,N4685,N4686,N4687,N4688,N4689,N4690,
  N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,N4699,N4700,N4701,N4702,N4703,N4704,
  N4705,N4706,N4707,N4708,N4709,N4710,N4711,N4712,N4713,N4714,N4715,N4716,N4717,
  N4718,N4719,N4720,N4721,N4722,N4723,N4724,N4725,N4726,N4727,N4728,N4729,N4730,
  N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,N4739,N4740,N4741,N4742,N4743,N4744,
  N4745,N4746,N4747,N4748,N4749,N4750,N4751,N4752,N4753,N4754,N4755,N4756,N4757,
  N4758,N4759,N4760,N4761,N4762,N4763,N4764,N4765,N4766,N4767,N4768,N4769,N4770,
  N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,N4779,N4780,N4781,N4782,N4783,N4784,
  N4785,N4786,N4787,N4788,N4789,N4790,N4791,N4792,N4793,N4794,N4795,N4796,N4797,
  N4798,N4799,N4800,N4801,N4802,N4803,N4804,N4805,N4806,N4807,N4808,N4809,N4810,
  N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,N4819,N4820,N4821,N4822,N4823,N4824,
  N4825,N4826,N4827,N4828,N4829,N4830,N4831,N4832,N4833,N4834,N4835,N4836,N4837,
  N4838,N4839,N4840,N4841,N4842,N4843,N4844,N4845,N4846,N4847,N4848,N4849,N4850,
  N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,N4859,N4860,N4861,N4862,N4863,N4864,
  N4865,N4866,N4867,N4868,N4869,N4870,N4871,N4872,N4873,N4874,N4875,N4876,N4877,
  N4878,N4879,N4880,N4881,N4882,N4883,N4884,N4885,N4886,N4887,N4888,N4889,N4890,
  N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4903,N4904,
  N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912,N4913,N4914,N4915,N4916,N4917,
  N4918,N4919,N4920,N4921,N4922,N4923,N4924,N4925,N4926,N4927,N4928,N4929,N4930,
  N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,N4939,N4940,N4941,N4942,N4943,N4944,
  N4945,N4946,N4947,N4948,N4949,N4950,N4951,N4952,N4953,N4954,N4955,N4956,N4957,
  N4958,N4959,N4960,N4961,N4962,N4963,N4964,N4965,N4966,N4967,N4968,N4969,N4970,
  N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,N4979,N4980,N4981,N4982,N4983,N4984,
  N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4992,N4993,N4994,N4995,N4996,N4997,
  N4998,N4999,N5000,N5001,N5002,N5003,N5004,N5005,N5006,N5007,N5008,N5009,N5010,
  N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,N5019,N5020,N5021,N5022,N5023,N5024,
  N5025,N5026,N5027,N5028,N5029,N5030,N5031,N5032,N5033,N5034,N5035,N5036,N5037,
  N5038,N5039,N5040,N5041,N5042,N5043,N5044,N5045,N5046,N5047,N5048,N5049,N5050,
  N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060,N5061,N5062,N5063,N5064,
  N5065,N5066,N5067,N5068,N5069,N5070,N5071,N5072,N5073,N5074,N5075,N5076,N5077,
  N5078,N5079,N5080,N5081,N5082,N5083,N5084,N5085,N5086,N5087,N5088,N5089,N5090,
  N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,N5099,N5100,N5101,N5102,N5103,N5104,
  N5105,N5106,N5107,N5108,N5109,N5110,N5111,N5112,N5113,N5114,N5115,N5116,N5117,
  N5118,N5119,N5120,N5121,N5122,N5123,N5124,N5125,N5126,N5127,N5128,N5129,N5130,
  N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,N5139,N5140,N5141,N5142,N5143,N5144,
  N5145,N5146,N5147,N5148,N5149,N5150,N5151,N5152,N5153,N5154,N5155,N5156,N5157,
  N5158,N5159,N5160,N5161,N5162,N5163,N5164,N5165,N5166,N5167,N5168,N5169,N5170,
  N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,N5179,N5180,N5181,N5182,N5183,N5184,
  N5185,N5186,N5187,N5188,N5189,N5190,N5191,N5192,N5193,N5194,N5195,N5196,N5197,
  N5198,N5199,N5200,N5201,N5202,N5203,N5204,N5205,N5206,N5207,N5208,N5209,N5210,
  N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,N5219,N5220,N5221,N5222,N5223,N5224,
  N5225,N5226,N5227,N5228,N5229,N5230,N5231,N5232,N5233,N5234,N5235,N5236,N5237,
  N5238,N5239,N5240,N5241,N5242,N5243,N5244,N5245,N5246,N5247,N5248,N5249,N5250,
  N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,N5259,N5260,N5261,N5262,N5263,N5264,
  N5265,N5266,N5267,N5268,N5269,N5270,N5271,N5272,N5273,N5274,N5275,N5276,N5277,
  N5278,N5279,N5280,N5281,N5282,N5283,N5284,N5285,N5286,N5287,N5288,N5289,N5290,
  N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,N5299,N5300,N5301,N5302,N5303,N5304,
  N5305,N5306,N5307,N5308,N5309,N5310,N5311,N5312,N5313,N5314,N5315,N5316,N5317,
  N5318,N5319,N5320,N5321,N5322,N5323,N5324,N5325,N5326,N5327,N5328,N5329,N5330,
  N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,N5339,N5340,N5341,N5342,N5343,N5344,
  N5345,N5346,N5347,N5348,N5349,N5350,N5351,N5352,N5353,N5354,N5355,N5356,N5357,
  N5358,N5359,N5360,N5361,N5362,N5363,N5364,N5365,N5366,N5367,N5368,N5369,N5370,
  N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,N5379,N5380,N5381,N5382,N5383,N5384,
  N5385,N5386,N5387,N5388,N5389,N5390,N5391,N5392,N5393,N5394,N5395,N5396,N5397,
  N5398,N5399,N5400,N5401,N5402,N5403,N5404,N5405,N5406,N5407,N5408,N5409,N5410,
  N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,N5419,N5420,N5421,N5422,N5423,N5424,
  N5425,N5426,N5427,N5428,N5429,N5430,N5431,N5432,N5433,N5434,N5435,N5436,N5437,
  N5438,N5439,N5440,N5441,N5442,N5443,N5444,N5445,N5446,N5447,N5448,N5449,N5450,
  N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,N5459,N5460,N5461,N5462,N5463,N5464,
  N5465,N5466,N5467,N5468,N5469,N5470,N5471,N5472,N5473,N5474,N5475,N5476,N5477,
  N5478,N5479,N5480,N5481,N5482,N5483,N5484,N5485,N5486,N5487,N5488,N5489,N5490,
  N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,N5499,N5500,N5501,N5502,N5503,N5504,
  N5505,N5506,N5507,N5508,N5509,N5510,N5511,N5512,N5513,N5514,N5515,N5516,N5517,
  N5518,N5519,N5520,N5521,N5522,N5523,N5524,N5525,N5526,N5527,N5528,N5529,N5530,
  N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,N5539,N5540,N5541,N5542,N5543,N5544,
  N5545,N5546,N5547,N5548,N5549,N5550,N5551,N5552,N5553,N5554,N5555,N5556,N5557,
  N5558,N5559,N5560,N5561,N5562,N5563,N5564,N5565,N5566,N5567,N5568,N5569,N5570,
  N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,N5579,N5580,N5581,N5582,N5583,N5584,
  N5585,N5586,N5587,N5588,N5589,N5590,N5591,N5592,N5593,N5594,N5595,N5596,N5597,
  N5598,N5599,N5600,N5601,N5602,N5603,N5604,N5605,N5606,N5607,N5608,N5609,N5610,
  N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,N5619,N5620,N5621,N5622,N5623,N5624,
  N5625,N5626,N5627,N5628,N5629,N5630,N5631,N5632,N5633,N5634,N5635,N5636,N5637,
  N5638,N5639,N5640,N5641,N5642,N5643,N5644,N5645,N5646,N5647,N5648,N5649,N5650,
  N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,N5659,N5660,N5661,N5662,N5663,N5664,
  N5665,N5666,N5667,N5668,N5669,N5670,N5671,N5672,N5673,N5674,N5675,N5676,N5677,
  N5678,N5679,N5680,N5681,N5682,N5683,N5684,N5685,N5686,N5687,N5688,N5689,N5690,
  N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,N5699,N5700,N5701,N5702,N5703,N5704,
  N5705,N5706,N5707,N5708,N5709,N5710,N5711,N5712,N5713,N5714,N5715,N5716,N5717,
  N5718,N5719,N5720,N5721,N5722,N5723,N5724,N5725,N5726,N5727,N5728,N5729,N5730,
  N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,N5739,N5740,N5741,N5742,N5743,N5744,
  N5745,N5746,N5747,N5748,N5749,N5750,N5751,N5752,N5753,N5754,N5755,N5756,N5757,
  N5758,N5759,N5760,N5761,N5762,N5763,N5764,N5765,N5766,N5767,N5768,N5769,N5770,
  N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,N5779,N5780,N5781,N5782,N5783,N5784,
  N5785,N5786,N5787,N5788,N5789,N5790,N5791,N5792,N5793,N5794,N5795,N5796,N5797,
  N5798,N5799,N5800,N5801,N5802,N5803,N5804,N5805,N5806,N5807,N5808,N5809,N5810,
  N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,N5819,N5820,N5821,N5822,N5823,N5824,
  N5825,N5826,N5827,N5828,N5829,N5830,N5831,N5832,N5833,N5834,N5835,N5836,N5837,
  N5838,N5839,N5840,N5841,N5842,N5843,N5844,N5845,N5846,N5847,N5848,N5849,N5850,
  N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,N5859,N5860,N5861,N5862,N5863,N5864,
  N5865,N5866,N5867,N5868,N5869,N5870,N5871,N5872,N5873,N5874,N5875,N5876,N5877,
  N5878,N5879,N5880,N5881,N5882,N5883,N5884,N5885,N5886,N5887,N5888,N5889,N5890,
  N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,N5899,N5900,N5901,N5902,N5903,N5904,
  N5905,N5906,N5907,N5908,N5909,N5910,N5911,N5912,N5913,N5914,N5915,N5916,N5917,
  N5918,N5919,N5920,N5921,N5922,N5923,N5924,N5925,N5926,N5927,N5928,N5929,N5930,
  N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,N5939,N5940,N5941,N5942,N5943,N5944,
  N5945,N5946,N5947,N5948,N5949,N5950,N5951,N5952,N5953,N5954,N5955,N5956,N5957,
  N5958,N5959,N5960,N5961,N5962,N5963,N5964,N5965,N5966,N5967,N5968,N5969,N5970,
  N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,N5979,N5980,N5981,N5982,N5983,N5984,
  N5985,N5986,N5987,N5988,N5989,N5990,N5991,N5992,N5993,N5994,N5995,N5996,N5997,
  N5998,N5999,N6000,N6001,N6002,N6003,N6004,N6005,N6006,N6007,N6008,N6009,N6010,
  N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,N6019,N6020,N6021,N6022,N6023,N6024,
  N6025,N6026,N6027,N6028,N6029,N6030,N6031,N6032,N6033,N6034,N6035,N6036,N6037,
  N6038,N6039,N6040,N6041,N6042,N6043,N6044,N6045,N6046,N6047,N6048,N6049,N6050,
  N6051,N6052,N6053,N6054,N6055,N6056,N6057,N6058,N6059,N6060,N6061,N6062,N6063,N6064,
  N6065,N6066,N6067,N6068,N6069,N6070,N6071,N6072,N6073,N6074,N6075,N6076,N6077,
  N6078,N6079,N6080,N6081,N6082,N6083,N6084,N6085,N6086,N6087,N6088,N6089,N6090,
  N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,N6099,N6100,N6101,N6102,N6103,N6104,
  N6105,N6106,N6107,N6108,N6109,N6110,N6111,N6112,N6113,N6114,N6115,N6116,N6117,
  N6118,N6119,N6120,N6121,N6122,N6123,N6124,N6125,N6126,N6127,N6128,N6129,N6130,
  N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,N6139,N6140,N6141,N6142,N6143,N6144,
  N6145,N6146,N6147,N6148,N6149,N6150,N6151,N6152,N6153,N6154,N6155,N6156,N6157,
  N6158,N6159,N6160,N6161,N6162,N6163,N6164,N6165,N6166,N6167,N6168,N6169,N6170,
  N6171,N6172,N6173,N6174,N6175,N6176,N6177,N6178,N6179,N6180,N6181,N6182,N6183,N6184,
  N6185,N6186,N6187,N6188,N6189,N6190,N6191,N6192,N6193,N6194,N6195,N6196,N6197,
  N6198,N6199,N6200,N6201,N6202,N6203,N6204,N6205,N6206,N6207,N6208,N6209,N6210,
  N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218,N6219,N6220,N6221,N6222,N6223,N6224,
  N6225,N6226,N6227,N6228,N6229,N6230,N6231,N6232,N6233,N6234,N6235,N6236,N6237,
  N6238,N6239,N6240,N6241,N6242,N6243,N6244,N6245,N6246,N6247,N6248,N6249,N6250,
  N6251,N6252,N6253,N6254,N6255,N6256,N6257,N6258,N6259,N6260,N6261,N6262,N6263,N6264,
  N6265,N6266,N6267,N6268,N6269,N6270,N6271,N6272,N6273,N6274,N6275,N6276,N6277,
  N6278,N6279,N6280,N6281,N6282,N6283,N6284,N6285,N6286,N6287,N6288,N6289,N6290,
  N6291,N6292,N6293,N6294,N6295,N6296,N6297,N6298,N6299,N6300,N6301,N6302,N6303,N6304,
  N6305,N6306,N6307,N6308,N6309,N6310,N6311,N6312,N6313,N6314,N6315,N6316,N6317,
  N6318,N6319,N6320,N6321,N6322,N6323,N6324,N6325,N6326,N6327,N6328,N6329,N6330,
  N6331,N6332,N6333,N6334,N6335,N6336,N6337,N6338,N6339,N6340,N6341,N6342,N6343,N6344,
  N6345,N6346,N6347,N6348,N6349,N6350,N6351,N6352,N6353,N6354,N6355,N6356,N6357,
  N6358,N6359,N6360,N6361,N6362,N6363,N6364,N6365,N6366,N6367,N6368,N6369,N6370,
  N6371,N6372,N6373,N6374,N6375,N6376,N6377,N6378,N6379,N6380,N6381,N6382,N6383,N6384,
  N6385,N6386,N6387,N6388,N6389,N6390,N6391,N6392,N6393,N6394,N6395,N6396,N6397,
  N6398,N6399,N6400,N6401,N6402,N6403,N6404,N6405,N6406,N6407,N6408,N6409,N6410,
  N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6418,N6419,N6420,N6421,N6422,N6423,N6424,
  N6425,N6426,N6427,N6428,N6429,N6430,N6431,N6432,N6433,N6434,N6435,N6436,N6437,
  N6438,N6439,N6440,N6441,N6442,N6443,N6444,N6445,N6446,N6447,N6448,N6449,N6450,
  N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458,N6459,N6460,N6461,N6462,N6463,N6464,
  N6465,N6466,N6467,N6468,N6469,N6470,N6471,N6472,N6473,N6474,N6475,N6476,N6477,
  N6478,N6479,N6480,N6481,N6482,N6483,N6484,N6485,N6486,N6487,N6488,N6489,N6490,
  N6491,N6492,N6493,N6494,N6495,N6496,N6497,N6498,N6499,N6500,N6501,N6502,N6503,N6504,
  N6505,N6506,N6507,N6508,N6509,N6510,N6511,N6512,N6513,N6514,N6515,N6516,N6517,
  N6518,N6519,N6520,N6521,N6522,N6523,N6524,N6525,N6526,N6527,N6528,N6529,N6530,
  N6531,N6532,N6533,N6534,N6535,N6536,N6537,N6538,N6539,N6540,N6541,N6542,N6543,N6544,
  N6545,N6546,N6547,N6548,N6549,N6550,N6551,N6552,N6553,N6554,N6555,N6556,N6557,
  N6558,N6559,N6560,N6561,N6562,N6563,N6564,N6565,N6566,N6567,N6568,N6569,N6570,
  N6571,N6572,N6573,N6574,N6575,N6576,N6577,N6578,N6579,N6580,N6581,N6582,N6583,N6584,
  N6585,N6586,N6587,N6588,N6589,N6590,N6591,N6592,N6593,N6594,N6595,N6596,N6597,
  N6598,N6599,N6600,N6601,N6602,N6603,N6604,N6605,N6606,N6607,N6608,N6609,N6610,
  N6611,N6612,N6613,N6614,N6615,N6616,N6617,N6618,N6619,N6620,N6621,N6622,N6623,N6624,
  N6625,N6626,N6627,N6628,N6629,N6630,N6631,N6632,N6633,N6634,N6635,N6636,N6637,
  N6638,N6639,N6640,N6641,N6642,N6643,N6644,N6645,N6646,N6647,N6648,N6649,N6650,
  N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,N6659,N6660,N6661,N6662,N6663,N6664,
  N6665,N6666,N6667,N6668,N6669,N6670,N6671,N6672,N6673,N6674,N6675,N6676,N6677,
  N6678,N6679,N6680,N6681,N6682,N6683,N6684,N6685,N6686,N6687,N6688,N6689,N6690,
  N6691,N6692,N6693,N6694,N6695,N6696,N6697,N6698,N6699,N6700,N6701,N6702,N6703,N6704,
  N6705,N6706,N6707,N6708,N6709,N6710,N6711,N6712,N6713,N6714,N6715,N6716,N6717,
  N6718,N6719,N6720,N6721,N6722,N6723,N6724,N6725,N6726,N6727,N6728,N6729,N6730,
  N6731,N6732,N6733,N6734,N6735,N6736,N6737,N6738,N6739,N6740,N6741,N6742,N6743,N6744,
  N6745,N6746,N6747,N6748,N6749,N6750,N6751,N6752,N6753,N6754,N6755,N6756,N6757,
  N6758,N6759,N6760,N6761,N6762,N6763,N6764,N6765,N6766,N6767,N6768,N6769,N6770,
  N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,N6779,N6780,N6781,N6782,N6783,N6784,
  N6785,N6786,N6787,N6788,N6789,N6790,N6791,N6792,N6793,N6794,N6795,N6796,N6797,
  N6798,N6799,N6800,N6801,N6802,N6803,N6804,N6805,N6806,N6807,N6808,N6809,N6810,
  N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6818,N6819,N6820,N6821,N6822,N6823,N6824,
  N6825,N6826,N6827,N6828,N6829,N6830,N6831,N6832,N6833,N6834,N6835,N6836,N6837,
  N6838,N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6846,N6847,N6848,N6849,N6850,
  N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,N6859,N6860,N6861,N6862,N6863,N6864,
  N6865,N6866,N6867,N6868,N6869,N6870,N6871,N6872,N6873,N6874,N6875,N6876,N6877,
  N6878,N6879,N6880,N6881,N6882,N6883,N6884,N6885,N6886,N6887,N6888,N6889,N6890,
  N6891,N6892,N6893,N6894,N6895,N6896,N6897,N6898,N6899,N6900,N6901,N6902,N6903,N6904,
  N6905,N6906,N6907,N6908,N6909,N6910,N6911,N6912,N6913,N6914,N6915,N6916,N6917,
  N6918,N6919,N6920,N6921,N6922,N6923,N6924,N6925,N6926,N6927,N6928,N6929,N6930,
  N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6938,N6939,N6940,N6941,N6942,N6943,N6944,
  N6945,N6946,N6947,N6948,N6949,N6950,N6951,N6952,N6953,N6954,N6955,N6956,N6957,
  N6958,N6959,N6960,N6961,N6962,N6963,N6964,N6965,N6966,N6967,N6968,N6969,N6970,
  N6971,N6972,N6973,N6974,N6975,N6976,N6977,N6978,N6979,N6980,N6981,N6982,N6983,N6984,
  N6985,N6986,N6987,N6988,N6989,N6990,N6991,N6992,N6993,N6994,N6995,N6996,N6997,
  N6998,N6999,N7000,N7001,N7002,N7003,N7004,N7005,N7006,N7007,N7008,N7009,N7010,
  N7011,N7012,N7013,N7014,N7015,N7016,N7017,N7018,N7019,N7020,N7021,N7022,N7023,N7024,
  N7025,N7026,N7027,N7028,N7029,N7030,N7031,N7032,N7033,N7034,N7035,N7036,N7037,
  N7038,N7039,N7040,N7041,N7042,N7043,N7044,N7045,N7046,N7047,N7048,N7049,N7050,
  N7051,N7052,N7053,N7054,N7055,N7056,N7057,N7058,N7059,N7060,N7061,N7062,N7063,N7064,
  N7065,N7066,N7067,N7068,N7069,N7070,N7071,N7072,N7073,N7074,N7075,N7076,N7077,
  N7078,N7079,N7080,N7081,N7082,N7083,N7084,N7085,N7086,N7087,N7088,N7089,N7090,
  N7091,N7092,N7093,N7094,N7095,N7096,N7097,N7098,N7099,N7100,N7101,N7102,N7103,N7104,
  N7105,N7106,N7107,N7108,N7109,N7110,N7111,N7112,N7113,N7114,N7115,N7116,N7117,
  N7118,N7119,N7120,N7121,N7122,N7123,N7124,N7125,N7126,N7127,N7128,N7129,N7130,
  N7131,N7132,N7133,N7134,N7135,N7136,N7137,N7138,N7139,N7140,N7141,N7142,N7143,N7144,
  N7145,N7146,N7147,N7148,N7149,N7150,N7151,N7152,N7153,N7154,N7155,N7156,N7157,
  N7158,N7159,N7160,N7161,N7162,N7163,N7164,N7165,N7166,N7167,N7168,N7169,N7170,
  N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,N7179,N7180,N7181,N7182,N7183,N7184,
  N7185,N7186,N7187,N7188,N7189,N7190,N7191,N7192,N7193,N7194,N7195,N7196,N7197,
  N7198,N7199,N7200,N7201,N7202,N7203,N7204,N7205,N7206,N7207,N7208,N7209,N7210,
  N7211,N7212,N7213,N7214,N7215,N7216,N7217,N7218,N7219,N7220,N7221,N7222,N7223,N7224,
  N7225,N7226,N7227,N7228,N7229,N7230,N7231,N7232,N7233,N7234,N7235,N7236,N7237,
  N7238,N7239,N7240,N7241,N7242,N7243,N7244,N7245,N7246,N7247,N7248,N7249,N7250,
  N7251,N7252,N7253,N7254,N7255,N7256,N7257,N7258,N7259,N7260,N7261,N7262,N7263,N7264,
  N7265,N7266,N7267,N7268,N7269,N7270,N7271,N7272,N7273,N7274,N7275,N7276,N7277,
  N7278,N7279,N7280,N7281,N7282,N7283,N7284,N7285,N7286,N7287,N7288,N7289,N7290,
  N7291,N7292,N7293,N7294,N7295,N7296,N7297,N7298,N7299,N7300,N7301,N7302,N7303,N7304,
  N7305,N7306,N7307,N7308,N7309,N7310,N7311,N7312,N7313,N7314,N7315,N7316,N7317,
  N7318,N7319,N7320,N7321,N7322,N7323,N7324,N7325,N7326,N7327,N7328,N7329,N7330,
  N7331,N7332,N7333,N7334,N7335,N7336,N7337,N7338,N7339,N7340,N7341,N7342,N7343,N7344,
  N7345,N7346,N7347,N7348,N7349,N7350,N7351,N7352,N7353,N7354,N7355,N7356,N7357,
  N7358,N7359,N7360,N7361,N7362,N7363,N7364,N7365,N7366,N7367,N7368,N7369,N7370,
  N7371,N7372,N7373,N7374,N7375,N7376,N7377,N7378,N7379,N7380,N7381,N7382,N7383,N7384,
  N7385,N7386,N7387,N7388,N7389,N7390,N7391,N7392,N7393,N7394,N7395,N7396,N7397,
  N7398,N7399,N7400,N7401,N7402,N7403,N7404,N7405,N7406,N7407,N7408,N7409,N7410,
  N7411,N7412,N7413,N7414,N7415,N7416,N7417,N7418,N7419,N7420,N7421,N7422,N7423,N7424,
  N7425,N7426,N7427,N7428,N7429,N7430,N7431,N7432,N7433,N7434,N7435,N7436,N7437,
  N7438,N7439,N7440,N7441,N7442,N7443,N7444,N7445,N7446,N7447,N7448,N7449,N7450,
  N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,N7459,N7460,N7461,N7462,N7463,N7464,
  N7465,N7466,N7467,N7468,N7469,N7470,N7471,N7472,N7473,N7474,N7475,N7476,N7477,
  N7478,N7479,N7480,N7481,N7482,N7483,N7484,N7485,N7486,N7487,N7488,N7489,N7490,
  N7491,N7492,N7493,N7494,N7495,N7496,N7497,N7498,N7499,N7500,N7501,N7502,N7503,N7504,
  N7505,N7506,N7507,N7508,N7509,N7510,N7511,N7512,N7513,N7514,N7515,N7516,N7517,
  N7518,N7519,N7520,N7521,N7522,N7523,N7524,N7525,N7526,N7527,N7528,N7529,N7530,
  N7531,N7532,N7533,N7534,N7535,N7536,N7537,N7538,N7539,N7540,N7541,N7542,N7543,N7544,
  N7545,N7546,N7547,N7548,N7549,N7550,N7551,N7552,N7553,N7554,N7555,N7556,N7557,
  N7558,N7559,N7560,N7561,N7562,N7563,N7564,N7565,N7566,N7567,N7568,N7569,N7570,
  N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578,N7579,N7580,N7581,N7582,N7583,N7584,
  N7585,N7586,N7587,N7588,N7589,N7590,N7591,N7592,N7593,N7594,N7595,N7596,N7597,
  N7598,N7599,N7600,N7601,N7602,N7603,N7604,N7605,N7606,N7607,N7608,N7609,N7610,
  N7611,N7612,N7613,N7614,N7615,N7616,N7617,N7618,N7619,N7620,N7621,N7622,N7623,N7624,
  N7625,N7626,N7627,N7628,N7629,N7630,N7631,N7632,N7633,N7634,N7635,N7636,N7637,
  N7638,N7639,N7640,N7641,N7642,N7643,N7644,N7645,N7646,N7647,N7648,N7649,N7650,
  N7651,N7652,N7653,N7654,N7655,N7656,N7657,N7658,N7659,N7660,N7661,N7662,N7663,N7664,
  N7665,N7666,N7667,N7668,N7669,N7670,N7671,N7672,N7673,N7674,N7675,N7676,N7677,
  N7678,N7679,N7680,N7681,N7682,N7683,N7684,N7685,N7686,N7687,N7688,N7689,N7690,
  N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698,N7699,N7700,N7701,N7702,N7703,N7704,
  N7705,N7706,N7707,N7708,N7709,N7710,N7711,N7712,N7713,N7714,N7715,N7716,N7717,
  N7718,N7719,N7720,N7721,N7722,N7723,N7724,N7725,N7726,N7727,N7728,N7729,N7730,
  N7731,N7732,N7733,N7734,N7735,N7736,N7737,N7738,N7739,N7740,N7741,N7742,N7743,N7744,
  N7745,N7746,N7747,N7748,N7749,N7750,N7751,N7752,N7753,N7754,N7755,N7756,N7757,
  N7758,N7759,N7760,N7761,N7762,N7763,N7764,N7765,N7766,N7767,N7768,N7769,N7770,
  N7771,N7772,N7773,N7774,N7775,N7776,N7777,N7778,N7779,N7780,N7781,N7782,N7783,N7784,
  N7785,N7786,N7787,N7788,N7789,N7790,N7791,N7792,N7793,N7794,N7795,N7796,N7797,
  N7798,N7799,N7800,N7801,N7802,N7803,N7804,N7805,N7806,N7807,N7808,N7809,N7810,
  N7811,N7812,N7813,N7814,N7815,N7816,N7817,N7818,N7819,N7820,N7821,N7822,N7823,N7824,
  N7825,N7826,N7827,N7828,N7829,N7830,N7831,N7832,N7833,N7834,N7835,N7836,N7837,
  N7838,N7839,N7840,N7841,N7842,N7843,N7844,N7845,N7846,N7847,N7848,N7849,N7850,
  N7851,N7852,N7853,N7854,N7855,N7856,N7857,N7858,N7859,N7860,N7861,N7862,N7863,N7864,
  N7865,N7866,N7867,N7868,N7869,N7870,N7871,N7872,N7873,N7874,N7875,N7876,N7877,
  N7878,N7879,N7880,N7881,N7882,N7883,N7884,N7885,N7886,N7887,N7888,N7889,N7890,
  N7891,N7892,N7893,N7894,N7895,N7896,N7897,N7898,N7899,N7900,N7901,N7902,N7903,N7904,
  N7905,N7906,N7907,N7908,N7909,N7910,N7911,N7912,N7913,N7914,N7915,N7916,N7917,
  N7918,N7919,N7920,N7921,N7922,N7923,N7924,N7925,N7926,N7927,N7928,N7929,N7930,
  N7931,N7932,N7933,N7934,N7935;
  wire [8191:0] data_masked;
  assign data_masked[127] = data_i[127] & sel_one_hot_i[0];
  assign data_masked[126] = data_i[126] & sel_one_hot_i[0];
  assign data_masked[125] = data_i[125] & sel_one_hot_i[0];
  assign data_masked[124] = data_i[124] & sel_one_hot_i[0];
  assign data_masked[123] = data_i[123] & sel_one_hot_i[0];
  assign data_masked[122] = data_i[122] & sel_one_hot_i[0];
  assign data_masked[121] = data_i[121] & sel_one_hot_i[0];
  assign data_masked[120] = data_i[120] & sel_one_hot_i[0];
  assign data_masked[119] = data_i[119] & sel_one_hot_i[0];
  assign data_masked[118] = data_i[118] & sel_one_hot_i[0];
  assign data_masked[117] = data_i[117] & sel_one_hot_i[0];
  assign data_masked[116] = data_i[116] & sel_one_hot_i[0];
  assign data_masked[115] = data_i[115] & sel_one_hot_i[0];
  assign data_masked[114] = data_i[114] & sel_one_hot_i[0];
  assign data_masked[113] = data_i[113] & sel_one_hot_i[0];
  assign data_masked[112] = data_i[112] & sel_one_hot_i[0];
  assign data_masked[111] = data_i[111] & sel_one_hot_i[0];
  assign data_masked[110] = data_i[110] & sel_one_hot_i[0];
  assign data_masked[109] = data_i[109] & sel_one_hot_i[0];
  assign data_masked[108] = data_i[108] & sel_one_hot_i[0];
  assign data_masked[107] = data_i[107] & sel_one_hot_i[0];
  assign data_masked[106] = data_i[106] & sel_one_hot_i[0];
  assign data_masked[105] = data_i[105] & sel_one_hot_i[0];
  assign data_masked[104] = data_i[104] & sel_one_hot_i[0];
  assign data_masked[103] = data_i[103] & sel_one_hot_i[0];
  assign data_masked[102] = data_i[102] & sel_one_hot_i[0];
  assign data_masked[101] = data_i[101] & sel_one_hot_i[0];
  assign data_masked[100] = data_i[100] & sel_one_hot_i[0];
  assign data_masked[99] = data_i[99] & sel_one_hot_i[0];
  assign data_masked[98] = data_i[98] & sel_one_hot_i[0];
  assign data_masked[97] = data_i[97] & sel_one_hot_i[0];
  assign data_masked[96] = data_i[96] & sel_one_hot_i[0];
  assign data_masked[95] = data_i[95] & sel_one_hot_i[0];
  assign data_masked[94] = data_i[94] & sel_one_hot_i[0];
  assign data_masked[93] = data_i[93] & sel_one_hot_i[0];
  assign data_masked[92] = data_i[92] & sel_one_hot_i[0];
  assign data_masked[91] = data_i[91] & sel_one_hot_i[0];
  assign data_masked[90] = data_i[90] & sel_one_hot_i[0];
  assign data_masked[89] = data_i[89] & sel_one_hot_i[0];
  assign data_masked[88] = data_i[88] & sel_one_hot_i[0];
  assign data_masked[87] = data_i[87] & sel_one_hot_i[0];
  assign data_masked[86] = data_i[86] & sel_one_hot_i[0];
  assign data_masked[85] = data_i[85] & sel_one_hot_i[0];
  assign data_masked[84] = data_i[84] & sel_one_hot_i[0];
  assign data_masked[83] = data_i[83] & sel_one_hot_i[0];
  assign data_masked[82] = data_i[82] & sel_one_hot_i[0];
  assign data_masked[81] = data_i[81] & sel_one_hot_i[0];
  assign data_masked[80] = data_i[80] & sel_one_hot_i[0];
  assign data_masked[79] = data_i[79] & sel_one_hot_i[0];
  assign data_masked[78] = data_i[78] & sel_one_hot_i[0];
  assign data_masked[77] = data_i[77] & sel_one_hot_i[0];
  assign data_masked[76] = data_i[76] & sel_one_hot_i[0];
  assign data_masked[75] = data_i[75] & sel_one_hot_i[0];
  assign data_masked[74] = data_i[74] & sel_one_hot_i[0];
  assign data_masked[73] = data_i[73] & sel_one_hot_i[0];
  assign data_masked[72] = data_i[72] & sel_one_hot_i[0];
  assign data_masked[71] = data_i[71] & sel_one_hot_i[0];
  assign data_masked[70] = data_i[70] & sel_one_hot_i[0];
  assign data_masked[69] = data_i[69] & sel_one_hot_i[0];
  assign data_masked[68] = data_i[68] & sel_one_hot_i[0];
  assign data_masked[67] = data_i[67] & sel_one_hot_i[0];
  assign data_masked[66] = data_i[66] & sel_one_hot_i[0];
  assign data_masked[65] = data_i[65] & sel_one_hot_i[0];
  assign data_masked[64] = data_i[64] & sel_one_hot_i[0];
  assign data_masked[63] = data_i[63] & sel_one_hot_i[0];
  assign data_masked[62] = data_i[62] & sel_one_hot_i[0];
  assign data_masked[61] = data_i[61] & sel_one_hot_i[0];
  assign data_masked[60] = data_i[60] & sel_one_hot_i[0];
  assign data_masked[59] = data_i[59] & sel_one_hot_i[0];
  assign data_masked[58] = data_i[58] & sel_one_hot_i[0];
  assign data_masked[57] = data_i[57] & sel_one_hot_i[0];
  assign data_masked[56] = data_i[56] & sel_one_hot_i[0];
  assign data_masked[55] = data_i[55] & sel_one_hot_i[0];
  assign data_masked[54] = data_i[54] & sel_one_hot_i[0];
  assign data_masked[53] = data_i[53] & sel_one_hot_i[0];
  assign data_masked[52] = data_i[52] & sel_one_hot_i[0];
  assign data_masked[51] = data_i[51] & sel_one_hot_i[0];
  assign data_masked[50] = data_i[50] & sel_one_hot_i[0];
  assign data_masked[49] = data_i[49] & sel_one_hot_i[0];
  assign data_masked[48] = data_i[48] & sel_one_hot_i[0];
  assign data_masked[47] = data_i[47] & sel_one_hot_i[0];
  assign data_masked[46] = data_i[46] & sel_one_hot_i[0];
  assign data_masked[45] = data_i[45] & sel_one_hot_i[0];
  assign data_masked[44] = data_i[44] & sel_one_hot_i[0];
  assign data_masked[43] = data_i[43] & sel_one_hot_i[0];
  assign data_masked[42] = data_i[42] & sel_one_hot_i[0];
  assign data_masked[41] = data_i[41] & sel_one_hot_i[0];
  assign data_masked[40] = data_i[40] & sel_one_hot_i[0];
  assign data_masked[39] = data_i[39] & sel_one_hot_i[0];
  assign data_masked[38] = data_i[38] & sel_one_hot_i[0];
  assign data_masked[37] = data_i[37] & sel_one_hot_i[0];
  assign data_masked[36] = data_i[36] & sel_one_hot_i[0];
  assign data_masked[35] = data_i[35] & sel_one_hot_i[0];
  assign data_masked[34] = data_i[34] & sel_one_hot_i[0];
  assign data_masked[33] = data_i[33] & sel_one_hot_i[0];
  assign data_masked[32] = data_i[32] & sel_one_hot_i[0];
  assign data_masked[31] = data_i[31] & sel_one_hot_i[0];
  assign data_masked[30] = data_i[30] & sel_one_hot_i[0];
  assign data_masked[29] = data_i[29] & sel_one_hot_i[0];
  assign data_masked[28] = data_i[28] & sel_one_hot_i[0];
  assign data_masked[27] = data_i[27] & sel_one_hot_i[0];
  assign data_masked[26] = data_i[26] & sel_one_hot_i[0];
  assign data_masked[25] = data_i[25] & sel_one_hot_i[0];
  assign data_masked[24] = data_i[24] & sel_one_hot_i[0];
  assign data_masked[23] = data_i[23] & sel_one_hot_i[0];
  assign data_masked[22] = data_i[22] & sel_one_hot_i[0];
  assign data_masked[21] = data_i[21] & sel_one_hot_i[0];
  assign data_masked[20] = data_i[20] & sel_one_hot_i[0];
  assign data_masked[19] = data_i[19] & sel_one_hot_i[0];
  assign data_masked[18] = data_i[18] & sel_one_hot_i[0];
  assign data_masked[17] = data_i[17] & sel_one_hot_i[0];
  assign data_masked[16] = data_i[16] & sel_one_hot_i[0];
  assign data_masked[15] = data_i[15] & sel_one_hot_i[0];
  assign data_masked[14] = data_i[14] & sel_one_hot_i[0];
  assign data_masked[13] = data_i[13] & sel_one_hot_i[0];
  assign data_masked[12] = data_i[12] & sel_one_hot_i[0];
  assign data_masked[11] = data_i[11] & sel_one_hot_i[0];
  assign data_masked[10] = data_i[10] & sel_one_hot_i[0];
  assign data_masked[9] = data_i[9] & sel_one_hot_i[0];
  assign data_masked[8] = data_i[8] & sel_one_hot_i[0];
  assign data_masked[7] = data_i[7] & sel_one_hot_i[0];
  assign data_masked[6] = data_i[6] & sel_one_hot_i[0];
  assign data_masked[5] = data_i[5] & sel_one_hot_i[0];
  assign data_masked[4] = data_i[4] & sel_one_hot_i[0];
  assign data_masked[3] = data_i[3] & sel_one_hot_i[0];
  assign data_masked[2] = data_i[2] & sel_one_hot_i[0];
  assign data_masked[1] = data_i[1] & sel_one_hot_i[0];
  assign data_masked[0] = data_i[0] & sel_one_hot_i[0];
  assign data_masked[255] = data_i[255] & sel_one_hot_i[1];
  assign data_masked[254] = data_i[254] & sel_one_hot_i[1];
  assign data_masked[253] = data_i[253] & sel_one_hot_i[1];
  assign data_masked[252] = data_i[252] & sel_one_hot_i[1];
  assign data_masked[251] = data_i[251] & sel_one_hot_i[1];
  assign data_masked[250] = data_i[250] & sel_one_hot_i[1];
  assign data_masked[249] = data_i[249] & sel_one_hot_i[1];
  assign data_masked[248] = data_i[248] & sel_one_hot_i[1];
  assign data_masked[247] = data_i[247] & sel_one_hot_i[1];
  assign data_masked[246] = data_i[246] & sel_one_hot_i[1];
  assign data_masked[245] = data_i[245] & sel_one_hot_i[1];
  assign data_masked[244] = data_i[244] & sel_one_hot_i[1];
  assign data_masked[243] = data_i[243] & sel_one_hot_i[1];
  assign data_masked[242] = data_i[242] & sel_one_hot_i[1];
  assign data_masked[241] = data_i[241] & sel_one_hot_i[1];
  assign data_masked[240] = data_i[240] & sel_one_hot_i[1];
  assign data_masked[239] = data_i[239] & sel_one_hot_i[1];
  assign data_masked[238] = data_i[238] & sel_one_hot_i[1];
  assign data_masked[237] = data_i[237] & sel_one_hot_i[1];
  assign data_masked[236] = data_i[236] & sel_one_hot_i[1];
  assign data_masked[235] = data_i[235] & sel_one_hot_i[1];
  assign data_masked[234] = data_i[234] & sel_one_hot_i[1];
  assign data_masked[233] = data_i[233] & sel_one_hot_i[1];
  assign data_masked[232] = data_i[232] & sel_one_hot_i[1];
  assign data_masked[231] = data_i[231] & sel_one_hot_i[1];
  assign data_masked[230] = data_i[230] & sel_one_hot_i[1];
  assign data_masked[229] = data_i[229] & sel_one_hot_i[1];
  assign data_masked[228] = data_i[228] & sel_one_hot_i[1];
  assign data_masked[227] = data_i[227] & sel_one_hot_i[1];
  assign data_masked[226] = data_i[226] & sel_one_hot_i[1];
  assign data_masked[225] = data_i[225] & sel_one_hot_i[1];
  assign data_masked[224] = data_i[224] & sel_one_hot_i[1];
  assign data_masked[223] = data_i[223] & sel_one_hot_i[1];
  assign data_masked[222] = data_i[222] & sel_one_hot_i[1];
  assign data_masked[221] = data_i[221] & sel_one_hot_i[1];
  assign data_masked[220] = data_i[220] & sel_one_hot_i[1];
  assign data_masked[219] = data_i[219] & sel_one_hot_i[1];
  assign data_masked[218] = data_i[218] & sel_one_hot_i[1];
  assign data_masked[217] = data_i[217] & sel_one_hot_i[1];
  assign data_masked[216] = data_i[216] & sel_one_hot_i[1];
  assign data_masked[215] = data_i[215] & sel_one_hot_i[1];
  assign data_masked[214] = data_i[214] & sel_one_hot_i[1];
  assign data_masked[213] = data_i[213] & sel_one_hot_i[1];
  assign data_masked[212] = data_i[212] & sel_one_hot_i[1];
  assign data_masked[211] = data_i[211] & sel_one_hot_i[1];
  assign data_masked[210] = data_i[210] & sel_one_hot_i[1];
  assign data_masked[209] = data_i[209] & sel_one_hot_i[1];
  assign data_masked[208] = data_i[208] & sel_one_hot_i[1];
  assign data_masked[207] = data_i[207] & sel_one_hot_i[1];
  assign data_masked[206] = data_i[206] & sel_one_hot_i[1];
  assign data_masked[205] = data_i[205] & sel_one_hot_i[1];
  assign data_masked[204] = data_i[204] & sel_one_hot_i[1];
  assign data_masked[203] = data_i[203] & sel_one_hot_i[1];
  assign data_masked[202] = data_i[202] & sel_one_hot_i[1];
  assign data_masked[201] = data_i[201] & sel_one_hot_i[1];
  assign data_masked[200] = data_i[200] & sel_one_hot_i[1];
  assign data_masked[199] = data_i[199] & sel_one_hot_i[1];
  assign data_masked[198] = data_i[198] & sel_one_hot_i[1];
  assign data_masked[197] = data_i[197] & sel_one_hot_i[1];
  assign data_masked[196] = data_i[196] & sel_one_hot_i[1];
  assign data_masked[195] = data_i[195] & sel_one_hot_i[1];
  assign data_masked[194] = data_i[194] & sel_one_hot_i[1];
  assign data_masked[193] = data_i[193] & sel_one_hot_i[1];
  assign data_masked[192] = data_i[192] & sel_one_hot_i[1];
  assign data_masked[191] = data_i[191] & sel_one_hot_i[1];
  assign data_masked[190] = data_i[190] & sel_one_hot_i[1];
  assign data_masked[189] = data_i[189] & sel_one_hot_i[1];
  assign data_masked[188] = data_i[188] & sel_one_hot_i[1];
  assign data_masked[187] = data_i[187] & sel_one_hot_i[1];
  assign data_masked[186] = data_i[186] & sel_one_hot_i[1];
  assign data_masked[185] = data_i[185] & sel_one_hot_i[1];
  assign data_masked[184] = data_i[184] & sel_one_hot_i[1];
  assign data_masked[183] = data_i[183] & sel_one_hot_i[1];
  assign data_masked[182] = data_i[182] & sel_one_hot_i[1];
  assign data_masked[181] = data_i[181] & sel_one_hot_i[1];
  assign data_masked[180] = data_i[180] & sel_one_hot_i[1];
  assign data_masked[179] = data_i[179] & sel_one_hot_i[1];
  assign data_masked[178] = data_i[178] & sel_one_hot_i[1];
  assign data_masked[177] = data_i[177] & sel_one_hot_i[1];
  assign data_masked[176] = data_i[176] & sel_one_hot_i[1];
  assign data_masked[175] = data_i[175] & sel_one_hot_i[1];
  assign data_masked[174] = data_i[174] & sel_one_hot_i[1];
  assign data_masked[173] = data_i[173] & sel_one_hot_i[1];
  assign data_masked[172] = data_i[172] & sel_one_hot_i[1];
  assign data_masked[171] = data_i[171] & sel_one_hot_i[1];
  assign data_masked[170] = data_i[170] & sel_one_hot_i[1];
  assign data_masked[169] = data_i[169] & sel_one_hot_i[1];
  assign data_masked[168] = data_i[168] & sel_one_hot_i[1];
  assign data_masked[167] = data_i[167] & sel_one_hot_i[1];
  assign data_masked[166] = data_i[166] & sel_one_hot_i[1];
  assign data_masked[165] = data_i[165] & sel_one_hot_i[1];
  assign data_masked[164] = data_i[164] & sel_one_hot_i[1];
  assign data_masked[163] = data_i[163] & sel_one_hot_i[1];
  assign data_masked[162] = data_i[162] & sel_one_hot_i[1];
  assign data_masked[161] = data_i[161] & sel_one_hot_i[1];
  assign data_masked[160] = data_i[160] & sel_one_hot_i[1];
  assign data_masked[159] = data_i[159] & sel_one_hot_i[1];
  assign data_masked[158] = data_i[158] & sel_one_hot_i[1];
  assign data_masked[157] = data_i[157] & sel_one_hot_i[1];
  assign data_masked[156] = data_i[156] & sel_one_hot_i[1];
  assign data_masked[155] = data_i[155] & sel_one_hot_i[1];
  assign data_masked[154] = data_i[154] & sel_one_hot_i[1];
  assign data_masked[153] = data_i[153] & sel_one_hot_i[1];
  assign data_masked[152] = data_i[152] & sel_one_hot_i[1];
  assign data_masked[151] = data_i[151] & sel_one_hot_i[1];
  assign data_masked[150] = data_i[150] & sel_one_hot_i[1];
  assign data_masked[149] = data_i[149] & sel_one_hot_i[1];
  assign data_masked[148] = data_i[148] & sel_one_hot_i[1];
  assign data_masked[147] = data_i[147] & sel_one_hot_i[1];
  assign data_masked[146] = data_i[146] & sel_one_hot_i[1];
  assign data_masked[145] = data_i[145] & sel_one_hot_i[1];
  assign data_masked[144] = data_i[144] & sel_one_hot_i[1];
  assign data_masked[143] = data_i[143] & sel_one_hot_i[1];
  assign data_masked[142] = data_i[142] & sel_one_hot_i[1];
  assign data_masked[141] = data_i[141] & sel_one_hot_i[1];
  assign data_masked[140] = data_i[140] & sel_one_hot_i[1];
  assign data_masked[139] = data_i[139] & sel_one_hot_i[1];
  assign data_masked[138] = data_i[138] & sel_one_hot_i[1];
  assign data_masked[137] = data_i[137] & sel_one_hot_i[1];
  assign data_masked[136] = data_i[136] & sel_one_hot_i[1];
  assign data_masked[135] = data_i[135] & sel_one_hot_i[1];
  assign data_masked[134] = data_i[134] & sel_one_hot_i[1];
  assign data_masked[133] = data_i[133] & sel_one_hot_i[1];
  assign data_masked[132] = data_i[132] & sel_one_hot_i[1];
  assign data_masked[131] = data_i[131] & sel_one_hot_i[1];
  assign data_masked[130] = data_i[130] & sel_one_hot_i[1];
  assign data_masked[129] = data_i[129] & sel_one_hot_i[1];
  assign data_masked[128] = data_i[128] & sel_one_hot_i[1];
  assign data_masked[383] = data_i[383] & sel_one_hot_i[2];
  assign data_masked[382] = data_i[382] & sel_one_hot_i[2];
  assign data_masked[381] = data_i[381] & sel_one_hot_i[2];
  assign data_masked[380] = data_i[380] & sel_one_hot_i[2];
  assign data_masked[379] = data_i[379] & sel_one_hot_i[2];
  assign data_masked[378] = data_i[378] & sel_one_hot_i[2];
  assign data_masked[377] = data_i[377] & sel_one_hot_i[2];
  assign data_masked[376] = data_i[376] & sel_one_hot_i[2];
  assign data_masked[375] = data_i[375] & sel_one_hot_i[2];
  assign data_masked[374] = data_i[374] & sel_one_hot_i[2];
  assign data_masked[373] = data_i[373] & sel_one_hot_i[2];
  assign data_masked[372] = data_i[372] & sel_one_hot_i[2];
  assign data_masked[371] = data_i[371] & sel_one_hot_i[2];
  assign data_masked[370] = data_i[370] & sel_one_hot_i[2];
  assign data_masked[369] = data_i[369] & sel_one_hot_i[2];
  assign data_masked[368] = data_i[368] & sel_one_hot_i[2];
  assign data_masked[367] = data_i[367] & sel_one_hot_i[2];
  assign data_masked[366] = data_i[366] & sel_one_hot_i[2];
  assign data_masked[365] = data_i[365] & sel_one_hot_i[2];
  assign data_masked[364] = data_i[364] & sel_one_hot_i[2];
  assign data_masked[363] = data_i[363] & sel_one_hot_i[2];
  assign data_masked[362] = data_i[362] & sel_one_hot_i[2];
  assign data_masked[361] = data_i[361] & sel_one_hot_i[2];
  assign data_masked[360] = data_i[360] & sel_one_hot_i[2];
  assign data_masked[359] = data_i[359] & sel_one_hot_i[2];
  assign data_masked[358] = data_i[358] & sel_one_hot_i[2];
  assign data_masked[357] = data_i[357] & sel_one_hot_i[2];
  assign data_masked[356] = data_i[356] & sel_one_hot_i[2];
  assign data_masked[355] = data_i[355] & sel_one_hot_i[2];
  assign data_masked[354] = data_i[354] & sel_one_hot_i[2];
  assign data_masked[353] = data_i[353] & sel_one_hot_i[2];
  assign data_masked[352] = data_i[352] & sel_one_hot_i[2];
  assign data_masked[351] = data_i[351] & sel_one_hot_i[2];
  assign data_masked[350] = data_i[350] & sel_one_hot_i[2];
  assign data_masked[349] = data_i[349] & sel_one_hot_i[2];
  assign data_masked[348] = data_i[348] & sel_one_hot_i[2];
  assign data_masked[347] = data_i[347] & sel_one_hot_i[2];
  assign data_masked[346] = data_i[346] & sel_one_hot_i[2];
  assign data_masked[345] = data_i[345] & sel_one_hot_i[2];
  assign data_masked[344] = data_i[344] & sel_one_hot_i[2];
  assign data_masked[343] = data_i[343] & sel_one_hot_i[2];
  assign data_masked[342] = data_i[342] & sel_one_hot_i[2];
  assign data_masked[341] = data_i[341] & sel_one_hot_i[2];
  assign data_masked[340] = data_i[340] & sel_one_hot_i[2];
  assign data_masked[339] = data_i[339] & sel_one_hot_i[2];
  assign data_masked[338] = data_i[338] & sel_one_hot_i[2];
  assign data_masked[337] = data_i[337] & sel_one_hot_i[2];
  assign data_masked[336] = data_i[336] & sel_one_hot_i[2];
  assign data_masked[335] = data_i[335] & sel_one_hot_i[2];
  assign data_masked[334] = data_i[334] & sel_one_hot_i[2];
  assign data_masked[333] = data_i[333] & sel_one_hot_i[2];
  assign data_masked[332] = data_i[332] & sel_one_hot_i[2];
  assign data_masked[331] = data_i[331] & sel_one_hot_i[2];
  assign data_masked[330] = data_i[330] & sel_one_hot_i[2];
  assign data_masked[329] = data_i[329] & sel_one_hot_i[2];
  assign data_masked[328] = data_i[328] & sel_one_hot_i[2];
  assign data_masked[327] = data_i[327] & sel_one_hot_i[2];
  assign data_masked[326] = data_i[326] & sel_one_hot_i[2];
  assign data_masked[325] = data_i[325] & sel_one_hot_i[2];
  assign data_masked[324] = data_i[324] & sel_one_hot_i[2];
  assign data_masked[323] = data_i[323] & sel_one_hot_i[2];
  assign data_masked[322] = data_i[322] & sel_one_hot_i[2];
  assign data_masked[321] = data_i[321] & sel_one_hot_i[2];
  assign data_masked[320] = data_i[320] & sel_one_hot_i[2];
  assign data_masked[319] = data_i[319] & sel_one_hot_i[2];
  assign data_masked[318] = data_i[318] & sel_one_hot_i[2];
  assign data_masked[317] = data_i[317] & sel_one_hot_i[2];
  assign data_masked[316] = data_i[316] & sel_one_hot_i[2];
  assign data_masked[315] = data_i[315] & sel_one_hot_i[2];
  assign data_masked[314] = data_i[314] & sel_one_hot_i[2];
  assign data_masked[313] = data_i[313] & sel_one_hot_i[2];
  assign data_masked[312] = data_i[312] & sel_one_hot_i[2];
  assign data_masked[311] = data_i[311] & sel_one_hot_i[2];
  assign data_masked[310] = data_i[310] & sel_one_hot_i[2];
  assign data_masked[309] = data_i[309] & sel_one_hot_i[2];
  assign data_masked[308] = data_i[308] & sel_one_hot_i[2];
  assign data_masked[307] = data_i[307] & sel_one_hot_i[2];
  assign data_masked[306] = data_i[306] & sel_one_hot_i[2];
  assign data_masked[305] = data_i[305] & sel_one_hot_i[2];
  assign data_masked[304] = data_i[304] & sel_one_hot_i[2];
  assign data_masked[303] = data_i[303] & sel_one_hot_i[2];
  assign data_masked[302] = data_i[302] & sel_one_hot_i[2];
  assign data_masked[301] = data_i[301] & sel_one_hot_i[2];
  assign data_masked[300] = data_i[300] & sel_one_hot_i[2];
  assign data_masked[299] = data_i[299] & sel_one_hot_i[2];
  assign data_masked[298] = data_i[298] & sel_one_hot_i[2];
  assign data_masked[297] = data_i[297] & sel_one_hot_i[2];
  assign data_masked[296] = data_i[296] & sel_one_hot_i[2];
  assign data_masked[295] = data_i[295] & sel_one_hot_i[2];
  assign data_masked[294] = data_i[294] & sel_one_hot_i[2];
  assign data_masked[293] = data_i[293] & sel_one_hot_i[2];
  assign data_masked[292] = data_i[292] & sel_one_hot_i[2];
  assign data_masked[291] = data_i[291] & sel_one_hot_i[2];
  assign data_masked[290] = data_i[290] & sel_one_hot_i[2];
  assign data_masked[289] = data_i[289] & sel_one_hot_i[2];
  assign data_masked[288] = data_i[288] & sel_one_hot_i[2];
  assign data_masked[287] = data_i[287] & sel_one_hot_i[2];
  assign data_masked[286] = data_i[286] & sel_one_hot_i[2];
  assign data_masked[285] = data_i[285] & sel_one_hot_i[2];
  assign data_masked[284] = data_i[284] & sel_one_hot_i[2];
  assign data_masked[283] = data_i[283] & sel_one_hot_i[2];
  assign data_masked[282] = data_i[282] & sel_one_hot_i[2];
  assign data_masked[281] = data_i[281] & sel_one_hot_i[2];
  assign data_masked[280] = data_i[280] & sel_one_hot_i[2];
  assign data_masked[279] = data_i[279] & sel_one_hot_i[2];
  assign data_masked[278] = data_i[278] & sel_one_hot_i[2];
  assign data_masked[277] = data_i[277] & sel_one_hot_i[2];
  assign data_masked[276] = data_i[276] & sel_one_hot_i[2];
  assign data_masked[275] = data_i[275] & sel_one_hot_i[2];
  assign data_masked[274] = data_i[274] & sel_one_hot_i[2];
  assign data_masked[273] = data_i[273] & sel_one_hot_i[2];
  assign data_masked[272] = data_i[272] & sel_one_hot_i[2];
  assign data_masked[271] = data_i[271] & sel_one_hot_i[2];
  assign data_masked[270] = data_i[270] & sel_one_hot_i[2];
  assign data_masked[269] = data_i[269] & sel_one_hot_i[2];
  assign data_masked[268] = data_i[268] & sel_one_hot_i[2];
  assign data_masked[267] = data_i[267] & sel_one_hot_i[2];
  assign data_masked[266] = data_i[266] & sel_one_hot_i[2];
  assign data_masked[265] = data_i[265] & sel_one_hot_i[2];
  assign data_masked[264] = data_i[264] & sel_one_hot_i[2];
  assign data_masked[263] = data_i[263] & sel_one_hot_i[2];
  assign data_masked[262] = data_i[262] & sel_one_hot_i[2];
  assign data_masked[261] = data_i[261] & sel_one_hot_i[2];
  assign data_masked[260] = data_i[260] & sel_one_hot_i[2];
  assign data_masked[259] = data_i[259] & sel_one_hot_i[2];
  assign data_masked[258] = data_i[258] & sel_one_hot_i[2];
  assign data_masked[257] = data_i[257] & sel_one_hot_i[2];
  assign data_masked[256] = data_i[256] & sel_one_hot_i[2];
  assign data_masked[511] = data_i[511] & sel_one_hot_i[3];
  assign data_masked[510] = data_i[510] & sel_one_hot_i[3];
  assign data_masked[509] = data_i[509] & sel_one_hot_i[3];
  assign data_masked[508] = data_i[508] & sel_one_hot_i[3];
  assign data_masked[507] = data_i[507] & sel_one_hot_i[3];
  assign data_masked[506] = data_i[506] & sel_one_hot_i[3];
  assign data_masked[505] = data_i[505] & sel_one_hot_i[3];
  assign data_masked[504] = data_i[504] & sel_one_hot_i[3];
  assign data_masked[503] = data_i[503] & sel_one_hot_i[3];
  assign data_masked[502] = data_i[502] & sel_one_hot_i[3];
  assign data_masked[501] = data_i[501] & sel_one_hot_i[3];
  assign data_masked[500] = data_i[500] & sel_one_hot_i[3];
  assign data_masked[499] = data_i[499] & sel_one_hot_i[3];
  assign data_masked[498] = data_i[498] & sel_one_hot_i[3];
  assign data_masked[497] = data_i[497] & sel_one_hot_i[3];
  assign data_masked[496] = data_i[496] & sel_one_hot_i[3];
  assign data_masked[495] = data_i[495] & sel_one_hot_i[3];
  assign data_masked[494] = data_i[494] & sel_one_hot_i[3];
  assign data_masked[493] = data_i[493] & sel_one_hot_i[3];
  assign data_masked[492] = data_i[492] & sel_one_hot_i[3];
  assign data_masked[491] = data_i[491] & sel_one_hot_i[3];
  assign data_masked[490] = data_i[490] & sel_one_hot_i[3];
  assign data_masked[489] = data_i[489] & sel_one_hot_i[3];
  assign data_masked[488] = data_i[488] & sel_one_hot_i[3];
  assign data_masked[487] = data_i[487] & sel_one_hot_i[3];
  assign data_masked[486] = data_i[486] & sel_one_hot_i[3];
  assign data_masked[485] = data_i[485] & sel_one_hot_i[3];
  assign data_masked[484] = data_i[484] & sel_one_hot_i[3];
  assign data_masked[483] = data_i[483] & sel_one_hot_i[3];
  assign data_masked[482] = data_i[482] & sel_one_hot_i[3];
  assign data_masked[481] = data_i[481] & sel_one_hot_i[3];
  assign data_masked[480] = data_i[480] & sel_one_hot_i[3];
  assign data_masked[479] = data_i[479] & sel_one_hot_i[3];
  assign data_masked[478] = data_i[478] & sel_one_hot_i[3];
  assign data_masked[477] = data_i[477] & sel_one_hot_i[3];
  assign data_masked[476] = data_i[476] & sel_one_hot_i[3];
  assign data_masked[475] = data_i[475] & sel_one_hot_i[3];
  assign data_masked[474] = data_i[474] & sel_one_hot_i[3];
  assign data_masked[473] = data_i[473] & sel_one_hot_i[3];
  assign data_masked[472] = data_i[472] & sel_one_hot_i[3];
  assign data_masked[471] = data_i[471] & sel_one_hot_i[3];
  assign data_masked[470] = data_i[470] & sel_one_hot_i[3];
  assign data_masked[469] = data_i[469] & sel_one_hot_i[3];
  assign data_masked[468] = data_i[468] & sel_one_hot_i[3];
  assign data_masked[467] = data_i[467] & sel_one_hot_i[3];
  assign data_masked[466] = data_i[466] & sel_one_hot_i[3];
  assign data_masked[465] = data_i[465] & sel_one_hot_i[3];
  assign data_masked[464] = data_i[464] & sel_one_hot_i[3];
  assign data_masked[463] = data_i[463] & sel_one_hot_i[3];
  assign data_masked[462] = data_i[462] & sel_one_hot_i[3];
  assign data_masked[461] = data_i[461] & sel_one_hot_i[3];
  assign data_masked[460] = data_i[460] & sel_one_hot_i[3];
  assign data_masked[459] = data_i[459] & sel_one_hot_i[3];
  assign data_masked[458] = data_i[458] & sel_one_hot_i[3];
  assign data_masked[457] = data_i[457] & sel_one_hot_i[3];
  assign data_masked[456] = data_i[456] & sel_one_hot_i[3];
  assign data_masked[455] = data_i[455] & sel_one_hot_i[3];
  assign data_masked[454] = data_i[454] & sel_one_hot_i[3];
  assign data_masked[453] = data_i[453] & sel_one_hot_i[3];
  assign data_masked[452] = data_i[452] & sel_one_hot_i[3];
  assign data_masked[451] = data_i[451] & sel_one_hot_i[3];
  assign data_masked[450] = data_i[450] & sel_one_hot_i[3];
  assign data_masked[449] = data_i[449] & sel_one_hot_i[3];
  assign data_masked[448] = data_i[448] & sel_one_hot_i[3];
  assign data_masked[447] = data_i[447] & sel_one_hot_i[3];
  assign data_masked[446] = data_i[446] & sel_one_hot_i[3];
  assign data_masked[445] = data_i[445] & sel_one_hot_i[3];
  assign data_masked[444] = data_i[444] & sel_one_hot_i[3];
  assign data_masked[443] = data_i[443] & sel_one_hot_i[3];
  assign data_masked[442] = data_i[442] & sel_one_hot_i[3];
  assign data_masked[441] = data_i[441] & sel_one_hot_i[3];
  assign data_masked[440] = data_i[440] & sel_one_hot_i[3];
  assign data_masked[439] = data_i[439] & sel_one_hot_i[3];
  assign data_masked[438] = data_i[438] & sel_one_hot_i[3];
  assign data_masked[437] = data_i[437] & sel_one_hot_i[3];
  assign data_masked[436] = data_i[436] & sel_one_hot_i[3];
  assign data_masked[435] = data_i[435] & sel_one_hot_i[3];
  assign data_masked[434] = data_i[434] & sel_one_hot_i[3];
  assign data_masked[433] = data_i[433] & sel_one_hot_i[3];
  assign data_masked[432] = data_i[432] & sel_one_hot_i[3];
  assign data_masked[431] = data_i[431] & sel_one_hot_i[3];
  assign data_masked[430] = data_i[430] & sel_one_hot_i[3];
  assign data_masked[429] = data_i[429] & sel_one_hot_i[3];
  assign data_masked[428] = data_i[428] & sel_one_hot_i[3];
  assign data_masked[427] = data_i[427] & sel_one_hot_i[3];
  assign data_masked[426] = data_i[426] & sel_one_hot_i[3];
  assign data_masked[425] = data_i[425] & sel_one_hot_i[3];
  assign data_masked[424] = data_i[424] & sel_one_hot_i[3];
  assign data_masked[423] = data_i[423] & sel_one_hot_i[3];
  assign data_masked[422] = data_i[422] & sel_one_hot_i[3];
  assign data_masked[421] = data_i[421] & sel_one_hot_i[3];
  assign data_masked[420] = data_i[420] & sel_one_hot_i[3];
  assign data_masked[419] = data_i[419] & sel_one_hot_i[3];
  assign data_masked[418] = data_i[418] & sel_one_hot_i[3];
  assign data_masked[417] = data_i[417] & sel_one_hot_i[3];
  assign data_masked[416] = data_i[416] & sel_one_hot_i[3];
  assign data_masked[415] = data_i[415] & sel_one_hot_i[3];
  assign data_masked[414] = data_i[414] & sel_one_hot_i[3];
  assign data_masked[413] = data_i[413] & sel_one_hot_i[3];
  assign data_masked[412] = data_i[412] & sel_one_hot_i[3];
  assign data_masked[411] = data_i[411] & sel_one_hot_i[3];
  assign data_masked[410] = data_i[410] & sel_one_hot_i[3];
  assign data_masked[409] = data_i[409] & sel_one_hot_i[3];
  assign data_masked[408] = data_i[408] & sel_one_hot_i[3];
  assign data_masked[407] = data_i[407] & sel_one_hot_i[3];
  assign data_masked[406] = data_i[406] & sel_one_hot_i[3];
  assign data_masked[405] = data_i[405] & sel_one_hot_i[3];
  assign data_masked[404] = data_i[404] & sel_one_hot_i[3];
  assign data_masked[403] = data_i[403] & sel_one_hot_i[3];
  assign data_masked[402] = data_i[402] & sel_one_hot_i[3];
  assign data_masked[401] = data_i[401] & sel_one_hot_i[3];
  assign data_masked[400] = data_i[400] & sel_one_hot_i[3];
  assign data_masked[399] = data_i[399] & sel_one_hot_i[3];
  assign data_masked[398] = data_i[398] & sel_one_hot_i[3];
  assign data_masked[397] = data_i[397] & sel_one_hot_i[3];
  assign data_masked[396] = data_i[396] & sel_one_hot_i[3];
  assign data_masked[395] = data_i[395] & sel_one_hot_i[3];
  assign data_masked[394] = data_i[394] & sel_one_hot_i[3];
  assign data_masked[393] = data_i[393] & sel_one_hot_i[3];
  assign data_masked[392] = data_i[392] & sel_one_hot_i[3];
  assign data_masked[391] = data_i[391] & sel_one_hot_i[3];
  assign data_masked[390] = data_i[390] & sel_one_hot_i[3];
  assign data_masked[389] = data_i[389] & sel_one_hot_i[3];
  assign data_masked[388] = data_i[388] & sel_one_hot_i[3];
  assign data_masked[387] = data_i[387] & sel_one_hot_i[3];
  assign data_masked[386] = data_i[386] & sel_one_hot_i[3];
  assign data_masked[385] = data_i[385] & sel_one_hot_i[3];
  assign data_masked[384] = data_i[384] & sel_one_hot_i[3];
  assign data_masked[639] = data_i[639] & sel_one_hot_i[4];
  assign data_masked[638] = data_i[638] & sel_one_hot_i[4];
  assign data_masked[637] = data_i[637] & sel_one_hot_i[4];
  assign data_masked[636] = data_i[636] & sel_one_hot_i[4];
  assign data_masked[635] = data_i[635] & sel_one_hot_i[4];
  assign data_masked[634] = data_i[634] & sel_one_hot_i[4];
  assign data_masked[633] = data_i[633] & sel_one_hot_i[4];
  assign data_masked[632] = data_i[632] & sel_one_hot_i[4];
  assign data_masked[631] = data_i[631] & sel_one_hot_i[4];
  assign data_masked[630] = data_i[630] & sel_one_hot_i[4];
  assign data_masked[629] = data_i[629] & sel_one_hot_i[4];
  assign data_masked[628] = data_i[628] & sel_one_hot_i[4];
  assign data_masked[627] = data_i[627] & sel_one_hot_i[4];
  assign data_masked[626] = data_i[626] & sel_one_hot_i[4];
  assign data_masked[625] = data_i[625] & sel_one_hot_i[4];
  assign data_masked[624] = data_i[624] & sel_one_hot_i[4];
  assign data_masked[623] = data_i[623] & sel_one_hot_i[4];
  assign data_masked[622] = data_i[622] & sel_one_hot_i[4];
  assign data_masked[621] = data_i[621] & sel_one_hot_i[4];
  assign data_masked[620] = data_i[620] & sel_one_hot_i[4];
  assign data_masked[619] = data_i[619] & sel_one_hot_i[4];
  assign data_masked[618] = data_i[618] & sel_one_hot_i[4];
  assign data_masked[617] = data_i[617] & sel_one_hot_i[4];
  assign data_masked[616] = data_i[616] & sel_one_hot_i[4];
  assign data_masked[615] = data_i[615] & sel_one_hot_i[4];
  assign data_masked[614] = data_i[614] & sel_one_hot_i[4];
  assign data_masked[613] = data_i[613] & sel_one_hot_i[4];
  assign data_masked[612] = data_i[612] & sel_one_hot_i[4];
  assign data_masked[611] = data_i[611] & sel_one_hot_i[4];
  assign data_masked[610] = data_i[610] & sel_one_hot_i[4];
  assign data_masked[609] = data_i[609] & sel_one_hot_i[4];
  assign data_masked[608] = data_i[608] & sel_one_hot_i[4];
  assign data_masked[607] = data_i[607] & sel_one_hot_i[4];
  assign data_masked[606] = data_i[606] & sel_one_hot_i[4];
  assign data_masked[605] = data_i[605] & sel_one_hot_i[4];
  assign data_masked[604] = data_i[604] & sel_one_hot_i[4];
  assign data_masked[603] = data_i[603] & sel_one_hot_i[4];
  assign data_masked[602] = data_i[602] & sel_one_hot_i[4];
  assign data_masked[601] = data_i[601] & sel_one_hot_i[4];
  assign data_masked[600] = data_i[600] & sel_one_hot_i[4];
  assign data_masked[599] = data_i[599] & sel_one_hot_i[4];
  assign data_masked[598] = data_i[598] & sel_one_hot_i[4];
  assign data_masked[597] = data_i[597] & sel_one_hot_i[4];
  assign data_masked[596] = data_i[596] & sel_one_hot_i[4];
  assign data_masked[595] = data_i[595] & sel_one_hot_i[4];
  assign data_masked[594] = data_i[594] & sel_one_hot_i[4];
  assign data_masked[593] = data_i[593] & sel_one_hot_i[4];
  assign data_masked[592] = data_i[592] & sel_one_hot_i[4];
  assign data_masked[591] = data_i[591] & sel_one_hot_i[4];
  assign data_masked[590] = data_i[590] & sel_one_hot_i[4];
  assign data_masked[589] = data_i[589] & sel_one_hot_i[4];
  assign data_masked[588] = data_i[588] & sel_one_hot_i[4];
  assign data_masked[587] = data_i[587] & sel_one_hot_i[4];
  assign data_masked[586] = data_i[586] & sel_one_hot_i[4];
  assign data_masked[585] = data_i[585] & sel_one_hot_i[4];
  assign data_masked[584] = data_i[584] & sel_one_hot_i[4];
  assign data_masked[583] = data_i[583] & sel_one_hot_i[4];
  assign data_masked[582] = data_i[582] & sel_one_hot_i[4];
  assign data_masked[581] = data_i[581] & sel_one_hot_i[4];
  assign data_masked[580] = data_i[580] & sel_one_hot_i[4];
  assign data_masked[579] = data_i[579] & sel_one_hot_i[4];
  assign data_masked[578] = data_i[578] & sel_one_hot_i[4];
  assign data_masked[577] = data_i[577] & sel_one_hot_i[4];
  assign data_masked[576] = data_i[576] & sel_one_hot_i[4];
  assign data_masked[575] = data_i[575] & sel_one_hot_i[4];
  assign data_masked[574] = data_i[574] & sel_one_hot_i[4];
  assign data_masked[573] = data_i[573] & sel_one_hot_i[4];
  assign data_masked[572] = data_i[572] & sel_one_hot_i[4];
  assign data_masked[571] = data_i[571] & sel_one_hot_i[4];
  assign data_masked[570] = data_i[570] & sel_one_hot_i[4];
  assign data_masked[569] = data_i[569] & sel_one_hot_i[4];
  assign data_masked[568] = data_i[568] & sel_one_hot_i[4];
  assign data_masked[567] = data_i[567] & sel_one_hot_i[4];
  assign data_masked[566] = data_i[566] & sel_one_hot_i[4];
  assign data_masked[565] = data_i[565] & sel_one_hot_i[4];
  assign data_masked[564] = data_i[564] & sel_one_hot_i[4];
  assign data_masked[563] = data_i[563] & sel_one_hot_i[4];
  assign data_masked[562] = data_i[562] & sel_one_hot_i[4];
  assign data_masked[561] = data_i[561] & sel_one_hot_i[4];
  assign data_masked[560] = data_i[560] & sel_one_hot_i[4];
  assign data_masked[559] = data_i[559] & sel_one_hot_i[4];
  assign data_masked[558] = data_i[558] & sel_one_hot_i[4];
  assign data_masked[557] = data_i[557] & sel_one_hot_i[4];
  assign data_masked[556] = data_i[556] & sel_one_hot_i[4];
  assign data_masked[555] = data_i[555] & sel_one_hot_i[4];
  assign data_masked[554] = data_i[554] & sel_one_hot_i[4];
  assign data_masked[553] = data_i[553] & sel_one_hot_i[4];
  assign data_masked[552] = data_i[552] & sel_one_hot_i[4];
  assign data_masked[551] = data_i[551] & sel_one_hot_i[4];
  assign data_masked[550] = data_i[550] & sel_one_hot_i[4];
  assign data_masked[549] = data_i[549] & sel_one_hot_i[4];
  assign data_masked[548] = data_i[548] & sel_one_hot_i[4];
  assign data_masked[547] = data_i[547] & sel_one_hot_i[4];
  assign data_masked[546] = data_i[546] & sel_one_hot_i[4];
  assign data_masked[545] = data_i[545] & sel_one_hot_i[4];
  assign data_masked[544] = data_i[544] & sel_one_hot_i[4];
  assign data_masked[543] = data_i[543] & sel_one_hot_i[4];
  assign data_masked[542] = data_i[542] & sel_one_hot_i[4];
  assign data_masked[541] = data_i[541] & sel_one_hot_i[4];
  assign data_masked[540] = data_i[540] & sel_one_hot_i[4];
  assign data_masked[539] = data_i[539] & sel_one_hot_i[4];
  assign data_masked[538] = data_i[538] & sel_one_hot_i[4];
  assign data_masked[537] = data_i[537] & sel_one_hot_i[4];
  assign data_masked[536] = data_i[536] & sel_one_hot_i[4];
  assign data_masked[535] = data_i[535] & sel_one_hot_i[4];
  assign data_masked[534] = data_i[534] & sel_one_hot_i[4];
  assign data_masked[533] = data_i[533] & sel_one_hot_i[4];
  assign data_masked[532] = data_i[532] & sel_one_hot_i[4];
  assign data_masked[531] = data_i[531] & sel_one_hot_i[4];
  assign data_masked[530] = data_i[530] & sel_one_hot_i[4];
  assign data_masked[529] = data_i[529] & sel_one_hot_i[4];
  assign data_masked[528] = data_i[528] & sel_one_hot_i[4];
  assign data_masked[527] = data_i[527] & sel_one_hot_i[4];
  assign data_masked[526] = data_i[526] & sel_one_hot_i[4];
  assign data_masked[525] = data_i[525] & sel_one_hot_i[4];
  assign data_masked[524] = data_i[524] & sel_one_hot_i[4];
  assign data_masked[523] = data_i[523] & sel_one_hot_i[4];
  assign data_masked[522] = data_i[522] & sel_one_hot_i[4];
  assign data_masked[521] = data_i[521] & sel_one_hot_i[4];
  assign data_masked[520] = data_i[520] & sel_one_hot_i[4];
  assign data_masked[519] = data_i[519] & sel_one_hot_i[4];
  assign data_masked[518] = data_i[518] & sel_one_hot_i[4];
  assign data_masked[517] = data_i[517] & sel_one_hot_i[4];
  assign data_masked[516] = data_i[516] & sel_one_hot_i[4];
  assign data_masked[515] = data_i[515] & sel_one_hot_i[4];
  assign data_masked[514] = data_i[514] & sel_one_hot_i[4];
  assign data_masked[513] = data_i[513] & sel_one_hot_i[4];
  assign data_masked[512] = data_i[512] & sel_one_hot_i[4];
  assign data_masked[767] = data_i[767] & sel_one_hot_i[5];
  assign data_masked[766] = data_i[766] & sel_one_hot_i[5];
  assign data_masked[765] = data_i[765] & sel_one_hot_i[5];
  assign data_masked[764] = data_i[764] & sel_one_hot_i[5];
  assign data_masked[763] = data_i[763] & sel_one_hot_i[5];
  assign data_masked[762] = data_i[762] & sel_one_hot_i[5];
  assign data_masked[761] = data_i[761] & sel_one_hot_i[5];
  assign data_masked[760] = data_i[760] & sel_one_hot_i[5];
  assign data_masked[759] = data_i[759] & sel_one_hot_i[5];
  assign data_masked[758] = data_i[758] & sel_one_hot_i[5];
  assign data_masked[757] = data_i[757] & sel_one_hot_i[5];
  assign data_masked[756] = data_i[756] & sel_one_hot_i[5];
  assign data_masked[755] = data_i[755] & sel_one_hot_i[5];
  assign data_masked[754] = data_i[754] & sel_one_hot_i[5];
  assign data_masked[753] = data_i[753] & sel_one_hot_i[5];
  assign data_masked[752] = data_i[752] & sel_one_hot_i[5];
  assign data_masked[751] = data_i[751] & sel_one_hot_i[5];
  assign data_masked[750] = data_i[750] & sel_one_hot_i[5];
  assign data_masked[749] = data_i[749] & sel_one_hot_i[5];
  assign data_masked[748] = data_i[748] & sel_one_hot_i[5];
  assign data_masked[747] = data_i[747] & sel_one_hot_i[5];
  assign data_masked[746] = data_i[746] & sel_one_hot_i[5];
  assign data_masked[745] = data_i[745] & sel_one_hot_i[5];
  assign data_masked[744] = data_i[744] & sel_one_hot_i[5];
  assign data_masked[743] = data_i[743] & sel_one_hot_i[5];
  assign data_masked[742] = data_i[742] & sel_one_hot_i[5];
  assign data_masked[741] = data_i[741] & sel_one_hot_i[5];
  assign data_masked[740] = data_i[740] & sel_one_hot_i[5];
  assign data_masked[739] = data_i[739] & sel_one_hot_i[5];
  assign data_masked[738] = data_i[738] & sel_one_hot_i[5];
  assign data_masked[737] = data_i[737] & sel_one_hot_i[5];
  assign data_masked[736] = data_i[736] & sel_one_hot_i[5];
  assign data_masked[735] = data_i[735] & sel_one_hot_i[5];
  assign data_masked[734] = data_i[734] & sel_one_hot_i[5];
  assign data_masked[733] = data_i[733] & sel_one_hot_i[5];
  assign data_masked[732] = data_i[732] & sel_one_hot_i[5];
  assign data_masked[731] = data_i[731] & sel_one_hot_i[5];
  assign data_masked[730] = data_i[730] & sel_one_hot_i[5];
  assign data_masked[729] = data_i[729] & sel_one_hot_i[5];
  assign data_masked[728] = data_i[728] & sel_one_hot_i[5];
  assign data_masked[727] = data_i[727] & sel_one_hot_i[5];
  assign data_masked[726] = data_i[726] & sel_one_hot_i[5];
  assign data_masked[725] = data_i[725] & sel_one_hot_i[5];
  assign data_masked[724] = data_i[724] & sel_one_hot_i[5];
  assign data_masked[723] = data_i[723] & sel_one_hot_i[5];
  assign data_masked[722] = data_i[722] & sel_one_hot_i[5];
  assign data_masked[721] = data_i[721] & sel_one_hot_i[5];
  assign data_masked[720] = data_i[720] & sel_one_hot_i[5];
  assign data_masked[719] = data_i[719] & sel_one_hot_i[5];
  assign data_masked[718] = data_i[718] & sel_one_hot_i[5];
  assign data_masked[717] = data_i[717] & sel_one_hot_i[5];
  assign data_masked[716] = data_i[716] & sel_one_hot_i[5];
  assign data_masked[715] = data_i[715] & sel_one_hot_i[5];
  assign data_masked[714] = data_i[714] & sel_one_hot_i[5];
  assign data_masked[713] = data_i[713] & sel_one_hot_i[5];
  assign data_masked[712] = data_i[712] & sel_one_hot_i[5];
  assign data_masked[711] = data_i[711] & sel_one_hot_i[5];
  assign data_masked[710] = data_i[710] & sel_one_hot_i[5];
  assign data_masked[709] = data_i[709] & sel_one_hot_i[5];
  assign data_masked[708] = data_i[708] & sel_one_hot_i[5];
  assign data_masked[707] = data_i[707] & sel_one_hot_i[5];
  assign data_masked[706] = data_i[706] & sel_one_hot_i[5];
  assign data_masked[705] = data_i[705] & sel_one_hot_i[5];
  assign data_masked[704] = data_i[704] & sel_one_hot_i[5];
  assign data_masked[703] = data_i[703] & sel_one_hot_i[5];
  assign data_masked[702] = data_i[702] & sel_one_hot_i[5];
  assign data_masked[701] = data_i[701] & sel_one_hot_i[5];
  assign data_masked[700] = data_i[700] & sel_one_hot_i[5];
  assign data_masked[699] = data_i[699] & sel_one_hot_i[5];
  assign data_masked[698] = data_i[698] & sel_one_hot_i[5];
  assign data_masked[697] = data_i[697] & sel_one_hot_i[5];
  assign data_masked[696] = data_i[696] & sel_one_hot_i[5];
  assign data_masked[695] = data_i[695] & sel_one_hot_i[5];
  assign data_masked[694] = data_i[694] & sel_one_hot_i[5];
  assign data_masked[693] = data_i[693] & sel_one_hot_i[5];
  assign data_masked[692] = data_i[692] & sel_one_hot_i[5];
  assign data_masked[691] = data_i[691] & sel_one_hot_i[5];
  assign data_masked[690] = data_i[690] & sel_one_hot_i[5];
  assign data_masked[689] = data_i[689] & sel_one_hot_i[5];
  assign data_masked[688] = data_i[688] & sel_one_hot_i[5];
  assign data_masked[687] = data_i[687] & sel_one_hot_i[5];
  assign data_masked[686] = data_i[686] & sel_one_hot_i[5];
  assign data_masked[685] = data_i[685] & sel_one_hot_i[5];
  assign data_masked[684] = data_i[684] & sel_one_hot_i[5];
  assign data_masked[683] = data_i[683] & sel_one_hot_i[5];
  assign data_masked[682] = data_i[682] & sel_one_hot_i[5];
  assign data_masked[681] = data_i[681] & sel_one_hot_i[5];
  assign data_masked[680] = data_i[680] & sel_one_hot_i[5];
  assign data_masked[679] = data_i[679] & sel_one_hot_i[5];
  assign data_masked[678] = data_i[678] & sel_one_hot_i[5];
  assign data_masked[677] = data_i[677] & sel_one_hot_i[5];
  assign data_masked[676] = data_i[676] & sel_one_hot_i[5];
  assign data_masked[675] = data_i[675] & sel_one_hot_i[5];
  assign data_masked[674] = data_i[674] & sel_one_hot_i[5];
  assign data_masked[673] = data_i[673] & sel_one_hot_i[5];
  assign data_masked[672] = data_i[672] & sel_one_hot_i[5];
  assign data_masked[671] = data_i[671] & sel_one_hot_i[5];
  assign data_masked[670] = data_i[670] & sel_one_hot_i[5];
  assign data_masked[669] = data_i[669] & sel_one_hot_i[5];
  assign data_masked[668] = data_i[668] & sel_one_hot_i[5];
  assign data_masked[667] = data_i[667] & sel_one_hot_i[5];
  assign data_masked[666] = data_i[666] & sel_one_hot_i[5];
  assign data_masked[665] = data_i[665] & sel_one_hot_i[5];
  assign data_masked[664] = data_i[664] & sel_one_hot_i[5];
  assign data_masked[663] = data_i[663] & sel_one_hot_i[5];
  assign data_masked[662] = data_i[662] & sel_one_hot_i[5];
  assign data_masked[661] = data_i[661] & sel_one_hot_i[5];
  assign data_masked[660] = data_i[660] & sel_one_hot_i[5];
  assign data_masked[659] = data_i[659] & sel_one_hot_i[5];
  assign data_masked[658] = data_i[658] & sel_one_hot_i[5];
  assign data_masked[657] = data_i[657] & sel_one_hot_i[5];
  assign data_masked[656] = data_i[656] & sel_one_hot_i[5];
  assign data_masked[655] = data_i[655] & sel_one_hot_i[5];
  assign data_masked[654] = data_i[654] & sel_one_hot_i[5];
  assign data_masked[653] = data_i[653] & sel_one_hot_i[5];
  assign data_masked[652] = data_i[652] & sel_one_hot_i[5];
  assign data_masked[651] = data_i[651] & sel_one_hot_i[5];
  assign data_masked[650] = data_i[650] & sel_one_hot_i[5];
  assign data_masked[649] = data_i[649] & sel_one_hot_i[5];
  assign data_masked[648] = data_i[648] & sel_one_hot_i[5];
  assign data_masked[647] = data_i[647] & sel_one_hot_i[5];
  assign data_masked[646] = data_i[646] & sel_one_hot_i[5];
  assign data_masked[645] = data_i[645] & sel_one_hot_i[5];
  assign data_masked[644] = data_i[644] & sel_one_hot_i[5];
  assign data_masked[643] = data_i[643] & sel_one_hot_i[5];
  assign data_masked[642] = data_i[642] & sel_one_hot_i[5];
  assign data_masked[641] = data_i[641] & sel_one_hot_i[5];
  assign data_masked[640] = data_i[640] & sel_one_hot_i[5];
  assign data_masked[895] = data_i[895] & sel_one_hot_i[6];
  assign data_masked[894] = data_i[894] & sel_one_hot_i[6];
  assign data_masked[893] = data_i[893] & sel_one_hot_i[6];
  assign data_masked[892] = data_i[892] & sel_one_hot_i[6];
  assign data_masked[891] = data_i[891] & sel_one_hot_i[6];
  assign data_masked[890] = data_i[890] & sel_one_hot_i[6];
  assign data_masked[889] = data_i[889] & sel_one_hot_i[6];
  assign data_masked[888] = data_i[888] & sel_one_hot_i[6];
  assign data_masked[887] = data_i[887] & sel_one_hot_i[6];
  assign data_masked[886] = data_i[886] & sel_one_hot_i[6];
  assign data_masked[885] = data_i[885] & sel_one_hot_i[6];
  assign data_masked[884] = data_i[884] & sel_one_hot_i[6];
  assign data_masked[883] = data_i[883] & sel_one_hot_i[6];
  assign data_masked[882] = data_i[882] & sel_one_hot_i[6];
  assign data_masked[881] = data_i[881] & sel_one_hot_i[6];
  assign data_masked[880] = data_i[880] & sel_one_hot_i[6];
  assign data_masked[879] = data_i[879] & sel_one_hot_i[6];
  assign data_masked[878] = data_i[878] & sel_one_hot_i[6];
  assign data_masked[877] = data_i[877] & sel_one_hot_i[6];
  assign data_masked[876] = data_i[876] & sel_one_hot_i[6];
  assign data_masked[875] = data_i[875] & sel_one_hot_i[6];
  assign data_masked[874] = data_i[874] & sel_one_hot_i[6];
  assign data_masked[873] = data_i[873] & sel_one_hot_i[6];
  assign data_masked[872] = data_i[872] & sel_one_hot_i[6];
  assign data_masked[871] = data_i[871] & sel_one_hot_i[6];
  assign data_masked[870] = data_i[870] & sel_one_hot_i[6];
  assign data_masked[869] = data_i[869] & sel_one_hot_i[6];
  assign data_masked[868] = data_i[868] & sel_one_hot_i[6];
  assign data_masked[867] = data_i[867] & sel_one_hot_i[6];
  assign data_masked[866] = data_i[866] & sel_one_hot_i[6];
  assign data_masked[865] = data_i[865] & sel_one_hot_i[6];
  assign data_masked[864] = data_i[864] & sel_one_hot_i[6];
  assign data_masked[863] = data_i[863] & sel_one_hot_i[6];
  assign data_masked[862] = data_i[862] & sel_one_hot_i[6];
  assign data_masked[861] = data_i[861] & sel_one_hot_i[6];
  assign data_masked[860] = data_i[860] & sel_one_hot_i[6];
  assign data_masked[859] = data_i[859] & sel_one_hot_i[6];
  assign data_masked[858] = data_i[858] & sel_one_hot_i[6];
  assign data_masked[857] = data_i[857] & sel_one_hot_i[6];
  assign data_masked[856] = data_i[856] & sel_one_hot_i[6];
  assign data_masked[855] = data_i[855] & sel_one_hot_i[6];
  assign data_masked[854] = data_i[854] & sel_one_hot_i[6];
  assign data_masked[853] = data_i[853] & sel_one_hot_i[6];
  assign data_masked[852] = data_i[852] & sel_one_hot_i[6];
  assign data_masked[851] = data_i[851] & sel_one_hot_i[6];
  assign data_masked[850] = data_i[850] & sel_one_hot_i[6];
  assign data_masked[849] = data_i[849] & sel_one_hot_i[6];
  assign data_masked[848] = data_i[848] & sel_one_hot_i[6];
  assign data_masked[847] = data_i[847] & sel_one_hot_i[6];
  assign data_masked[846] = data_i[846] & sel_one_hot_i[6];
  assign data_masked[845] = data_i[845] & sel_one_hot_i[6];
  assign data_masked[844] = data_i[844] & sel_one_hot_i[6];
  assign data_masked[843] = data_i[843] & sel_one_hot_i[6];
  assign data_masked[842] = data_i[842] & sel_one_hot_i[6];
  assign data_masked[841] = data_i[841] & sel_one_hot_i[6];
  assign data_masked[840] = data_i[840] & sel_one_hot_i[6];
  assign data_masked[839] = data_i[839] & sel_one_hot_i[6];
  assign data_masked[838] = data_i[838] & sel_one_hot_i[6];
  assign data_masked[837] = data_i[837] & sel_one_hot_i[6];
  assign data_masked[836] = data_i[836] & sel_one_hot_i[6];
  assign data_masked[835] = data_i[835] & sel_one_hot_i[6];
  assign data_masked[834] = data_i[834] & sel_one_hot_i[6];
  assign data_masked[833] = data_i[833] & sel_one_hot_i[6];
  assign data_masked[832] = data_i[832] & sel_one_hot_i[6];
  assign data_masked[831] = data_i[831] & sel_one_hot_i[6];
  assign data_masked[830] = data_i[830] & sel_one_hot_i[6];
  assign data_masked[829] = data_i[829] & sel_one_hot_i[6];
  assign data_masked[828] = data_i[828] & sel_one_hot_i[6];
  assign data_masked[827] = data_i[827] & sel_one_hot_i[6];
  assign data_masked[826] = data_i[826] & sel_one_hot_i[6];
  assign data_masked[825] = data_i[825] & sel_one_hot_i[6];
  assign data_masked[824] = data_i[824] & sel_one_hot_i[6];
  assign data_masked[823] = data_i[823] & sel_one_hot_i[6];
  assign data_masked[822] = data_i[822] & sel_one_hot_i[6];
  assign data_masked[821] = data_i[821] & sel_one_hot_i[6];
  assign data_masked[820] = data_i[820] & sel_one_hot_i[6];
  assign data_masked[819] = data_i[819] & sel_one_hot_i[6];
  assign data_masked[818] = data_i[818] & sel_one_hot_i[6];
  assign data_masked[817] = data_i[817] & sel_one_hot_i[6];
  assign data_masked[816] = data_i[816] & sel_one_hot_i[6];
  assign data_masked[815] = data_i[815] & sel_one_hot_i[6];
  assign data_masked[814] = data_i[814] & sel_one_hot_i[6];
  assign data_masked[813] = data_i[813] & sel_one_hot_i[6];
  assign data_masked[812] = data_i[812] & sel_one_hot_i[6];
  assign data_masked[811] = data_i[811] & sel_one_hot_i[6];
  assign data_masked[810] = data_i[810] & sel_one_hot_i[6];
  assign data_masked[809] = data_i[809] & sel_one_hot_i[6];
  assign data_masked[808] = data_i[808] & sel_one_hot_i[6];
  assign data_masked[807] = data_i[807] & sel_one_hot_i[6];
  assign data_masked[806] = data_i[806] & sel_one_hot_i[6];
  assign data_masked[805] = data_i[805] & sel_one_hot_i[6];
  assign data_masked[804] = data_i[804] & sel_one_hot_i[6];
  assign data_masked[803] = data_i[803] & sel_one_hot_i[6];
  assign data_masked[802] = data_i[802] & sel_one_hot_i[6];
  assign data_masked[801] = data_i[801] & sel_one_hot_i[6];
  assign data_masked[800] = data_i[800] & sel_one_hot_i[6];
  assign data_masked[799] = data_i[799] & sel_one_hot_i[6];
  assign data_masked[798] = data_i[798] & sel_one_hot_i[6];
  assign data_masked[797] = data_i[797] & sel_one_hot_i[6];
  assign data_masked[796] = data_i[796] & sel_one_hot_i[6];
  assign data_masked[795] = data_i[795] & sel_one_hot_i[6];
  assign data_masked[794] = data_i[794] & sel_one_hot_i[6];
  assign data_masked[793] = data_i[793] & sel_one_hot_i[6];
  assign data_masked[792] = data_i[792] & sel_one_hot_i[6];
  assign data_masked[791] = data_i[791] & sel_one_hot_i[6];
  assign data_masked[790] = data_i[790] & sel_one_hot_i[6];
  assign data_masked[789] = data_i[789] & sel_one_hot_i[6];
  assign data_masked[788] = data_i[788] & sel_one_hot_i[6];
  assign data_masked[787] = data_i[787] & sel_one_hot_i[6];
  assign data_masked[786] = data_i[786] & sel_one_hot_i[6];
  assign data_masked[785] = data_i[785] & sel_one_hot_i[6];
  assign data_masked[784] = data_i[784] & sel_one_hot_i[6];
  assign data_masked[783] = data_i[783] & sel_one_hot_i[6];
  assign data_masked[782] = data_i[782] & sel_one_hot_i[6];
  assign data_masked[781] = data_i[781] & sel_one_hot_i[6];
  assign data_masked[780] = data_i[780] & sel_one_hot_i[6];
  assign data_masked[779] = data_i[779] & sel_one_hot_i[6];
  assign data_masked[778] = data_i[778] & sel_one_hot_i[6];
  assign data_masked[777] = data_i[777] & sel_one_hot_i[6];
  assign data_masked[776] = data_i[776] & sel_one_hot_i[6];
  assign data_masked[775] = data_i[775] & sel_one_hot_i[6];
  assign data_masked[774] = data_i[774] & sel_one_hot_i[6];
  assign data_masked[773] = data_i[773] & sel_one_hot_i[6];
  assign data_masked[772] = data_i[772] & sel_one_hot_i[6];
  assign data_masked[771] = data_i[771] & sel_one_hot_i[6];
  assign data_masked[770] = data_i[770] & sel_one_hot_i[6];
  assign data_masked[769] = data_i[769] & sel_one_hot_i[6];
  assign data_masked[768] = data_i[768] & sel_one_hot_i[6];
  assign data_masked[1023] = data_i[1023] & sel_one_hot_i[7];
  assign data_masked[1022] = data_i[1022] & sel_one_hot_i[7];
  assign data_masked[1021] = data_i[1021] & sel_one_hot_i[7];
  assign data_masked[1020] = data_i[1020] & sel_one_hot_i[7];
  assign data_masked[1019] = data_i[1019] & sel_one_hot_i[7];
  assign data_masked[1018] = data_i[1018] & sel_one_hot_i[7];
  assign data_masked[1017] = data_i[1017] & sel_one_hot_i[7];
  assign data_masked[1016] = data_i[1016] & sel_one_hot_i[7];
  assign data_masked[1015] = data_i[1015] & sel_one_hot_i[7];
  assign data_masked[1014] = data_i[1014] & sel_one_hot_i[7];
  assign data_masked[1013] = data_i[1013] & sel_one_hot_i[7];
  assign data_masked[1012] = data_i[1012] & sel_one_hot_i[7];
  assign data_masked[1011] = data_i[1011] & sel_one_hot_i[7];
  assign data_masked[1010] = data_i[1010] & sel_one_hot_i[7];
  assign data_masked[1009] = data_i[1009] & sel_one_hot_i[7];
  assign data_masked[1008] = data_i[1008] & sel_one_hot_i[7];
  assign data_masked[1007] = data_i[1007] & sel_one_hot_i[7];
  assign data_masked[1006] = data_i[1006] & sel_one_hot_i[7];
  assign data_masked[1005] = data_i[1005] & sel_one_hot_i[7];
  assign data_masked[1004] = data_i[1004] & sel_one_hot_i[7];
  assign data_masked[1003] = data_i[1003] & sel_one_hot_i[7];
  assign data_masked[1002] = data_i[1002] & sel_one_hot_i[7];
  assign data_masked[1001] = data_i[1001] & sel_one_hot_i[7];
  assign data_masked[1000] = data_i[1000] & sel_one_hot_i[7];
  assign data_masked[999] = data_i[999] & sel_one_hot_i[7];
  assign data_masked[998] = data_i[998] & sel_one_hot_i[7];
  assign data_masked[997] = data_i[997] & sel_one_hot_i[7];
  assign data_masked[996] = data_i[996] & sel_one_hot_i[7];
  assign data_masked[995] = data_i[995] & sel_one_hot_i[7];
  assign data_masked[994] = data_i[994] & sel_one_hot_i[7];
  assign data_masked[993] = data_i[993] & sel_one_hot_i[7];
  assign data_masked[992] = data_i[992] & sel_one_hot_i[7];
  assign data_masked[991] = data_i[991] & sel_one_hot_i[7];
  assign data_masked[990] = data_i[990] & sel_one_hot_i[7];
  assign data_masked[989] = data_i[989] & sel_one_hot_i[7];
  assign data_masked[988] = data_i[988] & sel_one_hot_i[7];
  assign data_masked[987] = data_i[987] & sel_one_hot_i[7];
  assign data_masked[986] = data_i[986] & sel_one_hot_i[7];
  assign data_masked[985] = data_i[985] & sel_one_hot_i[7];
  assign data_masked[984] = data_i[984] & sel_one_hot_i[7];
  assign data_masked[983] = data_i[983] & sel_one_hot_i[7];
  assign data_masked[982] = data_i[982] & sel_one_hot_i[7];
  assign data_masked[981] = data_i[981] & sel_one_hot_i[7];
  assign data_masked[980] = data_i[980] & sel_one_hot_i[7];
  assign data_masked[979] = data_i[979] & sel_one_hot_i[7];
  assign data_masked[978] = data_i[978] & sel_one_hot_i[7];
  assign data_masked[977] = data_i[977] & sel_one_hot_i[7];
  assign data_masked[976] = data_i[976] & sel_one_hot_i[7];
  assign data_masked[975] = data_i[975] & sel_one_hot_i[7];
  assign data_masked[974] = data_i[974] & sel_one_hot_i[7];
  assign data_masked[973] = data_i[973] & sel_one_hot_i[7];
  assign data_masked[972] = data_i[972] & sel_one_hot_i[7];
  assign data_masked[971] = data_i[971] & sel_one_hot_i[7];
  assign data_masked[970] = data_i[970] & sel_one_hot_i[7];
  assign data_masked[969] = data_i[969] & sel_one_hot_i[7];
  assign data_masked[968] = data_i[968] & sel_one_hot_i[7];
  assign data_masked[967] = data_i[967] & sel_one_hot_i[7];
  assign data_masked[966] = data_i[966] & sel_one_hot_i[7];
  assign data_masked[965] = data_i[965] & sel_one_hot_i[7];
  assign data_masked[964] = data_i[964] & sel_one_hot_i[7];
  assign data_masked[963] = data_i[963] & sel_one_hot_i[7];
  assign data_masked[962] = data_i[962] & sel_one_hot_i[7];
  assign data_masked[961] = data_i[961] & sel_one_hot_i[7];
  assign data_masked[960] = data_i[960] & sel_one_hot_i[7];
  assign data_masked[959] = data_i[959] & sel_one_hot_i[7];
  assign data_masked[958] = data_i[958] & sel_one_hot_i[7];
  assign data_masked[957] = data_i[957] & sel_one_hot_i[7];
  assign data_masked[956] = data_i[956] & sel_one_hot_i[7];
  assign data_masked[955] = data_i[955] & sel_one_hot_i[7];
  assign data_masked[954] = data_i[954] & sel_one_hot_i[7];
  assign data_masked[953] = data_i[953] & sel_one_hot_i[7];
  assign data_masked[952] = data_i[952] & sel_one_hot_i[7];
  assign data_masked[951] = data_i[951] & sel_one_hot_i[7];
  assign data_masked[950] = data_i[950] & sel_one_hot_i[7];
  assign data_masked[949] = data_i[949] & sel_one_hot_i[7];
  assign data_masked[948] = data_i[948] & sel_one_hot_i[7];
  assign data_masked[947] = data_i[947] & sel_one_hot_i[7];
  assign data_masked[946] = data_i[946] & sel_one_hot_i[7];
  assign data_masked[945] = data_i[945] & sel_one_hot_i[7];
  assign data_masked[944] = data_i[944] & sel_one_hot_i[7];
  assign data_masked[943] = data_i[943] & sel_one_hot_i[7];
  assign data_masked[942] = data_i[942] & sel_one_hot_i[7];
  assign data_masked[941] = data_i[941] & sel_one_hot_i[7];
  assign data_masked[940] = data_i[940] & sel_one_hot_i[7];
  assign data_masked[939] = data_i[939] & sel_one_hot_i[7];
  assign data_masked[938] = data_i[938] & sel_one_hot_i[7];
  assign data_masked[937] = data_i[937] & sel_one_hot_i[7];
  assign data_masked[936] = data_i[936] & sel_one_hot_i[7];
  assign data_masked[935] = data_i[935] & sel_one_hot_i[7];
  assign data_masked[934] = data_i[934] & sel_one_hot_i[7];
  assign data_masked[933] = data_i[933] & sel_one_hot_i[7];
  assign data_masked[932] = data_i[932] & sel_one_hot_i[7];
  assign data_masked[931] = data_i[931] & sel_one_hot_i[7];
  assign data_masked[930] = data_i[930] & sel_one_hot_i[7];
  assign data_masked[929] = data_i[929] & sel_one_hot_i[7];
  assign data_masked[928] = data_i[928] & sel_one_hot_i[7];
  assign data_masked[927] = data_i[927] & sel_one_hot_i[7];
  assign data_masked[926] = data_i[926] & sel_one_hot_i[7];
  assign data_masked[925] = data_i[925] & sel_one_hot_i[7];
  assign data_masked[924] = data_i[924] & sel_one_hot_i[7];
  assign data_masked[923] = data_i[923] & sel_one_hot_i[7];
  assign data_masked[922] = data_i[922] & sel_one_hot_i[7];
  assign data_masked[921] = data_i[921] & sel_one_hot_i[7];
  assign data_masked[920] = data_i[920] & sel_one_hot_i[7];
  assign data_masked[919] = data_i[919] & sel_one_hot_i[7];
  assign data_masked[918] = data_i[918] & sel_one_hot_i[7];
  assign data_masked[917] = data_i[917] & sel_one_hot_i[7];
  assign data_masked[916] = data_i[916] & sel_one_hot_i[7];
  assign data_masked[915] = data_i[915] & sel_one_hot_i[7];
  assign data_masked[914] = data_i[914] & sel_one_hot_i[7];
  assign data_masked[913] = data_i[913] & sel_one_hot_i[7];
  assign data_masked[912] = data_i[912] & sel_one_hot_i[7];
  assign data_masked[911] = data_i[911] & sel_one_hot_i[7];
  assign data_masked[910] = data_i[910] & sel_one_hot_i[7];
  assign data_masked[909] = data_i[909] & sel_one_hot_i[7];
  assign data_masked[908] = data_i[908] & sel_one_hot_i[7];
  assign data_masked[907] = data_i[907] & sel_one_hot_i[7];
  assign data_masked[906] = data_i[906] & sel_one_hot_i[7];
  assign data_masked[905] = data_i[905] & sel_one_hot_i[7];
  assign data_masked[904] = data_i[904] & sel_one_hot_i[7];
  assign data_masked[903] = data_i[903] & sel_one_hot_i[7];
  assign data_masked[902] = data_i[902] & sel_one_hot_i[7];
  assign data_masked[901] = data_i[901] & sel_one_hot_i[7];
  assign data_masked[900] = data_i[900] & sel_one_hot_i[7];
  assign data_masked[899] = data_i[899] & sel_one_hot_i[7];
  assign data_masked[898] = data_i[898] & sel_one_hot_i[7];
  assign data_masked[897] = data_i[897] & sel_one_hot_i[7];
  assign data_masked[896] = data_i[896] & sel_one_hot_i[7];
  assign data_masked[1151] = data_i[1151] & sel_one_hot_i[8];
  assign data_masked[1150] = data_i[1150] & sel_one_hot_i[8];
  assign data_masked[1149] = data_i[1149] & sel_one_hot_i[8];
  assign data_masked[1148] = data_i[1148] & sel_one_hot_i[8];
  assign data_masked[1147] = data_i[1147] & sel_one_hot_i[8];
  assign data_masked[1146] = data_i[1146] & sel_one_hot_i[8];
  assign data_masked[1145] = data_i[1145] & sel_one_hot_i[8];
  assign data_masked[1144] = data_i[1144] & sel_one_hot_i[8];
  assign data_masked[1143] = data_i[1143] & sel_one_hot_i[8];
  assign data_masked[1142] = data_i[1142] & sel_one_hot_i[8];
  assign data_masked[1141] = data_i[1141] & sel_one_hot_i[8];
  assign data_masked[1140] = data_i[1140] & sel_one_hot_i[8];
  assign data_masked[1139] = data_i[1139] & sel_one_hot_i[8];
  assign data_masked[1138] = data_i[1138] & sel_one_hot_i[8];
  assign data_masked[1137] = data_i[1137] & sel_one_hot_i[8];
  assign data_masked[1136] = data_i[1136] & sel_one_hot_i[8];
  assign data_masked[1135] = data_i[1135] & sel_one_hot_i[8];
  assign data_masked[1134] = data_i[1134] & sel_one_hot_i[8];
  assign data_masked[1133] = data_i[1133] & sel_one_hot_i[8];
  assign data_masked[1132] = data_i[1132] & sel_one_hot_i[8];
  assign data_masked[1131] = data_i[1131] & sel_one_hot_i[8];
  assign data_masked[1130] = data_i[1130] & sel_one_hot_i[8];
  assign data_masked[1129] = data_i[1129] & sel_one_hot_i[8];
  assign data_masked[1128] = data_i[1128] & sel_one_hot_i[8];
  assign data_masked[1127] = data_i[1127] & sel_one_hot_i[8];
  assign data_masked[1126] = data_i[1126] & sel_one_hot_i[8];
  assign data_masked[1125] = data_i[1125] & sel_one_hot_i[8];
  assign data_masked[1124] = data_i[1124] & sel_one_hot_i[8];
  assign data_masked[1123] = data_i[1123] & sel_one_hot_i[8];
  assign data_masked[1122] = data_i[1122] & sel_one_hot_i[8];
  assign data_masked[1121] = data_i[1121] & sel_one_hot_i[8];
  assign data_masked[1120] = data_i[1120] & sel_one_hot_i[8];
  assign data_masked[1119] = data_i[1119] & sel_one_hot_i[8];
  assign data_masked[1118] = data_i[1118] & sel_one_hot_i[8];
  assign data_masked[1117] = data_i[1117] & sel_one_hot_i[8];
  assign data_masked[1116] = data_i[1116] & sel_one_hot_i[8];
  assign data_masked[1115] = data_i[1115] & sel_one_hot_i[8];
  assign data_masked[1114] = data_i[1114] & sel_one_hot_i[8];
  assign data_masked[1113] = data_i[1113] & sel_one_hot_i[8];
  assign data_masked[1112] = data_i[1112] & sel_one_hot_i[8];
  assign data_masked[1111] = data_i[1111] & sel_one_hot_i[8];
  assign data_masked[1110] = data_i[1110] & sel_one_hot_i[8];
  assign data_masked[1109] = data_i[1109] & sel_one_hot_i[8];
  assign data_masked[1108] = data_i[1108] & sel_one_hot_i[8];
  assign data_masked[1107] = data_i[1107] & sel_one_hot_i[8];
  assign data_masked[1106] = data_i[1106] & sel_one_hot_i[8];
  assign data_masked[1105] = data_i[1105] & sel_one_hot_i[8];
  assign data_masked[1104] = data_i[1104] & sel_one_hot_i[8];
  assign data_masked[1103] = data_i[1103] & sel_one_hot_i[8];
  assign data_masked[1102] = data_i[1102] & sel_one_hot_i[8];
  assign data_masked[1101] = data_i[1101] & sel_one_hot_i[8];
  assign data_masked[1100] = data_i[1100] & sel_one_hot_i[8];
  assign data_masked[1099] = data_i[1099] & sel_one_hot_i[8];
  assign data_masked[1098] = data_i[1098] & sel_one_hot_i[8];
  assign data_masked[1097] = data_i[1097] & sel_one_hot_i[8];
  assign data_masked[1096] = data_i[1096] & sel_one_hot_i[8];
  assign data_masked[1095] = data_i[1095] & sel_one_hot_i[8];
  assign data_masked[1094] = data_i[1094] & sel_one_hot_i[8];
  assign data_masked[1093] = data_i[1093] & sel_one_hot_i[8];
  assign data_masked[1092] = data_i[1092] & sel_one_hot_i[8];
  assign data_masked[1091] = data_i[1091] & sel_one_hot_i[8];
  assign data_masked[1090] = data_i[1090] & sel_one_hot_i[8];
  assign data_masked[1089] = data_i[1089] & sel_one_hot_i[8];
  assign data_masked[1088] = data_i[1088] & sel_one_hot_i[8];
  assign data_masked[1087] = data_i[1087] & sel_one_hot_i[8];
  assign data_masked[1086] = data_i[1086] & sel_one_hot_i[8];
  assign data_masked[1085] = data_i[1085] & sel_one_hot_i[8];
  assign data_masked[1084] = data_i[1084] & sel_one_hot_i[8];
  assign data_masked[1083] = data_i[1083] & sel_one_hot_i[8];
  assign data_masked[1082] = data_i[1082] & sel_one_hot_i[8];
  assign data_masked[1081] = data_i[1081] & sel_one_hot_i[8];
  assign data_masked[1080] = data_i[1080] & sel_one_hot_i[8];
  assign data_masked[1079] = data_i[1079] & sel_one_hot_i[8];
  assign data_masked[1078] = data_i[1078] & sel_one_hot_i[8];
  assign data_masked[1077] = data_i[1077] & sel_one_hot_i[8];
  assign data_masked[1076] = data_i[1076] & sel_one_hot_i[8];
  assign data_masked[1075] = data_i[1075] & sel_one_hot_i[8];
  assign data_masked[1074] = data_i[1074] & sel_one_hot_i[8];
  assign data_masked[1073] = data_i[1073] & sel_one_hot_i[8];
  assign data_masked[1072] = data_i[1072] & sel_one_hot_i[8];
  assign data_masked[1071] = data_i[1071] & sel_one_hot_i[8];
  assign data_masked[1070] = data_i[1070] & sel_one_hot_i[8];
  assign data_masked[1069] = data_i[1069] & sel_one_hot_i[8];
  assign data_masked[1068] = data_i[1068] & sel_one_hot_i[8];
  assign data_masked[1067] = data_i[1067] & sel_one_hot_i[8];
  assign data_masked[1066] = data_i[1066] & sel_one_hot_i[8];
  assign data_masked[1065] = data_i[1065] & sel_one_hot_i[8];
  assign data_masked[1064] = data_i[1064] & sel_one_hot_i[8];
  assign data_masked[1063] = data_i[1063] & sel_one_hot_i[8];
  assign data_masked[1062] = data_i[1062] & sel_one_hot_i[8];
  assign data_masked[1061] = data_i[1061] & sel_one_hot_i[8];
  assign data_masked[1060] = data_i[1060] & sel_one_hot_i[8];
  assign data_masked[1059] = data_i[1059] & sel_one_hot_i[8];
  assign data_masked[1058] = data_i[1058] & sel_one_hot_i[8];
  assign data_masked[1057] = data_i[1057] & sel_one_hot_i[8];
  assign data_masked[1056] = data_i[1056] & sel_one_hot_i[8];
  assign data_masked[1055] = data_i[1055] & sel_one_hot_i[8];
  assign data_masked[1054] = data_i[1054] & sel_one_hot_i[8];
  assign data_masked[1053] = data_i[1053] & sel_one_hot_i[8];
  assign data_masked[1052] = data_i[1052] & sel_one_hot_i[8];
  assign data_masked[1051] = data_i[1051] & sel_one_hot_i[8];
  assign data_masked[1050] = data_i[1050] & sel_one_hot_i[8];
  assign data_masked[1049] = data_i[1049] & sel_one_hot_i[8];
  assign data_masked[1048] = data_i[1048] & sel_one_hot_i[8];
  assign data_masked[1047] = data_i[1047] & sel_one_hot_i[8];
  assign data_masked[1046] = data_i[1046] & sel_one_hot_i[8];
  assign data_masked[1045] = data_i[1045] & sel_one_hot_i[8];
  assign data_masked[1044] = data_i[1044] & sel_one_hot_i[8];
  assign data_masked[1043] = data_i[1043] & sel_one_hot_i[8];
  assign data_masked[1042] = data_i[1042] & sel_one_hot_i[8];
  assign data_masked[1041] = data_i[1041] & sel_one_hot_i[8];
  assign data_masked[1040] = data_i[1040] & sel_one_hot_i[8];
  assign data_masked[1039] = data_i[1039] & sel_one_hot_i[8];
  assign data_masked[1038] = data_i[1038] & sel_one_hot_i[8];
  assign data_masked[1037] = data_i[1037] & sel_one_hot_i[8];
  assign data_masked[1036] = data_i[1036] & sel_one_hot_i[8];
  assign data_masked[1035] = data_i[1035] & sel_one_hot_i[8];
  assign data_masked[1034] = data_i[1034] & sel_one_hot_i[8];
  assign data_masked[1033] = data_i[1033] & sel_one_hot_i[8];
  assign data_masked[1032] = data_i[1032] & sel_one_hot_i[8];
  assign data_masked[1031] = data_i[1031] & sel_one_hot_i[8];
  assign data_masked[1030] = data_i[1030] & sel_one_hot_i[8];
  assign data_masked[1029] = data_i[1029] & sel_one_hot_i[8];
  assign data_masked[1028] = data_i[1028] & sel_one_hot_i[8];
  assign data_masked[1027] = data_i[1027] & sel_one_hot_i[8];
  assign data_masked[1026] = data_i[1026] & sel_one_hot_i[8];
  assign data_masked[1025] = data_i[1025] & sel_one_hot_i[8];
  assign data_masked[1024] = data_i[1024] & sel_one_hot_i[8];
  assign data_masked[1279] = data_i[1279] & sel_one_hot_i[9];
  assign data_masked[1278] = data_i[1278] & sel_one_hot_i[9];
  assign data_masked[1277] = data_i[1277] & sel_one_hot_i[9];
  assign data_masked[1276] = data_i[1276] & sel_one_hot_i[9];
  assign data_masked[1275] = data_i[1275] & sel_one_hot_i[9];
  assign data_masked[1274] = data_i[1274] & sel_one_hot_i[9];
  assign data_masked[1273] = data_i[1273] & sel_one_hot_i[9];
  assign data_masked[1272] = data_i[1272] & sel_one_hot_i[9];
  assign data_masked[1271] = data_i[1271] & sel_one_hot_i[9];
  assign data_masked[1270] = data_i[1270] & sel_one_hot_i[9];
  assign data_masked[1269] = data_i[1269] & sel_one_hot_i[9];
  assign data_masked[1268] = data_i[1268] & sel_one_hot_i[9];
  assign data_masked[1267] = data_i[1267] & sel_one_hot_i[9];
  assign data_masked[1266] = data_i[1266] & sel_one_hot_i[9];
  assign data_masked[1265] = data_i[1265] & sel_one_hot_i[9];
  assign data_masked[1264] = data_i[1264] & sel_one_hot_i[9];
  assign data_masked[1263] = data_i[1263] & sel_one_hot_i[9];
  assign data_masked[1262] = data_i[1262] & sel_one_hot_i[9];
  assign data_masked[1261] = data_i[1261] & sel_one_hot_i[9];
  assign data_masked[1260] = data_i[1260] & sel_one_hot_i[9];
  assign data_masked[1259] = data_i[1259] & sel_one_hot_i[9];
  assign data_masked[1258] = data_i[1258] & sel_one_hot_i[9];
  assign data_masked[1257] = data_i[1257] & sel_one_hot_i[9];
  assign data_masked[1256] = data_i[1256] & sel_one_hot_i[9];
  assign data_masked[1255] = data_i[1255] & sel_one_hot_i[9];
  assign data_masked[1254] = data_i[1254] & sel_one_hot_i[9];
  assign data_masked[1253] = data_i[1253] & sel_one_hot_i[9];
  assign data_masked[1252] = data_i[1252] & sel_one_hot_i[9];
  assign data_masked[1251] = data_i[1251] & sel_one_hot_i[9];
  assign data_masked[1250] = data_i[1250] & sel_one_hot_i[9];
  assign data_masked[1249] = data_i[1249] & sel_one_hot_i[9];
  assign data_masked[1248] = data_i[1248] & sel_one_hot_i[9];
  assign data_masked[1247] = data_i[1247] & sel_one_hot_i[9];
  assign data_masked[1246] = data_i[1246] & sel_one_hot_i[9];
  assign data_masked[1245] = data_i[1245] & sel_one_hot_i[9];
  assign data_masked[1244] = data_i[1244] & sel_one_hot_i[9];
  assign data_masked[1243] = data_i[1243] & sel_one_hot_i[9];
  assign data_masked[1242] = data_i[1242] & sel_one_hot_i[9];
  assign data_masked[1241] = data_i[1241] & sel_one_hot_i[9];
  assign data_masked[1240] = data_i[1240] & sel_one_hot_i[9];
  assign data_masked[1239] = data_i[1239] & sel_one_hot_i[9];
  assign data_masked[1238] = data_i[1238] & sel_one_hot_i[9];
  assign data_masked[1237] = data_i[1237] & sel_one_hot_i[9];
  assign data_masked[1236] = data_i[1236] & sel_one_hot_i[9];
  assign data_masked[1235] = data_i[1235] & sel_one_hot_i[9];
  assign data_masked[1234] = data_i[1234] & sel_one_hot_i[9];
  assign data_masked[1233] = data_i[1233] & sel_one_hot_i[9];
  assign data_masked[1232] = data_i[1232] & sel_one_hot_i[9];
  assign data_masked[1231] = data_i[1231] & sel_one_hot_i[9];
  assign data_masked[1230] = data_i[1230] & sel_one_hot_i[9];
  assign data_masked[1229] = data_i[1229] & sel_one_hot_i[9];
  assign data_masked[1228] = data_i[1228] & sel_one_hot_i[9];
  assign data_masked[1227] = data_i[1227] & sel_one_hot_i[9];
  assign data_masked[1226] = data_i[1226] & sel_one_hot_i[9];
  assign data_masked[1225] = data_i[1225] & sel_one_hot_i[9];
  assign data_masked[1224] = data_i[1224] & sel_one_hot_i[9];
  assign data_masked[1223] = data_i[1223] & sel_one_hot_i[9];
  assign data_masked[1222] = data_i[1222] & sel_one_hot_i[9];
  assign data_masked[1221] = data_i[1221] & sel_one_hot_i[9];
  assign data_masked[1220] = data_i[1220] & sel_one_hot_i[9];
  assign data_masked[1219] = data_i[1219] & sel_one_hot_i[9];
  assign data_masked[1218] = data_i[1218] & sel_one_hot_i[9];
  assign data_masked[1217] = data_i[1217] & sel_one_hot_i[9];
  assign data_masked[1216] = data_i[1216] & sel_one_hot_i[9];
  assign data_masked[1215] = data_i[1215] & sel_one_hot_i[9];
  assign data_masked[1214] = data_i[1214] & sel_one_hot_i[9];
  assign data_masked[1213] = data_i[1213] & sel_one_hot_i[9];
  assign data_masked[1212] = data_i[1212] & sel_one_hot_i[9];
  assign data_masked[1211] = data_i[1211] & sel_one_hot_i[9];
  assign data_masked[1210] = data_i[1210] & sel_one_hot_i[9];
  assign data_masked[1209] = data_i[1209] & sel_one_hot_i[9];
  assign data_masked[1208] = data_i[1208] & sel_one_hot_i[9];
  assign data_masked[1207] = data_i[1207] & sel_one_hot_i[9];
  assign data_masked[1206] = data_i[1206] & sel_one_hot_i[9];
  assign data_masked[1205] = data_i[1205] & sel_one_hot_i[9];
  assign data_masked[1204] = data_i[1204] & sel_one_hot_i[9];
  assign data_masked[1203] = data_i[1203] & sel_one_hot_i[9];
  assign data_masked[1202] = data_i[1202] & sel_one_hot_i[9];
  assign data_masked[1201] = data_i[1201] & sel_one_hot_i[9];
  assign data_masked[1200] = data_i[1200] & sel_one_hot_i[9];
  assign data_masked[1199] = data_i[1199] & sel_one_hot_i[9];
  assign data_masked[1198] = data_i[1198] & sel_one_hot_i[9];
  assign data_masked[1197] = data_i[1197] & sel_one_hot_i[9];
  assign data_masked[1196] = data_i[1196] & sel_one_hot_i[9];
  assign data_masked[1195] = data_i[1195] & sel_one_hot_i[9];
  assign data_masked[1194] = data_i[1194] & sel_one_hot_i[9];
  assign data_masked[1193] = data_i[1193] & sel_one_hot_i[9];
  assign data_masked[1192] = data_i[1192] & sel_one_hot_i[9];
  assign data_masked[1191] = data_i[1191] & sel_one_hot_i[9];
  assign data_masked[1190] = data_i[1190] & sel_one_hot_i[9];
  assign data_masked[1189] = data_i[1189] & sel_one_hot_i[9];
  assign data_masked[1188] = data_i[1188] & sel_one_hot_i[9];
  assign data_masked[1187] = data_i[1187] & sel_one_hot_i[9];
  assign data_masked[1186] = data_i[1186] & sel_one_hot_i[9];
  assign data_masked[1185] = data_i[1185] & sel_one_hot_i[9];
  assign data_masked[1184] = data_i[1184] & sel_one_hot_i[9];
  assign data_masked[1183] = data_i[1183] & sel_one_hot_i[9];
  assign data_masked[1182] = data_i[1182] & sel_one_hot_i[9];
  assign data_masked[1181] = data_i[1181] & sel_one_hot_i[9];
  assign data_masked[1180] = data_i[1180] & sel_one_hot_i[9];
  assign data_masked[1179] = data_i[1179] & sel_one_hot_i[9];
  assign data_masked[1178] = data_i[1178] & sel_one_hot_i[9];
  assign data_masked[1177] = data_i[1177] & sel_one_hot_i[9];
  assign data_masked[1176] = data_i[1176] & sel_one_hot_i[9];
  assign data_masked[1175] = data_i[1175] & sel_one_hot_i[9];
  assign data_masked[1174] = data_i[1174] & sel_one_hot_i[9];
  assign data_masked[1173] = data_i[1173] & sel_one_hot_i[9];
  assign data_masked[1172] = data_i[1172] & sel_one_hot_i[9];
  assign data_masked[1171] = data_i[1171] & sel_one_hot_i[9];
  assign data_masked[1170] = data_i[1170] & sel_one_hot_i[9];
  assign data_masked[1169] = data_i[1169] & sel_one_hot_i[9];
  assign data_masked[1168] = data_i[1168] & sel_one_hot_i[9];
  assign data_masked[1167] = data_i[1167] & sel_one_hot_i[9];
  assign data_masked[1166] = data_i[1166] & sel_one_hot_i[9];
  assign data_masked[1165] = data_i[1165] & sel_one_hot_i[9];
  assign data_masked[1164] = data_i[1164] & sel_one_hot_i[9];
  assign data_masked[1163] = data_i[1163] & sel_one_hot_i[9];
  assign data_masked[1162] = data_i[1162] & sel_one_hot_i[9];
  assign data_masked[1161] = data_i[1161] & sel_one_hot_i[9];
  assign data_masked[1160] = data_i[1160] & sel_one_hot_i[9];
  assign data_masked[1159] = data_i[1159] & sel_one_hot_i[9];
  assign data_masked[1158] = data_i[1158] & sel_one_hot_i[9];
  assign data_masked[1157] = data_i[1157] & sel_one_hot_i[9];
  assign data_masked[1156] = data_i[1156] & sel_one_hot_i[9];
  assign data_masked[1155] = data_i[1155] & sel_one_hot_i[9];
  assign data_masked[1154] = data_i[1154] & sel_one_hot_i[9];
  assign data_masked[1153] = data_i[1153] & sel_one_hot_i[9];
  assign data_masked[1152] = data_i[1152] & sel_one_hot_i[9];
  assign data_masked[1407] = data_i[1407] & sel_one_hot_i[10];
  assign data_masked[1406] = data_i[1406] & sel_one_hot_i[10];
  assign data_masked[1405] = data_i[1405] & sel_one_hot_i[10];
  assign data_masked[1404] = data_i[1404] & sel_one_hot_i[10];
  assign data_masked[1403] = data_i[1403] & sel_one_hot_i[10];
  assign data_masked[1402] = data_i[1402] & sel_one_hot_i[10];
  assign data_masked[1401] = data_i[1401] & sel_one_hot_i[10];
  assign data_masked[1400] = data_i[1400] & sel_one_hot_i[10];
  assign data_masked[1399] = data_i[1399] & sel_one_hot_i[10];
  assign data_masked[1398] = data_i[1398] & sel_one_hot_i[10];
  assign data_masked[1397] = data_i[1397] & sel_one_hot_i[10];
  assign data_masked[1396] = data_i[1396] & sel_one_hot_i[10];
  assign data_masked[1395] = data_i[1395] & sel_one_hot_i[10];
  assign data_masked[1394] = data_i[1394] & sel_one_hot_i[10];
  assign data_masked[1393] = data_i[1393] & sel_one_hot_i[10];
  assign data_masked[1392] = data_i[1392] & sel_one_hot_i[10];
  assign data_masked[1391] = data_i[1391] & sel_one_hot_i[10];
  assign data_masked[1390] = data_i[1390] & sel_one_hot_i[10];
  assign data_masked[1389] = data_i[1389] & sel_one_hot_i[10];
  assign data_masked[1388] = data_i[1388] & sel_one_hot_i[10];
  assign data_masked[1387] = data_i[1387] & sel_one_hot_i[10];
  assign data_masked[1386] = data_i[1386] & sel_one_hot_i[10];
  assign data_masked[1385] = data_i[1385] & sel_one_hot_i[10];
  assign data_masked[1384] = data_i[1384] & sel_one_hot_i[10];
  assign data_masked[1383] = data_i[1383] & sel_one_hot_i[10];
  assign data_masked[1382] = data_i[1382] & sel_one_hot_i[10];
  assign data_masked[1381] = data_i[1381] & sel_one_hot_i[10];
  assign data_masked[1380] = data_i[1380] & sel_one_hot_i[10];
  assign data_masked[1379] = data_i[1379] & sel_one_hot_i[10];
  assign data_masked[1378] = data_i[1378] & sel_one_hot_i[10];
  assign data_masked[1377] = data_i[1377] & sel_one_hot_i[10];
  assign data_masked[1376] = data_i[1376] & sel_one_hot_i[10];
  assign data_masked[1375] = data_i[1375] & sel_one_hot_i[10];
  assign data_masked[1374] = data_i[1374] & sel_one_hot_i[10];
  assign data_masked[1373] = data_i[1373] & sel_one_hot_i[10];
  assign data_masked[1372] = data_i[1372] & sel_one_hot_i[10];
  assign data_masked[1371] = data_i[1371] & sel_one_hot_i[10];
  assign data_masked[1370] = data_i[1370] & sel_one_hot_i[10];
  assign data_masked[1369] = data_i[1369] & sel_one_hot_i[10];
  assign data_masked[1368] = data_i[1368] & sel_one_hot_i[10];
  assign data_masked[1367] = data_i[1367] & sel_one_hot_i[10];
  assign data_masked[1366] = data_i[1366] & sel_one_hot_i[10];
  assign data_masked[1365] = data_i[1365] & sel_one_hot_i[10];
  assign data_masked[1364] = data_i[1364] & sel_one_hot_i[10];
  assign data_masked[1363] = data_i[1363] & sel_one_hot_i[10];
  assign data_masked[1362] = data_i[1362] & sel_one_hot_i[10];
  assign data_masked[1361] = data_i[1361] & sel_one_hot_i[10];
  assign data_masked[1360] = data_i[1360] & sel_one_hot_i[10];
  assign data_masked[1359] = data_i[1359] & sel_one_hot_i[10];
  assign data_masked[1358] = data_i[1358] & sel_one_hot_i[10];
  assign data_masked[1357] = data_i[1357] & sel_one_hot_i[10];
  assign data_masked[1356] = data_i[1356] & sel_one_hot_i[10];
  assign data_masked[1355] = data_i[1355] & sel_one_hot_i[10];
  assign data_masked[1354] = data_i[1354] & sel_one_hot_i[10];
  assign data_masked[1353] = data_i[1353] & sel_one_hot_i[10];
  assign data_masked[1352] = data_i[1352] & sel_one_hot_i[10];
  assign data_masked[1351] = data_i[1351] & sel_one_hot_i[10];
  assign data_masked[1350] = data_i[1350] & sel_one_hot_i[10];
  assign data_masked[1349] = data_i[1349] & sel_one_hot_i[10];
  assign data_masked[1348] = data_i[1348] & sel_one_hot_i[10];
  assign data_masked[1347] = data_i[1347] & sel_one_hot_i[10];
  assign data_masked[1346] = data_i[1346] & sel_one_hot_i[10];
  assign data_masked[1345] = data_i[1345] & sel_one_hot_i[10];
  assign data_masked[1344] = data_i[1344] & sel_one_hot_i[10];
  assign data_masked[1343] = data_i[1343] & sel_one_hot_i[10];
  assign data_masked[1342] = data_i[1342] & sel_one_hot_i[10];
  assign data_masked[1341] = data_i[1341] & sel_one_hot_i[10];
  assign data_masked[1340] = data_i[1340] & sel_one_hot_i[10];
  assign data_masked[1339] = data_i[1339] & sel_one_hot_i[10];
  assign data_masked[1338] = data_i[1338] & sel_one_hot_i[10];
  assign data_masked[1337] = data_i[1337] & sel_one_hot_i[10];
  assign data_masked[1336] = data_i[1336] & sel_one_hot_i[10];
  assign data_masked[1335] = data_i[1335] & sel_one_hot_i[10];
  assign data_masked[1334] = data_i[1334] & sel_one_hot_i[10];
  assign data_masked[1333] = data_i[1333] & sel_one_hot_i[10];
  assign data_masked[1332] = data_i[1332] & sel_one_hot_i[10];
  assign data_masked[1331] = data_i[1331] & sel_one_hot_i[10];
  assign data_masked[1330] = data_i[1330] & sel_one_hot_i[10];
  assign data_masked[1329] = data_i[1329] & sel_one_hot_i[10];
  assign data_masked[1328] = data_i[1328] & sel_one_hot_i[10];
  assign data_masked[1327] = data_i[1327] & sel_one_hot_i[10];
  assign data_masked[1326] = data_i[1326] & sel_one_hot_i[10];
  assign data_masked[1325] = data_i[1325] & sel_one_hot_i[10];
  assign data_masked[1324] = data_i[1324] & sel_one_hot_i[10];
  assign data_masked[1323] = data_i[1323] & sel_one_hot_i[10];
  assign data_masked[1322] = data_i[1322] & sel_one_hot_i[10];
  assign data_masked[1321] = data_i[1321] & sel_one_hot_i[10];
  assign data_masked[1320] = data_i[1320] & sel_one_hot_i[10];
  assign data_masked[1319] = data_i[1319] & sel_one_hot_i[10];
  assign data_masked[1318] = data_i[1318] & sel_one_hot_i[10];
  assign data_masked[1317] = data_i[1317] & sel_one_hot_i[10];
  assign data_masked[1316] = data_i[1316] & sel_one_hot_i[10];
  assign data_masked[1315] = data_i[1315] & sel_one_hot_i[10];
  assign data_masked[1314] = data_i[1314] & sel_one_hot_i[10];
  assign data_masked[1313] = data_i[1313] & sel_one_hot_i[10];
  assign data_masked[1312] = data_i[1312] & sel_one_hot_i[10];
  assign data_masked[1311] = data_i[1311] & sel_one_hot_i[10];
  assign data_masked[1310] = data_i[1310] & sel_one_hot_i[10];
  assign data_masked[1309] = data_i[1309] & sel_one_hot_i[10];
  assign data_masked[1308] = data_i[1308] & sel_one_hot_i[10];
  assign data_masked[1307] = data_i[1307] & sel_one_hot_i[10];
  assign data_masked[1306] = data_i[1306] & sel_one_hot_i[10];
  assign data_masked[1305] = data_i[1305] & sel_one_hot_i[10];
  assign data_masked[1304] = data_i[1304] & sel_one_hot_i[10];
  assign data_masked[1303] = data_i[1303] & sel_one_hot_i[10];
  assign data_masked[1302] = data_i[1302] & sel_one_hot_i[10];
  assign data_masked[1301] = data_i[1301] & sel_one_hot_i[10];
  assign data_masked[1300] = data_i[1300] & sel_one_hot_i[10];
  assign data_masked[1299] = data_i[1299] & sel_one_hot_i[10];
  assign data_masked[1298] = data_i[1298] & sel_one_hot_i[10];
  assign data_masked[1297] = data_i[1297] & sel_one_hot_i[10];
  assign data_masked[1296] = data_i[1296] & sel_one_hot_i[10];
  assign data_masked[1295] = data_i[1295] & sel_one_hot_i[10];
  assign data_masked[1294] = data_i[1294] & sel_one_hot_i[10];
  assign data_masked[1293] = data_i[1293] & sel_one_hot_i[10];
  assign data_masked[1292] = data_i[1292] & sel_one_hot_i[10];
  assign data_masked[1291] = data_i[1291] & sel_one_hot_i[10];
  assign data_masked[1290] = data_i[1290] & sel_one_hot_i[10];
  assign data_masked[1289] = data_i[1289] & sel_one_hot_i[10];
  assign data_masked[1288] = data_i[1288] & sel_one_hot_i[10];
  assign data_masked[1287] = data_i[1287] & sel_one_hot_i[10];
  assign data_masked[1286] = data_i[1286] & sel_one_hot_i[10];
  assign data_masked[1285] = data_i[1285] & sel_one_hot_i[10];
  assign data_masked[1284] = data_i[1284] & sel_one_hot_i[10];
  assign data_masked[1283] = data_i[1283] & sel_one_hot_i[10];
  assign data_masked[1282] = data_i[1282] & sel_one_hot_i[10];
  assign data_masked[1281] = data_i[1281] & sel_one_hot_i[10];
  assign data_masked[1280] = data_i[1280] & sel_one_hot_i[10];
  assign data_masked[1535] = data_i[1535] & sel_one_hot_i[11];
  assign data_masked[1534] = data_i[1534] & sel_one_hot_i[11];
  assign data_masked[1533] = data_i[1533] & sel_one_hot_i[11];
  assign data_masked[1532] = data_i[1532] & sel_one_hot_i[11];
  assign data_masked[1531] = data_i[1531] & sel_one_hot_i[11];
  assign data_masked[1530] = data_i[1530] & sel_one_hot_i[11];
  assign data_masked[1529] = data_i[1529] & sel_one_hot_i[11];
  assign data_masked[1528] = data_i[1528] & sel_one_hot_i[11];
  assign data_masked[1527] = data_i[1527] & sel_one_hot_i[11];
  assign data_masked[1526] = data_i[1526] & sel_one_hot_i[11];
  assign data_masked[1525] = data_i[1525] & sel_one_hot_i[11];
  assign data_masked[1524] = data_i[1524] & sel_one_hot_i[11];
  assign data_masked[1523] = data_i[1523] & sel_one_hot_i[11];
  assign data_masked[1522] = data_i[1522] & sel_one_hot_i[11];
  assign data_masked[1521] = data_i[1521] & sel_one_hot_i[11];
  assign data_masked[1520] = data_i[1520] & sel_one_hot_i[11];
  assign data_masked[1519] = data_i[1519] & sel_one_hot_i[11];
  assign data_masked[1518] = data_i[1518] & sel_one_hot_i[11];
  assign data_masked[1517] = data_i[1517] & sel_one_hot_i[11];
  assign data_masked[1516] = data_i[1516] & sel_one_hot_i[11];
  assign data_masked[1515] = data_i[1515] & sel_one_hot_i[11];
  assign data_masked[1514] = data_i[1514] & sel_one_hot_i[11];
  assign data_masked[1513] = data_i[1513] & sel_one_hot_i[11];
  assign data_masked[1512] = data_i[1512] & sel_one_hot_i[11];
  assign data_masked[1511] = data_i[1511] & sel_one_hot_i[11];
  assign data_masked[1510] = data_i[1510] & sel_one_hot_i[11];
  assign data_masked[1509] = data_i[1509] & sel_one_hot_i[11];
  assign data_masked[1508] = data_i[1508] & sel_one_hot_i[11];
  assign data_masked[1507] = data_i[1507] & sel_one_hot_i[11];
  assign data_masked[1506] = data_i[1506] & sel_one_hot_i[11];
  assign data_masked[1505] = data_i[1505] & sel_one_hot_i[11];
  assign data_masked[1504] = data_i[1504] & sel_one_hot_i[11];
  assign data_masked[1503] = data_i[1503] & sel_one_hot_i[11];
  assign data_masked[1502] = data_i[1502] & sel_one_hot_i[11];
  assign data_masked[1501] = data_i[1501] & sel_one_hot_i[11];
  assign data_masked[1500] = data_i[1500] & sel_one_hot_i[11];
  assign data_masked[1499] = data_i[1499] & sel_one_hot_i[11];
  assign data_masked[1498] = data_i[1498] & sel_one_hot_i[11];
  assign data_masked[1497] = data_i[1497] & sel_one_hot_i[11];
  assign data_masked[1496] = data_i[1496] & sel_one_hot_i[11];
  assign data_masked[1495] = data_i[1495] & sel_one_hot_i[11];
  assign data_masked[1494] = data_i[1494] & sel_one_hot_i[11];
  assign data_masked[1493] = data_i[1493] & sel_one_hot_i[11];
  assign data_masked[1492] = data_i[1492] & sel_one_hot_i[11];
  assign data_masked[1491] = data_i[1491] & sel_one_hot_i[11];
  assign data_masked[1490] = data_i[1490] & sel_one_hot_i[11];
  assign data_masked[1489] = data_i[1489] & sel_one_hot_i[11];
  assign data_masked[1488] = data_i[1488] & sel_one_hot_i[11];
  assign data_masked[1487] = data_i[1487] & sel_one_hot_i[11];
  assign data_masked[1486] = data_i[1486] & sel_one_hot_i[11];
  assign data_masked[1485] = data_i[1485] & sel_one_hot_i[11];
  assign data_masked[1484] = data_i[1484] & sel_one_hot_i[11];
  assign data_masked[1483] = data_i[1483] & sel_one_hot_i[11];
  assign data_masked[1482] = data_i[1482] & sel_one_hot_i[11];
  assign data_masked[1481] = data_i[1481] & sel_one_hot_i[11];
  assign data_masked[1480] = data_i[1480] & sel_one_hot_i[11];
  assign data_masked[1479] = data_i[1479] & sel_one_hot_i[11];
  assign data_masked[1478] = data_i[1478] & sel_one_hot_i[11];
  assign data_masked[1477] = data_i[1477] & sel_one_hot_i[11];
  assign data_masked[1476] = data_i[1476] & sel_one_hot_i[11];
  assign data_masked[1475] = data_i[1475] & sel_one_hot_i[11];
  assign data_masked[1474] = data_i[1474] & sel_one_hot_i[11];
  assign data_masked[1473] = data_i[1473] & sel_one_hot_i[11];
  assign data_masked[1472] = data_i[1472] & sel_one_hot_i[11];
  assign data_masked[1471] = data_i[1471] & sel_one_hot_i[11];
  assign data_masked[1470] = data_i[1470] & sel_one_hot_i[11];
  assign data_masked[1469] = data_i[1469] & sel_one_hot_i[11];
  assign data_masked[1468] = data_i[1468] & sel_one_hot_i[11];
  assign data_masked[1467] = data_i[1467] & sel_one_hot_i[11];
  assign data_masked[1466] = data_i[1466] & sel_one_hot_i[11];
  assign data_masked[1465] = data_i[1465] & sel_one_hot_i[11];
  assign data_masked[1464] = data_i[1464] & sel_one_hot_i[11];
  assign data_masked[1463] = data_i[1463] & sel_one_hot_i[11];
  assign data_masked[1462] = data_i[1462] & sel_one_hot_i[11];
  assign data_masked[1461] = data_i[1461] & sel_one_hot_i[11];
  assign data_masked[1460] = data_i[1460] & sel_one_hot_i[11];
  assign data_masked[1459] = data_i[1459] & sel_one_hot_i[11];
  assign data_masked[1458] = data_i[1458] & sel_one_hot_i[11];
  assign data_masked[1457] = data_i[1457] & sel_one_hot_i[11];
  assign data_masked[1456] = data_i[1456] & sel_one_hot_i[11];
  assign data_masked[1455] = data_i[1455] & sel_one_hot_i[11];
  assign data_masked[1454] = data_i[1454] & sel_one_hot_i[11];
  assign data_masked[1453] = data_i[1453] & sel_one_hot_i[11];
  assign data_masked[1452] = data_i[1452] & sel_one_hot_i[11];
  assign data_masked[1451] = data_i[1451] & sel_one_hot_i[11];
  assign data_masked[1450] = data_i[1450] & sel_one_hot_i[11];
  assign data_masked[1449] = data_i[1449] & sel_one_hot_i[11];
  assign data_masked[1448] = data_i[1448] & sel_one_hot_i[11];
  assign data_masked[1447] = data_i[1447] & sel_one_hot_i[11];
  assign data_masked[1446] = data_i[1446] & sel_one_hot_i[11];
  assign data_masked[1445] = data_i[1445] & sel_one_hot_i[11];
  assign data_masked[1444] = data_i[1444] & sel_one_hot_i[11];
  assign data_masked[1443] = data_i[1443] & sel_one_hot_i[11];
  assign data_masked[1442] = data_i[1442] & sel_one_hot_i[11];
  assign data_masked[1441] = data_i[1441] & sel_one_hot_i[11];
  assign data_masked[1440] = data_i[1440] & sel_one_hot_i[11];
  assign data_masked[1439] = data_i[1439] & sel_one_hot_i[11];
  assign data_masked[1438] = data_i[1438] & sel_one_hot_i[11];
  assign data_masked[1437] = data_i[1437] & sel_one_hot_i[11];
  assign data_masked[1436] = data_i[1436] & sel_one_hot_i[11];
  assign data_masked[1435] = data_i[1435] & sel_one_hot_i[11];
  assign data_masked[1434] = data_i[1434] & sel_one_hot_i[11];
  assign data_masked[1433] = data_i[1433] & sel_one_hot_i[11];
  assign data_masked[1432] = data_i[1432] & sel_one_hot_i[11];
  assign data_masked[1431] = data_i[1431] & sel_one_hot_i[11];
  assign data_masked[1430] = data_i[1430] & sel_one_hot_i[11];
  assign data_masked[1429] = data_i[1429] & sel_one_hot_i[11];
  assign data_masked[1428] = data_i[1428] & sel_one_hot_i[11];
  assign data_masked[1427] = data_i[1427] & sel_one_hot_i[11];
  assign data_masked[1426] = data_i[1426] & sel_one_hot_i[11];
  assign data_masked[1425] = data_i[1425] & sel_one_hot_i[11];
  assign data_masked[1424] = data_i[1424] & sel_one_hot_i[11];
  assign data_masked[1423] = data_i[1423] & sel_one_hot_i[11];
  assign data_masked[1422] = data_i[1422] & sel_one_hot_i[11];
  assign data_masked[1421] = data_i[1421] & sel_one_hot_i[11];
  assign data_masked[1420] = data_i[1420] & sel_one_hot_i[11];
  assign data_masked[1419] = data_i[1419] & sel_one_hot_i[11];
  assign data_masked[1418] = data_i[1418] & sel_one_hot_i[11];
  assign data_masked[1417] = data_i[1417] & sel_one_hot_i[11];
  assign data_masked[1416] = data_i[1416] & sel_one_hot_i[11];
  assign data_masked[1415] = data_i[1415] & sel_one_hot_i[11];
  assign data_masked[1414] = data_i[1414] & sel_one_hot_i[11];
  assign data_masked[1413] = data_i[1413] & sel_one_hot_i[11];
  assign data_masked[1412] = data_i[1412] & sel_one_hot_i[11];
  assign data_masked[1411] = data_i[1411] & sel_one_hot_i[11];
  assign data_masked[1410] = data_i[1410] & sel_one_hot_i[11];
  assign data_masked[1409] = data_i[1409] & sel_one_hot_i[11];
  assign data_masked[1408] = data_i[1408] & sel_one_hot_i[11];
  assign data_masked[1663] = data_i[1663] & sel_one_hot_i[12];
  assign data_masked[1662] = data_i[1662] & sel_one_hot_i[12];
  assign data_masked[1661] = data_i[1661] & sel_one_hot_i[12];
  assign data_masked[1660] = data_i[1660] & sel_one_hot_i[12];
  assign data_masked[1659] = data_i[1659] & sel_one_hot_i[12];
  assign data_masked[1658] = data_i[1658] & sel_one_hot_i[12];
  assign data_masked[1657] = data_i[1657] & sel_one_hot_i[12];
  assign data_masked[1656] = data_i[1656] & sel_one_hot_i[12];
  assign data_masked[1655] = data_i[1655] & sel_one_hot_i[12];
  assign data_masked[1654] = data_i[1654] & sel_one_hot_i[12];
  assign data_masked[1653] = data_i[1653] & sel_one_hot_i[12];
  assign data_masked[1652] = data_i[1652] & sel_one_hot_i[12];
  assign data_masked[1651] = data_i[1651] & sel_one_hot_i[12];
  assign data_masked[1650] = data_i[1650] & sel_one_hot_i[12];
  assign data_masked[1649] = data_i[1649] & sel_one_hot_i[12];
  assign data_masked[1648] = data_i[1648] & sel_one_hot_i[12];
  assign data_masked[1647] = data_i[1647] & sel_one_hot_i[12];
  assign data_masked[1646] = data_i[1646] & sel_one_hot_i[12];
  assign data_masked[1645] = data_i[1645] & sel_one_hot_i[12];
  assign data_masked[1644] = data_i[1644] & sel_one_hot_i[12];
  assign data_masked[1643] = data_i[1643] & sel_one_hot_i[12];
  assign data_masked[1642] = data_i[1642] & sel_one_hot_i[12];
  assign data_masked[1641] = data_i[1641] & sel_one_hot_i[12];
  assign data_masked[1640] = data_i[1640] & sel_one_hot_i[12];
  assign data_masked[1639] = data_i[1639] & sel_one_hot_i[12];
  assign data_masked[1638] = data_i[1638] & sel_one_hot_i[12];
  assign data_masked[1637] = data_i[1637] & sel_one_hot_i[12];
  assign data_masked[1636] = data_i[1636] & sel_one_hot_i[12];
  assign data_masked[1635] = data_i[1635] & sel_one_hot_i[12];
  assign data_masked[1634] = data_i[1634] & sel_one_hot_i[12];
  assign data_masked[1633] = data_i[1633] & sel_one_hot_i[12];
  assign data_masked[1632] = data_i[1632] & sel_one_hot_i[12];
  assign data_masked[1631] = data_i[1631] & sel_one_hot_i[12];
  assign data_masked[1630] = data_i[1630] & sel_one_hot_i[12];
  assign data_masked[1629] = data_i[1629] & sel_one_hot_i[12];
  assign data_masked[1628] = data_i[1628] & sel_one_hot_i[12];
  assign data_masked[1627] = data_i[1627] & sel_one_hot_i[12];
  assign data_masked[1626] = data_i[1626] & sel_one_hot_i[12];
  assign data_masked[1625] = data_i[1625] & sel_one_hot_i[12];
  assign data_masked[1624] = data_i[1624] & sel_one_hot_i[12];
  assign data_masked[1623] = data_i[1623] & sel_one_hot_i[12];
  assign data_masked[1622] = data_i[1622] & sel_one_hot_i[12];
  assign data_masked[1621] = data_i[1621] & sel_one_hot_i[12];
  assign data_masked[1620] = data_i[1620] & sel_one_hot_i[12];
  assign data_masked[1619] = data_i[1619] & sel_one_hot_i[12];
  assign data_masked[1618] = data_i[1618] & sel_one_hot_i[12];
  assign data_masked[1617] = data_i[1617] & sel_one_hot_i[12];
  assign data_masked[1616] = data_i[1616] & sel_one_hot_i[12];
  assign data_masked[1615] = data_i[1615] & sel_one_hot_i[12];
  assign data_masked[1614] = data_i[1614] & sel_one_hot_i[12];
  assign data_masked[1613] = data_i[1613] & sel_one_hot_i[12];
  assign data_masked[1612] = data_i[1612] & sel_one_hot_i[12];
  assign data_masked[1611] = data_i[1611] & sel_one_hot_i[12];
  assign data_masked[1610] = data_i[1610] & sel_one_hot_i[12];
  assign data_masked[1609] = data_i[1609] & sel_one_hot_i[12];
  assign data_masked[1608] = data_i[1608] & sel_one_hot_i[12];
  assign data_masked[1607] = data_i[1607] & sel_one_hot_i[12];
  assign data_masked[1606] = data_i[1606] & sel_one_hot_i[12];
  assign data_masked[1605] = data_i[1605] & sel_one_hot_i[12];
  assign data_masked[1604] = data_i[1604] & sel_one_hot_i[12];
  assign data_masked[1603] = data_i[1603] & sel_one_hot_i[12];
  assign data_masked[1602] = data_i[1602] & sel_one_hot_i[12];
  assign data_masked[1601] = data_i[1601] & sel_one_hot_i[12];
  assign data_masked[1600] = data_i[1600] & sel_one_hot_i[12];
  assign data_masked[1599] = data_i[1599] & sel_one_hot_i[12];
  assign data_masked[1598] = data_i[1598] & sel_one_hot_i[12];
  assign data_masked[1597] = data_i[1597] & sel_one_hot_i[12];
  assign data_masked[1596] = data_i[1596] & sel_one_hot_i[12];
  assign data_masked[1595] = data_i[1595] & sel_one_hot_i[12];
  assign data_masked[1594] = data_i[1594] & sel_one_hot_i[12];
  assign data_masked[1593] = data_i[1593] & sel_one_hot_i[12];
  assign data_masked[1592] = data_i[1592] & sel_one_hot_i[12];
  assign data_masked[1591] = data_i[1591] & sel_one_hot_i[12];
  assign data_masked[1590] = data_i[1590] & sel_one_hot_i[12];
  assign data_masked[1589] = data_i[1589] & sel_one_hot_i[12];
  assign data_masked[1588] = data_i[1588] & sel_one_hot_i[12];
  assign data_masked[1587] = data_i[1587] & sel_one_hot_i[12];
  assign data_masked[1586] = data_i[1586] & sel_one_hot_i[12];
  assign data_masked[1585] = data_i[1585] & sel_one_hot_i[12];
  assign data_masked[1584] = data_i[1584] & sel_one_hot_i[12];
  assign data_masked[1583] = data_i[1583] & sel_one_hot_i[12];
  assign data_masked[1582] = data_i[1582] & sel_one_hot_i[12];
  assign data_masked[1581] = data_i[1581] & sel_one_hot_i[12];
  assign data_masked[1580] = data_i[1580] & sel_one_hot_i[12];
  assign data_masked[1579] = data_i[1579] & sel_one_hot_i[12];
  assign data_masked[1578] = data_i[1578] & sel_one_hot_i[12];
  assign data_masked[1577] = data_i[1577] & sel_one_hot_i[12];
  assign data_masked[1576] = data_i[1576] & sel_one_hot_i[12];
  assign data_masked[1575] = data_i[1575] & sel_one_hot_i[12];
  assign data_masked[1574] = data_i[1574] & sel_one_hot_i[12];
  assign data_masked[1573] = data_i[1573] & sel_one_hot_i[12];
  assign data_masked[1572] = data_i[1572] & sel_one_hot_i[12];
  assign data_masked[1571] = data_i[1571] & sel_one_hot_i[12];
  assign data_masked[1570] = data_i[1570] & sel_one_hot_i[12];
  assign data_masked[1569] = data_i[1569] & sel_one_hot_i[12];
  assign data_masked[1568] = data_i[1568] & sel_one_hot_i[12];
  assign data_masked[1567] = data_i[1567] & sel_one_hot_i[12];
  assign data_masked[1566] = data_i[1566] & sel_one_hot_i[12];
  assign data_masked[1565] = data_i[1565] & sel_one_hot_i[12];
  assign data_masked[1564] = data_i[1564] & sel_one_hot_i[12];
  assign data_masked[1563] = data_i[1563] & sel_one_hot_i[12];
  assign data_masked[1562] = data_i[1562] & sel_one_hot_i[12];
  assign data_masked[1561] = data_i[1561] & sel_one_hot_i[12];
  assign data_masked[1560] = data_i[1560] & sel_one_hot_i[12];
  assign data_masked[1559] = data_i[1559] & sel_one_hot_i[12];
  assign data_masked[1558] = data_i[1558] & sel_one_hot_i[12];
  assign data_masked[1557] = data_i[1557] & sel_one_hot_i[12];
  assign data_masked[1556] = data_i[1556] & sel_one_hot_i[12];
  assign data_masked[1555] = data_i[1555] & sel_one_hot_i[12];
  assign data_masked[1554] = data_i[1554] & sel_one_hot_i[12];
  assign data_masked[1553] = data_i[1553] & sel_one_hot_i[12];
  assign data_masked[1552] = data_i[1552] & sel_one_hot_i[12];
  assign data_masked[1551] = data_i[1551] & sel_one_hot_i[12];
  assign data_masked[1550] = data_i[1550] & sel_one_hot_i[12];
  assign data_masked[1549] = data_i[1549] & sel_one_hot_i[12];
  assign data_masked[1548] = data_i[1548] & sel_one_hot_i[12];
  assign data_masked[1547] = data_i[1547] & sel_one_hot_i[12];
  assign data_masked[1546] = data_i[1546] & sel_one_hot_i[12];
  assign data_masked[1545] = data_i[1545] & sel_one_hot_i[12];
  assign data_masked[1544] = data_i[1544] & sel_one_hot_i[12];
  assign data_masked[1543] = data_i[1543] & sel_one_hot_i[12];
  assign data_masked[1542] = data_i[1542] & sel_one_hot_i[12];
  assign data_masked[1541] = data_i[1541] & sel_one_hot_i[12];
  assign data_masked[1540] = data_i[1540] & sel_one_hot_i[12];
  assign data_masked[1539] = data_i[1539] & sel_one_hot_i[12];
  assign data_masked[1538] = data_i[1538] & sel_one_hot_i[12];
  assign data_masked[1537] = data_i[1537] & sel_one_hot_i[12];
  assign data_masked[1536] = data_i[1536] & sel_one_hot_i[12];
  assign data_masked[1791] = data_i[1791] & sel_one_hot_i[13];
  assign data_masked[1790] = data_i[1790] & sel_one_hot_i[13];
  assign data_masked[1789] = data_i[1789] & sel_one_hot_i[13];
  assign data_masked[1788] = data_i[1788] & sel_one_hot_i[13];
  assign data_masked[1787] = data_i[1787] & sel_one_hot_i[13];
  assign data_masked[1786] = data_i[1786] & sel_one_hot_i[13];
  assign data_masked[1785] = data_i[1785] & sel_one_hot_i[13];
  assign data_masked[1784] = data_i[1784] & sel_one_hot_i[13];
  assign data_masked[1783] = data_i[1783] & sel_one_hot_i[13];
  assign data_masked[1782] = data_i[1782] & sel_one_hot_i[13];
  assign data_masked[1781] = data_i[1781] & sel_one_hot_i[13];
  assign data_masked[1780] = data_i[1780] & sel_one_hot_i[13];
  assign data_masked[1779] = data_i[1779] & sel_one_hot_i[13];
  assign data_masked[1778] = data_i[1778] & sel_one_hot_i[13];
  assign data_masked[1777] = data_i[1777] & sel_one_hot_i[13];
  assign data_masked[1776] = data_i[1776] & sel_one_hot_i[13];
  assign data_masked[1775] = data_i[1775] & sel_one_hot_i[13];
  assign data_masked[1774] = data_i[1774] & sel_one_hot_i[13];
  assign data_masked[1773] = data_i[1773] & sel_one_hot_i[13];
  assign data_masked[1772] = data_i[1772] & sel_one_hot_i[13];
  assign data_masked[1771] = data_i[1771] & sel_one_hot_i[13];
  assign data_masked[1770] = data_i[1770] & sel_one_hot_i[13];
  assign data_masked[1769] = data_i[1769] & sel_one_hot_i[13];
  assign data_masked[1768] = data_i[1768] & sel_one_hot_i[13];
  assign data_masked[1767] = data_i[1767] & sel_one_hot_i[13];
  assign data_masked[1766] = data_i[1766] & sel_one_hot_i[13];
  assign data_masked[1765] = data_i[1765] & sel_one_hot_i[13];
  assign data_masked[1764] = data_i[1764] & sel_one_hot_i[13];
  assign data_masked[1763] = data_i[1763] & sel_one_hot_i[13];
  assign data_masked[1762] = data_i[1762] & sel_one_hot_i[13];
  assign data_masked[1761] = data_i[1761] & sel_one_hot_i[13];
  assign data_masked[1760] = data_i[1760] & sel_one_hot_i[13];
  assign data_masked[1759] = data_i[1759] & sel_one_hot_i[13];
  assign data_masked[1758] = data_i[1758] & sel_one_hot_i[13];
  assign data_masked[1757] = data_i[1757] & sel_one_hot_i[13];
  assign data_masked[1756] = data_i[1756] & sel_one_hot_i[13];
  assign data_masked[1755] = data_i[1755] & sel_one_hot_i[13];
  assign data_masked[1754] = data_i[1754] & sel_one_hot_i[13];
  assign data_masked[1753] = data_i[1753] & sel_one_hot_i[13];
  assign data_masked[1752] = data_i[1752] & sel_one_hot_i[13];
  assign data_masked[1751] = data_i[1751] & sel_one_hot_i[13];
  assign data_masked[1750] = data_i[1750] & sel_one_hot_i[13];
  assign data_masked[1749] = data_i[1749] & sel_one_hot_i[13];
  assign data_masked[1748] = data_i[1748] & sel_one_hot_i[13];
  assign data_masked[1747] = data_i[1747] & sel_one_hot_i[13];
  assign data_masked[1746] = data_i[1746] & sel_one_hot_i[13];
  assign data_masked[1745] = data_i[1745] & sel_one_hot_i[13];
  assign data_masked[1744] = data_i[1744] & sel_one_hot_i[13];
  assign data_masked[1743] = data_i[1743] & sel_one_hot_i[13];
  assign data_masked[1742] = data_i[1742] & sel_one_hot_i[13];
  assign data_masked[1741] = data_i[1741] & sel_one_hot_i[13];
  assign data_masked[1740] = data_i[1740] & sel_one_hot_i[13];
  assign data_masked[1739] = data_i[1739] & sel_one_hot_i[13];
  assign data_masked[1738] = data_i[1738] & sel_one_hot_i[13];
  assign data_masked[1737] = data_i[1737] & sel_one_hot_i[13];
  assign data_masked[1736] = data_i[1736] & sel_one_hot_i[13];
  assign data_masked[1735] = data_i[1735] & sel_one_hot_i[13];
  assign data_masked[1734] = data_i[1734] & sel_one_hot_i[13];
  assign data_masked[1733] = data_i[1733] & sel_one_hot_i[13];
  assign data_masked[1732] = data_i[1732] & sel_one_hot_i[13];
  assign data_masked[1731] = data_i[1731] & sel_one_hot_i[13];
  assign data_masked[1730] = data_i[1730] & sel_one_hot_i[13];
  assign data_masked[1729] = data_i[1729] & sel_one_hot_i[13];
  assign data_masked[1728] = data_i[1728] & sel_one_hot_i[13];
  assign data_masked[1727] = data_i[1727] & sel_one_hot_i[13];
  assign data_masked[1726] = data_i[1726] & sel_one_hot_i[13];
  assign data_masked[1725] = data_i[1725] & sel_one_hot_i[13];
  assign data_masked[1724] = data_i[1724] & sel_one_hot_i[13];
  assign data_masked[1723] = data_i[1723] & sel_one_hot_i[13];
  assign data_masked[1722] = data_i[1722] & sel_one_hot_i[13];
  assign data_masked[1721] = data_i[1721] & sel_one_hot_i[13];
  assign data_masked[1720] = data_i[1720] & sel_one_hot_i[13];
  assign data_masked[1719] = data_i[1719] & sel_one_hot_i[13];
  assign data_masked[1718] = data_i[1718] & sel_one_hot_i[13];
  assign data_masked[1717] = data_i[1717] & sel_one_hot_i[13];
  assign data_masked[1716] = data_i[1716] & sel_one_hot_i[13];
  assign data_masked[1715] = data_i[1715] & sel_one_hot_i[13];
  assign data_masked[1714] = data_i[1714] & sel_one_hot_i[13];
  assign data_masked[1713] = data_i[1713] & sel_one_hot_i[13];
  assign data_masked[1712] = data_i[1712] & sel_one_hot_i[13];
  assign data_masked[1711] = data_i[1711] & sel_one_hot_i[13];
  assign data_masked[1710] = data_i[1710] & sel_one_hot_i[13];
  assign data_masked[1709] = data_i[1709] & sel_one_hot_i[13];
  assign data_masked[1708] = data_i[1708] & sel_one_hot_i[13];
  assign data_masked[1707] = data_i[1707] & sel_one_hot_i[13];
  assign data_masked[1706] = data_i[1706] & sel_one_hot_i[13];
  assign data_masked[1705] = data_i[1705] & sel_one_hot_i[13];
  assign data_masked[1704] = data_i[1704] & sel_one_hot_i[13];
  assign data_masked[1703] = data_i[1703] & sel_one_hot_i[13];
  assign data_masked[1702] = data_i[1702] & sel_one_hot_i[13];
  assign data_masked[1701] = data_i[1701] & sel_one_hot_i[13];
  assign data_masked[1700] = data_i[1700] & sel_one_hot_i[13];
  assign data_masked[1699] = data_i[1699] & sel_one_hot_i[13];
  assign data_masked[1698] = data_i[1698] & sel_one_hot_i[13];
  assign data_masked[1697] = data_i[1697] & sel_one_hot_i[13];
  assign data_masked[1696] = data_i[1696] & sel_one_hot_i[13];
  assign data_masked[1695] = data_i[1695] & sel_one_hot_i[13];
  assign data_masked[1694] = data_i[1694] & sel_one_hot_i[13];
  assign data_masked[1693] = data_i[1693] & sel_one_hot_i[13];
  assign data_masked[1692] = data_i[1692] & sel_one_hot_i[13];
  assign data_masked[1691] = data_i[1691] & sel_one_hot_i[13];
  assign data_masked[1690] = data_i[1690] & sel_one_hot_i[13];
  assign data_masked[1689] = data_i[1689] & sel_one_hot_i[13];
  assign data_masked[1688] = data_i[1688] & sel_one_hot_i[13];
  assign data_masked[1687] = data_i[1687] & sel_one_hot_i[13];
  assign data_masked[1686] = data_i[1686] & sel_one_hot_i[13];
  assign data_masked[1685] = data_i[1685] & sel_one_hot_i[13];
  assign data_masked[1684] = data_i[1684] & sel_one_hot_i[13];
  assign data_masked[1683] = data_i[1683] & sel_one_hot_i[13];
  assign data_masked[1682] = data_i[1682] & sel_one_hot_i[13];
  assign data_masked[1681] = data_i[1681] & sel_one_hot_i[13];
  assign data_masked[1680] = data_i[1680] & sel_one_hot_i[13];
  assign data_masked[1679] = data_i[1679] & sel_one_hot_i[13];
  assign data_masked[1678] = data_i[1678] & sel_one_hot_i[13];
  assign data_masked[1677] = data_i[1677] & sel_one_hot_i[13];
  assign data_masked[1676] = data_i[1676] & sel_one_hot_i[13];
  assign data_masked[1675] = data_i[1675] & sel_one_hot_i[13];
  assign data_masked[1674] = data_i[1674] & sel_one_hot_i[13];
  assign data_masked[1673] = data_i[1673] & sel_one_hot_i[13];
  assign data_masked[1672] = data_i[1672] & sel_one_hot_i[13];
  assign data_masked[1671] = data_i[1671] & sel_one_hot_i[13];
  assign data_masked[1670] = data_i[1670] & sel_one_hot_i[13];
  assign data_masked[1669] = data_i[1669] & sel_one_hot_i[13];
  assign data_masked[1668] = data_i[1668] & sel_one_hot_i[13];
  assign data_masked[1667] = data_i[1667] & sel_one_hot_i[13];
  assign data_masked[1666] = data_i[1666] & sel_one_hot_i[13];
  assign data_masked[1665] = data_i[1665] & sel_one_hot_i[13];
  assign data_masked[1664] = data_i[1664] & sel_one_hot_i[13];
  assign data_masked[1919] = data_i[1919] & sel_one_hot_i[14];
  assign data_masked[1918] = data_i[1918] & sel_one_hot_i[14];
  assign data_masked[1917] = data_i[1917] & sel_one_hot_i[14];
  assign data_masked[1916] = data_i[1916] & sel_one_hot_i[14];
  assign data_masked[1915] = data_i[1915] & sel_one_hot_i[14];
  assign data_masked[1914] = data_i[1914] & sel_one_hot_i[14];
  assign data_masked[1913] = data_i[1913] & sel_one_hot_i[14];
  assign data_masked[1912] = data_i[1912] & sel_one_hot_i[14];
  assign data_masked[1911] = data_i[1911] & sel_one_hot_i[14];
  assign data_masked[1910] = data_i[1910] & sel_one_hot_i[14];
  assign data_masked[1909] = data_i[1909] & sel_one_hot_i[14];
  assign data_masked[1908] = data_i[1908] & sel_one_hot_i[14];
  assign data_masked[1907] = data_i[1907] & sel_one_hot_i[14];
  assign data_masked[1906] = data_i[1906] & sel_one_hot_i[14];
  assign data_masked[1905] = data_i[1905] & sel_one_hot_i[14];
  assign data_masked[1904] = data_i[1904] & sel_one_hot_i[14];
  assign data_masked[1903] = data_i[1903] & sel_one_hot_i[14];
  assign data_masked[1902] = data_i[1902] & sel_one_hot_i[14];
  assign data_masked[1901] = data_i[1901] & sel_one_hot_i[14];
  assign data_masked[1900] = data_i[1900] & sel_one_hot_i[14];
  assign data_masked[1899] = data_i[1899] & sel_one_hot_i[14];
  assign data_masked[1898] = data_i[1898] & sel_one_hot_i[14];
  assign data_masked[1897] = data_i[1897] & sel_one_hot_i[14];
  assign data_masked[1896] = data_i[1896] & sel_one_hot_i[14];
  assign data_masked[1895] = data_i[1895] & sel_one_hot_i[14];
  assign data_masked[1894] = data_i[1894] & sel_one_hot_i[14];
  assign data_masked[1893] = data_i[1893] & sel_one_hot_i[14];
  assign data_masked[1892] = data_i[1892] & sel_one_hot_i[14];
  assign data_masked[1891] = data_i[1891] & sel_one_hot_i[14];
  assign data_masked[1890] = data_i[1890] & sel_one_hot_i[14];
  assign data_masked[1889] = data_i[1889] & sel_one_hot_i[14];
  assign data_masked[1888] = data_i[1888] & sel_one_hot_i[14];
  assign data_masked[1887] = data_i[1887] & sel_one_hot_i[14];
  assign data_masked[1886] = data_i[1886] & sel_one_hot_i[14];
  assign data_masked[1885] = data_i[1885] & sel_one_hot_i[14];
  assign data_masked[1884] = data_i[1884] & sel_one_hot_i[14];
  assign data_masked[1883] = data_i[1883] & sel_one_hot_i[14];
  assign data_masked[1882] = data_i[1882] & sel_one_hot_i[14];
  assign data_masked[1881] = data_i[1881] & sel_one_hot_i[14];
  assign data_masked[1880] = data_i[1880] & sel_one_hot_i[14];
  assign data_masked[1879] = data_i[1879] & sel_one_hot_i[14];
  assign data_masked[1878] = data_i[1878] & sel_one_hot_i[14];
  assign data_masked[1877] = data_i[1877] & sel_one_hot_i[14];
  assign data_masked[1876] = data_i[1876] & sel_one_hot_i[14];
  assign data_masked[1875] = data_i[1875] & sel_one_hot_i[14];
  assign data_masked[1874] = data_i[1874] & sel_one_hot_i[14];
  assign data_masked[1873] = data_i[1873] & sel_one_hot_i[14];
  assign data_masked[1872] = data_i[1872] & sel_one_hot_i[14];
  assign data_masked[1871] = data_i[1871] & sel_one_hot_i[14];
  assign data_masked[1870] = data_i[1870] & sel_one_hot_i[14];
  assign data_masked[1869] = data_i[1869] & sel_one_hot_i[14];
  assign data_masked[1868] = data_i[1868] & sel_one_hot_i[14];
  assign data_masked[1867] = data_i[1867] & sel_one_hot_i[14];
  assign data_masked[1866] = data_i[1866] & sel_one_hot_i[14];
  assign data_masked[1865] = data_i[1865] & sel_one_hot_i[14];
  assign data_masked[1864] = data_i[1864] & sel_one_hot_i[14];
  assign data_masked[1863] = data_i[1863] & sel_one_hot_i[14];
  assign data_masked[1862] = data_i[1862] & sel_one_hot_i[14];
  assign data_masked[1861] = data_i[1861] & sel_one_hot_i[14];
  assign data_masked[1860] = data_i[1860] & sel_one_hot_i[14];
  assign data_masked[1859] = data_i[1859] & sel_one_hot_i[14];
  assign data_masked[1858] = data_i[1858] & sel_one_hot_i[14];
  assign data_masked[1857] = data_i[1857] & sel_one_hot_i[14];
  assign data_masked[1856] = data_i[1856] & sel_one_hot_i[14];
  assign data_masked[1855] = data_i[1855] & sel_one_hot_i[14];
  assign data_masked[1854] = data_i[1854] & sel_one_hot_i[14];
  assign data_masked[1853] = data_i[1853] & sel_one_hot_i[14];
  assign data_masked[1852] = data_i[1852] & sel_one_hot_i[14];
  assign data_masked[1851] = data_i[1851] & sel_one_hot_i[14];
  assign data_masked[1850] = data_i[1850] & sel_one_hot_i[14];
  assign data_masked[1849] = data_i[1849] & sel_one_hot_i[14];
  assign data_masked[1848] = data_i[1848] & sel_one_hot_i[14];
  assign data_masked[1847] = data_i[1847] & sel_one_hot_i[14];
  assign data_masked[1846] = data_i[1846] & sel_one_hot_i[14];
  assign data_masked[1845] = data_i[1845] & sel_one_hot_i[14];
  assign data_masked[1844] = data_i[1844] & sel_one_hot_i[14];
  assign data_masked[1843] = data_i[1843] & sel_one_hot_i[14];
  assign data_masked[1842] = data_i[1842] & sel_one_hot_i[14];
  assign data_masked[1841] = data_i[1841] & sel_one_hot_i[14];
  assign data_masked[1840] = data_i[1840] & sel_one_hot_i[14];
  assign data_masked[1839] = data_i[1839] & sel_one_hot_i[14];
  assign data_masked[1838] = data_i[1838] & sel_one_hot_i[14];
  assign data_masked[1837] = data_i[1837] & sel_one_hot_i[14];
  assign data_masked[1836] = data_i[1836] & sel_one_hot_i[14];
  assign data_masked[1835] = data_i[1835] & sel_one_hot_i[14];
  assign data_masked[1834] = data_i[1834] & sel_one_hot_i[14];
  assign data_masked[1833] = data_i[1833] & sel_one_hot_i[14];
  assign data_masked[1832] = data_i[1832] & sel_one_hot_i[14];
  assign data_masked[1831] = data_i[1831] & sel_one_hot_i[14];
  assign data_masked[1830] = data_i[1830] & sel_one_hot_i[14];
  assign data_masked[1829] = data_i[1829] & sel_one_hot_i[14];
  assign data_masked[1828] = data_i[1828] & sel_one_hot_i[14];
  assign data_masked[1827] = data_i[1827] & sel_one_hot_i[14];
  assign data_masked[1826] = data_i[1826] & sel_one_hot_i[14];
  assign data_masked[1825] = data_i[1825] & sel_one_hot_i[14];
  assign data_masked[1824] = data_i[1824] & sel_one_hot_i[14];
  assign data_masked[1823] = data_i[1823] & sel_one_hot_i[14];
  assign data_masked[1822] = data_i[1822] & sel_one_hot_i[14];
  assign data_masked[1821] = data_i[1821] & sel_one_hot_i[14];
  assign data_masked[1820] = data_i[1820] & sel_one_hot_i[14];
  assign data_masked[1819] = data_i[1819] & sel_one_hot_i[14];
  assign data_masked[1818] = data_i[1818] & sel_one_hot_i[14];
  assign data_masked[1817] = data_i[1817] & sel_one_hot_i[14];
  assign data_masked[1816] = data_i[1816] & sel_one_hot_i[14];
  assign data_masked[1815] = data_i[1815] & sel_one_hot_i[14];
  assign data_masked[1814] = data_i[1814] & sel_one_hot_i[14];
  assign data_masked[1813] = data_i[1813] & sel_one_hot_i[14];
  assign data_masked[1812] = data_i[1812] & sel_one_hot_i[14];
  assign data_masked[1811] = data_i[1811] & sel_one_hot_i[14];
  assign data_masked[1810] = data_i[1810] & sel_one_hot_i[14];
  assign data_masked[1809] = data_i[1809] & sel_one_hot_i[14];
  assign data_masked[1808] = data_i[1808] & sel_one_hot_i[14];
  assign data_masked[1807] = data_i[1807] & sel_one_hot_i[14];
  assign data_masked[1806] = data_i[1806] & sel_one_hot_i[14];
  assign data_masked[1805] = data_i[1805] & sel_one_hot_i[14];
  assign data_masked[1804] = data_i[1804] & sel_one_hot_i[14];
  assign data_masked[1803] = data_i[1803] & sel_one_hot_i[14];
  assign data_masked[1802] = data_i[1802] & sel_one_hot_i[14];
  assign data_masked[1801] = data_i[1801] & sel_one_hot_i[14];
  assign data_masked[1800] = data_i[1800] & sel_one_hot_i[14];
  assign data_masked[1799] = data_i[1799] & sel_one_hot_i[14];
  assign data_masked[1798] = data_i[1798] & sel_one_hot_i[14];
  assign data_masked[1797] = data_i[1797] & sel_one_hot_i[14];
  assign data_masked[1796] = data_i[1796] & sel_one_hot_i[14];
  assign data_masked[1795] = data_i[1795] & sel_one_hot_i[14];
  assign data_masked[1794] = data_i[1794] & sel_one_hot_i[14];
  assign data_masked[1793] = data_i[1793] & sel_one_hot_i[14];
  assign data_masked[1792] = data_i[1792] & sel_one_hot_i[14];
  assign data_masked[2047] = data_i[2047] & sel_one_hot_i[15];
  assign data_masked[2046] = data_i[2046] & sel_one_hot_i[15];
  assign data_masked[2045] = data_i[2045] & sel_one_hot_i[15];
  assign data_masked[2044] = data_i[2044] & sel_one_hot_i[15];
  assign data_masked[2043] = data_i[2043] & sel_one_hot_i[15];
  assign data_masked[2042] = data_i[2042] & sel_one_hot_i[15];
  assign data_masked[2041] = data_i[2041] & sel_one_hot_i[15];
  assign data_masked[2040] = data_i[2040] & sel_one_hot_i[15];
  assign data_masked[2039] = data_i[2039] & sel_one_hot_i[15];
  assign data_masked[2038] = data_i[2038] & sel_one_hot_i[15];
  assign data_masked[2037] = data_i[2037] & sel_one_hot_i[15];
  assign data_masked[2036] = data_i[2036] & sel_one_hot_i[15];
  assign data_masked[2035] = data_i[2035] & sel_one_hot_i[15];
  assign data_masked[2034] = data_i[2034] & sel_one_hot_i[15];
  assign data_masked[2033] = data_i[2033] & sel_one_hot_i[15];
  assign data_masked[2032] = data_i[2032] & sel_one_hot_i[15];
  assign data_masked[2031] = data_i[2031] & sel_one_hot_i[15];
  assign data_masked[2030] = data_i[2030] & sel_one_hot_i[15];
  assign data_masked[2029] = data_i[2029] & sel_one_hot_i[15];
  assign data_masked[2028] = data_i[2028] & sel_one_hot_i[15];
  assign data_masked[2027] = data_i[2027] & sel_one_hot_i[15];
  assign data_masked[2026] = data_i[2026] & sel_one_hot_i[15];
  assign data_masked[2025] = data_i[2025] & sel_one_hot_i[15];
  assign data_masked[2024] = data_i[2024] & sel_one_hot_i[15];
  assign data_masked[2023] = data_i[2023] & sel_one_hot_i[15];
  assign data_masked[2022] = data_i[2022] & sel_one_hot_i[15];
  assign data_masked[2021] = data_i[2021] & sel_one_hot_i[15];
  assign data_masked[2020] = data_i[2020] & sel_one_hot_i[15];
  assign data_masked[2019] = data_i[2019] & sel_one_hot_i[15];
  assign data_masked[2018] = data_i[2018] & sel_one_hot_i[15];
  assign data_masked[2017] = data_i[2017] & sel_one_hot_i[15];
  assign data_masked[2016] = data_i[2016] & sel_one_hot_i[15];
  assign data_masked[2015] = data_i[2015] & sel_one_hot_i[15];
  assign data_masked[2014] = data_i[2014] & sel_one_hot_i[15];
  assign data_masked[2013] = data_i[2013] & sel_one_hot_i[15];
  assign data_masked[2012] = data_i[2012] & sel_one_hot_i[15];
  assign data_masked[2011] = data_i[2011] & sel_one_hot_i[15];
  assign data_masked[2010] = data_i[2010] & sel_one_hot_i[15];
  assign data_masked[2009] = data_i[2009] & sel_one_hot_i[15];
  assign data_masked[2008] = data_i[2008] & sel_one_hot_i[15];
  assign data_masked[2007] = data_i[2007] & sel_one_hot_i[15];
  assign data_masked[2006] = data_i[2006] & sel_one_hot_i[15];
  assign data_masked[2005] = data_i[2005] & sel_one_hot_i[15];
  assign data_masked[2004] = data_i[2004] & sel_one_hot_i[15];
  assign data_masked[2003] = data_i[2003] & sel_one_hot_i[15];
  assign data_masked[2002] = data_i[2002] & sel_one_hot_i[15];
  assign data_masked[2001] = data_i[2001] & sel_one_hot_i[15];
  assign data_masked[2000] = data_i[2000] & sel_one_hot_i[15];
  assign data_masked[1999] = data_i[1999] & sel_one_hot_i[15];
  assign data_masked[1998] = data_i[1998] & sel_one_hot_i[15];
  assign data_masked[1997] = data_i[1997] & sel_one_hot_i[15];
  assign data_masked[1996] = data_i[1996] & sel_one_hot_i[15];
  assign data_masked[1995] = data_i[1995] & sel_one_hot_i[15];
  assign data_masked[1994] = data_i[1994] & sel_one_hot_i[15];
  assign data_masked[1993] = data_i[1993] & sel_one_hot_i[15];
  assign data_masked[1992] = data_i[1992] & sel_one_hot_i[15];
  assign data_masked[1991] = data_i[1991] & sel_one_hot_i[15];
  assign data_masked[1990] = data_i[1990] & sel_one_hot_i[15];
  assign data_masked[1989] = data_i[1989] & sel_one_hot_i[15];
  assign data_masked[1988] = data_i[1988] & sel_one_hot_i[15];
  assign data_masked[1987] = data_i[1987] & sel_one_hot_i[15];
  assign data_masked[1986] = data_i[1986] & sel_one_hot_i[15];
  assign data_masked[1985] = data_i[1985] & sel_one_hot_i[15];
  assign data_masked[1984] = data_i[1984] & sel_one_hot_i[15];
  assign data_masked[1983] = data_i[1983] & sel_one_hot_i[15];
  assign data_masked[1982] = data_i[1982] & sel_one_hot_i[15];
  assign data_masked[1981] = data_i[1981] & sel_one_hot_i[15];
  assign data_masked[1980] = data_i[1980] & sel_one_hot_i[15];
  assign data_masked[1979] = data_i[1979] & sel_one_hot_i[15];
  assign data_masked[1978] = data_i[1978] & sel_one_hot_i[15];
  assign data_masked[1977] = data_i[1977] & sel_one_hot_i[15];
  assign data_masked[1976] = data_i[1976] & sel_one_hot_i[15];
  assign data_masked[1975] = data_i[1975] & sel_one_hot_i[15];
  assign data_masked[1974] = data_i[1974] & sel_one_hot_i[15];
  assign data_masked[1973] = data_i[1973] & sel_one_hot_i[15];
  assign data_masked[1972] = data_i[1972] & sel_one_hot_i[15];
  assign data_masked[1971] = data_i[1971] & sel_one_hot_i[15];
  assign data_masked[1970] = data_i[1970] & sel_one_hot_i[15];
  assign data_masked[1969] = data_i[1969] & sel_one_hot_i[15];
  assign data_masked[1968] = data_i[1968] & sel_one_hot_i[15];
  assign data_masked[1967] = data_i[1967] & sel_one_hot_i[15];
  assign data_masked[1966] = data_i[1966] & sel_one_hot_i[15];
  assign data_masked[1965] = data_i[1965] & sel_one_hot_i[15];
  assign data_masked[1964] = data_i[1964] & sel_one_hot_i[15];
  assign data_masked[1963] = data_i[1963] & sel_one_hot_i[15];
  assign data_masked[1962] = data_i[1962] & sel_one_hot_i[15];
  assign data_masked[1961] = data_i[1961] & sel_one_hot_i[15];
  assign data_masked[1960] = data_i[1960] & sel_one_hot_i[15];
  assign data_masked[1959] = data_i[1959] & sel_one_hot_i[15];
  assign data_masked[1958] = data_i[1958] & sel_one_hot_i[15];
  assign data_masked[1957] = data_i[1957] & sel_one_hot_i[15];
  assign data_masked[1956] = data_i[1956] & sel_one_hot_i[15];
  assign data_masked[1955] = data_i[1955] & sel_one_hot_i[15];
  assign data_masked[1954] = data_i[1954] & sel_one_hot_i[15];
  assign data_masked[1953] = data_i[1953] & sel_one_hot_i[15];
  assign data_masked[1952] = data_i[1952] & sel_one_hot_i[15];
  assign data_masked[1951] = data_i[1951] & sel_one_hot_i[15];
  assign data_masked[1950] = data_i[1950] & sel_one_hot_i[15];
  assign data_masked[1949] = data_i[1949] & sel_one_hot_i[15];
  assign data_masked[1948] = data_i[1948] & sel_one_hot_i[15];
  assign data_masked[1947] = data_i[1947] & sel_one_hot_i[15];
  assign data_masked[1946] = data_i[1946] & sel_one_hot_i[15];
  assign data_masked[1945] = data_i[1945] & sel_one_hot_i[15];
  assign data_masked[1944] = data_i[1944] & sel_one_hot_i[15];
  assign data_masked[1943] = data_i[1943] & sel_one_hot_i[15];
  assign data_masked[1942] = data_i[1942] & sel_one_hot_i[15];
  assign data_masked[1941] = data_i[1941] & sel_one_hot_i[15];
  assign data_masked[1940] = data_i[1940] & sel_one_hot_i[15];
  assign data_masked[1939] = data_i[1939] & sel_one_hot_i[15];
  assign data_masked[1938] = data_i[1938] & sel_one_hot_i[15];
  assign data_masked[1937] = data_i[1937] & sel_one_hot_i[15];
  assign data_masked[1936] = data_i[1936] & sel_one_hot_i[15];
  assign data_masked[1935] = data_i[1935] & sel_one_hot_i[15];
  assign data_masked[1934] = data_i[1934] & sel_one_hot_i[15];
  assign data_masked[1933] = data_i[1933] & sel_one_hot_i[15];
  assign data_masked[1932] = data_i[1932] & sel_one_hot_i[15];
  assign data_masked[1931] = data_i[1931] & sel_one_hot_i[15];
  assign data_masked[1930] = data_i[1930] & sel_one_hot_i[15];
  assign data_masked[1929] = data_i[1929] & sel_one_hot_i[15];
  assign data_masked[1928] = data_i[1928] & sel_one_hot_i[15];
  assign data_masked[1927] = data_i[1927] & sel_one_hot_i[15];
  assign data_masked[1926] = data_i[1926] & sel_one_hot_i[15];
  assign data_masked[1925] = data_i[1925] & sel_one_hot_i[15];
  assign data_masked[1924] = data_i[1924] & sel_one_hot_i[15];
  assign data_masked[1923] = data_i[1923] & sel_one_hot_i[15];
  assign data_masked[1922] = data_i[1922] & sel_one_hot_i[15];
  assign data_masked[1921] = data_i[1921] & sel_one_hot_i[15];
  assign data_masked[1920] = data_i[1920] & sel_one_hot_i[15];
  assign data_masked[2175] = data_i[2175] & sel_one_hot_i[16];
  assign data_masked[2174] = data_i[2174] & sel_one_hot_i[16];
  assign data_masked[2173] = data_i[2173] & sel_one_hot_i[16];
  assign data_masked[2172] = data_i[2172] & sel_one_hot_i[16];
  assign data_masked[2171] = data_i[2171] & sel_one_hot_i[16];
  assign data_masked[2170] = data_i[2170] & sel_one_hot_i[16];
  assign data_masked[2169] = data_i[2169] & sel_one_hot_i[16];
  assign data_masked[2168] = data_i[2168] & sel_one_hot_i[16];
  assign data_masked[2167] = data_i[2167] & sel_one_hot_i[16];
  assign data_masked[2166] = data_i[2166] & sel_one_hot_i[16];
  assign data_masked[2165] = data_i[2165] & sel_one_hot_i[16];
  assign data_masked[2164] = data_i[2164] & sel_one_hot_i[16];
  assign data_masked[2163] = data_i[2163] & sel_one_hot_i[16];
  assign data_masked[2162] = data_i[2162] & sel_one_hot_i[16];
  assign data_masked[2161] = data_i[2161] & sel_one_hot_i[16];
  assign data_masked[2160] = data_i[2160] & sel_one_hot_i[16];
  assign data_masked[2159] = data_i[2159] & sel_one_hot_i[16];
  assign data_masked[2158] = data_i[2158] & sel_one_hot_i[16];
  assign data_masked[2157] = data_i[2157] & sel_one_hot_i[16];
  assign data_masked[2156] = data_i[2156] & sel_one_hot_i[16];
  assign data_masked[2155] = data_i[2155] & sel_one_hot_i[16];
  assign data_masked[2154] = data_i[2154] & sel_one_hot_i[16];
  assign data_masked[2153] = data_i[2153] & sel_one_hot_i[16];
  assign data_masked[2152] = data_i[2152] & sel_one_hot_i[16];
  assign data_masked[2151] = data_i[2151] & sel_one_hot_i[16];
  assign data_masked[2150] = data_i[2150] & sel_one_hot_i[16];
  assign data_masked[2149] = data_i[2149] & sel_one_hot_i[16];
  assign data_masked[2148] = data_i[2148] & sel_one_hot_i[16];
  assign data_masked[2147] = data_i[2147] & sel_one_hot_i[16];
  assign data_masked[2146] = data_i[2146] & sel_one_hot_i[16];
  assign data_masked[2145] = data_i[2145] & sel_one_hot_i[16];
  assign data_masked[2144] = data_i[2144] & sel_one_hot_i[16];
  assign data_masked[2143] = data_i[2143] & sel_one_hot_i[16];
  assign data_masked[2142] = data_i[2142] & sel_one_hot_i[16];
  assign data_masked[2141] = data_i[2141] & sel_one_hot_i[16];
  assign data_masked[2140] = data_i[2140] & sel_one_hot_i[16];
  assign data_masked[2139] = data_i[2139] & sel_one_hot_i[16];
  assign data_masked[2138] = data_i[2138] & sel_one_hot_i[16];
  assign data_masked[2137] = data_i[2137] & sel_one_hot_i[16];
  assign data_masked[2136] = data_i[2136] & sel_one_hot_i[16];
  assign data_masked[2135] = data_i[2135] & sel_one_hot_i[16];
  assign data_masked[2134] = data_i[2134] & sel_one_hot_i[16];
  assign data_masked[2133] = data_i[2133] & sel_one_hot_i[16];
  assign data_masked[2132] = data_i[2132] & sel_one_hot_i[16];
  assign data_masked[2131] = data_i[2131] & sel_one_hot_i[16];
  assign data_masked[2130] = data_i[2130] & sel_one_hot_i[16];
  assign data_masked[2129] = data_i[2129] & sel_one_hot_i[16];
  assign data_masked[2128] = data_i[2128] & sel_one_hot_i[16];
  assign data_masked[2127] = data_i[2127] & sel_one_hot_i[16];
  assign data_masked[2126] = data_i[2126] & sel_one_hot_i[16];
  assign data_masked[2125] = data_i[2125] & sel_one_hot_i[16];
  assign data_masked[2124] = data_i[2124] & sel_one_hot_i[16];
  assign data_masked[2123] = data_i[2123] & sel_one_hot_i[16];
  assign data_masked[2122] = data_i[2122] & sel_one_hot_i[16];
  assign data_masked[2121] = data_i[2121] & sel_one_hot_i[16];
  assign data_masked[2120] = data_i[2120] & sel_one_hot_i[16];
  assign data_masked[2119] = data_i[2119] & sel_one_hot_i[16];
  assign data_masked[2118] = data_i[2118] & sel_one_hot_i[16];
  assign data_masked[2117] = data_i[2117] & sel_one_hot_i[16];
  assign data_masked[2116] = data_i[2116] & sel_one_hot_i[16];
  assign data_masked[2115] = data_i[2115] & sel_one_hot_i[16];
  assign data_masked[2114] = data_i[2114] & sel_one_hot_i[16];
  assign data_masked[2113] = data_i[2113] & sel_one_hot_i[16];
  assign data_masked[2112] = data_i[2112] & sel_one_hot_i[16];
  assign data_masked[2111] = data_i[2111] & sel_one_hot_i[16];
  assign data_masked[2110] = data_i[2110] & sel_one_hot_i[16];
  assign data_masked[2109] = data_i[2109] & sel_one_hot_i[16];
  assign data_masked[2108] = data_i[2108] & sel_one_hot_i[16];
  assign data_masked[2107] = data_i[2107] & sel_one_hot_i[16];
  assign data_masked[2106] = data_i[2106] & sel_one_hot_i[16];
  assign data_masked[2105] = data_i[2105] & sel_one_hot_i[16];
  assign data_masked[2104] = data_i[2104] & sel_one_hot_i[16];
  assign data_masked[2103] = data_i[2103] & sel_one_hot_i[16];
  assign data_masked[2102] = data_i[2102] & sel_one_hot_i[16];
  assign data_masked[2101] = data_i[2101] & sel_one_hot_i[16];
  assign data_masked[2100] = data_i[2100] & sel_one_hot_i[16];
  assign data_masked[2099] = data_i[2099] & sel_one_hot_i[16];
  assign data_masked[2098] = data_i[2098] & sel_one_hot_i[16];
  assign data_masked[2097] = data_i[2097] & sel_one_hot_i[16];
  assign data_masked[2096] = data_i[2096] & sel_one_hot_i[16];
  assign data_masked[2095] = data_i[2095] & sel_one_hot_i[16];
  assign data_masked[2094] = data_i[2094] & sel_one_hot_i[16];
  assign data_masked[2093] = data_i[2093] & sel_one_hot_i[16];
  assign data_masked[2092] = data_i[2092] & sel_one_hot_i[16];
  assign data_masked[2091] = data_i[2091] & sel_one_hot_i[16];
  assign data_masked[2090] = data_i[2090] & sel_one_hot_i[16];
  assign data_masked[2089] = data_i[2089] & sel_one_hot_i[16];
  assign data_masked[2088] = data_i[2088] & sel_one_hot_i[16];
  assign data_masked[2087] = data_i[2087] & sel_one_hot_i[16];
  assign data_masked[2086] = data_i[2086] & sel_one_hot_i[16];
  assign data_masked[2085] = data_i[2085] & sel_one_hot_i[16];
  assign data_masked[2084] = data_i[2084] & sel_one_hot_i[16];
  assign data_masked[2083] = data_i[2083] & sel_one_hot_i[16];
  assign data_masked[2082] = data_i[2082] & sel_one_hot_i[16];
  assign data_masked[2081] = data_i[2081] & sel_one_hot_i[16];
  assign data_masked[2080] = data_i[2080] & sel_one_hot_i[16];
  assign data_masked[2079] = data_i[2079] & sel_one_hot_i[16];
  assign data_masked[2078] = data_i[2078] & sel_one_hot_i[16];
  assign data_masked[2077] = data_i[2077] & sel_one_hot_i[16];
  assign data_masked[2076] = data_i[2076] & sel_one_hot_i[16];
  assign data_masked[2075] = data_i[2075] & sel_one_hot_i[16];
  assign data_masked[2074] = data_i[2074] & sel_one_hot_i[16];
  assign data_masked[2073] = data_i[2073] & sel_one_hot_i[16];
  assign data_masked[2072] = data_i[2072] & sel_one_hot_i[16];
  assign data_masked[2071] = data_i[2071] & sel_one_hot_i[16];
  assign data_masked[2070] = data_i[2070] & sel_one_hot_i[16];
  assign data_masked[2069] = data_i[2069] & sel_one_hot_i[16];
  assign data_masked[2068] = data_i[2068] & sel_one_hot_i[16];
  assign data_masked[2067] = data_i[2067] & sel_one_hot_i[16];
  assign data_masked[2066] = data_i[2066] & sel_one_hot_i[16];
  assign data_masked[2065] = data_i[2065] & sel_one_hot_i[16];
  assign data_masked[2064] = data_i[2064] & sel_one_hot_i[16];
  assign data_masked[2063] = data_i[2063] & sel_one_hot_i[16];
  assign data_masked[2062] = data_i[2062] & sel_one_hot_i[16];
  assign data_masked[2061] = data_i[2061] & sel_one_hot_i[16];
  assign data_masked[2060] = data_i[2060] & sel_one_hot_i[16];
  assign data_masked[2059] = data_i[2059] & sel_one_hot_i[16];
  assign data_masked[2058] = data_i[2058] & sel_one_hot_i[16];
  assign data_masked[2057] = data_i[2057] & sel_one_hot_i[16];
  assign data_masked[2056] = data_i[2056] & sel_one_hot_i[16];
  assign data_masked[2055] = data_i[2055] & sel_one_hot_i[16];
  assign data_masked[2054] = data_i[2054] & sel_one_hot_i[16];
  assign data_masked[2053] = data_i[2053] & sel_one_hot_i[16];
  assign data_masked[2052] = data_i[2052] & sel_one_hot_i[16];
  assign data_masked[2051] = data_i[2051] & sel_one_hot_i[16];
  assign data_masked[2050] = data_i[2050] & sel_one_hot_i[16];
  assign data_masked[2049] = data_i[2049] & sel_one_hot_i[16];
  assign data_masked[2048] = data_i[2048] & sel_one_hot_i[16];
  assign data_masked[2303] = data_i[2303] & sel_one_hot_i[17];
  assign data_masked[2302] = data_i[2302] & sel_one_hot_i[17];
  assign data_masked[2301] = data_i[2301] & sel_one_hot_i[17];
  assign data_masked[2300] = data_i[2300] & sel_one_hot_i[17];
  assign data_masked[2299] = data_i[2299] & sel_one_hot_i[17];
  assign data_masked[2298] = data_i[2298] & sel_one_hot_i[17];
  assign data_masked[2297] = data_i[2297] & sel_one_hot_i[17];
  assign data_masked[2296] = data_i[2296] & sel_one_hot_i[17];
  assign data_masked[2295] = data_i[2295] & sel_one_hot_i[17];
  assign data_masked[2294] = data_i[2294] & sel_one_hot_i[17];
  assign data_masked[2293] = data_i[2293] & sel_one_hot_i[17];
  assign data_masked[2292] = data_i[2292] & sel_one_hot_i[17];
  assign data_masked[2291] = data_i[2291] & sel_one_hot_i[17];
  assign data_masked[2290] = data_i[2290] & sel_one_hot_i[17];
  assign data_masked[2289] = data_i[2289] & sel_one_hot_i[17];
  assign data_masked[2288] = data_i[2288] & sel_one_hot_i[17];
  assign data_masked[2287] = data_i[2287] & sel_one_hot_i[17];
  assign data_masked[2286] = data_i[2286] & sel_one_hot_i[17];
  assign data_masked[2285] = data_i[2285] & sel_one_hot_i[17];
  assign data_masked[2284] = data_i[2284] & sel_one_hot_i[17];
  assign data_masked[2283] = data_i[2283] & sel_one_hot_i[17];
  assign data_masked[2282] = data_i[2282] & sel_one_hot_i[17];
  assign data_masked[2281] = data_i[2281] & sel_one_hot_i[17];
  assign data_masked[2280] = data_i[2280] & sel_one_hot_i[17];
  assign data_masked[2279] = data_i[2279] & sel_one_hot_i[17];
  assign data_masked[2278] = data_i[2278] & sel_one_hot_i[17];
  assign data_masked[2277] = data_i[2277] & sel_one_hot_i[17];
  assign data_masked[2276] = data_i[2276] & sel_one_hot_i[17];
  assign data_masked[2275] = data_i[2275] & sel_one_hot_i[17];
  assign data_masked[2274] = data_i[2274] & sel_one_hot_i[17];
  assign data_masked[2273] = data_i[2273] & sel_one_hot_i[17];
  assign data_masked[2272] = data_i[2272] & sel_one_hot_i[17];
  assign data_masked[2271] = data_i[2271] & sel_one_hot_i[17];
  assign data_masked[2270] = data_i[2270] & sel_one_hot_i[17];
  assign data_masked[2269] = data_i[2269] & sel_one_hot_i[17];
  assign data_masked[2268] = data_i[2268] & sel_one_hot_i[17];
  assign data_masked[2267] = data_i[2267] & sel_one_hot_i[17];
  assign data_masked[2266] = data_i[2266] & sel_one_hot_i[17];
  assign data_masked[2265] = data_i[2265] & sel_one_hot_i[17];
  assign data_masked[2264] = data_i[2264] & sel_one_hot_i[17];
  assign data_masked[2263] = data_i[2263] & sel_one_hot_i[17];
  assign data_masked[2262] = data_i[2262] & sel_one_hot_i[17];
  assign data_masked[2261] = data_i[2261] & sel_one_hot_i[17];
  assign data_masked[2260] = data_i[2260] & sel_one_hot_i[17];
  assign data_masked[2259] = data_i[2259] & sel_one_hot_i[17];
  assign data_masked[2258] = data_i[2258] & sel_one_hot_i[17];
  assign data_masked[2257] = data_i[2257] & sel_one_hot_i[17];
  assign data_masked[2256] = data_i[2256] & sel_one_hot_i[17];
  assign data_masked[2255] = data_i[2255] & sel_one_hot_i[17];
  assign data_masked[2254] = data_i[2254] & sel_one_hot_i[17];
  assign data_masked[2253] = data_i[2253] & sel_one_hot_i[17];
  assign data_masked[2252] = data_i[2252] & sel_one_hot_i[17];
  assign data_masked[2251] = data_i[2251] & sel_one_hot_i[17];
  assign data_masked[2250] = data_i[2250] & sel_one_hot_i[17];
  assign data_masked[2249] = data_i[2249] & sel_one_hot_i[17];
  assign data_masked[2248] = data_i[2248] & sel_one_hot_i[17];
  assign data_masked[2247] = data_i[2247] & sel_one_hot_i[17];
  assign data_masked[2246] = data_i[2246] & sel_one_hot_i[17];
  assign data_masked[2245] = data_i[2245] & sel_one_hot_i[17];
  assign data_masked[2244] = data_i[2244] & sel_one_hot_i[17];
  assign data_masked[2243] = data_i[2243] & sel_one_hot_i[17];
  assign data_masked[2242] = data_i[2242] & sel_one_hot_i[17];
  assign data_masked[2241] = data_i[2241] & sel_one_hot_i[17];
  assign data_masked[2240] = data_i[2240] & sel_one_hot_i[17];
  assign data_masked[2239] = data_i[2239] & sel_one_hot_i[17];
  assign data_masked[2238] = data_i[2238] & sel_one_hot_i[17];
  assign data_masked[2237] = data_i[2237] & sel_one_hot_i[17];
  assign data_masked[2236] = data_i[2236] & sel_one_hot_i[17];
  assign data_masked[2235] = data_i[2235] & sel_one_hot_i[17];
  assign data_masked[2234] = data_i[2234] & sel_one_hot_i[17];
  assign data_masked[2233] = data_i[2233] & sel_one_hot_i[17];
  assign data_masked[2232] = data_i[2232] & sel_one_hot_i[17];
  assign data_masked[2231] = data_i[2231] & sel_one_hot_i[17];
  assign data_masked[2230] = data_i[2230] & sel_one_hot_i[17];
  assign data_masked[2229] = data_i[2229] & sel_one_hot_i[17];
  assign data_masked[2228] = data_i[2228] & sel_one_hot_i[17];
  assign data_masked[2227] = data_i[2227] & sel_one_hot_i[17];
  assign data_masked[2226] = data_i[2226] & sel_one_hot_i[17];
  assign data_masked[2225] = data_i[2225] & sel_one_hot_i[17];
  assign data_masked[2224] = data_i[2224] & sel_one_hot_i[17];
  assign data_masked[2223] = data_i[2223] & sel_one_hot_i[17];
  assign data_masked[2222] = data_i[2222] & sel_one_hot_i[17];
  assign data_masked[2221] = data_i[2221] & sel_one_hot_i[17];
  assign data_masked[2220] = data_i[2220] & sel_one_hot_i[17];
  assign data_masked[2219] = data_i[2219] & sel_one_hot_i[17];
  assign data_masked[2218] = data_i[2218] & sel_one_hot_i[17];
  assign data_masked[2217] = data_i[2217] & sel_one_hot_i[17];
  assign data_masked[2216] = data_i[2216] & sel_one_hot_i[17];
  assign data_masked[2215] = data_i[2215] & sel_one_hot_i[17];
  assign data_masked[2214] = data_i[2214] & sel_one_hot_i[17];
  assign data_masked[2213] = data_i[2213] & sel_one_hot_i[17];
  assign data_masked[2212] = data_i[2212] & sel_one_hot_i[17];
  assign data_masked[2211] = data_i[2211] & sel_one_hot_i[17];
  assign data_masked[2210] = data_i[2210] & sel_one_hot_i[17];
  assign data_masked[2209] = data_i[2209] & sel_one_hot_i[17];
  assign data_masked[2208] = data_i[2208] & sel_one_hot_i[17];
  assign data_masked[2207] = data_i[2207] & sel_one_hot_i[17];
  assign data_masked[2206] = data_i[2206] & sel_one_hot_i[17];
  assign data_masked[2205] = data_i[2205] & sel_one_hot_i[17];
  assign data_masked[2204] = data_i[2204] & sel_one_hot_i[17];
  assign data_masked[2203] = data_i[2203] & sel_one_hot_i[17];
  assign data_masked[2202] = data_i[2202] & sel_one_hot_i[17];
  assign data_masked[2201] = data_i[2201] & sel_one_hot_i[17];
  assign data_masked[2200] = data_i[2200] & sel_one_hot_i[17];
  assign data_masked[2199] = data_i[2199] & sel_one_hot_i[17];
  assign data_masked[2198] = data_i[2198] & sel_one_hot_i[17];
  assign data_masked[2197] = data_i[2197] & sel_one_hot_i[17];
  assign data_masked[2196] = data_i[2196] & sel_one_hot_i[17];
  assign data_masked[2195] = data_i[2195] & sel_one_hot_i[17];
  assign data_masked[2194] = data_i[2194] & sel_one_hot_i[17];
  assign data_masked[2193] = data_i[2193] & sel_one_hot_i[17];
  assign data_masked[2192] = data_i[2192] & sel_one_hot_i[17];
  assign data_masked[2191] = data_i[2191] & sel_one_hot_i[17];
  assign data_masked[2190] = data_i[2190] & sel_one_hot_i[17];
  assign data_masked[2189] = data_i[2189] & sel_one_hot_i[17];
  assign data_masked[2188] = data_i[2188] & sel_one_hot_i[17];
  assign data_masked[2187] = data_i[2187] & sel_one_hot_i[17];
  assign data_masked[2186] = data_i[2186] & sel_one_hot_i[17];
  assign data_masked[2185] = data_i[2185] & sel_one_hot_i[17];
  assign data_masked[2184] = data_i[2184] & sel_one_hot_i[17];
  assign data_masked[2183] = data_i[2183] & sel_one_hot_i[17];
  assign data_masked[2182] = data_i[2182] & sel_one_hot_i[17];
  assign data_masked[2181] = data_i[2181] & sel_one_hot_i[17];
  assign data_masked[2180] = data_i[2180] & sel_one_hot_i[17];
  assign data_masked[2179] = data_i[2179] & sel_one_hot_i[17];
  assign data_masked[2178] = data_i[2178] & sel_one_hot_i[17];
  assign data_masked[2177] = data_i[2177] & sel_one_hot_i[17];
  assign data_masked[2176] = data_i[2176] & sel_one_hot_i[17];
  assign data_masked[2431] = data_i[2431] & sel_one_hot_i[18];
  assign data_masked[2430] = data_i[2430] & sel_one_hot_i[18];
  assign data_masked[2429] = data_i[2429] & sel_one_hot_i[18];
  assign data_masked[2428] = data_i[2428] & sel_one_hot_i[18];
  assign data_masked[2427] = data_i[2427] & sel_one_hot_i[18];
  assign data_masked[2426] = data_i[2426] & sel_one_hot_i[18];
  assign data_masked[2425] = data_i[2425] & sel_one_hot_i[18];
  assign data_masked[2424] = data_i[2424] & sel_one_hot_i[18];
  assign data_masked[2423] = data_i[2423] & sel_one_hot_i[18];
  assign data_masked[2422] = data_i[2422] & sel_one_hot_i[18];
  assign data_masked[2421] = data_i[2421] & sel_one_hot_i[18];
  assign data_masked[2420] = data_i[2420] & sel_one_hot_i[18];
  assign data_masked[2419] = data_i[2419] & sel_one_hot_i[18];
  assign data_masked[2418] = data_i[2418] & sel_one_hot_i[18];
  assign data_masked[2417] = data_i[2417] & sel_one_hot_i[18];
  assign data_masked[2416] = data_i[2416] & sel_one_hot_i[18];
  assign data_masked[2415] = data_i[2415] & sel_one_hot_i[18];
  assign data_masked[2414] = data_i[2414] & sel_one_hot_i[18];
  assign data_masked[2413] = data_i[2413] & sel_one_hot_i[18];
  assign data_masked[2412] = data_i[2412] & sel_one_hot_i[18];
  assign data_masked[2411] = data_i[2411] & sel_one_hot_i[18];
  assign data_masked[2410] = data_i[2410] & sel_one_hot_i[18];
  assign data_masked[2409] = data_i[2409] & sel_one_hot_i[18];
  assign data_masked[2408] = data_i[2408] & sel_one_hot_i[18];
  assign data_masked[2407] = data_i[2407] & sel_one_hot_i[18];
  assign data_masked[2406] = data_i[2406] & sel_one_hot_i[18];
  assign data_masked[2405] = data_i[2405] & sel_one_hot_i[18];
  assign data_masked[2404] = data_i[2404] & sel_one_hot_i[18];
  assign data_masked[2403] = data_i[2403] & sel_one_hot_i[18];
  assign data_masked[2402] = data_i[2402] & sel_one_hot_i[18];
  assign data_masked[2401] = data_i[2401] & sel_one_hot_i[18];
  assign data_masked[2400] = data_i[2400] & sel_one_hot_i[18];
  assign data_masked[2399] = data_i[2399] & sel_one_hot_i[18];
  assign data_masked[2398] = data_i[2398] & sel_one_hot_i[18];
  assign data_masked[2397] = data_i[2397] & sel_one_hot_i[18];
  assign data_masked[2396] = data_i[2396] & sel_one_hot_i[18];
  assign data_masked[2395] = data_i[2395] & sel_one_hot_i[18];
  assign data_masked[2394] = data_i[2394] & sel_one_hot_i[18];
  assign data_masked[2393] = data_i[2393] & sel_one_hot_i[18];
  assign data_masked[2392] = data_i[2392] & sel_one_hot_i[18];
  assign data_masked[2391] = data_i[2391] & sel_one_hot_i[18];
  assign data_masked[2390] = data_i[2390] & sel_one_hot_i[18];
  assign data_masked[2389] = data_i[2389] & sel_one_hot_i[18];
  assign data_masked[2388] = data_i[2388] & sel_one_hot_i[18];
  assign data_masked[2387] = data_i[2387] & sel_one_hot_i[18];
  assign data_masked[2386] = data_i[2386] & sel_one_hot_i[18];
  assign data_masked[2385] = data_i[2385] & sel_one_hot_i[18];
  assign data_masked[2384] = data_i[2384] & sel_one_hot_i[18];
  assign data_masked[2383] = data_i[2383] & sel_one_hot_i[18];
  assign data_masked[2382] = data_i[2382] & sel_one_hot_i[18];
  assign data_masked[2381] = data_i[2381] & sel_one_hot_i[18];
  assign data_masked[2380] = data_i[2380] & sel_one_hot_i[18];
  assign data_masked[2379] = data_i[2379] & sel_one_hot_i[18];
  assign data_masked[2378] = data_i[2378] & sel_one_hot_i[18];
  assign data_masked[2377] = data_i[2377] & sel_one_hot_i[18];
  assign data_masked[2376] = data_i[2376] & sel_one_hot_i[18];
  assign data_masked[2375] = data_i[2375] & sel_one_hot_i[18];
  assign data_masked[2374] = data_i[2374] & sel_one_hot_i[18];
  assign data_masked[2373] = data_i[2373] & sel_one_hot_i[18];
  assign data_masked[2372] = data_i[2372] & sel_one_hot_i[18];
  assign data_masked[2371] = data_i[2371] & sel_one_hot_i[18];
  assign data_masked[2370] = data_i[2370] & sel_one_hot_i[18];
  assign data_masked[2369] = data_i[2369] & sel_one_hot_i[18];
  assign data_masked[2368] = data_i[2368] & sel_one_hot_i[18];
  assign data_masked[2367] = data_i[2367] & sel_one_hot_i[18];
  assign data_masked[2366] = data_i[2366] & sel_one_hot_i[18];
  assign data_masked[2365] = data_i[2365] & sel_one_hot_i[18];
  assign data_masked[2364] = data_i[2364] & sel_one_hot_i[18];
  assign data_masked[2363] = data_i[2363] & sel_one_hot_i[18];
  assign data_masked[2362] = data_i[2362] & sel_one_hot_i[18];
  assign data_masked[2361] = data_i[2361] & sel_one_hot_i[18];
  assign data_masked[2360] = data_i[2360] & sel_one_hot_i[18];
  assign data_masked[2359] = data_i[2359] & sel_one_hot_i[18];
  assign data_masked[2358] = data_i[2358] & sel_one_hot_i[18];
  assign data_masked[2357] = data_i[2357] & sel_one_hot_i[18];
  assign data_masked[2356] = data_i[2356] & sel_one_hot_i[18];
  assign data_masked[2355] = data_i[2355] & sel_one_hot_i[18];
  assign data_masked[2354] = data_i[2354] & sel_one_hot_i[18];
  assign data_masked[2353] = data_i[2353] & sel_one_hot_i[18];
  assign data_masked[2352] = data_i[2352] & sel_one_hot_i[18];
  assign data_masked[2351] = data_i[2351] & sel_one_hot_i[18];
  assign data_masked[2350] = data_i[2350] & sel_one_hot_i[18];
  assign data_masked[2349] = data_i[2349] & sel_one_hot_i[18];
  assign data_masked[2348] = data_i[2348] & sel_one_hot_i[18];
  assign data_masked[2347] = data_i[2347] & sel_one_hot_i[18];
  assign data_masked[2346] = data_i[2346] & sel_one_hot_i[18];
  assign data_masked[2345] = data_i[2345] & sel_one_hot_i[18];
  assign data_masked[2344] = data_i[2344] & sel_one_hot_i[18];
  assign data_masked[2343] = data_i[2343] & sel_one_hot_i[18];
  assign data_masked[2342] = data_i[2342] & sel_one_hot_i[18];
  assign data_masked[2341] = data_i[2341] & sel_one_hot_i[18];
  assign data_masked[2340] = data_i[2340] & sel_one_hot_i[18];
  assign data_masked[2339] = data_i[2339] & sel_one_hot_i[18];
  assign data_masked[2338] = data_i[2338] & sel_one_hot_i[18];
  assign data_masked[2337] = data_i[2337] & sel_one_hot_i[18];
  assign data_masked[2336] = data_i[2336] & sel_one_hot_i[18];
  assign data_masked[2335] = data_i[2335] & sel_one_hot_i[18];
  assign data_masked[2334] = data_i[2334] & sel_one_hot_i[18];
  assign data_masked[2333] = data_i[2333] & sel_one_hot_i[18];
  assign data_masked[2332] = data_i[2332] & sel_one_hot_i[18];
  assign data_masked[2331] = data_i[2331] & sel_one_hot_i[18];
  assign data_masked[2330] = data_i[2330] & sel_one_hot_i[18];
  assign data_masked[2329] = data_i[2329] & sel_one_hot_i[18];
  assign data_masked[2328] = data_i[2328] & sel_one_hot_i[18];
  assign data_masked[2327] = data_i[2327] & sel_one_hot_i[18];
  assign data_masked[2326] = data_i[2326] & sel_one_hot_i[18];
  assign data_masked[2325] = data_i[2325] & sel_one_hot_i[18];
  assign data_masked[2324] = data_i[2324] & sel_one_hot_i[18];
  assign data_masked[2323] = data_i[2323] & sel_one_hot_i[18];
  assign data_masked[2322] = data_i[2322] & sel_one_hot_i[18];
  assign data_masked[2321] = data_i[2321] & sel_one_hot_i[18];
  assign data_masked[2320] = data_i[2320] & sel_one_hot_i[18];
  assign data_masked[2319] = data_i[2319] & sel_one_hot_i[18];
  assign data_masked[2318] = data_i[2318] & sel_one_hot_i[18];
  assign data_masked[2317] = data_i[2317] & sel_one_hot_i[18];
  assign data_masked[2316] = data_i[2316] & sel_one_hot_i[18];
  assign data_masked[2315] = data_i[2315] & sel_one_hot_i[18];
  assign data_masked[2314] = data_i[2314] & sel_one_hot_i[18];
  assign data_masked[2313] = data_i[2313] & sel_one_hot_i[18];
  assign data_masked[2312] = data_i[2312] & sel_one_hot_i[18];
  assign data_masked[2311] = data_i[2311] & sel_one_hot_i[18];
  assign data_masked[2310] = data_i[2310] & sel_one_hot_i[18];
  assign data_masked[2309] = data_i[2309] & sel_one_hot_i[18];
  assign data_masked[2308] = data_i[2308] & sel_one_hot_i[18];
  assign data_masked[2307] = data_i[2307] & sel_one_hot_i[18];
  assign data_masked[2306] = data_i[2306] & sel_one_hot_i[18];
  assign data_masked[2305] = data_i[2305] & sel_one_hot_i[18];
  assign data_masked[2304] = data_i[2304] & sel_one_hot_i[18];
  assign data_masked[2559] = data_i[2559] & sel_one_hot_i[19];
  assign data_masked[2558] = data_i[2558] & sel_one_hot_i[19];
  assign data_masked[2557] = data_i[2557] & sel_one_hot_i[19];
  assign data_masked[2556] = data_i[2556] & sel_one_hot_i[19];
  assign data_masked[2555] = data_i[2555] & sel_one_hot_i[19];
  assign data_masked[2554] = data_i[2554] & sel_one_hot_i[19];
  assign data_masked[2553] = data_i[2553] & sel_one_hot_i[19];
  assign data_masked[2552] = data_i[2552] & sel_one_hot_i[19];
  assign data_masked[2551] = data_i[2551] & sel_one_hot_i[19];
  assign data_masked[2550] = data_i[2550] & sel_one_hot_i[19];
  assign data_masked[2549] = data_i[2549] & sel_one_hot_i[19];
  assign data_masked[2548] = data_i[2548] & sel_one_hot_i[19];
  assign data_masked[2547] = data_i[2547] & sel_one_hot_i[19];
  assign data_masked[2546] = data_i[2546] & sel_one_hot_i[19];
  assign data_masked[2545] = data_i[2545] & sel_one_hot_i[19];
  assign data_masked[2544] = data_i[2544] & sel_one_hot_i[19];
  assign data_masked[2543] = data_i[2543] & sel_one_hot_i[19];
  assign data_masked[2542] = data_i[2542] & sel_one_hot_i[19];
  assign data_masked[2541] = data_i[2541] & sel_one_hot_i[19];
  assign data_masked[2540] = data_i[2540] & sel_one_hot_i[19];
  assign data_masked[2539] = data_i[2539] & sel_one_hot_i[19];
  assign data_masked[2538] = data_i[2538] & sel_one_hot_i[19];
  assign data_masked[2537] = data_i[2537] & sel_one_hot_i[19];
  assign data_masked[2536] = data_i[2536] & sel_one_hot_i[19];
  assign data_masked[2535] = data_i[2535] & sel_one_hot_i[19];
  assign data_masked[2534] = data_i[2534] & sel_one_hot_i[19];
  assign data_masked[2533] = data_i[2533] & sel_one_hot_i[19];
  assign data_masked[2532] = data_i[2532] & sel_one_hot_i[19];
  assign data_masked[2531] = data_i[2531] & sel_one_hot_i[19];
  assign data_masked[2530] = data_i[2530] & sel_one_hot_i[19];
  assign data_masked[2529] = data_i[2529] & sel_one_hot_i[19];
  assign data_masked[2528] = data_i[2528] & sel_one_hot_i[19];
  assign data_masked[2527] = data_i[2527] & sel_one_hot_i[19];
  assign data_masked[2526] = data_i[2526] & sel_one_hot_i[19];
  assign data_masked[2525] = data_i[2525] & sel_one_hot_i[19];
  assign data_masked[2524] = data_i[2524] & sel_one_hot_i[19];
  assign data_masked[2523] = data_i[2523] & sel_one_hot_i[19];
  assign data_masked[2522] = data_i[2522] & sel_one_hot_i[19];
  assign data_masked[2521] = data_i[2521] & sel_one_hot_i[19];
  assign data_masked[2520] = data_i[2520] & sel_one_hot_i[19];
  assign data_masked[2519] = data_i[2519] & sel_one_hot_i[19];
  assign data_masked[2518] = data_i[2518] & sel_one_hot_i[19];
  assign data_masked[2517] = data_i[2517] & sel_one_hot_i[19];
  assign data_masked[2516] = data_i[2516] & sel_one_hot_i[19];
  assign data_masked[2515] = data_i[2515] & sel_one_hot_i[19];
  assign data_masked[2514] = data_i[2514] & sel_one_hot_i[19];
  assign data_masked[2513] = data_i[2513] & sel_one_hot_i[19];
  assign data_masked[2512] = data_i[2512] & sel_one_hot_i[19];
  assign data_masked[2511] = data_i[2511] & sel_one_hot_i[19];
  assign data_masked[2510] = data_i[2510] & sel_one_hot_i[19];
  assign data_masked[2509] = data_i[2509] & sel_one_hot_i[19];
  assign data_masked[2508] = data_i[2508] & sel_one_hot_i[19];
  assign data_masked[2507] = data_i[2507] & sel_one_hot_i[19];
  assign data_masked[2506] = data_i[2506] & sel_one_hot_i[19];
  assign data_masked[2505] = data_i[2505] & sel_one_hot_i[19];
  assign data_masked[2504] = data_i[2504] & sel_one_hot_i[19];
  assign data_masked[2503] = data_i[2503] & sel_one_hot_i[19];
  assign data_masked[2502] = data_i[2502] & sel_one_hot_i[19];
  assign data_masked[2501] = data_i[2501] & sel_one_hot_i[19];
  assign data_masked[2500] = data_i[2500] & sel_one_hot_i[19];
  assign data_masked[2499] = data_i[2499] & sel_one_hot_i[19];
  assign data_masked[2498] = data_i[2498] & sel_one_hot_i[19];
  assign data_masked[2497] = data_i[2497] & sel_one_hot_i[19];
  assign data_masked[2496] = data_i[2496] & sel_one_hot_i[19];
  assign data_masked[2495] = data_i[2495] & sel_one_hot_i[19];
  assign data_masked[2494] = data_i[2494] & sel_one_hot_i[19];
  assign data_masked[2493] = data_i[2493] & sel_one_hot_i[19];
  assign data_masked[2492] = data_i[2492] & sel_one_hot_i[19];
  assign data_masked[2491] = data_i[2491] & sel_one_hot_i[19];
  assign data_masked[2490] = data_i[2490] & sel_one_hot_i[19];
  assign data_masked[2489] = data_i[2489] & sel_one_hot_i[19];
  assign data_masked[2488] = data_i[2488] & sel_one_hot_i[19];
  assign data_masked[2487] = data_i[2487] & sel_one_hot_i[19];
  assign data_masked[2486] = data_i[2486] & sel_one_hot_i[19];
  assign data_masked[2485] = data_i[2485] & sel_one_hot_i[19];
  assign data_masked[2484] = data_i[2484] & sel_one_hot_i[19];
  assign data_masked[2483] = data_i[2483] & sel_one_hot_i[19];
  assign data_masked[2482] = data_i[2482] & sel_one_hot_i[19];
  assign data_masked[2481] = data_i[2481] & sel_one_hot_i[19];
  assign data_masked[2480] = data_i[2480] & sel_one_hot_i[19];
  assign data_masked[2479] = data_i[2479] & sel_one_hot_i[19];
  assign data_masked[2478] = data_i[2478] & sel_one_hot_i[19];
  assign data_masked[2477] = data_i[2477] & sel_one_hot_i[19];
  assign data_masked[2476] = data_i[2476] & sel_one_hot_i[19];
  assign data_masked[2475] = data_i[2475] & sel_one_hot_i[19];
  assign data_masked[2474] = data_i[2474] & sel_one_hot_i[19];
  assign data_masked[2473] = data_i[2473] & sel_one_hot_i[19];
  assign data_masked[2472] = data_i[2472] & sel_one_hot_i[19];
  assign data_masked[2471] = data_i[2471] & sel_one_hot_i[19];
  assign data_masked[2470] = data_i[2470] & sel_one_hot_i[19];
  assign data_masked[2469] = data_i[2469] & sel_one_hot_i[19];
  assign data_masked[2468] = data_i[2468] & sel_one_hot_i[19];
  assign data_masked[2467] = data_i[2467] & sel_one_hot_i[19];
  assign data_masked[2466] = data_i[2466] & sel_one_hot_i[19];
  assign data_masked[2465] = data_i[2465] & sel_one_hot_i[19];
  assign data_masked[2464] = data_i[2464] & sel_one_hot_i[19];
  assign data_masked[2463] = data_i[2463] & sel_one_hot_i[19];
  assign data_masked[2462] = data_i[2462] & sel_one_hot_i[19];
  assign data_masked[2461] = data_i[2461] & sel_one_hot_i[19];
  assign data_masked[2460] = data_i[2460] & sel_one_hot_i[19];
  assign data_masked[2459] = data_i[2459] & sel_one_hot_i[19];
  assign data_masked[2458] = data_i[2458] & sel_one_hot_i[19];
  assign data_masked[2457] = data_i[2457] & sel_one_hot_i[19];
  assign data_masked[2456] = data_i[2456] & sel_one_hot_i[19];
  assign data_masked[2455] = data_i[2455] & sel_one_hot_i[19];
  assign data_masked[2454] = data_i[2454] & sel_one_hot_i[19];
  assign data_masked[2453] = data_i[2453] & sel_one_hot_i[19];
  assign data_masked[2452] = data_i[2452] & sel_one_hot_i[19];
  assign data_masked[2451] = data_i[2451] & sel_one_hot_i[19];
  assign data_masked[2450] = data_i[2450] & sel_one_hot_i[19];
  assign data_masked[2449] = data_i[2449] & sel_one_hot_i[19];
  assign data_masked[2448] = data_i[2448] & sel_one_hot_i[19];
  assign data_masked[2447] = data_i[2447] & sel_one_hot_i[19];
  assign data_masked[2446] = data_i[2446] & sel_one_hot_i[19];
  assign data_masked[2445] = data_i[2445] & sel_one_hot_i[19];
  assign data_masked[2444] = data_i[2444] & sel_one_hot_i[19];
  assign data_masked[2443] = data_i[2443] & sel_one_hot_i[19];
  assign data_masked[2442] = data_i[2442] & sel_one_hot_i[19];
  assign data_masked[2441] = data_i[2441] & sel_one_hot_i[19];
  assign data_masked[2440] = data_i[2440] & sel_one_hot_i[19];
  assign data_masked[2439] = data_i[2439] & sel_one_hot_i[19];
  assign data_masked[2438] = data_i[2438] & sel_one_hot_i[19];
  assign data_masked[2437] = data_i[2437] & sel_one_hot_i[19];
  assign data_masked[2436] = data_i[2436] & sel_one_hot_i[19];
  assign data_masked[2435] = data_i[2435] & sel_one_hot_i[19];
  assign data_masked[2434] = data_i[2434] & sel_one_hot_i[19];
  assign data_masked[2433] = data_i[2433] & sel_one_hot_i[19];
  assign data_masked[2432] = data_i[2432] & sel_one_hot_i[19];
  assign data_masked[2687] = data_i[2687] & sel_one_hot_i[20];
  assign data_masked[2686] = data_i[2686] & sel_one_hot_i[20];
  assign data_masked[2685] = data_i[2685] & sel_one_hot_i[20];
  assign data_masked[2684] = data_i[2684] & sel_one_hot_i[20];
  assign data_masked[2683] = data_i[2683] & sel_one_hot_i[20];
  assign data_masked[2682] = data_i[2682] & sel_one_hot_i[20];
  assign data_masked[2681] = data_i[2681] & sel_one_hot_i[20];
  assign data_masked[2680] = data_i[2680] & sel_one_hot_i[20];
  assign data_masked[2679] = data_i[2679] & sel_one_hot_i[20];
  assign data_masked[2678] = data_i[2678] & sel_one_hot_i[20];
  assign data_masked[2677] = data_i[2677] & sel_one_hot_i[20];
  assign data_masked[2676] = data_i[2676] & sel_one_hot_i[20];
  assign data_masked[2675] = data_i[2675] & sel_one_hot_i[20];
  assign data_masked[2674] = data_i[2674] & sel_one_hot_i[20];
  assign data_masked[2673] = data_i[2673] & sel_one_hot_i[20];
  assign data_masked[2672] = data_i[2672] & sel_one_hot_i[20];
  assign data_masked[2671] = data_i[2671] & sel_one_hot_i[20];
  assign data_masked[2670] = data_i[2670] & sel_one_hot_i[20];
  assign data_masked[2669] = data_i[2669] & sel_one_hot_i[20];
  assign data_masked[2668] = data_i[2668] & sel_one_hot_i[20];
  assign data_masked[2667] = data_i[2667] & sel_one_hot_i[20];
  assign data_masked[2666] = data_i[2666] & sel_one_hot_i[20];
  assign data_masked[2665] = data_i[2665] & sel_one_hot_i[20];
  assign data_masked[2664] = data_i[2664] & sel_one_hot_i[20];
  assign data_masked[2663] = data_i[2663] & sel_one_hot_i[20];
  assign data_masked[2662] = data_i[2662] & sel_one_hot_i[20];
  assign data_masked[2661] = data_i[2661] & sel_one_hot_i[20];
  assign data_masked[2660] = data_i[2660] & sel_one_hot_i[20];
  assign data_masked[2659] = data_i[2659] & sel_one_hot_i[20];
  assign data_masked[2658] = data_i[2658] & sel_one_hot_i[20];
  assign data_masked[2657] = data_i[2657] & sel_one_hot_i[20];
  assign data_masked[2656] = data_i[2656] & sel_one_hot_i[20];
  assign data_masked[2655] = data_i[2655] & sel_one_hot_i[20];
  assign data_masked[2654] = data_i[2654] & sel_one_hot_i[20];
  assign data_masked[2653] = data_i[2653] & sel_one_hot_i[20];
  assign data_masked[2652] = data_i[2652] & sel_one_hot_i[20];
  assign data_masked[2651] = data_i[2651] & sel_one_hot_i[20];
  assign data_masked[2650] = data_i[2650] & sel_one_hot_i[20];
  assign data_masked[2649] = data_i[2649] & sel_one_hot_i[20];
  assign data_masked[2648] = data_i[2648] & sel_one_hot_i[20];
  assign data_masked[2647] = data_i[2647] & sel_one_hot_i[20];
  assign data_masked[2646] = data_i[2646] & sel_one_hot_i[20];
  assign data_masked[2645] = data_i[2645] & sel_one_hot_i[20];
  assign data_masked[2644] = data_i[2644] & sel_one_hot_i[20];
  assign data_masked[2643] = data_i[2643] & sel_one_hot_i[20];
  assign data_masked[2642] = data_i[2642] & sel_one_hot_i[20];
  assign data_masked[2641] = data_i[2641] & sel_one_hot_i[20];
  assign data_masked[2640] = data_i[2640] & sel_one_hot_i[20];
  assign data_masked[2639] = data_i[2639] & sel_one_hot_i[20];
  assign data_masked[2638] = data_i[2638] & sel_one_hot_i[20];
  assign data_masked[2637] = data_i[2637] & sel_one_hot_i[20];
  assign data_masked[2636] = data_i[2636] & sel_one_hot_i[20];
  assign data_masked[2635] = data_i[2635] & sel_one_hot_i[20];
  assign data_masked[2634] = data_i[2634] & sel_one_hot_i[20];
  assign data_masked[2633] = data_i[2633] & sel_one_hot_i[20];
  assign data_masked[2632] = data_i[2632] & sel_one_hot_i[20];
  assign data_masked[2631] = data_i[2631] & sel_one_hot_i[20];
  assign data_masked[2630] = data_i[2630] & sel_one_hot_i[20];
  assign data_masked[2629] = data_i[2629] & sel_one_hot_i[20];
  assign data_masked[2628] = data_i[2628] & sel_one_hot_i[20];
  assign data_masked[2627] = data_i[2627] & sel_one_hot_i[20];
  assign data_masked[2626] = data_i[2626] & sel_one_hot_i[20];
  assign data_masked[2625] = data_i[2625] & sel_one_hot_i[20];
  assign data_masked[2624] = data_i[2624] & sel_one_hot_i[20];
  assign data_masked[2623] = data_i[2623] & sel_one_hot_i[20];
  assign data_masked[2622] = data_i[2622] & sel_one_hot_i[20];
  assign data_masked[2621] = data_i[2621] & sel_one_hot_i[20];
  assign data_masked[2620] = data_i[2620] & sel_one_hot_i[20];
  assign data_masked[2619] = data_i[2619] & sel_one_hot_i[20];
  assign data_masked[2618] = data_i[2618] & sel_one_hot_i[20];
  assign data_masked[2617] = data_i[2617] & sel_one_hot_i[20];
  assign data_masked[2616] = data_i[2616] & sel_one_hot_i[20];
  assign data_masked[2615] = data_i[2615] & sel_one_hot_i[20];
  assign data_masked[2614] = data_i[2614] & sel_one_hot_i[20];
  assign data_masked[2613] = data_i[2613] & sel_one_hot_i[20];
  assign data_masked[2612] = data_i[2612] & sel_one_hot_i[20];
  assign data_masked[2611] = data_i[2611] & sel_one_hot_i[20];
  assign data_masked[2610] = data_i[2610] & sel_one_hot_i[20];
  assign data_masked[2609] = data_i[2609] & sel_one_hot_i[20];
  assign data_masked[2608] = data_i[2608] & sel_one_hot_i[20];
  assign data_masked[2607] = data_i[2607] & sel_one_hot_i[20];
  assign data_masked[2606] = data_i[2606] & sel_one_hot_i[20];
  assign data_masked[2605] = data_i[2605] & sel_one_hot_i[20];
  assign data_masked[2604] = data_i[2604] & sel_one_hot_i[20];
  assign data_masked[2603] = data_i[2603] & sel_one_hot_i[20];
  assign data_masked[2602] = data_i[2602] & sel_one_hot_i[20];
  assign data_masked[2601] = data_i[2601] & sel_one_hot_i[20];
  assign data_masked[2600] = data_i[2600] & sel_one_hot_i[20];
  assign data_masked[2599] = data_i[2599] & sel_one_hot_i[20];
  assign data_masked[2598] = data_i[2598] & sel_one_hot_i[20];
  assign data_masked[2597] = data_i[2597] & sel_one_hot_i[20];
  assign data_masked[2596] = data_i[2596] & sel_one_hot_i[20];
  assign data_masked[2595] = data_i[2595] & sel_one_hot_i[20];
  assign data_masked[2594] = data_i[2594] & sel_one_hot_i[20];
  assign data_masked[2593] = data_i[2593] & sel_one_hot_i[20];
  assign data_masked[2592] = data_i[2592] & sel_one_hot_i[20];
  assign data_masked[2591] = data_i[2591] & sel_one_hot_i[20];
  assign data_masked[2590] = data_i[2590] & sel_one_hot_i[20];
  assign data_masked[2589] = data_i[2589] & sel_one_hot_i[20];
  assign data_masked[2588] = data_i[2588] & sel_one_hot_i[20];
  assign data_masked[2587] = data_i[2587] & sel_one_hot_i[20];
  assign data_masked[2586] = data_i[2586] & sel_one_hot_i[20];
  assign data_masked[2585] = data_i[2585] & sel_one_hot_i[20];
  assign data_masked[2584] = data_i[2584] & sel_one_hot_i[20];
  assign data_masked[2583] = data_i[2583] & sel_one_hot_i[20];
  assign data_masked[2582] = data_i[2582] & sel_one_hot_i[20];
  assign data_masked[2581] = data_i[2581] & sel_one_hot_i[20];
  assign data_masked[2580] = data_i[2580] & sel_one_hot_i[20];
  assign data_masked[2579] = data_i[2579] & sel_one_hot_i[20];
  assign data_masked[2578] = data_i[2578] & sel_one_hot_i[20];
  assign data_masked[2577] = data_i[2577] & sel_one_hot_i[20];
  assign data_masked[2576] = data_i[2576] & sel_one_hot_i[20];
  assign data_masked[2575] = data_i[2575] & sel_one_hot_i[20];
  assign data_masked[2574] = data_i[2574] & sel_one_hot_i[20];
  assign data_masked[2573] = data_i[2573] & sel_one_hot_i[20];
  assign data_masked[2572] = data_i[2572] & sel_one_hot_i[20];
  assign data_masked[2571] = data_i[2571] & sel_one_hot_i[20];
  assign data_masked[2570] = data_i[2570] & sel_one_hot_i[20];
  assign data_masked[2569] = data_i[2569] & sel_one_hot_i[20];
  assign data_masked[2568] = data_i[2568] & sel_one_hot_i[20];
  assign data_masked[2567] = data_i[2567] & sel_one_hot_i[20];
  assign data_masked[2566] = data_i[2566] & sel_one_hot_i[20];
  assign data_masked[2565] = data_i[2565] & sel_one_hot_i[20];
  assign data_masked[2564] = data_i[2564] & sel_one_hot_i[20];
  assign data_masked[2563] = data_i[2563] & sel_one_hot_i[20];
  assign data_masked[2562] = data_i[2562] & sel_one_hot_i[20];
  assign data_masked[2561] = data_i[2561] & sel_one_hot_i[20];
  assign data_masked[2560] = data_i[2560] & sel_one_hot_i[20];
  assign data_masked[2815] = data_i[2815] & sel_one_hot_i[21];
  assign data_masked[2814] = data_i[2814] & sel_one_hot_i[21];
  assign data_masked[2813] = data_i[2813] & sel_one_hot_i[21];
  assign data_masked[2812] = data_i[2812] & sel_one_hot_i[21];
  assign data_masked[2811] = data_i[2811] & sel_one_hot_i[21];
  assign data_masked[2810] = data_i[2810] & sel_one_hot_i[21];
  assign data_masked[2809] = data_i[2809] & sel_one_hot_i[21];
  assign data_masked[2808] = data_i[2808] & sel_one_hot_i[21];
  assign data_masked[2807] = data_i[2807] & sel_one_hot_i[21];
  assign data_masked[2806] = data_i[2806] & sel_one_hot_i[21];
  assign data_masked[2805] = data_i[2805] & sel_one_hot_i[21];
  assign data_masked[2804] = data_i[2804] & sel_one_hot_i[21];
  assign data_masked[2803] = data_i[2803] & sel_one_hot_i[21];
  assign data_masked[2802] = data_i[2802] & sel_one_hot_i[21];
  assign data_masked[2801] = data_i[2801] & sel_one_hot_i[21];
  assign data_masked[2800] = data_i[2800] & sel_one_hot_i[21];
  assign data_masked[2799] = data_i[2799] & sel_one_hot_i[21];
  assign data_masked[2798] = data_i[2798] & sel_one_hot_i[21];
  assign data_masked[2797] = data_i[2797] & sel_one_hot_i[21];
  assign data_masked[2796] = data_i[2796] & sel_one_hot_i[21];
  assign data_masked[2795] = data_i[2795] & sel_one_hot_i[21];
  assign data_masked[2794] = data_i[2794] & sel_one_hot_i[21];
  assign data_masked[2793] = data_i[2793] & sel_one_hot_i[21];
  assign data_masked[2792] = data_i[2792] & sel_one_hot_i[21];
  assign data_masked[2791] = data_i[2791] & sel_one_hot_i[21];
  assign data_masked[2790] = data_i[2790] & sel_one_hot_i[21];
  assign data_masked[2789] = data_i[2789] & sel_one_hot_i[21];
  assign data_masked[2788] = data_i[2788] & sel_one_hot_i[21];
  assign data_masked[2787] = data_i[2787] & sel_one_hot_i[21];
  assign data_masked[2786] = data_i[2786] & sel_one_hot_i[21];
  assign data_masked[2785] = data_i[2785] & sel_one_hot_i[21];
  assign data_masked[2784] = data_i[2784] & sel_one_hot_i[21];
  assign data_masked[2783] = data_i[2783] & sel_one_hot_i[21];
  assign data_masked[2782] = data_i[2782] & sel_one_hot_i[21];
  assign data_masked[2781] = data_i[2781] & sel_one_hot_i[21];
  assign data_masked[2780] = data_i[2780] & sel_one_hot_i[21];
  assign data_masked[2779] = data_i[2779] & sel_one_hot_i[21];
  assign data_masked[2778] = data_i[2778] & sel_one_hot_i[21];
  assign data_masked[2777] = data_i[2777] & sel_one_hot_i[21];
  assign data_masked[2776] = data_i[2776] & sel_one_hot_i[21];
  assign data_masked[2775] = data_i[2775] & sel_one_hot_i[21];
  assign data_masked[2774] = data_i[2774] & sel_one_hot_i[21];
  assign data_masked[2773] = data_i[2773] & sel_one_hot_i[21];
  assign data_masked[2772] = data_i[2772] & sel_one_hot_i[21];
  assign data_masked[2771] = data_i[2771] & sel_one_hot_i[21];
  assign data_masked[2770] = data_i[2770] & sel_one_hot_i[21];
  assign data_masked[2769] = data_i[2769] & sel_one_hot_i[21];
  assign data_masked[2768] = data_i[2768] & sel_one_hot_i[21];
  assign data_masked[2767] = data_i[2767] & sel_one_hot_i[21];
  assign data_masked[2766] = data_i[2766] & sel_one_hot_i[21];
  assign data_masked[2765] = data_i[2765] & sel_one_hot_i[21];
  assign data_masked[2764] = data_i[2764] & sel_one_hot_i[21];
  assign data_masked[2763] = data_i[2763] & sel_one_hot_i[21];
  assign data_masked[2762] = data_i[2762] & sel_one_hot_i[21];
  assign data_masked[2761] = data_i[2761] & sel_one_hot_i[21];
  assign data_masked[2760] = data_i[2760] & sel_one_hot_i[21];
  assign data_masked[2759] = data_i[2759] & sel_one_hot_i[21];
  assign data_masked[2758] = data_i[2758] & sel_one_hot_i[21];
  assign data_masked[2757] = data_i[2757] & sel_one_hot_i[21];
  assign data_masked[2756] = data_i[2756] & sel_one_hot_i[21];
  assign data_masked[2755] = data_i[2755] & sel_one_hot_i[21];
  assign data_masked[2754] = data_i[2754] & sel_one_hot_i[21];
  assign data_masked[2753] = data_i[2753] & sel_one_hot_i[21];
  assign data_masked[2752] = data_i[2752] & sel_one_hot_i[21];
  assign data_masked[2751] = data_i[2751] & sel_one_hot_i[21];
  assign data_masked[2750] = data_i[2750] & sel_one_hot_i[21];
  assign data_masked[2749] = data_i[2749] & sel_one_hot_i[21];
  assign data_masked[2748] = data_i[2748] & sel_one_hot_i[21];
  assign data_masked[2747] = data_i[2747] & sel_one_hot_i[21];
  assign data_masked[2746] = data_i[2746] & sel_one_hot_i[21];
  assign data_masked[2745] = data_i[2745] & sel_one_hot_i[21];
  assign data_masked[2744] = data_i[2744] & sel_one_hot_i[21];
  assign data_masked[2743] = data_i[2743] & sel_one_hot_i[21];
  assign data_masked[2742] = data_i[2742] & sel_one_hot_i[21];
  assign data_masked[2741] = data_i[2741] & sel_one_hot_i[21];
  assign data_masked[2740] = data_i[2740] & sel_one_hot_i[21];
  assign data_masked[2739] = data_i[2739] & sel_one_hot_i[21];
  assign data_masked[2738] = data_i[2738] & sel_one_hot_i[21];
  assign data_masked[2737] = data_i[2737] & sel_one_hot_i[21];
  assign data_masked[2736] = data_i[2736] & sel_one_hot_i[21];
  assign data_masked[2735] = data_i[2735] & sel_one_hot_i[21];
  assign data_masked[2734] = data_i[2734] & sel_one_hot_i[21];
  assign data_masked[2733] = data_i[2733] & sel_one_hot_i[21];
  assign data_masked[2732] = data_i[2732] & sel_one_hot_i[21];
  assign data_masked[2731] = data_i[2731] & sel_one_hot_i[21];
  assign data_masked[2730] = data_i[2730] & sel_one_hot_i[21];
  assign data_masked[2729] = data_i[2729] & sel_one_hot_i[21];
  assign data_masked[2728] = data_i[2728] & sel_one_hot_i[21];
  assign data_masked[2727] = data_i[2727] & sel_one_hot_i[21];
  assign data_masked[2726] = data_i[2726] & sel_one_hot_i[21];
  assign data_masked[2725] = data_i[2725] & sel_one_hot_i[21];
  assign data_masked[2724] = data_i[2724] & sel_one_hot_i[21];
  assign data_masked[2723] = data_i[2723] & sel_one_hot_i[21];
  assign data_masked[2722] = data_i[2722] & sel_one_hot_i[21];
  assign data_masked[2721] = data_i[2721] & sel_one_hot_i[21];
  assign data_masked[2720] = data_i[2720] & sel_one_hot_i[21];
  assign data_masked[2719] = data_i[2719] & sel_one_hot_i[21];
  assign data_masked[2718] = data_i[2718] & sel_one_hot_i[21];
  assign data_masked[2717] = data_i[2717] & sel_one_hot_i[21];
  assign data_masked[2716] = data_i[2716] & sel_one_hot_i[21];
  assign data_masked[2715] = data_i[2715] & sel_one_hot_i[21];
  assign data_masked[2714] = data_i[2714] & sel_one_hot_i[21];
  assign data_masked[2713] = data_i[2713] & sel_one_hot_i[21];
  assign data_masked[2712] = data_i[2712] & sel_one_hot_i[21];
  assign data_masked[2711] = data_i[2711] & sel_one_hot_i[21];
  assign data_masked[2710] = data_i[2710] & sel_one_hot_i[21];
  assign data_masked[2709] = data_i[2709] & sel_one_hot_i[21];
  assign data_masked[2708] = data_i[2708] & sel_one_hot_i[21];
  assign data_masked[2707] = data_i[2707] & sel_one_hot_i[21];
  assign data_masked[2706] = data_i[2706] & sel_one_hot_i[21];
  assign data_masked[2705] = data_i[2705] & sel_one_hot_i[21];
  assign data_masked[2704] = data_i[2704] & sel_one_hot_i[21];
  assign data_masked[2703] = data_i[2703] & sel_one_hot_i[21];
  assign data_masked[2702] = data_i[2702] & sel_one_hot_i[21];
  assign data_masked[2701] = data_i[2701] & sel_one_hot_i[21];
  assign data_masked[2700] = data_i[2700] & sel_one_hot_i[21];
  assign data_masked[2699] = data_i[2699] & sel_one_hot_i[21];
  assign data_masked[2698] = data_i[2698] & sel_one_hot_i[21];
  assign data_masked[2697] = data_i[2697] & sel_one_hot_i[21];
  assign data_masked[2696] = data_i[2696] & sel_one_hot_i[21];
  assign data_masked[2695] = data_i[2695] & sel_one_hot_i[21];
  assign data_masked[2694] = data_i[2694] & sel_one_hot_i[21];
  assign data_masked[2693] = data_i[2693] & sel_one_hot_i[21];
  assign data_masked[2692] = data_i[2692] & sel_one_hot_i[21];
  assign data_masked[2691] = data_i[2691] & sel_one_hot_i[21];
  assign data_masked[2690] = data_i[2690] & sel_one_hot_i[21];
  assign data_masked[2689] = data_i[2689] & sel_one_hot_i[21];
  assign data_masked[2688] = data_i[2688] & sel_one_hot_i[21];
  assign data_masked[2943] = data_i[2943] & sel_one_hot_i[22];
  assign data_masked[2942] = data_i[2942] & sel_one_hot_i[22];
  assign data_masked[2941] = data_i[2941] & sel_one_hot_i[22];
  assign data_masked[2940] = data_i[2940] & sel_one_hot_i[22];
  assign data_masked[2939] = data_i[2939] & sel_one_hot_i[22];
  assign data_masked[2938] = data_i[2938] & sel_one_hot_i[22];
  assign data_masked[2937] = data_i[2937] & sel_one_hot_i[22];
  assign data_masked[2936] = data_i[2936] & sel_one_hot_i[22];
  assign data_masked[2935] = data_i[2935] & sel_one_hot_i[22];
  assign data_masked[2934] = data_i[2934] & sel_one_hot_i[22];
  assign data_masked[2933] = data_i[2933] & sel_one_hot_i[22];
  assign data_masked[2932] = data_i[2932] & sel_one_hot_i[22];
  assign data_masked[2931] = data_i[2931] & sel_one_hot_i[22];
  assign data_masked[2930] = data_i[2930] & sel_one_hot_i[22];
  assign data_masked[2929] = data_i[2929] & sel_one_hot_i[22];
  assign data_masked[2928] = data_i[2928] & sel_one_hot_i[22];
  assign data_masked[2927] = data_i[2927] & sel_one_hot_i[22];
  assign data_masked[2926] = data_i[2926] & sel_one_hot_i[22];
  assign data_masked[2925] = data_i[2925] & sel_one_hot_i[22];
  assign data_masked[2924] = data_i[2924] & sel_one_hot_i[22];
  assign data_masked[2923] = data_i[2923] & sel_one_hot_i[22];
  assign data_masked[2922] = data_i[2922] & sel_one_hot_i[22];
  assign data_masked[2921] = data_i[2921] & sel_one_hot_i[22];
  assign data_masked[2920] = data_i[2920] & sel_one_hot_i[22];
  assign data_masked[2919] = data_i[2919] & sel_one_hot_i[22];
  assign data_masked[2918] = data_i[2918] & sel_one_hot_i[22];
  assign data_masked[2917] = data_i[2917] & sel_one_hot_i[22];
  assign data_masked[2916] = data_i[2916] & sel_one_hot_i[22];
  assign data_masked[2915] = data_i[2915] & sel_one_hot_i[22];
  assign data_masked[2914] = data_i[2914] & sel_one_hot_i[22];
  assign data_masked[2913] = data_i[2913] & sel_one_hot_i[22];
  assign data_masked[2912] = data_i[2912] & sel_one_hot_i[22];
  assign data_masked[2911] = data_i[2911] & sel_one_hot_i[22];
  assign data_masked[2910] = data_i[2910] & sel_one_hot_i[22];
  assign data_masked[2909] = data_i[2909] & sel_one_hot_i[22];
  assign data_masked[2908] = data_i[2908] & sel_one_hot_i[22];
  assign data_masked[2907] = data_i[2907] & sel_one_hot_i[22];
  assign data_masked[2906] = data_i[2906] & sel_one_hot_i[22];
  assign data_masked[2905] = data_i[2905] & sel_one_hot_i[22];
  assign data_masked[2904] = data_i[2904] & sel_one_hot_i[22];
  assign data_masked[2903] = data_i[2903] & sel_one_hot_i[22];
  assign data_masked[2902] = data_i[2902] & sel_one_hot_i[22];
  assign data_masked[2901] = data_i[2901] & sel_one_hot_i[22];
  assign data_masked[2900] = data_i[2900] & sel_one_hot_i[22];
  assign data_masked[2899] = data_i[2899] & sel_one_hot_i[22];
  assign data_masked[2898] = data_i[2898] & sel_one_hot_i[22];
  assign data_masked[2897] = data_i[2897] & sel_one_hot_i[22];
  assign data_masked[2896] = data_i[2896] & sel_one_hot_i[22];
  assign data_masked[2895] = data_i[2895] & sel_one_hot_i[22];
  assign data_masked[2894] = data_i[2894] & sel_one_hot_i[22];
  assign data_masked[2893] = data_i[2893] & sel_one_hot_i[22];
  assign data_masked[2892] = data_i[2892] & sel_one_hot_i[22];
  assign data_masked[2891] = data_i[2891] & sel_one_hot_i[22];
  assign data_masked[2890] = data_i[2890] & sel_one_hot_i[22];
  assign data_masked[2889] = data_i[2889] & sel_one_hot_i[22];
  assign data_masked[2888] = data_i[2888] & sel_one_hot_i[22];
  assign data_masked[2887] = data_i[2887] & sel_one_hot_i[22];
  assign data_masked[2886] = data_i[2886] & sel_one_hot_i[22];
  assign data_masked[2885] = data_i[2885] & sel_one_hot_i[22];
  assign data_masked[2884] = data_i[2884] & sel_one_hot_i[22];
  assign data_masked[2883] = data_i[2883] & sel_one_hot_i[22];
  assign data_masked[2882] = data_i[2882] & sel_one_hot_i[22];
  assign data_masked[2881] = data_i[2881] & sel_one_hot_i[22];
  assign data_masked[2880] = data_i[2880] & sel_one_hot_i[22];
  assign data_masked[2879] = data_i[2879] & sel_one_hot_i[22];
  assign data_masked[2878] = data_i[2878] & sel_one_hot_i[22];
  assign data_masked[2877] = data_i[2877] & sel_one_hot_i[22];
  assign data_masked[2876] = data_i[2876] & sel_one_hot_i[22];
  assign data_masked[2875] = data_i[2875] & sel_one_hot_i[22];
  assign data_masked[2874] = data_i[2874] & sel_one_hot_i[22];
  assign data_masked[2873] = data_i[2873] & sel_one_hot_i[22];
  assign data_masked[2872] = data_i[2872] & sel_one_hot_i[22];
  assign data_masked[2871] = data_i[2871] & sel_one_hot_i[22];
  assign data_masked[2870] = data_i[2870] & sel_one_hot_i[22];
  assign data_masked[2869] = data_i[2869] & sel_one_hot_i[22];
  assign data_masked[2868] = data_i[2868] & sel_one_hot_i[22];
  assign data_masked[2867] = data_i[2867] & sel_one_hot_i[22];
  assign data_masked[2866] = data_i[2866] & sel_one_hot_i[22];
  assign data_masked[2865] = data_i[2865] & sel_one_hot_i[22];
  assign data_masked[2864] = data_i[2864] & sel_one_hot_i[22];
  assign data_masked[2863] = data_i[2863] & sel_one_hot_i[22];
  assign data_masked[2862] = data_i[2862] & sel_one_hot_i[22];
  assign data_masked[2861] = data_i[2861] & sel_one_hot_i[22];
  assign data_masked[2860] = data_i[2860] & sel_one_hot_i[22];
  assign data_masked[2859] = data_i[2859] & sel_one_hot_i[22];
  assign data_masked[2858] = data_i[2858] & sel_one_hot_i[22];
  assign data_masked[2857] = data_i[2857] & sel_one_hot_i[22];
  assign data_masked[2856] = data_i[2856] & sel_one_hot_i[22];
  assign data_masked[2855] = data_i[2855] & sel_one_hot_i[22];
  assign data_masked[2854] = data_i[2854] & sel_one_hot_i[22];
  assign data_masked[2853] = data_i[2853] & sel_one_hot_i[22];
  assign data_masked[2852] = data_i[2852] & sel_one_hot_i[22];
  assign data_masked[2851] = data_i[2851] & sel_one_hot_i[22];
  assign data_masked[2850] = data_i[2850] & sel_one_hot_i[22];
  assign data_masked[2849] = data_i[2849] & sel_one_hot_i[22];
  assign data_masked[2848] = data_i[2848] & sel_one_hot_i[22];
  assign data_masked[2847] = data_i[2847] & sel_one_hot_i[22];
  assign data_masked[2846] = data_i[2846] & sel_one_hot_i[22];
  assign data_masked[2845] = data_i[2845] & sel_one_hot_i[22];
  assign data_masked[2844] = data_i[2844] & sel_one_hot_i[22];
  assign data_masked[2843] = data_i[2843] & sel_one_hot_i[22];
  assign data_masked[2842] = data_i[2842] & sel_one_hot_i[22];
  assign data_masked[2841] = data_i[2841] & sel_one_hot_i[22];
  assign data_masked[2840] = data_i[2840] & sel_one_hot_i[22];
  assign data_masked[2839] = data_i[2839] & sel_one_hot_i[22];
  assign data_masked[2838] = data_i[2838] & sel_one_hot_i[22];
  assign data_masked[2837] = data_i[2837] & sel_one_hot_i[22];
  assign data_masked[2836] = data_i[2836] & sel_one_hot_i[22];
  assign data_masked[2835] = data_i[2835] & sel_one_hot_i[22];
  assign data_masked[2834] = data_i[2834] & sel_one_hot_i[22];
  assign data_masked[2833] = data_i[2833] & sel_one_hot_i[22];
  assign data_masked[2832] = data_i[2832] & sel_one_hot_i[22];
  assign data_masked[2831] = data_i[2831] & sel_one_hot_i[22];
  assign data_masked[2830] = data_i[2830] & sel_one_hot_i[22];
  assign data_masked[2829] = data_i[2829] & sel_one_hot_i[22];
  assign data_masked[2828] = data_i[2828] & sel_one_hot_i[22];
  assign data_masked[2827] = data_i[2827] & sel_one_hot_i[22];
  assign data_masked[2826] = data_i[2826] & sel_one_hot_i[22];
  assign data_masked[2825] = data_i[2825] & sel_one_hot_i[22];
  assign data_masked[2824] = data_i[2824] & sel_one_hot_i[22];
  assign data_masked[2823] = data_i[2823] & sel_one_hot_i[22];
  assign data_masked[2822] = data_i[2822] & sel_one_hot_i[22];
  assign data_masked[2821] = data_i[2821] & sel_one_hot_i[22];
  assign data_masked[2820] = data_i[2820] & sel_one_hot_i[22];
  assign data_masked[2819] = data_i[2819] & sel_one_hot_i[22];
  assign data_masked[2818] = data_i[2818] & sel_one_hot_i[22];
  assign data_masked[2817] = data_i[2817] & sel_one_hot_i[22];
  assign data_masked[2816] = data_i[2816] & sel_one_hot_i[22];
  assign data_masked[3071] = data_i[3071] & sel_one_hot_i[23];
  assign data_masked[3070] = data_i[3070] & sel_one_hot_i[23];
  assign data_masked[3069] = data_i[3069] & sel_one_hot_i[23];
  assign data_masked[3068] = data_i[3068] & sel_one_hot_i[23];
  assign data_masked[3067] = data_i[3067] & sel_one_hot_i[23];
  assign data_masked[3066] = data_i[3066] & sel_one_hot_i[23];
  assign data_masked[3065] = data_i[3065] & sel_one_hot_i[23];
  assign data_masked[3064] = data_i[3064] & sel_one_hot_i[23];
  assign data_masked[3063] = data_i[3063] & sel_one_hot_i[23];
  assign data_masked[3062] = data_i[3062] & sel_one_hot_i[23];
  assign data_masked[3061] = data_i[3061] & sel_one_hot_i[23];
  assign data_masked[3060] = data_i[3060] & sel_one_hot_i[23];
  assign data_masked[3059] = data_i[3059] & sel_one_hot_i[23];
  assign data_masked[3058] = data_i[3058] & sel_one_hot_i[23];
  assign data_masked[3057] = data_i[3057] & sel_one_hot_i[23];
  assign data_masked[3056] = data_i[3056] & sel_one_hot_i[23];
  assign data_masked[3055] = data_i[3055] & sel_one_hot_i[23];
  assign data_masked[3054] = data_i[3054] & sel_one_hot_i[23];
  assign data_masked[3053] = data_i[3053] & sel_one_hot_i[23];
  assign data_masked[3052] = data_i[3052] & sel_one_hot_i[23];
  assign data_masked[3051] = data_i[3051] & sel_one_hot_i[23];
  assign data_masked[3050] = data_i[3050] & sel_one_hot_i[23];
  assign data_masked[3049] = data_i[3049] & sel_one_hot_i[23];
  assign data_masked[3048] = data_i[3048] & sel_one_hot_i[23];
  assign data_masked[3047] = data_i[3047] & sel_one_hot_i[23];
  assign data_masked[3046] = data_i[3046] & sel_one_hot_i[23];
  assign data_masked[3045] = data_i[3045] & sel_one_hot_i[23];
  assign data_masked[3044] = data_i[3044] & sel_one_hot_i[23];
  assign data_masked[3043] = data_i[3043] & sel_one_hot_i[23];
  assign data_masked[3042] = data_i[3042] & sel_one_hot_i[23];
  assign data_masked[3041] = data_i[3041] & sel_one_hot_i[23];
  assign data_masked[3040] = data_i[3040] & sel_one_hot_i[23];
  assign data_masked[3039] = data_i[3039] & sel_one_hot_i[23];
  assign data_masked[3038] = data_i[3038] & sel_one_hot_i[23];
  assign data_masked[3037] = data_i[3037] & sel_one_hot_i[23];
  assign data_masked[3036] = data_i[3036] & sel_one_hot_i[23];
  assign data_masked[3035] = data_i[3035] & sel_one_hot_i[23];
  assign data_masked[3034] = data_i[3034] & sel_one_hot_i[23];
  assign data_masked[3033] = data_i[3033] & sel_one_hot_i[23];
  assign data_masked[3032] = data_i[3032] & sel_one_hot_i[23];
  assign data_masked[3031] = data_i[3031] & sel_one_hot_i[23];
  assign data_masked[3030] = data_i[3030] & sel_one_hot_i[23];
  assign data_masked[3029] = data_i[3029] & sel_one_hot_i[23];
  assign data_masked[3028] = data_i[3028] & sel_one_hot_i[23];
  assign data_masked[3027] = data_i[3027] & sel_one_hot_i[23];
  assign data_masked[3026] = data_i[3026] & sel_one_hot_i[23];
  assign data_masked[3025] = data_i[3025] & sel_one_hot_i[23];
  assign data_masked[3024] = data_i[3024] & sel_one_hot_i[23];
  assign data_masked[3023] = data_i[3023] & sel_one_hot_i[23];
  assign data_masked[3022] = data_i[3022] & sel_one_hot_i[23];
  assign data_masked[3021] = data_i[3021] & sel_one_hot_i[23];
  assign data_masked[3020] = data_i[3020] & sel_one_hot_i[23];
  assign data_masked[3019] = data_i[3019] & sel_one_hot_i[23];
  assign data_masked[3018] = data_i[3018] & sel_one_hot_i[23];
  assign data_masked[3017] = data_i[3017] & sel_one_hot_i[23];
  assign data_masked[3016] = data_i[3016] & sel_one_hot_i[23];
  assign data_masked[3015] = data_i[3015] & sel_one_hot_i[23];
  assign data_masked[3014] = data_i[3014] & sel_one_hot_i[23];
  assign data_masked[3013] = data_i[3013] & sel_one_hot_i[23];
  assign data_masked[3012] = data_i[3012] & sel_one_hot_i[23];
  assign data_masked[3011] = data_i[3011] & sel_one_hot_i[23];
  assign data_masked[3010] = data_i[3010] & sel_one_hot_i[23];
  assign data_masked[3009] = data_i[3009] & sel_one_hot_i[23];
  assign data_masked[3008] = data_i[3008] & sel_one_hot_i[23];
  assign data_masked[3007] = data_i[3007] & sel_one_hot_i[23];
  assign data_masked[3006] = data_i[3006] & sel_one_hot_i[23];
  assign data_masked[3005] = data_i[3005] & sel_one_hot_i[23];
  assign data_masked[3004] = data_i[3004] & sel_one_hot_i[23];
  assign data_masked[3003] = data_i[3003] & sel_one_hot_i[23];
  assign data_masked[3002] = data_i[3002] & sel_one_hot_i[23];
  assign data_masked[3001] = data_i[3001] & sel_one_hot_i[23];
  assign data_masked[3000] = data_i[3000] & sel_one_hot_i[23];
  assign data_masked[2999] = data_i[2999] & sel_one_hot_i[23];
  assign data_masked[2998] = data_i[2998] & sel_one_hot_i[23];
  assign data_masked[2997] = data_i[2997] & sel_one_hot_i[23];
  assign data_masked[2996] = data_i[2996] & sel_one_hot_i[23];
  assign data_masked[2995] = data_i[2995] & sel_one_hot_i[23];
  assign data_masked[2994] = data_i[2994] & sel_one_hot_i[23];
  assign data_masked[2993] = data_i[2993] & sel_one_hot_i[23];
  assign data_masked[2992] = data_i[2992] & sel_one_hot_i[23];
  assign data_masked[2991] = data_i[2991] & sel_one_hot_i[23];
  assign data_masked[2990] = data_i[2990] & sel_one_hot_i[23];
  assign data_masked[2989] = data_i[2989] & sel_one_hot_i[23];
  assign data_masked[2988] = data_i[2988] & sel_one_hot_i[23];
  assign data_masked[2987] = data_i[2987] & sel_one_hot_i[23];
  assign data_masked[2986] = data_i[2986] & sel_one_hot_i[23];
  assign data_masked[2985] = data_i[2985] & sel_one_hot_i[23];
  assign data_masked[2984] = data_i[2984] & sel_one_hot_i[23];
  assign data_masked[2983] = data_i[2983] & sel_one_hot_i[23];
  assign data_masked[2982] = data_i[2982] & sel_one_hot_i[23];
  assign data_masked[2981] = data_i[2981] & sel_one_hot_i[23];
  assign data_masked[2980] = data_i[2980] & sel_one_hot_i[23];
  assign data_masked[2979] = data_i[2979] & sel_one_hot_i[23];
  assign data_masked[2978] = data_i[2978] & sel_one_hot_i[23];
  assign data_masked[2977] = data_i[2977] & sel_one_hot_i[23];
  assign data_masked[2976] = data_i[2976] & sel_one_hot_i[23];
  assign data_masked[2975] = data_i[2975] & sel_one_hot_i[23];
  assign data_masked[2974] = data_i[2974] & sel_one_hot_i[23];
  assign data_masked[2973] = data_i[2973] & sel_one_hot_i[23];
  assign data_masked[2972] = data_i[2972] & sel_one_hot_i[23];
  assign data_masked[2971] = data_i[2971] & sel_one_hot_i[23];
  assign data_masked[2970] = data_i[2970] & sel_one_hot_i[23];
  assign data_masked[2969] = data_i[2969] & sel_one_hot_i[23];
  assign data_masked[2968] = data_i[2968] & sel_one_hot_i[23];
  assign data_masked[2967] = data_i[2967] & sel_one_hot_i[23];
  assign data_masked[2966] = data_i[2966] & sel_one_hot_i[23];
  assign data_masked[2965] = data_i[2965] & sel_one_hot_i[23];
  assign data_masked[2964] = data_i[2964] & sel_one_hot_i[23];
  assign data_masked[2963] = data_i[2963] & sel_one_hot_i[23];
  assign data_masked[2962] = data_i[2962] & sel_one_hot_i[23];
  assign data_masked[2961] = data_i[2961] & sel_one_hot_i[23];
  assign data_masked[2960] = data_i[2960] & sel_one_hot_i[23];
  assign data_masked[2959] = data_i[2959] & sel_one_hot_i[23];
  assign data_masked[2958] = data_i[2958] & sel_one_hot_i[23];
  assign data_masked[2957] = data_i[2957] & sel_one_hot_i[23];
  assign data_masked[2956] = data_i[2956] & sel_one_hot_i[23];
  assign data_masked[2955] = data_i[2955] & sel_one_hot_i[23];
  assign data_masked[2954] = data_i[2954] & sel_one_hot_i[23];
  assign data_masked[2953] = data_i[2953] & sel_one_hot_i[23];
  assign data_masked[2952] = data_i[2952] & sel_one_hot_i[23];
  assign data_masked[2951] = data_i[2951] & sel_one_hot_i[23];
  assign data_masked[2950] = data_i[2950] & sel_one_hot_i[23];
  assign data_masked[2949] = data_i[2949] & sel_one_hot_i[23];
  assign data_masked[2948] = data_i[2948] & sel_one_hot_i[23];
  assign data_masked[2947] = data_i[2947] & sel_one_hot_i[23];
  assign data_masked[2946] = data_i[2946] & sel_one_hot_i[23];
  assign data_masked[2945] = data_i[2945] & sel_one_hot_i[23];
  assign data_masked[2944] = data_i[2944] & sel_one_hot_i[23];
  assign data_masked[3199] = data_i[3199] & sel_one_hot_i[24];
  assign data_masked[3198] = data_i[3198] & sel_one_hot_i[24];
  assign data_masked[3197] = data_i[3197] & sel_one_hot_i[24];
  assign data_masked[3196] = data_i[3196] & sel_one_hot_i[24];
  assign data_masked[3195] = data_i[3195] & sel_one_hot_i[24];
  assign data_masked[3194] = data_i[3194] & sel_one_hot_i[24];
  assign data_masked[3193] = data_i[3193] & sel_one_hot_i[24];
  assign data_masked[3192] = data_i[3192] & sel_one_hot_i[24];
  assign data_masked[3191] = data_i[3191] & sel_one_hot_i[24];
  assign data_masked[3190] = data_i[3190] & sel_one_hot_i[24];
  assign data_masked[3189] = data_i[3189] & sel_one_hot_i[24];
  assign data_masked[3188] = data_i[3188] & sel_one_hot_i[24];
  assign data_masked[3187] = data_i[3187] & sel_one_hot_i[24];
  assign data_masked[3186] = data_i[3186] & sel_one_hot_i[24];
  assign data_masked[3185] = data_i[3185] & sel_one_hot_i[24];
  assign data_masked[3184] = data_i[3184] & sel_one_hot_i[24];
  assign data_masked[3183] = data_i[3183] & sel_one_hot_i[24];
  assign data_masked[3182] = data_i[3182] & sel_one_hot_i[24];
  assign data_masked[3181] = data_i[3181] & sel_one_hot_i[24];
  assign data_masked[3180] = data_i[3180] & sel_one_hot_i[24];
  assign data_masked[3179] = data_i[3179] & sel_one_hot_i[24];
  assign data_masked[3178] = data_i[3178] & sel_one_hot_i[24];
  assign data_masked[3177] = data_i[3177] & sel_one_hot_i[24];
  assign data_masked[3176] = data_i[3176] & sel_one_hot_i[24];
  assign data_masked[3175] = data_i[3175] & sel_one_hot_i[24];
  assign data_masked[3174] = data_i[3174] & sel_one_hot_i[24];
  assign data_masked[3173] = data_i[3173] & sel_one_hot_i[24];
  assign data_masked[3172] = data_i[3172] & sel_one_hot_i[24];
  assign data_masked[3171] = data_i[3171] & sel_one_hot_i[24];
  assign data_masked[3170] = data_i[3170] & sel_one_hot_i[24];
  assign data_masked[3169] = data_i[3169] & sel_one_hot_i[24];
  assign data_masked[3168] = data_i[3168] & sel_one_hot_i[24];
  assign data_masked[3167] = data_i[3167] & sel_one_hot_i[24];
  assign data_masked[3166] = data_i[3166] & sel_one_hot_i[24];
  assign data_masked[3165] = data_i[3165] & sel_one_hot_i[24];
  assign data_masked[3164] = data_i[3164] & sel_one_hot_i[24];
  assign data_masked[3163] = data_i[3163] & sel_one_hot_i[24];
  assign data_masked[3162] = data_i[3162] & sel_one_hot_i[24];
  assign data_masked[3161] = data_i[3161] & sel_one_hot_i[24];
  assign data_masked[3160] = data_i[3160] & sel_one_hot_i[24];
  assign data_masked[3159] = data_i[3159] & sel_one_hot_i[24];
  assign data_masked[3158] = data_i[3158] & sel_one_hot_i[24];
  assign data_masked[3157] = data_i[3157] & sel_one_hot_i[24];
  assign data_masked[3156] = data_i[3156] & sel_one_hot_i[24];
  assign data_masked[3155] = data_i[3155] & sel_one_hot_i[24];
  assign data_masked[3154] = data_i[3154] & sel_one_hot_i[24];
  assign data_masked[3153] = data_i[3153] & sel_one_hot_i[24];
  assign data_masked[3152] = data_i[3152] & sel_one_hot_i[24];
  assign data_masked[3151] = data_i[3151] & sel_one_hot_i[24];
  assign data_masked[3150] = data_i[3150] & sel_one_hot_i[24];
  assign data_masked[3149] = data_i[3149] & sel_one_hot_i[24];
  assign data_masked[3148] = data_i[3148] & sel_one_hot_i[24];
  assign data_masked[3147] = data_i[3147] & sel_one_hot_i[24];
  assign data_masked[3146] = data_i[3146] & sel_one_hot_i[24];
  assign data_masked[3145] = data_i[3145] & sel_one_hot_i[24];
  assign data_masked[3144] = data_i[3144] & sel_one_hot_i[24];
  assign data_masked[3143] = data_i[3143] & sel_one_hot_i[24];
  assign data_masked[3142] = data_i[3142] & sel_one_hot_i[24];
  assign data_masked[3141] = data_i[3141] & sel_one_hot_i[24];
  assign data_masked[3140] = data_i[3140] & sel_one_hot_i[24];
  assign data_masked[3139] = data_i[3139] & sel_one_hot_i[24];
  assign data_masked[3138] = data_i[3138] & sel_one_hot_i[24];
  assign data_masked[3137] = data_i[3137] & sel_one_hot_i[24];
  assign data_masked[3136] = data_i[3136] & sel_one_hot_i[24];
  assign data_masked[3135] = data_i[3135] & sel_one_hot_i[24];
  assign data_masked[3134] = data_i[3134] & sel_one_hot_i[24];
  assign data_masked[3133] = data_i[3133] & sel_one_hot_i[24];
  assign data_masked[3132] = data_i[3132] & sel_one_hot_i[24];
  assign data_masked[3131] = data_i[3131] & sel_one_hot_i[24];
  assign data_masked[3130] = data_i[3130] & sel_one_hot_i[24];
  assign data_masked[3129] = data_i[3129] & sel_one_hot_i[24];
  assign data_masked[3128] = data_i[3128] & sel_one_hot_i[24];
  assign data_masked[3127] = data_i[3127] & sel_one_hot_i[24];
  assign data_masked[3126] = data_i[3126] & sel_one_hot_i[24];
  assign data_masked[3125] = data_i[3125] & sel_one_hot_i[24];
  assign data_masked[3124] = data_i[3124] & sel_one_hot_i[24];
  assign data_masked[3123] = data_i[3123] & sel_one_hot_i[24];
  assign data_masked[3122] = data_i[3122] & sel_one_hot_i[24];
  assign data_masked[3121] = data_i[3121] & sel_one_hot_i[24];
  assign data_masked[3120] = data_i[3120] & sel_one_hot_i[24];
  assign data_masked[3119] = data_i[3119] & sel_one_hot_i[24];
  assign data_masked[3118] = data_i[3118] & sel_one_hot_i[24];
  assign data_masked[3117] = data_i[3117] & sel_one_hot_i[24];
  assign data_masked[3116] = data_i[3116] & sel_one_hot_i[24];
  assign data_masked[3115] = data_i[3115] & sel_one_hot_i[24];
  assign data_masked[3114] = data_i[3114] & sel_one_hot_i[24];
  assign data_masked[3113] = data_i[3113] & sel_one_hot_i[24];
  assign data_masked[3112] = data_i[3112] & sel_one_hot_i[24];
  assign data_masked[3111] = data_i[3111] & sel_one_hot_i[24];
  assign data_masked[3110] = data_i[3110] & sel_one_hot_i[24];
  assign data_masked[3109] = data_i[3109] & sel_one_hot_i[24];
  assign data_masked[3108] = data_i[3108] & sel_one_hot_i[24];
  assign data_masked[3107] = data_i[3107] & sel_one_hot_i[24];
  assign data_masked[3106] = data_i[3106] & sel_one_hot_i[24];
  assign data_masked[3105] = data_i[3105] & sel_one_hot_i[24];
  assign data_masked[3104] = data_i[3104] & sel_one_hot_i[24];
  assign data_masked[3103] = data_i[3103] & sel_one_hot_i[24];
  assign data_masked[3102] = data_i[3102] & sel_one_hot_i[24];
  assign data_masked[3101] = data_i[3101] & sel_one_hot_i[24];
  assign data_masked[3100] = data_i[3100] & sel_one_hot_i[24];
  assign data_masked[3099] = data_i[3099] & sel_one_hot_i[24];
  assign data_masked[3098] = data_i[3098] & sel_one_hot_i[24];
  assign data_masked[3097] = data_i[3097] & sel_one_hot_i[24];
  assign data_masked[3096] = data_i[3096] & sel_one_hot_i[24];
  assign data_masked[3095] = data_i[3095] & sel_one_hot_i[24];
  assign data_masked[3094] = data_i[3094] & sel_one_hot_i[24];
  assign data_masked[3093] = data_i[3093] & sel_one_hot_i[24];
  assign data_masked[3092] = data_i[3092] & sel_one_hot_i[24];
  assign data_masked[3091] = data_i[3091] & sel_one_hot_i[24];
  assign data_masked[3090] = data_i[3090] & sel_one_hot_i[24];
  assign data_masked[3089] = data_i[3089] & sel_one_hot_i[24];
  assign data_masked[3088] = data_i[3088] & sel_one_hot_i[24];
  assign data_masked[3087] = data_i[3087] & sel_one_hot_i[24];
  assign data_masked[3086] = data_i[3086] & sel_one_hot_i[24];
  assign data_masked[3085] = data_i[3085] & sel_one_hot_i[24];
  assign data_masked[3084] = data_i[3084] & sel_one_hot_i[24];
  assign data_masked[3083] = data_i[3083] & sel_one_hot_i[24];
  assign data_masked[3082] = data_i[3082] & sel_one_hot_i[24];
  assign data_masked[3081] = data_i[3081] & sel_one_hot_i[24];
  assign data_masked[3080] = data_i[3080] & sel_one_hot_i[24];
  assign data_masked[3079] = data_i[3079] & sel_one_hot_i[24];
  assign data_masked[3078] = data_i[3078] & sel_one_hot_i[24];
  assign data_masked[3077] = data_i[3077] & sel_one_hot_i[24];
  assign data_masked[3076] = data_i[3076] & sel_one_hot_i[24];
  assign data_masked[3075] = data_i[3075] & sel_one_hot_i[24];
  assign data_masked[3074] = data_i[3074] & sel_one_hot_i[24];
  assign data_masked[3073] = data_i[3073] & sel_one_hot_i[24];
  assign data_masked[3072] = data_i[3072] & sel_one_hot_i[24];
  assign data_masked[3327] = data_i[3327] & sel_one_hot_i[25];
  assign data_masked[3326] = data_i[3326] & sel_one_hot_i[25];
  assign data_masked[3325] = data_i[3325] & sel_one_hot_i[25];
  assign data_masked[3324] = data_i[3324] & sel_one_hot_i[25];
  assign data_masked[3323] = data_i[3323] & sel_one_hot_i[25];
  assign data_masked[3322] = data_i[3322] & sel_one_hot_i[25];
  assign data_masked[3321] = data_i[3321] & sel_one_hot_i[25];
  assign data_masked[3320] = data_i[3320] & sel_one_hot_i[25];
  assign data_masked[3319] = data_i[3319] & sel_one_hot_i[25];
  assign data_masked[3318] = data_i[3318] & sel_one_hot_i[25];
  assign data_masked[3317] = data_i[3317] & sel_one_hot_i[25];
  assign data_masked[3316] = data_i[3316] & sel_one_hot_i[25];
  assign data_masked[3315] = data_i[3315] & sel_one_hot_i[25];
  assign data_masked[3314] = data_i[3314] & sel_one_hot_i[25];
  assign data_masked[3313] = data_i[3313] & sel_one_hot_i[25];
  assign data_masked[3312] = data_i[3312] & sel_one_hot_i[25];
  assign data_masked[3311] = data_i[3311] & sel_one_hot_i[25];
  assign data_masked[3310] = data_i[3310] & sel_one_hot_i[25];
  assign data_masked[3309] = data_i[3309] & sel_one_hot_i[25];
  assign data_masked[3308] = data_i[3308] & sel_one_hot_i[25];
  assign data_masked[3307] = data_i[3307] & sel_one_hot_i[25];
  assign data_masked[3306] = data_i[3306] & sel_one_hot_i[25];
  assign data_masked[3305] = data_i[3305] & sel_one_hot_i[25];
  assign data_masked[3304] = data_i[3304] & sel_one_hot_i[25];
  assign data_masked[3303] = data_i[3303] & sel_one_hot_i[25];
  assign data_masked[3302] = data_i[3302] & sel_one_hot_i[25];
  assign data_masked[3301] = data_i[3301] & sel_one_hot_i[25];
  assign data_masked[3300] = data_i[3300] & sel_one_hot_i[25];
  assign data_masked[3299] = data_i[3299] & sel_one_hot_i[25];
  assign data_masked[3298] = data_i[3298] & sel_one_hot_i[25];
  assign data_masked[3297] = data_i[3297] & sel_one_hot_i[25];
  assign data_masked[3296] = data_i[3296] & sel_one_hot_i[25];
  assign data_masked[3295] = data_i[3295] & sel_one_hot_i[25];
  assign data_masked[3294] = data_i[3294] & sel_one_hot_i[25];
  assign data_masked[3293] = data_i[3293] & sel_one_hot_i[25];
  assign data_masked[3292] = data_i[3292] & sel_one_hot_i[25];
  assign data_masked[3291] = data_i[3291] & sel_one_hot_i[25];
  assign data_masked[3290] = data_i[3290] & sel_one_hot_i[25];
  assign data_masked[3289] = data_i[3289] & sel_one_hot_i[25];
  assign data_masked[3288] = data_i[3288] & sel_one_hot_i[25];
  assign data_masked[3287] = data_i[3287] & sel_one_hot_i[25];
  assign data_masked[3286] = data_i[3286] & sel_one_hot_i[25];
  assign data_masked[3285] = data_i[3285] & sel_one_hot_i[25];
  assign data_masked[3284] = data_i[3284] & sel_one_hot_i[25];
  assign data_masked[3283] = data_i[3283] & sel_one_hot_i[25];
  assign data_masked[3282] = data_i[3282] & sel_one_hot_i[25];
  assign data_masked[3281] = data_i[3281] & sel_one_hot_i[25];
  assign data_masked[3280] = data_i[3280] & sel_one_hot_i[25];
  assign data_masked[3279] = data_i[3279] & sel_one_hot_i[25];
  assign data_masked[3278] = data_i[3278] & sel_one_hot_i[25];
  assign data_masked[3277] = data_i[3277] & sel_one_hot_i[25];
  assign data_masked[3276] = data_i[3276] & sel_one_hot_i[25];
  assign data_masked[3275] = data_i[3275] & sel_one_hot_i[25];
  assign data_masked[3274] = data_i[3274] & sel_one_hot_i[25];
  assign data_masked[3273] = data_i[3273] & sel_one_hot_i[25];
  assign data_masked[3272] = data_i[3272] & sel_one_hot_i[25];
  assign data_masked[3271] = data_i[3271] & sel_one_hot_i[25];
  assign data_masked[3270] = data_i[3270] & sel_one_hot_i[25];
  assign data_masked[3269] = data_i[3269] & sel_one_hot_i[25];
  assign data_masked[3268] = data_i[3268] & sel_one_hot_i[25];
  assign data_masked[3267] = data_i[3267] & sel_one_hot_i[25];
  assign data_masked[3266] = data_i[3266] & sel_one_hot_i[25];
  assign data_masked[3265] = data_i[3265] & sel_one_hot_i[25];
  assign data_masked[3264] = data_i[3264] & sel_one_hot_i[25];
  assign data_masked[3263] = data_i[3263] & sel_one_hot_i[25];
  assign data_masked[3262] = data_i[3262] & sel_one_hot_i[25];
  assign data_masked[3261] = data_i[3261] & sel_one_hot_i[25];
  assign data_masked[3260] = data_i[3260] & sel_one_hot_i[25];
  assign data_masked[3259] = data_i[3259] & sel_one_hot_i[25];
  assign data_masked[3258] = data_i[3258] & sel_one_hot_i[25];
  assign data_masked[3257] = data_i[3257] & sel_one_hot_i[25];
  assign data_masked[3256] = data_i[3256] & sel_one_hot_i[25];
  assign data_masked[3255] = data_i[3255] & sel_one_hot_i[25];
  assign data_masked[3254] = data_i[3254] & sel_one_hot_i[25];
  assign data_masked[3253] = data_i[3253] & sel_one_hot_i[25];
  assign data_masked[3252] = data_i[3252] & sel_one_hot_i[25];
  assign data_masked[3251] = data_i[3251] & sel_one_hot_i[25];
  assign data_masked[3250] = data_i[3250] & sel_one_hot_i[25];
  assign data_masked[3249] = data_i[3249] & sel_one_hot_i[25];
  assign data_masked[3248] = data_i[3248] & sel_one_hot_i[25];
  assign data_masked[3247] = data_i[3247] & sel_one_hot_i[25];
  assign data_masked[3246] = data_i[3246] & sel_one_hot_i[25];
  assign data_masked[3245] = data_i[3245] & sel_one_hot_i[25];
  assign data_masked[3244] = data_i[3244] & sel_one_hot_i[25];
  assign data_masked[3243] = data_i[3243] & sel_one_hot_i[25];
  assign data_masked[3242] = data_i[3242] & sel_one_hot_i[25];
  assign data_masked[3241] = data_i[3241] & sel_one_hot_i[25];
  assign data_masked[3240] = data_i[3240] & sel_one_hot_i[25];
  assign data_masked[3239] = data_i[3239] & sel_one_hot_i[25];
  assign data_masked[3238] = data_i[3238] & sel_one_hot_i[25];
  assign data_masked[3237] = data_i[3237] & sel_one_hot_i[25];
  assign data_masked[3236] = data_i[3236] & sel_one_hot_i[25];
  assign data_masked[3235] = data_i[3235] & sel_one_hot_i[25];
  assign data_masked[3234] = data_i[3234] & sel_one_hot_i[25];
  assign data_masked[3233] = data_i[3233] & sel_one_hot_i[25];
  assign data_masked[3232] = data_i[3232] & sel_one_hot_i[25];
  assign data_masked[3231] = data_i[3231] & sel_one_hot_i[25];
  assign data_masked[3230] = data_i[3230] & sel_one_hot_i[25];
  assign data_masked[3229] = data_i[3229] & sel_one_hot_i[25];
  assign data_masked[3228] = data_i[3228] & sel_one_hot_i[25];
  assign data_masked[3227] = data_i[3227] & sel_one_hot_i[25];
  assign data_masked[3226] = data_i[3226] & sel_one_hot_i[25];
  assign data_masked[3225] = data_i[3225] & sel_one_hot_i[25];
  assign data_masked[3224] = data_i[3224] & sel_one_hot_i[25];
  assign data_masked[3223] = data_i[3223] & sel_one_hot_i[25];
  assign data_masked[3222] = data_i[3222] & sel_one_hot_i[25];
  assign data_masked[3221] = data_i[3221] & sel_one_hot_i[25];
  assign data_masked[3220] = data_i[3220] & sel_one_hot_i[25];
  assign data_masked[3219] = data_i[3219] & sel_one_hot_i[25];
  assign data_masked[3218] = data_i[3218] & sel_one_hot_i[25];
  assign data_masked[3217] = data_i[3217] & sel_one_hot_i[25];
  assign data_masked[3216] = data_i[3216] & sel_one_hot_i[25];
  assign data_masked[3215] = data_i[3215] & sel_one_hot_i[25];
  assign data_masked[3214] = data_i[3214] & sel_one_hot_i[25];
  assign data_masked[3213] = data_i[3213] & sel_one_hot_i[25];
  assign data_masked[3212] = data_i[3212] & sel_one_hot_i[25];
  assign data_masked[3211] = data_i[3211] & sel_one_hot_i[25];
  assign data_masked[3210] = data_i[3210] & sel_one_hot_i[25];
  assign data_masked[3209] = data_i[3209] & sel_one_hot_i[25];
  assign data_masked[3208] = data_i[3208] & sel_one_hot_i[25];
  assign data_masked[3207] = data_i[3207] & sel_one_hot_i[25];
  assign data_masked[3206] = data_i[3206] & sel_one_hot_i[25];
  assign data_masked[3205] = data_i[3205] & sel_one_hot_i[25];
  assign data_masked[3204] = data_i[3204] & sel_one_hot_i[25];
  assign data_masked[3203] = data_i[3203] & sel_one_hot_i[25];
  assign data_masked[3202] = data_i[3202] & sel_one_hot_i[25];
  assign data_masked[3201] = data_i[3201] & sel_one_hot_i[25];
  assign data_masked[3200] = data_i[3200] & sel_one_hot_i[25];
  assign data_masked[3455] = data_i[3455] & sel_one_hot_i[26];
  assign data_masked[3454] = data_i[3454] & sel_one_hot_i[26];
  assign data_masked[3453] = data_i[3453] & sel_one_hot_i[26];
  assign data_masked[3452] = data_i[3452] & sel_one_hot_i[26];
  assign data_masked[3451] = data_i[3451] & sel_one_hot_i[26];
  assign data_masked[3450] = data_i[3450] & sel_one_hot_i[26];
  assign data_masked[3449] = data_i[3449] & sel_one_hot_i[26];
  assign data_masked[3448] = data_i[3448] & sel_one_hot_i[26];
  assign data_masked[3447] = data_i[3447] & sel_one_hot_i[26];
  assign data_masked[3446] = data_i[3446] & sel_one_hot_i[26];
  assign data_masked[3445] = data_i[3445] & sel_one_hot_i[26];
  assign data_masked[3444] = data_i[3444] & sel_one_hot_i[26];
  assign data_masked[3443] = data_i[3443] & sel_one_hot_i[26];
  assign data_masked[3442] = data_i[3442] & sel_one_hot_i[26];
  assign data_masked[3441] = data_i[3441] & sel_one_hot_i[26];
  assign data_masked[3440] = data_i[3440] & sel_one_hot_i[26];
  assign data_masked[3439] = data_i[3439] & sel_one_hot_i[26];
  assign data_masked[3438] = data_i[3438] & sel_one_hot_i[26];
  assign data_masked[3437] = data_i[3437] & sel_one_hot_i[26];
  assign data_masked[3436] = data_i[3436] & sel_one_hot_i[26];
  assign data_masked[3435] = data_i[3435] & sel_one_hot_i[26];
  assign data_masked[3434] = data_i[3434] & sel_one_hot_i[26];
  assign data_masked[3433] = data_i[3433] & sel_one_hot_i[26];
  assign data_masked[3432] = data_i[3432] & sel_one_hot_i[26];
  assign data_masked[3431] = data_i[3431] & sel_one_hot_i[26];
  assign data_masked[3430] = data_i[3430] & sel_one_hot_i[26];
  assign data_masked[3429] = data_i[3429] & sel_one_hot_i[26];
  assign data_masked[3428] = data_i[3428] & sel_one_hot_i[26];
  assign data_masked[3427] = data_i[3427] & sel_one_hot_i[26];
  assign data_masked[3426] = data_i[3426] & sel_one_hot_i[26];
  assign data_masked[3425] = data_i[3425] & sel_one_hot_i[26];
  assign data_masked[3424] = data_i[3424] & sel_one_hot_i[26];
  assign data_masked[3423] = data_i[3423] & sel_one_hot_i[26];
  assign data_masked[3422] = data_i[3422] & sel_one_hot_i[26];
  assign data_masked[3421] = data_i[3421] & sel_one_hot_i[26];
  assign data_masked[3420] = data_i[3420] & sel_one_hot_i[26];
  assign data_masked[3419] = data_i[3419] & sel_one_hot_i[26];
  assign data_masked[3418] = data_i[3418] & sel_one_hot_i[26];
  assign data_masked[3417] = data_i[3417] & sel_one_hot_i[26];
  assign data_masked[3416] = data_i[3416] & sel_one_hot_i[26];
  assign data_masked[3415] = data_i[3415] & sel_one_hot_i[26];
  assign data_masked[3414] = data_i[3414] & sel_one_hot_i[26];
  assign data_masked[3413] = data_i[3413] & sel_one_hot_i[26];
  assign data_masked[3412] = data_i[3412] & sel_one_hot_i[26];
  assign data_masked[3411] = data_i[3411] & sel_one_hot_i[26];
  assign data_masked[3410] = data_i[3410] & sel_one_hot_i[26];
  assign data_masked[3409] = data_i[3409] & sel_one_hot_i[26];
  assign data_masked[3408] = data_i[3408] & sel_one_hot_i[26];
  assign data_masked[3407] = data_i[3407] & sel_one_hot_i[26];
  assign data_masked[3406] = data_i[3406] & sel_one_hot_i[26];
  assign data_masked[3405] = data_i[3405] & sel_one_hot_i[26];
  assign data_masked[3404] = data_i[3404] & sel_one_hot_i[26];
  assign data_masked[3403] = data_i[3403] & sel_one_hot_i[26];
  assign data_masked[3402] = data_i[3402] & sel_one_hot_i[26];
  assign data_masked[3401] = data_i[3401] & sel_one_hot_i[26];
  assign data_masked[3400] = data_i[3400] & sel_one_hot_i[26];
  assign data_masked[3399] = data_i[3399] & sel_one_hot_i[26];
  assign data_masked[3398] = data_i[3398] & sel_one_hot_i[26];
  assign data_masked[3397] = data_i[3397] & sel_one_hot_i[26];
  assign data_masked[3396] = data_i[3396] & sel_one_hot_i[26];
  assign data_masked[3395] = data_i[3395] & sel_one_hot_i[26];
  assign data_masked[3394] = data_i[3394] & sel_one_hot_i[26];
  assign data_masked[3393] = data_i[3393] & sel_one_hot_i[26];
  assign data_masked[3392] = data_i[3392] & sel_one_hot_i[26];
  assign data_masked[3391] = data_i[3391] & sel_one_hot_i[26];
  assign data_masked[3390] = data_i[3390] & sel_one_hot_i[26];
  assign data_masked[3389] = data_i[3389] & sel_one_hot_i[26];
  assign data_masked[3388] = data_i[3388] & sel_one_hot_i[26];
  assign data_masked[3387] = data_i[3387] & sel_one_hot_i[26];
  assign data_masked[3386] = data_i[3386] & sel_one_hot_i[26];
  assign data_masked[3385] = data_i[3385] & sel_one_hot_i[26];
  assign data_masked[3384] = data_i[3384] & sel_one_hot_i[26];
  assign data_masked[3383] = data_i[3383] & sel_one_hot_i[26];
  assign data_masked[3382] = data_i[3382] & sel_one_hot_i[26];
  assign data_masked[3381] = data_i[3381] & sel_one_hot_i[26];
  assign data_masked[3380] = data_i[3380] & sel_one_hot_i[26];
  assign data_masked[3379] = data_i[3379] & sel_one_hot_i[26];
  assign data_masked[3378] = data_i[3378] & sel_one_hot_i[26];
  assign data_masked[3377] = data_i[3377] & sel_one_hot_i[26];
  assign data_masked[3376] = data_i[3376] & sel_one_hot_i[26];
  assign data_masked[3375] = data_i[3375] & sel_one_hot_i[26];
  assign data_masked[3374] = data_i[3374] & sel_one_hot_i[26];
  assign data_masked[3373] = data_i[3373] & sel_one_hot_i[26];
  assign data_masked[3372] = data_i[3372] & sel_one_hot_i[26];
  assign data_masked[3371] = data_i[3371] & sel_one_hot_i[26];
  assign data_masked[3370] = data_i[3370] & sel_one_hot_i[26];
  assign data_masked[3369] = data_i[3369] & sel_one_hot_i[26];
  assign data_masked[3368] = data_i[3368] & sel_one_hot_i[26];
  assign data_masked[3367] = data_i[3367] & sel_one_hot_i[26];
  assign data_masked[3366] = data_i[3366] & sel_one_hot_i[26];
  assign data_masked[3365] = data_i[3365] & sel_one_hot_i[26];
  assign data_masked[3364] = data_i[3364] & sel_one_hot_i[26];
  assign data_masked[3363] = data_i[3363] & sel_one_hot_i[26];
  assign data_masked[3362] = data_i[3362] & sel_one_hot_i[26];
  assign data_masked[3361] = data_i[3361] & sel_one_hot_i[26];
  assign data_masked[3360] = data_i[3360] & sel_one_hot_i[26];
  assign data_masked[3359] = data_i[3359] & sel_one_hot_i[26];
  assign data_masked[3358] = data_i[3358] & sel_one_hot_i[26];
  assign data_masked[3357] = data_i[3357] & sel_one_hot_i[26];
  assign data_masked[3356] = data_i[3356] & sel_one_hot_i[26];
  assign data_masked[3355] = data_i[3355] & sel_one_hot_i[26];
  assign data_masked[3354] = data_i[3354] & sel_one_hot_i[26];
  assign data_masked[3353] = data_i[3353] & sel_one_hot_i[26];
  assign data_masked[3352] = data_i[3352] & sel_one_hot_i[26];
  assign data_masked[3351] = data_i[3351] & sel_one_hot_i[26];
  assign data_masked[3350] = data_i[3350] & sel_one_hot_i[26];
  assign data_masked[3349] = data_i[3349] & sel_one_hot_i[26];
  assign data_masked[3348] = data_i[3348] & sel_one_hot_i[26];
  assign data_masked[3347] = data_i[3347] & sel_one_hot_i[26];
  assign data_masked[3346] = data_i[3346] & sel_one_hot_i[26];
  assign data_masked[3345] = data_i[3345] & sel_one_hot_i[26];
  assign data_masked[3344] = data_i[3344] & sel_one_hot_i[26];
  assign data_masked[3343] = data_i[3343] & sel_one_hot_i[26];
  assign data_masked[3342] = data_i[3342] & sel_one_hot_i[26];
  assign data_masked[3341] = data_i[3341] & sel_one_hot_i[26];
  assign data_masked[3340] = data_i[3340] & sel_one_hot_i[26];
  assign data_masked[3339] = data_i[3339] & sel_one_hot_i[26];
  assign data_masked[3338] = data_i[3338] & sel_one_hot_i[26];
  assign data_masked[3337] = data_i[3337] & sel_one_hot_i[26];
  assign data_masked[3336] = data_i[3336] & sel_one_hot_i[26];
  assign data_masked[3335] = data_i[3335] & sel_one_hot_i[26];
  assign data_masked[3334] = data_i[3334] & sel_one_hot_i[26];
  assign data_masked[3333] = data_i[3333] & sel_one_hot_i[26];
  assign data_masked[3332] = data_i[3332] & sel_one_hot_i[26];
  assign data_masked[3331] = data_i[3331] & sel_one_hot_i[26];
  assign data_masked[3330] = data_i[3330] & sel_one_hot_i[26];
  assign data_masked[3329] = data_i[3329] & sel_one_hot_i[26];
  assign data_masked[3328] = data_i[3328] & sel_one_hot_i[26];
  assign data_masked[3583] = data_i[3583] & sel_one_hot_i[27];
  assign data_masked[3582] = data_i[3582] & sel_one_hot_i[27];
  assign data_masked[3581] = data_i[3581] & sel_one_hot_i[27];
  assign data_masked[3580] = data_i[3580] & sel_one_hot_i[27];
  assign data_masked[3579] = data_i[3579] & sel_one_hot_i[27];
  assign data_masked[3578] = data_i[3578] & sel_one_hot_i[27];
  assign data_masked[3577] = data_i[3577] & sel_one_hot_i[27];
  assign data_masked[3576] = data_i[3576] & sel_one_hot_i[27];
  assign data_masked[3575] = data_i[3575] & sel_one_hot_i[27];
  assign data_masked[3574] = data_i[3574] & sel_one_hot_i[27];
  assign data_masked[3573] = data_i[3573] & sel_one_hot_i[27];
  assign data_masked[3572] = data_i[3572] & sel_one_hot_i[27];
  assign data_masked[3571] = data_i[3571] & sel_one_hot_i[27];
  assign data_masked[3570] = data_i[3570] & sel_one_hot_i[27];
  assign data_masked[3569] = data_i[3569] & sel_one_hot_i[27];
  assign data_masked[3568] = data_i[3568] & sel_one_hot_i[27];
  assign data_masked[3567] = data_i[3567] & sel_one_hot_i[27];
  assign data_masked[3566] = data_i[3566] & sel_one_hot_i[27];
  assign data_masked[3565] = data_i[3565] & sel_one_hot_i[27];
  assign data_masked[3564] = data_i[3564] & sel_one_hot_i[27];
  assign data_masked[3563] = data_i[3563] & sel_one_hot_i[27];
  assign data_masked[3562] = data_i[3562] & sel_one_hot_i[27];
  assign data_masked[3561] = data_i[3561] & sel_one_hot_i[27];
  assign data_masked[3560] = data_i[3560] & sel_one_hot_i[27];
  assign data_masked[3559] = data_i[3559] & sel_one_hot_i[27];
  assign data_masked[3558] = data_i[3558] & sel_one_hot_i[27];
  assign data_masked[3557] = data_i[3557] & sel_one_hot_i[27];
  assign data_masked[3556] = data_i[3556] & sel_one_hot_i[27];
  assign data_masked[3555] = data_i[3555] & sel_one_hot_i[27];
  assign data_masked[3554] = data_i[3554] & sel_one_hot_i[27];
  assign data_masked[3553] = data_i[3553] & sel_one_hot_i[27];
  assign data_masked[3552] = data_i[3552] & sel_one_hot_i[27];
  assign data_masked[3551] = data_i[3551] & sel_one_hot_i[27];
  assign data_masked[3550] = data_i[3550] & sel_one_hot_i[27];
  assign data_masked[3549] = data_i[3549] & sel_one_hot_i[27];
  assign data_masked[3548] = data_i[3548] & sel_one_hot_i[27];
  assign data_masked[3547] = data_i[3547] & sel_one_hot_i[27];
  assign data_masked[3546] = data_i[3546] & sel_one_hot_i[27];
  assign data_masked[3545] = data_i[3545] & sel_one_hot_i[27];
  assign data_masked[3544] = data_i[3544] & sel_one_hot_i[27];
  assign data_masked[3543] = data_i[3543] & sel_one_hot_i[27];
  assign data_masked[3542] = data_i[3542] & sel_one_hot_i[27];
  assign data_masked[3541] = data_i[3541] & sel_one_hot_i[27];
  assign data_masked[3540] = data_i[3540] & sel_one_hot_i[27];
  assign data_masked[3539] = data_i[3539] & sel_one_hot_i[27];
  assign data_masked[3538] = data_i[3538] & sel_one_hot_i[27];
  assign data_masked[3537] = data_i[3537] & sel_one_hot_i[27];
  assign data_masked[3536] = data_i[3536] & sel_one_hot_i[27];
  assign data_masked[3535] = data_i[3535] & sel_one_hot_i[27];
  assign data_masked[3534] = data_i[3534] & sel_one_hot_i[27];
  assign data_masked[3533] = data_i[3533] & sel_one_hot_i[27];
  assign data_masked[3532] = data_i[3532] & sel_one_hot_i[27];
  assign data_masked[3531] = data_i[3531] & sel_one_hot_i[27];
  assign data_masked[3530] = data_i[3530] & sel_one_hot_i[27];
  assign data_masked[3529] = data_i[3529] & sel_one_hot_i[27];
  assign data_masked[3528] = data_i[3528] & sel_one_hot_i[27];
  assign data_masked[3527] = data_i[3527] & sel_one_hot_i[27];
  assign data_masked[3526] = data_i[3526] & sel_one_hot_i[27];
  assign data_masked[3525] = data_i[3525] & sel_one_hot_i[27];
  assign data_masked[3524] = data_i[3524] & sel_one_hot_i[27];
  assign data_masked[3523] = data_i[3523] & sel_one_hot_i[27];
  assign data_masked[3522] = data_i[3522] & sel_one_hot_i[27];
  assign data_masked[3521] = data_i[3521] & sel_one_hot_i[27];
  assign data_masked[3520] = data_i[3520] & sel_one_hot_i[27];
  assign data_masked[3519] = data_i[3519] & sel_one_hot_i[27];
  assign data_masked[3518] = data_i[3518] & sel_one_hot_i[27];
  assign data_masked[3517] = data_i[3517] & sel_one_hot_i[27];
  assign data_masked[3516] = data_i[3516] & sel_one_hot_i[27];
  assign data_masked[3515] = data_i[3515] & sel_one_hot_i[27];
  assign data_masked[3514] = data_i[3514] & sel_one_hot_i[27];
  assign data_masked[3513] = data_i[3513] & sel_one_hot_i[27];
  assign data_masked[3512] = data_i[3512] & sel_one_hot_i[27];
  assign data_masked[3511] = data_i[3511] & sel_one_hot_i[27];
  assign data_masked[3510] = data_i[3510] & sel_one_hot_i[27];
  assign data_masked[3509] = data_i[3509] & sel_one_hot_i[27];
  assign data_masked[3508] = data_i[3508] & sel_one_hot_i[27];
  assign data_masked[3507] = data_i[3507] & sel_one_hot_i[27];
  assign data_masked[3506] = data_i[3506] & sel_one_hot_i[27];
  assign data_masked[3505] = data_i[3505] & sel_one_hot_i[27];
  assign data_masked[3504] = data_i[3504] & sel_one_hot_i[27];
  assign data_masked[3503] = data_i[3503] & sel_one_hot_i[27];
  assign data_masked[3502] = data_i[3502] & sel_one_hot_i[27];
  assign data_masked[3501] = data_i[3501] & sel_one_hot_i[27];
  assign data_masked[3500] = data_i[3500] & sel_one_hot_i[27];
  assign data_masked[3499] = data_i[3499] & sel_one_hot_i[27];
  assign data_masked[3498] = data_i[3498] & sel_one_hot_i[27];
  assign data_masked[3497] = data_i[3497] & sel_one_hot_i[27];
  assign data_masked[3496] = data_i[3496] & sel_one_hot_i[27];
  assign data_masked[3495] = data_i[3495] & sel_one_hot_i[27];
  assign data_masked[3494] = data_i[3494] & sel_one_hot_i[27];
  assign data_masked[3493] = data_i[3493] & sel_one_hot_i[27];
  assign data_masked[3492] = data_i[3492] & sel_one_hot_i[27];
  assign data_masked[3491] = data_i[3491] & sel_one_hot_i[27];
  assign data_masked[3490] = data_i[3490] & sel_one_hot_i[27];
  assign data_masked[3489] = data_i[3489] & sel_one_hot_i[27];
  assign data_masked[3488] = data_i[3488] & sel_one_hot_i[27];
  assign data_masked[3487] = data_i[3487] & sel_one_hot_i[27];
  assign data_masked[3486] = data_i[3486] & sel_one_hot_i[27];
  assign data_masked[3485] = data_i[3485] & sel_one_hot_i[27];
  assign data_masked[3484] = data_i[3484] & sel_one_hot_i[27];
  assign data_masked[3483] = data_i[3483] & sel_one_hot_i[27];
  assign data_masked[3482] = data_i[3482] & sel_one_hot_i[27];
  assign data_masked[3481] = data_i[3481] & sel_one_hot_i[27];
  assign data_masked[3480] = data_i[3480] & sel_one_hot_i[27];
  assign data_masked[3479] = data_i[3479] & sel_one_hot_i[27];
  assign data_masked[3478] = data_i[3478] & sel_one_hot_i[27];
  assign data_masked[3477] = data_i[3477] & sel_one_hot_i[27];
  assign data_masked[3476] = data_i[3476] & sel_one_hot_i[27];
  assign data_masked[3475] = data_i[3475] & sel_one_hot_i[27];
  assign data_masked[3474] = data_i[3474] & sel_one_hot_i[27];
  assign data_masked[3473] = data_i[3473] & sel_one_hot_i[27];
  assign data_masked[3472] = data_i[3472] & sel_one_hot_i[27];
  assign data_masked[3471] = data_i[3471] & sel_one_hot_i[27];
  assign data_masked[3470] = data_i[3470] & sel_one_hot_i[27];
  assign data_masked[3469] = data_i[3469] & sel_one_hot_i[27];
  assign data_masked[3468] = data_i[3468] & sel_one_hot_i[27];
  assign data_masked[3467] = data_i[3467] & sel_one_hot_i[27];
  assign data_masked[3466] = data_i[3466] & sel_one_hot_i[27];
  assign data_masked[3465] = data_i[3465] & sel_one_hot_i[27];
  assign data_masked[3464] = data_i[3464] & sel_one_hot_i[27];
  assign data_masked[3463] = data_i[3463] & sel_one_hot_i[27];
  assign data_masked[3462] = data_i[3462] & sel_one_hot_i[27];
  assign data_masked[3461] = data_i[3461] & sel_one_hot_i[27];
  assign data_masked[3460] = data_i[3460] & sel_one_hot_i[27];
  assign data_masked[3459] = data_i[3459] & sel_one_hot_i[27];
  assign data_masked[3458] = data_i[3458] & sel_one_hot_i[27];
  assign data_masked[3457] = data_i[3457] & sel_one_hot_i[27];
  assign data_masked[3456] = data_i[3456] & sel_one_hot_i[27];
  assign data_masked[3711] = data_i[3711] & sel_one_hot_i[28];
  assign data_masked[3710] = data_i[3710] & sel_one_hot_i[28];
  assign data_masked[3709] = data_i[3709] & sel_one_hot_i[28];
  assign data_masked[3708] = data_i[3708] & sel_one_hot_i[28];
  assign data_masked[3707] = data_i[3707] & sel_one_hot_i[28];
  assign data_masked[3706] = data_i[3706] & sel_one_hot_i[28];
  assign data_masked[3705] = data_i[3705] & sel_one_hot_i[28];
  assign data_masked[3704] = data_i[3704] & sel_one_hot_i[28];
  assign data_masked[3703] = data_i[3703] & sel_one_hot_i[28];
  assign data_masked[3702] = data_i[3702] & sel_one_hot_i[28];
  assign data_masked[3701] = data_i[3701] & sel_one_hot_i[28];
  assign data_masked[3700] = data_i[3700] & sel_one_hot_i[28];
  assign data_masked[3699] = data_i[3699] & sel_one_hot_i[28];
  assign data_masked[3698] = data_i[3698] & sel_one_hot_i[28];
  assign data_masked[3697] = data_i[3697] & sel_one_hot_i[28];
  assign data_masked[3696] = data_i[3696] & sel_one_hot_i[28];
  assign data_masked[3695] = data_i[3695] & sel_one_hot_i[28];
  assign data_masked[3694] = data_i[3694] & sel_one_hot_i[28];
  assign data_masked[3693] = data_i[3693] & sel_one_hot_i[28];
  assign data_masked[3692] = data_i[3692] & sel_one_hot_i[28];
  assign data_masked[3691] = data_i[3691] & sel_one_hot_i[28];
  assign data_masked[3690] = data_i[3690] & sel_one_hot_i[28];
  assign data_masked[3689] = data_i[3689] & sel_one_hot_i[28];
  assign data_masked[3688] = data_i[3688] & sel_one_hot_i[28];
  assign data_masked[3687] = data_i[3687] & sel_one_hot_i[28];
  assign data_masked[3686] = data_i[3686] & sel_one_hot_i[28];
  assign data_masked[3685] = data_i[3685] & sel_one_hot_i[28];
  assign data_masked[3684] = data_i[3684] & sel_one_hot_i[28];
  assign data_masked[3683] = data_i[3683] & sel_one_hot_i[28];
  assign data_masked[3682] = data_i[3682] & sel_one_hot_i[28];
  assign data_masked[3681] = data_i[3681] & sel_one_hot_i[28];
  assign data_masked[3680] = data_i[3680] & sel_one_hot_i[28];
  assign data_masked[3679] = data_i[3679] & sel_one_hot_i[28];
  assign data_masked[3678] = data_i[3678] & sel_one_hot_i[28];
  assign data_masked[3677] = data_i[3677] & sel_one_hot_i[28];
  assign data_masked[3676] = data_i[3676] & sel_one_hot_i[28];
  assign data_masked[3675] = data_i[3675] & sel_one_hot_i[28];
  assign data_masked[3674] = data_i[3674] & sel_one_hot_i[28];
  assign data_masked[3673] = data_i[3673] & sel_one_hot_i[28];
  assign data_masked[3672] = data_i[3672] & sel_one_hot_i[28];
  assign data_masked[3671] = data_i[3671] & sel_one_hot_i[28];
  assign data_masked[3670] = data_i[3670] & sel_one_hot_i[28];
  assign data_masked[3669] = data_i[3669] & sel_one_hot_i[28];
  assign data_masked[3668] = data_i[3668] & sel_one_hot_i[28];
  assign data_masked[3667] = data_i[3667] & sel_one_hot_i[28];
  assign data_masked[3666] = data_i[3666] & sel_one_hot_i[28];
  assign data_masked[3665] = data_i[3665] & sel_one_hot_i[28];
  assign data_masked[3664] = data_i[3664] & sel_one_hot_i[28];
  assign data_masked[3663] = data_i[3663] & sel_one_hot_i[28];
  assign data_masked[3662] = data_i[3662] & sel_one_hot_i[28];
  assign data_masked[3661] = data_i[3661] & sel_one_hot_i[28];
  assign data_masked[3660] = data_i[3660] & sel_one_hot_i[28];
  assign data_masked[3659] = data_i[3659] & sel_one_hot_i[28];
  assign data_masked[3658] = data_i[3658] & sel_one_hot_i[28];
  assign data_masked[3657] = data_i[3657] & sel_one_hot_i[28];
  assign data_masked[3656] = data_i[3656] & sel_one_hot_i[28];
  assign data_masked[3655] = data_i[3655] & sel_one_hot_i[28];
  assign data_masked[3654] = data_i[3654] & sel_one_hot_i[28];
  assign data_masked[3653] = data_i[3653] & sel_one_hot_i[28];
  assign data_masked[3652] = data_i[3652] & sel_one_hot_i[28];
  assign data_masked[3651] = data_i[3651] & sel_one_hot_i[28];
  assign data_masked[3650] = data_i[3650] & sel_one_hot_i[28];
  assign data_masked[3649] = data_i[3649] & sel_one_hot_i[28];
  assign data_masked[3648] = data_i[3648] & sel_one_hot_i[28];
  assign data_masked[3647] = data_i[3647] & sel_one_hot_i[28];
  assign data_masked[3646] = data_i[3646] & sel_one_hot_i[28];
  assign data_masked[3645] = data_i[3645] & sel_one_hot_i[28];
  assign data_masked[3644] = data_i[3644] & sel_one_hot_i[28];
  assign data_masked[3643] = data_i[3643] & sel_one_hot_i[28];
  assign data_masked[3642] = data_i[3642] & sel_one_hot_i[28];
  assign data_masked[3641] = data_i[3641] & sel_one_hot_i[28];
  assign data_masked[3640] = data_i[3640] & sel_one_hot_i[28];
  assign data_masked[3639] = data_i[3639] & sel_one_hot_i[28];
  assign data_masked[3638] = data_i[3638] & sel_one_hot_i[28];
  assign data_masked[3637] = data_i[3637] & sel_one_hot_i[28];
  assign data_masked[3636] = data_i[3636] & sel_one_hot_i[28];
  assign data_masked[3635] = data_i[3635] & sel_one_hot_i[28];
  assign data_masked[3634] = data_i[3634] & sel_one_hot_i[28];
  assign data_masked[3633] = data_i[3633] & sel_one_hot_i[28];
  assign data_masked[3632] = data_i[3632] & sel_one_hot_i[28];
  assign data_masked[3631] = data_i[3631] & sel_one_hot_i[28];
  assign data_masked[3630] = data_i[3630] & sel_one_hot_i[28];
  assign data_masked[3629] = data_i[3629] & sel_one_hot_i[28];
  assign data_masked[3628] = data_i[3628] & sel_one_hot_i[28];
  assign data_masked[3627] = data_i[3627] & sel_one_hot_i[28];
  assign data_masked[3626] = data_i[3626] & sel_one_hot_i[28];
  assign data_masked[3625] = data_i[3625] & sel_one_hot_i[28];
  assign data_masked[3624] = data_i[3624] & sel_one_hot_i[28];
  assign data_masked[3623] = data_i[3623] & sel_one_hot_i[28];
  assign data_masked[3622] = data_i[3622] & sel_one_hot_i[28];
  assign data_masked[3621] = data_i[3621] & sel_one_hot_i[28];
  assign data_masked[3620] = data_i[3620] & sel_one_hot_i[28];
  assign data_masked[3619] = data_i[3619] & sel_one_hot_i[28];
  assign data_masked[3618] = data_i[3618] & sel_one_hot_i[28];
  assign data_masked[3617] = data_i[3617] & sel_one_hot_i[28];
  assign data_masked[3616] = data_i[3616] & sel_one_hot_i[28];
  assign data_masked[3615] = data_i[3615] & sel_one_hot_i[28];
  assign data_masked[3614] = data_i[3614] & sel_one_hot_i[28];
  assign data_masked[3613] = data_i[3613] & sel_one_hot_i[28];
  assign data_masked[3612] = data_i[3612] & sel_one_hot_i[28];
  assign data_masked[3611] = data_i[3611] & sel_one_hot_i[28];
  assign data_masked[3610] = data_i[3610] & sel_one_hot_i[28];
  assign data_masked[3609] = data_i[3609] & sel_one_hot_i[28];
  assign data_masked[3608] = data_i[3608] & sel_one_hot_i[28];
  assign data_masked[3607] = data_i[3607] & sel_one_hot_i[28];
  assign data_masked[3606] = data_i[3606] & sel_one_hot_i[28];
  assign data_masked[3605] = data_i[3605] & sel_one_hot_i[28];
  assign data_masked[3604] = data_i[3604] & sel_one_hot_i[28];
  assign data_masked[3603] = data_i[3603] & sel_one_hot_i[28];
  assign data_masked[3602] = data_i[3602] & sel_one_hot_i[28];
  assign data_masked[3601] = data_i[3601] & sel_one_hot_i[28];
  assign data_masked[3600] = data_i[3600] & sel_one_hot_i[28];
  assign data_masked[3599] = data_i[3599] & sel_one_hot_i[28];
  assign data_masked[3598] = data_i[3598] & sel_one_hot_i[28];
  assign data_masked[3597] = data_i[3597] & sel_one_hot_i[28];
  assign data_masked[3596] = data_i[3596] & sel_one_hot_i[28];
  assign data_masked[3595] = data_i[3595] & sel_one_hot_i[28];
  assign data_masked[3594] = data_i[3594] & sel_one_hot_i[28];
  assign data_masked[3593] = data_i[3593] & sel_one_hot_i[28];
  assign data_masked[3592] = data_i[3592] & sel_one_hot_i[28];
  assign data_masked[3591] = data_i[3591] & sel_one_hot_i[28];
  assign data_masked[3590] = data_i[3590] & sel_one_hot_i[28];
  assign data_masked[3589] = data_i[3589] & sel_one_hot_i[28];
  assign data_masked[3588] = data_i[3588] & sel_one_hot_i[28];
  assign data_masked[3587] = data_i[3587] & sel_one_hot_i[28];
  assign data_masked[3586] = data_i[3586] & sel_one_hot_i[28];
  assign data_masked[3585] = data_i[3585] & sel_one_hot_i[28];
  assign data_masked[3584] = data_i[3584] & sel_one_hot_i[28];
  assign data_masked[3839] = data_i[3839] & sel_one_hot_i[29];
  assign data_masked[3838] = data_i[3838] & sel_one_hot_i[29];
  assign data_masked[3837] = data_i[3837] & sel_one_hot_i[29];
  assign data_masked[3836] = data_i[3836] & sel_one_hot_i[29];
  assign data_masked[3835] = data_i[3835] & sel_one_hot_i[29];
  assign data_masked[3834] = data_i[3834] & sel_one_hot_i[29];
  assign data_masked[3833] = data_i[3833] & sel_one_hot_i[29];
  assign data_masked[3832] = data_i[3832] & sel_one_hot_i[29];
  assign data_masked[3831] = data_i[3831] & sel_one_hot_i[29];
  assign data_masked[3830] = data_i[3830] & sel_one_hot_i[29];
  assign data_masked[3829] = data_i[3829] & sel_one_hot_i[29];
  assign data_masked[3828] = data_i[3828] & sel_one_hot_i[29];
  assign data_masked[3827] = data_i[3827] & sel_one_hot_i[29];
  assign data_masked[3826] = data_i[3826] & sel_one_hot_i[29];
  assign data_masked[3825] = data_i[3825] & sel_one_hot_i[29];
  assign data_masked[3824] = data_i[3824] & sel_one_hot_i[29];
  assign data_masked[3823] = data_i[3823] & sel_one_hot_i[29];
  assign data_masked[3822] = data_i[3822] & sel_one_hot_i[29];
  assign data_masked[3821] = data_i[3821] & sel_one_hot_i[29];
  assign data_masked[3820] = data_i[3820] & sel_one_hot_i[29];
  assign data_masked[3819] = data_i[3819] & sel_one_hot_i[29];
  assign data_masked[3818] = data_i[3818] & sel_one_hot_i[29];
  assign data_masked[3817] = data_i[3817] & sel_one_hot_i[29];
  assign data_masked[3816] = data_i[3816] & sel_one_hot_i[29];
  assign data_masked[3815] = data_i[3815] & sel_one_hot_i[29];
  assign data_masked[3814] = data_i[3814] & sel_one_hot_i[29];
  assign data_masked[3813] = data_i[3813] & sel_one_hot_i[29];
  assign data_masked[3812] = data_i[3812] & sel_one_hot_i[29];
  assign data_masked[3811] = data_i[3811] & sel_one_hot_i[29];
  assign data_masked[3810] = data_i[3810] & sel_one_hot_i[29];
  assign data_masked[3809] = data_i[3809] & sel_one_hot_i[29];
  assign data_masked[3808] = data_i[3808] & sel_one_hot_i[29];
  assign data_masked[3807] = data_i[3807] & sel_one_hot_i[29];
  assign data_masked[3806] = data_i[3806] & sel_one_hot_i[29];
  assign data_masked[3805] = data_i[3805] & sel_one_hot_i[29];
  assign data_masked[3804] = data_i[3804] & sel_one_hot_i[29];
  assign data_masked[3803] = data_i[3803] & sel_one_hot_i[29];
  assign data_masked[3802] = data_i[3802] & sel_one_hot_i[29];
  assign data_masked[3801] = data_i[3801] & sel_one_hot_i[29];
  assign data_masked[3800] = data_i[3800] & sel_one_hot_i[29];
  assign data_masked[3799] = data_i[3799] & sel_one_hot_i[29];
  assign data_masked[3798] = data_i[3798] & sel_one_hot_i[29];
  assign data_masked[3797] = data_i[3797] & sel_one_hot_i[29];
  assign data_masked[3796] = data_i[3796] & sel_one_hot_i[29];
  assign data_masked[3795] = data_i[3795] & sel_one_hot_i[29];
  assign data_masked[3794] = data_i[3794] & sel_one_hot_i[29];
  assign data_masked[3793] = data_i[3793] & sel_one_hot_i[29];
  assign data_masked[3792] = data_i[3792] & sel_one_hot_i[29];
  assign data_masked[3791] = data_i[3791] & sel_one_hot_i[29];
  assign data_masked[3790] = data_i[3790] & sel_one_hot_i[29];
  assign data_masked[3789] = data_i[3789] & sel_one_hot_i[29];
  assign data_masked[3788] = data_i[3788] & sel_one_hot_i[29];
  assign data_masked[3787] = data_i[3787] & sel_one_hot_i[29];
  assign data_masked[3786] = data_i[3786] & sel_one_hot_i[29];
  assign data_masked[3785] = data_i[3785] & sel_one_hot_i[29];
  assign data_masked[3784] = data_i[3784] & sel_one_hot_i[29];
  assign data_masked[3783] = data_i[3783] & sel_one_hot_i[29];
  assign data_masked[3782] = data_i[3782] & sel_one_hot_i[29];
  assign data_masked[3781] = data_i[3781] & sel_one_hot_i[29];
  assign data_masked[3780] = data_i[3780] & sel_one_hot_i[29];
  assign data_masked[3779] = data_i[3779] & sel_one_hot_i[29];
  assign data_masked[3778] = data_i[3778] & sel_one_hot_i[29];
  assign data_masked[3777] = data_i[3777] & sel_one_hot_i[29];
  assign data_masked[3776] = data_i[3776] & sel_one_hot_i[29];
  assign data_masked[3775] = data_i[3775] & sel_one_hot_i[29];
  assign data_masked[3774] = data_i[3774] & sel_one_hot_i[29];
  assign data_masked[3773] = data_i[3773] & sel_one_hot_i[29];
  assign data_masked[3772] = data_i[3772] & sel_one_hot_i[29];
  assign data_masked[3771] = data_i[3771] & sel_one_hot_i[29];
  assign data_masked[3770] = data_i[3770] & sel_one_hot_i[29];
  assign data_masked[3769] = data_i[3769] & sel_one_hot_i[29];
  assign data_masked[3768] = data_i[3768] & sel_one_hot_i[29];
  assign data_masked[3767] = data_i[3767] & sel_one_hot_i[29];
  assign data_masked[3766] = data_i[3766] & sel_one_hot_i[29];
  assign data_masked[3765] = data_i[3765] & sel_one_hot_i[29];
  assign data_masked[3764] = data_i[3764] & sel_one_hot_i[29];
  assign data_masked[3763] = data_i[3763] & sel_one_hot_i[29];
  assign data_masked[3762] = data_i[3762] & sel_one_hot_i[29];
  assign data_masked[3761] = data_i[3761] & sel_one_hot_i[29];
  assign data_masked[3760] = data_i[3760] & sel_one_hot_i[29];
  assign data_masked[3759] = data_i[3759] & sel_one_hot_i[29];
  assign data_masked[3758] = data_i[3758] & sel_one_hot_i[29];
  assign data_masked[3757] = data_i[3757] & sel_one_hot_i[29];
  assign data_masked[3756] = data_i[3756] & sel_one_hot_i[29];
  assign data_masked[3755] = data_i[3755] & sel_one_hot_i[29];
  assign data_masked[3754] = data_i[3754] & sel_one_hot_i[29];
  assign data_masked[3753] = data_i[3753] & sel_one_hot_i[29];
  assign data_masked[3752] = data_i[3752] & sel_one_hot_i[29];
  assign data_masked[3751] = data_i[3751] & sel_one_hot_i[29];
  assign data_masked[3750] = data_i[3750] & sel_one_hot_i[29];
  assign data_masked[3749] = data_i[3749] & sel_one_hot_i[29];
  assign data_masked[3748] = data_i[3748] & sel_one_hot_i[29];
  assign data_masked[3747] = data_i[3747] & sel_one_hot_i[29];
  assign data_masked[3746] = data_i[3746] & sel_one_hot_i[29];
  assign data_masked[3745] = data_i[3745] & sel_one_hot_i[29];
  assign data_masked[3744] = data_i[3744] & sel_one_hot_i[29];
  assign data_masked[3743] = data_i[3743] & sel_one_hot_i[29];
  assign data_masked[3742] = data_i[3742] & sel_one_hot_i[29];
  assign data_masked[3741] = data_i[3741] & sel_one_hot_i[29];
  assign data_masked[3740] = data_i[3740] & sel_one_hot_i[29];
  assign data_masked[3739] = data_i[3739] & sel_one_hot_i[29];
  assign data_masked[3738] = data_i[3738] & sel_one_hot_i[29];
  assign data_masked[3737] = data_i[3737] & sel_one_hot_i[29];
  assign data_masked[3736] = data_i[3736] & sel_one_hot_i[29];
  assign data_masked[3735] = data_i[3735] & sel_one_hot_i[29];
  assign data_masked[3734] = data_i[3734] & sel_one_hot_i[29];
  assign data_masked[3733] = data_i[3733] & sel_one_hot_i[29];
  assign data_masked[3732] = data_i[3732] & sel_one_hot_i[29];
  assign data_masked[3731] = data_i[3731] & sel_one_hot_i[29];
  assign data_masked[3730] = data_i[3730] & sel_one_hot_i[29];
  assign data_masked[3729] = data_i[3729] & sel_one_hot_i[29];
  assign data_masked[3728] = data_i[3728] & sel_one_hot_i[29];
  assign data_masked[3727] = data_i[3727] & sel_one_hot_i[29];
  assign data_masked[3726] = data_i[3726] & sel_one_hot_i[29];
  assign data_masked[3725] = data_i[3725] & sel_one_hot_i[29];
  assign data_masked[3724] = data_i[3724] & sel_one_hot_i[29];
  assign data_masked[3723] = data_i[3723] & sel_one_hot_i[29];
  assign data_masked[3722] = data_i[3722] & sel_one_hot_i[29];
  assign data_masked[3721] = data_i[3721] & sel_one_hot_i[29];
  assign data_masked[3720] = data_i[3720] & sel_one_hot_i[29];
  assign data_masked[3719] = data_i[3719] & sel_one_hot_i[29];
  assign data_masked[3718] = data_i[3718] & sel_one_hot_i[29];
  assign data_masked[3717] = data_i[3717] & sel_one_hot_i[29];
  assign data_masked[3716] = data_i[3716] & sel_one_hot_i[29];
  assign data_masked[3715] = data_i[3715] & sel_one_hot_i[29];
  assign data_masked[3714] = data_i[3714] & sel_one_hot_i[29];
  assign data_masked[3713] = data_i[3713] & sel_one_hot_i[29];
  assign data_masked[3712] = data_i[3712] & sel_one_hot_i[29];
  assign data_masked[3967] = data_i[3967] & sel_one_hot_i[30];
  assign data_masked[3966] = data_i[3966] & sel_one_hot_i[30];
  assign data_masked[3965] = data_i[3965] & sel_one_hot_i[30];
  assign data_masked[3964] = data_i[3964] & sel_one_hot_i[30];
  assign data_masked[3963] = data_i[3963] & sel_one_hot_i[30];
  assign data_masked[3962] = data_i[3962] & sel_one_hot_i[30];
  assign data_masked[3961] = data_i[3961] & sel_one_hot_i[30];
  assign data_masked[3960] = data_i[3960] & sel_one_hot_i[30];
  assign data_masked[3959] = data_i[3959] & sel_one_hot_i[30];
  assign data_masked[3958] = data_i[3958] & sel_one_hot_i[30];
  assign data_masked[3957] = data_i[3957] & sel_one_hot_i[30];
  assign data_masked[3956] = data_i[3956] & sel_one_hot_i[30];
  assign data_masked[3955] = data_i[3955] & sel_one_hot_i[30];
  assign data_masked[3954] = data_i[3954] & sel_one_hot_i[30];
  assign data_masked[3953] = data_i[3953] & sel_one_hot_i[30];
  assign data_masked[3952] = data_i[3952] & sel_one_hot_i[30];
  assign data_masked[3951] = data_i[3951] & sel_one_hot_i[30];
  assign data_masked[3950] = data_i[3950] & sel_one_hot_i[30];
  assign data_masked[3949] = data_i[3949] & sel_one_hot_i[30];
  assign data_masked[3948] = data_i[3948] & sel_one_hot_i[30];
  assign data_masked[3947] = data_i[3947] & sel_one_hot_i[30];
  assign data_masked[3946] = data_i[3946] & sel_one_hot_i[30];
  assign data_masked[3945] = data_i[3945] & sel_one_hot_i[30];
  assign data_masked[3944] = data_i[3944] & sel_one_hot_i[30];
  assign data_masked[3943] = data_i[3943] & sel_one_hot_i[30];
  assign data_masked[3942] = data_i[3942] & sel_one_hot_i[30];
  assign data_masked[3941] = data_i[3941] & sel_one_hot_i[30];
  assign data_masked[3940] = data_i[3940] & sel_one_hot_i[30];
  assign data_masked[3939] = data_i[3939] & sel_one_hot_i[30];
  assign data_masked[3938] = data_i[3938] & sel_one_hot_i[30];
  assign data_masked[3937] = data_i[3937] & sel_one_hot_i[30];
  assign data_masked[3936] = data_i[3936] & sel_one_hot_i[30];
  assign data_masked[3935] = data_i[3935] & sel_one_hot_i[30];
  assign data_masked[3934] = data_i[3934] & sel_one_hot_i[30];
  assign data_masked[3933] = data_i[3933] & sel_one_hot_i[30];
  assign data_masked[3932] = data_i[3932] & sel_one_hot_i[30];
  assign data_masked[3931] = data_i[3931] & sel_one_hot_i[30];
  assign data_masked[3930] = data_i[3930] & sel_one_hot_i[30];
  assign data_masked[3929] = data_i[3929] & sel_one_hot_i[30];
  assign data_masked[3928] = data_i[3928] & sel_one_hot_i[30];
  assign data_masked[3927] = data_i[3927] & sel_one_hot_i[30];
  assign data_masked[3926] = data_i[3926] & sel_one_hot_i[30];
  assign data_masked[3925] = data_i[3925] & sel_one_hot_i[30];
  assign data_masked[3924] = data_i[3924] & sel_one_hot_i[30];
  assign data_masked[3923] = data_i[3923] & sel_one_hot_i[30];
  assign data_masked[3922] = data_i[3922] & sel_one_hot_i[30];
  assign data_masked[3921] = data_i[3921] & sel_one_hot_i[30];
  assign data_masked[3920] = data_i[3920] & sel_one_hot_i[30];
  assign data_masked[3919] = data_i[3919] & sel_one_hot_i[30];
  assign data_masked[3918] = data_i[3918] & sel_one_hot_i[30];
  assign data_masked[3917] = data_i[3917] & sel_one_hot_i[30];
  assign data_masked[3916] = data_i[3916] & sel_one_hot_i[30];
  assign data_masked[3915] = data_i[3915] & sel_one_hot_i[30];
  assign data_masked[3914] = data_i[3914] & sel_one_hot_i[30];
  assign data_masked[3913] = data_i[3913] & sel_one_hot_i[30];
  assign data_masked[3912] = data_i[3912] & sel_one_hot_i[30];
  assign data_masked[3911] = data_i[3911] & sel_one_hot_i[30];
  assign data_masked[3910] = data_i[3910] & sel_one_hot_i[30];
  assign data_masked[3909] = data_i[3909] & sel_one_hot_i[30];
  assign data_masked[3908] = data_i[3908] & sel_one_hot_i[30];
  assign data_masked[3907] = data_i[3907] & sel_one_hot_i[30];
  assign data_masked[3906] = data_i[3906] & sel_one_hot_i[30];
  assign data_masked[3905] = data_i[3905] & sel_one_hot_i[30];
  assign data_masked[3904] = data_i[3904] & sel_one_hot_i[30];
  assign data_masked[3903] = data_i[3903] & sel_one_hot_i[30];
  assign data_masked[3902] = data_i[3902] & sel_one_hot_i[30];
  assign data_masked[3901] = data_i[3901] & sel_one_hot_i[30];
  assign data_masked[3900] = data_i[3900] & sel_one_hot_i[30];
  assign data_masked[3899] = data_i[3899] & sel_one_hot_i[30];
  assign data_masked[3898] = data_i[3898] & sel_one_hot_i[30];
  assign data_masked[3897] = data_i[3897] & sel_one_hot_i[30];
  assign data_masked[3896] = data_i[3896] & sel_one_hot_i[30];
  assign data_masked[3895] = data_i[3895] & sel_one_hot_i[30];
  assign data_masked[3894] = data_i[3894] & sel_one_hot_i[30];
  assign data_masked[3893] = data_i[3893] & sel_one_hot_i[30];
  assign data_masked[3892] = data_i[3892] & sel_one_hot_i[30];
  assign data_masked[3891] = data_i[3891] & sel_one_hot_i[30];
  assign data_masked[3890] = data_i[3890] & sel_one_hot_i[30];
  assign data_masked[3889] = data_i[3889] & sel_one_hot_i[30];
  assign data_masked[3888] = data_i[3888] & sel_one_hot_i[30];
  assign data_masked[3887] = data_i[3887] & sel_one_hot_i[30];
  assign data_masked[3886] = data_i[3886] & sel_one_hot_i[30];
  assign data_masked[3885] = data_i[3885] & sel_one_hot_i[30];
  assign data_masked[3884] = data_i[3884] & sel_one_hot_i[30];
  assign data_masked[3883] = data_i[3883] & sel_one_hot_i[30];
  assign data_masked[3882] = data_i[3882] & sel_one_hot_i[30];
  assign data_masked[3881] = data_i[3881] & sel_one_hot_i[30];
  assign data_masked[3880] = data_i[3880] & sel_one_hot_i[30];
  assign data_masked[3879] = data_i[3879] & sel_one_hot_i[30];
  assign data_masked[3878] = data_i[3878] & sel_one_hot_i[30];
  assign data_masked[3877] = data_i[3877] & sel_one_hot_i[30];
  assign data_masked[3876] = data_i[3876] & sel_one_hot_i[30];
  assign data_masked[3875] = data_i[3875] & sel_one_hot_i[30];
  assign data_masked[3874] = data_i[3874] & sel_one_hot_i[30];
  assign data_masked[3873] = data_i[3873] & sel_one_hot_i[30];
  assign data_masked[3872] = data_i[3872] & sel_one_hot_i[30];
  assign data_masked[3871] = data_i[3871] & sel_one_hot_i[30];
  assign data_masked[3870] = data_i[3870] & sel_one_hot_i[30];
  assign data_masked[3869] = data_i[3869] & sel_one_hot_i[30];
  assign data_masked[3868] = data_i[3868] & sel_one_hot_i[30];
  assign data_masked[3867] = data_i[3867] & sel_one_hot_i[30];
  assign data_masked[3866] = data_i[3866] & sel_one_hot_i[30];
  assign data_masked[3865] = data_i[3865] & sel_one_hot_i[30];
  assign data_masked[3864] = data_i[3864] & sel_one_hot_i[30];
  assign data_masked[3863] = data_i[3863] & sel_one_hot_i[30];
  assign data_masked[3862] = data_i[3862] & sel_one_hot_i[30];
  assign data_masked[3861] = data_i[3861] & sel_one_hot_i[30];
  assign data_masked[3860] = data_i[3860] & sel_one_hot_i[30];
  assign data_masked[3859] = data_i[3859] & sel_one_hot_i[30];
  assign data_masked[3858] = data_i[3858] & sel_one_hot_i[30];
  assign data_masked[3857] = data_i[3857] & sel_one_hot_i[30];
  assign data_masked[3856] = data_i[3856] & sel_one_hot_i[30];
  assign data_masked[3855] = data_i[3855] & sel_one_hot_i[30];
  assign data_masked[3854] = data_i[3854] & sel_one_hot_i[30];
  assign data_masked[3853] = data_i[3853] & sel_one_hot_i[30];
  assign data_masked[3852] = data_i[3852] & sel_one_hot_i[30];
  assign data_masked[3851] = data_i[3851] & sel_one_hot_i[30];
  assign data_masked[3850] = data_i[3850] & sel_one_hot_i[30];
  assign data_masked[3849] = data_i[3849] & sel_one_hot_i[30];
  assign data_masked[3848] = data_i[3848] & sel_one_hot_i[30];
  assign data_masked[3847] = data_i[3847] & sel_one_hot_i[30];
  assign data_masked[3846] = data_i[3846] & sel_one_hot_i[30];
  assign data_masked[3845] = data_i[3845] & sel_one_hot_i[30];
  assign data_masked[3844] = data_i[3844] & sel_one_hot_i[30];
  assign data_masked[3843] = data_i[3843] & sel_one_hot_i[30];
  assign data_masked[3842] = data_i[3842] & sel_one_hot_i[30];
  assign data_masked[3841] = data_i[3841] & sel_one_hot_i[30];
  assign data_masked[3840] = data_i[3840] & sel_one_hot_i[30];
  assign data_masked[4095] = data_i[4095] & sel_one_hot_i[31];
  assign data_masked[4094] = data_i[4094] & sel_one_hot_i[31];
  assign data_masked[4093] = data_i[4093] & sel_one_hot_i[31];
  assign data_masked[4092] = data_i[4092] & sel_one_hot_i[31];
  assign data_masked[4091] = data_i[4091] & sel_one_hot_i[31];
  assign data_masked[4090] = data_i[4090] & sel_one_hot_i[31];
  assign data_masked[4089] = data_i[4089] & sel_one_hot_i[31];
  assign data_masked[4088] = data_i[4088] & sel_one_hot_i[31];
  assign data_masked[4087] = data_i[4087] & sel_one_hot_i[31];
  assign data_masked[4086] = data_i[4086] & sel_one_hot_i[31];
  assign data_masked[4085] = data_i[4085] & sel_one_hot_i[31];
  assign data_masked[4084] = data_i[4084] & sel_one_hot_i[31];
  assign data_masked[4083] = data_i[4083] & sel_one_hot_i[31];
  assign data_masked[4082] = data_i[4082] & sel_one_hot_i[31];
  assign data_masked[4081] = data_i[4081] & sel_one_hot_i[31];
  assign data_masked[4080] = data_i[4080] & sel_one_hot_i[31];
  assign data_masked[4079] = data_i[4079] & sel_one_hot_i[31];
  assign data_masked[4078] = data_i[4078] & sel_one_hot_i[31];
  assign data_masked[4077] = data_i[4077] & sel_one_hot_i[31];
  assign data_masked[4076] = data_i[4076] & sel_one_hot_i[31];
  assign data_masked[4075] = data_i[4075] & sel_one_hot_i[31];
  assign data_masked[4074] = data_i[4074] & sel_one_hot_i[31];
  assign data_masked[4073] = data_i[4073] & sel_one_hot_i[31];
  assign data_masked[4072] = data_i[4072] & sel_one_hot_i[31];
  assign data_masked[4071] = data_i[4071] & sel_one_hot_i[31];
  assign data_masked[4070] = data_i[4070] & sel_one_hot_i[31];
  assign data_masked[4069] = data_i[4069] & sel_one_hot_i[31];
  assign data_masked[4068] = data_i[4068] & sel_one_hot_i[31];
  assign data_masked[4067] = data_i[4067] & sel_one_hot_i[31];
  assign data_masked[4066] = data_i[4066] & sel_one_hot_i[31];
  assign data_masked[4065] = data_i[4065] & sel_one_hot_i[31];
  assign data_masked[4064] = data_i[4064] & sel_one_hot_i[31];
  assign data_masked[4063] = data_i[4063] & sel_one_hot_i[31];
  assign data_masked[4062] = data_i[4062] & sel_one_hot_i[31];
  assign data_masked[4061] = data_i[4061] & sel_one_hot_i[31];
  assign data_masked[4060] = data_i[4060] & sel_one_hot_i[31];
  assign data_masked[4059] = data_i[4059] & sel_one_hot_i[31];
  assign data_masked[4058] = data_i[4058] & sel_one_hot_i[31];
  assign data_masked[4057] = data_i[4057] & sel_one_hot_i[31];
  assign data_masked[4056] = data_i[4056] & sel_one_hot_i[31];
  assign data_masked[4055] = data_i[4055] & sel_one_hot_i[31];
  assign data_masked[4054] = data_i[4054] & sel_one_hot_i[31];
  assign data_masked[4053] = data_i[4053] & sel_one_hot_i[31];
  assign data_masked[4052] = data_i[4052] & sel_one_hot_i[31];
  assign data_masked[4051] = data_i[4051] & sel_one_hot_i[31];
  assign data_masked[4050] = data_i[4050] & sel_one_hot_i[31];
  assign data_masked[4049] = data_i[4049] & sel_one_hot_i[31];
  assign data_masked[4048] = data_i[4048] & sel_one_hot_i[31];
  assign data_masked[4047] = data_i[4047] & sel_one_hot_i[31];
  assign data_masked[4046] = data_i[4046] & sel_one_hot_i[31];
  assign data_masked[4045] = data_i[4045] & sel_one_hot_i[31];
  assign data_masked[4044] = data_i[4044] & sel_one_hot_i[31];
  assign data_masked[4043] = data_i[4043] & sel_one_hot_i[31];
  assign data_masked[4042] = data_i[4042] & sel_one_hot_i[31];
  assign data_masked[4041] = data_i[4041] & sel_one_hot_i[31];
  assign data_masked[4040] = data_i[4040] & sel_one_hot_i[31];
  assign data_masked[4039] = data_i[4039] & sel_one_hot_i[31];
  assign data_masked[4038] = data_i[4038] & sel_one_hot_i[31];
  assign data_masked[4037] = data_i[4037] & sel_one_hot_i[31];
  assign data_masked[4036] = data_i[4036] & sel_one_hot_i[31];
  assign data_masked[4035] = data_i[4035] & sel_one_hot_i[31];
  assign data_masked[4034] = data_i[4034] & sel_one_hot_i[31];
  assign data_masked[4033] = data_i[4033] & sel_one_hot_i[31];
  assign data_masked[4032] = data_i[4032] & sel_one_hot_i[31];
  assign data_masked[4031] = data_i[4031] & sel_one_hot_i[31];
  assign data_masked[4030] = data_i[4030] & sel_one_hot_i[31];
  assign data_masked[4029] = data_i[4029] & sel_one_hot_i[31];
  assign data_masked[4028] = data_i[4028] & sel_one_hot_i[31];
  assign data_masked[4027] = data_i[4027] & sel_one_hot_i[31];
  assign data_masked[4026] = data_i[4026] & sel_one_hot_i[31];
  assign data_masked[4025] = data_i[4025] & sel_one_hot_i[31];
  assign data_masked[4024] = data_i[4024] & sel_one_hot_i[31];
  assign data_masked[4023] = data_i[4023] & sel_one_hot_i[31];
  assign data_masked[4022] = data_i[4022] & sel_one_hot_i[31];
  assign data_masked[4021] = data_i[4021] & sel_one_hot_i[31];
  assign data_masked[4020] = data_i[4020] & sel_one_hot_i[31];
  assign data_masked[4019] = data_i[4019] & sel_one_hot_i[31];
  assign data_masked[4018] = data_i[4018] & sel_one_hot_i[31];
  assign data_masked[4017] = data_i[4017] & sel_one_hot_i[31];
  assign data_masked[4016] = data_i[4016] & sel_one_hot_i[31];
  assign data_masked[4015] = data_i[4015] & sel_one_hot_i[31];
  assign data_masked[4014] = data_i[4014] & sel_one_hot_i[31];
  assign data_masked[4013] = data_i[4013] & sel_one_hot_i[31];
  assign data_masked[4012] = data_i[4012] & sel_one_hot_i[31];
  assign data_masked[4011] = data_i[4011] & sel_one_hot_i[31];
  assign data_masked[4010] = data_i[4010] & sel_one_hot_i[31];
  assign data_masked[4009] = data_i[4009] & sel_one_hot_i[31];
  assign data_masked[4008] = data_i[4008] & sel_one_hot_i[31];
  assign data_masked[4007] = data_i[4007] & sel_one_hot_i[31];
  assign data_masked[4006] = data_i[4006] & sel_one_hot_i[31];
  assign data_masked[4005] = data_i[4005] & sel_one_hot_i[31];
  assign data_masked[4004] = data_i[4004] & sel_one_hot_i[31];
  assign data_masked[4003] = data_i[4003] & sel_one_hot_i[31];
  assign data_masked[4002] = data_i[4002] & sel_one_hot_i[31];
  assign data_masked[4001] = data_i[4001] & sel_one_hot_i[31];
  assign data_masked[4000] = data_i[4000] & sel_one_hot_i[31];
  assign data_masked[3999] = data_i[3999] & sel_one_hot_i[31];
  assign data_masked[3998] = data_i[3998] & sel_one_hot_i[31];
  assign data_masked[3997] = data_i[3997] & sel_one_hot_i[31];
  assign data_masked[3996] = data_i[3996] & sel_one_hot_i[31];
  assign data_masked[3995] = data_i[3995] & sel_one_hot_i[31];
  assign data_masked[3994] = data_i[3994] & sel_one_hot_i[31];
  assign data_masked[3993] = data_i[3993] & sel_one_hot_i[31];
  assign data_masked[3992] = data_i[3992] & sel_one_hot_i[31];
  assign data_masked[3991] = data_i[3991] & sel_one_hot_i[31];
  assign data_masked[3990] = data_i[3990] & sel_one_hot_i[31];
  assign data_masked[3989] = data_i[3989] & sel_one_hot_i[31];
  assign data_masked[3988] = data_i[3988] & sel_one_hot_i[31];
  assign data_masked[3987] = data_i[3987] & sel_one_hot_i[31];
  assign data_masked[3986] = data_i[3986] & sel_one_hot_i[31];
  assign data_masked[3985] = data_i[3985] & sel_one_hot_i[31];
  assign data_masked[3984] = data_i[3984] & sel_one_hot_i[31];
  assign data_masked[3983] = data_i[3983] & sel_one_hot_i[31];
  assign data_masked[3982] = data_i[3982] & sel_one_hot_i[31];
  assign data_masked[3981] = data_i[3981] & sel_one_hot_i[31];
  assign data_masked[3980] = data_i[3980] & sel_one_hot_i[31];
  assign data_masked[3979] = data_i[3979] & sel_one_hot_i[31];
  assign data_masked[3978] = data_i[3978] & sel_one_hot_i[31];
  assign data_masked[3977] = data_i[3977] & sel_one_hot_i[31];
  assign data_masked[3976] = data_i[3976] & sel_one_hot_i[31];
  assign data_masked[3975] = data_i[3975] & sel_one_hot_i[31];
  assign data_masked[3974] = data_i[3974] & sel_one_hot_i[31];
  assign data_masked[3973] = data_i[3973] & sel_one_hot_i[31];
  assign data_masked[3972] = data_i[3972] & sel_one_hot_i[31];
  assign data_masked[3971] = data_i[3971] & sel_one_hot_i[31];
  assign data_masked[3970] = data_i[3970] & sel_one_hot_i[31];
  assign data_masked[3969] = data_i[3969] & sel_one_hot_i[31];
  assign data_masked[3968] = data_i[3968] & sel_one_hot_i[31];
  assign data_masked[4223] = data_i[4223] & sel_one_hot_i[32];
  assign data_masked[4222] = data_i[4222] & sel_one_hot_i[32];
  assign data_masked[4221] = data_i[4221] & sel_one_hot_i[32];
  assign data_masked[4220] = data_i[4220] & sel_one_hot_i[32];
  assign data_masked[4219] = data_i[4219] & sel_one_hot_i[32];
  assign data_masked[4218] = data_i[4218] & sel_one_hot_i[32];
  assign data_masked[4217] = data_i[4217] & sel_one_hot_i[32];
  assign data_masked[4216] = data_i[4216] & sel_one_hot_i[32];
  assign data_masked[4215] = data_i[4215] & sel_one_hot_i[32];
  assign data_masked[4214] = data_i[4214] & sel_one_hot_i[32];
  assign data_masked[4213] = data_i[4213] & sel_one_hot_i[32];
  assign data_masked[4212] = data_i[4212] & sel_one_hot_i[32];
  assign data_masked[4211] = data_i[4211] & sel_one_hot_i[32];
  assign data_masked[4210] = data_i[4210] & sel_one_hot_i[32];
  assign data_masked[4209] = data_i[4209] & sel_one_hot_i[32];
  assign data_masked[4208] = data_i[4208] & sel_one_hot_i[32];
  assign data_masked[4207] = data_i[4207] & sel_one_hot_i[32];
  assign data_masked[4206] = data_i[4206] & sel_one_hot_i[32];
  assign data_masked[4205] = data_i[4205] & sel_one_hot_i[32];
  assign data_masked[4204] = data_i[4204] & sel_one_hot_i[32];
  assign data_masked[4203] = data_i[4203] & sel_one_hot_i[32];
  assign data_masked[4202] = data_i[4202] & sel_one_hot_i[32];
  assign data_masked[4201] = data_i[4201] & sel_one_hot_i[32];
  assign data_masked[4200] = data_i[4200] & sel_one_hot_i[32];
  assign data_masked[4199] = data_i[4199] & sel_one_hot_i[32];
  assign data_masked[4198] = data_i[4198] & sel_one_hot_i[32];
  assign data_masked[4197] = data_i[4197] & sel_one_hot_i[32];
  assign data_masked[4196] = data_i[4196] & sel_one_hot_i[32];
  assign data_masked[4195] = data_i[4195] & sel_one_hot_i[32];
  assign data_masked[4194] = data_i[4194] & sel_one_hot_i[32];
  assign data_masked[4193] = data_i[4193] & sel_one_hot_i[32];
  assign data_masked[4192] = data_i[4192] & sel_one_hot_i[32];
  assign data_masked[4191] = data_i[4191] & sel_one_hot_i[32];
  assign data_masked[4190] = data_i[4190] & sel_one_hot_i[32];
  assign data_masked[4189] = data_i[4189] & sel_one_hot_i[32];
  assign data_masked[4188] = data_i[4188] & sel_one_hot_i[32];
  assign data_masked[4187] = data_i[4187] & sel_one_hot_i[32];
  assign data_masked[4186] = data_i[4186] & sel_one_hot_i[32];
  assign data_masked[4185] = data_i[4185] & sel_one_hot_i[32];
  assign data_masked[4184] = data_i[4184] & sel_one_hot_i[32];
  assign data_masked[4183] = data_i[4183] & sel_one_hot_i[32];
  assign data_masked[4182] = data_i[4182] & sel_one_hot_i[32];
  assign data_masked[4181] = data_i[4181] & sel_one_hot_i[32];
  assign data_masked[4180] = data_i[4180] & sel_one_hot_i[32];
  assign data_masked[4179] = data_i[4179] & sel_one_hot_i[32];
  assign data_masked[4178] = data_i[4178] & sel_one_hot_i[32];
  assign data_masked[4177] = data_i[4177] & sel_one_hot_i[32];
  assign data_masked[4176] = data_i[4176] & sel_one_hot_i[32];
  assign data_masked[4175] = data_i[4175] & sel_one_hot_i[32];
  assign data_masked[4174] = data_i[4174] & sel_one_hot_i[32];
  assign data_masked[4173] = data_i[4173] & sel_one_hot_i[32];
  assign data_masked[4172] = data_i[4172] & sel_one_hot_i[32];
  assign data_masked[4171] = data_i[4171] & sel_one_hot_i[32];
  assign data_masked[4170] = data_i[4170] & sel_one_hot_i[32];
  assign data_masked[4169] = data_i[4169] & sel_one_hot_i[32];
  assign data_masked[4168] = data_i[4168] & sel_one_hot_i[32];
  assign data_masked[4167] = data_i[4167] & sel_one_hot_i[32];
  assign data_masked[4166] = data_i[4166] & sel_one_hot_i[32];
  assign data_masked[4165] = data_i[4165] & sel_one_hot_i[32];
  assign data_masked[4164] = data_i[4164] & sel_one_hot_i[32];
  assign data_masked[4163] = data_i[4163] & sel_one_hot_i[32];
  assign data_masked[4162] = data_i[4162] & sel_one_hot_i[32];
  assign data_masked[4161] = data_i[4161] & sel_one_hot_i[32];
  assign data_masked[4160] = data_i[4160] & sel_one_hot_i[32];
  assign data_masked[4159] = data_i[4159] & sel_one_hot_i[32];
  assign data_masked[4158] = data_i[4158] & sel_one_hot_i[32];
  assign data_masked[4157] = data_i[4157] & sel_one_hot_i[32];
  assign data_masked[4156] = data_i[4156] & sel_one_hot_i[32];
  assign data_masked[4155] = data_i[4155] & sel_one_hot_i[32];
  assign data_masked[4154] = data_i[4154] & sel_one_hot_i[32];
  assign data_masked[4153] = data_i[4153] & sel_one_hot_i[32];
  assign data_masked[4152] = data_i[4152] & sel_one_hot_i[32];
  assign data_masked[4151] = data_i[4151] & sel_one_hot_i[32];
  assign data_masked[4150] = data_i[4150] & sel_one_hot_i[32];
  assign data_masked[4149] = data_i[4149] & sel_one_hot_i[32];
  assign data_masked[4148] = data_i[4148] & sel_one_hot_i[32];
  assign data_masked[4147] = data_i[4147] & sel_one_hot_i[32];
  assign data_masked[4146] = data_i[4146] & sel_one_hot_i[32];
  assign data_masked[4145] = data_i[4145] & sel_one_hot_i[32];
  assign data_masked[4144] = data_i[4144] & sel_one_hot_i[32];
  assign data_masked[4143] = data_i[4143] & sel_one_hot_i[32];
  assign data_masked[4142] = data_i[4142] & sel_one_hot_i[32];
  assign data_masked[4141] = data_i[4141] & sel_one_hot_i[32];
  assign data_masked[4140] = data_i[4140] & sel_one_hot_i[32];
  assign data_masked[4139] = data_i[4139] & sel_one_hot_i[32];
  assign data_masked[4138] = data_i[4138] & sel_one_hot_i[32];
  assign data_masked[4137] = data_i[4137] & sel_one_hot_i[32];
  assign data_masked[4136] = data_i[4136] & sel_one_hot_i[32];
  assign data_masked[4135] = data_i[4135] & sel_one_hot_i[32];
  assign data_masked[4134] = data_i[4134] & sel_one_hot_i[32];
  assign data_masked[4133] = data_i[4133] & sel_one_hot_i[32];
  assign data_masked[4132] = data_i[4132] & sel_one_hot_i[32];
  assign data_masked[4131] = data_i[4131] & sel_one_hot_i[32];
  assign data_masked[4130] = data_i[4130] & sel_one_hot_i[32];
  assign data_masked[4129] = data_i[4129] & sel_one_hot_i[32];
  assign data_masked[4128] = data_i[4128] & sel_one_hot_i[32];
  assign data_masked[4127] = data_i[4127] & sel_one_hot_i[32];
  assign data_masked[4126] = data_i[4126] & sel_one_hot_i[32];
  assign data_masked[4125] = data_i[4125] & sel_one_hot_i[32];
  assign data_masked[4124] = data_i[4124] & sel_one_hot_i[32];
  assign data_masked[4123] = data_i[4123] & sel_one_hot_i[32];
  assign data_masked[4122] = data_i[4122] & sel_one_hot_i[32];
  assign data_masked[4121] = data_i[4121] & sel_one_hot_i[32];
  assign data_masked[4120] = data_i[4120] & sel_one_hot_i[32];
  assign data_masked[4119] = data_i[4119] & sel_one_hot_i[32];
  assign data_masked[4118] = data_i[4118] & sel_one_hot_i[32];
  assign data_masked[4117] = data_i[4117] & sel_one_hot_i[32];
  assign data_masked[4116] = data_i[4116] & sel_one_hot_i[32];
  assign data_masked[4115] = data_i[4115] & sel_one_hot_i[32];
  assign data_masked[4114] = data_i[4114] & sel_one_hot_i[32];
  assign data_masked[4113] = data_i[4113] & sel_one_hot_i[32];
  assign data_masked[4112] = data_i[4112] & sel_one_hot_i[32];
  assign data_masked[4111] = data_i[4111] & sel_one_hot_i[32];
  assign data_masked[4110] = data_i[4110] & sel_one_hot_i[32];
  assign data_masked[4109] = data_i[4109] & sel_one_hot_i[32];
  assign data_masked[4108] = data_i[4108] & sel_one_hot_i[32];
  assign data_masked[4107] = data_i[4107] & sel_one_hot_i[32];
  assign data_masked[4106] = data_i[4106] & sel_one_hot_i[32];
  assign data_masked[4105] = data_i[4105] & sel_one_hot_i[32];
  assign data_masked[4104] = data_i[4104] & sel_one_hot_i[32];
  assign data_masked[4103] = data_i[4103] & sel_one_hot_i[32];
  assign data_masked[4102] = data_i[4102] & sel_one_hot_i[32];
  assign data_masked[4101] = data_i[4101] & sel_one_hot_i[32];
  assign data_masked[4100] = data_i[4100] & sel_one_hot_i[32];
  assign data_masked[4099] = data_i[4099] & sel_one_hot_i[32];
  assign data_masked[4098] = data_i[4098] & sel_one_hot_i[32];
  assign data_masked[4097] = data_i[4097] & sel_one_hot_i[32];
  assign data_masked[4096] = data_i[4096] & sel_one_hot_i[32];
  assign data_masked[4351] = data_i[4351] & sel_one_hot_i[33];
  assign data_masked[4350] = data_i[4350] & sel_one_hot_i[33];
  assign data_masked[4349] = data_i[4349] & sel_one_hot_i[33];
  assign data_masked[4348] = data_i[4348] & sel_one_hot_i[33];
  assign data_masked[4347] = data_i[4347] & sel_one_hot_i[33];
  assign data_masked[4346] = data_i[4346] & sel_one_hot_i[33];
  assign data_masked[4345] = data_i[4345] & sel_one_hot_i[33];
  assign data_masked[4344] = data_i[4344] & sel_one_hot_i[33];
  assign data_masked[4343] = data_i[4343] & sel_one_hot_i[33];
  assign data_masked[4342] = data_i[4342] & sel_one_hot_i[33];
  assign data_masked[4341] = data_i[4341] & sel_one_hot_i[33];
  assign data_masked[4340] = data_i[4340] & sel_one_hot_i[33];
  assign data_masked[4339] = data_i[4339] & sel_one_hot_i[33];
  assign data_masked[4338] = data_i[4338] & sel_one_hot_i[33];
  assign data_masked[4337] = data_i[4337] & sel_one_hot_i[33];
  assign data_masked[4336] = data_i[4336] & sel_one_hot_i[33];
  assign data_masked[4335] = data_i[4335] & sel_one_hot_i[33];
  assign data_masked[4334] = data_i[4334] & sel_one_hot_i[33];
  assign data_masked[4333] = data_i[4333] & sel_one_hot_i[33];
  assign data_masked[4332] = data_i[4332] & sel_one_hot_i[33];
  assign data_masked[4331] = data_i[4331] & sel_one_hot_i[33];
  assign data_masked[4330] = data_i[4330] & sel_one_hot_i[33];
  assign data_masked[4329] = data_i[4329] & sel_one_hot_i[33];
  assign data_masked[4328] = data_i[4328] & sel_one_hot_i[33];
  assign data_masked[4327] = data_i[4327] & sel_one_hot_i[33];
  assign data_masked[4326] = data_i[4326] & sel_one_hot_i[33];
  assign data_masked[4325] = data_i[4325] & sel_one_hot_i[33];
  assign data_masked[4324] = data_i[4324] & sel_one_hot_i[33];
  assign data_masked[4323] = data_i[4323] & sel_one_hot_i[33];
  assign data_masked[4322] = data_i[4322] & sel_one_hot_i[33];
  assign data_masked[4321] = data_i[4321] & sel_one_hot_i[33];
  assign data_masked[4320] = data_i[4320] & sel_one_hot_i[33];
  assign data_masked[4319] = data_i[4319] & sel_one_hot_i[33];
  assign data_masked[4318] = data_i[4318] & sel_one_hot_i[33];
  assign data_masked[4317] = data_i[4317] & sel_one_hot_i[33];
  assign data_masked[4316] = data_i[4316] & sel_one_hot_i[33];
  assign data_masked[4315] = data_i[4315] & sel_one_hot_i[33];
  assign data_masked[4314] = data_i[4314] & sel_one_hot_i[33];
  assign data_masked[4313] = data_i[4313] & sel_one_hot_i[33];
  assign data_masked[4312] = data_i[4312] & sel_one_hot_i[33];
  assign data_masked[4311] = data_i[4311] & sel_one_hot_i[33];
  assign data_masked[4310] = data_i[4310] & sel_one_hot_i[33];
  assign data_masked[4309] = data_i[4309] & sel_one_hot_i[33];
  assign data_masked[4308] = data_i[4308] & sel_one_hot_i[33];
  assign data_masked[4307] = data_i[4307] & sel_one_hot_i[33];
  assign data_masked[4306] = data_i[4306] & sel_one_hot_i[33];
  assign data_masked[4305] = data_i[4305] & sel_one_hot_i[33];
  assign data_masked[4304] = data_i[4304] & sel_one_hot_i[33];
  assign data_masked[4303] = data_i[4303] & sel_one_hot_i[33];
  assign data_masked[4302] = data_i[4302] & sel_one_hot_i[33];
  assign data_masked[4301] = data_i[4301] & sel_one_hot_i[33];
  assign data_masked[4300] = data_i[4300] & sel_one_hot_i[33];
  assign data_masked[4299] = data_i[4299] & sel_one_hot_i[33];
  assign data_masked[4298] = data_i[4298] & sel_one_hot_i[33];
  assign data_masked[4297] = data_i[4297] & sel_one_hot_i[33];
  assign data_masked[4296] = data_i[4296] & sel_one_hot_i[33];
  assign data_masked[4295] = data_i[4295] & sel_one_hot_i[33];
  assign data_masked[4294] = data_i[4294] & sel_one_hot_i[33];
  assign data_masked[4293] = data_i[4293] & sel_one_hot_i[33];
  assign data_masked[4292] = data_i[4292] & sel_one_hot_i[33];
  assign data_masked[4291] = data_i[4291] & sel_one_hot_i[33];
  assign data_masked[4290] = data_i[4290] & sel_one_hot_i[33];
  assign data_masked[4289] = data_i[4289] & sel_one_hot_i[33];
  assign data_masked[4288] = data_i[4288] & sel_one_hot_i[33];
  assign data_masked[4287] = data_i[4287] & sel_one_hot_i[33];
  assign data_masked[4286] = data_i[4286] & sel_one_hot_i[33];
  assign data_masked[4285] = data_i[4285] & sel_one_hot_i[33];
  assign data_masked[4284] = data_i[4284] & sel_one_hot_i[33];
  assign data_masked[4283] = data_i[4283] & sel_one_hot_i[33];
  assign data_masked[4282] = data_i[4282] & sel_one_hot_i[33];
  assign data_masked[4281] = data_i[4281] & sel_one_hot_i[33];
  assign data_masked[4280] = data_i[4280] & sel_one_hot_i[33];
  assign data_masked[4279] = data_i[4279] & sel_one_hot_i[33];
  assign data_masked[4278] = data_i[4278] & sel_one_hot_i[33];
  assign data_masked[4277] = data_i[4277] & sel_one_hot_i[33];
  assign data_masked[4276] = data_i[4276] & sel_one_hot_i[33];
  assign data_masked[4275] = data_i[4275] & sel_one_hot_i[33];
  assign data_masked[4274] = data_i[4274] & sel_one_hot_i[33];
  assign data_masked[4273] = data_i[4273] & sel_one_hot_i[33];
  assign data_masked[4272] = data_i[4272] & sel_one_hot_i[33];
  assign data_masked[4271] = data_i[4271] & sel_one_hot_i[33];
  assign data_masked[4270] = data_i[4270] & sel_one_hot_i[33];
  assign data_masked[4269] = data_i[4269] & sel_one_hot_i[33];
  assign data_masked[4268] = data_i[4268] & sel_one_hot_i[33];
  assign data_masked[4267] = data_i[4267] & sel_one_hot_i[33];
  assign data_masked[4266] = data_i[4266] & sel_one_hot_i[33];
  assign data_masked[4265] = data_i[4265] & sel_one_hot_i[33];
  assign data_masked[4264] = data_i[4264] & sel_one_hot_i[33];
  assign data_masked[4263] = data_i[4263] & sel_one_hot_i[33];
  assign data_masked[4262] = data_i[4262] & sel_one_hot_i[33];
  assign data_masked[4261] = data_i[4261] & sel_one_hot_i[33];
  assign data_masked[4260] = data_i[4260] & sel_one_hot_i[33];
  assign data_masked[4259] = data_i[4259] & sel_one_hot_i[33];
  assign data_masked[4258] = data_i[4258] & sel_one_hot_i[33];
  assign data_masked[4257] = data_i[4257] & sel_one_hot_i[33];
  assign data_masked[4256] = data_i[4256] & sel_one_hot_i[33];
  assign data_masked[4255] = data_i[4255] & sel_one_hot_i[33];
  assign data_masked[4254] = data_i[4254] & sel_one_hot_i[33];
  assign data_masked[4253] = data_i[4253] & sel_one_hot_i[33];
  assign data_masked[4252] = data_i[4252] & sel_one_hot_i[33];
  assign data_masked[4251] = data_i[4251] & sel_one_hot_i[33];
  assign data_masked[4250] = data_i[4250] & sel_one_hot_i[33];
  assign data_masked[4249] = data_i[4249] & sel_one_hot_i[33];
  assign data_masked[4248] = data_i[4248] & sel_one_hot_i[33];
  assign data_masked[4247] = data_i[4247] & sel_one_hot_i[33];
  assign data_masked[4246] = data_i[4246] & sel_one_hot_i[33];
  assign data_masked[4245] = data_i[4245] & sel_one_hot_i[33];
  assign data_masked[4244] = data_i[4244] & sel_one_hot_i[33];
  assign data_masked[4243] = data_i[4243] & sel_one_hot_i[33];
  assign data_masked[4242] = data_i[4242] & sel_one_hot_i[33];
  assign data_masked[4241] = data_i[4241] & sel_one_hot_i[33];
  assign data_masked[4240] = data_i[4240] & sel_one_hot_i[33];
  assign data_masked[4239] = data_i[4239] & sel_one_hot_i[33];
  assign data_masked[4238] = data_i[4238] & sel_one_hot_i[33];
  assign data_masked[4237] = data_i[4237] & sel_one_hot_i[33];
  assign data_masked[4236] = data_i[4236] & sel_one_hot_i[33];
  assign data_masked[4235] = data_i[4235] & sel_one_hot_i[33];
  assign data_masked[4234] = data_i[4234] & sel_one_hot_i[33];
  assign data_masked[4233] = data_i[4233] & sel_one_hot_i[33];
  assign data_masked[4232] = data_i[4232] & sel_one_hot_i[33];
  assign data_masked[4231] = data_i[4231] & sel_one_hot_i[33];
  assign data_masked[4230] = data_i[4230] & sel_one_hot_i[33];
  assign data_masked[4229] = data_i[4229] & sel_one_hot_i[33];
  assign data_masked[4228] = data_i[4228] & sel_one_hot_i[33];
  assign data_masked[4227] = data_i[4227] & sel_one_hot_i[33];
  assign data_masked[4226] = data_i[4226] & sel_one_hot_i[33];
  assign data_masked[4225] = data_i[4225] & sel_one_hot_i[33];
  assign data_masked[4224] = data_i[4224] & sel_one_hot_i[33];
  assign data_masked[4479] = data_i[4479] & sel_one_hot_i[34];
  assign data_masked[4478] = data_i[4478] & sel_one_hot_i[34];
  assign data_masked[4477] = data_i[4477] & sel_one_hot_i[34];
  assign data_masked[4476] = data_i[4476] & sel_one_hot_i[34];
  assign data_masked[4475] = data_i[4475] & sel_one_hot_i[34];
  assign data_masked[4474] = data_i[4474] & sel_one_hot_i[34];
  assign data_masked[4473] = data_i[4473] & sel_one_hot_i[34];
  assign data_masked[4472] = data_i[4472] & sel_one_hot_i[34];
  assign data_masked[4471] = data_i[4471] & sel_one_hot_i[34];
  assign data_masked[4470] = data_i[4470] & sel_one_hot_i[34];
  assign data_masked[4469] = data_i[4469] & sel_one_hot_i[34];
  assign data_masked[4468] = data_i[4468] & sel_one_hot_i[34];
  assign data_masked[4467] = data_i[4467] & sel_one_hot_i[34];
  assign data_masked[4466] = data_i[4466] & sel_one_hot_i[34];
  assign data_masked[4465] = data_i[4465] & sel_one_hot_i[34];
  assign data_masked[4464] = data_i[4464] & sel_one_hot_i[34];
  assign data_masked[4463] = data_i[4463] & sel_one_hot_i[34];
  assign data_masked[4462] = data_i[4462] & sel_one_hot_i[34];
  assign data_masked[4461] = data_i[4461] & sel_one_hot_i[34];
  assign data_masked[4460] = data_i[4460] & sel_one_hot_i[34];
  assign data_masked[4459] = data_i[4459] & sel_one_hot_i[34];
  assign data_masked[4458] = data_i[4458] & sel_one_hot_i[34];
  assign data_masked[4457] = data_i[4457] & sel_one_hot_i[34];
  assign data_masked[4456] = data_i[4456] & sel_one_hot_i[34];
  assign data_masked[4455] = data_i[4455] & sel_one_hot_i[34];
  assign data_masked[4454] = data_i[4454] & sel_one_hot_i[34];
  assign data_masked[4453] = data_i[4453] & sel_one_hot_i[34];
  assign data_masked[4452] = data_i[4452] & sel_one_hot_i[34];
  assign data_masked[4451] = data_i[4451] & sel_one_hot_i[34];
  assign data_masked[4450] = data_i[4450] & sel_one_hot_i[34];
  assign data_masked[4449] = data_i[4449] & sel_one_hot_i[34];
  assign data_masked[4448] = data_i[4448] & sel_one_hot_i[34];
  assign data_masked[4447] = data_i[4447] & sel_one_hot_i[34];
  assign data_masked[4446] = data_i[4446] & sel_one_hot_i[34];
  assign data_masked[4445] = data_i[4445] & sel_one_hot_i[34];
  assign data_masked[4444] = data_i[4444] & sel_one_hot_i[34];
  assign data_masked[4443] = data_i[4443] & sel_one_hot_i[34];
  assign data_masked[4442] = data_i[4442] & sel_one_hot_i[34];
  assign data_masked[4441] = data_i[4441] & sel_one_hot_i[34];
  assign data_masked[4440] = data_i[4440] & sel_one_hot_i[34];
  assign data_masked[4439] = data_i[4439] & sel_one_hot_i[34];
  assign data_masked[4438] = data_i[4438] & sel_one_hot_i[34];
  assign data_masked[4437] = data_i[4437] & sel_one_hot_i[34];
  assign data_masked[4436] = data_i[4436] & sel_one_hot_i[34];
  assign data_masked[4435] = data_i[4435] & sel_one_hot_i[34];
  assign data_masked[4434] = data_i[4434] & sel_one_hot_i[34];
  assign data_masked[4433] = data_i[4433] & sel_one_hot_i[34];
  assign data_masked[4432] = data_i[4432] & sel_one_hot_i[34];
  assign data_masked[4431] = data_i[4431] & sel_one_hot_i[34];
  assign data_masked[4430] = data_i[4430] & sel_one_hot_i[34];
  assign data_masked[4429] = data_i[4429] & sel_one_hot_i[34];
  assign data_masked[4428] = data_i[4428] & sel_one_hot_i[34];
  assign data_masked[4427] = data_i[4427] & sel_one_hot_i[34];
  assign data_masked[4426] = data_i[4426] & sel_one_hot_i[34];
  assign data_masked[4425] = data_i[4425] & sel_one_hot_i[34];
  assign data_masked[4424] = data_i[4424] & sel_one_hot_i[34];
  assign data_masked[4423] = data_i[4423] & sel_one_hot_i[34];
  assign data_masked[4422] = data_i[4422] & sel_one_hot_i[34];
  assign data_masked[4421] = data_i[4421] & sel_one_hot_i[34];
  assign data_masked[4420] = data_i[4420] & sel_one_hot_i[34];
  assign data_masked[4419] = data_i[4419] & sel_one_hot_i[34];
  assign data_masked[4418] = data_i[4418] & sel_one_hot_i[34];
  assign data_masked[4417] = data_i[4417] & sel_one_hot_i[34];
  assign data_masked[4416] = data_i[4416] & sel_one_hot_i[34];
  assign data_masked[4415] = data_i[4415] & sel_one_hot_i[34];
  assign data_masked[4414] = data_i[4414] & sel_one_hot_i[34];
  assign data_masked[4413] = data_i[4413] & sel_one_hot_i[34];
  assign data_masked[4412] = data_i[4412] & sel_one_hot_i[34];
  assign data_masked[4411] = data_i[4411] & sel_one_hot_i[34];
  assign data_masked[4410] = data_i[4410] & sel_one_hot_i[34];
  assign data_masked[4409] = data_i[4409] & sel_one_hot_i[34];
  assign data_masked[4408] = data_i[4408] & sel_one_hot_i[34];
  assign data_masked[4407] = data_i[4407] & sel_one_hot_i[34];
  assign data_masked[4406] = data_i[4406] & sel_one_hot_i[34];
  assign data_masked[4405] = data_i[4405] & sel_one_hot_i[34];
  assign data_masked[4404] = data_i[4404] & sel_one_hot_i[34];
  assign data_masked[4403] = data_i[4403] & sel_one_hot_i[34];
  assign data_masked[4402] = data_i[4402] & sel_one_hot_i[34];
  assign data_masked[4401] = data_i[4401] & sel_one_hot_i[34];
  assign data_masked[4400] = data_i[4400] & sel_one_hot_i[34];
  assign data_masked[4399] = data_i[4399] & sel_one_hot_i[34];
  assign data_masked[4398] = data_i[4398] & sel_one_hot_i[34];
  assign data_masked[4397] = data_i[4397] & sel_one_hot_i[34];
  assign data_masked[4396] = data_i[4396] & sel_one_hot_i[34];
  assign data_masked[4395] = data_i[4395] & sel_one_hot_i[34];
  assign data_masked[4394] = data_i[4394] & sel_one_hot_i[34];
  assign data_masked[4393] = data_i[4393] & sel_one_hot_i[34];
  assign data_masked[4392] = data_i[4392] & sel_one_hot_i[34];
  assign data_masked[4391] = data_i[4391] & sel_one_hot_i[34];
  assign data_masked[4390] = data_i[4390] & sel_one_hot_i[34];
  assign data_masked[4389] = data_i[4389] & sel_one_hot_i[34];
  assign data_masked[4388] = data_i[4388] & sel_one_hot_i[34];
  assign data_masked[4387] = data_i[4387] & sel_one_hot_i[34];
  assign data_masked[4386] = data_i[4386] & sel_one_hot_i[34];
  assign data_masked[4385] = data_i[4385] & sel_one_hot_i[34];
  assign data_masked[4384] = data_i[4384] & sel_one_hot_i[34];
  assign data_masked[4383] = data_i[4383] & sel_one_hot_i[34];
  assign data_masked[4382] = data_i[4382] & sel_one_hot_i[34];
  assign data_masked[4381] = data_i[4381] & sel_one_hot_i[34];
  assign data_masked[4380] = data_i[4380] & sel_one_hot_i[34];
  assign data_masked[4379] = data_i[4379] & sel_one_hot_i[34];
  assign data_masked[4378] = data_i[4378] & sel_one_hot_i[34];
  assign data_masked[4377] = data_i[4377] & sel_one_hot_i[34];
  assign data_masked[4376] = data_i[4376] & sel_one_hot_i[34];
  assign data_masked[4375] = data_i[4375] & sel_one_hot_i[34];
  assign data_masked[4374] = data_i[4374] & sel_one_hot_i[34];
  assign data_masked[4373] = data_i[4373] & sel_one_hot_i[34];
  assign data_masked[4372] = data_i[4372] & sel_one_hot_i[34];
  assign data_masked[4371] = data_i[4371] & sel_one_hot_i[34];
  assign data_masked[4370] = data_i[4370] & sel_one_hot_i[34];
  assign data_masked[4369] = data_i[4369] & sel_one_hot_i[34];
  assign data_masked[4368] = data_i[4368] & sel_one_hot_i[34];
  assign data_masked[4367] = data_i[4367] & sel_one_hot_i[34];
  assign data_masked[4366] = data_i[4366] & sel_one_hot_i[34];
  assign data_masked[4365] = data_i[4365] & sel_one_hot_i[34];
  assign data_masked[4364] = data_i[4364] & sel_one_hot_i[34];
  assign data_masked[4363] = data_i[4363] & sel_one_hot_i[34];
  assign data_masked[4362] = data_i[4362] & sel_one_hot_i[34];
  assign data_masked[4361] = data_i[4361] & sel_one_hot_i[34];
  assign data_masked[4360] = data_i[4360] & sel_one_hot_i[34];
  assign data_masked[4359] = data_i[4359] & sel_one_hot_i[34];
  assign data_masked[4358] = data_i[4358] & sel_one_hot_i[34];
  assign data_masked[4357] = data_i[4357] & sel_one_hot_i[34];
  assign data_masked[4356] = data_i[4356] & sel_one_hot_i[34];
  assign data_masked[4355] = data_i[4355] & sel_one_hot_i[34];
  assign data_masked[4354] = data_i[4354] & sel_one_hot_i[34];
  assign data_masked[4353] = data_i[4353] & sel_one_hot_i[34];
  assign data_masked[4352] = data_i[4352] & sel_one_hot_i[34];
  assign data_masked[4607] = data_i[4607] & sel_one_hot_i[35];
  assign data_masked[4606] = data_i[4606] & sel_one_hot_i[35];
  assign data_masked[4605] = data_i[4605] & sel_one_hot_i[35];
  assign data_masked[4604] = data_i[4604] & sel_one_hot_i[35];
  assign data_masked[4603] = data_i[4603] & sel_one_hot_i[35];
  assign data_masked[4602] = data_i[4602] & sel_one_hot_i[35];
  assign data_masked[4601] = data_i[4601] & sel_one_hot_i[35];
  assign data_masked[4600] = data_i[4600] & sel_one_hot_i[35];
  assign data_masked[4599] = data_i[4599] & sel_one_hot_i[35];
  assign data_masked[4598] = data_i[4598] & sel_one_hot_i[35];
  assign data_masked[4597] = data_i[4597] & sel_one_hot_i[35];
  assign data_masked[4596] = data_i[4596] & sel_one_hot_i[35];
  assign data_masked[4595] = data_i[4595] & sel_one_hot_i[35];
  assign data_masked[4594] = data_i[4594] & sel_one_hot_i[35];
  assign data_masked[4593] = data_i[4593] & sel_one_hot_i[35];
  assign data_masked[4592] = data_i[4592] & sel_one_hot_i[35];
  assign data_masked[4591] = data_i[4591] & sel_one_hot_i[35];
  assign data_masked[4590] = data_i[4590] & sel_one_hot_i[35];
  assign data_masked[4589] = data_i[4589] & sel_one_hot_i[35];
  assign data_masked[4588] = data_i[4588] & sel_one_hot_i[35];
  assign data_masked[4587] = data_i[4587] & sel_one_hot_i[35];
  assign data_masked[4586] = data_i[4586] & sel_one_hot_i[35];
  assign data_masked[4585] = data_i[4585] & sel_one_hot_i[35];
  assign data_masked[4584] = data_i[4584] & sel_one_hot_i[35];
  assign data_masked[4583] = data_i[4583] & sel_one_hot_i[35];
  assign data_masked[4582] = data_i[4582] & sel_one_hot_i[35];
  assign data_masked[4581] = data_i[4581] & sel_one_hot_i[35];
  assign data_masked[4580] = data_i[4580] & sel_one_hot_i[35];
  assign data_masked[4579] = data_i[4579] & sel_one_hot_i[35];
  assign data_masked[4578] = data_i[4578] & sel_one_hot_i[35];
  assign data_masked[4577] = data_i[4577] & sel_one_hot_i[35];
  assign data_masked[4576] = data_i[4576] & sel_one_hot_i[35];
  assign data_masked[4575] = data_i[4575] & sel_one_hot_i[35];
  assign data_masked[4574] = data_i[4574] & sel_one_hot_i[35];
  assign data_masked[4573] = data_i[4573] & sel_one_hot_i[35];
  assign data_masked[4572] = data_i[4572] & sel_one_hot_i[35];
  assign data_masked[4571] = data_i[4571] & sel_one_hot_i[35];
  assign data_masked[4570] = data_i[4570] & sel_one_hot_i[35];
  assign data_masked[4569] = data_i[4569] & sel_one_hot_i[35];
  assign data_masked[4568] = data_i[4568] & sel_one_hot_i[35];
  assign data_masked[4567] = data_i[4567] & sel_one_hot_i[35];
  assign data_masked[4566] = data_i[4566] & sel_one_hot_i[35];
  assign data_masked[4565] = data_i[4565] & sel_one_hot_i[35];
  assign data_masked[4564] = data_i[4564] & sel_one_hot_i[35];
  assign data_masked[4563] = data_i[4563] & sel_one_hot_i[35];
  assign data_masked[4562] = data_i[4562] & sel_one_hot_i[35];
  assign data_masked[4561] = data_i[4561] & sel_one_hot_i[35];
  assign data_masked[4560] = data_i[4560] & sel_one_hot_i[35];
  assign data_masked[4559] = data_i[4559] & sel_one_hot_i[35];
  assign data_masked[4558] = data_i[4558] & sel_one_hot_i[35];
  assign data_masked[4557] = data_i[4557] & sel_one_hot_i[35];
  assign data_masked[4556] = data_i[4556] & sel_one_hot_i[35];
  assign data_masked[4555] = data_i[4555] & sel_one_hot_i[35];
  assign data_masked[4554] = data_i[4554] & sel_one_hot_i[35];
  assign data_masked[4553] = data_i[4553] & sel_one_hot_i[35];
  assign data_masked[4552] = data_i[4552] & sel_one_hot_i[35];
  assign data_masked[4551] = data_i[4551] & sel_one_hot_i[35];
  assign data_masked[4550] = data_i[4550] & sel_one_hot_i[35];
  assign data_masked[4549] = data_i[4549] & sel_one_hot_i[35];
  assign data_masked[4548] = data_i[4548] & sel_one_hot_i[35];
  assign data_masked[4547] = data_i[4547] & sel_one_hot_i[35];
  assign data_masked[4546] = data_i[4546] & sel_one_hot_i[35];
  assign data_masked[4545] = data_i[4545] & sel_one_hot_i[35];
  assign data_masked[4544] = data_i[4544] & sel_one_hot_i[35];
  assign data_masked[4543] = data_i[4543] & sel_one_hot_i[35];
  assign data_masked[4542] = data_i[4542] & sel_one_hot_i[35];
  assign data_masked[4541] = data_i[4541] & sel_one_hot_i[35];
  assign data_masked[4540] = data_i[4540] & sel_one_hot_i[35];
  assign data_masked[4539] = data_i[4539] & sel_one_hot_i[35];
  assign data_masked[4538] = data_i[4538] & sel_one_hot_i[35];
  assign data_masked[4537] = data_i[4537] & sel_one_hot_i[35];
  assign data_masked[4536] = data_i[4536] & sel_one_hot_i[35];
  assign data_masked[4535] = data_i[4535] & sel_one_hot_i[35];
  assign data_masked[4534] = data_i[4534] & sel_one_hot_i[35];
  assign data_masked[4533] = data_i[4533] & sel_one_hot_i[35];
  assign data_masked[4532] = data_i[4532] & sel_one_hot_i[35];
  assign data_masked[4531] = data_i[4531] & sel_one_hot_i[35];
  assign data_masked[4530] = data_i[4530] & sel_one_hot_i[35];
  assign data_masked[4529] = data_i[4529] & sel_one_hot_i[35];
  assign data_masked[4528] = data_i[4528] & sel_one_hot_i[35];
  assign data_masked[4527] = data_i[4527] & sel_one_hot_i[35];
  assign data_masked[4526] = data_i[4526] & sel_one_hot_i[35];
  assign data_masked[4525] = data_i[4525] & sel_one_hot_i[35];
  assign data_masked[4524] = data_i[4524] & sel_one_hot_i[35];
  assign data_masked[4523] = data_i[4523] & sel_one_hot_i[35];
  assign data_masked[4522] = data_i[4522] & sel_one_hot_i[35];
  assign data_masked[4521] = data_i[4521] & sel_one_hot_i[35];
  assign data_masked[4520] = data_i[4520] & sel_one_hot_i[35];
  assign data_masked[4519] = data_i[4519] & sel_one_hot_i[35];
  assign data_masked[4518] = data_i[4518] & sel_one_hot_i[35];
  assign data_masked[4517] = data_i[4517] & sel_one_hot_i[35];
  assign data_masked[4516] = data_i[4516] & sel_one_hot_i[35];
  assign data_masked[4515] = data_i[4515] & sel_one_hot_i[35];
  assign data_masked[4514] = data_i[4514] & sel_one_hot_i[35];
  assign data_masked[4513] = data_i[4513] & sel_one_hot_i[35];
  assign data_masked[4512] = data_i[4512] & sel_one_hot_i[35];
  assign data_masked[4511] = data_i[4511] & sel_one_hot_i[35];
  assign data_masked[4510] = data_i[4510] & sel_one_hot_i[35];
  assign data_masked[4509] = data_i[4509] & sel_one_hot_i[35];
  assign data_masked[4508] = data_i[4508] & sel_one_hot_i[35];
  assign data_masked[4507] = data_i[4507] & sel_one_hot_i[35];
  assign data_masked[4506] = data_i[4506] & sel_one_hot_i[35];
  assign data_masked[4505] = data_i[4505] & sel_one_hot_i[35];
  assign data_masked[4504] = data_i[4504] & sel_one_hot_i[35];
  assign data_masked[4503] = data_i[4503] & sel_one_hot_i[35];
  assign data_masked[4502] = data_i[4502] & sel_one_hot_i[35];
  assign data_masked[4501] = data_i[4501] & sel_one_hot_i[35];
  assign data_masked[4500] = data_i[4500] & sel_one_hot_i[35];
  assign data_masked[4499] = data_i[4499] & sel_one_hot_i[35];
  assign data_masked[4498] = data_i[4498] & sel_one_hot_i[35];
  assign data_masked[4497] = data_i[4497] & sel_one_hot_i[35];
  assign data_masked[4496] = data_i[4496] & sel_one_hot_i[35];
  assign data_masked[4495] = data_i[4495] & sel_one_hot_i[35];
  assign data_masked[4494] = data_i[4494] & sel_one_hot_i[35];
  assign data_masked[4493] = data_i[4493] & sel_one_hot_i[35];
  assign data_masked[4492] = data_i[4492] & sel_one_hot_i[35];
  assign data_masked[4491] = data_i[4491] & sel_one_hot_i[35];
  assign data_masked[4490] = data_i[4490] & sel_one_hot_i[35];
  assign data_masked[4489] = data_i[4489] & sel_one_hot_i[35];
  assign data_masked[4488] = data_i[4488] & sel_one_hot_i[35];
  assign data_masked[4487] = data_i[4487] & sel_one_hot_i[35];
  assign data_masked[4486] = data_i[4486] & sel_one_hot_i[35];
  assign data_masked[4485] = data_i[4485] & sel_one_hot_i[35];
  assign data_masked[4484] = data_i[4484] & sel_one_hot_i[35];
  assign data_masked[4483] = data_i[4483] & sel_one_hot_i[35];
  assign data_masked[4482] = data_i[4482] & sel_one_hot_i[35];
  assign data_masked[4481] = data_i[4481] & sel_one_hot_i[35];
  assign data_masked[4480] = data_i[4480] & sel_one_hot_i[35];
  assign data_masked[4735] = data_i[4735] & sel_one_hot_i[36];
  assign data_masked[4734] = data_i[4734] & sel_one_hot_i[36];
  assign data_masked[4733] = data_i[4733] & sel_one_hot_i[36];
  assign data_masked[4732] = data_i[4732] & sel_one_hot_i[36];
  assign data_masked[4731] = data_i[4731] & sel_one_hot_i[36];
  assign data_masked[4730] = data_i[4730] & sel_one_hot_i[36];
  assign data_masked[4729] = data_i[4729] & sel_one_hot_i[36];
  assign data_masked[4728] = data_i[4728] & sel_one_hot_i[36];
  assign data_masked[4727] = data_i[4727] & sel_one_hot_i[36];
  assign data_masked[4726] = data_i[4726] & sel_one_hot_i[36];
  assign data_masked[4725] = data_i[4725] & sel_one_hot_i[36];
  assign data_masked[4724] = data_i[4724] & sel_one_hot_i[36];
  assign data_masked[4723] = data_i[4723] & sel_one_hot_i[36];
  assign data_masked[4722] = data_i[4722] & sel_one_hot_i[36];
  assign data_masked[4721] = data_i[4721] & sel_one_hot_i[36];
  assign data_masked[4720] = data_i[4720] & sel_one_hot_i[36];
  assign data_masked[4719] = data_i[4719] & sel_one_hot_i[36];
  assign data_masked[4718] = data_i[4718] & sel_one_hot_i[36];
  assign data_masked[4717] = data_i[4717] & sel_one_hot_i[36];
  assign data_masked[4716] = data_i[4716] & sel_one_hot_i[36];
  assign data_masked[4715] = data_i[4715] & sel_one_hot_i[36];
  assign data_masked[4714] = data_i[4714] & sel_one_hot_i[36];
  assign data_masked[4713] = data_i[4713] & sel_one_hot_i[36];
  assign data_masked[4712] = data_i[4712] & sel_one_hot_i[36];
  assign data_masked[4711] = data_i[4711] & sel_one_hot_i[36];
  assign data_masked[4710] = data_i[4710] & sel_one_hot_i[36];
  assign data_masked[4709] = data_i[4709] & sel_one_hot_i[36];
  assign data_masked[4708] = data_i[4708] & sel_one_hot_i[36];
  assign data_masked[4707] = data_i[4707] & sel_one_hot_i[36];
  assign data_masked[4706] = data_i[4706] & sel_one_hot_i[36];
  assign data_masked[4705] = data_i[4705] & sel_one_hot_i[36];
  assign data_masked[4704] = data_i[4704] & sel_one_hot_i[36];
  assign data_masked[4703] = data_i[4703] & sel_one_hot_i[36];
  assign data_masked[4702] = data_i[4702] & sel_one_hot_i[36];
  assign data_masked[4701] = data_i[4701] & sel_one_hot_i[36];
  assign data_masked[4700] = data_i[4700] & sel_one_hot_i[36];
  assign data_masked[4699] = data_i[4699] & sel_one_hot_i[36];
  assign data_masked[4698] = data_i[4698] & sel_one_hot_i[36];
  assign data_masked[4697] = data_i[4697] & sel_one_hot_i[36];
  assign data_masked[4696] = data_i[4696] & sel_one_hot_i[36];
  assign data_masked[4695] = data_i[4695] & sel_one_hot_i[36];
  assign data_masked[4694] = data_i[4694] & sel_one_hot_i[36];
  assign data_masked[4693] = data_i[4693] & sel_one_hot_i[36];
  assign data_masked[4692] = data_i[4692] & sel_one_hot_i[36];
  assign data_masked[4691] = data_i[4691] & sel_one_hot_i[36];
  assign data_masked[4690] = data_i[4690] & sel_one_hot_i[36];
  assign data_masked[4689] = data_i[4689] & sel_one_hot_i[36];
  assign data_masked[4688] = data_i[4688] & sel_one_hot_i[36];
  assign data_masked[4687] = data_i[4687] & sel_one_hot_i[36];
  assign data_masked[4686] = data_i[4686] & sel_one_hot_i[36];
  assign data_masked[4685] = data_i[4685] & sel_one_hot_i[36];
  assign data_masked[4684] = data_i[4684] & sel_one_hot_i[36];
  assign data_masked[4683] = data_i[4683] & sel_one_hot_i[36];
  assign data_masked[4682] = data_i[4682] & sel_one_hot_i[36];
  assign data_masked[4681] = data_i[4681] & sel_one_hot_i[36];
  assign data_masked[4680] = data_i[4680] & sel_one_hot_i[36];
  assign data_masked[4679] = data_i[4679] & sel_one_hot_i[36];
  assign data_masked[4678] = data_i[4678] & sel_one_hot_i[36];
  assign data_masked[4677] = data_i[4677] & sel_one_hot_i[36];
  assign data_masked[4676] = data_i[4676] & sel_one_hot_i[36];
  assign data_masked[4675] = data_i[4675] & sel_one_hot_i[36];
  assign data_masked[4674] = data_i[4674] & sel_one_hot_i[36];
  assign data_masked[4673] = data_i[4673] & sel_one_hot_i[36];
  assign data_masked[4672] = data_i[4672] & sel_one_hot_i[36];
  assign data_masked[4671] = data_i[4671] & sel_one_hot_i[36];
  assign data_masked[4670] = data_i[4670] & sel_one_hot_i[36];
  assign data_masked[4669] = data_i[4669] & sel_one_hot_i[36];
  assign data_masked[4668] = data_i[4668] & sel_one_hot_i[36];
  assign data_masked[4667] = data_i[4667] & sel_one_hot_i[36];
  assign data_masked[4666] = data_i[4666] & sel_one_hot_i[36];
  assign data_masked[4665] = data_i[4665] & sel_one_hot_i[36];
  assign data_masked[4664] = data_i[4664] & sel_one_hot_i[36];
  assign data_masked[4663] = data_i[4663] & sel_one_hot_i[36];
  assign data_masked[4662] = data_i[4662] & sel_one_hot_i[36];
  assign data_masked[4661] = data_i[4661] & sel_one_hot_i[36];
  assign data_masked[4660] = data_i[4660] & sel_one_hot_i[36];
  assign data_masked[4659] = data_i[4659] & sel_one_hot_i[36];
  assign data_masked[4658] = data_i[4658] & sel_one_hot_i[36];
  assign data_masked[4657] = data_i[4657] & sel_one_hot_i[36];
  assign data_masked[4656] = data_i[4656] & sel_one_hot_i[36];
  assign data_masked[4655] = data_i[4655] & sel_one_hot_i[36];
  assign data_masked[4654] = data_i[4654] & sel_one_hot_i[36];
  assign data_masked[4653] = data_i[4653] & sel_one_hot_i[36];
  assign data_masked[4652] = data_i[4652] & sel_one_hot_i[36];
  assign data_masked[4651] = data_i[4651] & sel_one_hot_i[36];
  assign data_masked[4650] = data_i[4650] & sel_one_hot_i[36];
  assign data_masked[4649] = data_i[4649] & sel_one_hot_i[36];
  assign data_masked[4648] = data_i[4648] & sel_one_hot_i[36];
  assign data_masked[4647] = data_i[4647] & sel_one_hot_i[36];
  assign data_masked[4646] = data_i[4646] & sel_one_hot_i[36];
  assign data_masked[4645] = data_i[4645] & sel_one_hot_i[36];
  assign data_masked[4644] = data_i[4644] & sel_one_hot_i[36];
  assign data_masked[4643] = data_i[4643] & sel_one_hot_i[36];
  assign data_masked[4642] = data_i[4642] & sel_one_hot_i[36];
  assign data_masked[4641] = data_i[4641] & sel_one_hot_i[36];
  assign data_masked[4640] = data_i[4640] & sel_one_hot_i[36];
  assign data_masked[4639] = data_i[4639] & sel_one_hot_i[36];
  assign data_masked[4638] = data_i[4638] & sel_one_hot_i[36];
  assign data_masked[4637] = data_i[4637] & sel_one_hot_i[36];
  assign data_masked[4636] = data_i[4636] & sel_one_hot_i[36];
  assign data_masked[4635] = data_i[4635] & sel_one_hot_i[36];
  assign data_masked[4634] = data_i[4634] & sel_one_hot_i[36];
  assign data_masked[4633] = data_i[4633] & sel_one_hot_i[36];
  assign data_masked[4632] = data_i[4632] & sel_one_hot_i[36];
  assign data_masked[4631] = data_i[4631] & sel_one_hot_i[36];
  assign data_masked[4630] = data_i[4630] & sel_one_hot_i[36];
  assign data_masked[4629] = data_i[4629] & sel_one_hot_i[36];
  assign data_masked[4628] = data_i[4628] & sel_one_hot_i[36];
  assign data_masked[4627] = data_i[4627] & sel_one_hot_i[36];
  assign data_masked[4626] = data_i[4626] & sel_one_hot_i[36];
  assign data_masked[4625] = data_i[4625] & sel_one_hot_i[36];
  assign data_masked[4624] = data_i[4624] & sel_one_hot_i[36];
  assign data_masked[4623] = data_i[4623] & sel_one_hot_i[36];
  assign data_masked[4622] = data_i[4622] & sel_one_hot_i[36];
  assign data_masked[4621] = data_i[4621] & sel_one_hot_i[36];
  assign data_masked[4620] = data_i[4620] & sel_one_hot_i[36];
  assign data_masked[4619] = data_i[4619] & sel_one_hot_i[36];
  assign data_masked[4618] = data_i[4618] & sel_one_hot_i[36];
  assign data_masked[4617] = data_i[4617] & sel_one_hot_i[36];
  assign data_masked[4616] = data_i[4616] & sel_one_hot_i[36];
  assign data_masked[4615] = data_i[4615] & sel_one_hot_i[36];
  assign data_masked[4614] = data_i[4614] & sel_one_hot_i[36];
  assign data_masked[4613] = data_i[4613] & sel_one_hot_i[36];
  assign data_masked[4612] = data_i[4612] & sel_one_hot_i[36];
  assign data_masked[4611] = data_i[4611] & sel_one_hot_i[36];
  assign data_masked[4610] = data_i[4610] & sel_one_hot_i[36];
  assign data_masked[4609] = data_i[4609] & sel_one_hot_i[36];
  assign data_masked[4608] = data_i[4608] & sel_one_hot_i[36];
  assign data_masked[4863] = data_i[4863] & sel_one_hot_i[37];
  assign data_masked[4862] = data_i[4862] & sel_one_hot_i[37];
  assign data_masked[4861] = data_i[4861] & sel_one_hot_i[37];
  assign data_masked[4860] = data_i[4860] & sel_one_hot_i[37];
  assign data_masked[4859] = data_i[4859] & sel_one_hot_i[37];
  assign data_masked[4858] = data_i[4858] & sel_one_hot_i[37];
  assign data_masked[4857] = data_i[4857] & sel_one_hot_i[37];
  assign data_masked[4856] = data_i[4856] & sel_one_hot_i[37];
  assign data_masked[4855] = data_i[4855] & sel_one_hot_i[37];
  assign data_masked[4854] = data_i[4854] & sel_one_hot_i[37];
  assign data_masked[4853] = data_i[4853] & sel_one_hot_i[37];
  assign data_masked[4852] = data_i[4852] & sel_one_hot_i[37];
  assign data_masked[4851] = data_i[4851] & sel_one_hot_i[37];
  assign data_masked[4850] = data_i[4850] & sel_one_hot_i[37];
  assign data_masked[4849] = data_i[4849] & sel_one_hot_i[37];
  assign data_masked[4848] = data_i[4848] & sel_one_hot_i[37];
  assign data_masked[4847] = data_i[4847] & sel_one_hot_i[37];
  assign data_masked[4846] = data_i[4846] & sel_one_hot_i[37];
  assign data_masked[4845] = data_i[4845] & sel_one_hot_i[37];
  assign data_masked[4844] = data_i[4844] & sel_one_hot_i[37];
  assign data_masked[4843] = data_i[4843] & sel_one_hot_i[37];
  assign data_masked[4842] = data_i[4842] & sel_one_hot_i[37];
  assign data_masked[4841] = data_i[4841] & sel_one_hot_i[37];
  assign data_masked[4840] = data_i[4840] & sel_one_hot_i[37];
  assign data_masked[4839] = data_i[4839] & sel_one_hot_i[37];
  assign data_masked[4838] = data_i[4838] & sel_one_hot_i[37];
  assign data_masked[4837] = data_i[4837] & sel_one_hot_i[37];
  assign data_masked[4836] = data_i[4836] & sel_one_hot_i[37];
  assign data_masked[4835] = data_i[4835] & sel_one_hot_i[37];
  assign data_masked[4834] = data_i[4834] & sel_one_hot_i[37];
  assign data_masked[4833] = data_i[4833] & sel_one_hot_i[37];
  assign data_masked[4832] = data_i[4832] & sel_one_hot_i[37];
  assign data_masked[4831] = data_i[4831] & sel_one_hot_i[37];
  assign data_masked[4830] = data_i[4830] & sel_one_hot_i[37];
  assign data_masked[4829] = data_i[4829] & sel_one_hot_i[37];
  assign data_masked[4828] = data_i[4828] & sel_one_hot_i[37];
  assign data_masked[4827] = data_i[4827] & sel_one_hot_i[37];
  assign data_masked[4826] = data_i[4826] & sel_one_hot_i[37];
  assign data_masked[4825] = data_i[4825] & sel_one_hot_i[37];
  assign data_masked[4824] = data_i[4824] & sel_one_hot_i[37];
  assign data_masked[4823] = data_i[4823] & sel_one_hot_i[37];
  assign data_masked[4822] = data_i[4822] & sel_one_hot_i[37];
  assign data_masked[4821] = data_i[4821] & sel_one_hot_i[37];
  assign data_masked[4820] = data_i[4820] & sel_one_hot_i[37];
  assign data_masked[4819] = data_i[4819] & sel_one_hot_i[37];
  assign data_masked[4818] = data_i[4818] & sel_one_hot_i[37];
  assign data_masked[4817] = data_i[4817] & sel_one_hot_i[37];
  assign data_masked[4816] = data_i[4816] & sel_one_hot_i[37];
  assign data_masked[4815] = data_i[4815] & sel_one_hot_i[37];
  assign data_masked[4814] = data_i[4814] & sel_one_hot_i[37];
  assign data_masked[4813] = data_i[4813] & sel_one_hot_i[37];
  assign data_masked[4812] = data_i[4812] & sel_one_hot_i[37];
  assign data_masked[4811] = data_i[4811] & sel_one_hot_i[37];
  assign data_masked[4810] = data_i[4810] & sel_one_hot_i[37];
  assign data_masked[4809] = data_i[4809] & sel_one_hot_i[37];
  assign data_masked[4808] = data_i[4808] & sel_one_hot_i[37];
  assign data_masked[4807] = data_i[4807] & sel_one_hot_i[37];
  assign data_masked[4806] = data_i[4806] & sel_one_hot_i[37];
  assign data_masked[4805] = data_i[4805] & sel_one_hot_i[37];
  assign data_masked[4804] = data_i[4804] & sel_one_hot_i[37];
  assign data_masked[4803] = data_i[4803] & sel_one_hot_i[37];
  assign data_masked[4802] = data_i[4802] & sel_one_hot_i[37];
  assign data_masked[4801] = data_i[4801] & sel_one_hot_i[37];
  assign data_masked[4800] = data_i[4800] & sel_one_hot_i[37];
  assign data_masked[4799] = data_i[4799] & sel_one_hot_i[37];
  assign data_masked[4798] = data_i[4798] & sel_one_hot_i[37];
  assign data_masked[4797] = data_i[4797] & sel_one_hot_i[37];
  assign data_masked[4796] = data_i[4796] & sel_one_hot_i[37];
  assign data_masked[4795] = data_i[4795] & sel_one_hot_i[37];
  assign data_masked[4794] = data_i[4794] & sel_one_hot_i[37];
  assign data_masked[4793] = data_i[4793] & sel_one_hot_i[37];
  assign data_masked[4792] = data_i[4792] & sel_one_hot_i[37];
  assign data_masked[4791] = data_i[4791] & sel_one_hot_i[37];
  assign data_masked[4790] = data_i[4790] & sel_one_hot_i[37];
  assign data_masked[4789] = data_i[4789] & sel_one_hot_i[37];
  assign data_masked[4788] = data_i[4788] & sel_one_hot_i[37];
  assign data_masked[4787] = data_i[4787] & sel_one_hot_i[37];
  assign data_masked[4786] = data_i[4786] & sel_one_hot_i[37];
  assign data_masked[4785] = data_i[4785] & sel_one_hot_i[37];
  assign data_masked[4784] = data_i[4784] & sel_one_hot_i[37];
  assign data_masked[4783] = data_i[4783] & sel_one_hot_i[37];
  assign data_masked[4782] = data_i[4782] & sel_one_hot_i[37];
  assign data_masked[4781] = data_i[4781] & sel_one_hot_i[37];
  assign data_masked[4780] = data_i[4780] & sel_one_hot_i[37];
  assign data_masked[4779] = data_i[4779] & sel_one_hot_i[37];
  assign data_masked[4778] = data_i[4778] & sel_one_hot_i[37];
  assign data_masked[4777] = data_i[4777] & sel_one_hot_i[37];
  assign data_masked[4776] = data_i[4776] & sel_one_hot_i[37];
  assign data_masked[4775] = data_i[4775] & sel_one_hot_i[37];
  assign data_masked[4774] = data_i[4774] & sel_one_hot_i[37];
  assign data_masked[4773] = data_i[4773] & sel_one_hot_i[37];
  assign data_masked[4772] = data_i[4772] & sel_one_hot_i[37];
  assign data_masked[4771] = data_i[4771] & sel_one_hot_i[37];
  assign data_masked[4770] = data_i[4770] & sel_one_hot_i[37];
  assign data_masked[4769] = data_i[4769] & sel_one_hot_i[37];
  assign data_masked[4768] = data_i[4768] & sel_one_hot_i[37];
  assign data_masked[4767] = data_i[4767] & sel_one_hot_i[37];
  assign data_masked[4766] = data_i[4766] & sel_one_hot_i[37];
  assign data_masked[4765] = data_i[4765] & sel_one_hot_i[37];
  assign data_masked[4764] = data_i[4764] & sel_one_hot_i[37];
  assign data_masked[4763] = data_i[4763] & sel_one_hot_i[37];
  assign data_masked[4762] = data_i[4762] & sel_one_hot_i[37];
  assign data_masked[4761] = data_i[4761] & sel_one_hot_i[37];
  assign data_masked[4760] = data_i[4760] & sel_one_hot_i[37];
  assign data_masked[4759] = data_i[4759] & sel_one_hot_i[37];
  assign data_masked[4758] = data_i[4758] & sel_one_hot_i[37];
  assign data_masked[4757] = data_i[4757] & sel_one_hot_i[37];
  assign data_masked[4756] = data_i[4756] & sel_one_hot_i[37];
  assign data_masked[4755] = data_i[4755] & sel_one_hot_i[37];
  assign data_masked[4754] = data_i[4754] & sel_one_hot_i[37];
  assign data_masked[4753] = data_i[4753] & sel_one_hot_i[37];
  assign data_masked[4752] = data_i[4752] & sel_one_hot_i[37];
  assign data_masked[4751] = data_i[4751] & sel_one_hot_i[37];
  assign data_masked[4750] = data_i[4750] & sel_one_hot_i[37];
  assign data_masked[4749] = data_i[4749] & sel_one_hot_i[37];
  assign data_masked[4748] = data_i[4748] & sel_one_hot_i[37];
  assign data_masked[4747] = data_i[4747] & sel_one_hot_i[37];
  assign data_masked[4746] = data_i[4746] & sel_one_hot_i[37];
  assign data_masked[4745] = data_i[4745] & sel_one_hot_i[37];
  assign data_masked[4744] = data_i[4744] & sel_one_hot_i[37];
  assign data_masked[4743] = data_i[4743] & sel_one_hot_i[37];
  assign data_masked[4742] = data_i[4742] & sel_one_hot_i[37];
  assign data_masked[4741] = data_i[4741] & sel_one_hot_i[37];
  assign data_masked[4740] = data_i[4740] & sel_one_hot_i[37];
  assign data_masked[4739] = data_i[4739] & sel_one_hot_i[37];
  assign data_masked[4738] = data_i[4738] & sel_one_hot_i[37];
  assign data_masked[4737] = data_i[4737] & sel_one_hot_i[37];
  assign data_masked[4736] = data_i[4736] & sel_one_hot_i[37];
  assign data_masked[4991] = data_i[4991] & sel_one_hot_i[38];
  assign data_masked[4990] = data_i[4990] & sel_one_hot_i[38];
  assign data_masked[4989] = data_i[4989] & sel_one_hot_i[38];
  assign data_masked[4988] = data_i[4988] & sel_one_hot_i[38];
  assign data_masked[4987] = data_i[4987] & sel_one_hot_i[38];
  assign data_masked[4986] = data_i[4986] & sel_one_hot_i[38];
  assign data_masked[4985] = data_i[4985] & sel_one_hot_i[38];
  assign data_masked[4984] = data_i[4984] & sel_one_hot_i[38];
  assign data_masked[4983] = data_i[4983] & sel_one_hot_i[38];
  assign data_masked[4982] = data_i[4982] & sel_one_hot_i[38];
  assign data_masked[4981] = data_i[4981] & sel_one_hot_i[38];
  assign data_masked[4980] = data_i[4980] & sel_one_hot_i[38];
  assign data_masked[4979] = data_i[4979] & sel_one_hot_i[38];
  assign data_masked[4978] = data_i[4978] & sel_one_hot_i[38];
  assign data_masked[4977] = data_i[4977] & sel_one_hot_i[38];
  assign data_masked[4976] = data_i[4976] & sel_one_hot_i[38];
  assign data_masked[4975] = data_i[4975] & sel_one_hot_i[38];
  assign data_masked[4974] = data_i[4974] & sel_one_hot_i[38];
  assign data_masked[4973] = data_i[4973] & sel_one_hot_i[38];
  assign data_masked[4972] = data_i[4972] & sel_one_hot_i[38];
  assign data_masked[4971] = data_i[4971] & sel_one_hot_i[38];
  assign data_masked[4970] = data_i[4970] & sel_one_hot_i[38];
  assign data_masked[4969] = data_i[4969] & sel_one_hot_i[38];
  assign data_masked[4968] = data_i[4968] & sel_one_hot_i[38];
  assign data_masked[4967] = data_i[4967] & sel_one_hot_i[38];
  assign data_masked[4966] = data_i[4966] & sel_one_hot_i[38];
  assign data_masked[4965] = data_i[4965] & sel_one_hot_i[38];
  assign data_masked[4964] = data_i[4964] & sel_one_hot_i[38];
  assign data_masked[4963] = data_i[4963] & sel_one_hot_i[38];
  assign data_masked[4962] = data_i[4962] & sel_one_hot_i[38];
  assign data_masked[4961] = data_i[4961] & sel_one_hot_i[38];
  assign data_masked[4960] = data_i[4960] & sel_one_hot_i[38];
  assign data_masked[4959] = data_i[4959] & sel_one_hot_i[38];
  assign data_masked[4958] = data_i[4958] & sel_one_hot_i[38];
  assign data_masked[4957] = data_i[4957] & sel_one_hot_i[38];
  assign data_masked[4956] = data_i[4956] & sel_one_hot_i[38];
  assign data_masked[4955] = data_i[4955] & sel_one_hot_i[38];
  assign data_masked[4954] = data_i[4954] & sel_one_hot_i[38];
  assign data_masked[4953] = data_i[4953] & sel_one_hot_i[38];
  assign data_masked[4952] = data_i[4952] & sel_one_hot_i[38];
  assign data_masked[4951] = data_i[4951] & sel_one_hot_i[38];
  assign data_masked[4950] = data_i[4950] & sel_one_hot_i[38];
  assign data_masked[4949] = data_i[4949] & sel_one_hot_i[38];
  assign data_masked[4948] = data_i[4948] & sel_one_hot_i[38];
  assign data_masked[4947] = data_i[4947] & sel_one_hot_i[38];
  assign data_masked[4946] = data_i[4946] & sel_one_hot_i[38];
  assign data_masked[4945] = data_i[4945] & sel_one_hot_i[38];
  assign data_masked[4944] = data_i[4944] & sel_one_hot_i[38];
  assign data_masked[4943] = data_i[4943] & sel_one_hot_i[38];
  assign data_masked[4942] = data_i[4942] & sel_one_hot_i[38];
  assign data_masked[4941] = data_i[4941] & sel_one_hot_i[38];
  assign data_masked[4940] = data_i[4940] & sel_one_hot_i[38];
  assign data_masked[4939] = data_i[4939] & sel_one_hot_i[38];
  assign data_masked[4938] = data_i[4938] & sel_one_hot_i[38];
  assign data_masked[4937] = data_i[4937] & sel_one_hot_i[38];
  assign data_masked[4936] = data_i[4936] & sel_one_hot_i[38];
  assign data_masked[4935] = data_i[4935] & sel_one_hot_i[38];
  assign data_masked[4934] = data_i[4934] & sel_one_hot_i[38];
  assign data_masked[4933] = data_i[4933] & sel_one_hot_i[38];
  assign data_masked[4932] = data_i[4932] & sel_one_hot_i[38];
  assign data_masked[4931] = data_i[4931] & sel_one_hot_i[38];
  assign data_masked[4930] = data_i[4930] & sel_one_hot_i[38];
  assign data_masked[4929] = data_i[4929] & sel_one_hot_i[38];
  assign data_masked[4928] = data_i[4928] & sel_one_hot_i[38];
  assign data_masked[4927] = data_i[4927] & sel_one_hot_i[38];
  assign data_masked[4926] = data_i[4926] & sel_one_hot_i[38];
  assign data_masked[4925] = data_i[4925] & sel_one_hot_i[38];
  assign data_masked[4924] = data_i[4924] & sel_one_hot_i[38];
  assign data_masked[4923] = data_i[4923] & sel_one_hot_i[38];
  assign data_masked[4922] = data_i[4922] & sel_one_hot_i[38];
  assign data_masked[4921] = data_i[4921] & sel_one_hot_i[38];
  assign data_masked[4920] = data_i[4920] & sel_one_hot_i[38];
  assign data_masked[4919] = data_i[4919] & sel_one_hot_i[38];
  assign data_masked[4918] = data_i[4918] & sel_one_hot_i[38];
  assign data_masked[4917] = data_i[4917] & sel_one_hot_i[38];
  assign data_masked[4916] = data_i[4916] & sel_one_hot_i[38];
  assign data_masked[4915] = data_i[4915] & sel_one_hot_i[38];
  assign data_masked[4914] = data_i[4914] & sel_one_hot_i[38];
  assign data_masked[4913] = data_i[4913] & sel_one_hot_i[38];
  assign data_masked[4912] = data_i[4912] & sel_one_hot_i[38];
  assign data_masked[4911] = data_i[4911] & sel_one_hot_i[38];
  assign data_masked[4910] = data_i[4910] & sel_one_hot_i[38];
  assign data_masked[4909] = data_i[4909] & sel_one_hot_i[38];
  assign data_masked[4908] = data_i[4908] & sel_one_hot_i[38];
  assign data_masked[4907] = data_i[4907] & sel_one_hot_i[38];
  assign data_masked[4906] = data_i[4906] & sel_one_hot_i[38];
  assign data_masked[4905] = data_i[4905] & sel_one_hot_i[38];
  assign data_masked[4904] = data_i[4904] & sel_one_hot_i[38];
  assign data_masked[4903] = data_i[4903] & sel_one_hot_i[38];
  assign data_masked[4902] = data_i[4902] & sel_one_hot_i[38];
  assign data_masked[4901] = data_i[4901] & sel_one_hot_i[38];
  assign data_masked[4900] = data_i[4900] & sel_one_hot_i[38];
  assign data_masked[4899] = data_i[4899] & sel_one_hot_i[38];
  assign data_masked[4898] = data_i[4898] & sel_one_hot_i[38];
  assign data_masked[4897] = data_i[4897] & sel_one_hot_i[38];
  assign data_masked[4896] = data_i[4896] & sel_one_hot_i[38];
  assign data_masked[4895] = data_i[4895] & sel_one_hot_i[38];
  assign data_masked[4894] = data_i[4894] & sel_one_hot_i[38];
  assign data_masked[4893] = data_i[4893] & sel_one_hot_i[38];
  assign data_masked[4892] = data_i[4892] & sel_one_hot_i[38];
  assign data_masked[4891] = data_i[4891] & sel_one_hot_i[38];
  assign data_masked[4890] = data_i[4890] & sel_one_hot_i[38];
  assign data_masked[4889] = data_i[4889] & sel_one_hot_i[38];
  assign data_masked[4888] = data_i[4888] & sel_one_hot_i[38];
  assign data_masked[4887] = data_i[4887] & sel_one_hot_i[38];
  assign data_masked[4886] = data_i[4886] & sel_one_hot_i[38];
  assign data_masked[4885] = data_i[4885] & sel_one_hot_i[38];
  assign data_masked[4884] = data_i[4884] & sel_one_hot_i[38];
  assign data_masked[4883] = data_i[4883] & sel_one_hot_i[38];
  assign data_masked[4882] = data_i[4882] & sel_one_hot_i[38];
  assign data_masked[4881] = data_i[4881] & sel_one_hot_i[38];
  assign data_masked[4880] = data_i[4880] & sel_one_hot_i[38];
  assign data_masked[4879] = data_i[4879] & sel_one_hot_i[38];
  assign data_masked[4878] = data_i[4878] & sel_one_hot_i[38];
  assign data_masked[4877] = data_i[4877] & sel_one_hot_i[38];
  assign data_masked[4876] = data_i[4876] & sel_one_hot_i[38];
  assign data_masked[4875] = data_i[4875] & sel_one_hot_i[38];
  assign data_masked[4874] = data_i[4874] & sel_one_hot_i[38];
  assign data_masked[4873] = data_i[4873] & sel_one_hot_i[38];
  assign data_masked[4872] = data_i[4872] & sel_one_hot_i[38];
  assign data_masked[4871] = data_i[4871] & sel_one_hot_i[38];
  assign data_masked[4870] = data_i[4870] & sel_one_hot_i[38];
  assign data_masked[4869] = data_i[4869] & sel_one_hot_i[38];
  assign data_masked[4868] = data_i[4868] & sel_one_hot_i[38];
  assign data_masked[4867] = data_i[4867] & sel_one_hot_i[38];
  assign data_masked[4866] = data_i[4866] & sel_one_hot_i[38];
  assign data_masked[4865] = data_i[4865] & sel_one_hot_i[38];
  assign data_masked[4864] = data_i[4864] & sel_one_hot_i[38];
  assign data_masked[5119] = data_i[5119] & sel_one_hot_i[39];
  assign data_masked[5118] = data_i[5118] & sel_one_hot_i[39];
  assign data_masked[5117] = data_i[5117] & sel_one_hot_i[39];
  assign data_masked[5116] = data_i[5116] & sel_one_hot_i[39];
  assign data_masked[5115] = data_i[5115] & sel_one_hot_i[39];
  assign data_masked[5114] = data_i[5114] & sel_one_hot_i[39];
  assign data_masked[5113] = data_i[5113] & sel_one_hot_i[39];
  assign data_masked[5112] = data_i[5112] & sel_one_hot_i[39];
  assign data_masked[5111] = data_i[5111] & sel_one_hot_i[39];
  assign data_masked[5110] = data_i[5110] & sel_one_hot_i[39];
  assign data_masked[5109] = data_i[5109] & sel_one_hot_i[39];
  assign data_masked[5108] = data_i[5108] & sel_one_hot_i[39];
  assign data_masked[5107] = data_i[5107] & sel_one_hot_i[39];
  assign data_masked[5106] = data_i[5106] & sel_one_hot_i[39];
  assign data_masked[5105] = data_i[5105] & sel_one_hot_i[39];
  assign data_masked[5104] = data_i[5104] & sel_one_hot_i[39];
  assign data_masked[5103] = data_i[5103] & sel_one_hot_i[39];
  assign data_masked[5102] = data_i[5102] & sel_one_hot_i[39];
  assign data_masked[5101] = data_i[5101] & sel_one_hot_i[39];
  assign data_masked[5100] = data_i[5100] & sel_one_hot_i[39];
  assign data_masked[5099] = data_i[5099] & sel_one_hot_i[39];
  assign data_masked[5098] = data_i[5098] & sel_one_hot_i[39];
  assign data_masked[5097] = data_i[5097] & sel_one_hot_i[39];
  assign data_masked[5096] = data_i[5096] & sel_one_hot_i[39];
  assign data_masked[5095] = data_i[5095] & sel_one_hot_i[39];
  assign data_masked[5094] = data_i[5094] & sel_one_hot_i[39];
  assign data_masked[5093] = data_i[5093] & sel_one_hot_i[39];
  assign data_masked[5092] = data_i[5092] & sel_one_hot_i[39];
  assign data_masked[5091] = data_i[5091] & sel_one_hot_i[39];
  assign data_masked[5090] = data_i[5090] & sel_one_hot_i[39];
  assign data_masked[5089] = data_i[5089] & sel_one_hot_i[39];
  assign data_masked[5088] = data_i[5088] & sel_one_hot_i[39];
  assign data_masked[5087] = data_i[5087] & sel_one_hot_i[39];
  assign data_masked[5086] = data_i[5086] & sel_one_hot_i[39];
  assign data_masked[5085] = data_i[5085] & sel_one_hot_i[39];
  assign data_masked[5084] = data_i[5084] & sel_one_hot_i[39];
  assign data_masked[5083] = data_i[5083] & sel_one_hot_i[39];
  assign data_masked[5082] = data_i[5082] & sel_one_hot_i[39];
  assign data_masked[5081] = data_i[5081] & sel_one_hot_i[39];
  assign data_masked[5080] = data_i[5080] & sel_one_hot_i[39];
  assign data_masked[5079] = data_i[5079] & sel_one_hot_i[39];
  assign data_masked[5078] = data_i[5078] & sel_one_hot_i[39];
  assign data_masked[5077] = data_i[5077] & sel_one_hot_i[39];
  assign data_masked[5076] = data_i[5076] & sel_one_hot_i[39];
  assign data_masked[5075] = data_i[5075] & sel_one_hot_i[39];
  assign data_masked[5074] = data_i[5074] & sel_one_hot_i[39];
  assign data_masked[5073] = data_i[5073] & sel_one_hot_i[39];
  assign data_masked[5072] = data_i[5072] & sel_one_hot_i[39];
  assign data_masked[5071] = data_i[5071] & sel_one_hot_i[39];
  assign data_masked[5070] = data_i[5070] & sel_one_hot_i[39];
  assign data_masked[5069] = data_i[5069] & sel_one_hot_i[39];
  assign data_masked[5068] = data_i[5068] & sel_one_hot_i[39];
  assign data_masked[5067] = data_i[5067] & sel_one_hot_i[39];
  assign data_masked[5066] = data_i[5066] & sel_one_hot_i[39];
  assign data_masked[5065] = data_i[5065] & sel_one_hot_i[39];
  assign data_masked[5064] = data_i[5064] & sel_one_hot_i[39];
  assign data_masked[5063] = data_i[5063] & sel_one_hot_i[39];
  assign data_masked[5062] = data_i[5062] & sel_one_hot_i[39];
  assign data_masked[5061] = data_i[5061] & sel_one_hot_i[39];
  assign data_masked[5060] = data_i[5060] & sel_one_hot_i[39];
  assign data_masked[5059] = data_i[5059] & sel_one_hot_i[39];
  assign data_masked[5058] = data_i[5058] & sel_one_hot_i[39];
  assign data_masked[5057] = data_i[5057] & sel_one_hot_i[39];
  assign data_masked[5056] = data_i[5056] & sel_one_hot_i[39];
  assign data_masked[5055] = data_i[5055] & sel_one_hot_i[39];
  assign data_masked[5054] = data_i[5054] & sel_one_hot_i[39];
  assign data_masked[5053] = data_i[5053] & sel_one_hot_i[39];
  assign data_masked[5052] = data_i[5052] & sel_one_hot_i[39];
  assign data_masked[5051] = data_i[5051] & sel_one_hot_i[39];
  assign data_masked[5050] = data_i[5050] & sel_one_hot_i[39];
  assign data_masked[5049] = data_i[5049] & sel_one_hot_i[39];
  assign data_masked[5048] = data_i[5048] & sel_one_hot_i[39];
  assign data_masked[5047] = data_i[5047] & sel_one_hot_i[39];
  assign data_masked[5046] = data_i[5046] & sel_one_hot_i[39];
  assign data_masked[5045] = data_i[5045] & sel_one_hot_i[39];
  assign data_masked[5044] = data_i[5044] & sel_one_hot_i[39];
  assign data_masked[5043] = data_i[5043] & sel_one_hot_i[39];
  assign data_masked[5042] = data_i[5042] & sel_one_hot_i[39];
  assign data_masked[5041] = data_i[5041] & sel_one_hot_i[39];
  assign data_masked[5040] = data_i[5040] & sel_one_hot_i[39];
  assign data_masked[5039] = data_i[5039] & sel_one_hot_i[39];
  assign data_masked[5038] = data_i[5038] & sel_one_hot_i[39];
  assign data_masked[5037] = data_i[5037] & sel_one_hot_i[39];
  assign data_masked[5036] = data_i[5036] & sel_one_hot_i[39];
  assign data_masked[5035] = data_i[5035] & sel_one_hot_i[39];
  assign data_masked[5034] = data_i[5034] & sel_one_hot_i[39];
  assign data_masked[5033] = data_i[5033] & sel_one_hot_i[39];
  assign data_masked[5032] = data_i[5032] & sel_one_hot_i[39];
  assign data_masked[5031] = data_i[5031] & sel_one_hot_i[39];
  assign data_masked[5030] = data_i[5030] & sel_one_hot_i[39];
  assign data_masked[5029] = data_i[5029] & sel_one_hot_i[39];
  assign data_masked[5028] = data_i[5028] & sel_one_hot_i[39];
  assign data_masked[5027] = data_i[5027] & sel_one_hot_i[39];
  assign data_masked[5026] = data_i[5026] & sel_one_hot_i[39];
  assign data_masked[5025] = data_i[5025] & sel_one_hot_i[39];
  assign data_masked[5024] = data_i[5024] & sel_one_hot_i[39];
  assign data_masked[5023] = data_i[5023] & sel_one_hot_i[39];
  assign data_masked[5022] = data_i[5022] & sel_one_hot_i[39];
  assign data_masked[5021] = data_i[5021] & sel_one_hot_i[39];
  assign data_masked[5020] = data_i[5020] & sel_one_hot_i[39];
  assign data_masked[5019] = data_i[5019] & sel_one_hot_i[39];
  assign data_masked[5018] = data_i[5018] & sel_one_hot_i[39];
  assign data_masked[5017] = data_i[5017] & sel_one_hot_i[39];
  assign data_masked[5016] = data_i[5016] & sel_one_hot_i[39];
  assign data_masked[5015] = data_i[5015] & sel_one_hot_i[39];
  assign data_masked[5014] = data_i[5014] & sel_one_hot_i[39];
  assign data_masked[5013] = data_i[5013] & sel_one_hot_i[39];
  assign data_masked[5012] = data_i[5012] & sel_one_hot_i[39];
  assign data_masked[5011] = data_i[5011] & sel_one_hot_i[39];
  assign data_masked[5010] = data_i[5010] & sel_one_hot_i[39];
  assign data_masked[5009] = data_i[5009] & sel_one_hot_i[39];
  assign data_masked[5008] = data_i[5008] & sel_one_hot_i[39];
  assign data_masked[5007] = data_i[5007] & sel_one_hot_i[39];
  assign data_masked[5006] = data_i[5006] & sel_one_hot_i[39];
  assign data_masked[5005] = data_i[5005] & sel_one_hot_i[39];
  assign data_masked[5004] = data_i[5004] & sel_one_hot_i[39];
  assign data_masked[5003] = data_i[5003] & sel_one_hot_i[39];
  assign data_masked[5002] = data_i[5002] & sel_one_hot_i[39];
  assign data_masked[5001] = data_i[5001] & sel_one_hot_i[39];
  assign data_masked[5000] = data_i[5000] & sel_one_hot_i[39];
  assign data_masked[4999] = data_i[4999] & sel_one_hot_i[39];
  assign data_masked[4998] = data_i[4998] & sel_one_hot_i[39];
  assign data_masked[4997] = data_i[4997] & sel_one_hot_i[39];
  assign data_masked[4996] = data_i[4996] & sel_one_hot_i[39];
  assign data_masked[4995] = data_i[4995] & sel_one_hot_i[39];
  assign data_masked[4994] = data_i[4994] & sel_one_hot_i[39];
  assign data_masked[4993] = data_i[4993] & sel_one_hot_i[39];
  assign data_masked[4992] = data_i[4992] & sel_one_hot_i[39];
  assign data_masked[5247] = data_i[5247] & sel_one_hot_i[40];
  assign data_masked[5246] = data_i[5246] & sel_one_hot_i[40];
  assign data_masked[5245] = data_i[5245] & sel_one_hot_i[40];
  assign data_masked[5244] = data_i[5244] & sel_one_hot_i[40];
  assign data_masked[5243] = data_i[5243] & sel_one_hot_i[40];
  assign data_masked[5242] = data_i[5242] & sel_one_hot_i[40];
  assign data_masked[5241] = data_i[5241] & sel_one_hot_i[40];
  assign data_masked[5240] = data_i[5240] & sel_one_hot_i[40];
  assign data_masked[5239] = data_i[5239] & sel_one_hot_i[40];
  assign data_masked[5238] = data_i[5238] & sel_one_hot_i[40];
  assign data_masked[5237] = data_i[5237] & sel_one_hot_i[40];
  assign data_masked[5236] = data_i[5236] & sel_one_hot_i[40];
  assign data_masked[5235] = data_i[5235] & sel_one_hot_i[40];
  assign data_masked[5234] = data_i[5234] & sel_one_hot_i[40];
  assign data_masked[5233] = data_i[5233] & sel_one_hot_i[40];
  assign data_masked[5232] = data_i[5232] & sel_one_hot_i[40];
  assign data_masked[5231] = data_i[5231] & sel_one_hot_i[40];
  assign data_masked[5230] = data_i[5230] & sel_one_hot_i[40];
  assign data_masked[5229] = data_i[5229] & sel_one_hot_i[40];
  assign data_masked[5228] = data_i[5228] & sel_one_hot_i[40];
  assign data_masked[5227] = data_i[5227] & sel_one_hot_i[40];
  assign data_masked[5226] = data_i[5226] & sel_one_hot_i[40];
  assign data_masked[5225] = data_i[5225] & sel_one_hot_i[40];
  assign data_masked[5224] = data_i[5224] & sel_one_hot_i[40];
  assign data_masked[5223] = data_i[5223] & sel_one_hot_i[40];
  assign data_masked[5222] = data_i[5222] & sel_one_hot_i[40];
  assign data_masked[5221] = data_i[5221] & sel_one_hot_i[40];
  assign data_masked[5220] = data_i[5220] & sel_one_hot_i[40];
  assign data_masked[5219] = data_i[5219] & sel_one_hot_i[40];
  assign data_masked[5218] = data_i[5218] & sel_one_hot_i[40];
  assign data_masked[5217] = data_i[5217] & sel_one_hot_i[40];
  assign data_masked[5216] = data_i[5216] & sel_one_hot_i[40];
  assign data_masked[5215] = data_i[5215] & sel_one_hot_i[40];
  assign data_masked[5214] = data_i[5214] & sel_one_hot_i[40];
  assign data_masked[5213] = data_i[5213] & sel_one_hot_i[40];
  assign data_masked[5212] = data_i[5212] & sel_one_hot_i[40];
  assign data_masked[5211] = data_i[5211] & sel_one_hot_i[40];
  assign data_masked[5210] = data_i[5210] & sel_one_hot_i[40];
  assign data_masked[5209] = data_i[5209] & sel_one_hot_i[40];
  assign data_masked[5208] = data_i[5208] & sel_one_hot_i[40];
  assign data_masked[5207] = data_i[5207] & sel_one_hot_i[40];
  assign data_masked[5206] = data_i[5206] & sel_one_hot_i[40];
  assign data_masked[5205] = data_i[5205] & sel_one_hot_i[40];
  assign data_masked[5204] = data_i[5204] & sel_one_hot_i[40];
  assign data_masked[5203] = data_i[5203] & sel_one_hot_i[40];
  assign data_masked[5202] = data_i[5202] & sel_one_hot_i[40];
  assign data_masked[5201] = data_i[5201] & sel_one_hot_i[40];
  assign data_masked[5200] = data_i[5200] & sel_one_hot_i[40];
  assign data_masked[5199] = data_i[5199] & sel_one_hot_i[40];
  assign data_masked[5198] = data_i[5198] & sel_one_hot_i[40];
  assign data_masked[5197] = data_i[5197] & sel_one_hot_i[40];
  assign data_masked[5196] = data_i[5196] & sel_one_hot_i[40];
  assign data_masked[5195] = data_i[5195] & sel_one_hot_i[40];
  assign data_masked[5194] = data_i[5194] & sel_one_hot_i[40];
  assign data_masked[5193] = data_i[5193] & sel_one_hot_i[40];
  assign data_masked[5192] = data_i[5192] & sel_one_hot_i[40];
  assign data_masked[5191] = data_i[5191] & sel_one_hot_i[40];
  assign data_masked[5190] = data_i[5190] & sel_one_hot_i[40];
  assign data_masked[5189] = data_i[5189] & sel_one_hot_i[40];
  assign data_masked[5188] = data_i[5188] & sel_one_hot_i[40];
  assign data_masked[5187] = data_i[5187] & sel_one_hot_i[40];
  assign data_masked[5186] = data_i[5186] & sel_one_hot_i[40];
  assign data_masked[5185] = data_i[5185] & sel_one_hot_i[40];
  assign data_masked[5184] = data_i[5184] & sel_one_hot_i[40];
  assign data_masked[5183] = data_i[5183] & sel_one_hot_i[40];
  assign data_masked[5182] = data_i[5182] & sel_one_hot_i[40];
  assign data_masked[5181] = data_i[5181] & sel_one_hot_i[40];
  assign data_masked[5180] = data_i[5180] & sel_one_hot_i[40];
  assign data_masked[5179] = data_i[5179] & sel_one_hot_i[40];
  assign data_masked[5178] = data_i[5178] & sel_one_hot_i[40];
  assign data_masked[5177] = data_i[5177] & sel_one_hot_i[40];
  assign data_masked[5176] = data_i[5176] & sel_one_hot_i[40];
  assign data_masked[5175] = data_i[5175] & sel_one_hot_i[40];
  assign data_masked[5174] = data_i[5174] & sel_one_hot_i[40];
  assign data_masked[5173] = data_i[5173] & sel_one_hot_i[40];
  assign data_masked[5172] = data_i[5172] & sel_one_hot_i[40];
  assign data_masked[5171] = data_i[5171] & sel_one_hot_i[40];
  assign data_masked[5170] = data_i[5170] & sel_one_hot_i[40];
  assign data_masked[5169] = data_i[5169] & sel_one_hot_i[40];
  assign data_masked[5168] = data_i[5168] & sel_one_hot_i[40];
  assign data_masked[5167] = data_i[5167] & sel_one_hot_i[40];
  assign data_masked[5166] = data_i[5166] & sel_one_hot_i[40];
  assign data_masked[5165] = data_i[5165] & sel_one_hot_i[40];
  assign data_masked[5164] = data_i[5164] & sel_one_hot_i[40];
  assign data_masked[5163] = data_i[5163] & sel_one_hot_i[40];
  assign data_masked[5162] = data_i[5162] & sel_one_hot_i[40];
  assign data_masked[5161] = data_i[5161] & sel_one_hot_i[40];
  assign data_masked[5160] = data_i[5160] & sel_one_hot_i[40];
  assign data_masked[5159] = data_i[5159] & sel_one_hot_i[40];
  assign data_masked[5158] = data_i[5158] & sel_one_hot_i[40];
  assign data_masked[5157] = data_i[5157] & sel_one_hot_i[40];
  assign data_masked[5156] = data_i[5156] & sel_one_hot_i[40];
  assign data_masked[5155] = data_i[5155] & sel_one_hot_i[40];
  assign data_masked[5154] = data_i[5154] & sel_one_hot_i[40];
  assign data_masked[5153] = data_i[5153] & sel_one_hot_i[40];
  assign data_masked[5152] = data_i[5152] & sel_one_hot_i[40];
  assign data_masked[5151] = data_i[5151] & sel_one_hot_i[40];
  assign data_masked[5150] = data_i[5150] & sel_one_hot_i[40];
  assign data_masked[5149] = data_i[5149] & sel_one_hot_i[40];
  assign data_masked[5148] = data_i[5148] & sel_one_hot_i[40];
  assign data_masked[5147] = data_i[5147] & sel_one_hot_i[40];
  assign data_masked[5146] = data_i[5146] & sel_one_hot_i[40];
  assign data_masked[5145] = data_i[5145] & sel_one_hot_i[40];
  assign data_masked[5144] = data_i[5144] & sel_one_hot_i[40];
  assign data_masked[5143] = data_i[5143] & sel_one_hot_i[40];
  assign data_masked[5142] = data_i[5142] & sel_one_hot_i[40];
  assign data_masked[5141] = data_i[5141] & sel_one_hot_i[40];
  assign data_masked[5140] = data_i[5140] & sel_one_hot_i[40];
  assign data_masked[5139] = data_i[5139] & sel_one_hot_i[40];
  assign data_masked[5138] = data_i[5138] & sel_one_hot_i[40];
  assign data_masked[5137] = data_i[5137] & sel_one_hot_i[40];
  assign data_masked[5136] = data_i[5136] & sel_one_hot_i[40];
  assign data_masked[5135] = data_i[5135] & sel_one_hot_i[40];
  assign data_masked[5134] = data_i[5134] & sel_one_hot_i[40];
  assign data_masked[5133] = data_i[5133] & sel_one_hot_i[40];
  assign data_masked[5132] = data_i[5132] & sel_one_hot_i[40];
  assign data_masked[5131] = data_i[5131] & sel_one_hot_i[40];
  assign data_masked[5130] = data_i[5130] & sel_one_hot_i[40];
  assign data_masked[5129] = data_i[5129] & sel_one_hot_i[40];
  assign data_masked[5128] = data_i[5128] & sel_one_hot_i[40];
  assign data_masked[5127] = data_i[5127] & sel_one_hot_i[40];
  assign data_masked[5126] = data_i[5126] & sel_one_hot_i[40];
  assign data_masked[5125] = data_i[5125] & sel_one_hot_i[40];
  assign data_masked[5124] = data_i[5124] & sel_one_hot_i[40];
  assign data_masked[5123] = data_i[5123] & sel_one_hot_i[40];
  assign data_masked[5122] = data_i[5122] & sel_one_hot_i[40];
  assign data_masked[5121] = data_i[5121] & sel_one_hot_i[40];
  assign data_masked[5120] = data_i[5120] & sel_one_hot_i[40];
  assign data_masked[5375] = data_i[5375] & sel_one_hot_i[41];
  assign data_masked[5374] = data_i[5374] & sel_one_hot_i[41];
  assign data_masked[5373] = data_i[5373] & sel_one_hot_i[41];
  assign data_masked[5372] = data_i[5372] & sel_one_hot_i[41];
  assign data_masked[5371] = data_i[5371] & sel_one_hot_i[41];
  assign data_masked[5370] = data_i[5370] & sel_one_hot_i[41];
  assign data_masked[5369] = data_i[5369] & sel_one_hot_i[41];
  assign data_masked[5368] = data_i[5368] & sel_one_hot_i[41];
  assign data_masked[5367] = data_i[5367] & sel_one_hot_i[41];
  assign data_masked[5366] = data_i[5366] & sel_one_hot_i[41];
  assign data_masked[5365] = data_i[5365] & sel_one_hot_i[41];
  assign data_masked[5364] = data_i[5364] & sel_one_hot_i[41];
  assign data_masked[5363] = data_i[5363] & sel_one_hot_i[41];
  assign data_masked[5362] = data_i[5362] & sel_one_hot_i[41];
  assign data_masked[5361] = data_i[5361] & sel_one_hot_i[41];
  assign data_masked[5360] = data_i[5360] & sel_one_hot_i[41];
  assign data_masked[5359] = data_i[5359] & sel_one_hot_i[41];
  assign data_masked[5358] = data_i[5358] & sel_one_hot_i[41];
  assign data_masked[5357] = data_i[5357] & sel_one_hot_i[41];
  assign data_masked[5356] = data_i[5356] & sel_one_hot_i[41];
  assign data_masked[5355] = data_i[5355] & sel_one_hot_i[41];
  assign data_masked[5354] = data_i[5354] & sel_one_hot_i[41];
  assign data_masked[5353] = data_i[5353] & sel_one_hot_i[41];
  assign data_masked[5352] = data_i[5352] & sel_one_hot_i[41];
  assign data_masked[5351] = data_i[5351] & sel_one_hot_i[41];
  assign data_masked[5350] = data_i[5350] & sel_one_hot_i[41];
  assign data_masked[5349] = data_i[5349] & sel_one_hot_i[41];
  assign data_masked[5348] = data_i[5348] & sel_one_hot_i[41];
  assign data_masked[5347] = data_i[5347] & sel_one_hot_i[41];
  assign data_masked[5346] = data_i[5346] & sel_one_hot_i[41];
  assign data_masked[5345] = data_i[5345] & sel_one_hot_i[41];
  assign data_masked[5344] = data_i[5344] & sel_one_hot_i[41];
  assign data_masked[5343] = data_i[5343] & sel_one_hot_i[41];
  assign data_masked[5342] = data_i[5342] & sel_one_hot_i[41];
  assign data_masked[5341] = data_i[5341] & sel_one_hot_i[41];
  assign data_masked[5340] = data_i[5340] & sel_one_hot_i[41];
  assign data_masked[5339] = data_i[5339] & sel_one_hot_i[41];
  assign data_masked[5338] = data_i[5338] & sel_one_hot_i[41];
  assign data_masked[5337] = data_i[5337] & sel_one_hot_i[41];
  assign data_masked[5336] = data_i[5336] & sel_one_hot_i[41];
  assign data_masked[5335] = data_i[5335] & sel_one_hot_i[41];
  assign data_masked[5334] = data_i[5334] & sel_one_hot_i[41];
  assign data_masked[5333] = data_i[5333] & sel_one_hot_i[41];
  assign data_masked[5332] = data_i[5332] & sel_one_hot_i[41];
  assign data_masked[5331] = data_i[5331] & sel_one_hot_i[41];
  assign data_masked[5330] = data_i[5330] & sel_one_hot_i[41];
  assign data_masked[5329] = data_i[5329] & sel_one_hot_i[41];
  assign data_masked[5328] = data_i[5328] & sel_one_hot_i[41];
  assign data_masked[5327] = data_i[5327] & sel_one_hot_i[41];
  assign data_masked[5326] = data_i[5326] & sel_one_hot_i[41];
  assign data_masked[5325] = data_i[5325] & sel_one_hot_i[41];
  assign data_masked[5324] = data_i[5324] & sel_one_hot_i[41];
  assign data_masked[5323] = data_i[5323] & sel_one_hot_i[41];
  assign data_masked[5322] = data_i[5322] & sel_one_hot_i[41];
  assign data_masked[5321] = data_i[5321] & sel_one_hot_i[41];
  assign data_masked[5320] = data_i[5320] & sel_one_hot_i[41];
  assign data_masked[5319] = data_i[5319] & sel_one_hot_i[41];
  assign data_masked[5318] = data_i[5318] & sel_one_hot_i[41];
  assign data_masked[5317] = data_i[5317] & sel_one_hot_i[41];
  assign data_masked[5316] = data_i[5316] & sel_one_hot_i[41];
  assign data_masked[5315] = data_i[5315] & sel_one_hot_i[41];
  assign data_masked[5314] = data_i[5314] & sel_one_hot_i[41];
  assign data_masked[5313] = data_i[5313] & sel_one_hot_i[41];
  assign data_masked[5312] = data_i[5312] & sel_one_hot_i[41];
  assign data_masked[5311] = data_i[5311] & sel_one_hot_i[41];
  assign data_masked[5310] = data_i[5310] & sel_one_hot_i[41];
  assign data_masked[5309] = data_i[5309] & sel_one_hot_i[41];
  assign data_masked[5308] = data_i[5308] & sel_one_hot_i[41];
  assign data_masked[5307] = data_i[5307] & sel_one_hot_i[41];
  assign data_masked[5306] = data_i[5306] & sel_one_hot_i[41];
  assign data_masked[5305] = data_i[5305] & sel_one_hot_i[41];
  assign data_masked[5304] = data_i[5304] & sel_one_hot_i[41];
  assign data_masked[5303] = data_i[5303] & sel_one_hot_i[41];
  assign data_masked[5302] = data_i[5302] & sel_one_hot_i[41];
  assign data_masked[5301] = data_i[5301] & sel_one_hot_i[41];
  assign data_masked[5300] = data_i[5300] & sel_one_hot_i[41];
  assign data_masked[5299] = data_i[5299] & sel_one_hot_i[41];
  assign data_masked[5298] = data_i[5298] & sel_one_hot_i[41];
  assign data_masked[5297] = data_i[5297] & sel_one_hot_i[41];
  assign data_masked[5296] = data_i[5296] & sel_one_hot_i[41];
  assign data_masked[5295] = data_i[5295] & sel_one_hot_i[41];
  assign data_masked[5294] = data_i[5294] & sel_one_hot_i[41];
  assign data_masked[5293] = data_i[5293] & sel_one_hot_i[41];
  assign data_masked[5292] = data_i[5292] & sel_one_hot_i[41];
  assign data_masked[5291] = data_i[5291] & sel_one_hot_i[41];
  assign data_masked[5290] = data_i[5290] & sel_one_hot_i[41];
  assign data_masked[5289] = data_i[5289] & sel_one_hot_i[41];
  assign data_masked[5288] = data_i[5288] & sel_one_hot_i[41];
  assign data_masked[5287] = data_i[5287] & sel_one_hot_i[41];
  assign data_masked[5286] = data_i[5286] & sel_one_hot_i[41];
  assign data_masked[5285] = data_i[5285] & sel_one_hot_i[41];
  assign data_masked[5284] = data_i[5284] & sel_one_hot_i[41];
  assign data_masked[5283] = data_i[5283] & sel_one_hot_i[41];
  assign data_masked[5282] = data_i[5282] & sel_one_hot_i[41];
  assign data_masked[5281] = data_i[5281] & sel_one_hot_i[41];
  assign data_masked[5280] = data_i[5280] & sel_one_hot_i[41];
  assign data_masked[5279] = data_i[5279] & sel_one_hot_i[41];
  assign data_masked[5278] = data_i[5278] & sel_one_hot_i[41];
  assign data_masked[5277] = data_i[5277] & sel_one_hot_i[41];
  assign data_masked[5276] = data_i[5276] & sel_one_hot_i[41];
  assign data_masked[5275] = data_i[5275] & sel_one_hot_i[41];
  assign data_masked[5274] = data_i[5274] & sel_one_hot_i[41];
  assign data_masked[5273] = data_i[5273] & sel_one_hot_i[41];
  assign data_masked[5272] = data_i[5272] & sel_one_hot_i[41];
  assign data_masked[5271] = data_i[5271] & sel_one_hot_i[41];
  assign data_masked[5270] = data_i[5270] & sel_one_hot_i[41];
  assign data_masked[5269] = data_i[5269] & sel_one_hot_i[41];
  assign data_masked[5268] = data_i[5268] & sel_one_hot_i[41];
  assign data_masked[5267] = data_i[5267] & sel_one_hot_i[41];
  assign data_masked[5266] = data_i[5266] & sel_one_hot_i[41];
  assign data_masked[5265] = data_i[5265] & sel_one_hot_i[41];
  assign data_masked[5264] = data_i[5264] & sel_one_hot_i[41];
  assign data_masked[5263] = data_i[5263] & sel_one_hot_i[41];
  assign data_masked[5262] = data_i[5262] & sel_one_hot_i[41];
  assign data_masked[5261] = data_i[5261] & sel_one_hot_i[41];
  assign data_masked[5260] = data_i[5260] & sel_one_hot_i[41];
  assign data_masked[5259] = data_i[5259] & sel_one_hot_i[41];
  assign data_masked[5258] = data_i[5258] & sel_one_hot_i[41];
  assign data_masked[5257] = data_i[5257] & sel_one_hot_i[41];
  assign data_masked[5256] = data_i[5256] & sel_one_hot_i[41];
  assign data_masked[5255] = data_i[5255] & sel_one_hot_i[41];
  assign data_masked[5254] = data_i[5254] & sel_one_hot_i[41];
  assign data_masked[5253] = data_i[5253] & sel_one_hot_i[41];
  assign data_masked[5252] = data_i[5252] & sel_one_hot_i[41];
  assign data_masked[5251] = data_i[5251] & sel_one_hot_i[41];
  assign data_masked[5250] = data_i[5250] & sel_one_hot_i[41];
  assign data_masked[5249] = data_i[5249] & sel_one_hot_i[41];
  assign data_masked[5248] = data_i[5248] & sel_one_hot_i[41];
  assign data_masked[5503] = data_i[5503] & sel_one_hot_i[42];
  assign data_masked[5502] = data_i[5502] & sel_one_hot_i[42];
  assign data_masked[5501] = data_i[5501] & sel_one_hot_i[42];
  assign data_masked[5500] = data_i[5500] & sel_one_hot_i[42];
  assign data_masked[5499] = data_i[5499] & sel_one_hot_i[42];
  assign data_masked[5498] = data_i[5498] & sel_one_hot_i[42];
  assign data_masked[5497] = data_i[5497] & sel_one_hot_i[42];
  assign data_masked[5496] = data_i[5496] & sel_one_hot_i[42];
  assign data_masked[5495] = data_i[5495] & sel_one_hot_i[42];
  assign data_masked[5494] = data_i[5494] & sel_one_hot_i[42];
  assign data_masked[5493] = data_i[5493] & sel_one_hot_i[42];
  assign data_masked[5492] = data_i[5492] & sel_one_hot_i[42];
  assign data_masked[5491] = data_i[5491] & sel_one_hot_i[42];
  assign data_masked[5490] = data_i[5490] & sel_one_hot_i[42];
  assign data_masked[5489] = data_i[5489] & sel_one_hot_i[42];
  assign data_masked[5488] = data_i[5488] & sel_one_hot_i[42];
  assign data_masked[5487] = data_i[5487] & sel_one_hot_i[42];
  assign data_masked[5486] = data_i[5486] & sel_one_hot_i[42];
  assign data_masked[5485] = data_i[5485] & sel_one_hot_i[42];
  assign data_masked[5484] = data_i[5484] & sel_one_hot_i[42];
  assign data_masked[5483] = data_i[5483] & sel_one_hot_i[42];
  assign data_masked[5482] = data_i[5482] & sel_one_hot_i[42];
  assign data_masked[5481] = data_i[5481] & sel_one_hot_i[42];
  assign data_masked[5480] = data_i[5480] & sel_one_hot_i[42];
  assign data_masked[5479] = data_i[5479] & sel_one_hot_i[42];
  assign data_masked[5478] = data_i[5478] & sel_one_hot_i[42];
  assign data_masked[5477] = data_i[5477] & sel_one_hot_i[42];
  assign data_masked[5476] = data_i[5476] & sel_one_hot_i[42];
  assign data_masked[5475] = data_i[5475] & sel_one_hot_i[42];
  assign data_masked[5474] = data_i[5474] & sel_one_hot_i[42];
  assign data_masked[5473] = data_i[5473] & sel_one_hot_i[42];
  assign data_masked[5472] = data_i[5472] & sel_one_hot_i[42];
  assign data_masked[5471] = data_i[5471] & sel_one_hot_i[42];
  assign data_masked[5470] = data_i[5470] & sel_one_hot_i[42];
  assign data_masked[5469] = data_i[5469] & sel_one_hot_i[42];
  assign data_masked[5468] = data_i[5468] & sel_one_hot_i[42];
  assign data_masked[5467] = data_i[5467] & sel_one_hot_i[42];
  assign data_masked[5466] = data_i[5466] & sel_one_hot_i[42];
  assign data_masked[5465] = data_i[5465] & sel_one_hot_i[42];
  assign data_masked[5464] = data_i[5464] & sel_one_hot_i[42];
  assign data_masked[5463] = data_i[5463] & sel_one_hot_i[42];
  assign data_masked[5462] = data_i[5462] & sel_one_hot_i[42];
  assign data_masked[5461] = data_i[5461] & sel_one_hot_i[42];
  assign data_masked[5460] = data_i[5460] & sel_one_hot_i[42];
  assign data_masked[5459] = data_i[5459] & sel_one_hot_i[42];
  assign data_masked[5458] = data_i[5458] & sel_one_hot_i[42];
  assign data_masked[5457] = data_i[5457] & sel_one_hot_i[42];
  assign data_masked[5456] = data_i[5456] & sel_one_hot_i[42];
  assign data_masked[5455] = data_i[5455] & sel_one_hot_i[42];
  assign data_masked[5454] = data_i[5454] & sel_one_hot_i[42];
  assign data_masked[5453] = data_i[5453] & sel_one_hot_i[42];
  assign data_masked[5452] = data_i[5452] & sel_one_hot_i[42];
  assign data_masked[5451] = data_i[5451] & sel_one_hot_i[42];
  assign data_masked[5450] = data_i[5450] & sel_one_hot_i[42];
  assign data_masked[5449] = data_i[5449] & sel_one_hot_i[42];
  assign data_masked[5448] = data_i[5448] & sel_one_hot_i[42];
  assign data_masked[5447] = data_i[5447] & sel_one_hot_i[42];
  assign data_masked[5446] = data_i[5446] & sel_one_hot_i[42];
  assign data_masked[5445] = data_i[5445] & sel_one_hot_i[42];
  assign data_masked[5444] = data_i[5444] & sel_one_hot_i[42];
  assign data_masked[5443] = data_i[5443] & sel_one_hot_i[42];
  assign data_masked[5442] = data_i[5442] & sel_one_hot_i[42];
  assign data_masked[5441] = data_i[5441] & sel_one_hot_i[42];
  assign data_masked[5440] = data_i[5440] & sel_one_hot_i[42];
  assign data_masked[5439] = data_i[5439] & sel_one_hot_i[42];
  assign data_masked[5438] = data_i[5438] & sel_one_hot_i[42];
  assign data_masked[5437] = data_i[5437] & sel_one_hot_i[42];
  assign data_masked[5436] = data_i[5436] & sel_one_hot_i[42];
  assign data_masked[5435] = data_i[5435] & sel_one_hot_i[42];
  assign data_masked[5434] = data_i[5434] & sel_one_hot_i[42];
  assign data_masked[5433] = data_i[5433] & sel_one_hot_i[42];
  assign data_masked[5432] = data_i[5432] & sel_one_hot_i[42];
  assign data_masked[5431] = data_i[5431] & sel_one_hot_i[42];
  assign data_masked[5430] = data_i[5430] & sel_one_hot_i[42];
  assign data_masked[5429] = data_i[5429] & sel_one_hot_i[42];
  assign data_masked[5428] = data_i[5428] & sel_one_hot_i[42];
  assign data_masked[5427] = data_i[5427] & sel_one_hot_i[42];
  assign data_masked[5426] = data_i[5426] & sel_one_hot_i[42];
  assign data_masked[5425] = data_i[5425] & sel_one_hot_i[42];
  assign data_masked[5424] = data_i[5424] & sel_one_hot_i[42];
  assign data_masked[5423] = data_i[5423] & sel_one_hot_i[42];
  assign data_masked[5422] = data_i[5422] & sel_one_hot_i[42];
  assign data_masked[5421] = data_i[5421] & sel_one_hot_i[42];
  assign data_masked[5420] = data_i[5420] & sel_one_hot_i[42];
  assign data_masked[5419] = data_i[5419] & sel_one_hot_i[42];
  assign data_masked[5418] = data_i[5418] & sel_one_hot_i[42];
  assign data_masked[5417] = data_i[5417] & sel_one_hot_i[42];
  assign data_masked[5416] = data_i[5416] & sel_one_hot_i[42];
  assign data_masked[5415] = data_i[5415] & sel_one_hot_i[42];
  assign data_masked[5414] = data_i[5414] & sel_one_hot_i[42];
  assign data_masked[5413] = data_i[5413] & sel_one_hot_i[42];
  assign data_masked[5412] = data_i[5412] & sel_one_hot_i[42];
  assign data_masked[5411] = data_i[5411] & sel_one_hot_i[42];
  assign data_masked[5410] = data_i[5410] & sel_one_hot_i[42];
  assign data_masked[5409] = data_i[5409] & sel_one_hot_i[42];
  assign data_masked[5408] = data_i[5408] & sel_one_hot_i[42];
  assign data_masked[5407] = data_i[5407] & sel_one_hot_i[42];
  assign data_masked[5406] = data_i[5406] & sel_one_hot_i[42];
  assign data_masked[5405] = data_i[5405] & sel_one_hot_i[42];
  assign data_masked[5404] = data_i[5404] & sel_one_hot_i[42];
  assign data_masked[5403] = data_i[5403] & sel_one_hot_i[42];
  assign data_masked[5402] = data_i[5402] & sel_one_hot_i[42];
  assign data_masked[5401] = data_i[5401] & sel_one_hot_i[42];
  assign data_masked[5400] = data_i[5400] & sel_one_hot_i[42];
  assign data_masked[5399] = data_i[5399] & sel_one_hot_i[42];
  assign data_masked[5398] = data_i[5398] & sel_one_hot_i[42];
  assign data_masked[5397] = data_i[5397] & sel_one_hot_i[42];
  assign data_masked[5396] = data_i[5396] & sel_one_hot_i[42];
  assign data_masked[5395] = data_i[5395] & sel_one_hot_i[42];
  assign data_masked[5394] = data_i[5394] & sel_one_hot_i[42];
  assign data_masked[5393] = data_i[5393] & sel_one_hot_i[42];
  assign data_masked[5392] = data_i[5392] & sel_one_hot_i[42];
  assign data_masked[5391] = data_i[5391] & sel_one_hot_i[42];
  assign data_masked[5390] = data_i[5390] & sel_one_hot_i[42];
  assign data_masked[5389] = data_i[5389] & sel_one_hot_i[42];
  assign data_masked[5388] = data_i[5388] & sel_one_hot_i[42];
  assign data_masked[5387] = data_i[5387] & sel_one_hot_i[42];
  assign data_masked[5386] = data_i[5386] & sel_one_hot_i[42];
  assign data_masked[5385] = data_i[5385] & sel_one_hot_i[42];
  assign data_masked[5384] = data_i[5384] & sel_one_hot_i[42];
  assign data_masked[5383] = data_i[5383] & sel_one_hot_i[42];
  assign data_masked[5382] = data_i[5382] & sel_one_hot_i[42];
  assign data_masked[5381] = data_i[5381] & sel_one_hot_i[42];
  assign data_masked[5380] = data_i[5380] & sel_one_hot_i[42];
  assign data_masked[5379] = data_i[5379] & sel_one_hot_i[42];
  assign data_masked[5378] = data_i[5378] & sel_one_hot_i[42];
  assign data_masked[5377] = data_i[5377] & sel_one_hot_i[42];
  assign data_masked[5376] = data_i[5376] & sel_one_hot_i[42];
  assign data_masked[5631] = data_i[5631] & sel_one_hot_i[43];
  assign data_masked[5630] = data_i[5630] & sel_one_hot_i[43];
  assign data_masked[5629] = data_i[5629] & sel_one_hot_i[43];
  assign data_masked[5628] = data_i[5628] & sel_one_hot_i[43];
  assign data_masked[5627] = data_i[5627] & sel_one_hot_i[43];
  assign data_masked[5626] = data_i[5626] & sel_one_hot_i[43];
  assign data_masked[5625] = data_i[5625] & sel_one_hot_i[43];
  assign data_masked[5624] = data_i[5624] & sel_one_hot_i[43];
  assign data_masked[5623] = data_i[5623] & sel_one_hot_i[43];
  assign data_masked[5622] = data_i[5622] & sel_one_hot_i[43];
  assign data_masked[5621] = data_i[5621] & sel_one_hot_i[43];
  assign data_masked[5620] = data_i[5620] & sel_one_hot_i[43];
  assign data_masked[5619] = data_i[5619] & sel_one_hot_i[43];
  assign data_masked[5618] = data_i[5618] & sel_one_hot_i[43];
  assign data_masked[5617] = data_i[5617] & sel_one_hot_i[43];
  assign data_masked[5616] = data_i[5616] & sel_one_hot_i[43];
  assign data_masked[5615] = data_i[5615] & sel_one_hot_i[43];
  assign data_masked[5614] = data_i[5614] & sel_one_hot_i[43];
  assign data_masked[5613] = data_i[5613] & sel_one_hot_i[43];
  assign data_masked[5612] = data_i[5612] & sel_one_hot_i[43];
  assign data_masked[5611] = data_i[5611] & sel_one_hot_i[43];
  assign data_masked[5610] = data_i[5610] & sel_one_hot_i[43];
  assign data_masked[5609] = data_i[5609] & sel_one_hot_i[43];
  assign data_masked[5608] = data_i[5608] & sel_one_hot_i[43];
  assign data_masked[5607] = data_i[5607] & sel_one_hot_i[43];
  assign data_masked[5606] = data_i[5606] & sel_one_hot_i[43];
  assign data_masked[5605] = data_i[5605] & sel_one_hot_i[43];
  assign data_masked[5604] = data_i[5604] & sel_one_hot_i[43];
  assign data_masked[5603] = data_i[5603] & sel_one_hot_i[43];
  assign data_masked[5602] = data_i[5602] & sel_one_hot_i[43];
  assign data_masked[5601] = data_i[5601] & sel_one_hot_i[43];
  assign data_masked[5600] = data_i[5600] & sel_one_hot_i[43];
  assign data_masked[5599] = data_i[5599] & sel_one_hot_i[43];
  assign data_masked[5598] = data_i[5598] & sel_one_hot_i[43];
  assign data_masked[5597] = data_i[5597] & sel_one_hot_i[43];
  assign data_masked[5596] = data_i[5596] & sel_one_hot_i[43];
  assign data_masked[5595] = data_i[5595] & sel_one_hot_i[43];
  assign data_masked[5594] = data_i[5594] & sel_one_hot_i[43];
  assign data_masked[5593] = data_i[5593] & sel_one_hot_i[43];
  assign data_masked[5592] = data_i[5592] & sel_one_hot_i[43];
  assign data_masked[5591] = data_i[5591] & sel_one_hot_i[43];
  assign data_masked[5590] = data_i[5590] & sel_one_hot_i[43];
  assign data_masked[5589] = data_i[5589] & sel_one_hot_i[43];
  assign data_masked[5588] = data_i[5588] & sel_one_hot_i[43];
  assign data_masked[5587] = data_i[5587] & sel_one_hot_i[43];
  assign data_masked[5586] = data_i[5586] & sel_one_hot_i[43];
  assign data_masked[5585] = data_i[5585] & sel_one_hot_i[43];
  assign data_masked[5584] = data_i[5584] & sel_one_hot_i[43];
  assign data_masked[5583] = data_i[5583] & sel_one_hot_i[43];
  assign data_masked[5582] = data_i[5582] & sel_one_hot_i[43];
  assign data_masked[5581] = data_i[5581] & sel_one_hot_i[43];
  assign data_masked[5580] = data_i[5580] & sel_one_hot_i[43];
  assign data_masked[5579] = data_i[5579] & sel_one_hot_i[43];
  assign data_masked[5578] = data_i[5578] & sel_one_hot_i[43];
  assign data_masked[5577] = data_i[5577] & sel_one_hot_i[43];
  assign data_masked[5576] = data_i[5576] & sel_one_hot_i[43];
  assign data_masked[5575] = data_i[5575] & sel_one_hot_i[43];
  assign data_masked[5574] = data_i[5574] & sel_one_hot_i[43];
  assign data_masked[5573] = data_i[5573] & sel_one_hot_i[43];
  assign data_masked[5572] = data_i[5572] & sel_one_hot_i[43];
  assign data_masked[5571] = data_i[5571] & sel_one_hot_i[43];
  assign data_masked[5570] = data_i[5570] & sel_one_hot_i[43];
  assign data_masked[5569] = data_i[5569] & sel_one_hot_i[43];
  assign data_masked[5568] = data_i[5568] & sel_one_hot_i[43];
  assign data_masked[5567] = data_i[5567] & sel_one_hot_i[43];
  assign data_masked[5566] = data_i[5566] & sel_one_hot_i[43];
  assign data_masked[5565] = data_i[5565] & sel_one_hot_i[43];
  assign data_masked[5564] = data_i[5564] & sel_one_hot_i[43];
  assign data_masked[5563] = data_i[5563] & sel_one_hot_i[43];
  assign data_masked[5562] = data_i[5562] & sel_one_hot_i[43];
  assign data_masked[5561] = data_i[5561] & sel_one_hot_i[43];
  assign data_masked[5560] = data_i[5560] & sel_one_hot_i[43];
  assign data_masked[5559] = data_i[5559] & sel_one_hot_i[43];
  assign data_masked[5558] = data_i[5558] & sel_one_hot_i[43];
  assign data_masked[5557] = data_i[5557] & sel_one_hot_i[43];
  assign data_masked[5556] = data_i[5556] & sel_one_hot_i[43];
  assign data_masked[5555] = data_i[5555] & sel_one_hot_i[43];
  assign data_masked[5554] = data_i[5554] & sel_one_hot_i[43];
  assign data_masked[5553] = data_i[5553] & sel_one_hot_i[43];
  assign data_masked[5552] = data_i[5552] & sel_one_hot_i[43];
  assign data_masked[5551] = data_i[5551] & sel_one_hot_i[43];
  assign data_masked[5550] = data_i[5550] & sel_one_hot_i[43];
  assign data_masked[5549] = data_i[5549] & sel_one_hot_i[43];
  assign data_masked[5548] = data_i[5548] & sel_one_hot_i[43];
  assign data_masked[5547] = data_i[5547] & sel_one_hot_i[43];
  assign data_masked[5546] = data_i[5546] & sel_one_hot_i[43];
  assign data_masked[5545] = data_i[5545] & sel_one_hot_i[43];
  assign data_masked[5544] = data_i[5544] & sel_one_hot_i[43];
  assign data_masked[5543] = data_i[5543] & sel_one_hot_i[43];
  assign data_masked[5542] = data_i[5542] & sel_one_hot_i[43];
  assign data_masked[5541] = data_i[5541] & sel_one_hot_i[43];
  assign data_masked[5540] = data_i[5540] & sel_one_hot_i[43];
  assign data_masked[5539] = data_i[5539] & sel_one_hot_i[43];
  assign data_masked[5538] = data_i[5538] & sel_one_hot_i[43];
  assign data_masked[5537] = data_i[5537] & sel_one_hot_i[43];
  assign data_masked[5536] = data_i[5536] & sel_one_hot_i[43];
  assign data_masked[5535] = data_i[5535] & sel_one_hot_i[43];
  assign data_masked[5534] = data_i[5534] & sel_one_hot_i[43];
  assign data_masked[5533] = data_i[5533] & sel_one_hot_i[43];
  assign data_masked[5532] = data_i[5532] & sel_one_hot_i[43];
  assign data_masked[5531] = data_i[5531] & sel_one_hot_i[43];
  assign data_masked[5530] = data_i[5530] & sel_one_hot_i[43];
  assign data_masked[5529] = data_i[5529] & sel_one_hot_i[43];
  assign data_masked[5528] = data_i[5528] & sel_one_hot_i[43];
  assign data_masked[5527] = data_i[5527] & sel_one_hot_i[43];
  assign data_masked[5526] = data_i[5526] & sel_one_hot_i[43];
  assign data_masked[5525] = data_i[5525] & sel_one_hot_i[43];
  assign data_masked[5524] = data_i[5524] & sel_one_hot_i[43];
  assign data_masked[5523] = data_i[5523] & sel_one_hot_i[43];
  assign data_masked[5522] = data_i[5522] & sel_one_hot_i[43];
  assign data_masked[5521] = data_i[5521] & sel_one_hot_i[43];
  assign data_masked[5520] = data_i[5520] & sel_one_hot_i[43];
  assign data_masked[5519] = data_i[5519] & sel_one_hot_i[43];
  assign data_masked[5518] = data_i[5518] & sel_one_hot_i[43];
  assign data_masked[5517] = data_i[5517] & sel_one_hot_i[43];
  assign data_masked[5516] = data_i[5516] & sel_one_hot_i[43];
  assign data_masked[5515] = data_i[5515] & sel_one_hot_i[43];
  assign data_masked[5514] = data_i[5514] & sel_one_hot_i[43];
  assign data_masked[5513] = data_i[5513] & sel_one_hot_i[43];
  assign data_masked[5512] = data_i[5512] & sel_one_hot_i[43];
  assign data_masked[5511] = data_i[5511] & sel_one_hot_i[43];
  assign data_masked[5510] = data_i[5510] & sel_one_hot_i[43];
  assign data_masked[5509] = data_i[5509] & sel_one_hot_i[43];
  assign data_masked[5508] = data_i[5508] & sel_one_hot_i[43];
  assign data_masked[5507] = data_i[5507] & sel_one_hot_i[43];
  assign data_masked[5506] = data_i[5506] & sel_one_hot_i[43];
  assign data_masked[5505] = data_i[5505] & sel_one_hot_i[43];
  assign data_masked[5504] = data_i[5504] & sel_one_hot_i[43];
  assign data_masked[5759] = data_i[5759] & sel_one_hot_i[44];
  assign data_masked[5758] = data_i[5758] & sel_one_hot_i[44];
  assign data_masked[5757] = data_i[5757] & sel_one_hot_i[44];
  assign data_masked[5756] = data_i[5756] & sel_one_hot_i[44];
  assign data_masked[5755] = data_i[5755] & sel_one_hot_i[44];
  assign data_masked[5754] = data_i[5754] & sel_one_hot_i[44];
  assign data_masked[5753] = data_i[5753] & sel_one_hot_i[44];
  assign data_masked[5752] = data_i[5752] & sel_one_hot_i[44];
  assign data_masked[5751] = data_i[5751] & sel_one_hot_i[44];
  assign data_masked[5750] = data_i[5750] & sel_one_hot_i[44];
  assign data_masked[5749] = data_i[5749] & sel_one_hot_i[44];
  assign data_masked[5748] = data_i[5748] & sel_one_hot_i[44];
  assign data_masked[5747] = data_i[5747] & sel_one_hot_i[44];
  assign data_masked[5746] = data_i[5746] & sel_one_hot_i[44];
  assign data_masked[5745] = data_i[5745] & sel_one_hot_i[44];
  assign data_masked[5744] = data_i[5744] & sel_one_hot_i[44];
  assign data_masked[5743] = data_i[5743] & sel_one_hot_i[44];
  assign data_masked[5742] = data_i[5742] & sel_one_hot_i[44];
  assign data_masked[5741] = data_i[5741] & sel_one_hot_i[44];
  assign data_masked[5740] = data_i[5740] & sel_one_hot_i[44];
  assign data_masked[5739] = data_i[5739] & sel_one_hot_i[44];
  assign data_masked[5738] = data_i[5738] & sel_one_hot_i[44];
  assign data_masked[5737] = data_i[5737] & sel_one_hot_i[44];
  assign data_masked[5736] = data_i[5736] & sel_one_hot_i[44];
  assign data_masked[5735] = data_i[5735] & sel_one_hot_i[44];
  assign data_masked[5734] = data_i[5734] & sel_one_hot_i[44];
  assign data_masked[5733] = data_i[5733] & sel_one_hot_i[44];
  assign data_masked[5732] = data_i[5732] & sel_one_hot_i[44];
  assign data_masked[5731] = data_i[5731] & sel_one_hot_i[44];
  assign data_masked[5730] = data_i[5730] & sel_one_hot_i[44];
  assign data_masked[5729] = data_i[5729] & sel_one_hot_i[44];
  assign data_masked[5728] = data_i[5728] & sel_one_hot_i[44];
  assign data_masked[5727] = data_i[5727] & sel_one_hot_i[44];
  assign data_masked[5726] = data_i[5726] & sel_one_hot_i[44];
  assign data_masked[5725] = data_i[5725] & sel_one_hot_i[44];
  assign data_masked[5724] = data_i[5724] & sel_one_hot_i[44];
  assign data_masked[5723] = data_i[5723] & sel_one_hot_i[44];
  assign data_masked[5722] = data_i[5722] & sel_one_hot_i[44];
  assign data_masked[5721] = data_i[5721] & sel_one_hot_i[44];
  assign data_masked[5720] = data_i[5720] & sel_one_hot_i[44];
  assign data_masked[5719] = data_i[5719] & sel_one_hot_i[44];
  assign data_masked[5718] = data_i[5718] & sel_one_hot_i[44];
  assign data_masked[5717] = data_i[5717] & sel_one_hot_i[44];
  assign data_masked[5716] = data_i[5716] & sel_one_hot_i[44];
  assign data_masked[5715] = data_i[5715] & sel_one_hot_i[44];
  assign data_masked[5714] = data_i[5714] & sel_one_hot_i[44];
  assign data_masked[5713] = data_i[5713] & sel_one_hot_i[44];
  assign data_masked[5712] = data_i[5712] & sel_one_hot_i[44];
  assign data_masked[5711] = data_i[5711] & sel_one_hot_i[44];
  assign data_masked[5710] = data_i[5710] & sel_one_hot_i[44];
  assign data_masked[5709] = data_i[5709] & sel_one_hot_i[44];
  assign data_masked[5708] = data_i[5708] & sel_one_hot_i[44];
  assign data_masked[5707] = data_i[5707] & sel_one_hot_i[44];
  assign data_masked[5706] = data_i[5706] & sel_one_hot_i[44];
  assign data_masked[5705] = data_i[5705] & sel_one_hot_i[44];
  assign data_masked[5704] = data_i[5704] & sel_one_hot_i[44];
  assign data_masked[5703] = data_i[5703] & sel_one_hot_i[44];
  assign data_masked[5702] = data_i[5702] & sel_one_hot_i[44];
  assign data_masked[5701] = data_i[5701] & sel_one_hot_i[44];
  assign data_masked[5700] = data_i[5700] & sel_one_hot_i[44];
  assign data_masked[5699] = data_i[5699] & sel_one_hot_i[44];
  assign data_masked[5698] = data_i[5698] & sel_one_hot_i[44];
  assign data_masked[5697] = data_i[5697] & sel_one_hot_i[44];
  assign data_masked[5696] = data_i[5696] & sel_one_hot_i[44];
  assign data_masked[5695] = data_i[5695] & sel_one_hot_i[44];
  assign data_masked[5694] = data_i[5694] & sel_one_hot_i[44];
  assign data_masked[5693] = data_i[5693] & sel_one_hot_i[44];
  assign data_masked[5692] = data_i[5692] & sel_one_hot_i[44];
  assign data_masked[5691] = data_i[5691] & sel_one_hot_i[44];
  assign data_masked[5690] = data_i[5690] & sel_one_hot_i[44];
  assign data_masked[5689] = data_i[5689] & sel_one_hot_i[44];
  assign data_masked[5688] = data_i[5688] & sel_one_hot_i[44];
  assign data_masked[5687] = data_i[5687] & sel_one_hot_i[44];
  assign data_masked[5686] = data_i[5686] & sel_one_hot_i[44];
  assign data_masked[5685] = data_i[5685] & sel_one_hot_i[44];
  assign data_masked[5684] = data_i[5684] & sel_one_hot_i[44];
  assign data_masked[5683] = data_i[5683] & sel_one_hot_i[44];
  assign data_masked[5682] = data_i[5682] & sel_one_hot_i[44];
  assign data_masked[5681] = data_i[5681] & sel_one_hot_i[44];
  assign data_masked[5680] = data_i[5680] & sel_one_hot_i[44];
  assign data_masked[5679] = data_i[5679] & sel_one_hot_i[44];
  assign data_masked[5678] = data_i[5678] & sel_one_hot_i[44];
  assign data_masked[5677] = data_i[5677] & sel_one_hot_i[44];
  assign data_masked[5676] = data_i[5676] & sel_one_hot_i[44];
  assign data_masked[5675] = data_i[5675] & sel_one_hot_i[44];
  assign data_masked[5674] = data_i[5674] & sel_one_hot_i[44];
  assign data_masked[5673] = data_i[5673] & sel_one_hot_i[44];
  assign data_masked[5672] = data_i[5672] & sel_one_hot_i[44];
  assign data_masked[5671] = data_i[5671] & sel_one_hot_i[44];
  assign data_masked[5670] = data_i[5670] & sel_one_hot_i[44];
  assign data_masked[5669] = data_i[5669] & sel_one_hot_i[44];
  assign data_masked[5668] = data_i[5668] & sel_one_hot_i[44];
  assign data_masked[5667] = data_i[5667] & sel_one_hot_i[44];
  assign data_masked[5666] = data_i[5666] & sel_one_hot_i[44];
  assign data_masked[5665] = data_i[5665] & sel_one_hot_i[44];
  assign data_masked[5664] = data_i[5664] & sel_one_hot_i[44];
  assign data_masked[5663] = data_i[5663] & sel_one_hot_i[44];
  assign data_masked[5662] = data_i[5662] & sel_one_hot_i[44];
  assign data_masked[5661] = data_i[5661] & sel_one_hot_i[44];
  assign data_masked[5660] = data_i[5660] & sel_one_hot_i[44];
  assign data_masked[5659] = data_i[5659] & sel_one_hot_i[44];
  assign data_masked[5658] = data_i[5658] & sel_one_hot_i[44];
  assign data_masked[5657] = data_i[5657] & sel_one_hot_i[44];
  assign data_masked[5656] = data_i[5656] & sel_one_hot_i[44];
  assign data_masked[5655] = data_i[5655] & sel_one_hot_i[44];
  assign data_masked[5654] = data_i[5654] & sel_one_hot_i[44];
  assign data_masked[5653] = data_i[5653] & sel_one_hot_i[44];
  assign data_masked[5652] = data_i[5652] & sel_one_hot_i[44];
  assign data_masked[5651] = data_i[5651] & sel_one_hot_i[44];
  assign data_masked[5650] = data_i[5650] & sel_one_hot_i[44];
  assign data_masked[5649] = data_i[5649] & sel_one_hot_i[44];
  assign data_masked[5648] = data_i[5648] & sel_one_hot_i[44];
  assign data_masked[5647] = data_i[5647] & sel_one_hot_i[44];
  assign data_masked[5646] = data_i[5646] & sel_one_hot_i[44];
  assign data_masked[5645] = data_i[5645] & sel_one_hot_i[44];
  assign data_masked[5644] = data_i[5644] & sel_one_hot_i[44];
  assign data_masked[5643] = data_i[5643] & sel_one_hot_i[44];
  assign data_masked[5642] = data_i[5642] & sel_one_hot_i[44];
  assign data_masked[5641] = data_i[5641] & sel_one_hot_i[44];
  assign data_masked[5640] = data_i[5640] & sel_one_hot_i[44];
  assign data_masked[5639] = data_i[5639] & sel_one_hot_i[44];
  assign data_masked[5638] = data_i[5638] & sel_one_hot_i[44];
  assign data_masked[5637] = data_i[5637] & sel_one_hot_i[44];
  assign data_masked[5636] = data_i[5636] & sel_one_hot_i[44];
  assign data_masked[5635] = data_i[5635] & sel_one_hot_i[44];
  assign data_masked[5634] = data_i[5634] & sel_one_hot_i[44];
  assign data_masked[5633] = data_i[5633] & sel_one_hot_i[44];
  assign data_masked[5632] = data_i[5632] & sel_one_hot_i[44];
  assign data_masked[5887] = data_i[5887] & sel_one_hot_i[45];
  assign data_masked[5886] = data_i[5886] & sel_one_hot_i[45];
  assign data_masked[5885] = data_i[5885] & sel_one_hot_i[45];
  assign data_masked[5884] = data_i[5884] & sel_one_hot_i[45];
  assign data_masked[5883] = data_i[5883] & sel_one_hot_i[45];
  assign data_masked[5882] = data_i[5882] & sel_one_hot_i[45];
  assign data_masked[5881] = data_i[5881] & sel_one_hot_i[45];
  assign data_masked[5880] = data_i[5880] & sel_one_hot_i[45];
  assign data_masked[5879] = data_i[5879] & sel_one_hot_i[45];
  assign data_masked[5878] = data_i[5878] & sel_one_hot_i[45];
  assign data_masked[5877] = data_i[5877] & sel_one_hot_i[45];
  assign data_masked[5876] = data_i[5876] & sel_one_hot_i[45];
  assign data_masked[5875] = data_i[5875] & sel_one_hot_i[45];
  assign data_masked[5874] = data_i[5874] & sel_one_hot_i[45];
  assign data_masked[5873] = data_i[5873] & sel_one_hot_i[45];
  assign data_masked[5872] = data_i[5872] & sel_one_hot_i[45];
  assign data_masked[5871] = data_i[5871] & sel_one_hot_i[45];
  assign data_masked[5870] = data_i[5870] & sel_one_hot_i[45];
  assign data_masked[5869] = data_i[5869] & sel_one_hot_i[45];
  assign data_masked[5868] = data_i[5868] & sel_one_hot_i[45];
  assign data_masked[5867] = data_i[5867] & sel_one_hot_i[45];
  assign data_masked[5866] = data_i[5866] & sel_one_hot_i[45];
  assign data_masked[5865] = data_i[5865] & sel_one_hot_i[45];
  assign data_masked[5864] = data_i[5864] & sel_one_hot_i[45];
  assign data_masked[5863] = data_i[5863] & sel_one_hot_i[45];
  assign data_masked[5862] = data_i[5862] & sel_one_hot_i[45];
  assign data_masked[5861] = data_i[5861] & sel_one_hot_i[45];
  assign data_masked[5860] = data_i[5860] & sel_one_hot_i[45];
  assign data_masked[5859] = data_i[5859] & sel_one_hot_i[45];
  assign data_masked[5858] = data_i[5858] & sel_one_hot_i[45];
  assign data_masked[5857] = data_i[5857] & sel_one_hot_i[45];
  assign data_masked[5856] = data_i[5856] & sel_one_hot_i[45];
  assign data_masked[5855] = data_i[5855] & sel_one_hot_i[45];
  assign data_masked[5854] = data_i[5854] & sel_one_hot_i[45];
  assign data_masked[5853] = data_i[5853] & sel_one_hot_i[45];
  assign data_masked[5852] = data_i[5852] & sel_one_hot_i[45];
  assign data_masked[5851] = data_i[5851] & sel_one_hot_i[45];
  assign data_masked[5850] = data_i[5850] & sel_one_hot_i[45];
  assign data_masked[5849] = data_i[5849] & sel_one_hot_i[45];
  assign data_masked[5848] = data_i[5848] & sel_one_hot_i[45];
  assign data_masked[5847] = data_i[5847] & sel_one_hot_i[45];
  assign data_masked[5846] = data_i[5846] & sel_one_hot_i[45];
  assign data_masked[5845] = data_i[5845] & sel_one_hot_i[45];
  assign data_masked[5844] = data_i[5844] & sel_one_hot_i[45];
  assign data_masked[5843] = data_i[5843] & sel_one_hot_i[45];
  assign data_masked[5842] = data_i[5842] & sel_one_hot_i[45];
  assign data_masked[5841] = data_i[5841] & sel_one_hot_i[45];
  assign data_masked[5840] = data_i[5840] & sel_one_hot_i[45];
  assign data_masked[5839] = data_i[5839] & sel_one_hot_i[45];
  assign data_masked[5838] = data_i[5838] & sel_one_hot_i[45];
  assign data_masked[5837] = data_i[5837] & sel_one_hot_i[45];
  assign data_masked[5836] = data_i[5836] & sel_one_hot_i[45];
  assign data_masked[5835] = data_i[5835] & sel_one_hot_i[45];
  assign data_masked[5834] = data_i[5834] & sel_one_hot_i[45];
  assign data_masked[5833] = data_i[5833] & sel_one_hot_i[45];
  assign data_masked[5832] = data_i[5832] & sel_one_hot_i[45];
  assign data_masked[5831] = data_i[5831] & sel_one_hot_i[45];
  assign data_masked[5830] = data_i[5830] & sel_one_hot_i[45];
  assign data_masked[5829] = data_i[5829] & sel_one_hot_i[45];
  assign data_masked[5828] = data_i[5828] & sel_one_hot_i[45];
  assign data_masked[5827] = data_i[5827] & sel_one_hot_i[45];
  assign data_masked[5826] = data_i[5826] & sel_one_hot_i[45];
  assign data_masked[5825] = data_i[5825] & sel_one_hot_i[45];
  assign data_masked[5824] = data_i[5824] & sel_one_hot_i[45];
  assign data_masked[5823] = data_i[5823] & sel_one_hot_i[45];
  assign data_masked[5822] = data_i[5822] & sel_one_hot_i[45];
  assign data_masked[5821] = data_i[5821] & sel_one_hot_i[45];
  assign data_masked[5820] = data_i[5820] & sel_one_hot_i[45];
  assign data_masked[5819] = data_i[5819] & sel_one_hot_i[45];
  assign data_masked[5818] = data_i[5818] & sel_one_hot_i[45];
  assign data_masked[5817] = data_i[5817] & sel_one_hot_i[45];
  assign data_masked[5816] = data_i[5816] & sel_one_hot_i[45];
  assign data_masked[5815] = data_i[5815] & sel_one_hot_i[45];
  assign data_masked[5814] = data_i[5814] & sel_one_hot_i[45];
  assign data_masked[5813] = data_i[5813] & sel_one_hot_i[45];
  assign data_masked[5812] = data_i[5812] & sel_one_hot_i[45];
  assign data_masked[5811] = data_i[5811] & sel_one_hot_i[45];
  assign data_masked[5810] = data_i[5810] & sel_one_hot_i[45];
  assign data_masked[5809] = data_i[5809] & sel_one_hot_i[45];
  assign data_masked[5808] = data_i[5808] & sel_one_hot_i[45];
  assign data_masked[5807] = data_i[5807] & sel_one_hot_i[45];
  assign data_masked[5806] = data_i[5806] & sel_one_hot_i[45];
  assign data_masked[5805] = data_i[5805] & sel_one_hot_i[45];
  assign data_masked[5804] = data_i[5804] & sel_one_hot_i[45];
  assign data_masked[5803] = data_i[5803] & sel_one_hot_i[45];
  assign data_masked[5802] = data_i[5802] & sel_one_hot_i[45];
  assign data_masked[5801] = data_i[5801] & sel_one_hot_i[45];
  assign data_masked[5800] = data_i[5800] & sel_one_hot_i[45];
  assign data_masked[5799] = data_i[5799] & sel_one_hot_i[45];
  assign data_masked[5798] = data_i[5798] & sel_one_hot_i[45];
  assign data_masked[5797] = data_i[5797] & sel_one_hot_i[45];
  assign data_masked[5796] = data_i[5796] & sel_one_hot_i[45];
  assign data_masked[5795] = data_i[5795] & sel_one_hot_i[45];
  assign data_masked[5794] = data_i[5794] & sel_one_hot_i[45];
  assign data_masked[5793] = data_i[5793] & sel_one_hot_i[45];
  assign data_masked[5792] = data_i[5792] & sel_one_hot_i[45];
  assign data_masked[5791] = data_i[5791] & sel_one_hot_i[45];
  assign data_masked[5790] = data_i[5790] & sel_one_hot_i[45];
  assign data_masked[5789] = data_i[5789] & sel_one_hot_i[45];
  assign data_masked[5788] = data_i[5788] & sel_one_hot_i[45];
  assign data_masked[5787] = data_i[5787] & sel_one_hot_i[45];
  assign data_masked[5786] = data_i[5786] & sel_one_hot_i[45];
  assign data_masked[5785] = data_i[5785] & sel_one_hot_i[45];
  assign data_masked[5784] = data_i[5784] & sel_one_hot_i[45];
  assign data_masked[5783] = data_i[5783] & sel_one_hot_i[45];
  assign data_masked[5782] = data_i[5782] & sel_one_hot_i[45];
  assign data_masked[5781] = data_i[5781] & sel_one_hot_i[45];
  assign data_masked[5780] = data_i[5780] & sel_one_hot_i[45];
  assign data_masked[5779] = data_i[5779] & sel_one_hot_i[45];
  assign data_masked[5778] = data_i[5778] & sel_one_hot_i[45];
  assign data_masked[5777] = data_i[5777] & sel_one_hot_i[45];
  assign data_masked[5776] = data_i[5776] & sel_one_hot_i[45];
  assign data_masked[5775] = data_i[5775] & sel_one_hot_i[45];
  assign data_masked[5774] = data_i[5774] & sel_one_hot_i[45];
  assign data_masked[5773] = data_i[5773] & sel_one_hot_i[45];
  assign data_masked[5772] = data_i[5772] & sel_one_hot_i[45];
  assign data_masked[5771] = data_i[5771] & sel_one_hot_i[45];
  assign data_masked[5770] = data_i[5770] & sel_one_hot_i[45];
  assign data_masked[5769] = data_i[5769] & sel_one_hot_i[45];
  assign data_masked[5768] = data_i[5768] & sel_one_hot_i[45];
  assign data_masked[5767] = data_i[5767] & sel_one_hot_i[45];
  assign data_masked[5766] = data_i[5766] & sel_one_hot_i[45];
  assign data_masked[5765] = data_i[5765] & sel_one_hot_i[45];
  assign data_masked[5764] = data_i[5764] & sel_one_hot_i[45];
  assign data_masked[5763] = data_i[5763] & sel_one_hot_i[45];
  assign data_masked[5762] = data_i[5762] & sel_one_hot_i[45];
  assign data_masked[5761] = data_i[5761] & sel_one_hot_i[45];
  assign data_masked[5760] = data_i[5760] & sel_one_hot_i[45];
  assign data_masked[6015] = data_i[6015] & sel_one_hot_i[46];
  assign data_masked[6014] = data_i[6014] & sel_one_hot_i[46];
  assign data_masked[6013] = data_i[6013] & sel_one_hot_i[46];
  assign data_masked[6012] = data_i[6012] & sel_one_hot_i[46];
  assign data_masked[6011] = data_i[6011] & sel_one_hot_i[46];
  assign data_masked[6010] = data_i[6010] & sel_one_hot_i[46];
  assign data_masked[6009] = data_i[6009] & sel_one_hot_i[46];
  assign data_masked[6008] = data_i[6008] & sel_one_hot_i[46];
  assign data_masked[6007] = data_i[6007] & sel_one_hot_i[46];
  assign data_masked[6006] = data_i[6006] & sel_one_hot_i[46];
  assign data_masked[6005] = data_i[6005] & sel_one_hot_i[46];
  assign data_masked[6004] = data_i[6004] & sel_one_hot_i[46];
  assign data_masked[6003] = data_i[6003] & sel_one_hot_i[46];
  assign data_masked[6002] = data_i[6002] & sel_one_hot_i[46];
  assign data_masked[6001] = data_i[6001] & sel_one_hot_i[46];
  assign data_masked[6000] = data_i[6000] & sel_one_hot_i[46];
  assign data_masked[5999] = data_i[5999] & sel_one_hot_i[46];
  assign data_masked[5998] = data_i[5998] & sel_one_hot_i[46];
  assign data_masked[5997] = data_i[5997] & sel_one_hot_i[46];
  assign data_masked[5996] = data_i[5996] & sel_one_hot_i[46];
  assign data_masked[5995] = data_i[5995] & sel_one_hot_i[46];
  assign data_masked[5994] = data_i[5994] & sel_one_hot_i[46];
  assign data_masked[5993] = data_i[5993] & sel_one_hot_i[46];
  assign data_masked[5992] = data_i[5992] & sel_one_hot_i[46];
  assign data_masked[5991] = data_i[5991] & sel_one_hot_i[46];
  assign data_masked[5990] = data_i[5990] & sel_one_hot_i[46];
  assign data_masked[5989] = data_i[5989] & sel_one_hot_i[46];
  assign data_masked[5988] = data_i[5988] & sel_one_hot_i[46];
  assign data_masked[5987] = data_i[5987] & sel_one_hot_i[46];
  assign data_masked[5986] = data_i[5986] & sel_one_hot_i[46];
  assign data_masked[5985] = data_i[5985] & sel_one_hot_i[46];
  assign data_masked[5984] = data_i[5984] & sel_one_hot_i[46];
  assign data_masked[5983] = data_i[5983] & sel_one_hot_i[46];
  assign data_masked[5982] = data_i[5982] & sel_one_hot_i[46];
  assign data_masked[5981] = data_i[5981] & sel_one_hot_i[46];
  assign data_masked[5980] = data_i[5980] & sel_one_hot_i[46];
  assign data_masked[5979] = data_i[5979] & sel_one_hot_i[46];
  assign data_masked[5978] = data_i[5978] & sel_one_hot_i[46];
  assign data_masked[5977] = data_i[5977] & sel_one_hot_i[46];
  assign data_masked[5976] = data_i[5976] & sel_one_hot_i[46];
  assign data_masked[5975] = data_i[5975] & sel_one_hot_i[46];
  assign data_masked[5974] = data_i[5974] & sel_one_hot_i[46];
  assign data_masked[5973] = data_i[5973] & sel_one_hot_i[46];
  assign data_masked[5972] = data_i[5972] & sel_one_hot_i[46];
  assign data_masked[5971] = data_i[5971] & sel_one_hot_i[46];
  assign data_masked[5970] = data_i[5970] & sel_one_hot_i[46];
  assign data_masked[5969] = data_i[5969] & sel_one_hot_i[46];
  assign data_masked[5968] = data_i[5968] & sel_one_hot_i[46];
  assign data_masked[5967] = data_i[5967] & sel_one_hot_i[46];
  assign data_masked[5966] = data_i[5966] & sel_one_hot_i[46];
  assign data_masked[5965] = data_i[5965] & sel_one_hot_i[46];
  assign data_masked[5964] = data_i[5964] & sel_one_hot_i[46];
  assign data_masked[5963] = data_i[5963] & sel_one_hot_i[46];
  assign data_masked[5962] = data_i[5962] & sel_one_hot_i[46];
  assign data_masked[5961] = data_i[5961] & sel_one_hot_i[46];
  assign data_masked[5960] = data_i[5960] & sel_one_hot_i[46];
  assign data_masked[5959] = data_i[5959] & sel_one_hot_i[46];
  assign data_masked[5958] = data_i[5958] & sel_one_hot_i[46];
  assign data_masked[5957] = data_i[5957] & sel_one_hot_i[46];
  assign data_masked[5956] = data_i[5956] & sel_one_hot_i[46];
  assign data_masked[5955] = data_i[5955] & sel_one_hot_i[46];
  assign data_masked[5954] = data_i[5954] & sel_one_hot_i[46];
  assign data_masked[5953] = data_i[5953] & sel_one_hot_i[46];
  assign data_masked[5952] = data_i[5952] & sel_one_hot_i[46];
  assign data_masked[5951] = data_i[5951] & sel_one_hot_i[46];
  assign data_masked[5950] = data_i[5950] & sel_one_hot_i[46];
  assign data_masked[5949] = data_i[5949] & sel_one_hot_i[46];
  assign data_masked[5948] = data_i[5948] & sel_one_hot_i[46];
  assign data_masked[5947] = data_i[5947] & sel_one_hot_i[46];
  assign data_masked[5946] = data_i[5946] & sel_one_hot_i[46];
  assign data_masked[5945] = data_i[5945] & sel_one_hot_i[46];
  assign data_masked[5944] = data_i[5944] & sel_one_hot_i[46];
  assign data_masked[5943] = data_i[5943] & sel_one_hot_i[46];
  assign data_masked[5942] = data_i[5942] & sel_one_hot_i[46];
  assign data_masked[5941] = data_i[5941] & sel_one_hot_i[46];
  assign data_masked[5940] = data_i[5940] & sel_one_hot_i[46];
  assign data_masked[5939] = data_i[5939] & sel_one_hot_i[46];
  assign data_masked[5938] = data_i[5938] & sel_one_hot_i[46];
  assign data_masked[5937] = data_i[5937] & sel_one_hot_i[46];
  assign data_masked[5936] = data_i[5936] & sel_one_hot_i[46];
  assign data_masked[5935] = data_i[5935] & sel_one_hot_i[46];
  assign data_masked[5934] = data_i[5934] & sel_one_hot_i[46];
  assign data_masked[5933] = data_i[5933] & sel_one_hot_i[46];
  assign data_masked[5932] = data_i[5932] & sel_one_hot_i[46];
  assign data_masked[5931] = data_i[5931] & sel_one_hot_i[46];
  assign data_masked[5930] = data_i[5930] & sel_one_hot_i[46];
  assign data_masked[5929] = data_i[5929] & sel_one_hot_i[46];
  assign data_masked[5928] = data_i[5928] & sel_one_hot_i[46];
  assign data_masked[5927] = data_i[5927] & sel_one_hot_i[46];
  assign data_masked[5926] = data_i[5926] & sel_one_hot_i[46];
  assign data_masked[5925] = data_i[5925] & sel_one_hot_i[46];
  assign data_masked[5924] = data_i[5924] & sel_one_hot_i[46];
  assign data_masked[5923] = data_i[5923] & sel_one_hot_i[46];
  assign data_masked[5922] = data_i[5922] & sel_one_hot_i[46];
  assign data_masked[5921] = data_i[5921] & sel_one_hot_i[46];
  assign data_masked[5920] = data_i[5920] & sel_one_hot_i[46];
  assign data_masked[5919] = data_i[5919] & sel_one_hot_i[46];
  assign data_masked[5918] = data_i[5918] & sel_one_hot_i[46];
  assign data_masked[5917] = data_i[5917] & sel_one_hot_i[46];
  assign data_masked[5916] = data_i[5916] & sel_one_hot_i[46];
  assign data_masked[5915] = data_i[5915] & sel_one_hot_i[46];
  assign data_masked[5914] = data_i[5914] & sel_one_hot_i[46];
  assign data_masked[5913] = data_i[5913] & sel_one_hot_i[46];
  assign data_masked[5912] = data_i[5912] & sel_one_hot_i[46];
  assign data_masked[5911] = data_i[5911] & sel_one_hot_i[46];
  assign data_masked[5910] = data_i[5910] & sel_one_hot_i[46];
  assign data_masked[5909] = data_i[5909] & sel_one_hot_i[46];
  assign data_masked[5908] = data_i[5908] & sel_one_hot_i[46];
  assign data_masked[5907] = data_i[5907] & sel_one_hot_i[46];
  assign data_masked[5906] = data_i[5906] & sel_one_hot_i[46];
  assign data_masked[5905] = data_i[5905] & sel_one_hot_i[46];
  assign data_masked[5904] = data_i[5904] & sel_one_hot_i[46];
  assign data_masked[5903] = data_i[5903] & sel_one_hot_i[46];
  assign data_masked[5902] = data_i[5902] & sel_one_hot_i[46];
  assign data_masked[5901] = data_i[5901] & sel_one_hot_i[46];
  assign data_masked[5900] = data_i[5900] & sel_one_hot_i[46];
  assign data_masked[5899] = data_i[5899] & sel_one_hot_i[46];
  assign data_masked[5898] = data_i[5898] & sel_one_hot_i[46];
  assign data_masked[5897] = data_i[5897] & sel_one_hot_i[46];
  assign data_masked[5896] = data_i[5896] & sel_one_hot_i[46];
  assign data_masked[5895] = data_i[5895] & sel_one_hot_i[46];
  assign data_masked[5894] = data_i[5894] & sel_one_hot_i[46];
  assign data_masked[5893] = data_i[5893] & sel_one_hot_i[46];
  assign data_masked[5892] = data_i[5892] & sel_one_hot_i[46];
  assign data_masked[5891] = data_i[5891] & sel_one_hot_i[46];
  assign data_masked[5890] = data_i[5890] & sel_one_hot_i[46];
  assign data_masked[5889] = data_i[5889] & sel_one_hot_i[46];
  assign data_masked[5888] = data_i[5888] & sel_one_hot_i[46];
  assign data_masked[6143] = data_i[6143] & sel_one_hot_i[47];
  assign data_masked[6142] = data_i[6142] & sel_one_hot_i[47];
  assign data_masked[6141] = data_i[6141] & sel_one_hot_i[47];
  assign data_masked[6140] = data_i[6140] & sel_one_hot_i[47];
  assign data_masked[6139] = data_i[6139] & sel_one_hot_i[47];
  assign data_masked[6138] = data_i[6138] & sel_one_hot_i[47];
  assign data_masked[6137] = data_i[6137] & sel_one_hot_i[47];
  assign data_masked[6136] = data_i[6136] & sel_one_hot_i[47];
  assign data_masked[6135] = data_i[6135] & sel_one_hot_i[47];
  assign data_masked[6134] = data_i[6134] & sel_one_hot_i[47];
  assign data_masked[6133] = data_i[6133] & sel_one_hot_i[47];
  assign data_masked[6132] = data_i[6132] & sel_one_hot_i[47];
  assign data_masked[6131] = data_i[6131] & sel_one_hot_i[47];
  assign data_masked[6130] = data_i[6130] & sel_one_hot_i[47];
  assign data_masked[6129] = data_i[6129] & sel_one_hot_i[47];
  assign data_masked[6128] = data_i[6128] & sel_one_hot_i[47];
  assign data_masked[6127] = data_i[6127] & sel_one_hot_i[47];
  assign data_masked[6126] = data_i[6126] & sel_one_hot_i[47];
  assign data_masked[6125] = data_i[6125] & sel_one_hot_i[47];
  assign data_masked[6124] = data_i[6124] & sel_one_hot_i[47];
  assign data_masked[6123] = data_i[6123] & sel_one_hot_i[47];
  assign data_masked[6122] = data_i[6122] & sel_one_hot_i[47];
  assign data_masked[6121] = data_i[6121] & sel_one_hot_i[47];
  assign data_masked[6120] = data_i[6120] & sel_one_hot_i[47];
  assign data_masked[6119] = data_i[6119] & sel_one_hot_i[47];
  assign data_masked[6118] = data_i[6118] & sel_one_hot_i[47];
  assign data_masked[6117] = data_i[6117] & sel_one_hot_i[47];
  assign data_masked[6116] = data_i[6116] & sel_one_hot_i[47];
  assign data_masked[6115] = data_i[6115] & sel_one_hot_i[47];
  assign data_masked[6114] = data_i[6114] & sel_one_hot_i[47];
  assign data_masked[6113] = data_i[6113] & sel_one_hot_i[47];
  assign data_masked[6112] = data_i[6112] & sel_one_hot_i[47];
  assign data_masked[6111] = data_i[6111] & sel_one_hot_i[47];
  assign data_masked[6110] = data_i[6110] & sel_one_hot_i[47];
  assign data_masked[6109] = data_i[6109] & sel_one_hot_i[47];
  assign data_masked[6108] = data_i[6108] & sel_one_hot_i[47];
  assign data_masked[6107] = data_i[6107] & sel_one_hot_i[47];
  assign data_masked[6106] = data_i[6106] & sel_one_hot_i[47];
  assign data_masked[6105] = data_i[6105] & sel_one_hot_i[47];
  assign data_masked[6104] = data_i[6104] & sel_one_hot_i[47];
  assign data_masked[6103] = data_i[6103] & sel_one_hot_i[47];
  assign data_masked[6102] = data_i[6102] & sel_one_hot_i[47];
  assign data_masked[6101] = data_i[6101] & sel_one_hot_i[47];
  assign data_masked[6100] = data_i[6100] & sel_one_hot_i[47];
  assign data_masked[6099] = data_i[6099] & sel_one_hot_i[47];
  assign data_masked[6098] = data_i[6098] & sel_one_hot_i[47];
  assign data_masked[6097] = data_i[6097] & sel_one_hot_i[47];
  assign data_masked[6096] = data_i[6096] & sel_one_hot_i[47];
  assign data_masked[6095] = data_i[6095] & sel_one_hot_i[47];
  assign data_masked[6094] = data_i[6094] & sel_one_hot_i[47];
  assign data_masked[6093] = data_i[6093] & sel_one_hot_i[47];
  assign data_masked[6092] = data_i[6092] & sel_one_hot_i[47];
  assign data_masked[6091] = data_i[6091] & sel_one_hot_i[47];
  assign data_masked[6090] = data_i[6090] & sel_one_hot_i[47];
  assign data_masked[6089] = data_i[6089] & sel_one_hot_i[47];
  assign data_masked[6088] = data_i[6088] & sel_one_hot_i[47];
  assign data_masked[6087] = data_i[6087] & sel_one_hot_i[47];
  assign data_masked[6086] = data_i[6086] & sel_one_hot_i[47];
  assign data_masked[6085] = data_i[6085] & sel_one_hot_i[47];
  assign data_masked[6084] = data_i[6084] & sel_one_hot_i[47];
  assign data_masked[6083] = data_i[6083] & sel_one_hot_i[47];
  assign data_masked[6082] = data_i[6082] & sel_one_hot_i[47];
  assign data_masked[6081] = data_i[6081] & sel_one_hot_i[47];
  assign data_masked[6080] = data_i[6080] & sel_one_hot_i[47];
  assign data_masked[6079] = data_i[6079] & sel_one_hot_i[47];
  assign data_masked[6078] = data_i[6078] & sel_one_hot_i[47];
  assign data_masked[6077] = data_i[6077] & sel_one_hot_i[47];
  assign data_masked[6076] = data_i[6076] & sel_one_hot_i[47];
  assign data_masked[6075] = data_i[6075] & sel_one_hot_i[47];
  assign data_masked[6074] = data_i[6074] & sel_one_hot_i[47];
  assign data_masked[6073] = data_i[6073] & sel_one_hot_i[47];
  assign data_masked[6072] = data_i[6072] & sel_one_hot_i[47];
  assign data_masked[6071] = data_i[6071] & sel_one_hot_i[47];
  assign data_masked[6070] = data_i[6070] & sel_one_hot_i[47];
  assign data_masked[6069] = data_i[6069] & sel_one_hot_i[47];
  assign data_masked[6068] = data_i[6068] & sel_one_hot_i[47];
  assign data_masked[6067] = data_i[6067] & sel_one_hot_i[47];
  assign data_masked[6066] = data_i[6066] & sel_one_hot_i[47];
  assign data_masked[6065] = data_i[6065] & sel_one_hot_i[47];
  assign data_masked[6064] = data_i[6064] & sel_one_hot_i[47];
  assign data_masked[6063] = data_i[6063] & sel_one_hot_i[47];
  assign data_masked[6062] = data_i[6062] & sel_one_hot_i[47];
  assign data_masked[6061] = data_i[6061] & sel_one_hot_i[47];
  assign data_masked[6060] = data_i[6060] & sel_one_hot_i[47];
  assign data_masked[6059] = data_i[6059] & sel_one_hot_i[47];
  assign data_masked[6058] = data_i[6058] & sel_one_hot_i[47];
  assign data_masked[6057] = data_i[6057] & sel_one_hot_i[47];
  assign data_masked[6056] = data_i[6056] & sel_one_hot_i[47];
  assign data_masked[6055] = data_i[6055] & sel_one_hot_i[47];
  assign data_masked[6054] = data_i[6054] & sel_one_hot_i[47];
  assign data_masked[6053] = data_i[6053] & sel_one_hot_i[47];
  assign data_masked[6052] = data_i[6052] & sel_one_hot_i[47];
  assign data_masked[6051] = data_i[6051] & sel_one_hot_i[47];
  assign data_masked[6050] = data_i[6050] & sel_one_hot_i[47];
  assign data_masked[6049] = data_i[6049] & sel_one_hot_i[47];
  assign data_masked[6048] = data_i[6048] & sel_one_hot_i[47];
  assign data_masked[6047] = data_i[6047] & sel_one_hot_i[47];
  assign data_masked[6046] = data_i[6046] & sel_one_hot_i[47];
  assign data_masked[6045] = data_i[6045] & sel_one_hot_i[47];
  assign data_masked[6044] = data_i[6044] & sel_one_hot_i[47];
  assign data_masked[6043] = data_i[6043] & sel_one_hot_i[47];
  assign data_masked[6042] = data_i[6042] & sel_one_hot_i[47];
  assign data_masked[6041] = data_i[6041] & sel_one_hot_i[47];
  assign data_masked[6040] = data_i[6040] & sel_one_hot_i[47];
  assign data_masked[6039] = data_i[6039] & sel_one_hot_i[47];
  assign data_masked[6038] = data_i[6038] & sel_one_hot_i[47];
  assign data_masked[6037] = data_i[6037] & sel_one_hot_i[47];
  assign data_masked[6036] = data_i[6036] & sel_one_hot_i[47];
  assign data_masked[6035] = data_i[6035] & sel_one_hot_i[47];
  assign data_masked[6034] = data_i[6034] & sel_one_hot_i[47];
  assign data_masked[6033] = data_i[6033] & sel_one_hot_i[47];
  assign data_masked[6032] = data_i[6032] & sel_one_hot_i[47];
  assign data_masked[6031] = data_i[6031] & sel_one_hot_i[47];
  assign data_masked[6030] = data_i[6030] & sel_one_hot_i[47];
  assign data_masked[6029] = data_i[6029] & sel_one_hot_i[47];
  assign data_masked[6028] = data_i[6028] & sel_one_hot_i[47];
  assign data_masked[6027] = data_i[6027] & sel_one_hot_i[47];
  assign data_masked[6026] = data_i[6026] & sel_one_hot_i[47];
  assign data_masked[6025] = data_i[6025] & sel_one_hot_i[47];
  assign data_masked[6024] = data_i[6024] & sel_one_hot_i[47];
  assign data_masked[6023] = data_i[6023] & sel_one_hot_i[47];
  assign data_masked[6022] = data_i[6022] & sel_one_hot_i[47];
  assign data_masked[6021] = data_i[6021] & sel_one_hot_i[47];
  assign data_masked[6020] = data_i[6020] & sel_one_hot_i[47];
  assign data_masked[6019] = data_i[6019] & sel_one_hot_i[47];
  assign data_masked[6018] = data_i[6018] & sel_one_hot_i[47];
  assign data_masked[6017] = data_i[6017] & sel_one_hot_i[47];
  assign data_masked[6016] = data_i[6016] & sel_one_hot_i[47];
  assign data_masked[6271] = data_i[6271] & sel_one_hot_i[48];
  assign data_masked[6270] = data_i[6270] & sel_one_hot_i[48];
  assign data_masked[6269] = data_i[6269] & sel_one_hot_i[48];
  assign data_masked[6268] = data_i[6268] & sel_one_hot_i[48];
  assign data_masked[6267] = data_i[6267] & sel_one_hot_i[48];
  assign data_masked[6266] = data_i[6266] & sel_one_hot_i[48];
  assign data_masked[6265] = data_i[6265] & sel_one_hot_i[48];
  assign data_masked[6264] = data_i[6264] & sel_one_hot_i[48];
  assign data_masked[6263] = data_i[6263] & sel_one_hot_i[48];
  assign data_masked[6262] = data_i[6262] & sel_one_hot_i[48];
  assign data_masked[6261] = data_i[6261] & sel_one_hot_i[48];
  assign data_masked[6260] = data_i[6260] & sel_one_hot_i[48];
  assign data_masked[6259] = data_i[6259] & sel_one_hot_i[48];
  assign data_masked[6258] = data_i[6258] & sel_one_hot_i[48];
  assign data_masked[6257] = data_i[6257] & sel_one_hot_i[48];
  assign data_masked[6256] = data_i[6256] & sel_one_hot_i[48];
  assign data_masked[6255] = data_i[6255] & sel_one_hot_i[48];
  assign data_masked[6254] = data_i[6254] & sel_one_hot_i[48];
  assign data_masked[6253] = data_i[6253] & sel_one_hot_i[48];
  assign data_masked[6252] = data_i[6252] & sel_one_hot_i[48];
  assign data_masked[6251] = data_i[6251] & sel_one_hot_i[48];
  assign data_masked[6250] = data_i[6250] & sel_one_hot_i[48];
  assign data_masked[6249] = data_i[6249] & sel_one_hot_i[48];
  assign data_masked[6248] = data_i[6248] & sel_one_hot_i[48];
  assign data_masked[6247] = data_i[6247] & sel_one_hot_i[48];
  assign data_masked[6246] = data_i[6246] & sel_one_hot_i[48];
  assign data_masked[6245] = data_i[6245] & sel_one_hot_i[48];
  assign data_masked[6244] = data_i[6244] & sel_one_hot_i[48];
  assign data_masked[6243] = data_i[6243] & sel_one_hot_i[48];
  assign data_masked[6242] = data_i[6242] & sel_one_hot_i[48];
  assign data_masked[6241] = data_i[6241] & sel_one_hot_i[48];
  assign data_masked[6240] = data_i[6240] & sel_one_hot_i[48];
  assign data_masked[6239] = data_i[6239] & sel_one_hot_i[48];
  assign data_masked[6238] = data_i[6238] & sel_one_hot_i[48];
  assign data_masked[6237] = data_i[6237] & sel_one_hot_i[48];
  assign data_masked[6236] = data_i[6236] & sel_one_hot_i[48];
  assign data_masked[6235] = data_i[6235] & sel_one_hot_i[48];
  assign data_masked[6234] = data_i[6234] & sel_one_hot_i[48];
  assign data_masked[6233] = data_i[6233] & sel_one_hot_i[48];
  assign data_masked[6232] = data_i[6232] & sel_one_hot_i[48];
  assign data_masked[6231] = data_i[6231] & sel_one_hot_i[48];
  assign data_masked[6230] = data_i[6230] & sel_one_hot_i[48];
  assign data_masked[6229] = data_i[6229] & sel_one_hot_i[48];
  assign data_masked[6228] = data_i[6228] & sel_one_hot_i[48];
  assign data_masked[6227] = data_i[6227] & sel_one_hot_i[48];
  assign data_masked[6226] = data_i[6226] & sel_one_hot_i[48];
  assign data_masked[6225] = data_i[6225] & sel_one_hot_i[48];
  assign data_masked[6224] = data_i[6224] & sel_one_hot_i[48];
  assign data_masked[6223] = data_i[6223] & sel_one_hot_i[48];
  assign data_masked[6222] = data_i[6222] & sel_one_hot_i[48];
  assign data_masked[6221] = data_i[6221] & sel_one_hot_i[48];
  assign data_masked[6220] = data_i[6220] & sel_one_hot_i[48];
  assign data_masked[6219] = data_i[6219] & sel_one_hot_i[48];
  assign data_masked[6218] = data_i[6218] & sel_one_hot_i[48];
  assign data_masked[6217] = data_i[6217] & sel_one_hot_i[48];
  assign data_masked[6216] = data_i[6216] & sel_one_hot_i[48];
  assign data_masked[6215] = data_i[6215] & sel_one_hot_i[48];
  assign data_masked[6214] = data_i[6214] & sel_one_hot_i[48];
  assign data_masked[6213] = data_i[6213] & sel_one_hot_i[48];
  assign data_masked[6212] = data_i[6212] & sel_one_hot_i[48];
  assign data_masked[6211] = data_i[6211] & sel_one_hot_i[48];
  assign data_masked[6210] = data_i[6210] & sel_one_hot_i[48];
  assign data_masked[6209] = data_i[6209] & sel_one_hot_i[48];
  assign data_masked[6208] = data_i[6208] & sel_one_hot_i[48];
  assign data_masked[6207] = data_i[6207] & sel_one_hot_i[48];
  assign data_masked[6206] = data_i[6206] & sel_one_hot_i[48];
  assign data_masked[6205] = data_i[6205] & sel_one_hot_i[48];
  assign data_masked[6204] = data_i[6204] & sel_one_hot_i[48];
  assign data_masked[6203] = data_i[6203] & sel_one_hot_i[48];
  assign data_masked[6202] = data_i[6202] & sel_one_hot_i[48];
  assign data_masked[6201] = data_i[6201] & sel_one_hot_i[48];
  assign data_masked[6200] = data_i[6200] & sel_one_hot_i[48];
  assign data_masked[6199] = data_i[6199] & sel_one_hot_i[48];
  assign data_masked[6198] = data_i[6198] & sel_one_hot_i[48];
  assign data_masked[6197] = data_i[6197] & sel_one_hot_i[48];
  assign data_masked[6196] = data_i[6196] & sel_one_hot_i[48];
  assign data_masked[6195] = data_i[6195] & sel_one_hot_i[48];
  assign data_masked[6194] = data_i[6194] & sel_one_hot_i[48];
  assign data_masked[6193] = data_i[6193] & sel_one_hot_i[48];
  assign data_masked[6192] = data_i[6192] & sel_one_hot_i[48];
  assign data_masked[6191] = data_i[6191] & sel_one_hot_i[48];
  assign data_masked[6190] = data_i[6190] & sel_one_hot_i[48];
  assign data_masked[6189] = data_i[6189] & sel_one_hot_i[48];
  assign data_masked[6188] = data_i[6188] & sel_one_hot_i[48];
  assign data_masked[6187] = data_i[6187] & sel_one_hot_i[48];
  assign data_masked[6186] = data_i[6186] & sel_one_hot_i[48];
  assign data_masked[6185] = data_i[6185] & sel_one_hot_i[48];
  assign data_masked[6184] = data_i[6184] & sel_one_hot_i[48];
  assign data_masked[6183] = data_i[6183] & sel_one_hot_i[48];
  assign data_masked[6182] = data_i[6182] & sel_one_hot_i[48];
  assign data_masked[6181] = data_i[6181] & sel_one_hot_i[48];
  assign data_masked[6180] = data_i[6180] & sel_one_hot_i[48];
  assign data_masked[6179] = data_i[6179] & sel_one_hot_i[48];
  assign data_masked[6178] = data_i[6178] & sel_one_hot_i[48];
  assign data_masked[6177] = data_i[6177] & sel_one_hot_i[48];
  assign data_masked[6176] = data_i[6176] & sel_one_hot_i[48];
  assign data_masked[6175] = data_i[6175] & sel_one_hot_i[48];
  assign data_masked[6174] = data_i[6174] & sel_one_hot_i[48];
  assign data_masked[6173] = data_i[6173] & sel_one_hot_i[48];
  assign data_masked[6172] = data_i[6172] & sel_one_hot_i[48];
  assign data_masked[6171] = data_i[6171] & sel_one_hot_i[48];
  assign data_masked[6170] = data_i[6170] & sel_one_hot_i[48];
  assign data_masked[6169] = data_i[6169] & sel_one_hot_i[48];
  assign data_masked[6168] = data_i[6168] & sel_one_hot_i[48];
  assign data_masked[6167] = data_i[6167] & sel_one_hot_i[48];
  assign data_masked[6166] = data_i[6166] & sel_one_hot_i[48];
  assign data_masked[6165] = data_i[6165] & sel_one_hot_i[48];
  assign data_masked[6164] = data_i[6164] & sel_one_hot_i[48];
  assign data_masked[6163] = data_i[6163] & sel_one_hot_i[48];
  assign data_masked[6162] = data_i[6162] & sel_one_hot_i[48];
  assign data_masked[6161] = data_i[6161] & sel_one_hot_i[48];
  assign data_masked[6160] = data_i[6160] & sel_one_hot_i[48];
  assign data_masked[6159] = data_i[6159] & sel_one_hot_i[48];
  assign data_masked[6158] = data_i[6158] & sel_one_hot_i[48];
  assign data_masked[6157] = data_i[6157] & sel_one_hot_i[48];
  assign data_masked[6156] = data_i[6156] & sel_one_hot_i[48];
  assign data_masked[6155] = data_i[6155] & sel_one_hot_i[48];
  assign data_masked[6154] = data_i[6154] & sel_one_hot_i[48];
  assign data_masked[6153] = data_i[6153] & sel_one_hot_i[48];
  assign data_masked[6152] = data_i[6152] & sel_one_hot_i[48];
  assign data_masked[6151] = data_i[6151] & sel_one_hot_i[48];
  assign data_masked[6150] = data_i[6150] & sel_one_hot_i[48];
  assign data_masked[6149] = data_i[6149] & sel_one_hot_i[48];
  assign data_masked[6148] = data_i[6148] & sel_one_hot_i[48];
  assign data_masked[6147] = data_i[6147] & sel_one_hot_i[48];
  assign data_masked[6146] = data_i[6146] & sel_one_hot_i[48];
  assign data_masked[6145] = data_i[6145] & sel_one_hot_i[48];
  assign data_masked[6144] = data_i[6144] & sel_one_hot_i[48];
  assign data_masked[6399] = data_i[6399] & sel_one_hot_i[49];
  assign data_masked[6398] = data_i[6398] & sel_one_hot_i[49];
  assign data_masked[6397] = data_i[6397] & sel_one_hot_i[49];
  assign data_masked[6396] = data_i[6396] & sel_one_hot_i[49];
  assign data_masked[6395] = data_i[6395] & sel_one_hot_i[49];
  assign data_masked[6394] = data_i[6394] & sel_one_hot_i[49];
  assign data_masked[6393] = data_i[6393] & sel_one_hot_i[49];
  assign data_masked[6392] = data_i[6392] & sel_one_hot_i[49];
  assign data_masked[6391] = data_i[6391] & sel_one_hot_i[49];
  assign data_masked[6390] = data_i[6390] & sel_one_hot_i[49];
  assign data_masked[6389] = data_i[6389] & sel_one_hot_i[49];
  assign data_masked[6388] = data_i[6388] & sel_one_hot_i[49];
  assign data_masked[6387] = data_i[6387] & sel_one_hot_i[49];
  assign data_masked[6386] = data_i[6386] & sel_one_hot_i[49];
  assign data_masked[6385] = data_i[6385] & sel_one_hot_i[49];
  assign data_masked[6384] = data_i[6384] & sel_one_hot_i[49];
  assign data_masked[6383] = data_i[6383] & sel_one_hot_i[49];
  assign data_masked[6382] = data_i[6382] & sel_one_hot_i[49];
  assign data_masked[6381] = data_i[6381] & sel_one_hot_i[49];
  assign data_masked[6380] = data_i[6380] & sel_one_hot_i[49];
  assign data_masked[6379] = data_i[6379] & sel_one_hot_i[49];
  assign data_masked[6378] = data_i[6378] & sel_one_hot_i[49];
  assign data_masked[6377] = data_i[6377] & sel_one_hot_i[49];
  assign data_masked[6376] = data_i[6376] & sel_one_hot_i[49];
  assign data_masked[6375] = data_i[6375] & sel_one_hot_i[49];
  assign data_masked[6374] = data_i[6374] & sel_one_hot_i[49];
  assign data_masked[6373] = data_i[6373] & sel_one_hot_i[49];
  assign data_masked[6372] = data_i[6372] & sel_one_hot_i[49];
  assign data_masked[6371] = data_i[6371] & sel_one_hot_i[49];
  assign data_masked[6370] = data_i[6370] & sel_one_hot_i[49];
  assign data_masked[6369] = data_i[6369] & sel_one_hot_i[49];
  assign data_masked[6368] = data_i[6368] & sel_one_hot_i[49];
  assign data_masked[6367] = data_i[6367] & sel_one_hot_i[49];
  assign data_masked[6366] = data_i[6366] & sel_one_hot_i[49];
  assign data_masked[6365] = data_i[6365] & sel_one_hot_i[49];
  assign data_masked[6364] = data_i[6364] & sel_one_hot_i[49];
  assign data_masked[6363] = data_i[6363] & sel_one_hot_i[49];
  assign data_masked[6362] = data_i[6362] & sel_one_hot_i[49];
  assign data_masked[6361] = data_i[6361] & sel_one_hot_i[49];
  assign data_masked[6360] = data_i[6360] & sel_one_hot_i[49];
  assign data_masked[6359] = data_i[6359] & sel_one_hot_i[49];
  assign data_masked[6358] = data_i[6358] & sel_one_hot_i[49];
  assign data_masked[6357] = data_i[6357] & sel_one_hot_i[49];
  assign data_masked[6356] = data_i[6356] & sel_one_hot_i[49];
  assign data_masked[6355] = data_i[6355] & sel_one_hot_i[49];
  assign data_masked[6354] = data_i[6354] & sel_one_hot_i[49];
  assign data_masked[6353] = data_i[6353] & sel_one_hot_i[49];
  assign data_masked[6352] = data_i[6352] & sel_one_hot_i[49];
  assign data_masked[6351] = data_i[6351] & sel_one_hot_i[49];
  assign data_masked[6350] = data_i[6350] & sel_one_hot_i[49];
  assign data_masked[6349] = data_i[6349] & sel_one_hot_i[49];
  assign data_masked[6348] = data_i[6348] & sel_one_hot_i[49];
  assign data_masked[6347] = data_i[6347] & sel_one_hot_i[49];
  assign data_masked[6346] = data_i[6346] & sel_one_hot_i[49];
  assign data_masked[6345] = data_i[6345] & sel_one_hot_i[49];
  assign data_masked[6344] = data_i[6344] & sel_one_hot_i[49];
  assign data_masked[6343] = data_i[6343] & sel_one_hot_i[49];
  assign data_masked[6342] = data_i[6342] & sel_one_hot_i[49];
  assign data_masked[6341] = data_i[6341] & sel_one_hot_i[49];
  assign data_masked[6340] = data_i[6340] & sel_one_hot_i[49];
  assign data_masked[6339] = data_i[6339] & sel_one_hot_i[49];
  assign data_masked[6338] = data_i[6338] & sel_one_hot_i[49];
  assign data_masked[6337] = data_i[6337] & sel_one_hot_i[49];
  assign data_masked[6336] = data_i[6336] & sel_one_hot_i[49];
  assign data_masked[6335] = data_i[6335] & sel_one_hot_i[49];
  assign data_masked[6334] = data_i[6334] & sel_one_hot_i[49];
  assign data_masked[6333] = data_i[6333] & sel_one_hot_i[49];
  assign data_masked[6332] = data_i[6332] & sel_one_hot_i[49];
  assign data_masked[6331] = data_i[6331] & sel_one_hot_i[49];
  assign data_masked[6330] = data_i[6330] & sel_one_hot_i[49];
  assign data_masked[6329] = data_i[6329] & sel_one_hot_i[49];
  assign data_masked[6328] = data_i[6328] & sel_one_hot_i[49];
  assign data_masked[6327] = data_i[6327] & sel_one_hot_i[49];
  assign data_masked[6326] = data_i[6326] & sel_one_hot_i[49];
  assign data_masked[6325] = data_i[6325] & sel_one_hot_i[49];
  assign data_masked[6324] = data_i[6324] & sel_one_hot_i[49];
  assign data_masked[6323] = data_i[6323] & sel_one_hot_i[49];
  assign data_masked[6322] = data_i[6322] & sel_one_hot_i[49];
  assign data_masked[6321] = data_i[6321] & sel_one_hot_i[49];
  assign data_masked[6320] = data_i[6320] & sel_one_hot_i[49];
  assign data_masked[6319] = data_i[6319] & sel_one_hot_i[49];
  assign data_masked[6318] = data_i[6318] & sel_one_hot_i[49];
  assign data_masked[6317] = data_i[6317] & sel_one_hot_i[49];
  assign data_masked[6316] = data_i[6316] & sel_one_hot_i[49];
  assign data_masked[6315] = data_i[6315] & sel_one_hot_i[49];
  assign data_masked[6314] = data_i[6314] & sel_one_hot_i[49];
  assign data_masked[6313] = data_i[6313] & sel_one_hot_i[49];
  assign data_masked[6312] = data_i[6312] & sel_one_hot_i[49];
  assign data_masked[6311] = data_i[6311] & sel_one_hot_i[49];
  assign data_masked[6310] = data_i[6310] & sel_one_hot_i[49];
  assign data_masked[6309] = data_i[6309] & sel_one_hot_i[49];
  assign data_masked[6308] = data_i[6308] & sel_one_hot_i[49];
  assign data_masked[6307] = data_i[6307] & sel_one_hot_i[49];
  assign data_masked[6306] = data_i[6306] & sel_one_hot_i[49];
  assign data_masked[6305] = data_i[6305] & sel_one_hot_i[49];
  assign data_masked[6304] = data_i[6304] & sel_one_hot_i[49];
  assign data_masked[6303] = data_i[6303] & sel_one_hot_i[49];
  assign data_masked[6302] = data_i[6302] & sel_one_hot_i[49];
  assign data_masked[6301] = data_i[6301] & sel_one_hot_i[49];
  assign data_masked[6300] = data_i[6300] & sel_one_hot_i[49];
  assign data_masked[6299] = data_i[6299] & sel_one_hot_i[49];
  assign data_masked[6298] = data_i[6298] & sel_one_hot_i[49];
  assign data_masked[6297] = data_i[6297] & sel_one_hot_i[49];
  assign data_masked[6296] = data_i[6296] & sel_one_hot_i[49];
  assign data_masked[6295] = data_i[6295] & sel_one_hot_i[49];
  assign data_masked[6294] = data_i[6294] & sel_one_hot_i[49];
  assign data_masked[6293] = data_i[6293] & sel_one_hot_i[49];
  assign data_masked[6292] = data_i[6292] & sel_one_hot_i[49];
  assign data_masked[6291] = data_i[6291] & sel_one_hot_i[49];
  assign data_masked[6290] = data_i[6290] & sel_one_hot_i[49];
  assign data_masked[6289] = data_i[6289] & sel_one_hot_i[49];
  assign data_masked[6288] = data_i[6288] & sel_one_hot_i[49];
  assign data_masked[6287] = data_i[6287] & sel_one_hot_i[49];
  assign data_masked[6286] = data_i[6286] & sel_one_hot_i[49];
  assign data_masked[6285] = data_i[6285] & sel_one_hot_i[49];
  assign data_masked[6284] = data_i[6284] & sel_one_hot_i[49];
  assign data_masked[6283] = data_i[6283] & sel_one_hot_i[49];
  assign data_masked[6282] = data_i[6282] & sel_one_hot_i[49];
  assign data_masked[6281] = data_i[6281] & sel_one_hot_i[49];
  assign data_masked[6280] = data_i[6280] & sel_one_hot_i[49];
  assign data_masked[6279] = data_i[6279] & sel_one_hot_i[49];
  assign data_masked[6278] = data_i[6278] & sel_one_hot_i[49];
  assign data_masked[6277] = data_i[6277] & sel_one_hot_i[49];
  assign data_masked[6276] = data_i[6276] & sel_one_hot_i[49];
  assign data_masked[6275] = data_i[6275] & sel_one_hot_i[49];
  assign data_masked[6274] = data_i[6274] & sel_one_hot_i[49];
  assign data_masked[6273] = data_i[6273] & sel_one_hot_i[49];
  assign data_masked[6272] = data_i[6272] & sel_one_hot_i[49];
  assign data_masked[6527] = data_i[6527] & sel_one_hot_i[50];
  assign data_masked[6526] = data_i[6526] & sel_one_hot_i[50];
  assign data_masked[6525] = data_i[6525] & sel_one_hot_i[50];
  assign data_masked[6524] = data_i[6524] & sel_one_hot_i[50];
  assign data_masked[6523] = data_i[6523] & sel_one_hot_i[50];
  assign data_masked[6522] = data_i[6522] & sel_one_hot_i[50];
  assign data_masked[6521] = data_i[6521] & sel_one_hot_i[50];
  assign data_masked[6520] = data_i[6520] & sel_one_hot_i[50];
  assign data_masked[6519] = data_i[6519] & sel_one_hot_i[50];
  assign data_masked[6518] = data_i[6518] & sel_one_hot_i[50];
  assign data_masked[6517] = data_i[6517] & sel_one_hot_i[50];
  assign data_masked[6516] = data_i[6516] & sel_one_hot_i[50];
  assign data_masked[6515] = data_i[6515] & sel_one_hot_i[50];
  assign data_masked[6514] = data_i[6514] & sel_one_hot_i[50];
  assign data_masked[6513] = data_i[6513] & sel_one_hot_i[50];
  assign data_masked[6512] = data_i[6512] & sel_one_hot_i[50];
  assign data_masked[6511] = data_i[6511] & sel_one_hot_i[50];
  assign data_masked[6510] = data_i[6510] & sel_one_hot_i[50];
  assign data_masked[6509] = data_i[6509] & sel_one_hot_i[50];
  assign data_masked[6508] = data_i[6508] & sel_one_hot_i[50];
  assign data_masked[6507] = data_i[6507] & sel_one_hot_i[50];
  assign data_masked[6506] = data_i[6506] & sel_one_hot_i[50];
  assign data_masked[6505] = data_i[6505] & sel_one_hot_i[50];
  assign data_masked[6504] = data_i[6504] & sel_one_hot_i[50];
  assign data_masked[6503] = data_i[6503] & sel_one_hot_i[50];
  assign data_masked[6502] = data_i[6502] & sel_one_hot_i[50];
  assign data_masked[6501] = data_i[6501] & sel_one_hot_i[50];
  assign data_masked[6500] = data_i[6500] & sel_one_hot_i[50];
  assign data_masked[6499] = data_i[6499] & sel_one_hot_i[50];
  assign data_masked[6498] = data_i[6498] & sel_one_hot_i[50];
  assign data_masked[6497] = data_i[6497] & sel_one_hot_i[50];
  assign data_masked[6496] = data_i[6496] & sel_one_hot_i[50];
  assign data_masked[6495] = data_i[6495] & sel_one_hot_i[50];
  assign data_masked[6494] = data_i[6494] & sel_one_hot_i[50];
  assign data_masked[6493] = data_i[6493] & sel_one_hot_i[50];
  assign data_masked[6492] = data_i[6492] & sel_one_hot_i[50];
  assign data_masked[6491] = data_i[6491] & sel_one_hot_i[50];
  assign data_masked[6490] = data_i[6490] & sel_one_hot_i[50];
  assign data_masked[6489] = data_i[6489] & sel_one_hot_i[50];
  assign data_masked[6488] = data_i[6488] & sel_one_hot_i[50];
  assign data_masked[6487] = data_i[6487] & sel_one_hot_i[50];
  assign data_masked[6486] = data_i[6486] & sel_one_hot_i[50];
  assign data_masked[6485] = data_i[6485] & sel_one_hot_i[50];
  assign data_masked[6484] = data_i[6484] & sel_one_hot_i[50];
  assign data_masked[6483] = data_i[6483] & sel_one_hot_i[50];
  assign data_masked[6482] = data_i[6482] & sel_one_hot_i[50];
  assign data_masked[6481] = data_i[6481] & sel_one_hot_i[50];
  assign data_masked[6480] = data_i[6480] & sel_one_hot_i[50];
  assign data_masked[6479] = data_i[6479] & sel_one_hot_i[50];
  assign data_masked[6478] = data_i[6478] & sel_one_hot_i[50];
  assign data_masked[6477] = data_i[6477] & sel_one_hot_i[50];
  assign data_masked[6476] = data_i[6476] & sel_one_hot_i[50];
  assign data_masked[6475] = data_i[6475] & sel_one_hot_i[50];
  assign data_masked[6474] = data_i[6474] & sel_one_hot_i[50];
  assign data_masked[6473] = data_i[6473] & sel_one_hot_i[50];
  assign data_masked[6472] = data_i[6472] & sel_one_hot_i[50];
  assign data_masked[6471] = data_i[6471] & sel_one_hot_i[50];
  assign data_masked[6470] = data_i[6470] & sel_one_hot_i[50];
  assign data_masked[6469] = data_i[6469] & sel_one_hot_i[50];
  assign data_masked[6468] = data_i[6468] & sel_one_hot_i[50];
  assign data_masked[6467] = data_i[6467] & sel_one_hot_i[50];
  assign data_masked[6466] = data_i[6466] & sel_one_hot_i[50];
  assign data_masked[6465] = data_i[6465] & sel_one_hot_i[50];
  assign data_masked[6464] = data_i[6464] & sel_one_hot_i[50];
  assign data_masked[6463] = data_i[6463] & sel_one_hot_i[50];
  assign data_masked[6462] = data_i[6462] & sel_one_hot_i[50];
  assign data_masked[6461] = data_i[6461] & sel_one_hot_i[50];
  assign data_masked[6460] = data_i[6460] & sel_one_hot_i[50];
  assign data_masked[6459] = data_i[6459] & sel_one_hot_i[50];
  assign data_masked[6458] = data_i[6458] & sel_one_hot_i[50];
  assign data_masked[6457] = data_i[6457] & sel_one_hot_i[50];
  assign data_masked[6456] = data_i[6456] & sel_one_hot_i[50];
  assign data_masked[6455] = data_i[6455] & sel_one_hot_i[50];
  assign data_masked[6454] = data_i[6454] & sel_one_hot_i[50];
  assign data_masked[6453] = data_i[6453] & sel_one_hot_i[50];
  assign data_masked[6452] = data_i[6452] & sel_one_hot_i[50];
  assign data_masked[6451] = data_i[6451] & sel_one_hot_i[50];
  assign data_masked[6450] = data_i[6450] & sel_one_hot_i[50];
  assign data_masked[6449] = data_i[6449] & sel_one_hot_i[50];
  assign data_masked[6448] = data_i[6448] & sel_one_hot_i[50];
  assign data_masked[6447] = data_i[6447] & sel_one_hot_i[50];
  assign data_masked[6446] = data_i[6446] & sel_one_hot_i[50];
  assign data_masked[6445] = data_i[6445] & sel_one_hot_i[50];
  assign data_masked[6444] = data_i[6444] & sel_one_hot_i[50];
  assign data_masked[6443] = data_i[6443] & sel_one_hot_i[50];
  assign data_masked[6442] = data_i[6442] & sel_one_hot_i[50];
  assign data_masked[6441] = data_i[6441] & sel_one_hot_i[50];
  assign data_masked[6440] = data_i[6440] & sel_one_hot_i[50];
  assign data_masked[6439] = data_i[6439] & sel_one_hot_i[50];
  assign data_masked[6438] = data_i[6438] & sel_one_hot_i[50];
  assign data_masked[6437] = data_i[6437] & sel_one_hot_i[50];
  assign data_masked[6436] = data_i[6436] & sel_one_hot_i[50];
  assign data_masked[6435] = data_i[6435] & sel_one_hot_i[50];
  assign data_masked[6434] = data_i[6434] & sel_one_hot_i[50];
  assign data_masked[6433] = data_i[6433] & sel_one_hot_i[50];
  assign data_masked[6432] = data_i[6432] & sel_one_hot_i[50];
  assign data_masked[6431] = data_i[6431] & sel_one_hot_i[50];
  assign data_masked[6430] = data_i[6430] & sel_one_hot_i[50];
  assign data_masked[6429] = data_i[6429] & sel_one_hot_i[50];
  assign data_masked[6428] = data_i[6428] & sel_one_hot_i[50];
  assign data_masked[6427] = data_i[6427] & sel_one_hot_i[50];
  assign data_masked[6426] = data_i[6426] & sel_one_hot_i[50];
  assign data_masked[6425] = data_i[6425] & sel_one_hot_i[50];
  assign data_masked[6424] = data_i[6424] & sel_one_hot_i[50];
  assign data_masked[6423] = data_i[6423] & sel_one_hot_i[50];
  assign data_masked[6422] = data_i[6422] & sel_one_hot_i[50];
  assign data_masked[6421] = data_i[6421] & sel_one_hot_i[50];
  assign data_masked[6420] = data_i[6420] & sel_one_hot_i[50];
  assign data_masked[6419] = data_i[6419] & sel_one_hot_i[50];
  assign data_masked[6418] = data_i[6418] & sel_one_hot_i[50];
  assign data_masked[6417] = data_i[6417] & sel_one_hot_i[50];
  assign data_masked[6416] = data_i[6416] & sel_one_hot_i[50];
  assign data_masked[6415] = data_i[6415] & sel_one_hot_i[50];
  assign data_masked[6414] = data_i[6414] & sel_one_hot_i[50];
  assign data_masked[6413] = data_i[6413] & sel_one_hot_i[50];
  assign data_masked[6412] = data_i[6412] & sel_one_hot_i[50];
  assign data_masked[6411] = data_i[6411] & sel_one_hot_i[50];
  assign data_masked[6410] = data_i[6410] & sel_one_hot_i[50];
  assign data_masked[6409] = data_i[6409] & sel_one_hot_i[50];
  assign data_masked[6408] = data_i[6408] & sel_one_hot_i[50];
  assign data_masked[6407] = data_i[6407] & sel_one_hot_i[50];
  assign data_masked[6406] = data_i[6406] & sel_one_hot_i[50];
  assign data_masked[6405] = data_i[6405] & sel_one_hot_i[50];
  assign data_masked[6404] = data_i[6404] & sel_one_hot_i[50];
  assign data_masked[6403] = data_i[6403] & sel_one_hot_i[50];
  assign data_masked[6402] = data_i[6402] & sel_one_hot_i[50];
  assign data_masked[6401] = data_i[6401] & sel_one_hot_i[50];
  assign data_masked[6400] = data_i[6400] & sel_one_hot_i[50];
  assign data_masked[6655] = data_i[6655] & sel_one_hot_i[51];
  assign data_masked[6654] = data_i[6654] & sel_one_hot_i[51];
  assign data_masked[6653] = data_i[6653] & sel_one_hot_i[51];
  assign data_masked[6652] = data_i[6652] & sel_one_hot_i[51];
  assign data_masked[6651] = data_i[6651] & sel_one_hot_i[51];
  assign data_masked[6650] = data_i[6650] & sel_one_hot_i[51];
  assign data_masked[6649] = data_i[6649] & sel_one_hot_i[51];
  assign data_masked[6648] = data_i[6648] & sel_one_hot_i[51];
  assign data_masked[6647] = data_i[6647] & sel_one_hot_i[51];
  assign data_masked[6646] = data_i[6646] & sel_one_hot_i[51];
  assign data_masked[6645] = data_i[6645] & sel_one_hot_i[51];
  assign data_masked[6644] = data_i[6644] & sel_one_hot_i[51];
  assign data_masked[6643] = data_i[6643] & sel_one_hot_i[51];
  assign data_masked[6642] = data_i[6642] & sel_one_hot_i[51];
  assign data_masked[6641] = data_i[6641] & sel_one_hot_i[51];
  assign data_masked[6640] = data_i[6640] & sel_one_hot_i[51];
  assign data_masked[6639] = data_i[6639] & sel_one_hot_i[51];
  assign data_masked[6638] = data_i[6638] & sel_one_hot_i[51];
  assign data_masked[6637] = data_i[6637] & sel_one_hot_i[51];
  assign data_masked[6636] = data_i[6636] & sel_one_hot_i[51];
  assign data_masked[6635] = data_i[6635] & sel_one_hot_i[51];
  assign data_masked[6634] = data_i[6634] & sel_one_hot_i[51];
  assign data_masked[6633] = data_i[6633] & sel_one_hot_i[51];
  assign data_masked[6632] = data_i[6632] & sel_one_hot_i[51];
  assign data_masked[6631] = data_i[6631] & sel_one_hot_i[51];
  assign data_masked[6630] = data_i[6630] & sel_one_hot_i[51];
  assign data_masked[6629] = data_i[6629] & sel_one_hot_i[51];
  assign data_masked[6628] = data_i[6628] & sel_one_hot_i[51];
  assign data_masked[6627] = data_i[6627] & sel_one_hot_i[51];
  assign data_masked[6626] = data_i[6626] & sel_one_hot_i[51];
  assign data_masked[6625] = data_i[6625] & sel_one_hot_i[51];
  assign data_masked[6624] = data_i[6624] & sel_one_hot_i[51];
  assign data_masked[6623] = data_i[6623] & sel_one_hot_i[51];
  assign data_masked[6622] = data_i[6622] & sel_one_hot_i[51];
  assign data_masked[6621] = data_i[6621] & sel_one_hot_i[51];
  assign data_masked[6620] = data_i[6620] & sel_one_hot_i[51];
  assign data_masked[6619] = data_i[6619] & sel_one_hot_i[51];
  assign data_masked[6618] = data_i[6618] & sel_one_hot_i[51];
  assign data_masked[6617] = data_i[6617] & sel_one_hot_i[51];
  assign data_masked[6616] = data_i[6616] & sel_one_hot_i[51];
  assign data_masked[6615] = data_i[6615] & sel_one_hot_i[51];
  assign data_masked[6614] = data_i[6614] & sel_one_hot_i[51];
  assign data_masked[6613] = data_i[6613] & sel_one_hot_i[51];
  assign data_masked[6612] = data_i[6612] & sel_one_hot_i[51];
  assign data_masked[6611] = data_i[6611] & sel_one_hot_i[51];
  assign data_masked[6610] = data_i[6610] & sel_one_hot_i[51];
  assign data_masked[6609] = data_i[6609] & sel_one_hot_i[51];
  assign data_masked[6608] = data_i[6608] & sel_one_hot_i[51];
  assign data_masked[6607] = data_i[6607] & sel_one_hot_i[51];
  assign data_masked[6606] = data_i[6606] & sel_one_hot_i[51];
  assign data_masked[6605] = data_i[6605] & sel_one_hot_i[51];
  assign data_masked[6604] = data_i[6604] & sel_one_hot_i[51];
  assign data_masked[6603] = data_i[6603] & sel_one_hot_i[51];
  assign data_masked[6602] = data_i[6602] & sel_one_hot_i[51];
  assign data_masked[6601] = data_i[6601] & sel_one_hot_i[51];
  assign data_masked[6600] = data_i[6600] & sel_one_hot_i[51];
  assign data_masked[6599] = data_i[6599] & sel_one_hot_i[51];
  assign data_masked[6598] = data_i[6598] & sel_one_hot_i[51];
  assign data_masked[6597] = data_i[6597] & sel_one_hot_i[51];
  assign data_masked[6596] = data_i[6596] & sel_one_hot_i[51];
  assign data_masked[6595] = data_i[6595] & sel_one_hot_i[51];
  assign data_masked[6594] = data_i[6594] & sel_one_hot_i[51];
  assign data_masked[6593] = data_i[6593] & sel_one_hot_i[51];
  assign data_masked[6592] = data_i[6592] & sel_one_hot_i[51];
  assign data_masked[6591] = data_i[6591] & sel_one_hot_i[51];
  assign data_masked[6590] = data_i[6590] & sel_one_hot_i[51];
  assign data_masked[6589] = data_i[6589] & sel_one_hot_i[51];
  assign data_masked[6588] = data_i[6588] & sel_one_hot_i[51];
  assign data_masked[6587] = data_i[6587] & sel_one_hot_i[51];
  assign data_masked[6586] = data_i[6586] & sel_one_hot_i[51];
  assign data_masked[6585] = data_i[6585] & sel_one_hot_i[51];
  assign data_masked[6584] = data_i[6584] & sel_one_hot_i[51];
  assign data_masked[6583] = data_i[6583] & sel_one_hot_i[51];
  assign data_masked[6582] = data_i[6582] & sel_one_hot_i[51];
  assign data_masked[6581] = data_i[6581] & sel_one_hot_i[51];
  assign data_masked[6580] = data_i[6580] & sel_one_hot_i[51];
  assign data_masked[6579] = data_i[6579] & sel_one_hot_i[51];
  assign data_masked[6578] = data_i[6578] & sel_one_hot_i[51];
  assign data_masked[6577] = data_i[6577] & sel_one_hot_i[51];
  assign data_masked[6576] = data_i[6576] & sel_one_hot_i[51];
  assign data_masked[6575] = data_i[6575] & sel_one_hot_i[51];
  assign data_masked[6574] = data_i[6574] & sel_one_hot_i[51];
  assign data_masked[6573] = data_i[6573] & sel_one_hot_i[51];
  assign data_masked[6572] = data_i[6572] & sel_one_hot_i[51];
  assign data_masked[6571] = data_i[6571] & sel_one_hot_i[51];
  assign data_masked[6570] = data_i[6570] & sel_one_hot_i[51];
  assign data_masked[6569] = data_i[6569] & sel_one_hot_i[51];
  assign data_masked[6568] = data_i[6568] & sel_one_hot_i[51];
  assign data_masked[6567] = data_i[6567] & sel_one_hot_i[51];
  assign data_masked[6566] = data_i[6566] & sel_one_hot_i[51];
  assign data_masked[6565] = data_i[6565] & sel_one_hot_i[51];
  assign data_masked[6564] = data_i[6564] & sel_one_hot_i[51];
  assign data_masked[6563] = data_i[6563] & sel_one_hot_i[51];
  assign data_masked[6562] = data_i[6562] & sel_one_hot_i[51];
  assign data_masked[6561] = data_i[6561] & sel_one_hot_i[51];
  assign data_masked[6560] = data_i[6560] & sel_one_hot_i[51];
  assign data_masked[6559] = data_i[6559] & sel_one_hot_i[51];
  assign data_masked[6558] = data_i[6558] & sel_one_hot_i[51];
  assign data_masked[6557] = data_i[6557] & sel_one_hot_i[51];
  assign data_masked[6556] = data_i[6556] & sel_one_hot_i[51];
  assign data_masked[6555] = data_i[6555] & sel_one_hot_i[51];
  assign data_masked[6554] = data_i[6554] & sel_one_hot_i[51];
  assign data_masked[6553] = data_i[6553] & sel_one_hot_i[51];
  assign data_masked[6552] = data_i[6552] & sel_one_hot_i[51];
  assign data_masked[6551] = data_i[6551] & sel_one_hot_i[51];
  assign data_masked[6550] = data_i[6550] & sel_one_hot_i[51];
  assign data_masked[6549] = data_i[6549] & sel_one_hot_i[51];
  assign data_masked[6548] = data_i[6548] & sel_one_hot_i[51];
  assign data_masked[6547] = data_i[6547] & sel_one_hot_i[51];
  assign data_masked[6546] = data_i[6546] & sel_one_hot_i[51];
  assign data_masked[6545] = data_i[6545] & sel_one_hot_i[51];
  assign data_masked[6544] = data_i[6544] & sel_one_hot_i[51];
  assign data_masked[6543] = data_i[6543] & sel_one_hot_i[51];
  assign data_masked[6542] = data_i[6542] & sel_one_hot_i[51];
  assign data_masked[6541] = data_i[6541] & sel_one_hot_i[51];
  assign data_masked[6540] = data_i[6540] & sel_one_hot_i[51];
  assign data_masked[6539] = data_i[6539] & sel_one_hot_i[51];
  assign data_masked[6538] = data_i[6538] & sel_one_hot_i[51];
  assign data_masked[6537] = data_i[6537] & sel_one_hot_i[51];
  assign data_masked[6536] = data_i[6536] & sel_one_hot_i[51];
  assign data_masked[6535] = data_i[6535] & sel_one_hot_i[51];
  assign data_masked[6534] = data_i[6534] & sel_one_hot_i[51];
  assign data_masked[6533] = data_i[6533] & sel_one_hot_i[51];
  assign data_masked[6532] = data_i[6532] & sel_one_hot_i[51];
  assign data_masked[6531] = data_i[6531] & sel_one_hot_i[51];
  assign data_masked[6530] = data_i[6530] & sel_one_hot_i[51];
  assign data_masked[6529] = data_i[6529] & sel_one_hot_i[51];
  assign data_masked[6528] = data_i[6528] & sel_one_hot_i[51];
  assign data_masked[6783] = data_i[6783] & sel_one_hot_i[52];
  assign data_masked[6782] = data_i[6782] & sel_one_hot_i[52];
  assign data_masked[6781] = data_i[6781] & sel_one_hot_i[52];
  assign data_masked[6780] = data_i[6780] & sel_one_hot_i[52];
  assign data_masked[6779] = data_i[6779] & sel_one_hot_i[52];
  assign data_masked[6778] = data_i[6778] & sel_one_hot_i[52];
  assign data_masked[6777] = data_i[6777] & sel_one_hot_i[52];
  assign data_masked[6776] = data_i[6776] & sel_one_hot_i[52];
  assign data_masked[6775] = data_i[6775] & sel_one_hot_i[52];
  assign data_masked[6774] = data_i[6774] & sel_one_hot_i[52];
  assign data_masked[6773] = data_i[6773] & sel_one_hot_i[52];
  assign data_masked[6772] = data_i[6772] & sel_one_hot_i[52];
  assign data_masked[6771] = data_i[6771] & sel_one_hot_i[52];
  assign data_masked[6770] = data_i[6770] & sel_one_hot_i[52];
  assign data_masked[6769] = data_i[6769] & sel_one_hot_i[52];
  assign data_masked[6768] = data_i[6768] & sel_one_hot_i[52];
  assign data_masked[6767] = data_i[6767] & sel_one_hot_i[52];
  assign data_masked[6766] = data_i[6766] & sel_one_hot_i[52];
  assign data_masked[6765] = data_i[6765] & sel_one_hot_i[52];
  assign data_masked[6764] = data_i[6764] & sel_one_hot_i[52];
  assign data_masked[6763] = data_i[6763] & sel_one_hot_i[52];
  assign data_masked[6762] = data_i[6762] & sel_one_hot_i[52];
  assign data_masked[6761] = data_i[6761] & sel_one_hot_i[52];
  assign data_masked[6760] = data_i[6760] & sel_one_hot_i[52];
  assign data_masked[6759] = data_i[6759] & sel_one_hot_i[52];
  assign data_masked[6758] = data_i[6758] & sel_one_hot_i[52];
  assign data_masked[6757] = data_i[6757] & sel_one_hot_i[52];
  assign data_masked[6756] = data_i[6756] & sel_one_hot_i[52];
  assign data_masked[6755] = data_i[6755] & sel_one_hot_i[52];
  assign data_masked[6754] = data_i[6754] & sel_one_hot_i[52];
  assign data_masked[6753] = data_i[6753] & sel_one_hot_i[52];
  assign data_masked[6752] = data_i[6752] & sel_one_hot_i[52];
  assign data_masked[6751] = data_i[6751] & sel_one_hot_i[52];
  assign data_masked[6750] = data_i[6750] & sel_one_hot_i[52];
  assign data_masked[6749] = data_i[6749] & sel_one_hot_i[52];
  assign data_masked[6748] = data_i[6748] & sel_one_hot_i[52];
  assign data_masked[6747] = data_i[6747] & sel_one_hot_i[52];
  assign data_masked[6746] = data_i[6746] & sel_one_hot_i[52];
  assign data_masked[6745] = data_i[6745] & sel_one_hot_i[52];
  assign data_masked[6744] = data_i[6744] & sel_one_hot_i[52];
  assign data_masked[6743] = data_i[6743] & sel_one_hot_i[52];
  assign data_masked[6742] = data_i[6742] & sel_one_hot_i[52];
  assign data_masked[6741] = data_i[6741] & sel_one_hot_i[52];
  assign data_masked[6740] = data_i[6740] & sel_one_hot_i[52];
  assign data_masked[6739] = data_i[6739] & sel_one_hot_i[52];
  assign data_masked[6738] = data_i[6738] & sel_one_hot_i[52];
  assign data_masked[6737] = data_i[6737] & sel_one_hot_i[52];
  assign data_masked[6736] = data_i[6736] & sel_one_hot_i[52];
  assign data_masked[6735] = data_i[6735] & sel_one_hot_i[52];
  assign data_masked[6734] = data_i[6734] & sel_one_hot_i[52];
  assign data_masked[6733] = data_i[6733] & sel_one_hot_i[52];
  assign data_masked[6732] = data_i[6732] & sel_one_hot_i[52];
  assign data_masked[6731] = data_i[6731] & sel_one_hot_i[52];
  assign data_masked[6730] = data_i[6730] & sel_one_hot_i[52];
  assign data_masked[6729] = data_i[6729] & sel_one_hot_i[52];
  assign data_masked[6728] = data_i[6728] & sel_one_hot_i[52];
  assign data_masked[6727] = data_i[6727] & sel_one_hot_i[52];
  assign data_masked[6726] = data_i[6726] & sel_one_hot_i[52];
  assign data_masked[6725] = data_i[6725] & sel_one_hot_i[52];
  assign data_masked[6724] = data_i[6724] & sel_one_hot_i[52];
  assign data_masked[6723] = data_i[6723] & sel_one_hot_i[52];
  assign data_masked[6722] = data_i[6722] & sel_one_hot_i[52];
  assign data_masked[6721] = data_i[6721] & sel_one_hot_i[52];
  assign data_masked[6720] = data_i[6720] & sel_one_hot_i[52];
  assign data_masked[6719] = data_i[6719] & sel_one_hot_i[52];
  assign data_masked[6718] = data_i[6718] & sel_one_hot_i[52];
  assign data_masked[6717] = data_i[6717] & sel_one_hot_i[52];
  assign data_masked[6716] = data_i[6716] & sel_one_hot_i[52];
  assign data_masked[6715] = data_i[6715] & sel_one_hot_i[52];
  assign data_masked[6714] = data_i[6714] & sel_one_hot_i[52];
  assign data_masked[6713] = data_i[6713] & sel_one_hot_i[52];
  assign data_masked[6712] = data_i[6712] & sel_one_hot_i[52];
  assign data_masked[6711] = data_i[6711] & sel_one_hot_i[52];
  assign data_masked[6710] = data_i[6710] & sel_one_hot_i[52];
  assign data_masked[6709] = data_i[6709] & sel_one_hot_i[52];
  assign data_masked[6708] = data_i[6708] & sel_one_hot_i[52];
  assign data_masked[6707] = data_i[6707] & sel_one_hot_i[52];
  assign data_masked[6706] = data_i[6706] & sel_one_hot_i[52];
  assign data_masked[6705] = data_i[6705] & sel_one_hot_i[52];
  assign data_masked[6704] = data_i[6704] & sel_one_hot_i[52];
  assign data_masked[6703] = data_i[6703] & sel_one_hot_i[52];
  assign data_masked[6702] = data_i[6702] & sel_one_hot_i[52];
  assign data_masked[6701] = data_i[6701] & sel_one_hot_i[52];
  assign data_masked[6700] = data_i[6700] & sel_one_hot_i[52];
  assign data_masked[6699] = data_i[6699] & sel_one_hot_i[52];
  assign data_masked[6698] = data_i[6698] & sel_one_hot_i[52];
  assign data_masked[6697] = data_i[6697] & sel_one_hot_i[52];
  assign data_masked[6696] = data_i[6696] & sel_one_hot_i[52];
  assign data_masked[6695] = data_i[6695] & sel_one_hot_i[52];
  assign data_masked[6694] = data_i[6694] & sel_one_hot_i[52];
  assign data_masked[6693] = data_i[6693] & sel_one_hot_i[52];
  assign data_masked[6692] = data_i[6692] & sel_one_hot_i[52];
  assign data_masked[6691] = data_i[6691] & sel_one_hot_i[52];
  assign data_masked[6690] = data_i[6690] & sel_one_hot_i[52];
  assign data_masked[6689] = data_i[6689] & sel_one_hot_i[52];
  assign data_masked[6688] = data_i[6688] & sel_one_hot_i[52];
  assign data_masked[6687] = data_i[6687] & sel_one_hot_i[52];
  assign data_masked[6686] = data_i[6686] & sel_one_hot_i[52];
  assign data_masked[6685] = data_i[6685] & sel_one_hot_i[52];
  assign data_masked[6684] = data_i[6684] & sel_one_hot_i[52];
  assign data_masked[6683] = data_i[6683] & sel_one_hot_i[52];
  assign data_masked[6682] = data_i[6682] & sel_one_hot_i[52];
  assign data_masked[6681] = data_i[6681] & sel_one_hot_i[52];
  assign data_masked[6680] = data_i[6680] & sel_one_hot_i[52];
  assign data_masked[6679] = data_i[6679] & sel_one_hot_i[52];
  assign data_masked[6678] = data_i[6678] & sel_one_hot_i[52];
  assign data_masked[6677] = data_i[6677] & sel_one_hot_i[52];
  assign data_masked[6676] = data_i[6676] & sel_one_hot_i[52];
  assign data_masked[6675] = data_i[6675] & sel_one_hot_i[52];
  assign data_masked[6674] = data_i[6674] & sel_one_hot_i[52];
  assign data_masked[6673] = data_i[6673] & sel_one_hot_i[52];
  assign data_masked[6672] = data_i[6672] & sel_one_hot_i[52];
  assign data_masked[6671] = data_i[6671] & sel_one_hot_i[52];
  assign data_masked[6670] = data_i[6670] & sel_one_hot_i[52];
  assign data_masked[6669] = data_i[6669] & sel_one_hot_i[52];
  assign data_masked[6668] = data_i[6668] & sel_one_hot_i[52];
  assign data_masked[6667] = data_i[6667] & sel_one_hot_i[52];
  assign data_masked[6666] = data_i[6666] & sel_one_hot_i[52];
  assign data_masked[6665] = data_i[6665] & sel_one_hot_i[52];
  assign data_masked[6664] = data_i[6664] & sel_one_hot_i[52];
  assign data_masked[6663] = data_i[6663] & sel_one_hot_i[52];
  assign data_masked[6662] = data_i[6662] & sel_one_hot_i[52];
  assign data_masked[6661] = data_i[6661] & sel_one_hot_i[52];
  assign data_masked[6660] = data_i[6660] & sel_one_hot_i[52];
  assign data_masked[6659] = data_i[6659] & sel_one_hot_i[52];
  assign data_masked[6658] = data_i[6658] & sel_one_hot_i[52];
  assign data_masked[6657] = data_i[6657] & sel_one_hot_i[52];
  assign data_masked[6656] = data_i[6656] & sel_one_hot_i[52];
  assign data_masked[6911] = data_i[6911] & sel_one_hot_i[53];
  assign data_masked[6910] = data_i[6910] & sel_one_hot_i[53];
  assign data_masked[6909] = data_i[6909] & sel_one_hot_i[53];
  assign data_masked[6908] = data_i[6908] & sel_one_hot_i[53];
  assign data_masked[6907] = data_i[6907] & sel_one_hot_i[53];
  assign data_masked[6906] = data_i[6906] & sel_one_hot_i[53];
  assign data_masked[6905] = data_i[6905] & sel_one_hot_i[53];
  assign data_masked[6904] = data_i[6904] & sel_one_hot_i[53];
  assign data_masked[6903] = data_i[6903] & sel_one_hot_i[53];
  assign data_masked[6902] = data_i[6902] & sel_one_hot_i[53];
  assign data_masked[6901] = data_i[6901] & sel_one_hot_i[53];
  assign data_masked[6900] = data_i[6900] & sel_one_hot_i[53];
  assign data_masked[6899] = data_i[6899] & sel_one_hot_i[53];
  assign data_masked[6898] = data_i[6898] & sel_one_hot_i[53];
  assign data_masked[6897] = data_i[6897] & sel_one_hot_i[53];
  assign data_masked[6896] = data_i[6896] & sel_one_hot_i[53];
  assign data_masked[6895] = data_i[6895] & sel_one_hot_i[53];
  assign data_masked[6894] = data_i[6894] & sel_one_hot_i[53];
  assign data_masked[6893] = data_i[6893] & sel_one_hot_i[53];
  assign data_masked[6892] = data_i[6892] & sel_one_hot_i[53];
  assign data_masked[6891] = data_i[6891] & sel_one_hot_i[53];
  assign data_masked[6890] = data_i[6890] & sel_one_hot_i[53];
  assign data_masked[6889] = data_i[6889] & sel_one_hot_i[53];
  assign data_masked[6888] = data_i[6888] & sel_one_hot_i[53];
  assign data_masked[6887] = data_i[6887] & sel_one_hot_i[53];
  assign data_masked[6886] = data_i[6886] & sel_one_hot_i[53];
  assign data_masked[6885] = data_i[6885] & sel_one_hot_i[53];
  assign data_masked[6884] = data_i[6884] & sel_one_hot_i[53];
  assign data_masked[6883] = data_i[6883] & sel_one_hot_i[53];
  assign data_masked[6882] = data_i[6882] & sel_one_hot_i[53];
  assign data_masked[6881] = data_i[6881] & sel_one_hot_i[53];
  assign data_masked[6880] = data_i[6880] & sel_one_hot_i[53];
  assign data_masked[6879] = data_i[6879] & sel_one_hot_i[53];
  assign data_masked[6878] = data_i[6878] & sel_one_hot_i[53];
  assign data_masked[6877] = data_i[6877] & sel_one_hot_i[53];
  assign data_masked[6876] = data_i[6876] & sel_one_hot_i[53];
  assign data_masked[6875] = data_i[6875] & sel_one_hot_i[53];
  assign data_masked[6874] = data_i[6874] & sel_one_hot_i[53];
  assign data_masked[6873] = data_i[6873] & sel_one_hot_i[53];
  assign data_masked[6872] = data_i[6872] & sel_one_hot_i[53];
  assign data_masked[6871] = data_i[6871] & sel_one_hot_i[53];
  assign data_masked[6870] = data_i[6870] & sel_one_hot_i[53];
  assign data_masked[6869] = data_i[6869] & sel_one_hot_i[53];
  assign data_masked[6868] = data_i[6868] & sel_one_hot_i[53];
  assign data_masked[6867] = data_i[6867] & sel_one_hot_i[53];
  assign data_masked[6866] = data_i[6866] & sel_one_hot_i[53];
  assign data_masked[6865] = data_i[6865] & sel_one_hot_i[53];
  assign data_masked[6864] = data_i[6864] & sel_one_hot_i[53];
  assign data_masked[6863] = data_i[6863] & sel_one_hot_i[53];
  assign data_masked[6862] = data_i[6862] & sel_one_hot_i[53];
  assign data_masked[6861] = data_i[6861] & sel_one_hot_i[53];
  assign data_masked[6860] = data_i[6860] & sel_one_hot_i[53];
  assign data_masked[6859] = data_i[6859] & sel_one_hot_i[53];
  assign data_masked[6858] = data_i[6858] & sel_one_hot_i[53];
  assign data_masked[6857] = data_i[6857] & sel_one_hot_i[53];
  assign data_masked[6856] = data_i[6856] & sel_one_hot_i[53];
  assign data_masked[6855] = data_i[6855] & sel_one_hot_i[53];
  assign data_masked[6854] = data_i[6854] & sel_one_hot_i[53];
  assign data_masked[6853] = data_i[6853] & sel_one_hot_i[53];
  assign data_masked[6852] = data_i[6852] & sel_one_hot_i[53];
  assign data_masked[6851] = data_i[6851] & sel_one_hot_i[53];
  assign data_masked[6850] = data_i[6850] & sel_one_hot_i[53];
  assign data_masked[6849] = data_i[6849] & sel_one_hot_i[53];
  assign data_masked[6848] = data_i[6848] & sel_one_hot_i[53];
  assign data_masked[6847] = data_i[6847] & sel_one_hot_i[53];
  assign data_masked[6846] = data_i[6846] & sel_one_hot_i[53];
  assign data_masked[6845] = data_i[6845] & sel_one_hot_i[53];
  assign data_masked[6844] = data_i[6844] & sel_one_hot_i[53];
  assign data_masked[6843] = data_i[6843] & sel_one_hot_i[53];
  assign data_masked[6842] = data_i[6842] & sel_one_hot_i[53];
  assign data_masked[6841] = data_i[6841] & sel_one_hot_i[53];
  assign data_masked[6840] = data_i[6840] & sel_one_hot_i[53];
  assign data_masked[6839] = data_i[6839] & sel_one_hot_i[53];
  assign data_masked[6838] = data_i[6838] & sel_one_hot_i[53];
  assign data_masked[6837] = data_i[6837] & sel_one_hot_i[53];
  assign data_masked[6836] = data_i[6836] & sel_one_hot_i[53];
  assign data_masked[6835] = data_i[6835] & sel_one_hot_i[53];
  assign data_masked[6834] = data_i[6834] & sel_one_hot_i[53];
  assign data_masked[6833] = data_i[6833] & sel_one_hot_i[53];
  assign data_masked[6832] = data_i[6832] & sel_one_hot_i[53];
  assign data_masked[6831] = data_i[6831] & sel_one_hot_i[53];
  assign data_masked[6830] = data_i[6830] & sel_one_hot_i[53];
  assign data_masked[6829] = data_i[6829] & sel_one_hot_i[53];
  assign data_masked[6828] = data_i[6828] & sel_one_hot_i[53];
  assign data_masked[6827] = data_i[6827] & sel_one_hot_i[53];
  assign data_masked[6826] = data_i[6826] & sel_one_hot_i[53];
  assign data_masked[6825] = data_i[6825] & sel_one_hot_i[53];
  assign data_masked[6824] = data_i[6824] & sel_one_hot_i[53];
  assign data_masked[6823] = data_i[6823] & sel_one_hot_i[53];
  assign data_masked[6822] = data_i[6822] & sel_one_hot_i[53];
  assign data_masked[6821] = data_i[6821] & sel_one_hot_i[53];
  assign data_masked[6820] = data_i[6820] & sel_one_hot_i[53];
  assign data_masked[6819] = data_i[6819] & sel_one_hot_i[53];
  assign data_masked[6818] = data_i[6818] & sel_one_hot_i[53];
  assign data_masked[6817] = data_i[6817] & sel_one_hot_i[53];
  assign data_masked[6816] = data_i[6816] & sel_one_hot_i[53];
  assign data_masked[6815] = data_i[6815] & sel_one_hot_i[53];
  assign data_masked[6814] = data_i[6814] & sel_one_hot_i[53];
  assign data_masked[6813] = data_i[6813] & sel_one_hot_i[53];
  assign data_masked[6812] = data_i[6812] & sel_one_hot_i[53];
  assign data_masked[6811] = data_i[6811] & sel_one_hot_i[53];
  assign data_masked[6810] = data_i[6810] & sel_one_hot_i[53];
  assign data_masked[6809] = data_i[6809] & sel_one_hot_i[53];
  assign data_masked[6808] = data_i[6808] & sel_one_hot_i[53];
  assign data_masked[6807] = data_i[6807] & sel_one_hot_i[53];
  assign data_masked[6806] = data_i[6806] & sel_one_hot_i[53];
  assign data_masked[6805] = data_i[6805] & sel_one_hot_i[53];
  assign data_masked[6804] = data_i[6804] & sel_one_hot_i[53];
  assign data_masked[6803] = data_i[6803] & sel_one_hot_i[53];
  assign data_masked[6802] = data_i[6802] & sel_one_hot_i[53];
  assign data_masked[6801] = data_i[6801] & sel_one_hot_i[53];
  assign data_masked[6800] = data_i[6800] & sel_one_hot_i[53];
  assign data_masked[6799] = data_i[6799] & sel_one_hot_i[53];
  assign data_masked[6798] = data_i[6798] & sel_one_hot_i[53];
  assign data_masked[6797] = data_i[6797] & sel_one_hot_i[53];
  assign data_masked[6796] = data_i[6796] & sel_one_hot_i[53];
  assign data_masked[6795] = data_i[6795] & sel_one_hot_i[53];
  assign data_masked[6794] = data_i[6794] & sel_one_hot_i[53];
  assign data_masked[6793] = data_i[6793] & sel_one_hot_i[53];
  assign data_masked[6792] = data_i[6792] & sel_one_hot_i[53];
  assign data_masked[6791] = data_i[6791] & sel_one_hot_i[53];
  assign data_masked[6790] = data_i[6790] & sel_one_hot_i[53];
  assign data_masked[6789] = data_i[6789] & sel_one_hot_i[53];
  assign data_masked[6788] = data_i[6788] & sel_one_hot_i[53];
  assign data_masked[6787] = data_i[6787] & sel_one_hot_i[53];
  assign data_masked[6786] = data_i[6786] & sel_one_hot_i[53];
  assign data_masked[6785] = data_i[6785] & sel_one_hot_i[53];
  assign data_masked[6784] = data_i[6784] & sel_one_hot_i[53];
  assign data_masked[7039] = data_i[7039] & sel_one_hot_i[54];
  assign data_masked[7038] = data_i[7038] & sel_one_hot_i[54];
  assign data_masked[7037] = data_i[7037] & sel_one_hot_i[54];
  assign data_masked[7036] = data_i[7036] & sel_one_hot_i[54];
  assign data_masked[7035] = data_i[7035] & sel_one_hot_i[54];
  assign data_masked[7034] = data_i[7034] & sel_one_hot_i[54];
  assign data_masked[7033] = data_i[7033] & sel_one_hot_i[54];
  assign data_masked[7032] = data_i[7032] & sel_one_hot_i[54];
  assign data_masked[7031] = data_i[7031] & sel_one_hot_i[54];
  assign data_masked[7030] = data_i[7030] & sel_one_hot_i[54];
  assign data_masked[7029] = data_i[7029] & sel_one_hot_i[54];
  assign data_masked[7028] = data_i[7028] & sel_one_hot_i[54];
  assign data_masked[7027] = data_i[7027] & sel_one_hot_i[54];
  assign data_masked[7026] = data_i[7026] & sel_one_hot_i[54];
  assign data_masked[7025] = data_i[7025] & sel_one_hot_i[54];
  assign data_masked[7024] = data_i[7024] & sel_one_hot_i[54];
  assign data_masked[7023] = data_i[7023] & sel_one_hot_i[54];
  assign data_masked[7022] = data_i[7022] & sel_one_hot_i[54];
  assign data_masked[7021] = data_i[7021] & sel_one_hot_i[54];
  assign data_masked[7020] = data_i[7020] & sel_one_hot_i[54];
  assign data_masked[7019] = data_i[7019] & sel_one_hot_i[54];
  assign data_masked[7018] = data_i[7018] & sel_one_hot_i[54];
  assign data_masked[7017] = data_i[7017] & sel_one_hot_i[54];
  assign data_masked[7016] = data_i[7016] & sel_one_hot_i[54];
  assign data_masked[7015] = data_i[7015] & sel_one_hot_i[54];
  assign data_masked[7014] = data_i[7014] & sel_one_hot_i[54];
  assign data_masked[7013] = data_i[7013] & sel_one_hot_i[54];
  assign data_masked[7012] = data_i[7012] & sel_one_hot_i[54];
  assign data_masked[7011] = data_i[7011] & sel_one_hot_i[54];
  assign data_masked[7010] = data_i[7010] & sel_one_hot_i[54];
  assign data_masked[7009] = data_i[7009] & sel_one_hot_i[54];
  assign data_masked[7008] = data_i[7008] & sel_one_hot_i[54];
  assign data_masked[7007] = data_i[7007] & sel_one_hot_i[54];
  assign data_masked[7006] = data_i[7006] & sel_one_hot_i[54];
  assign data_masked[7005] = data_i[7005] & sel_one_hot_i[54];
  assign data_masked[7004] = data_i[7004] & sel_one_hot_i[54];
  assign data_masked[7003] = data_i[7003] & sel_one_hot_i[54];
  assign data_masked[7002] = data_i[7002] & sel_one_hot_i[54];
  assign data_masked[7001] = data_i[7001] & sel_one_hot_i[54];
  assign data_masked[7000] = data_i[7000] & sel_one_hot_i[54];
  assign data_masked[6999] = data_i[6999] & sel_one_hot_i[54];
  assign data_masked[6998] = data_i[6998] & sel_one_hot_i[54];
  assign data_masked[6997] = data_i[6997] & sel_one_hot_i[54];
  assign data_masked[6996] = data_i[6996] & sel_one_hot_i[54];
  assign data_masked[6995] = data_i[6995] & sel_one_hot_i[54];
  assign data_masked[6994] = data_i[6994] & sel_one_hot_i[54];
  assign data_masked[6993] = data_i[6993] & sel_one_hot_i[54];
  assign data_masked[6992] = data_i[6992] & sel_one_hot_i[54];
  assign data_masked[6991] = data_i[6991] & sel_one_hot_i[54];
  assign data_masked[6990] = data_i[6990] & sel_one_hot_i[54];
  assign data_masked[6989] = data_i[6989] & sel_one_hot_i[54];
  assign data_masked[6988] = data_i[6988] & sel_one_hot_i[54];
  assign data_masked[6987] = data_i[6987] & sel_one_hot_i[54];
  assign data_masked[6986] = data_i[6986] & sel_one_hot_i[54];
  assign data_masked[6985] = data_i[6985] & sel_one_hot_i[54];
  assign data_masked[6984] = data_i[6984] & sel_one_hot_i[54];
  assign data_masked[6983] = data_i[6983] & sel_one_hot_i[54];
  assign data_masked[6982] = data_i[6982] & sel_one_hot_i[54];
  assign data_masked[6981] = data_i[6981] & sel_one_hot_i[54];
  assign data_masked[6980] = data_i[6980] & sel_one_hot_i[54];
  assign data_masked[6979] = data_i[6979] & sel_one_hot_i[54];
  assign data_masked[6978] = data_i[6978] & sel_one_hot_i[54];
  assign data_masked[6977] = data_i[6977] & sel_one_hot_i[54];
  assign data_masked[6976] = data_i[6976] & sel_one_hot_i[54];
  assign data_masked[6975] = data_i[6975] & sel_one_hot_i[54];
  assign data_masked[6974] = data_i[6974] & sel_one_hot_i[54];
  assign data_masked[6973] = data_i[6973] & sel_one_hot_i[54];
  assign data_masked[6972] = data_i[6972] & sel_one_hot_i[54];
  assign data_masked[6971] = data_i[6971] & sel_one_hot_i[54];
  assign data_masked[6970] = data_i[6970] & sel_one_hot_i[54];
  assign data_masked[6969] = data_i[6969] & sel_one_hot_i[54];
  assign data_masked[6968] = data_i[6968] & sel_one_hot_i[54];
  assign data_masked[6967] = data_i[6967] & sel_one_hot_i[54];
  assign data_masked[6966] = data_i[6966] & sel_one_hot_i[54];
  assign data_masked[6965] = data_i[6965] & sel_one_hot_i[54];
  assign data_masked[6964] = data_i[6964] & sel_one_hot_i[54];
  assign data_masked[6963] = data_i[6963] & sel_one_hot_i[54];
  assign data_masked[6962] = data_i[6962] & sel_one_hot_i[54];
  assign data_masked[6961] = data_i[6961] & sel_one_hot_i[54];
  assign data_masked[6960] = data_i[6960] & sel_one_hot_i[54];
  assign data_masked[6959] = data_i[6959] & sel_one_hot_i[54];
  assign data_masked[6958] = data_i[6958] & sel_one_hot_i[54];
  assign data_masked[6957] = data_i[6957] & sel_one_hot_i[54];
  assign data_masked[6956] = data_i[6956] & sel_one_hot_i[54];
  assign data_masked[6955] = data_i[6955] & sel_one_hot_i[54];
  assign data_masked[6954] = data_i[6954] & sel_one_hot_i[54];
  assign data_masked[6953] = data_i[6953] & sel_one_hot_i[54];
  assign data_masked[6952] = data_i[6952] & sel_one_hot_i[54];
  assign data_masked[6951] = data_i[6951] & sel_one_hot_i[54];
  assign data_masked[6950] = data_i[6950] & sel_one_hot_i[54];
  assign data_masked[6949] = data_i[6949] & sel_one_hot_i[54];
  assign data_masked[6948] = data_i[6948] & sel_one_hot_i[54];
  assign data_masked[6947] = data_i[6947] & sel_one_hot_i[54];
  assign data_masked[6946] = data_i[6946] & sel_one_hot_i[54];
  assign data_masked[6945] = data_i[6945] & sel_one_hot_i[54];
  assign data_masked[6944] = data_i[6944] & sel_one_hot_i[54];
  assign data_masked[6943] = data_i[6943] & sel_one_hot_i[54];
  assign data_masked[6942] = data_i[6942] & sel_one_hot_i[54];
  assign data_masked[6941] = data_i[6941] & sel_one_hot_i[54];
  assign data_masked[6940] = data_i[6940] & sel_one_hot_i[54];
  assign data_masked[6939] = data_i[6939] & sel_one_hot_i[54];
  assign data_masked[6938] = data_i[6938] & sel_one_hot_i[54];
  assign data_masked[6937] = data_i[6937] & sel_one_hot_i[54];
  assign data_masked[6936] = data_i[6936] & sel_one_hot_i[54];
  assign data_masked[6935] = data_i[6935] & sel_one_hot_i[54];
  assign data_masked[6934] = data_i[6934] & sel_one_hot_i[54];
  assign data_masked[6933] = data_i[6933] & sel_one_hot_i[54];
  assign data_masked[6932] = data_i[6932] & sel_one_hot_i[54];
  assign data_masked[6931] = data_i[6931] & sel_one_hot_i[54];
  assign data_masked[6930] = data_i[6930] & sel_one_hot_i[54];
  assign data_masked[6929] = data_i[6929] & sel_one_hot_i[54];
  assign data_masked[6928] = data_i[6928] & sel_one_hot_i[54];
  assign data_masked[6927] = data_i[6927] & sel_one_hot_i[54];
  assign data_masked[6926] = data_i[6926] & sel_one_hot_i[54];
  assign data_masked[6925] = data_i[6925] & sel_one_hot_i[54];
  assign data_masked[6924] = data_i[6924] & sel_one_hot_i[54];
  assign data_masked[6923] = data_i[6923] & sel_one_hot_i[54];
  assign data_masked[6922] = data_i[6922] & sel_one_hot_i[54];
  assign data_masked[6921] = data_i[6921] & sel_one_hot_i[54];
  assign data_masked[6920] = data_i[6920] & sel_one_hot_i[54];
  assign data_masked[6919] = data_i[6919] & sel_one_hot_i[54];
  assign data_masked[6918] = data_i[6918] & sel_one_hot_i[54];
  assign data_masked[6917] = data_i[6917] & sel_one_hot_i[54];
  assign data_masked[6916] = data_i[6916] & sel_one_hot_i[54];
  assign data_masked[6915] = data_i[6915] & sel_one_hot_i[54];
  assign data_masked[6914] = data_i[6914] & sel_one_hot_i[54];
  assign data_masked[6913] = data_i[6913] & sel_one_hot_i[54];
  assign data_masked[6912] = data_i[6912] & sel_one_hot_i[54];
  assign data_masked[7167] = data_i[7167] & sel_one_hot_i[55];
  assign data_masked[7166] = data_i[7166] & sel_one_hot_i[55];
  assign data_masked[7165] = data_i[7165] & sel_one_hot_i[55];
  assign data_masked[7164] = data_i[7164] & sel_one_hot_i[55];
  assign data_masked[7163] = data_i[7163] & sel_one_hot_i[55];
  assign data_masked[7162] = data_i[7162] & sel_one_hot_i[55];
  assign data_masked[7161] = data_i[7161] & sel_one_hot_i[55];
  assign data_masked[7160] = data_i[7160] & sel_one_hot_i[55];
  assign data_masked[7159] = data_i[7159] & sel_one_hot_i[55];
  assign data_masked[7158] = data_i[7158] & sel_one_hot_i[55];
  assign data_masked[7157] = data_i[7157] & sel_one_hot_i[55];
  assign data_masked[7156] = data_i[7156] & sel_one_hot_i[55];
  assign data_masked[7155] = data_i[7155] & sel_one_hot_i[55];
  assign data_masked[7154] = data_i[7154] & sel_one_hot_i[55];
  assign data_masked[7153] = data_i[7153] & sel_one_hot_i[55];
  assign data_masked[7152] = data_i[7152] & sel_one_hot_i[55];
  assign data_masked[7151] = data_i[7151] & sel_one_hot_i[55];
  assign data_masked[7150] = data_i[7150] & sel_one_hot_i[55];
  assign data_masked[7149] = data_i[7149] & sel_one_hot_i[55];
  assign data_masked[7148] = data_i[7148] & sel_one_hot_i[55];
  assign data_masked[7147] = data_i[7147] & sel_one_hot_i[55];
  assign data_masked[7146] = data_i[7146] & sel_one_hot_i[55];
  assign data_masked[7145] = data_i[7145] & sel_one_hot_i[55];
  assign data_masked[7144] = data_i[7144] & sel_one_hot_i[55];
  assign data_masked[7143] = data_i[7143] & sel_one_hot_i[55];
  assign data_masked[7142] = data_i[7142] & sel_one_hot_i[55];
  assign data_masked[7141] = data_i[7141] & sel_one_hot_i[55];
  assign data_masked[7140] = data_i[7140] & sel_one_hot_i[55];
  assign data_masked[7139] = data_i[7139] & sel_one_hot_i[55];
  assign data_masked[7138] = data_i[7138] & sel_one_hot_i[55];
  assign data_masked[7137] = data_i[7137] & sel_one_hot_i[55];
  assign data_masked[7136] = data_i[7136] & sel_one_hot_i[55];
  assign data_masked[7135] = data_i[7135] & sel_one_hot_i[55];
  assign data_masked[7134] = data_i[7134] & sel_one_hot_i[55];
  assign data_masked[7133] = data_i[7133] & sel_one_hot_i[55];
  assign data_masked[7132] = data_i[7132] & sel_one_hot_i[55];
  assign data_masked[7131] = data_i[7131] & sel_one_hot_i[55];
  assign data_masked[7130] = data_i[7130] & sel_one_hot_i[55];
  assign data_masked[7129] = data_i[7129] & sel_one_hot_i[55];
  assign data_masked[7128] = data_i[7128] & sel_one_hot_i[55];
  assign data_masked[7127] = data_i[7127] & sel_one_hot_i[55];
  assign data_masked[7126] = data_i[7126] & sel_one_hot_i[55];
  assign data_masked[7125] = data_i[7125] & sel_one_hot_i[55];
  assign data_masked[7124] = data_i[7124] & sel_one_hot_i[55];
  assign data_masked[7123] = data_i[7123] & sel_one_hot_i[55];
  assign data_masked[7122] = data_i[7122] & sel_one_hot_i[55];
  assign data_masked[7121] = data_i[7121] & sel_one_hot_i[55];
  assign data_masked[7120] = data_i[7120] & sel_one_hot_i[55];
  assign data_masked[7119] = data_i[7119] & sel_one_hot_i[55];
  assign data_masked[7118] = data_i[7118] & sel_one_hot_i[55];
  assign data_masked[7117] = data_i[7117] & sel_one_hot_i[55];
  assign data_masked[7116] = data_i[7116] & sel_one_hot_i[55];
  assign data_masked[7115] = data_i[7115] & sel_one_hot_i[55];
  assign data_masked[7114] = data_i[7114] & sel_one_hot_i[55];
  assign data_masked[7113] = data_i[7113] & sel_one_hot_i[55];
  assign data_masked[7112] = data_i[7112] & sel_one_hot_i[55];
  assign data_masked[7111] = data_i[7111] & sel_one_hot_i[55];
  assign data_masked[7110] = data_i[7110] & sel_one_hot_i[55];
  assign data_masked[7109] = data_i[7109] & sel_one_hot_i[55];
  assign data_masked[7108] = data_i[7108] & sel_one_hot_i[55];
  assign data_masked[7107] = data_i[7107] & sel_one_hot_i[55];
  assign data_masked[7106] = data_i[7106] & sel_one_hot_i[55];
  assign data_masked[7105] = data_i[7105] & sel_one_hot_i[55];
  assign data_masked[7104] = data_i[7104] & sel_one_hot_i[55];
  assign data_masked[7103] = data_i[7103] & sel_one_hot_i[55];
  assign data_masked[7102] = data_i[7102] & sel_one_hot_i[55];
  assign data_masked[7101] = data_i[7101] & sel_one_hot_i[55];
  assign data_masked[7100] = data_i[7100] & sel_one_hot_i[55];
  assign data_masked[7099] = data_i[7099] & sel_one_hot_i[55];
  assign data_masked[7098] = data_i[7098] & sel_one_hot_i[55];
  assign data_masked[7097] = data_i[7097] & sel_one_hot_i[55];
  assign data_masked[7096] = data_i[7096] & sel_one_hot_i[55];
  assign data_masked[7095] = data_i[7095] & sel_one_hot_i[55];
  assign data_masked[7094] = data_i[7094] & sel_one_hot_i[55];
  assign data_masked[7093] = data_i[7093] & sel_one_hot_i[55];
  assign data_masked[7092] = data_i[7092] & sel_one_hot_i[55];
  assign data_masked[7091] = data_i[7091] & sel_one_hot_i[55];
  assign data_masked[7090] = data_i[7090] & sel_one_hot_i[55];
  assign data_masked[7089] = data_i[7089] & sel_one_hot_i[55];
  assign data_masked[7088] = data_i[7088] & sel_one_hot_i[55];
  assign data_masked[7087] = data_i[7087] & sel_one_hot_i[55];
  assign data_masked[7086] = data_i[7086] & sel_one_hot_i[55];
  assign data_masked[7085] = data_i[7085] & sel_one_hot_i[55];
  assign data_masked[7084] = data_i[7084] & sel_one_hot_i[55];
  assign data_masked[7083] = data_i[7083] & sel_one_hot_i[55];
  assign data_masked[7082] = data_i[7082] & sel_one_hot_i[55];
  assign data_masked[7081] = data_i[7081] & sel_one_hot_i[55];
  assign data_masked[7080] = data_i[7080] & sel_one_hot_i[55];
  assign data_masked[7079] = data_i[7079] & sel_one_hot_i[55];
  assign data_masked[7078] = data_i[7078] & sel_one_hot_i[55];
  assign data_masked[7077] = data_i[7077] & sel_one_hot_i[55];
  assign data_masked[7076] = data_i[7076] & sel_one_hot_i[55];
  assign data_masked[7075] = data_i[7075] & sel_one_hot_i[55];
  assign data_masked[7074] = data_i[7074] & sel_one_hot_i[55];
  assign data_masked[7073] = data_i[7073] & sel_one_hot_i[55];
  assign data_masked[7072] = data_i[7072] & sel_one_hot_i[55];
  assign data_masked[7071] = data_i[7071] & sel_one_hot_i[55];
  assign data_masked[7070] = data_i[7070] & sel_one_hot_i[55];
  assign data_masked[7069] = data_i[7069] & sel_one_hot_i[55];
  assign data_masked[7068] = data_i[7068] & sel_one_hot_i[55];
  assign data_masked[7067] = data_i[7067] & sel_one_hot_i[55];
  assign data_masked[7066] = data_i[7066] & sel_one_hot_i[55];
  assign data_masked[7065] = data_i[7065] & sel_one_hot_i[55];
  assign data_masked[7064] = data_i[7064] & sel_one_hot_i[55];
  assign data_masked[7063] = data_i[7063] & sel_one_hot_i[55];
  assign data_masked[7062] = data_i[7062] & sel_one_hot_i[55];
  assign data_masked[7061] = data_i[7061] & sel_one_hot_i[55];
  assign data_masked[7060] = data_i[7060] & sel_one_hot_i[55];
  assign data_masked[7059] = data_i[7059] & sel_one_hot_i[55];
  assign data_masked[7058] = data_i[7058] & sel_one_hot_i[55];
  assign data_masked[7057] = data_i[7057] & sel_one_hot_i[55];
  assign data_masked[7056] = data_i[7056] & sel_one_hot_i[55];
  assign data_masked[7055] = data_i[7055] & sel_one_hot_i[55];
  assign data_masked[7054] = data_i[7054] & sel_one_hot_i[55];
  assign data_masked[7053] = data_i[7053] & sel_one_hot_i[55];
  assign data_masked[7052] = data_i[7052] & sel_one_hot_i[55];
  assign data_masked[7051] = data_i[7051] & sel_one_hot_i[55];
  assign data_masked[7050] = data_i[7050] & sel_one_hot_i[55];
  assign data_masked[7049] = data_i[7049] & sel_one_hot_i[55];
  assign data_masked[7048] = data_i[7048] & sel_one_hot_i[55];
  assign data_masked[7047] = data_i[7047] & sel_one_hot_i[55];
  assign data_masked[7046] = data_i[7046] & sel_one_hot_i[55];
  assign data_masked[7045] = data_i[7045] & sel_one_hot_i[55];
  assign data_masked[7044] = data_i[7044] & sel_one_hot_i[55];
  assign data_masked[7043] = data_i[7043] & sel_one_hot_i[55];
  assign data_masked[7042] = data_i[7042] & sel_one_hot_i[55];
  assign data_masked[7041] = data_i[7041] & sel_one_hot_i[55];
  assign data_masked[7040] = data_i[7040] & sel_one_hot_i[55];
  assign data_masked[7295] = data_i[7295] & sel_one_hot_i[56];
  assign data_masked[7294] = data_i[7294] & sel_one_hot_i[56];
  assign data_masked[7293] = data_i[7293] & sel_one_hot_i[56];
  assign data_masked[7292] = data_i[7292] & sel_one_hot_i[56];
  assign data_masked[7291] = data_i[7291] & sel_one_hot_i[56];
  assign data_masked[7290] = data_i[7290] & sel_one_hot_i[56];
  assign data_masked[7289] = data_i[7289] & sel_one_hot_i[56];
  assign data_masked[7288] = data_i[7288] & sel_one_hot_i[56];
  assign data_masked[7287] = data_i[7287] & sel_one_hot_i[56];
  assign data_masked[7286] = data_i[7286] & sel_one_hot_i[56];
  assign data_masked[7285] = data_i[7285] & sel_one_hot_i[56];
  assign data_masked[7284] = data_i[7284] & sel_one_hot_i[56];
  assign data_masked[7283] = data_i[7283] & sel_one_hot_i[56];
  assign data_masked[7282] = data_i[7282] & sel_one_hot_i[56];
  assign data_masked[7281] = data_i[7281] & sel_one_hot_i[56];
  assign data_masked[7280] = data_i[7280] & sel_one_hot_i[56];
  assign data_masked[7279] = data_i[7279] & sel_one_hot_i[56];
  assign data_masked[7278] = data_i[7278] & sel_one_hot_i[56];
  assign data_masked[7277] = data_i[7277] & sel_one_hot_i[56];
  assign data_masked[7276] = data_i[7276] & sel_one_hot_i[56];
  assign data_masked[7275] = data_i[7275] & sel_one_hot_i[56];
  assign data_masked[7274] = data_i[7274] & sel_one_hot_i[56];
  assign data_masked[7273] = data_i[7273] & sel_one_hot_i[56];
  assign data_masked[7272] = data_i[7272] & sel_one_hot_i[56];
  assign data_masked[7271] = data_i[7271] & sel_one_hot_i[56];
  assign data_masked[7270] = data_i[7270] & sel_one_hot_i[56];
  assign data_masked[7269] = data_i[7269] & sel_one_hot_i[56];
  assign data_masked[7268] = data_i[7268] & sel_one_hot_i[56];
  assign data_masked[7267] = data_i[7267] & sel_one_hot_i[56];
  assign data_masked[7266] = data_i[7266] & sel_one_hot_i[56];
  assign data_masked[7265] = data_i[7265] & sel_one_hot_i[56];
  assign data_masked[7264] = data_i[7264] & sel_one_hot_i[56];
  assign data_masked[7263] = data_i[7263] & sel_one_hot_i[56];
  assign data_masked[7262] = data_i[7262] & sel_one_hot_i[56];
  assign data_masked[7261] = data_i[7261] & sel_one_hot_i[56];
  assign data_masked[7260] = data_i[7260] & sel_one_hot_i[56];
  assign data_masked[7259] = data_i[7259] & sel_one_hot_i[56];
  assign data_masked[7258] = data_i[7258] & sel_one_hot_i[56];
  assign data_masked[7257] = data_i[7257] & sel_one_hot_i[56];
  assign data_masked[7256] = data_i[7256] & sel_one_hot_i[56];
  assign data_masked[7255] = data_i[7255] & sel_one_hot_i[56];
  assign data_masked[7254] = data_i[7254] & sel_one_hot_i[56];
  assign data_masked[7253] = data_i[7253] & sel_one_hot_i[56];
  assign data_masked[7252] = data_i[7252] & sel_one_hot_i[56];
  assign data_masked[7251] = data_i[7251] & sel_one_hot_i[56];
  assign data_masked[7250] = data_i[7250] & sel_one_hot_i[56];
  assign data_masked[7249] = data_i[7249] & sel_one_hot_i[56];
  assign data_masked[7248] = data_i[7248] & sel_one_hot_i[56];
  assign data_masked[7247] = data_i[7247] & sel_one_hot_i[56];
  assign data_masked[7246] = data_i[7246] & sel_one_hot_i[56];
  assign data_masked[7245] = data_i[7245] & sel_one_hot_i[56];
  assign data_masked[7244] = data_i[7244] & sel_one_hot_i[56];
  assign data_masked[7243] = data_i[7243] & sel_one_hot_i[56];
  assign data_masked[7242] = data_i[7242] & sel_one_hot_i[56];
  assign data_masked[7241] = data_i[7241] & sel_one_hot_i[56];
  assign data_masked[7240] = data_i[7240] & sel_one_hot_i[56];
  assign data_masked[7239] = data_i[7239] & sel_one_hot_i[56];
  assign data_masked[7238] = data_i[7238] & sel_one_hot_i[56];
  assign data_masked[7237] = data_i[7237] & sel_one_hot_i[56];
  assign data_masked[7236] = data_i[7236] & sel_one_hot_i[56];
  assign data_masked[7235] = data_i[7235] & sel_one_hot_i[56];
  assign data_masked[7234] = data_i[7234] & sel_one_hot_i[56];
  assign data_masked[7233] = data_i[7233] & sel_one_hot_i[56];
  assign data_masked[7232] = data_i[7232] & sel_one_hot_i[56];
  assign data_masked[7231] = data_i[7231] & sel_one_hot_i[56];
  assign data_masked[7230] = data_i[7230] & sel_one_hot_i[56];
  assign data_masked[7229] = data_i[7229] & sel_one_hot_i[56];
  assign data_masked[7228] = data_i[7228] & sel_one_hot_i[56];
  assign data_masked[7227] = data_i[7227] & sel_one_hot_i[56];
  assign data_masked[7226] = data_i[7226] & sel_one_hot_i[56];
  assign data_masked[7225] = data_i[7225] & sel_one_hot_i[56];
  assign data_masked[7224] = data_i[7224] & sel_one_hot_i[56];
  assign data_masked[7223] = data_i[7223] & sel_one_hot_i[56];
  assign data_masked[7222] = data_i[7222] & sel_one_hot_i[56];
  assign data_masked[7221] = data_i[7221] & sel_one_hot_i[56];
  assign data_masked[7220] = data_i[7220] & sel_one_hot_i[56];
  assign data_masked[7219] = data_i[7219] & sel_one_hot_i[56];
  assign data_masked[7218] = data_i[7218] & sel_one_hot_i[56];
  assign data_masked[7217] = data_i[7217] & sel_one_hot_i[56];
  assign data_masked[7216] = data_i[7216] & sel_one_hot_i[56];
  assign data_masked[7215] = data_i[7215] & sel_one_hot_i[56];
  assign data_masked[7214] = data_i[7214] & sel_one_hot_i[56];
  assign data_masked[7213] = data_i[7213] & sel_one_hot_i[56];
  assign data_masked[7212] = data_i[7212] & sel_one_hot_i[56];
  assign data_masked[7211] = data_i[7211] & sel_one_hot_i[56];
  assign data_masked[7210] = data_i[7210] & sel_one_hot_i[56];
  assign data_masked[7209] = data_i[7209] & sel_one_hot_i[56];
  assign data_masked[7208] = data_i[7208] & sel_one_hot_i[56];
  assign data_masked[7207] = data_i[7207] & sel_one_hot_i[56];
  assign data_masked[7206] = data_i[7206] & sel_one_hot_i[56];
  assign data_masked[7205] = data_i[7205] & sel_one_hot_i[56];
  assign data_masked[7204] = data_i[7204] & sel_one_hot_i[56];
  assign data_masked[7203] = data_i[7203] & sel_one_hot_i[56];
  assign data_masked[7202] = data_i[7202] & sel_one_hot_i[56];
  assign data_masked[7201] = data_i[7201] & sel_one_hot_i[56];
  assign data_masked[7200] = data_i[7200] & sel_one_hot_i[56];
  assign data_masked[7199] = data_i[7199] & sel_one_hot_i[56];
  assign data_masked[7198] = data_i[7198] & sel_one_hot_i[56];
  assign data_masked[7197] = data_i[7197] & sel_one_hot_i[56];
  assign data_masked[7196] = data_i[7196] & sel_one_hot_i[56];
  assign data_masked[7195] = data_i[7195] & sel_one_hot_i[56];
  assign data_masked[7194] = data_i[7194] & sel_one_hot_i[56];
  assign data_masked[7193] = data_i[7193] & sel_one_hot_i[56];
  assign data_masked[7192] = data_i[7192] & sel_one_hot_i[56];
  assign data_masked[7191] = data_i[7191] & sel_one_hot_i[56];
  assign data_masked[7190] = data_i[7190] & sel_one_hot_i[56];
  assign data_masked[7189] = data_i[7189] & sel_one_hot_i[56];
  assign data_masked[7188] = data_i[7188] & sel_one_hot_i[56];
  assign data_masked[7187] = data_i[7187] & sel_one_hot_i[56];
  assign data_masked[7186] = data_i[7186] & sel_one_hot_i[56];
  assign data_masked[7185] = data_i[7185] & sel_one_hot_i[56];
  assign data_masked[7184] = data_i[7184] & sel_one_hot_i[56];
  assign data_masked[7183] = data_i[7183] & sel_one_hot_i[56];
  assign data_masked[7182] = data_i[7182] & sel_one_hot_i[56];
  assign data_masked[7181] = data_i[7181] & sel_one_hot_i[56];
  assign data_masked[7180] = data_i[7180] & sel_one_hot_i[56];
  assign data_masked[7179] = data_i[7179] & sel_one_hot_i[56];
  assign data_masked[7178] = data_i[7178] & sel_one_hot_i[56];
  assign data_masked[7177] = data_i[7177] & sel_one_hot_i[56];
  assign data_masked[7176] = data_i[7176] & sel_one_hot_i[56];
  assign data_masked[7175] = data_i[7175] & sel_one_hot_i[56];
  assign data_masked[7174] = data_i[7174] & sel_one_hot_i[56];
  assign data_masked[7173] = data_i[7173] & sel_one_hot_i[56];
  assign data_masked[7172] = data_i[7172] & sel_one_hot_i[56];
  assign data_masked[7171] = data_i[7171] & sel_one_hot_i[56];
  assign data_masked[7170] = data_i[7170] & sel_one_hot_i[56];
  assign data_masked[7169] = data_i[7169] & sel_one_hot_i[56];
  assign data_masked[7168] = data_i[7168] & sel_one_hot_i[56];
  assign data_masked[7423] = data_i[7423] & sel_one_hot_i[57];
  assign data_masked[7422] = data_i[7422] & sel_one_hot_i[57];
  assign data_masked[7421] = data_i[7421] & sel_one_hot_i[57];
  assign data_masked[7420] = data_i[7420] & sel_one_hot_i[57];
  assign data_masked[7419] = data_i[7419] & sel_one_hot_i[57];
  assign data_masked[7418] = data_i[7418] & sel_one_hot_i[57];
  assign data_masked[7417] = data_i[7417] & sel_one_hot_i[57];
  assign data_masked[7416] = data_i[7416] & sel_one_hot_i[57];
  assign data_masked[7415] = data_i[7415] & sel_one_hot_i[57];
  assign data_masked[7414] = data_i[7414] & sel_one_hot_i[57];
  assign data_masked[7413] = data_i[7413] & sel_one_hot_i[57];
  assign data_masked[7412] = data_i[7412] & sel_one_hot_i[57];
  assign data_masked[7411] = data_i[7411] & sel_one_hot_i[57];
  assign data_masked[7410] = data_i[7410] & sel_one_hot_i[57];
  assign data_masked[7409] = data_i[7409] & sel_one_hot_i[57];
  assign data_masked[7408] = data_i[7408] & sel_one_hot_i[57];
  assign data_masked[7407] = data_i[7407] & sel_one_hot_i[57];
  assign data_masked[7406] = data_i[7406] & sel_one_hot_i[57];
  assign data_masked[7405] = data_i[7405] & sel_one_hot_i[57];
  assign data_masked[7404] = data_i[7404] & sel_one_hot_i[57];
  assign data_masked[7403] = data_i[7403] & sel_one_hot_i[57];
  assign data_masked[7402] = data_i[7402] & sel_one_hot_i[57];
  assign data_masked[7401] = data_i[7401] & sel_one_hot_i[57];
  assign data_masked[7400] = data_i[7400] & sel_one_hot_i[57];
  assign data_masked[7399] = data_i[7399] & sel_one_hot_i[57];
  assign data_masked[7398] = data_i[7398] & sel_one_hot_i[57];
  assign data_masked[7397] = data_i[7397] & sel_one_hot_i[57];
  assign data_masked[7396] = data_i[7396] & sel_one_hot_i[57];
  assign data_masked[7395] = data_i[7395] & sel_one_hot_i[57];
  assign data_masked[7394] = data_i[7394] & sel_one_hot_i[57];
  assign data_masked[7393] = data_i[7393] & sel_one_hot_i[57];
  assign data_masked[7392] = data_i[7392] & sel_one_hot_i[57];
  assign data_masked[7391] = data_i[7391] & sel_one_hot_i[57];
  assign data_masked[7390] = data_i[7390] & sel_one_hot_i[57];
  assign data_masked[7389] = data_i[7389] & sel_one_hot_i[57];
  assign data_masked[7388] = data_i[7388] & sel_one_hot_i[57];
  assign data_masked[7387] = data_i[7387] & sel_one_hot_i[57];
  assign data_masked[7386] = data_i[7386] & sel_one_hot_i[57];
  assign data_masked[7385] = data_i[7385] & sel_one_hot_i[57];
  assign data_masked[7384] = data_i[7384] & sel_one_hot_i[57];
  assign data_masked[7383] = data_i[7383] & sel_one_hot_i[57];
  assign data_masked[7382] = data_i[7382] & sel_one_hot_i[57];
  assign data_masked[7381] = data_i[7381] & sel_one_hot_i[57];
  assign data_masked[7380] = data_i[7380] & sel_one_hot_i[57];
  assign data_masked[7379] = data_i[7379] & sel_one_hot_i[57];
  assign data_masked[7378] = data_i[7378] & sel_one_hot_i[57];
  assign data_masked[7377] = data_i[7377] & sel_one_hot_i[57];
  assign data_masked[7376] = data_i[7376] & sel_one_hot_i[57];
  assign data_masked[7375] = data_i[7375] & sel_one_hot_i[57];
  assign data_masked[7374] = data_i[7374] & sel_one_hot_i[57];
  assign data_masked[7373] = data_i[7373] & sel_one_hot_i[57];
  assign data_masked[7372] = data_i[7372] & sel_one_hot_i[57];
  assign data_masked[7371] = data_i[7371] & sel_one_hot_i[57];
  assign data_masked[7370] = data_i[7370] & sel_one_hot_i[57];
  assign data_masked[7369] = data_i[7369] & sel_one_hot_i[57];
  assign data_masked[7368] = data_i[7368] & sel_one_hot_i[57];
  assign data_masked[7367] = data_i[7367] & sel_one_hot_i[57];
  assign data_masked[7366] = data_i[7366] & sel_one_hot_i[57];
  assign data_masked[7365] = data_i[7365] & sel_one_hot_i[57];
  assign data_masked[7364] = data_i[7364] & sel_one_hot_i[57];
  assign data_masked[7363] = data_i[7363] & sel_one_hot_i[57];
  assign data_masked[7362] = data_i[7362] & sel_one_hot_i[57];
  assign data_masked[7361] = data_i[7361] & sel_one_hot_i[57];
  assign data_masked[7360] = data_i[7360] & sel_one_hot_i[57];
  assign data_masked[7359] = data_i[7359] & sel_one_hot_i[57];
  assign data_masked[7358] = data_i[7358] & sel_one_hot_i[57];
  assign data_masked[7357] = data_i[7357] & sel_one_hot_i[57];
  assign data_masked[7356] = data_i[7356] & sel_one_hot_i[57];
  assign data_masked[7355] = data_i[7355] & sel_one_hot_i[57];
  assign data_masked[7354] = data_i[7354] & sel_one_hot_i[57];
  assign data_masked[7353] = data_i[7353] & sel_one_hot_i[57];
  assign data_masked[7352] = data_i[7352] & sel_one_hot_i[57];
  assign data_masked[7351] = data_i[7351] & sel_one_hot_i[57];
  assign data_masked[7350] = data_i[7350] & sel_one_hot_i[57];
  assign data_masked[7349] = data_i[7349] & sel_one_hot_i[57];
  assign data_masked[7348] = data_i[7348] & sel_one_hot_i[57];
  assign data_masked[7347] = data_i[7347] & sel_one_hot_i[57];
  assign data_masked[7346] = data_i[7346] & sel_one_hot_i[57];
  assign data_masked[7345] = data_i[7345] & sel_one_hot_i[57];
  assign data_masked[7344] = data_i[7344] & sel_one_hot_i[57];
  assign data_masked[7343] = data_i[7343] & sel_one_hot_i[57];
  assign data_masked[7342] = data_i[7342] & sel_one_hot_i[57];
  assign data_masked[7341] = data_i[7341] & sel_one_hot_i[57];
  assign data_masked[7340] = data_i[7340] & sel_one_hot_i[57];
  assign data_masked[7339] = data_i[7339] & sel_one_hot_i[57];
  assign data_masked[7338] = data_i[7338] & sel_one_hot_i[57];
  assign data_masked[7337] = data_i[7337] & sel_one_hot_i[57];
  assign data_masked[7336] = data_i[7336] & sel_one_hot_i[57];
  assign data_masked[7335] = data_i[7335] & sel_one_hot_i[57];
  assign data_masked[7334] = data_i[7334] & sel_one_hot_i[57];
  assign data_masked[7333] = data_i[7333] & sel_one_hot_i[57];
  assign data_masked[7332] = data_i[7332] & sel_one_hot_i[57];
  assign data_masked[7331] = data_i[7331] & sel_one_hot_i[57];
  assign data_masked[7330] = data_i[7330] & sel_one_hot_i[57];
  assign data_masked[7329] = data_i[7329] & sel_one_hot_i[57];
  assign data_masked[7328] = data_i[7328] & sel_one_hot_i[57];
  assign data_masked[7327] = data_i[7327] & sel_one_hot_i[57];
  assign data_masked[7326] = data_i[7326] & sel_one_hot_i[57];
  assign data_masked[7325] = data_i[7325] & sel_one_hot_i[57];
  assign data_masked[7324] = data_i[7324] & sel_one_hot_i[57];
  assign data_masked[7323] = data_i[7323] & sel_one_hot_i[57];
  assign data_masked[7322] = data_i[7322] & sel_one_hot_i[57];
  assign data_masked[7321] = data_i[7321] & sel_one_hot_i[57];
  assign data_masked[7320] = data_i[7320] & sel_one_hot_i[57];
  assign data_masked[7319] = data_i[7319] & sel_one_hot_i[57];
  assign data_masked[7318] = data_i[7318] & sel_one_hot_i[57];
  assign data_masked[7317] = data_i[7317] & sel_one_hot_i[57];
  assign data_masked[7316] = data_i[7316] & sel_one_hot_i[57];
  assign data_masked[7315] = data_i[7315] & sel_one_hot_i[57];
  assign data_masked[7314] = data_i[7314] & sel_one_hot_i[57];
  assign data_masked[7313] = data_i[7313] & sel_one_hot_i[57];
  assign data_masked[7312] = data_i[7312] & sel_one_hot_i[57];
  assign data_masked[7311] = data_i[7311] & sel_one_hot_i[57];
  assign data_masked[7310] = data_i[7310] & sel_one_hot_i[57];
  assign data_masked[7309] = data_i[7309] & sel_one_hot_i[57];
  assign data_masked[7308] = data_i[7308] & sel_one_hot_i[57];
  assign data_masked[7307] = data_i[7307] & sel_one_hot_i[57];
  assign data_masked[7306] = data_i[7306] & sel_one_hot_i[57];
  assign data_masked[7305] = data_i[7305] & sel_one_hot_i[57];
  assign data_masked[7304] = data_i[7304] & sel_one_hot_i[57];
  assign data_masked[7303] = data_i[7303] & sel_one_hot_i[57];
  assign data_masked[7302] = data_i[7302] & sel_one_hot_i[57];
  assign data_masked[7301] = data_i[7301] & sel_one_hot_i[57];
  assign data_masked[7300] = data_i[7300] & sel_one_hot_i[57];
  assign data_masked[7299] = data_i[7299] & sel_one_hot_i[57];
  assign data_masked[7298] = data_i[7298] & sel_one_hot_i[57];
  assign data_masked[7297] = data_i[7297] & sel_one_hot_i[57];
  assign data_masked[7296] = data_i[7296] & sel_one_hot_i[57];
  assign data_masked[7551] = data_i[7551] & sel_one_hot_i[58];
  assign data_masked[7550] = data_i[7550] & sel_one_hot_i[58];
  assign data_masked[7549] = data_i[7549] & sel_one_hot_i[58];
  assign data_masked[7548] = data_i[7548] & sel_one_hot_i[58];
  assign data_masked[7547] = data_i[7547] & sel_one_hot_i[58];
  assign data_masked[7546] = data_i[7546] & sel_one_hot_i[58];
  assign data_masked[7545] = data_i[7545] & sel_one_hot_i[58];
  assign data_masked[7544] = data_i[7544] & sel_one_hot_i[58];
  assign data_masked[7543] = data_i[7543] & sel_one_hot_i[58];
  assign data_masked[7542] = data_i[7542] & sel_one_hot_i[58];
  assign data_masked[7541] = data_i[7541] & sel_one_hot_i[58];
  assign data_masked[7540] = data_i[7540] & sel_one_hot_i[58];
  assign data_masked[7539] = data_i[7539] & sel_one_hot_i[58];
  assign data_masked[7538] = data_i[7538] & sel_one_hot_i[58];
  assign data_masked[7537] = data_i[7537] & sel_one_hot_i[58];
  assign data_masked[7536] = data_i[7536] & sel_one_hot_i[58];
  assign data_masked[7535] = data_i[7535] & sel_one_hot_i[58];
  assign data_masked[7534] = data_i[7534] & sel_one_hot_i[58];
  assign data_masked[7533] = data_i[7533] & sel_one_hot_i[58];
  assign data_masked[7532] = data_i[7532] & sel_one_hot_i[58];
  assign data_masked[7531] = data_i[7531] & sel_one_hot_i[58];
  assign data_masked[7530] = data_i[7530] & sel_one_hot_i[58];
  assign data_masked[7529] = data_i[7529] & sel_one_hot_i[58];
  assign data_masked[7528] = data_i[7528] & sel_one_hot_i[58];
  assign data_masked[7527] = data_i[7527] & sel_one_hot_i[58];
  assign data_masked[7526] = data_i[7526] & sel_one_hot_i[58];
  assign data_masked[7525] = data_i[7525] & sel_one_hot_i[58];
  assign data_masked[7524] = data_i[7524] & sel_one_hot_i[58];
  assign data_masked[7523] = data_i[7523] & sel_one_hot_i[58];
  assign data_masked[7522] = data_i[7522] & sel_one_hot_i[58];
  assign data_masked[7521] = data_i[7521] & sel_one_hot_i[58];
  assign data_masked[7520] = data_i[7520] & sel_one_hot_i[58];
  assign data_masked[7519] = data_i[7519] & sel_one_hot_i[58];
  assign data_masked[7518] = data_i[7518] & sel_one_hot_i[58];
  assign data_masked[7517] = data_i[7517] & sel_one_hot_i[58];
  assign data_masked[7516] = data_i[7516] & sel_one_hot_i[58];
  assign data_masked[7515] = data_i[7515] & sel_one_hot_i[58];
  assign data_masked[7514] = data_i[7514] & sel_one_hot_i[58];
  assign data_masked[7513] = data_i[7513] & sel_one_hot_i[58];
  assign data_masked[7512] = data_i[7512] & sel_one_hot_i[58];
  assign data_masked[7511] = data_i[7511] & sel_one_hot_i[58];
  assign data_masked[7510] = data_i[7510] & sel_one_hot_i[58];
  assign data_masked[7509] = data_i[7509] & sel_one_hot_i[58];
  assign data_masked[7508] = data_i[7508] & sel_one_hot_i[58];
  assign data_masked[7507] = data_i[7507] & sel_one_hot_i[58];
  assign data_masked[7506] = data_i[7506] & sel_one_hot_i[58];
  assign data_masked[7505] = data_i[7505] & sel_one_hot_i[58];
  assign data_masked[7504] = data_i[7504] & sel_one_hot_i[58];
  assign data_masked[7503] = data_i[7503] & sel_one_hot_i[58];
  assign data_masked[7502] = data_i[7502] & sel_one_hot_i[58];
  assign data_masked[7501] = data_i[7501] & sel_one_hot_i[58];
  assign data_masked[7500] = data_i[7500] & sel_one_hot_i[58];
  assign data_masked[7499] = data_i[7499] & sel_one_hot_i[58];
  assign data_masked[7498] = data_i[7498] & sel_one_hot_i[58];
  assign data_masked[7497] = data_i[7497] & sel_one_hot_i[58];
  assign data_masked[7496] = data_i[7496] & sel_one_hot_i[58];
  assign data_masked[7495] = data_i[7495] & sel_one_hot_i[58];
  assign data_masked[7494] = data_i[7494] & sel_one_hot_i[58];
  assign data_masked[7493] = data_i[7493] & sel_one_hot_i[58];
  assign data_masked[7492] = data_i[7492] & sel_one_hot_i[58];
  assign data_masked[7491] = data_i[7491] & sel_one_hot_i[58];
  assign data_masked[7490] = data_i[7490] & sel_one_hot_i[58];
  assign data_masked[7489] = data_i[7489] & sel_one_hot_i[58];
  assign data_masked[7488] = data_i[7488] & sel_one_hot_i[58];
  assign data_masked[7487] = data_i[7487] & sel_one_hot_i[58];
  assign data_masked[7486] = data_i[7486] & sel_one_hot_i[58];
  assign data_masked[7485] = data_i[7485] & sel_one_hot_i[58];
  assign data_masked[7484] = data_i[7484] & sel_one_hot_i[58];
  assign data_masked[7483] = data_i[7483] & sel_one_hot_i[58];
  assign data_masked[7482] = data_i[7482] & sel_one_hot_i[58];
  assign data_masked[7481] = data_i[7481] & sel_one_hot_i[58];
  assign data_masked[7480] = data_i[7480] & sel_one_hot_i[58];
  assign data_masked[7479] = data_i[7479] & sel_one_hot_i[58];
  assign data_masked[7478] = data_i[7478] & sel_one_hot_i[58];
  assign data_masked[7477] = data_i[7477] & sel_one_hot_i[58];
  assign data_masked[7476] = data_i[7476] & sel_one_hot_i[58];
  assign data_masked[7475] = data_i[7475] & sel_one_hot_i[58];
  assign data_masked[7474] = data_i[7474] & sel_one_hot_i[58];
  assign data_masked[7473] = data_i[7473] & sel_one_hot_i[58];
  assign data_masked[7472] = data_i[7472] & sel_one_hot_i[58];
  assign data_masked[7471] = data_i[7471] & sel_one_hot_i[58];
  assign data_masked[7470] = data_i[7470] & sel_one_hot_i[58];
  assign data_masked[7469] = data_i[7469] & sel_one_hot_i[58];
  assign data_masked[7468] = data_i[7468] & sel_one_hot_i[58];
  assign data_masked[7467] = data_i[7467] & sel_one_hot_i[58];
  assign data_masked[7466] = data_i[7466] & sel_one_hot_i[58];
  assign data_masked[7465] = data_i[7465] & sel_one_hot_i[58];
  assign data_masked[7464] = data_i[7464] & sel_one_hot_i[58];
  assign data_masked[7463] = data_i[7463] & sel_one_hot_i[58];
  assign data_masked[7462] = data_i[7462] & sel_one_hot_i[58];
  assign data_masked[7461] = data_i[7461] & sel_one_hot_i[58];
  assign data_masked[7460] = data_i[7460] & sel_one_hot_i[58];
  assign data_masked[7459] = data_i[7459] & sel_one_hot_i[58];
  assign data_masked[7458] = data_i[7458] & sel_one_hot_i[58];
  assign data_masked[7457] = data_i[7457] & sel_one_hot_i[58];
  assign data_masked[7456] = data_i[7456] & sel_one_hot_i[58];
  assign data_masked[7455] = data_i[7455] & sel_one_hot_i[58];
  assign data_masked[7454] = data_i[7454] & sel_one_hot_i[58];
  assign data_masked[7453] = data_i[7453] & sel_one_hot_i[58];
  assign data_masked[7452] = data_i[7452] & sel_one_hot_i[58];
  assign data_masked[7451] = data_i[7451] & sel_one_hot_i[58];
  assign data_masked[7450] = data_i[7450] & sel_one_hot_i[58];
  assign data_masked[7449] = data_i[7449] & sel_one_hot_i[58];
  assign data_masked[7448] = data_i[7448] & sel_one_hot_i[58];
  assign data_masked[7447] = data_i[7447] & sel_one_hot_i[58];
  assign data_masked[7446] = data_i[7446] & sel_one_hot_i[58];
  assign data_masked[7445] = data_i[7445] & sel_one_hot_i[58];
  assign data_masked[7444] = data_i[7444] & sel_one_hot_i[58];
  assign data_masked[7443] = data_i[7443] & sel_one_hot_i[58];
  assign data_masked[7442] = data_i[7442] & sel_one_hot_i[58];
  assign data_masked[7441] = data_i[7441] & sel_one_hot_i[58];
  assign data_masked[7440] = data_i[7440] & sel_one_hot_i[58];
  assign data_masked[7439] = data_i[7439] & sel_one_hot_i[58];
  assign data_masked[7438] = data_i[7438] & sel_one_hot_i[58];
  assign data_masked[7437] = data_i[7437] & sel_one_hot_i[58];
  assign data_masked[7436] = data_i[7436] & sel_one_hot_i[58];
  assign data_masked[7435] = data_i[7435] & sel_one_hot_i[58];
  assign data_masked[7434] = data_i[7434] & sel_one_hot_i[58];
  assign data_masked[7433] = data_i[7433] & sel_one_hot_i[58];
  assign data_masked[7432] = data_i[7432] & sel_one_hot_i[58];
  assign data_masked[7431] = data_i[7431] & sel_one_hot_i[58];
  assign data_masked[7430] = data_i[7430] & sel_one_hot_i[58];
  assign data_masked[7429] = data_i[7429] & sel_one_hot_i[58];
  assign data_masked[7428] = data_i[7428] & sel_one_hot_i[58];
  assign data_masked[7427] = data_i[7427] & sel_one_hot_i[58];
  assign data_masked[7426] = data_i[7426] & sel_one_hot_i[58];
  assign data_masked[7425] = data_i[7425] & sel_one_hot_i[58];
  assign data_masked[7424] = data_i[7424] & sel_one_hot_i[58];
  assign data_masked[7679] = data_i[7679] & sel_one_hot_i[59];
  assign data_masked[7678] = data_i[7678] & sel_one_hot_i[59];
  assign data_masked[7677] = data_i[7677] & sel_one_hot_i[59];
  assign data_masked[7676] = data_i[7676] & sel_one_hot_i[59];
  assign data_masked[7675] = data_i[7675] & sel_one_hot_i[59];
  assign data_masked[7674] = data_i[7674] & sel_one_hot_i[59];
  assign data_masked[7673] = data_i[7673] & sel_one_hot_i[59];
  assign data_masked[7672] = data_i[7672] & sel_one_hot_i[59];
  assign data_masked[7671] = data_i[7671] & sel_one_hot_i[59];
  assign data_masked[7670] = data_i[7670] & sel_one_hot_i[59];
  assign data_masked[7669] = data_i[7669] & sel_one_hot_i[59];
  assign data_masked[7668] = data_i[7668] & sel_one_hot_i[59];
  assign data_masked[7667] = data_i[7667] & sel_one_hot_i[59];
  assign data_masked[7666] = data_i[7666] & sel_one_hot_i[59];
  assign data_masked[7665] = data_i[7665] & sel_one_hot_i[59];
  assign data_masked[7664] = data_i[7664] & sel_one_hot_i[59];
  assign data_masked[7663] = data_i[7663] & sel_one_hot_i[59];
  assign data_masked[7662] = data_i[7662] & sel_one_hot_i[59];
  assign data_masked[7661] = data_i[7661] & sel_one_hot_i[59];
  assign data_masked[7660] = data_i[7660] & sel_one_hot_i[59];
  assign data_masked[7659] = data_i[7659] & sel_one_hot_i[59];
  assign data_masked[7658] = data_i[7658] & sel_one_hot_i[59];
  assign data_masked[7657] = data_i[7657] & sel_one_hot_i[59];
  assign data_masked[7656] = data_i[7656] & sel_one_hot_i[59];
  assign data_masked[7655] = data_i[7655] & sel_one_hot_i[59];
  assign data_masked[7654] = data_i[7654] & sel_one_hot_i[59];
  assign data_masked[7653] = data_i[7653] & sel_one_hot_i[59];
  assign data_masked[7652] = data_i[7652] & sel_one_hot_i[59];
  assign data_masked[7651] = data_i[7651] & sel_one_hot_i[59];
  assign data_masked[7650] = data_i[7650] & sel_one_hot_i[59];
  assign data_masked[7649] = data_i[7649] & sel_one_hot_i[59];
  assign data_masked[7648] = data_i[7648] & sel_one_hot_i[59];
  assign data_masked[7647] = data_i[7647] & sel_one_hot_i[59];
  assign data_masked[7646] = data_i[7646] & sel_one_hot_i[59];
  assign data_masked[7645] = data_i[7645] & sel_one_hot_i[59];
  assign data_masked[7644] = data_i[7644] & sel_one_hot_i[59];
  assign data_masked[7643] = data_i[7643] & sel_one_hot_i[59];
  assign data_masked[7642] = data_i[7642] & sel_one_hot_i[59];
  assign data_masked[7641] = data_i[7641] & sel_one_hot_i[59];
  assign data_masked[7640] = data_i[7640] & sel_one_hot_i[59];
  assign data_masked[7639] = data_i[7639] & sel_one_hot_i[59];
  assign data_masked[7638] = data_i[7638] & sel_one_hot_i[59];
  assign data_masked[7637] = data_i[7637] & sel_one_hot_i[59];
  assign data_masked[7636] = data_i[7636] & sel_one_hot_i[59];
  assign data_masked[7635] = data_i[7635] & sel_one_hot_i[59];
  assign data_masked[7634] = data_i[7634] & sel_one_hot_i[59];
  assign data_masked[7633] = data_i[7633] & sel_one_hot_i[59];
  assign data_masked[7632] = data_i[7632] & sel_one_hot_i[59];
  assign data_masked[7631] = data_i[7631] & sel_one_hot_i[59];
  assign data_masked[7630] = data_i[7630] & sel_one_hot_i[59];
  assign data_masked[7629] = data_i[7629] & sel_one_hot_i[59];
  assign data_masked[7628] = data_i[7628] & sel_one_hot_i[59];
  assign data_masked[7627] = data_i[7627] & sel_one_hot_i[59];
  assign data_masked[7626] = data_i[7626] & sel_one_hot_i[59];
  assign data_masked[7625] = data_i[7625] & sel_one_hot_i[59];
  assign data_masked[7624] = data_i[7624] & sel_one_hot_i[59];
  assign data_masked[7623] = data_i[7623] & sel_one_hot_i[59];
  assign data_masked[7622] = data_i[7622] & sel_one_hot_i[59];
  assign data_masked[7621] = data_i[7621] & sel_one_hot_i[59];
  assign data_masked[7620] = data_i[7620] & sel_one_hot_i[59];
  assign data_masked[7619] = data_i[7619] & sel_one_hot_i[59];
  assign data_masked[7618] = data_i[7618] & sel_one_hot_i[59];
  assign data_masked[7617] = data_i[7617] & sel_one_hot_i[59];
  assign data_masked[7616] = data_i[7616] & sel_one_hot_i[59];
  assign data_masked[7615] = data_i[7615] & sel_one_hot_i[59];
  assign data_masked[7614] = data_i[7614] & sel_one_hot_i[59];
  assign data_masked[7613] = data_i[7613] & sel_one_hot_i[59];
  assign data_masked[7612] = data_i[7612] & sel_one_hot_i[59];
  assign data_masked[7611] = data_i[7611] & sel_one_hot_i[59];
  assign data_masked[7610] = data_i[7610] & sel_one_hot_i[59];
  assign data_masked[7609] = data_i[7609] & sel_one_hot_i[59];
  assign data_masked[7608] = data_i[7608] & sel_one_hot_i[59];
  assign data_masked[7607] = data_i[7607] & sel_one_hot_i[59];
  assign data_masked[7606] = data_i[7606] & sel_one_hot_i[59];
  assign data_masked[7605] = data_i[7605] & sel_one_hot_i[59];
  assign data_masked[7604] = data_i[7604] & sel_one_hot_i[59];
  assign data_masked[7603] = data_i[7603] & sel_one_hot_i[59];
  assign data_masked[7602] = data_i[7602] & sel_one_hot_i[59];
  assign data_masked[7601] = data_i[7601] & sel_one_hot_i[59];
  assign data_masked[7600] = data_i[7600] & sel_one_hot_i[59];
  assign data_masked[7599] = data_i[7599] & sel_one_hot_i[59];
  assign data_masked[7598] = data_i[7598] & sel_one_hot_i[59];
  assign data_masked[7597] = data_i[7597] & sel_one_hot_i[59];
  assign data_masked[7596] = data_i[7596] & sel_one_hot_i[59];
  assign data_masked[7595] = data_i[7595] & sel_one_hot_i[59];
  assign data_masked[7594] = data_i[7594] & sel_one_hot_i[59];
  assign data_masked[7593] = data_i[7593] & sel_one_hot_i[59];
  assign data_masked[7592] = data_i[7592] & sel_one_hot_i[59];
  assign data_masked[7591] = data_i[7591] & sel_one_hot_i[59];
  assign data_masked[7590] = data_i[7590] & sel_one_hot_i[59];
  assign data_masked[7589] = data_i[7589] & sel_one_hot_i[59];
  assign data_masked[7588] = data_i[7588] & sel_one_hot_i[59];
  assign data_masked[7587] = data_i[7587] & sel_one_hot_i[59];
  assign data_masked[7586] = data_i[7586] & sel_one_hot_i[59];
  assign data_masked[7585] = data_i[7585] & sel_one_hot_i[59];
  assign data_masked[7584] = data_i[7584] & sel_one_hot_i[59];
  assign data_masked[7583] = data_i[7583] & sel_one_hot_i[59];
  assign data_masked[7582] = data_i[7582] & sel_one_hot_i[59];
  assign data_masked[7581] = data_i[7581] & sel_one_hot_i[59];
  assign data_masked[7580] = data_i[7580] & sel_one_hot_i[59];
  assign data_masked[7579] = data_i[7579] & sel_one_hot_i[59];
  assign data_masked[7578] = data_i[7578] & sel_one_hot_i[59];
  assign data_masked[7577] = data_i[7577] & sel_one_hot_i[59];
  assign data_masked[7576] = data_i[7576] & sel_one_hot_i[59];
  assign data_masked[7575] = data_i[7575] & sel_one_hot_i[59];
  assign data_masked[7574] = data_i[7574] & sel_one_hot_i[59];
  assign data_masked[7573] = data_i[7573] & sel_one_hot_i[59];
  assign data_masked[7572] = data_i[7572] & sel_one_hot_i[59];
  assign data_masked[7571] = data_i[7571] & sel_one_hot_i[59];
  assign data_masked[7570] = data_i[7570] & sel_one_hot_i[59];
  assign data_masked[7569] = data_i[7569] & sel_one_hot_i[59];
  assign data_masked[7568] = data_i[7568] & sel_one_hot_i[59];
  assign data_masked[7567] = data_i[7567] & sel_one_hot_i[59];
  assign data_masked[7566] = data_i[7566] & sel_one_hot_i[59];
  assign data_masked[7565] = data_i[7565] & sel_one_hot_i[59];
  assign data_masked[7564] = data_i[7564] & sel_one_hot_i[59];
  assign data_masked[7563] = data_i[7563] & sel_one_hot_i[59];
  assign data_masked[7562] = data_i[7562] & sel_one_hot_i[59];
  assign data_masked[7561] = data_i[7561] & sel_one_hot_i[59];
  assign data_masked[7560] = data_i[7560] & sel_one_hot_i[59];
  assign data_masked[7559] = data_i[7559] & sel_one_hot_i[59];
  assign data_masked[7558] = data_i[7558] & sel_one_hot_i[59];
  assign data_masked[7557] = data_i[7557] & sel_one_hot_i[59];
  assign data_masked[7556] = data_i[7556] & sel_one_hot_i[59];
  assign data_masked[7555] = data_i[7555] & sel_one_hot_i[59];
  assign data_masked[7554] = data_i[7554] & sel_one_hot_i[59];
  assign data_masked[7553] = data_i[7553] & sel_one_hot_i[59];
  assign data_masked[7552] = data_i[7552] & sel_one_hot_i[59];
  assign data_masked[7807] = data_i[7807] & sel_one_hot_i[60];
  assign data_masked[7806] = data_i[7806] & sel_one_hot_i[60];
  assign data_masked[7805] = data_i[7805] & sel_one_hot_i[60];
  assign data_masked[7804] = data_i[7804] & sel_one_hot_i[60];
  assign data_masked[7803] = data_i[7803] & sel_one_hot_i[60];
  assign data_masked[7802] = data_i[7802] & sel_one_hot_i[60];
  assign data_masked[7801] = data_i[7801] & sel_one_hot_i[60];
  assign data_masked[7800] = data_i[7800] & sel_one_hot_i[60];
  assign data_masked[7799] = data_i[7799] & sel_one_hot_i[60];
  assign data_masked[7798] = data_i[7798] & sel_one_hot_i[60];
  assign data_masked[7797] = data_i[7797] & sel_one_hot_i[60];
  assign data_masked[7796] = data_i[7796] & sel_one_hot_i[60];
  assign data_masked[7795] = data_i[7795] & sel_one_hot_i[60];
  assign data_masked[7794] = data_i[7794] & sel_one_hot_i[60];
  assign data_masked[7793] = data_i[7793] & sel_one_hot_i[60];
  assign data_masked[7792] = data_i[7792] & sel_one_hot_i[60];
  assign data_masked[7791] = data_i[7791] & sel_one_hot_i[60];
  assign data_masked[7790] = data_i[7790] & sel_one_hot_i[60];
  assign data_masked[7789] = data_i[7789] & sel_one_hot_i[60];
  assign data_masked[7788] = data_i[7788] & sel_one_hot_i[60];
  assign data_masked[7787] = data_i[7787] & sel_one_hot_i[60];
  assign data_masked[7786] = data_i[7786] & sel_one_hot_i[60];
  assign data_masked[7785] = data_i[7785] & sel_one_hot_i[60];
  assign data_masked[7784] = data_i[7784] & sel_one_hot_i[60];
  assign data_masked[7783] = data_i[7783] & sel_one_hot_i[60];
  assign data_masked[7782] = data_i[7782] & sel_one_hot_i[60];
  assign data_masked[7781] = data_i[7781] & sel_one_hot_i[60];
  assign data_masked[7780] = data_i[7780] & sel_one_hot_i[60];
  assign data_masked[7779] = data_i[7779] & sel_one_hot_i[60];
  assign data_masked[7778] = data_i[7778] & sel_one_hot_i[60];
  assign data_masked[7777] = data_i[7777] & sel_one_hot_i[60];
  assign data_masked[7776] = data_i[7776] & sel_one_hot_i[60];
  assign data_masked[7775] = data_i[7775] & sel_one_hot_i[60];
  assign data_masked[7774] = data_i[7774] & sel_one_hot_i[60];
  assign data_masked[7773] = data_i[7773] & sel_one_hot_i[60];
  assign data_masked[7772] = data_i[7772] & sel_one_hot_i[60];
  assign data_masked[7771] = data_i[7771] & sel_one_hot_i[60];
  assign data_masked[7770] = data_i[7770] & sel_one_hot_i[60];
  assign data_masked[7769] = data_i[7769] & sel_one_hot_i[60];
  assign data_masked[7768] = data_i[7768] & sel_one_hot_i[60];
  assign data_masked[7767] = data_i[7767] & sel_one_hot_i[60];
  assign data_masked[7766] = data_i[7766] & sel_one_hot_i[60];
  assign data_masked[7765] = data_i[7765] & sel_one_hot_i[60];
  assign data_masked[7764] = data_i[7764] & sel_one_hot_i[60];
  assign data_masked[7763] = data_i[7763] & sel_one_hot_i[60];
  assign data_masked[7762] = data_i[7762] & sel_one_hot_i[60];
  assign data_masked[7761] = data_i[7761] & sel_one_hot_i[60];
  assign data_masked[7760] = data_i[7760] & sel_one_hot_i[60];
  assign data_masked[7759] = data_i[7759] & sel_one_hot_i[60];
  assign data_masked[7758] = data_i[7758] & sel_one_hot_i[60];
  assign data_masked[7757] = data_i[7757] & sel_one_hot_i[60];
  assign data_masked[7756] = data_i[7756] & sel_one_hot_i[60];
  assign data_masked[7755] = data_i[7755] & sel_one_hot_i[60];
  assign data_masked[7754] = data_i[7754] & sel_one_hot_i[60];
  assign data_masked[7753] = data_i[7753] & sel_one_hot_i[60];
  assign data_masked[7752] = data_i[7752] & sel_one_hot_i[60];
  assign data_masked[7751] = data_i[7751] & sel_one_hot_i[60];
  assign data_masked[7750] = data_i[7750] & sel_one_hot_i[60];
  assign data_masked[7749] = data_i[7749] & sel_one_hot_i[60];
  assign data_masked[7748] = data_i[7748] & sel_one_hot_i[60];
  assign data_masked[7747] = data_i[7747] & sel_one_hot_i[60];
  assign data_masked[7746] = data_i[7746] & sel_one_hot_i[60];
  assign data_masked[7745] = data_i[7745] & sel_one_hot_i[60];
  assign data_masked[7744] = data_i[7744] & sel_one_hot_i[60];
  assign data_masked[7743] = data_i[7743] & sel_one_hot_i[60];
  assign data_masked[7742] = data_i[7742] & sel_one_hot_i[60];
  assign data_masked[7741] = data_i[7741] & sel_one_hot_i[60];
  assign data_masked[7740] = data_i[7740] & sel_one_hot_i[60];
  assign data_masked[7739] = data_i[7739] & sel_one_hot_i[60];
  assign data_masked[7738] = data_i[7738] & sel_one_hot_i[60];
  assign data_masked[7737] = data_i[7737] & sel_one_hot_i[60];
  assign data_masked[7736] = data_i[7736] & sel_one_hot_i[60];
  assign data_masked[7735] = data_i[7735] & sel_one_hot_i[60];
  assign data_masked[7734] = data_i[7734] & sel_one_hot_i[60];
  assign data_masked[7733] = data_i[7733] & sel_one_hot_i[60];
  assign data_masked[7732] = data_i[7732] & sel_one_hot_i[60];
  assign data_masked[7731] = data_i[7731] & sel_one_hot_i[60];
  assign data_masked[7730] = data_i[7730] & sel_one_hot_i[60];
  assign data_masked[7729] = data_i[7729] & sel_one_hot_i[60];
  assign data_masked[7728] = data_i[7728] & sel_one_hot_i[60];
  assign data_masked[7727] = data_i[7727] & sel_one_hot_i[60];
  assign data_masked[7726] = data_i[7726] & sel_one_hot_i[60];
  assign data_masked[7725] = data_i[7725] & sel_one_hot_i[60];
  assign data_masked[7724] = data_i[7724] & sel_one_hot_i[60];
  assign data_masked[7723] = data_i[7723] & sel_one_hot_i[60];
  assign data_masked[7722] = data_i[7722] & sel_one_hot_i[60];
  assign data_masked[7721] = data_i[7721] & sel_one_hot_i[60];
  assign data_masked[7720] = data_i[7720] & sel_one_hot_i[60];
  assign data_masked[7719] = data_i[7719] & sel_one_hot_i[60];
  assign data_masked[7718] = data_i[7718] & sel_one_hot_i[60];
  assign data_masked[7717] = data_i[7717] & sel_one_hot_i[60];
  assign data_masked[7716] = data_i[7716] & sel_one_hot_i[60];
  assign data_masked[7715] = data_i[7715] & sel_one_hot_i[60];
  assign data_masked[7714] = data_i[7714] & sel_one_hot_i[60];
  assign data_masked[7713] = data_i[7713] & sel_one_hot_i[60];
  assign data_masked[7712] = data_i[7712] & sel_one_hot_i[60];
  assign data_masked[7711] = data_i[7711] & sel_one_hot_i[60];
  assign data_masked[7710] = data_i[7710] & sel_one_hot_i[60];
  assign data_masked[7709] = data_i[7709] & sel_one_hot_i[60];
  assign data_masked[7708] = data_i[7708] & sel_one_hot_i[60];
  assign data_masked[7707] = data_i[7707] & sel_one_hot_i[60];
  assign data_masked[7706] = data_i[7706] & sel_one_hot_i[60];
  assign data_masked[7705] = data_i[7705] & sel_one_hot_i[60];
  assign data_masked[7704] = data_i[7704] & sel_one_hot_i[60];
  assign data_masked[7703] = data_i[7703] & sel_one_hot_i[60];
  assign data_masked[7702] = data_i[7702] & sel_one_hot_i[60];
  assign data_masked[7701] = data_i[7701] & sel_one_hot_i[60];
  assign data_masked[7700] = data_i[7700] & sel_one_hot_i[60];
  assign data_masked[7699] = data_i[7699] & sel_one_hot_i[60];
  assign data_masked[7698] = data_i[7698] & sel_one_hot_i[60];
  assign data_masked[7697] = data_i[7697] & sel_one_hot_i[60];
  assign data_masked[7696] = data_i[7696] & sel_one_hot_i[60];
  assign data_masked[7695] = data_i[7695] & sel_one_hot_i[60];
  assign data_masked[7694] = data_i[7694] & sel_one_hot_i[60];
  assign data_masked[7693] = data_i[7693] & sel_one_hot_i[60];
  assign data_masked[7692] = data_i[7692] & sel_one_hot_i[60];
  assign data_masked[7691] = data_i[7691] & sel_one_hot_i[60];
  assign data_masked[7690] = data_i[7690] & sel_one_hot_i[60];
  assign data_masked[7689] = data_i[7689] & sel_one_hot_i[60];
  assign data_masked[7688] = data_i[7688] & sel_one_hot_i[60];
  assign data_masked[7687] = data_i[7687] & sel_one_hot_i[60];
  assign data_masked[7686] = data_i[7686] & sel_one_hot_i[60];
  assign data_masked[7685] = data_i[7685] & sel_one_hot_i[60];
  assign data_masked[7684] = data_i[7684] & sel_one_hot_i[60];
  assign data_masked[7683] = data_i[7683] & sel_one_hot_i[60];
  assign data_masked[7682] = data_i[7682] & sel_one_hot_i[60];
  assign data_masked[7681] = data_i[7681] & sel_one_hot_i[60];
  assign data_masked[7680] = data_i[7680] & sel_one_hot_i[60];
  assign data_masked[7935] = data_i[7935] & sel_one_hot_i[61];
  assign data_masked[7934] = data_i[7934] & sel_one_hot_i[61];
  assign data_masked[7933] = data_i[7933] & sel_one_hot_i[61];
  assign data_masked[7932] = data_i[7932] & sel_one_hot_i[61];
  assign data_masked[7931] = data_i[7931] & sel_one_hot_i[61];
  assign data_masked[7930] = data_i[7930] & sel_one_hot_i[61];
  assign data_masked[7929] = data_i[7929] & sel_one_hot_i[61];
  assign data_masked[7928] = data_i[7928] & sel_one_hot_i[61];
  assign data_masked[7927] = data_i[7927] & sel_one_hot_i[61];
  assign data_masked[7926] = data_i[7926] & sel_one_hot_i[61];
  assign data_masked[7925] = data_i[7925] & sel_one_hot_i[61];
  assign data_masked[7924] = data_i[7924] & sel_one_hot_i[61];
  assign data_masked[7923] = data_i[7923] & sel_one_hot_i[61];
  assign data_masked[7922] = data_i[7922] & sel_one_hot_i[61];
  assign data_masked[7921] = data_i[7921] & sel_one_hot_i[61];
  assign data_masked[7920] = data_i[7920] & sel_one_hot_i[61];
  assign data_masked[7919] = data_i[7919] & sel_one_hot_i[61];
  assign data_masked[7918] = data_i[7918] & sel_one_hot_i[61];
  assign data_masked[7917] = data_i[7917] & sel_one_hot_i[61];
  assign data_masked[7916] = data_i[7916] & sel_one_hot_i[61];
  assign data_masked[7915] = data_i[7915] & sel_one_hot_i[61];
  assign data_masked[7914] = data_i[7914] & sel_one_hot_i[61];
  assign data_masked[7913] = data_i[7913] & sel_one_hot_i[61];
  assign data_masked[7912] = data_i[7912] & sel_one_hot_i[61];
  assign data_masked[7911] = data_i[7911] & sel_one_hot_i[61];
  assign data_masked[7910] = data_i[7910] & sel_one_hot_i[61];
  assign data_masked[7909] = data_i[7909] & sel_one_hot_i[61];
  assign data_masked[7908] = data_i[7908] & sel_one_hot_i[61];
  assign data_masked[7907] = data_i[7907] & sel_one_hot_i[61];
  assign data_masked[7906] = data_i[7906] & sel_one_hot_i[61];
  assign data_masked[7905] = data_i[7905] & sel_one_hot_i[61];
  assign data_masked[7904] = data_i[7904] & sel_one_hot_i[61];
  assign data_masked[7903] = data_i[7903] & sel_one_hot_i[61];
  assign data_masked[7902] = data_i[7902] & sel_one_hot_i[61];
  assign data_masked[7901] = data_i[7901] & sel_one_hot_i[61];
  assign data_masked[7900] = data_i[7900] & sel_one_hot_i[61];
  assign data_masked[7899] = data_i[7899] & sel_one_hot_i[61];
  assign data_masked[7898] = data_i[7898] & sel_one_hot_i[61];
  assign data_masked[7897] = data_i[7897] & sel_one_hot_i[61];
  assign data_masked[7896] = data_i[7896] & sel_one_hot_i[61];
  assign data_masked[7895] = data_i[7895] & sel_one_hot_i[61];
  assign data_masked[7894] = data_i[7894] & sel_one_hot_i[61];
  assign data_masked[7893] = data_i[7893] & sel_one_hot_i[61];
  assign data_masked[7892] = data_i[7892] & sel_one_hot_i[61];
  assign data_masked[7891] = data_i[7891] & sel_one_hot_i[61];
  assign data_masked[7890] = data_i[7890] & sel_one_hot_i[61];
  assign data_masked[7889] = data_i[7889] & sel_one_hot_i[61];
  assign data_masked[7888] = data_i[7888] & sel_one_hot_i[61];
  assign data_masked[7887] = data_i[7887] & sel_one_hot_i[61];
  assign data_masked[7886] = data_i[7886] & sel_one_hot_i[61];
  assign data_masked[7885] = data_i[7885] & sel_one_hot_i[61];
  assign data_masked[7884] = data_i[7884] & sel_one_hot_i[61];
  assign data_masked[7883] = data_i[7883] & sel_one_hot_i[61];
  assign data_masked[7882] = data_i[7882] & sel_one_hot_i[61];
  assign data_masked[7881] = data_i[7881] & sel_one_hot_i[61];
  assign data_masked[7880] = data_i[7880] & sel_one_hot_i[61];
  assign data_masked[7879] = data_i[7879] & sel_one_hot_i[61];
  assign data_masked[7878] = data_i[7878] & sel_one_hot_i[61];
  assign data_masked[7877] = data_i[7877] & sel_one_hot_i[61];
  assign data_masked[7876] = data_i[7876] & sel_one_hot_i[61];
  assign data_masked[7875] = data_i[7875] & sel_one_hot_i[61];
  assign data_masked[7874] = data_i[7874] & sel_one_hot_i[61];
  assign data_masked[7873] = data_i[7873] & sel_one_hot_i[61];
  assign data_masked[7872] = data_i[7872] & sel_one_hot_i[61];
  assign data_masked[7871] = data_i[7871] & sel_one_hot_i[61];
  assign data_masked[7870] = data_i[7870] & sel_one_hot_i[61];
  assign data_masked[7869] = data_i[7869] & sel_one_hot_i[61];
  assign data_masked[7868] = data_i[7868] & sel_one_hot_i[61];
  assign data_masked[7867] = data_i[7867] & sel_one_hot_i[61];
  assign data_masked[7866] = data_i[7866] & sel_one_hot_i[61];
  assign data_masked[7865] = data_i[7865] & sel_one_hot_i[61];
  assign data_masked[7864] = data_i[7864] & sel_one_hot_i[61];
  assign data_masked[7863] = data_i[7863] & sel_one_hot_i[61];
  assign data_masked[7862] = data_i[7862] & sel_one_hot_i[61];
  assign data_masked[7861] = data_i[7861] & sel_one_hot_i[61];
  assign data_masked[7860] = data_i[7860] & sel_one_hot_i[61];
  assign data_masked[7859] = data_i[7859] & sel_one_hot_i[61];
  assign data_masked[7858] = data_i[7858] & sel_one_hot_i[61];
  assign data_masked[7857] = data_i[7857] & sel_one_hot_i[61];
  assign data_masked[7856] = data_i[7856] & sel_one_hot_i[61];
  assign data_masked[7855] = data_i[7855] & sel_one_hot_i[61];
  assign data_masked[7854] = data_i[7854] & sel_one_hot_i[61];
  assign data_masked[7853] = data_i[7853] & sel_one_hot_i[61];
  assign data_masked[7852] = data_i[7852] & sel_one_hot_i[61];
  assign data_masked[7851] = data_i[7851] & sel_one_hot_i[61];
  assign data_masked[7850] = data_i[7850] & sel_one_hot_i[61];
  assign data_masked[7849] = data_i[7849] & sel_one_hot_i[61];
  assign data_masked[7848] = data_i[7848] & sel_one_hot_i[61];
  assign data_masked[7847] = data_i[7847] & sel_one_hot_i[61];
  assign data_masked[7846] = data_i[7846] & sel_one_hot_i[61];
  assign data_masked[7845] = data_i[7845] & sel_one_hot_i[61];
  assign data_masked[7844] = data_i[7844] & sel_one_hot_i[61];
  assign data_masked[7843] = data_i[7843] & sel_one_hot_i[61];
  assign data_masked[7842] = data_i[7842] & sel_one_hot_i[61];
  assign data_masked[7841] = data_i[7841] & sel_one_hot_i[61];
  assign data_masked[7840] = data_i[7840] & sel_one_hot_i[61];
  assign data_masked[7839] = data_i[7839] & sel_one_hot_i[61];
  assign data_masked[7838] = data_i[7838] & sel_one_hot_i[61];
  assign data_masked[7837] = data_i[7837] & sel_one_hot_i[61];
  assign data_masked[7836] = data_i[7836] & sel_one_hot_i[61];
  assign data_masked[7835] = data_i[7835] & sel_one_hot_i[61];
  assign data_masked[7834] = data_i[7834] & sel_one_hot_i[61];
  assign data_masked[7833] = data_i[7833] & sel_one_hot_i[61];
  assign data_masked[7832] = data_i[7832] & sel_one_hot_i[61];
  assign data_masked[7831] = data_i[7831] & sel_one_hot_i[61];
  assign data_masked[7830] = data_i[7830] & sel_one_hot_i[61];
  assign data_masked[7829] = data_i[7829] & sel_one_hot_i[61];
  assign data_masked[7828] = data_i[7828] & sel_one_hot_i[61];
  assign data_masked[7827] = data_i[7827] & sel_one_hot_i[61];
  assign data_masked[7826] = data_i[7826] & sel_one_hot_i[61];
  assign data_masked[7825] = data_i[7825] & sel_one_hot_i[61];
  assign data_masked[7824] = data_i[7824] & sel_one_hot_i[61];
  assign data_masked[7823] = data_i[7823] & sel_one_hot_i[61];
  assign data_masked[7822] = data_i[7822] & sel_one_hot_i[61];
  assign data_masked[7821] = data_i[7821] & sel_one_hot_i[61];
  assign data_masked[7820] = data_i[7820] & sel_one_hot_i[61];
  assign data_masked[7819] = data_i[7819] & sel_one_hot_i[61];
  assign data_masked[7818] = data_i[7818] & sel_one_hot_i[61];
  assign data_masked[7817] = data_i[7817] & sel_one_hot_i[61];
  assign data_masked[7816] = data_i[7816] & sel_one_hot_i[61];
  assign data_masked[7815] = data_i[7815] & sel_one_hot_i[61];
  assign data_masked[7814] = data_i[7814] & sel_one_hot_i[61];
  assign data_masked[7813] = data_i[7813] & sel_one_hot_i[61];
  assign data_masked[7812] = data_i[7812] & sel_one_hot_i[61];
  assign data_masked[7811] = data_i[7811] & sel_one_hot_i[61];
  assign data_masked[7810] = data_i[7810] & sel_one_hot_i[61];
  assign data_masked[7809] = data_i[7809] & sel_one_hot_i[61];
  assign data_masked[7808] = data_i[7808] & sel_one_hot_i[61];
  assign data_masked[8063] = data_i[8063] & sel_one_hot_i[62];
  assign data_masked[8062] = data_i[8062] & sel_one_hot_i[62];
  assign data_masked[8061] = data_i[8061] & sel_one_hot_i[62];
  assign data_masked[8060] = data_i[8060] & sel_one_hot_i[62];
  assign data_masked[8059] = data_i[8059] & sel_one_hot_i[62];
  assign data_masked[8058] = data_i[8058] & sel_one_hot_i[62];
  assign data_masked[8057] = data_i[8057] & sel_one_hot_i[62];
  assign data_masked[8056] = data_i[8056] & sel_one_hot_i[62];
  assign data_masked[8055] = data_i[8055] & sel_one_hot_i[62];
  assign data_masked[8054] = data_i[8054] & sel_one_hot_i[62];
  assign data_masked[8053] = data_i[8053] & sel_one_hot_i[62];
  assign data_masked[8052] = data_i[8052] & sel_one_hot_i[62];
  assign data_masked[8051] = data_i[8051] & sel_one_hot_i[62];
  assign data_masked[8050] = data_i[8050] & sel_one_hot_i[62];
  assign data_masked[8049] = data_i[8049] & sel_one_hot_i[62];
  assign data_masked[8048] = data_i[8048] & sel_one_hot_i[62];
  assign data_masked[8047] = data_i[8047] & sel_one_hot_i[62];
  assign data_masked[8046] = data_i[8046] & sel_one_hot_i[62];
  assign data_masked[8045] = data_i[8045] & sel_one_hot_i[62];
  assign data_masked[8044] = data_i[8044] & sel_one_hot_i[62];
  assign data_masked[8043] = data_i[8043] & sel_one_hot_i[62];
  assign data_masked[8042] = data_i[8042] & sel_one_hot_i[62];
  assign data_masked[8041] = data_i[8041] & sel_one_hot_i[62];
  assign data_masked[8040] = data_i[8040] & sel_one_hot_i[62];
  assign data_masked[8039] = data_i[8039] & sel_one_hot_i[62];
  assign data_masked[8038] = data_i[8038] & sel_one_hot_i[62];
  assign data_masked[8037] = data_i[8037] & sel_one_hot_i[62];
  assign data_masked[8036] = data_i[8036] & sel_one_hot_i[62];
  assign data_masked[8035] = data_i[8035] & sel_one_hot_i[62];
  assign data_masked[8034] = data_i[8034] & sel_one_hot_i[62];
  assign data_masked[8033] = data_i[8033] & sel_one_hot_i[62];
  assign data_masked[8032] = data_i[8032] & sel_one_hot_i[62];
  assign data_masked[8031] = data_i[8031] & sel_one_hot_i[62];
  assign data_masked[8030] = data_i[8030] & sel_one_hot_i[62];
  assign data_masked[8029] = data_i[8029] & sel_one_hot_i[62];
  assign data_masked[8028] = data_i[8028] & sel_one_hot_i[62];
  assign data_masked[8027] = data_i[8027] & sel_one_hot_i[62];
  assign data_masked[8026] = data_i[8026] & sel_one_hot_i[62];
  assign data_masked[8025] = data_i[8025] & sel_one_hot_i[62];
  assign data_masked[8024] = data_i[8024] & sel_one_hot_i[62];
  assign data_masked[8023] = data_i[8023] & sel_one_hot_i[62];
  assign data_masked[8022] = data_i[8022] & sel_one_hot_i[62];
  assign data_masked[8021] = data_i[8021] & sel_one_hot_i[62];
  assign data_masked[8020] = data_i[8020] & sel_one_hot_i[62];
  assign data_masked[8019] = data_i[8019] & sel_one_hot_i[62];
  assign data_masked[8018] = data_i[8018] & sel_one_hot_i[62];
  assign data_masked[8017] = data_i[8017] & sel_one_hot_i[62];
  assign data_masked[8016] = data_i[8016] & sel_one_hot_i[62];
  assign data_masked[8015] = data_i[8015] & sel_one_hot_i[62];
  assign data_masked[8014] = data_i[8014] & sel_one_hot_i[62];
  assign data_masked[8013] = data_i[8013] & sel_one_hot_i[62];
  assign data_masked[8012] = data_i[8012] & sel_one_hot_i[62];
  assign data_masked[8011] = data_i[8011] & sel_one_hot_i[62];
  assign data_masked[8010] = data_i[8010] & sel_one_hot_i[62];
  assign data_masked[8009] = data_i[8009] & sel_one_hot_i[62];
  assign data_masked[8008] = data_i[8008] & sel_one_hot_i[62];
  assign data_masked[8007] = data_i[8007] & sel_one_hot_i[62];
  assign data_masked[8006] = data_i[8006] & sel_one_hot_i[62];
  assign data_masked[8005] = data_i[8005] & sel_one_hot_i[62];
  assign data_masked[8004] = data_i[8004] & sel_one_hot_i[62];
  assign data_masked[8003] = data_i[8003] & sel_one_hot_i[62];
  assign data_masked[8002] = data_i[8002] & sel_one_hot_i[62];
  assign data_masked[8001] = data_i[8001] & sel_one_hot_i[62];
  assign data_masked[8000] = data_i[8000] & sel_one_hot_i[62];
  assign data_masked[7999] = data_i[7999] & sel_one_hot_i[62];
  assign data_masked[7998] = data_i[7998] & sel_one_hot_i[62];
  assign data_masked[7997] = data_i[7997] & sel_one_hot_i[62];
  assign data_masked[7996] = data_i[7996] & sel_one_hot_i[62];
  assign data_masked[7995] = data_i[7995] & sel_one_hot_i[62];
  assign data_masked[7994] = data_i[7994] & sel_one_hot_i[62];
  assign data_masked[7993] = data_i[7993] & sel_one_hot_i[62];
  assign data_masked[7992] = data_i[7992] & sel_one_hot_i[62];
  assign data_masked[7991] = data_i[7991] & sel_one_hot_i[62];
  assign data_masked[7990] = data_i[7990] & sel_one_hot_i[62];
  assign data_masked[7989] = data_i[7989] & sel_one_hot_i[62];
  assign data_masked[7988] = data_i[7988] & sel_one_hot_i[62];
  assign data_masked[7987] = data_i[7987] & sel_one_hot_i[62];
  assign data_masked[7986] = data_i[7986] & sel_one_hot_i[62];
  assign data_masked[7985] = data_i[7985] & sel_one_hot_i[62];
  assign data_masked[7984] = data_i[7984] & sel_one_hot_i[62];
  assign data_masked[7983] = data_i[7983] & sel_one_hot_i[62];
  assign data_masked[7982] = data_i[7982] & sel_one_hot_i[62];
  assign data_masked[7981] = data_i[7981] & sel_one_hot_i[62];
  assign data_masked[7980] = data_i[7980] & sel_one_hot_i[62];
  assign data_masked[7979] = data_i[7979] & sel_one_hot_i[62];
  assign data_masked[7978] = data_i[7978] & sel_one_hot_i[62];
  assign data_masked[7977] = data_i[7977] & sel_one_hot_i[62];
  assign data_masked[7976] = data_i[7976] & sel_one_hot_i[62];
  assign data_masked[7975] = data_i[7975] & sel_one_hot_i[62];
  assign data_masked[7974] = data_i[7974] & sel_one_hot_i[62];
  assign data_masked[7973] = data_i[7973] & sel_one_hot_i[62];
  assign data_masked[7972] = data_i[7972] & sel_one_hot_i[62];
  assign data_masked[7971] = data_i[7971] & sel_one_hot_i[62];
  assign data_masked[7970] = data_i[7970] & sel_one_hot_i[62];
  assign data_masked[7969] = data_i[7969] & sel_one_hot_i[62];
  assign data_masked[7968] = data_i[7968] & sel_one_hot_i[62];
  assign data_masked[7967] = data_i[7967] & sel_one_hot_i[62];
  assign data_masked[7966] = data_i[7966] & sel_one_hot_i[62];
  assign data_masked[7965] = data_i[7965] & sel_one_hot_i[62];
  assign data_masked[7964] = data_i[7964] & sel_one_hot_i[62];
  assign data_masked[7963] = data_i[7963] & sel_one_hot_i[62];
  assign data_masked[7962] = data_i[7962] & sel_one_hot_i[62];
  assign data_masked[7961] = data_i[7961] & sel_one_hot_i[62];
  assign data_masked[7960] = data_i[7960] & sel_one_hot_i[62];
  assign data_masked[7959] = data_i[7959] & sel_one_hot_i[62];
  assign data_masked[7958] = data_i[7958] & sel_one_hot_i[62];
  assign data_masked[7957] = data_i[7957] & sel_one_hot_i[62];
  assign data_masked[7956] = data_i[7956] & sel_one_hot_i[62];
  assign data_masked[7955] = data_i[7955] & sel_one_hot_i[62];
  assign data_masked[7954] = data_i[7954] & sel_one_hot_i[62];
  assign data_masked[7953] = data_i[7953] & sel_one_hot_i[62];
  assign data_masked[7952] = data_i[7952] & sel_one_hot_i[62];
  assign data_masked[7951] = data_i[7951] & sel_one_hot_i[62];
  assign data_masked[7950] = data_i[7950] & sel_one_hot_i[62];
  assign data_masked[7949] = data_i[7949] & sel_one_hot_i[62];
  assign data_masked[7948] = data_i[7948] & sel_one_hot_i[62];
  assign data_masked[7947] = data_i[7947] & sel_one_hot_i[62];
  assign data_masked[7946] = data_i[7946] & sel_one_hot_i[62];
  assign data_masked[7945] = data_i[7945] & sel_one_hot_i[62];
  assign data_masked[7944] = data_i[7944] & sel_one_hot_i[62];
  assign data_masked[7943] = data_i[7943] & sel_one_hot_i[62];
  assign data_masked[7942] = data_i[7942] & sel_one_hot_i[62];
  assign data_masked[7941] = data_i[7941] & sel_one_hot_i[62];
  assign data_masked[7940] = data_i[7940] & sel_one_hot_i[62];
  assign data_masked[7939] = data_i[7939] & sel_one_hot_i[62];
  assign data_masked[7938] = data_i[7938] & sel_one_hot_i[62];
  assign data_masked[7937] = data_i[7937] & sel_one_hot_i[62];
  assign data_masked[7936] = data_i[7936] & sel_one_hot_i[62];
  assign data_masked[8191] = data_i[8191] & sel_one_hot_i[63];
  assign data_masked[8190] = data_i[8190] & sel_one_hot_i[63];
  assign data_masked[8189] = data_i[8189] & sel_one_hot_i[63];
  assign data_masked[8188] = data_i[8188] & sel_one_hot_i[63];
  assign data_masked[8187] = data_i[8187] & sel_one_hot_i[63];
  assign data_masked[8186] = data_i[8186] & sel_one_hot_i[63];
  assign data_masked[8185] = data_i[8185] & sel_one_hot_i[63];
  assign data_masked[8184] = data_i[8184] & sel_one_hot_i[63];
  assign data_masked[8183] = data_i[8183] & sel_one_hot_i[63];
  assign data_masked[8182] = data_i[8182] & sel_one_hot_i[63];
  assign data_masked[8181] = data_i[8181] & sel_one_hot_i[63];
  assign data_masked[8180] = data_i[8180] & sel_one_hot_i[63];
  assign data_masked[8179] = data_i[8179] & sel_one_hot_i[63];
  assign data_masked[8178] = data_i[8178] & sel_one_hot_i[63];
  assign data_masked[8177] = data_i[8177] & sel_one_hot_i[63];
  assign data_masked[8176] = data_i[8176] & sel_one_hot_i[63];
  assign data_masked[8175] = data_i[8175] & sel_one_hot_i[63];
  assign data_masked[8174] = data_i[8174] & sel_one_hot_i[63];
  assign data_masked[8173] = data_i[8173] & sel_one_hot_i[63];
  assign data_masked[8172] = data_i[8172] & sel_one_hot_i[63];
  assign data_masked[8171] = data_i[8171] & sel_one_hot_i[63];
  assign data_masked[8170] = data_i[8170] & sel_one_hot_i[63];
  assign data_masked[8169] = data_i[8169] & sel_one_hot_i[63];
  assign data_masked[8168] = data_i[8168] & sel_one_hot_i[63];
  assign data_masked[8167] = data_i[8167] & sel_one_hot_i[63];
  assign data_masked[8166] = data_i[8166] & sel_one_hot_i[63];
  assign data_masked[8165] = data_i[8165] & sel_one_hot_i[63];
  assign data_masked[8164] = data_i[8164] & sel_one_hot_i[63];
  assign data_masked[8163] = data_i[8163] & sel_one_hot_i[63];
  assign data_masked[8162] = data_i[8162] & sel_one_hot_i[63];
  assign data_masked[8161] = data_i[8161] & sel_one_hot_i[63];
  assign data_masked[8160] = data_i[8160] & sel_one_hot_i[63];
  assign data_masked[8159] = data_i[8159] & sel_one_hot_i[63];
  assign data_masked[8158] = data_i[8158] & sel_one_hot_i[63];
  assign data_masked[8157] = data_i[8157] & sel_one_hot_i[63];
  assign data_masked[8156] = data_i[8156] & sel_one_hot_i[63];
  assign data_masked[8155] = data_i[8155] & sel_one_hot_i[63];
  assign data_masked[8154] = data_i[8154] & sel_one_hot_i[63];
  assign data_masked[8153] = data_i[8153] & sel_one_hot_i[63];
  assign data_masked[8152] = data_i[8152] & sel_one_hot_i[63];
  assign data_masked[8151] = data_i[8151] & sel_one_hot_i[63];
  assign data_masked[8150] = data_i[8150] & sel_one_hot_i[63];
  assign data_masked[8149] = data_i[8149] & sel_one_hot_i[63];
  assign data_masked[8148] = data_i[8148] & sel_one_hot_i[63];
  assign data_masked[8147] = data_i[8147] & sel_one_hot_i[63];
  assign data_masked[8146] = data_i[8146] & sel_one_hot_i[63];
  assign data_masked[8145] = data_i[8145] & sel_one_hot_i[63];
  assign data_masked[8144] = data_i[8144] & sel_one_hot_i[63];
  assign data_masked[8143] = data_i[8143] & sel_one_hot_i[63];
  assign data_masked[8142] = data_i[8142] & sel_one_hot_i[63];
  assign data_masked[8141] = data_i[8141] & sel_one_hot_i[63];
  assign data_masked[8140] = data_i[8140] & sel_one_hot_i[63];
  assign data_masked[8139] = data_i[8139] & sel_one_hot_i[63];
  assign data_masked[8138] = data_i[8138] & sel_one_hot_i[63];
  assign data_masked[8137] = data_i[8137] & sel_one_hot_i[63];
  assign data_masked[8136] = data_i[8136] & sel_one_hot_i[63];
  assign data_masked[8135] = data_i[8135] & sel_one_hot_i[63];
  assign data_masked[8134] = data_i[8134] & sel_one_hot_i[63];
  assign data_masked[8133] = data_i[8133] & sel_one_hot_i[63];
  assign data_masked[8132] = data_i[8132] & sel_one_hot_i[63];
  assign data_masked[8131] = data_i[8131] & sel_one_hot_i[63];
  assign data_masked[8130] = data_i[8130] & sel_one_hot_i[63];
  assign data_masked[8129] = data_i[8129] & sel_one_hot_i[63];
  assign data_masked[8128] = data_i[8128] & sel_one_hot_i[63];
  assign data_masked[8127] = data_i[8127] & sel_one_hot_i[63];
  assign data_masked[8126] = data_i[8126] & sel_one_hot_i[63];
  assign data_masked[8125] = data_i[8125] & sel_one_hot_i[63];
  assign data_masked[8124] = data_i[8124] & sel_one_hot_i[63];
  assign data_masked[8123] = data_i[8123] & sel_one_hot_i[63];
  assign data_masked[8122] = data_i[8122] & sel_one_hot_i[63];
  assign data_masked[8121] = data_i[8121] & sel_one_hot_i[63];
  assign data_masked[8120] = data_i[8120] & sel_one_hot_i[63];
  assign data_masked[8119] = data_i[8119] & sel_one_hot_i[63];
  assign data_masked[8118] = data_i[8118] & sel_one_hot_i[63];
  assign data_masked[8117] = data_i[8117] & sel_one_hot_i[63];
  assign data_masked[8116] = data_i[8116] & sel_one_hot_i[63];
  assign data_masked[8115] = data_i[8115] & sel_one_hot_i[63];
  assign data_masked[8114] = data_i[8114] & sel_one_hot_i[63];
  assign data_masked[8113] = data_i[8113] & sel_one_hot_i[63];
  assign data_masked[8112] = data_i[8112] & sel_one_hot_i[63];
  assign data_masked[8111] = data_i[8111] & sel_one_hot_i[63];
  assign data_masked[8110] = data_i[8110] & sel_one_hot_i[63];
  assign data_masked[8109] = data_i[8109] & sel_one_hot_i[63];
  assign data_masked[8108] = data_i[8108] & sel_one_hot_i[63];
  assign data_masked[8107] = data_i[8107] & sel_one_hot_i[63];
  assign data_masked[8106] = data_i[8106] & sel_one_hot_i[63];
  assign data_masked[8105] = data_i[8105] & sel_one_hot_i[63];
  assign data_masked[8104] = data_i[8104] & sel_one_hot_i[63];
  assign data_masked[8103] = data_i[8103] & sel_one_hot_i[63];
  assign data_masked[8102] = data_i[8102] & sel_one_hot_i[63];
  assign data_masked[8101] = data_i[8101] & sel_one_hot_i[63];
  assign data_masked[8100] = data_i[8100] & sel_one_hot_i[63];
  assign data_masked[8099] = data_i[8099] & sel_one_hot_i[63];
  assign data_masked[8098] = data_i[8098] & sel_one_hot_i[63];
  assign data_masked[8097] = data_i[8097] & sel_one_hot_i[63];
  assign data_masked[8096] = data_i[8096] & sel_one_hot_i[63];
  assign data_masked[8095] = data_i[8095] & sel_one_hot_i[63];
  assign data_masked[8094] = data_i[8094] & sel_one_hot_i[63];
  assign data_masked[8093] = data_i[8093] & sel_one_hot_i[63];
  assign data_masked[8092] = data_i[8092] & sel_one_hot_i[63];
  assign data_masked[8091] = data_i[8091] & sel_one_hot_i[63];
  assign data_masked[8090] = data_i[8090] & sel_one_hot_i[63];
  assign data_masked[8089] = data_i[8089] & sel_one_hot_i[63];
  assign data_masked[8088] = data_i[8088] & sel_one_hot_i[63];
  assign data_masked[8087] = data_i[8087] & sel_one_hot_i[63];
  assign data_masked[8086] = data_i[8086] & sel_one_hot_i[63];
  assign data_masked[8085] = data_i[8085] & sel_one_hot_i[63];
  assign data_masked[8084] = data_i[8084] & sel_one_hot_i[63];
  assign data_masked[8083] = data_i[8083] & sel_one_hot_i[63];
  assign data_masked[8082] = data_i[8082] & sel_one_hot_i[63];
  assign data_masked[8081] = data_i[8081] & sel_one_hot_i[63];
  assign data_masked[8080] = data_i[8080] & sel_one_hot_i[63];
  assign data_masked[8079] = data_i[8079] & sel_one_hot_i[63];
  assign data_masked[8078] = data_i[8078] & sel_one_hot_i[63];
  assign data_masked[8077] = data_i[8077] & sel_one_hot_i[63];
  assign data_masked[8076] = data_i[8076] & sel_one_hot_i[63];
  assign data_masked[8075] = data_i[8075] & sel_one_hot_i[63];
  assign data_masked[8074] = data_i[8074] & sel_one_hot_i[63];
  assign data_masked[8073] = data_i[8073] & sel_one_hot_i[63];
  assign data_masked[8072] = data_i[8072] & sel_one_hot_i[63];
  assign data_masked[8071] = data_i[8071] & sel_one_hot_i[63];
  assign data_masked[8070] = data_i[8070] & sel_one_hot_i[63];
  assign data_masked[8069] = data_i[8069] & sel_one_hot_i[63];
  assign data_masked[8068] = data_i[8068] & sel_one_hot_i[63];
  assign data_masked[8067] = data_i[8067] & sel_one_hot_i[63];
  assign data_masked[8066] = data_i[8066] & sel_one_hot_i[63];
  assign data_masked[8065] = data_i[8065] & sel_one_hot_i[63];
  assign data_masked[8064] = data_i[8064] & sel_one_hot_i[63];
  assign data_o[0] = N61 | data_masked[0];
  assign N61 = N60 | data_masked[128];
  assign N60 = N59 | data_masked[256];
  assign N59 = N58 | data_masked[384];
  assign N58 = N57 | data_masked[512];
  assign N57 = N56 | data_masked[640];
  assign N56 = N55 | data_masked[768];
  assign N55 = N54 | data_masked[896];
  assign N54 = N53 | data_masked[1024];
  assign N53 = N52 | data_masked[1152];
  assign N52 = N51 | data_masked[1280];
  assign N51 = N50 | data_masked[1408];
  assign N50 = N49 | data_masked[1536];
  assign N49 = N48 | data_masked[1664];
  assign N48 = N47 | data_masked[1792];
  assign N47 = N46 | data_masked[1920];
  assign N46 = N45 | data_masked[2048];
  assign N45 = N44 | data_masked[2176];
  assign N44 = N43 | data_masked[2304];
  assign N43 = N42 | data_masked[2432];
  assign N42 = N41 | data_masked[2560];
  assign N41 = N40 | data_masked[2688];
  assign N40 = N39 | data_masked[2816];
  assign N39 = N38 | data_masked[2944];
  assign N38 = N37 | data_masked[3072];
  assign N37 = N36 | data_masked[3200];
  assign N36 = N35 | data_masked[3328];
  assign N35 = N34 | data_masked[3456];
  assign N34 = N33 | data_masked[3584];
  assign N33 = N32 | data_masked[3712];
  assign N32 = N31 | data_masked[3840];
  assign N31 = N30 | data_masked[3968];
  assign N30 = N29 | data_masked[4096];
  assign N29 = N28 | data_masked[4224];
  assign N28 = N27 | data_masked[4352];
  assign N27 = N26 | data_masked[4480];
  assign N26 = N25 | data_masked[4608];
  assign N25 = N24 | data_masked[4736];
  assign N24 = N23 | data_masked[4864];
  assign N23 = N22 | data_masked[4992];
  assign N22 = N21 | data_masked[5120];
  assign N21 = N20 | data_masked[5248];
  assign N20 = N19 | data_masked[5376];
  assign N19 = N18 | data_masked[5504];
  assign N18 = N17 | data_masked[5632];
  assign N17 = N16 | data_masked[5760];
  assign N16 = N15 | data_masked[5888];
  assign N15 = N14 | data_masked[6016];
  assign N14 = N13 | data_masked[6144];
  assign N13 = N12 | data_masked[6272];
  assign N12 = N11 | data_masked[6400];
  assign N11 = N10 | data_masked[6528];
  assign N10 = N9 | data_masked[6656];
  assign N9 = N8 | data_masked[6784];
  assign N8 = N7 | data_masked[6912];
  assign N7 = N6 | data_masked[7040];
  assign N6 = N5 | data_masked[7168];
  assign N5 = N4 | data_masked[7296];
  assign N4 = N3 | data_masked[7424];
  assign N3 = N2 | data_masked[7552];
  assign N2 = N1 | data_masked[7680];
  assign N1 = N0 | data_masked[7808];
  assign N0 = data_masked[8064] | data_masked[7936];
  assign data_o[1] = N123 | data_masked[1];
  assign N123 = N122 | data_masked[129];
  assign N122 = N121 | data_masked[257];
  assign N121 = N120 | data_masked[385];
  assign N120 = N119 | data_masked[513];
  assign N119 = N118 | data_masked[641];
  assign N118 = N117 | data_masked[769];
  assign N117 = N116 | data_masked[897];
  assign N116 = N115 | data_masked[1025];
  assign N115 = N114 | data_masked[1153];
  assign N114 = N113 | data_masked[1281];
  assign N113 = N112 | data_masked[1409];
  assign N112 = N111 | data_masked[1537];
  assign N111 = N110 | data_masked[1665];
  assign N110 = N109 | data_masked[1793];
  assign N109 = N108 | data_masked[1921];
  assign N108 = N107 | data_masked[2049];
  assign N107 = N106 | data_masked[2177];
  assign N106 = N105 | data_masked[2305];
  assign N105 = N104 | data_masked[2433];
  assign N104 = N103 | data_masked[2561];
  assign N103 = N102 | data_masked[2689];
  assign N102 = N101 | data_masked[2817];
  assign N101 = N100 | data_masked[2945];
  assign N100 = N99 | data_masked[3073];
  assign N99 = N98 | data_masked[3201];
  assign N98 = N97 | data_masked[3329];
  assign N97 = N96 | data_masked[3457];
  assign N96 = N95 | data_masked[3585];
  assign N95 = N94 | data_masked[3713];
  assign N94 = N93 | data_masked[3841];
  assign N93 = N92 | data_masked[3969];
  assign N92 = N91 | data_masked[4097];
  assign N91 = N90 | data_masked[4225];
  assign N90 = N89 | data_masked[4353];
  assign N89 = N88 | data_masked[4481];
  assign N88 = N87 | data_masked[4609];
  assign N87 = N86 | data_masked[4737];
  assign N86 = N85 | data_masked[4865];
  assign N85 = N84 | data_masked[4993];
  assign N84 = N83 | data_masked[5121];
  assign N83 = N82 | data_masked[5249];
  assign N82 = N81 | data_masked[5377];
  assign N81 = N80 | data_masked[5505];
  assign N80 = N79 | data_masked[5633];
  assign N79 = N78 | data_masked[5761];
  assign N78 = N77 | data_masked[5889];
  assign N77 = N76 | data_masked[6017];
  assign N76 = N75 | data_masked[6145];
  assign N75 = N74 | data_masked[6273];
  assign N74 = N73 | data_masked[6401];
  assign N73 = N72 | data_masked[6529];
  assign N72 = N71 | data_masked[6657];
  assign N71 = N70 | data_masked[6785];
  assign N70 = N69 | data_masked[6913];
  assign N69 = N68 | data_masked[7041];
  assign N68 = N67 | data_masked[7169];
  assign N67 = N66 | data_masked[7297];
  assign N66 = N65 | data_masked[7425];
  assign N65 = N64 | data_masked[7553];
  assign N64 = N63 | data_masked[7681];
  assign N63 = N62 | data_masked[7809];
  assign N62 = data_masked[8065] | data_masked[7937];
  assign data_o[2] = N185 | data_masked[2];
  assign N185 = N184 | data_masked[130];
  assign N184 = N183 | data_masked[258];
  assign N183 = N182 | data_masked[386];
  assign N182 = N181 | data_masked[514];
  assign N181 = N180 | data_masked[642];
  assign N180 = N179 | data_masked[770];
  assign N179 = N178 | data_masked[898];
  assign N178 = N177 | data_masked[1026];
  assign N177 = N176 | data_masked[1154];
  assign N176 = N175 | data_masked[1282];
  assign N175 = N174 | data_masked[1410];
  assign N174 = N173 | data_masked[1538];
  assign N173 = N172 | data_masked[1666];
  assign N172 = N171 | data_masked[1794];
  assign N171 = N170 | data_masked[1922];
  assign N170 = N169 | data_masked[2050];
  assign N169 = N168 | data_masked[2178];
  assign N168 = N167 | data_masked[2306];
  assign N167 = N166 | data_masked[2434];
  assign N166 = N165 | data_masked[2562];
  assign N165 = N164 | data_masked[2690];
  assign N164 = N163 | data_masked[2818];
  assign N163 = N162 | data_masked[2946];
  assign N162 = N161 | data_masked[3074];
  assign N161 = N160 | data_masked[3202];
  assign N160 = N159 | data_masked[3330];
  assign N159 = N158 | data_masked[3458];
  assign N158 = N157 | data_masked[3586];
  assign N157 = N156 | data_masked[3714];
  assign N156 = N155 | data_masked[3842];
  assign N155 = N154 | data_masked[3970];
  assign N154 = N153 | data_masked[4098];
  assign N153 = N152 | data_masked[4226];
  assign N152 = N151 | data_masked[4354];
  assign N151 = N150 | data_masked[4482];
  assign N150 = N149 | data_masked[4610];
  assign N149 = N148 | data_masked[4738];
  assign N148 = N147 | data_masked[4866];
  assign N147 = N146 | data_masked[4994];
  assign N146 = N145 | data_masked[5122];
  assign N145 = N144 | data_masked[5250];
  assign N144 = N143 | data_masked[5378];
  assign N143 = N142 | data_masked[5506];
  assign N142 = N141 | data_masked[5634];
  assign N141 = N140 | data_masked[5762];
  assign N140 = N139 | data_masked[5890];
  assign N139 = N138 | data_masked[6018];
  assign N138 = N137 | data_masked[6146];
  assign N137 = N136 | data_masked[6274];
  assign N136 = N135 | data_masked[6402];
  assign N135 = N134 | data_masked[6530];
  assign N134 = N133 | data_masked[6658];
  assign N133 = N132 | data_masked[6786];
  assign N132 = N131 | data_masked[6914];
  assign N131 = N130 | data_masked[7042];
  assign N130 = N129 | data_masked[7170];
  assign N129 = N128 | data_masked[7298];
  assign N128 = N127 | data_masked[7426];
  assign N127 = N126 | data_masked[7554];
  assign N126 = N125 | data_masked[7682];
  assign N125 = N124 | data_masked[7810];
  assign N124 = data_masked[8066] | data_masked[7938];
  assign data_o[3] = N247 | data_masked[3];
  assign N247 = N246 | data_masked[131];
  assign N246 = N245 | data_masked[259];
  assign N245 = N244 | data_masked[387];
  assign N244 = N243 | data_masked[515];
  assign N243 = N242 | data_masked[643];
  assign N242 = N241 | data_masked[771];
  assign N241 = N240 | data_masked[899];
  assign N240 = N239 | data_masked[1027];
  assign N239 = N238 | data_masked[1155];
  assign N238 = N237 | data_masked[1283];
  assign N237 = N236 | data_masked[1411];
  assign N236 = N235 | data_masked[1539];
  assign N235 = N234 | data_masked[1667];
  assign N234 = N233 | data_masked[1795];
  assign N233 = N232 | data_masked[1923];
  assign N232 = N231 | data_masked[2051];
  assign N231 = N230 | data_masked[2179];
  assign N230 = N229 | data_masked[2307];
  assign N229 = N228 | data_masked[2435];
  assign N228 = N227 | data_masked[2563];
  assign N227 = N226 | data_masked[2691];
  assign N226 = N225 | data_masked[2819];
  assign N225 = N224 | data_masked[2947];
  assign N224 = N223 | data_masked[3075];
  assign N223 = N222 | data_masked[3203];
  assign N222 = N221 | data_masked[3331];
  assign N221 = N220 | data_masked[3459];
  assign N220 = N219 | data_masked[3587];
  assign N219 = N218 | data_masked[3715];
  assign N218 = N217 | data_masked[3843];
  assign N217 = N216 | data_masked[3971];
  assign N216 = N215 | data_masked[4099];
  assign N215 = N214 | data_masked[4227];
  assign N214 = N213 | data_masked[4355];
  assign N213 = N212 | data_masked[4483];
  assign N212 = N211 | data_masked[4611];
  assign N211 = N210 | data_masked[4739];
  assign N210 = N209 | data_masked[4867];
  assign N209 = N208 | data_masked[4995];
  assign N208 = N207 | data_masked[5123];
  assign N207 = N206 | data_masked[5251];
  assign N206 = N205 | data_masked[5379];
  assign N205 = N204 | data_masked[5507];
  assign N204 = N203 | data_masked[5635];
  assign N203 = N202 | data_masked[5763];
  assign N202 = N201 | data_masked[5891];
  assign N201 = N200 | data_masked[6019];
  assign N200 = N199 | data_masked[6147];
  assign N199 = N198 | data_masked[6275];
  assign N198 = N197 | data_masked[6403];
  assign N197 = N196 | data_masked[6531];
  assign N196 = N195 | data_masked[6659];
  assign N195 = N194 | data_masked[6787];
  assign N194 = N193 | data_masked[6915];
  assign N193 = N192 | data_masked[7043];
  assign N192 = N191 | data_masked[7171];
  assign N191 = N190 | data_masked[7299];
  assign N190 = N189 | data_masked[7427];
  assign N189 = N188 | data_masked[7555];
  assign N188 = N187 | data_masked[7683];
  assign N187 = N186 | data_masked[7811];
  assign N186 = data_masked[8067] | data_masked[7939];
  assign data_o[4] = N309 | data_masked[4];
  assign N309 = N308 | data_masked[132];
  assign N308 = N307 | data_masked[260];
  assign N307 = N306 | data_masked[388];
  assign N306 = N305 | data_masked[516];
  assign N305 = N304 | data_masked[644];
  assign N304 = N303 | data_masked[772];
  assign N303 = N302 | data_masked[900];
  assign N302 = N301 | data_masked[1028];
  assign N301 = N300 | data_masked[1156];
  assign N300 = N299 | data_masked[1284];
  assign N299 = N298 | data_masked[1412];
  assign N298 = N297 | data_masked[1540];
  assign N297 = N296 | data_masked[1668];
  assign N296 = N295 | data_masked[1796];
  assign N295 = N294 | data_masked[1924];
  assign N294 = N293 | data_masked[2052];
  assign N293 = N292 | data_masked[2180];
  assign N292 = N291 | data_masked[2308];
  assign N291 = N290 | data_masked[2436];
  assign N290 = N289 | data_masked[2564];
  assign N289 = N288 | data_masked[2692];
  assign N288 = N287 | data_masked[2820];
  assign N287 = N286 | data_masked[2948];
  assign N286 = N285 | data_masked[3076];
  assign N285 = N284 | data_masked[3204];
  assign N284 = N283 | data_masked[3332];
  assign N283 = N282 | data_masked[3460];
  assign N282 = N281 | data_masked[3588];
  assign N281 = N280 | data_masked[3716];
  assign N280 = N279 | data_masked[3844];
  assign N279 = N278 | data_masked[3972];
  assign N278 = N277 | data_masked[4100];
  assign N277 = N276 | data_masked[4228];
  assign N276 = N275 | data_masked[4356];
  assign N275 = N274 | data_masked[4484];
  assign N274 = N273 | data_masked[4612];
  assign N273 = N272 | data_masked[4740];
  assign N272 = N271 | data_masked[4868];
  assign N271 = N270 | data_masked[4996];
  assign N270 = N269 | data_masked[5124];
  assign N269 = N268 | data_masked[5252];
  assign N268 = N267 | data_masked[5380];
  assign N267 = N266 | data_masked[5508];
  assign N266 = N265 | data_masked[5636];
  assign N265 = N264 | data_masked[5764];
  assign N264 = N263 | data_masked[5892];
  assign N263 = N262 | data_masked[6020];
  assign N262 = N261 | data_masked[6148];
  assign N261 = N260 | data_masked[6276];
  assign N260 = N259 | data_masked[6404];
  assign N259 = N258 | data_masked[6532];
  assign N258 = N257 | data_masked[6660];
  assign N257 = N256 | data_masked[6788];
  assign N256 = N255 | data_masked[6916];
  assign N255 = N254 | data_masked[7044];
  assign N254 = N253 | data_masked[7172];
  assign N253 = N252 | data_masked[7300];
  assign N252 = N251 | data_masked[7428];
  assign N251 = N250 | data_masked[7556];
  assign N250 = N249 | data_masked[7684];
  assign N249 = N248 | data_masked[7812];
  assign N248 = data_masked[8068] | data_masked[7940];
  assign data_o[5] = N371 | data_masked[5];
  assign N371 = N370 | data_masked[133];
  assign N370 = N369 | data_masked[261];
  assign N369 = N368 | data_masked[389];
  assign N368 = N367 | data_masked[517];
  assign N367 = N366 | data_masked[645];
  assign N366 = N365 | data_masked[773];
  assign N365 = N364 | data_masked[901];
  assign N364 = N363 | data_masked[1029];
  assign N363 = N362 | data_masked[1157];
  assign N362 = N361 | data_masked[1285];
  assign N361 = N360 | data_masked[1413];
  assign N360 = N359 | data_masked[1541];
  assign N359 = N358 | data_masked[1669];
  assign N358 = N357 | data_masked[1797];
  assign N357 = N356 | data_masked[1925];
  assign N356 = N355 | data_masked[2053];
  assign N355 = N354 | data_masked[2181];
  assign N354 = N353 | data_masked[2309];
  assign N353 = N352 | data_masked[2437];
  assign N352 = N351 | data_masked[2565];
  assign N351 = N350 | data_masked[2693];
  assign N350 = N349 | data_masked[2821];
  assign N349 = N348 | data_masked[2949];
  assign N348 = N347 | data_masked[3077];
  assign N347 = N346 | data_masked[3205];
  assign N346 = N345 | data_masked[3333];
  assign N345 = N344 | data_masked[3461];
  assign N344 = N343 | data_masked[3589];
  assign N343 = N342 | data_masked[3717];
  assign N342 = N341 | data_masked[3845];
  assign N341 = N340 | data_masked[3973];
  assign N340 = N339 | data_masked[4101];
  assign N339 = N338 | data_masked[4229];
  assign N338 = N337 | data_masked[4357];
  assign N337 = N336 | data_masked[4485];
  assign N336 = N335 | data_masked[4613];
  assign N335 = N334 | data_masked[4741];
  assign N334 = N333 | data_masked[4869];
  assign N333 = N332 | data_masked[4997];
  assign N332 = N331 | data_masked[5125];
  assign N331 = N330 | data_masked[5253];
  assign N330 = N329 | data_masked[5381];
  assign N329 = N328 | data_masked[5509];
  assign N328 = N327 | data_masked[5637];
  assign N327 = N326 | data_masked[5765];
  assign N326 = N325 | data_masked[5893];
  assign N325 = N324 | data_masked[6021];
  assign N324 = N323 | data_masked[6149];
  assign N323 = N322 | data_masked[6277];
  assign N322 = N321 | data_masked[6405];
  assign N321 = N320 | data_masked[6533];
  assign N320 = N319 | data_masked[6661];
  assign N319 = N318 | data_masked[6789];
  assign N318 = N317 | data_masked[6917];
  assign N317 = N316 | data_masked[7045];
  assign N316 = N315 | data_masked[7173];
  assign N315 = N314 | data_masked[7301];
  assign N314 = N313 | data_masked[7429];
  assign N313 = N312 | data_masked[7557];
  assign N312 = N311 | data_masked[7685];
  assign N311 = N310 | data_masked[7813];
  assign N310 = data_masked[8069] | data_masked[7941];
  assign data_o[6] = N433 | data_masked[6];
  assign N433 = N432 | data_masked[134];
  assign N432 = N431 | data_masked[262];
  assign N431 = N430 | data_masked[390];
  assign N430 = N429 | data_masked[518];
  assign N429 = N428 | data_masked[646];
  assign N428 = N427 | data_masked[774];
  assign N427 = N426 | data_masked[902];
  assign N426 = N425 | data_masked[1030];
  assign N425 = N424 | data_masked[1158];
  assign N424 = N423 | data_masked[1286];
  assign N423 = N422 | data_masked[1414];
  assign N422 = N421 | data_masked[1542];
  assign N421 = N420 | data_masked[1670];
  assign N420 = N419 | data_masked[1798];
  assign N419 = N418 | data_masked[1926];
  assign N418 = N417 | data_masked[2054];
  assign N417 = N416 | data_masked[2182];
  assign N416 = N415 | data_masked[2310];
  assign N415 = N414 | data_masked[2438];
  assign N414 = N413 | data_masked[2566];
  assign N413 = N412 | data_masked[2694];
  assign N412 = N411 | data_masked[2822];
  assign N411 = N410 | data_masked[2950];
  assign N410 = N409 | data_masked[3078];
  assign N409 = N408 | data_masked[3206];
  assign N408 = N407 | data_masked[3334];
  assign N407 = N406 | data_masked[3462];
  assign N406 = N405 | data_masked[3590];
  assign N405 = N404 | data_masked[3718];
  assign N404 = N403 | data_masked[3846];
  assign N403 = N402 | data_masked[3974];
  assign N402 = N401 | data_masked[4102];
  assign N401 = N400 | data_masked[4230];
  assign N400 = N399 | data_masked[4358];
  assign N399 = N398 | data_masked[4486];
  assign N398 = N397 | data_masked[4614];
  assign N397 = N396 | data_masked[4742];
  assign N396 = N395 | data_masked[4870];
  assign N395 = N394 | data_masked[4998];
  assign N394 = N393 | data_masked[5126];
  assign N393 = N392 | data_masked[5254];
  assign N392 = N391 | data_masked[5382];
  assign N391 = N390 | data_masked[5510];
  assign N390 = N389 | data_masked[5638];
  assign N389 = N388 | data_masked[5766];
  assign N388 = N387 | data_masked[5894];
  assign N387 = N386 | data_masked[6022];
  assign N386 = N385 | data_masked[6150];
  assign N385 = N384 | data_masked[6278];
  assign N384 = N383 | data_masked[6406];
  assign N383 = N382 | data_masked[6534];
  assign N382 = N381 | data_masked[6662];
  assign N381 = N380 | data_masked[6790];
  assign N380 = N379 | data_masked[6918];
  assign N379 = N378 | data_masked[7046];
  assign N378 = N377 | data_masked[7174];
  assign N377 = N376 | data_masked[7302];
  assign N376 = N375 | data_masked[7430];
  assign N375 = N374 | data_masked[7558];
  assign N374 = N373 | data_masked[7686];
  assign N373 = N372 | data_masked[7814];
  assign N372 = data_masked[8070] | data_masked[7942];
  assign data_o[7] = N495 | data_masked[7];
  assign N495 = N494 | data_masked[135];
  assign N494 = N493 | data_masked[263];
  assign N493 = N492 | data_masked[391];
  assign N492 = N491 | data_masked[519];
  assign N491 = N490 | data_masked[647];
  assign N490 = N489 | data_masked[775];
  assign N489 = N488 | data_masked[903];
  assign N488 = N487 | data_masked[1031];
  assign N487 = N486 | data_masked[1159];
  assign N486 = N485 | data_masked[1287];
  assign N485 = N484 | data_masked[1415];
  assign N484 = N483 | data_masked[1543];
  assign N483 = N482 | data_masked[1671];
  assign N482 = N481 | data_masked[1799];
  assign N481 = N480 | data_masked[1927];
  assign N480 = N479 | data_masked[2055];
  assign N479 = N478 | data_masked[2183];
  assign N478 = N477 | data_masked[2311];
  assign N477 = N476 | data_masked[2439];
  assign N476 = N475 | data_masked[2567];
  assign N475 = N474 | data_masked[2695];
  assign N474 = N473 | data_masked[2823];
  assign N473 = N472 | data_masked[2951];
  assign N472 = N471 | data_masked[3079];
  assign N471 = N470 | data_masked[3207];
  assign N470 = N469 | data_masked[3335];
  assign N469 = N468 | data_masked[3463];
  assign N468 = N467 | data_masked[3591];
  assign N467 = N466 | data_masked[3719];
  assign N466 = N465 | data_masked[3847];
  assign N465 = N464 | data_masked[3975];
  assign N464 = N463 | data_masked[4103];
  assign N463 = N462 | data_masked[4231];
  assign N462 = N461 | data_masked[4359];
  assign N461 = N460 | data_masked[4487];
  assign N460 = N459 | data_masked[4615];
  assign N459 = N458 | data_masked[4743];
  assign N458 = N457 | data_masked[4871];
  assign N457 = N456 | data_masked[4999];
  assign N456 = N455 | data_masked[5127];
  assign N455 = N454 | data_masked[5255];
  assign N454 = N453 | data_masked[5383];
  assign N453 = N452 | data_masked[5511];
  assign N452 = N451 | data_masked[5639];
  assign N451 = N450 | data_masked[5767];
  assign N450 = N449 | data_masked[5895];
  assign N449 = N448 | data_masked[6023];
  assign N448 = N447 | data_masked[6151];
  assign N447 = N446 | data_masked[6279];
  assign N446 = N445 | data_masked[6407];
  assign N445 = N444 | data_masked[6535];
  assign N444 = N443 | data_masked[6663];
  assign N443 = N442 | data_masked[6791];
  assign N442 = N441 | data_masked[6919];
  assign N441 = N440 | data_masked[7047];
  assign N440 = N439 | data_masked[7175];
  assign N439 = N438 | data_masked[7303];
  assign N438 = N437 | data_masked[7431];
  assign N437 = N436 | data_masked[7559];
  assign N436 = N435 | data_masked[7687];
  assign N435 = N434 | data_masked[7815];
  assign N434 = data_masked[8071] | data_masked[7943];
  assign data_o[8] = N557 | data_masked[8];
  assign N557 = N556 | data_masked[136];
  assign N556 = N555 | data_masked[264];
  assign N555 = N554 | data_masked[392];
  assign N554 = N553 | data_masked[520];
  assign N553 = N552 | data_masked[648];
  assign N552 = N551 | data_masked[776];
  assign N551 = N550 | data_masked[904];
  assign N550 = N549 | data_masked[1032];
  assign N549 = N548 | data_masked[1160];
  assign N548 = N547 | data_masked[1288];
  assign N547 = N546 | data_masked[1416];
  assign N546 = N545 | data_masked[1544];
  assign N545 = N544 | data_masked[1672];
  assign N544 = N543 | data_masked[1800];
  assign N543 = N542 | data_masked[1928];
  assign N542 = N541 | data_masked[2056];
  assign N541 = N540 | data_masked[2184];
  assign N540 = N539 | data_masked[2312];
  assign N539 = N538 | data_masked[2440];
  assign N538 = N537 | data_masked[2568];
  assign N537 = N536 | data_masked[2696];
  assign N536 = N535 | data_masked[2824];
  assign N535 = N534 | data_masked[2952];
  assign N534 = N533 | data_masked[3080];
  assign N533 = N532 | data_masked[3208];
  assign N532 = N531 | data_masked[3336];
  assign N531 = N530 | data_masked[3464];
  assign N530 = N529 | data_masked[3592];
  assign N529 = N528 | data_masked[3720];
  assign N528 = N527 | data_masked[3848];
  assign N527 = N526 | data_masked[3976];
  assign N526 = N525 | data_masked[4104];
  assign N525 = N524 | data_masked[4232];
  assign N524 = N523 | data_masked[4360];
  assign N523 = N522 | data_masked[4488];
  assign N522 = N521 | data_masked[4616];
  assign N521 = N520 | data_masked[4744];
  assign N520 = N519 | data_masked[4872];
  assign N519 = N518 | data_masked[5000];
  assign N518 = N517 | data_masked[5128];
  assign N517 = N516 | data_masked[5256];
  assign N516 = N515 | data_masked[5384];
  assign N515 = N514 | data_masked[5512];
  assign N514 = N513 | data_masked[5640];
  assign N513 = N512 | data_masked[5768];
  assign N512 = N511 | data_masked[5896];
  assign N511 = N510 | data_masked[6024];
  assign N510 = N509 | data_masked[6152];
  assign N509 = N508 | data_masked[6280];
  assign N508 = N507 | data_masked[6408];
  assign N507 = N506 | data_masked[6536];
  assign N506 = N505 | data_masked[6664];
  assign N505 = N504 | data_masked[6792];
  assign N504 = N503 | data_masked[6920];
  assign N503 = N502 | data_masked[7048];
  assign N502 = N501 | data_masked[7176];
  assign N501 = N500 | data_masked[7304];
  assign N500 = N499 | data_masked[7432];
  assign N499 = N498 | data_masked[7560];
  assign N498 = N497 | data_masked[7688];
  assign N497 = N496 | data_masked[7816];
  assign N496 = data_masked[8072] | data_masked[7944];
  assign data_o[9] = N619 | data_masked[9];
  assign N619 = N618 | data_masked[137];
  assign N618 = N617 | data_masked[265];
  assign N617 = N616 | data_masked[393];
  assign N616 = N615 | data_masked[521];
  assign N615 = N614 | data_masked[649];
  assign N614 = N613 | data_masked[777];
  assign N613 = N612 | data_masked[905];
  assign N612 = N611 | data_masked[1033];
  assign N611 = N610 | data_masked[1161];
  assign N610 = N609 | data_masked[1289];
  assign N609 = N608 | data_masked[1417];
  assign N608 = N607 | data_masked[1545];
  assign N607 = N606 | data_masked[1673];
  assign N606 = N605 | data_masked[1801];
  assign N605 = N604 | data_masked[1929];
  assign N604 = N603 | data_masked[2057];
  assign N603 = N602 | data_masked[2185];
  assign N602 = N601 | data_masked[2313];
  assign N601 = N600 | data_masked[2441];
  assign N600 = N599 | data_masked[2569];
  assign N599 = N598 | data_masked[2697];
  assign N598 = N597 | data_masked[2825];
  assign N597 = N596 | data_masked[2953];
  assign N596 = N595 | data_masked[3081];
  assign N595 = N594 | data_masked[3209];
  assign N594 = N593 | data_masked[3337];
  assign N593 = N592 | data_masked[3465];
  assign N592 = N591 | data_masked[3593];
  assign N591 = N590 | data_masked[3721];
  assign N590 = N589 | data_masked[3849];
  assign N589 = N588 | data_masked[3977];
  assign N588 = N587 | data_masked[4105];
  assign N587 = N586 | data_masked[4233];
  assign N586 = N585 | data_masked[4361];
  assign N585 = N584 | data_masked[4489];
  assign N584 = N583 | data_masked[4617];
  assign N583 = N582 | data_masked[4745];
  assign N582 = N581 | data_masked[4873];
  assign N581 = N580 | data_masked[5001];
  assign N580 = N579 | data_masked[5129];
  assign N579 = N578 | data_masked[5257];
  assign N578 = N577 | data_masked[5385];
  assign N577 = N576 | data_masked[5513];
  assign N576 = N575 | data_masked[5641];
  assign N575 = N574 | data_masked[5769];
  assign N574 = N573 | data_masked[5897];
  assign N573 = N572 | data_masked[6025];
  assign N572 = N571 | data_masked[6153];
  assign N571 = N570 | data_masked[6281];
  assign N570 = N569 | data_masked[6409];
  assign N569 = N568 | data_masked[6537];
  assign N568 = N567 | data_masked[6665];
  assign N567 = N566 | data_masked[6793];
  assign N566 = N565 | data_masked[6921];
  assign N565 = N564 | data_masked[7049];
  assign N564 = N563 | data_masked[7177];
  assign N563 = N562 | data_masked[7305];
  assign N562 = N561 | data_masked[7433];
  assign N561 = N560 | data_masked[7561];
  assign N560 = N559 | data_masked[7689];
  assign N559 = N558 | data_masked[7817];
  assign N558 = data_masked[8073] | data_masked[7945];
  assign data_o[10] = N681 | data_masked[10];
  assign N681 = N680 | data_masked[138];
  assign N680 = N679 | data_masked[266];
  assign N679 = N678 | data_masked[394];
  assign N678 = N677 | data_masked[522];
  assign N677 = N676 | data_masked[650];
  assign N676 = N675 | data_masked[778];
  assign N675 = N674 | data_masked[906];
  assign N674 = N673 | data_masked[1034];
  assign N673 = N672 | data_masked[1162];
  assign N672 = N671 | data_masked[1290];
  assign N671 = N670 | data_masked[1418];
  assign N670 = N669 | data_masked[1546];
  assign N669 = N668 | data_masked[1674];
  assign N668 = N667 | data_masked[1802];
  assign N667 = N666 | data_masked[1930];
  assign N666 = N665 | data_masked[2058];
  assign N665 = N664 | data_masked[2186];
  assign N664 = N663 | data_masked[2314];
  assign N663 = N662 | data_masked[2442];
  assign N662 = N661 | data_masked[2570];
  assign N661 = N660 | data_masked[2698];
  assign N660 = N659 | data_masked[2826];
  assign N659 = N658 | data_masked[2954];
  assign N658 = N657 | data_masked[3082];
  assign N657 = N656 | data_masked[3210];
  assign N656 = N655 | data_masked[3338];
  assign N655 = N654 | data_masked[3466];
  assign N654 = N653 | data_masked[3594];
  assign N653 = N652 | data_masked[3722];
  assign N652 = N651 | data_masked[3850];
  assign N651 = N650 | data_masked[3978];
  assign N650 = N649 | data_masked[4106];
  assign N649 = N648 | data_masked[4234];
  assign N648 = N647 | data_masked[4362];
  assign N647 = N646 | data_masked[4490];
  assign N646 = N645 | data_masked[4618];
  assign N645 = N644 | data_masked[4746];
  assign N644 = N643 | data_masked[4874];
  assign N643 = N642 | data_masked[5002];
  assign N642 = N641 | data_masked[5130];
  assign N641 = N640 | data_masked[5258];
  assign N640 = N639 | data_masked[5386];
  assign N639 = N638 | data_masked[5514];
  assign N638 = N637 | data_masked[5642];
  assign N637 = N636 | data_masked[5770];
  assign N636 = N635 | data_masked[5898];
  assign N635 = N634 | data_masked[6026];
  assign N634 = N633 | data_masked[6154];
  assign N633 = N632 | data_masked[6282];
  assign N632 = N631 | data_masked[6410];
  assign N631 = N630 | data_masked[6538];
  assign N630 = N629 | data_masked[6666];
  assign N629 = N628 | data_masked[6794];
  assign N628 = N627 | data_masked[6922];
  assign N627 = N626 | data_masked[7050];
  assign N626 = N625 | data_masked[7178];
  assign N625 = N624 | data_masked[7306];
  assign N624 = N623 | data_masked[7434];
  assign N623 = N622 | data_masked[7562];
  assign N622 = N621 | data_masked[7690];
  assign N621 = N620 | data_masked[7818];
  assign N620 = data_masked[8074] | data_masked[7946];
  assign data_o[11] = N743 | data_masked[11];
  assign N743 = N742 | data_masked[139];
  assign N742 = N741 | data_masked[267];
  assign N741 = N740 | data_masked[395];
  assign N740 = N739 | data_masked[523];
  assign N739 = N738 | data_masked[651];
  assign N738 = N737 | data_masked[779];
  assign N737 = N736 | data_masked[907];
  assign N736 = N735 | data_masked[1035];
  assign N735 = N734 | data_masked[1163];
  assign N734 = N733 | data_masked[1291];
  assign N733 = N732 | data_masked[1419];
  assign N732 = N731 | data_masked[1547];
  assign N731 = N730 | data_masked[1675];
  assign N730 = N729 | data_masked[1803];
  assign N729 = N728 | data_masked[1931];
  assign N728 = N727 | data_masked[2059];
  assign N727 = N726 | data_masked[2187];
  assign N726 = N725 | data_masked[2315];
  assign N725 = N724 | data_masked[2443];
  assign N724 = N723 | data_masked[2571];
  assign N723 = N722 | data_masked[2699];
  assign N722 = N721 | data_masked[2827];
  assign N721 = N720 | data_masked[2955];
  assign N720 = N719 | data_masked[3083];
  assign N719 = N718 | data_masked[3211];
  assign N718 = N717 | data_masked[3339];
  assign N717 = N716 | data_masked[3467];
  assign N716 = N715 | data_masked[3595];
  assign N715 = N714 | data_masked[3723];
  assign N714 = N713 | data_masked[3851];
  assign N713 = N712 | data_masked[3979];
  assign N712 = N711 | data_masked[4107];
  assign N711 = N710 | data_masked[4235];
  assign N710 = N709 | data_masked[4363];
  assign N709 = N708 | data_masked[4491];
  assign N708 = N707 | data_masked[4619];
  assign N707 = N706 | data_masked[4747];
  assign N706 = N705 | data_masked[4875];
  assign N705 = N704 | data_masked[5003];
  assign N704 = N703 | data_masked[5131];
  assign N703 = N702 | data_masked[5259];
  assign N702 = N701 | data_masked[5387];
  assign N701 = N700 | data_masked[5515];
  assign N700 = N699 | data_masked[5643];
  assign N699 = N698 | data_masked[5771];
  assign N698 = N697 | data_masked[5899];
  assign N697 = N696 | data_masked[6027];
  assign N696 = N695 | data_masked[6155];
  assign N695 = N694 | data_masked[6283];
  assign N694 = N693 | data_masked[6411];
  assign N693 = N692 | data_masked[6539];
  assign N692 = N691 | data_masked[6667];
  assign N691 = N690 | data_masked[6795];
  assign N690 = N689 | data_masked[6923];
  assign N689 = N688 | data_masked[7051];
  assign N688 = N687 | data_masked[7179];
  assign N687 = N686 | data_masked[7307];
  assign N686 = N685 | data_masked[7435];
  assign N685 = N684 | data_masked[7563];
  assign N684 = N683 | data_masked[7691];
  assign N683 = N682 | data_masked[7819];
  assign N682 = data_masked[8075] | data_masked[7947];
  assign data_o[12] = N805 | data_masked[12];
  assign N805 = N804 | data_masked[140];
  assign N804 = N803 | data_masked[268];
  assign N803 = N802 | data_masked[396];
  assign N802 = N801 | data_masked[524];
  assign N801 = N800 | data_masked[652];
  assign N800 = N799 | data_masked[780];
  assign N799 = N798 | data_masked[908];
  assign N798 = N797 | data_masked[1036];
  assign N797 = N796 | data_masked[1164];
  assign N796 = N795 | data_masked[1292];
  assign N795 = N794 | data_masked[1420];
  assign N794 = N793 | data_masked[1548];
  assign N793 = N792 | data_masked[1676];
  assign N792 = N791 | data_masked[1804];
  assign N791 = N790 | data_masked[1932];
  assign N790 = N789 | data_masked[2060];
  assign N789 = N788 | data_masked[2188];
  assign N788 = N787 | data_masked[2316];
  assign N787 = N786 | data_masked[2444];
  assign N786 = N785 | data_masked[2572];
  assign N785 = N784 | data_masked[2700];
  assign N784 = N783 | data_masked[2828];
  assign N783 = N782 | data_masked[2956];
  assign N782 = N781 | data_masked[3084];
  assign N781 = N780 | data_masked[3212];
  assign N780 = N779 | data_masked[3340];
  assign N779 = N778 | data_masked[3468];
  assign N778 = N777 | data_masked[3596];
  assign N777 = N776 | data_masked[3724];
  assign N776 = N775 | data_masked[3852];
  assign N775 = N774 | data_masked[3980];
  assign N774 = N773 | data_masked[4108];
  assign N773 = N772 | data_masked[4236];
  assign N772 = N771 | data_masked[4364];
  assign N771 = N770 | data_masked[4492];
  assign N770 = N769 | data_masked[4620];
  assign N769 = N768 | data_masked[4748];
  assign N768 = N767 | data_masked[4876];
  assign N767 = N766 | data_masked[5004];
  assign N766 = N765 | data_masked[5132];
  assign N765 = N764 | data_masked[5260];
  assign N764 = N763 | data_masked[5388];
  assign N763 = N762 | data_masked[5516];
  assign N762 = N761 | data_masked[5644];
  assign N761 = N760 | data_masked[5772];
  assign N760 = N759 | data_masked[5900];
  assign N759 = N758 | data_masked[6028];
  assign N758 = N757 | data_masked[6156];
  assign N757 = N756 | data_masked[6284];
  assign N756 = N755 | data_masked[6412];
  assign N755 = N754 | data_masked[6540];
  assign N754 = N753 | data_masked[6668];
  assign N753 = N752 | data_masked[6796];
  assign N752 = N751 | data_masked[6924];
  assign N751 = N750 | data_masked[7052];
  assign N750 = N749 | data_masked[7180];
  assign N749 = N748 | data_masked[7308];
  assign N748 = N747 | data_masked[7436];
  assign N747 = N746 | data_masked[7564];
  assign N746 = N745 | data_masked[7692];
  assign N745 = N744 | data_masked[7820];
  assign N744 = data_masked[8076] | data_masked[7948];
  assign data_o[13] = N867 | data_masked[13];
  assign N867 = N866 | data_masked[141];
  assign N866 = N865 | data_masked[269];
  assign N865 = N864 | data_masked[397];
  assign N864 = N863 | data_masked[525];
  assign N863 = N862 | data_masked[653];
  assign N862 = N861 | data_masked[781];
  assign N861 = N860 | data_masked[909];
  assign N860 = N859 | data_masked[1037];
  assign N859 = N858 | data_masked[1165];
  assign N858 = N857 | data_masked[1293];
  assign N857 = N856 | data_masked[1421];
  assign N856 = N855 | data_masked[1549];
  assign N855 = N854 | data_masked[1677];
  assign N854 = N853 | data_masked[1805];
  assign N853 = N852 | data_masked[1933];
  assign N852 = N851 | data_masked[2061];
  assign N851 = N850 | data_masked[2189];
  assign N850 = N849 | data_masked[2317];
  assign N849 = N848 | data_masked[2445];
  assign N848 = N847 | data_masked[2573];
  assign N847 = N846 | data_masked[2701];
  assign N846 = N845 | data_masked[2829];
  assign N845 = N844 | data_masked[2957];
  assign N844 = N843 | data_masked[3085];
  assign N843 = N842 | data_masked[3213];
  assign N842 = N841 | data_masked[3341];
  assign N841 = N840 | data_masked[3469];
  assign N840 = N839 | data_masked[3597];
  assign N839 = N838 | data_masked[3725];
  assign N838 = N837 | data_masked[3853];
  assign N837 = N836 | data_masked[3981];
  assign N836 = N835 | data_masked[4109];
  assign N835 = N834 | data_masked[4237];
  assign N834 = N833 | data_masked[4365];
  assign N833 = N832 | data_masked[4493];
  assign N832 = N831 | data_masked[4621];
  assign N831 = N830 | data_masked[4749];
  assign N830 = N829 | data_masked[4877];
  assign N829 = N828 | data_masked[5005];
  assign N828 = N827 | data_masked[5133];
  assign N827 = N826 | data_masked[5261];
  assign N826 = N825 | data_masked[5389];
  assign N825 = N824 | data_masked[5517];
  assign N824 = N823 | data_masked[5645];
  assign N823 = N822 | data_masked[5773];
  assign N822 = N821 | data_masked[5901];
  assign N821 = N820 | data_masked[6029];
  assign N820 = N819 | data_masked[6157];
  assign N819 = N818 | data_masked[6285];
  assign N818 = N817 | data_masked[6413];
  assign N817 = N816 | data_masked[6541];
  assign N816 = N815 | data_masked[6669];
  assign N815 = N814 | data_masked[6797];
  assign N814 = N813 | data_masked[6925];
  assign N813 = N812 | data_masked[7053];
  assign N812 = N811 | data_masked[7181];
  assign N811 = N810 | data_masked[7309];
  assign N810 = N809 | data_masked[7437];
  assign N809 = N808 | data_masked[7565];
  assign N808 = N807 | data_masked[7693];
  assign N807 = N806 | data_masked[7821];
  assign N806 = data_masked[8077] | data_masked[7949];
  assign data_o[14] = N929 | data_masked[14];
  assign N929 = N928 | data_masked[142];
  assign N928 = N927 | data_masked[270];
  assign N927 = N926 | data_masked[398];
  assign N926 = N925 | data_masked[526];
  assign N925 = N924 | data_masked[654];
  assign N924 = N923 | data_masked[782];
  assign N923 = N922 | data_masked[910];
  assign N922 = N921 | data_masked[1038];
  assign N921 = N920 | data_masked[1166];
  assign N920 = N919 | data_masked[1294];
  assign N919 = N918 | data_masked[1422];
  assign N918 = N917 | data_masked[1550];
  assign N917 = N916 | data_masked[1678];
  assign N916 = N915 | data_masked[1806];
  assign N915 = N914 | data_masked[1934];
  assign N914 = N913 | data_masked[2062];
  assign N913 = N912 | data_masked[2190];
  assign N912 = N911 | data_masked[2318];
  assign N911 = N910 | data_masked[2446];
  assign N910 = N909 | data_masked[2574];
  assign N909 = N908 | data_masked[2702];
  assign N908 = N907 | data_masked[2830];
  assign N907 = N906 | data_masked[2958];
  assign N906 = N905 | data_masked[3086];
  assign N905 = N904 | data_masked[3214];
  assign N904 = N903 | data_masked[3342];
  assign N903 = N902 | data_masked[3470];
  assign N902 = N901 | data_masked[3598];
  assign N901 = N900 | data_masked[3726];
  assign N900 = N899 | data_masked[3854];
  assign N899 = N898 | data_masked[3982];
  assign N898 = N897 | data_masked[4110];
  assign N897 = N896 | data_masked[4238];
  assign N896 = N895 | data_masked[4366];
  assign N895 = N894 | data_masked[4494];
  assign N894 = N893 | data_masked[4622];
  assign N893 = N892 | data_masked[4750];
  assign N892 = N891 | data_masked[4878];
  assign N891 = N890 | data_masked[5006];
  assign N890 = N889 | data_masked[5134];
  assign N889 = N888 | data_masked[5262];
  assign N888 = N887 | data_masked[5390];
  assign N887 = N886 | data_masked[5518];
  assign N886 = N885 | data_masked[5646];
  assign N885 = N884 | data_masked[5774];
  assign N884 = N883 | data_masked[5902];
  assign N883 = N882 | data_masked[6030];
  assign N882 = N881 | data_masked[6158];
  assign N881 = N880 | data_masked[6286];
  assign N880 = N879 | data_masked[6414];
  assign N879 = N878 | data_masked[6542];
  assign N878 = N877 | data_masked[6670];
  assign N877 = N876 | data_masked[6798];
  assign N876 = N875 | data_masked[6926];
  assign N875 = N874 | data_masked[7054];
  assign N874 = N873 | data_masked[7182];
  assign N873 = N872 | data_masked[7310];
  assign N872 = N871 | data_masked[7438];
  assign N871 = N870 | data_masked[7566];
  assign N870 = N869 | data_masked[7694];
  assign N869 = N868 | data_masked[7822];
  assign N868 = data_masked[8078] | data_masked[7950];
  assign data_o[15] = N991 | data_masked[15];
  assign N991 = N990 | data_masked[143];
  assign N990 = N989 | data_masked[271];
  assign N989 = N988 | data_masked[399];
  assign N988 = N987 | data_masked[527];
  assign N987 = N986 | data_masked[655];
  assign N986 = N985 | data_masked[783];
  assign N985 = N984 | data_masked[911];
  assign N984 = N983 | data_masked[1039];
  assign N983 = N982 | data_masked[1167];
  assign N982 = N981 | data_masked[1295];
  assign N981 = N980 | data_masked[1423];
  assign N980 = N979 | data_masked[1551];
  assign N979 = N978 | data_masked[1679];
  assign N978 = N977 | data_masked[1807];
  assign N977 = N976 | data_masked[1935];
  assign N976 = N975 | data_masked[2063];
  assign N975 = N974 | data_masked[2191];
  assign N974 = N973 | data_masked[2319];
  assign N973 = N972 | data_masked[2447];
  assign N972 = N971 | data_masked[2575];
  assign N971 = N970 | data_masked[2703];
  assign N970 = N969 | data_masked[2831];
  assign N969 = N968 | data_masked[2959];
  assign N968 = N967 | data_masked[3087];
  assign N967 = N966 | data_masked[3215];
  assign N966 = N965 | data_masked[3343];
  assign N965 = N964 | data_masked[3471];
  assign N964 = N963 | data_masked[3599];
  assign N963 = N962 | data_masked[3727];
  assign N962 = N961 | data_masked[3855];
  assign N961 = N960 | data_masked[3983];
  assign N960 = N959 | data_masked[4111];
  assign N959 = N958 | data_masked[4239];
  assign N958 = N957 | data_masked[4367];
  assign N957 = N956 | data_masked[4495];
  assign N956 = N955 | data_masked[4623];
  assign N955 = N954 | data_masked[4751];
  assign N954 = N953 | data_masked[4879];
  assign N953 = N952 | data_masked[5007];
  assign N952 = N951 | data_masked[5135];
  assign N951 = N950 | data_masked[5263];
  assign N950 = N949 | data_masked[5391];
  assign N949 = N948 | data_masked[5519];
  assign N948 = N947 | data_masked[5647];
  assign N947 = N946 | data_masked[5775];
  assign N946 = N945 | data_masked[5903];
  assign N945 = N944 | data_masked[6031];
  assign N944 = N943 | data_masked[6159];
  assign N943 = N942 | data_masked[6287];
  assign N942 = N941 | data_masked[6415];
  assign N941 = N940 | data_masked[6543];
  assign N940 = N939 | data_masked[6671];
  assign N939 = N938 | data_masked[6799];
  assign N938 = N937 | data_masked[6927];
  assign N937 = N936 | data_masked[7055];
  assign N936 = N935 | data_masked[7183];
  assign N935 = N934 | data_masked[7311];
  assign N934 = N933 | data_masked[7439];
  assign N933 = N932 | data_masked[7567];
  assign N932 = N931 | data_masked[7695];
  assign N931 = N930 | data_masked[7823];
  assign N930 = data_masked[8079] | data_masked[7951];
  assign data_o[16] = N1053 | data_masked[16];
  assign N1053 = N1052 | data_masked[144];
  assign N1052 = N1051 | data_masked[272];
  assign N1051 = N1050 | data_masked[400];
  assign N1050 = N1049 | data_masked[528];
  assign N1049 = N1048 | data_masked[656];
  assign N1048 = N1047 | data_masked[784];
  assign N1047 = N1046 | data_masked[912];
  assign N1046 = N1045 | data_masked[1040];
  assign N1045 = N1044 | data_masked[1168];
  assign N1044 = N1043 | data_masked[1296];
  assign N1043 = N1042 | data_masked[1424];
  assign N1042 = N1041 | data_masked[1552];
  assign N1041 = N1040 | data_masked[1680];
  assign N1040 = N1039 | data_masked[1808];
  assign N1039 = N1038 | data_masked[1936];
  assign N1038 = N1037 | data_masked[2064];
  assign N1037 = N1036 | data_masked[2192];
  assign N1036 = N1035 | data_masked[2320];
  assign N1035 = N1034 | data_masked[2448];
  assign N1034 = N1033 | data_masked[2576];
  assign N1033 = N1032 | data_masked[2704];
  assign N1032 = N1031 | data_masked[2832];
  assign N1031 = N1030 | data_masked[2960];
  assign N1030 = N1029 | data_masked[3088];
  assign N1029 = N1028 | data_masked[3216];
  assign N1028 = N1027 | data_masked[3344];
  assign N1027 = N1026 | data_masked[3472];
  assign N1026 = N1025 | data_masked[3600];
  assign N1025 = N1024 | data_masked[3728];
  assign N1024 = N1023 | data_masked[3856];
  assign N1023 = N1022 | data_masked[3984];
  assign N1022 = N1021 | data_masked[4112];
  assign N1021 = N1020 | data_masked[4240];
  assign N1020 = N1019 | data_masked[4368];
  assign N1019 = N1018 | data_masked[4496];
  assign N1018 = N1017 | data_masked[4624];
  assign N1017 = N1016 | data_masked[4752];
  assign N1016 = N1015 | data_masked[4880];
  assign N1015 = N1014 | data_masked[5008];
  assign N1014 = N1013 | data_masked[5136];
  assign N1013 = N1012 | data_masked[5264];
  assign N1012 = N1011 | data_masked[5392];
  assign N1011 = N1010 | data_masked[5520];
  assign N1010 = N1009 | data_masked[5648];
  assign N1009 = N1008 | data_masked[5776];
  assign N1008 = N1007 | data_masked[5904];
  assign N1007 = N1006 | data_masked[6032];
  assign N1006 = N1005 | data_masked[6160];
  assign N1005 = N1004 | data_masked[6288];
  assign N1004 = N1003 | data_masked[6416];
  assign N1003 = N1002 | data_masked[6544];
  assign N1002 = N1001 | data_masked[6672];
  assign N1001 = N1000 | data_masked[6800];
  assign N1000 = N999 | data_masked[6928];
  assign N999 = N998 | data_masked[7056];
  assign N998 = N997 | data_masked[7184];
  assign N997 = N996 | data_masked[7312];
  assign N996 = N995 | data_masked[7440];
  assign N995 = N994 | data_masked[7568];
  assign N994 = N993 | data_masked[7696];
  assign N993 = N992 | data_masked[7824];
  assign N992 = data_masked[8080] | data_masked[7952];
  assign data_o[17] = N1115 | data_masked[17];
  assign N1115 = N1114 | data_masked[145];
  assign N1114 = N1113 | data_masked[273];
  assign N1113 = N1112 | data_masked[401];
  assign N1112 = N1111 | data_masked[529];
  assign N1111 = N1110 | data_masked[657];
  assign N1110 = N1109 | data_masked[785];
  assign N1109 = N1108 | data_masked[913];
  assign N1108 = N1107 | data_masked[1041];
  assign N1107 = N1106 | data_masked[1169];
  assign N1106 = N1105 | data_masked[1297];
  assign N1105 = N1104 | data_masked[1425];
  assign N1104 = N1103 | data_masked[1553];
  assign N1103 = N1102 | data_masked[1681];
  assign N1102 = N1101 | data_masked[1809];
  assign N1101 = N1100 | data_masked[1937];
  assign N1100 = N1099 | data_masked[2065];
  assign N1099 = N1098 | data_masked[2193];
  assign N1098 = N1097 | data_masked[2321];
  assign N1097 = N1096 | data_masked[2449];
  assign N1096 = N1095 | data_masked[2577];
  assign N1095 = N1094 | data_masked[2705];
  assign N1094 = N1093 | data_masked[2833];
  assign N1093 = N1092 | data_masked[2961];
  assign N1092 = N1091 | data_masked[3089];
  assign N1091 = N1090 | data_masked[3217];
  assign N1090 = N1089 | data_masked[3345];
  assign N1089 = N1088 | data_masked[3473];
  assign N1088 = N1087 | data_masked[3601];
  assign N1087 = N1086 | data_masked[3729];
  assign N1086 = N1085 | data_masked[3857];
  assign N1085 = N1084 | data_masked[3985];
  assign N1084 = N1083 | data_masked[4113];
  assign N1083 = N1082 | data_masked[4241];
  assign N1082 = N1081 | data_masked[4369];
  assign N1081 = N1080 | data_masked[4497];
  assign N1080 = N1079 | data_masked[4625];
  assign N1079 = N1078 | data_masked[4753];
  assign N1078 = N1077 | data_masked[4881];
  assign N1077 = N1076 | data_masked[5009];
  assign N1076 = N1075 | data_masked[5137];
  assign N1075 = N1074 | data_masked[5265];
  assign N1074 = N1073 | data_masked[5393];
  assign N1073 = N1072 | data_masked[5521];
  assign N1072 = N1071 | data_masked[5649];
  assign N1071 = N1070 | data_masked[5777];
  assign N1070 = N1069 | data_masked[5905];
  assign N1069 = N1068 | data_masked[6033];
  assign N1068 = N1067 | data_masked[6161];
  assign N1067 = N1066 | data_masked[6289];
  assign N1066 = N1065 | data_masked[6417];
  assign N1065 = N1064 | data_masked[6545];
  assign N1064 = N1063 | data_masked[6673];
  assign N1063 = N1062 | data_masked[6801];
  assign N1062 = N1061 | data_masked[6929];
  assign N1061 = N1060 | data_masked[7057];
  assign N1060 = N1059 | data_masked[7185];
  assign N1059 = N1058 | data_masked[7313];
  assign N1058 = N1057 | data_masked[7441];
  assign N1057 = N1056 | data_masked[7569];
  assign N1056 = N1055 | data_masked[7697];
  assign N1055 = N1054 | data_masked[7825];
  assign N1054 = data_masked[8081] | data_masked[7953];
  assign data_o[18] = N1177 | data_masked[18];
  assign N1177 = N1176 | data_masked[146];
  assign N1176 = N1175 | data_masked[274];
  assign N1175 = N1174 | data_masked[402];
  assign N1174 = N1173 | data_masked[530];
  assign N1173 = N1172 | data_masked[658];
  assign N1172 = N1171 | data_masked[786];
  assign N1171 = N1170 | data_masked[914];
  assign N1170 = N1169 | data_masked[1042];
  assign N1169 = N1168 | data_masked[1170];
  assign N1168 = N1167 | data_masked[1298];
  assign N1167 = N1166 | data_masked[1426];
  assign N1166 = N1165 | data_masked[1554];
  assign N1165 = N1164 | data_masked[1682];
  assign N1164 = N1163 | data_masked[1810];
  assign N1163 = N1162 | data_masked[1938];
  assign N1162 = N1161 | data_masked[2066];
  assign N1161 = N1160 | data_masked[2194];
  assign N1160 = N1159 | data_masked[2322];
  assign N1159 = N1158 | data_masked[2450];
  assign N1158 = N1157 | data_masked[2578];
  assign N1157 = N1156 | data_masked[2706];
  assign N1156 = N1155 | data_masked[2834];
  assign N1155 = N1154 | data_masked[2962];
  assign N1154 = N1153 | data_masked[3090];
  assign N1153 = N1152 | data_masked[3218];
  assign N1152 = N1151 | data_masked[3346];
  assign N1151 = N1150 | data_masked[3474];
  assign N1150 = N1149 | data_masked[3602];
  assign N1149 = N1148 | data_masked[3730];
  assign N1148 = N1147 | data_masked[3858];
  assign N1147 = N1146 | data_masked[3986];
  assign N1146 = N1145 | data_masked[4114];
  assign N1145 = N1144 | data_masked[4242];
  assign N1144 = N1143 | data_masked[4370];
  assign N1143 = N1142 | data_masked[4498];
  assign N1142 = N1141 | data_masked[4626];
  assign N1141 = N1140 | data_masked[4754];
  assign N1140 = N1139 | data_masked[4882];
  assign N1139 = N1138 | data_masked[5010];
  assign N1138 = N1137 | data_masked[5138];
  assign N1137 = N1136 | data_masked[5266];
  assign N1136 = N1135 | data_masked[5394];
  assign N1135 = N1134 | data_masked[5522];
  assign N1134 = N1133 | data_masked[5650];
  assign N1133 = N1132 | data_masked[5778];
  assign N1132 = N1131 | data_masked[5906];
  assign N1131 = N1130 | data_masked[6034];
  assign N1130 = N1129 | data_masked[6162];
  assign N1129 = N1128 | data_masked[6290];
  assign N1128 = N1127 | data_masked[6418];
  assign N1127 = N1126 | data_masked[6546];
  assign N1126 = N1125 | data_masked[6674];
  assign N1125 = N1124 | data_masked[6802];
  assign N1124 = N1123 | data_masked[6930];
  assign N1123 = N1122 | data_masked[7058];
  assign N1122 = N1121 | data_masked[7186];
  assign N1121 = N1120 | data_masked[7314];
  assign N1120 = N1119 | data_masked[7442];
  assign N1119 = N1118 | data_masked[7570];
  assign N1118 = N1117 | data_masked[7698];
  assign N1117 = N1116 | data_masked[7826];
  assign N1116 = data_masked[8082] | data_masked[7954];
  assign data_o[19] = N1239 | data_masked[19];
  assign N1239 = N1238 | data_masked[147];
  assign N1238 = N1237 | data_masked[275];
  assign N1237 = N1236 | data_masked[403];
  assign N1236 = N1235 | data_masked[531];
  assign N1235 = N1234 | data_masked[659];
  assign N1234 = N1233 | data_masked[787];
  assign N1233 = N1232 | data_masked[915];
  assign N1232 = N1231 | data_masked[1043];
  assign N1231 = N1230 | data_masked[1171];
  assign N1230 = N1229 | data_masked[1299];
  assign N1229 = N1228 | data_masked[1427];
  assign N1228 = N1227 | data_masked[1555];
  assign N1227 = N1226 | data_masked[1683];
  assign N1226 = N1225 | data_masked[1811];
  assign N1225 = N1224 | data_masked[1939];
  assign N1224 = N1223 | data_masked[2067];
  assign N1223 = N1222 | data_masked[2195];
  assign N1222 = N1221 | data_masked[2323];
  assign N1221 = N1220 | data_masked[2451];
  assign N1220 = N1219 | data_masked[2579];
  assign N1219 = N1218 | data_masked[2707];
  assign N1218 = N1217 | data_masked[2835];
  assign N1217 = N1216 | data_masked[2963];
  assign N1216 = N1215 | data_masked[3091];
  assign N1215 = N1214 | data_masked[3219];
  assign N1214 = N1213 | data_masked[3347];
  assign N1213 = N1212 | data_masked[3475];
  assign N1212 = N1211 | data_masked[3603];
  assign N1211 = N1210 | data_masked[3731];
  assign N1210 = N1209 | data_masked[3859];
  assign N1209 = N1208 | data_masked[3987];
  assign N1208 = N1207 | data_masked[4115];
  assign N1207 = N1206 | data_masked[4243];
  assign N1206 = N1205 | data_masked[4371];
  assign N1205 = N1204 | data_masked[4499];
  assign N1204 = N1203 | data_masked[4627];
  assign N1203 = N1202 | data_masked[4755];
  assign N1202 = N1201 | data_masked[4883];
  assign N1201 = N1200 | data_masked[5011];
  assign N1200 = N1199 | data_masked[5139];
  assign N1199 = N1198 | data_masked[5267];
  assign N1198 = N1197 | data_masked[5395];
  assign N1197 = N1196 | data_masked[5523];
  assign N1196 = N1195 | data_masked[5651];
  assign N1195 = N1194 | data_masked[5779];
  assign N1194 = N1193 | data_masked[5907];
  assign N1193 = N1192 | data_masked[6035];
  assign N1192 = N1191 | data_masked[6163];
  assign N1191 = N1190 | data_masked[6291];
  assign N1190 = N1189 | data_masked[6419];
  assign N1189 = N1188 | data_masked[6547];
  assign N1188 = N1187 | data_masked[6675];
  assign N1187 = N1186 | data_masked[6803];
  assign N1186 = N1185 | data_masked[6931];
  assign N1185 = N1184 | data_masked[7059];
  assign N1184 = N1183 | data_masked[7187];
  assign N1183 = N1182 | data_masked[7315];
  assign N1182 = N1181 | data_masked[7443];
  assign N1181 = N1180 | data_masked[7571];
  assign N1180 = N1179 | data_masked[7699];
  assign N1179 = N1178 | data_masked[7827];
  assign N1178 = data_masked[8083] | data_masked[7955];
  assign data_o[20] = N1301 | data_masked[20];
  assign N1301 = N1300 | data_masked[148];
  assign N1300 = N1299 | data_masked[276];
  assign N1299 = N1298 | data_masked[404];
  assign N1298 = N1297 | data_masked[532];
  assign N1297 = N1296 | data_masked[660];
  assign N1296 = N1295 | data_masked[788];
  assign N1295 = N1294 | data_masked[916];
  assign N1294 = N1293 | data_masked[1044];
  assign N1293 = N1292 | data_masked[1172];
  assign N1292 = N1291 | data_masked[1300];
  assign N1291 = N1290 | data_masked[1428];
  assign N1290 = N1289 | data_masked[1556];
  assign N1289 = N1288 | data_masked[1684];
  assign N1288 = N1287 | data_masked[1812];
  assign N1287 = N1286 | data_masked[1940];
  assign N1286 = N1285 | data_masked[2068];
  assign N1285 = N1284 | data_masked[2196];
  assign N1284 = N1283 | data_masked[2324];
  assign N1283 = N1282 | data_masked[2452];
  assign N1282 = N1281 | data_masked[2580];
  assign N1281 = N1280 | data_masked[2708];
  assign N1280 = N1279 | data_masked[2836];
  assign N1279 = N1278 | data_masked[2964];
  assign N1278 = N1277 | data_masked[3092];
  assign N1277 = N1276 | data_masked[3220];
  assign N1276 = N1275 | data_masked[3348];
  assign N1275 = N1274 | data_masked[3476];
  assign N1274 = N1273 | data_masked[3604];
  assign N1273 = N1272 | data_masked[3732];
  assign N1272 = N1271 | data_masked[3860];
  assign N1271 = N1270 | data_masked[3988];
  assign N1270 = N1269 | data_masked[4116];
  assign N1269 = N1268 | data_masked[4244];
  assign N1268 = N1267 | data_masked[4372];
  assign N1267 = N1266 | data_masked[4500];
  assign N1266 = N1265 | data_masked[4628];
  assign N1265 = N1264 | data_masked[4756];
  assign N1264 = N1263 | data_masked[4884];
  assign N1263 = N1262 | data_masked[5012];
  assign N1262 = N1261 | data_masked[5140];
  assign N1261 = N1260 | data_masked[5268];
  assign N1260 = N1259 | data_masked[5396];
  assign N1259 = N1258 | data_masked[5524];
  assign N1258 = N1257 | data_masked[5652];
  assign N1257 = N1256 | data_masked[5780];
  assign N1256 = N1255 | data_masked[5908];
  assign N1255 = N1254 | data_masked[6036];
  assign N1254 = N1253 | data_masked[6164];
  assign N1253 = N1252 | data_masked[6292];
  assign N1252 = N1251 | data_masked[6420];
  assign N1251 = N1250 | data_masked[6548];
  assign N1250 = N1249 | data_masked[6676];
  assign N1249 = N1248 | data_masked[6804];
  assign N1248 = N1247 | data_masked[6932];
  assign N1247 = N1246 | data_masked[7060];
  assign N1246 = N1245 | data_masked[7188];
  assign N1245 = N1244 | data_masked[7316];
  assign N1244 = N1243 | data_masked[7444];
  assign N1243 = N1242 | data_masked[7572];
  assign N1242 = N1241 | data_masked[7700];
  assign N1241 = N1240 | data_masked[7828];
  assign N1240 = data_masked[8084] | data_masked[7956];
  assign data_o[21] = N1363 | data_masked[21];
  assign N1363 = N1362 | data_masked[149];
  assign N1362 = N1361 | data_masked[277];
  assign N1361 = N1360 | data_masked[405];
  assign N1360 = N1359 | data_masked[533];
  assign N1359 = N1358 | data_masked[661];
  assign N1358 = N1357 | data_masked[789];
  assign N1357 = N1356 | data_masked[917];
  assign N1356 = N1355 | data_masked[1045];
  assign N1355 = N1354 | data_masked[1173];
  assign N1354 = N1353 | data_masked[1301];
  assign N1353 = N1352 | data_masked[1429];
  assign N1352 = N1351 | data_masked[1557];
  assign N1351 = N1350 | data_masked[1685];
  assign N1350 = N1349 | data_masked[1813];
  assign N1349 = N1348 | data_masked[1941];
  assign N1348 = N1347 | data_masked[2069];
  assign N1347 = N1346 | data_masked[2197];
  assign N1346 = N1345 | data_masked[2325];
  assign N1345 = N1344 | data_masked[2453];
  assign N1344 = N1343 | data_masked[2581];
  assign N1343 = N1342 | data_masked[2709];
  assign N1342 = N1341 | data_masked[2837];
  assign N1341 = N1340 | data_masked[2965];
  assign N1340 = N1339 | data_masked[3093];
  assign N1339 = N1338 | data_masked[3221];
  assign N1338 = N1337 | data_masked[3349];
  assign N1337 = N1336 | data_masked[3477];
  assign N1336 = N1335 | data_masked[3605];
  assign N1335 = N1334 | data_masked[3733];
  assign N1334 = N1333 | data_masked[3861];
  assign N1333 = N1332 | data_masked[3989];
  assign N1332 = N1331 | data_masked[4117];
  assign N1331 = N1330 | data_masked[4245];
  assign N1330 = N1329 | data_masked[4373];
  assign N1329 = N1328 | data_masked[4501];
  assign N1328 = N1327 | data_masked[4629];
  assign N1327 = N1326 | data_masked[4757];
  assign N1326 = N1325 | data_masked[4885];
  assign N1325 = N1324 | data_masked[5013];
  assign N1324 = N1323 | data_masked[5141];
  assign N1323 = N1322 | data_masked[5269];
  assign N1322 = N1321 | data_masked[5397];
  assign N1321 = N1320 | data_masked[5525];
  assign N1320 = N1319 | data_masked[5653];
  assign N1319 = N1318 | data_masked[5781];
  assign N1318 = N1317 | data_masked[5909];
  assign N1317 = N1316 | data_masked[6037];
  assign N1316 = N1315 | data_masked[6165];
  assign N1315 = N1314 | data_masked[6293];
  assign N1314 = N1313 | data_masked[6421];
  assign N1313 = N1312 | data_masked[6549];
  assign N1312 = N1311 | data_masked[6677];
  assign N1311 = N1310 | data_masked[6805];
  assign N1310 = N1309 | data_masked[6933];
  assign N1309 = N1308 | data_masked[7061];
  assign N1308 = N1307 | data_masked[7189];
  assign N1307 = N1306 | data_masked[7317];
  assign N1306 = N1305 | data_masked[7445];
  assign N1305 = N1304 | data_masked[7573];
  assign N1304 = N1303 | data_masked[7701];
  assign N1303 = N1302 | data_masked[7829];
  assign N1302 = data_masked[8085] | data_masked[7957];
  assign data_o[22] = N1425 | data_masked[22];
  assign N1425 = N1424 | data_masked[150];
  assign N1424 = N1423 | data_masked[278];
  assign N1423 = N1422 | data_masked[406];
  assign N1422 = N1421 | data_masked[534];
  assign N1421 = N1420 | data_masked[662];
  assign N1420 = N1419 | data_masked[790];
  assign N1419 = N1418 | data_masked[918];
  assign N1418 = N1417 | data_masked[1046];
  assign N1417 = N1416 | data_masked[1174];
  assign N1416 = N1415 | data_masked[1302];
  assign N1415 = N1414 | data_masked[1430];
  assign N1414 = N1413 | data_masked[1558];
  assign N1413 = N1412 | data_masked[1686];
  assign N1412 = N1411 | data_masked[1814];
  assign N1411 = N1410 | data_masked[1942];
  assign N1410 = N1409 | data_masked[2070];
  assign N1409 = N1408 | data_masked[2198];
  assign N1408 = N1407 | data_masked[2326];
  assign N1407 = N1406 | data_masked[2454];
  assign N1406 = N1405 | data_masked[2582];
  assign N1405 = N1404 | data_masked[2710];
  assign N1404 = N1403 | data_masked[2838];
  assign N1403 = N1402 | data_masked[2966];
  assign N1402 = N1401 | data_masked[3094];
  assign N1401 = N1400 | data_masked[3222];
  assign N1400 = N1399 | data_masked[3350];
  assign N1399 = N1398 | data_masked[3478];
  assign N1398 = N1397 | data_masked[3606];
  assign N1397 = N1396 | data_masked[3734];
  assign N1396 = N1395 | data_masked[3862];
  assign N1395 = N1394 | data_masked[3990];
  assign N1394 = N1393 | data_masked[4118];
  assign N1393 = N1392 | data_masked[4246];
  assign N1392 = N1391 | data_masked[4374];
  assign N1391 = N1390 | data_masked[4502];
  assign N1390 = N1389 | data_masked[4630];
  assign N1389 = N1388 | data_masked[4758];
  assign N1388 = N1387 | data_masked[4886];
  assign N1387 = N1386 | data_masked[5014];
  assign N1386 = N1385 | data_masked[5142];
  assign N1385 = N1384 | data_masked[5270];
  assign N1384 = N1383 | data_masked[5398];
  assign N1383 = N1382 | data_masked[5526];
  assign N1382 = N1381 | data_masked[5654];
  assign N1381 = N1380 | data_masked[5782];
  assign N1380 = N1379 | data_masked[5910];
  assign N1379 = N1378 | data_masked[6038];
  assign N1378 = N1377 | data_masked[6166];
  assign N1377 = N1376 | data_masked[6294];
  assign N1376 = N1375 | data_masked[6422];
  assign N1375 = N1374 | data_masked[6550];
  assign N1374 = N1373 | data_masked[6678];
  assign N1373 = N1372 | data_masked[6806];
  assign N1372 = N1371 | data_masked[6934];
  assign N1371 = N1370 | data_masked[7062];
  assign N1370 = N1369 | data_masked[7190];
  assign N1369 = N1368 | data_masked[7318];
  assign N1368 = N1367 | data_masked[7446];
  assign N1367 = N1366 | data_masked[7574];
  assign N1366 = N1365 | data_masked[7702];
  assign N1365 = N1364 | data_masked[7830];
  assign N1364 = data_masked[8086] | data_masked[7958];
  assign data_o[23] = N1487 | data_masked[23];
  assign N1487 = N1486 | data_masked[151];
  assign N1486 = N1485 | data_masked[279];
  assign N1485 = N1484 | data_masked[407];
  assign N1484 = N1483 | data_masked[535];
  assign N1483 = N1482 | data_masked[663];
  assign N1482 = N1481 | data_masked[791];
  assign N1481 = N1480 | data_masked[919];
  assign N1480 = N1479 | data_masked[1047];
  assign N1479 = N1478 | data_masked[1175];
  assign N1478 = N1477 | data_masked[1303];
  assign N1477 = N1476 | data_masked[1431];
  assign N1476 = N1475 | data_masked[1559];
  assign N1475 = N1474 | data_masked[1687];
  assign N1474 = N1473 | data_masked[1815];
  assign N1473 = N1472 | data_masked[1943];
  assign N1472 = N1471 | data_masked[2071];
  assign N1471 = N1470 | data_masked[2199];
  assign N1470 = N1469 | data_masked[2327];
  assign N1469 = N1468 | data_masked[2455];
  assign N1468 = N1467 | data_masked[2583];
  assign N1467 = N1466 | data_masked[2711];
  assign N1466 = N1465 | data_masked[2839];
  assign N1465 = N1464 | data_masked[2967];
  assign N1464 = N1463 | data_masked[3095];
  assign N1463 = N1462 | data_masked[3223];
  assign N1462 = N1461 | data_masked[3351];
  assign N1461 = N1460 | data_masked[3479];
  assign N1460 = N1459 | data_masked[3607];
  assign N1459 = N1458 | data_masked[3735];
  assign N1458 = N1457 | data_masked[3863];
  assign N1457 = N1456 | data_masked[3991];
  assign N1456 = N1455 | data_masked[4119];
  assign N1455 = N1454 | data_masked[4247];
  assign N1454 = N1453 | data_masked[4375];
  assign N1453 = N1452 | data_masked[4503];
  assign N1452 = N1451 | data_masked[4631];
  assign N1451 = N1450 | data_masked[4759];
  assign N1450 = N1449 | data_masked[4887];
  assign N1449 = N1448 | data_masked[5015];
  assign N1448 = N1447 | data_masked[5143];
  assign N1447 = N1446 | data_masked[5271];
  assign N1446 = N1445 | data_masked[5399];
  assign N1445 = N1444 | data_masked[5527];
  assign N1444 = N1443 | data_masked[5655];
  assign N1443 = N1442 | data_masked[5783];
  assign N1442 = N1441 | data_masked[5911];
  assign N1441 = N1440 | data_masked[6039];
  assign N1440 = N1439 | data_masked[6167];
  assign N1439 = N1438 | data_masked[6295];
  assign N1438 = N1437 | data_masked[6423];
  assign N1437 = N1436 | data_masked[6551];
  assign N1436 = N1435 | data_masked[6679];
  assign N1435 = N1434 | data_masked[6807];
  assign N1434 = N1433 | data_masked[6935];
  assign N1433 = N1432 | data_masked[7063];
  assign N1432 = N1431 | data_masked[7191];
  assign N1431 = N1430 | data_masked[7319];
  assign N1430 = N1429 | data_masked[7447];
  assign N1429 = N1428 | data_masked[7575];
  assign N1428 = N1427 | data_masked[7703];
  assign N1427 = N1426 | data_masked[7831];
  assign N1426 = data_masked[8087] | data_masked[7959];
  assign data_o[24] = N1549 | data_masked[24];
  assign N1549 = N1548 | data_masked[152];
  assign N1548 = N1547 | data_masked[280];
  assign N1547 = N1546 | data_masked[408];
  assign N1546 = N1545 | data_masked[536];
  assign N1545 = N1544 | data_masked[664];
  assign N1544 = N1543 | data_masked[792];
  assign N1543 = N1542 | data_masked[920];
  assign N1542 = N1541 | data_masked[1048];
  assign N1541 = N1540 | data_masked[1176];
  assign N1540 = N1539 | data_masked[1304];
  assign N1539 = N1538 | data_masked[1432];
  assign N1538 = N1537 | data_masked[1560];
  assign N1537 = N1536 | data_masked[1688];
  assign N1536 = N1535 | data_masked[1816];
  assign N1535 = N1534 | data_masked[1944];
  assign N1534 = N1533 | data_masked[2072];
  assign N1533 = N1532 | data_masked[2200];
  assign N1532 = N1531 | data_masked[2328];
  assign N1531 = N1530 | data_masked[2456];
  assign N1530 = N1529 | data_masked[2584];
  assign N1529 = N1528 | data_masked[2712];
  assign N1528 = N1527 | data_masked[2840];
  assign N1527 = N1526 | data_masked[2968];
  assign N1526 = N1525 | data_masked[3096];
  assign N1525 = N1524 | data_masked[3224];
  assign N1524 = N1523 | data_masked[3352];
  assign N1523 = N1522 | data_masked[3480];
  assign N1522 = N1521 | data_masked[3608];
  assign N1521 = N1520 | data_masked[3736];
  assign N1520 = N1519 | data_masked[3864];
  assign N1519 = N1518 | data_masked[3992];
  assign N1518 = N1517 | data_masked[4120];
  assign N1517 = N1516 | data_masked[4248];
  assign N1516 = N1515 | data_masked[4376];
  assign N1515 = N1514 | data_masked[4504];
  assign N1514 = N1513 | data_masked[4632];
  assign N1513 = N1512 | data_masked[4760];
  assign N1512 = N1511 | data_masked[4888];
  assign N1511 = N1510 | data_masked[5016];
  assign N1510 = N1509 | data_masked[5144];
  assign N1509 = N1508 | data_masked[5272];
  assign N1508 = N1507 | data_masked[5400];
  assign N1507 = N1506 | data_masked[5528];
  assign N1506 = N1505 | data_masked[5656];
  assign N1505 = N1504 | data_masked[5784];
  assign N1504 = N1503 | data_masked[5912];
  assign N1503 = N1502 | data_masked[6040];
  assign N1502 = N1501 | data_masked[6168];
  assign N1501 = N1500 | data_masked[6296];
  assign N1500 = N1499 | data_masked[6424];
  assign N1499 = N1498 | data_masked[6552];
  assign N1498 = N1497 | data_masked[6680];
  assign N1497 = N1496 | data_masked[6808];
  assign N1496 = N1495 | data_masked[6936];
  assign N1495 = N1494 | data_masked[7064];
  assign N1494 = N1493 | data_masked[7192];
  assign N1493 = N1492 | data_masked[7320];
  assign N1492 = N1491 | data_masked[7448];
  assign N1491 = N1490 | data_masked[7576];
  assign N1490 = N1489 | data_masked[7704];
  assign N1489 = N1488 | data_masked[7832];
  assign N1488 = data_masked[8088] | data_masked[7960];
  assign data_o[25] = N1611 | data_masked[25];
  assign N1611 = N1610 | data_masked[153];
  assign N1610 = N1609 | data_masked[281];
  assign N1609 = N1608 | data_masked[409];
  assign N1608 = N1607 | data_masked[537];
  assign N1607 = N1606 | data_masked[665];
  assign N1606 = N1605 | data_masked[793];
  assign N1605 = N1604 | data_masked[921];
  assign N1604 = N1603 | data_masked[1049];
  assign N1603 = N1602 | data_masked[1177];
  assign N1602 = N1601 | data_masked[1305];
  assign N1601 = N1600 | data_masked[1433];
  assign N1600 = N1599 | data_masked[1561];
  assign N1599 = N1598 | data_masked[1689];
  assign N1598 = N1597 | data_masked[1817];
  assign N1597 = N1596 | data_masked[1945];
  assign N1596 = N1595 | data_masked[2073];
  assign N1595 = N1594 | data_masked[2201];
  assign N1594 = N1593 | data_masked[2329];
  assign N1593 = N1592 | data_masked[2457];
  assign N1592 = N1591 | data_masked[2585];
  assign N1591 = N1590 | data_masked[2713];
  assign N1590 = N1589 | data_masked[2841];
  assign N1589 = N1588 | data_masked[2969];
  assign N1588 = N1587 | data_masked[3097];
  assign N1587 = N1586 | data_masked[3225];
  assign N1586 = N1585 | data_masked[3353];
  assign N1585 = N1584 | data_masked[3481];
  assign N1584 = N1583 | data_masked[3609];
  assign N1583 = N1582 | data_masked[3737];
  assign N1582 = N1581 | data_masked[3865];
  assign N1581 = N1580 | data_masked[3993];
  assign N1580 = N1579 | data_masked[4121];
  assign N1579 = N1578 | data_masked[4249];
  assign N1578 = N1577 | data_masked[4377];
  assign N1577 = N1576 | data_masked[4505];
  assign N1576 = N1575 | data_masked[4633];
  assign N1575 = N1574 | data_masked[4761];
  assign N1574 = N1573 | data_masked[4889];
  assign N1573 = N1572 | data_masked[5017];
  assign N1572 = N1571 | data_masked[5145];
  assign N1571 = N1570 | data_masked[5273];
  assign N1570 = N1569 | data_masked[5401];
  assign N1569 = N1568 | data_masked[5529];
  assign N1568 = N1567 | data_masked[5657];
  assign N1567 = N1566 | data_masked[5785];
  assign N1566 = N1565 | data_masked[5913];
  assign N1565 = N1564 | data_masked[6041];
  assign N1564 = N1563 | data_masked[6169];
  assign N1563 = N1562 | data_masked[6297];
  assign N1562 = N1561 | data_masked[6425];
  assign N1561 = N1560 | data_masked[6553];
  assign N1560 = N1559 | data_masked[6681];
  assign N1559 = N1558 | data_masked[6809];
  assign N1558 = N1557 | data_masked[6937];
  assign N1557 = N1556 | data_masked[7065];
  assign N1556 = N1555 | data_masked[7193];
  assign N1555 = N1554 | data_masked[7321];
  assign N1554 = N1553 | data_masked[7449];
  assign N1553 = N1552 | data_masked[7577];
  assign N1552 = N1551 | data_masked[7705];
  assign N1551 = N1550 | data_masked[7833];
  assign N1550 = data_masked[8089] | data_masked[7961];
  assign data_o[26] = N1673 | data_masked[26];
  assign N1673 = N1672 | data_masked[154];
  assign N1672 = N1671 | data_masked[282];
  assign N1671 = N1670 | data_masked[410];
  assign N1670 = N1669 | data_masked[538];
  assign N1669 = N1668 | data_masked[666];
  assign N1668 = N1667 | data_masked[794];
  assign N1667 = N1666 | data_masked[922];
  assign N1666 = N1665 | data_masked[1050];
  assign N1665 = N1664 | data_masked[1178];
  assign N1664 = N1663 | data_masked[1306];
  assign N1663 = N1662 | data_masked[1434];
  assign N1662 = N1661 | data_masked[1562];
  assign N1661 = N1660 | data_masked[1690];
  assign N1660 = N1659 | data_masked[1818];
  assign N1659 = N1658 | data_masked[1946];
  assign N1658 = N1657 | data_masked[2074];
  assign N1657 = N1656 | data_masked[2202];
  assign N1656 = N1655 | data_masked[2330];
  assign N1655 = N1654 | data_masked[2458];
  assign N1654 = N1653 | data_masked[2586];
  assign N1653 = N1652 | data_masked[2714];
  assign N1652 = N1651 | data_masked[2842];
  assign N1651 = N1650 | data_masked[2970];
  assign N1650 = N1649 | data_masked[3098];
  assign N1649 = N1648 | data_masked[3226];
  assign N1648 = N1647 | data_masked[3354];
  assign N1647 = N1646 | data_masked[3482];
  assign N1646 = N1645 | data_masked[3610];
  assign N1645 = N1644 | data_masked[3738];
  assign N1644 = N1643 | data_masked[3866];
  assign N1643 = N1642 | data_masked[3994];
  assign N1642 = N1641 | data_masked[4122];
  assign N1641 = N1640 | data_masked[4250];
  assign N1640 = N1639 | data_masked[4378];
  assign N1639 = N1638 | data_masked[4506];
  assign N1638 = N1637 | data_masked[4634];
  assign N1637 = N1636 | data_masked[4762];
  assign N1636 = N1635 | data_masked[4890];
  assign N1635 = N1634 | data_masked[5018];
  assign N1634 = N1633 | data_masked[5146];
  assign N1633 = N1632 | data_masked[5274];
  assign N1632 = N1631 | data_masked[5402];
  assign N1631 = N1630 | data_masked[5530];
  assign N1630 = N1629 | data_masked[5658];
  assign N1629 = N1628 | data_masked[5786];
  assign N1628 = N1627 | data_masked[5914];
  assign N1627 = N1626 | data_masked[6042];
  assign N1626 = N1625 | data_masked[6170];
  assign N1625 = N1624 | data_masked[6298];
  assign N1624 = N1623 | data_masked[6426];
  assign N1623 = N1622 | data_masked[6554];
  assign N1622 = N1621 | data_masked[6682];
  assign N1621 = N1620 | data_masked[6810];
  assign N1620 = N1619 | data_masked[6938];
  assign N1619 = N1618 | data_masked[7066];
  assign N1618 = N1617 | data_masked[7194];
  assign N1617 = N1616 | data_masked[7322];
  assign N1616 = N1615 | data_masked[7450];
  assign N1615 = N1614 | data_masked[7578];
  assign N1614 = N1613 | data_masked[7706];
  assign N1613 = N1612 | data_masked[7834];
  assign N1612 = data_masked[8090] | data_masked[7962];
  assign data_o[27] = N1735 | data_masked[27];
  assign N1735 = N1734 | data_masked[155];
  assign N1734 = N1733 | data_masked[283];
  assign N1733 = N1732 | data_masked[411];
  assign N1732 = N1731 | data_masked[539];
  assign N1731 = N1730 | data_masked[667];
  assign N1730 = N1729 | data_masked[795];
  assign N1729 = N1728 | data_masked[923];
  assign N1728 = N1727 | data_masked[1051];
  assign N1727 = N1726 | data_masked[1179];
  assign N1726 = N1725 | data_masked[1307];
  assign N1725 = N1724 | data_masked[1435];
  assign N1724 = N1723 | data_masked[1563];
  assign N1723 = N1722 | data_masked[1691];
  assign N1722 = N1721 | data_masked[1819];
  assign N1721 = N1720 | data_masked[1947];
  assign N1720 = N1719 | data_masked[2075];
  assign N1719 = N1718 | data_masked[2203];
  assign N1718 = N1717 | data_masked[2331];
  assign N1717 = N1716 | data_masked[2459];
  assign N1716 = N1715 | data_masked[2587];
  assign N1715 = N1714 | data_masked[2715];
  assign N1714 = N1713 | data_masked[2843];
  assign N1713 = N1712 | data_masked[2971];
  assign N1712 = N1711 | data_masked[3099];
  assign N1711 = N1710 | data_masked[3227];
  assign N1710 = N1709 | data_masked[3355];
  assign N1709 = N1708 | data_masked[3483];
  assign N1708 = N1707 | data_masked[3611];
  assign N1707 = N1706 | data_masked[3739];
  assign N1706 = N1705 | data_masked[3867];
  assign N1705 = N1704 | data_masked[3995];
  assign N1704 = N1703 | data_masked[4123];
  assign N1703 = N1702 | data_masked[4251];
  assign N1702 = N1701 | data_masked[4379];
  assign N1701 = N1700 | data_masked[4507];
  assign N1700 = N1699 | data_masked[4635];
  assign N1699 = N1698 | data_masked[4763];
  assign N1698 = N1697 | data_masked[4891];
  assign N1697 = N1696 | data_masked[5019];
  assign N1696 = N1695 | data_masked[5147];
  assign N1695 = N1694 | data_masked[5275];
  assign N1694 = N1693 | data_masked[5403];
  assign N1693 = N1692 | data_masked[5531];
  assign N1692 = N1691 | data_masked[5659];
  assign N1691 = N1690 | data_masked[5787];
  assign N1690 = N1689 | data_masked[5915];
  assign N1689 = N1688 | data_masked[6043];
  assign N1688 = N1687 | data_masked[6171];
  assign N1687 = N1686 | data_masked[6299];
  assign N1686 = N1685 | data_masked[6427];
  assign N1685 = N1684 | data_masked[6555];
  assign N1684 = N1683 | data_masked[6683];
  assign N1683 = N1682 | data_masked[6811];
  assign N1682 = N1681 | data_masked[6939];
  assign N1681 = N1680 | data_masked[7067];
  assign N1680 = N1679 | data_masked[7195];
  assign N1679 = N1678 | data_masked[7323];
  assign N1678 = N1677 | data_masked[7451];
  assign N1677 = N1676 | data_masked[7579];
  assign N1676 = N1675 | data_masked[7707];
  assign N1675 = N1674 | data_masked[7835];
  assign N1674 = data_masked[8091] | data_masked[7963];
  assign data_o[28] = N1797 | data_masked[28];
  assign N1797 = N1796 | data_masked[156];
  assign N1796 = N1795 | data_masked[284];
  assign N1795 = N1794 | data_masked[412];
  assign N1794 = N1793 | data_masked[540];
  assign N1793 = N1792 | data_masked[668];
  assign N1792 = N1791 | data_masked[796];
  assign N1791 = N1790 | data_masked[924];
  assign N1790 = N1789 | data_masked[1052];
  assign N1789 = N1788 | data_masked[1180];
  assign N1788 = N1787 | data_masked[1308];
  assign N1787 = N1786 | data_masked[1436];
  assign N1786 = N1785 | data_masked[1564];
  assign N1785 = N1784 | data_masked[1692];
  assign N1784 = N1783 | data_masked[1820];
  assign N1783 = N1782 | data_masked[1948];
  assign N1782 = N1781 | data_masked[2076];
  assign N1781 = N1780 | data_masked[2204];
  assign N1780 = N1779 | data_masked[2332];
  assign N1779 = N1778 | data_masked[2460];
  assign N1778 = N1777 | data_masked[2588];
  assign N1777 = N1776 | data_masked[2716];
  assign N1776 = N1775 | data_masked[2844];
  assign N1775 = N1774 | data_masked[2972];
  assign N1774 = N1773 | data_masked[3100];
  assign N1773 = N1772 | data_masked[3228];
  assign N1772 = N1771 | data_masked[3356];
  assign N1771 = N1770 | data_masked[3484];
  assign N1770 = N1769 | data_masked[3612];
  assign N1769 = N1768 | data_masked[3740];
  assign N1768 = N1767 | data_masked[3868];
  assign N1767 = N1766 | data_masked[3996];
  assign N1766 = N1765 | data_masked[4124];
  assign N1765 = N1764 | data_masked[4252];
  assign N1764 = N1763 | data_masked[4380];
  assign N1763 = N1762 | data_masked[4508];
  assign N1762 = N1761 | data_masked[4636];
  assign N1761 = N1760 | data_masked[4764];
  assign N1760 = N1759 | data_masked[4892];
  assign N1759 = N1758 | data_masked[5020];
  assign N1758 = N1757 | data_masked[5148];
  assign N1757 = N1756 | data_masked[5276];
  assign N1756 = N1755 | data_masked[5404];
  assign N1755 = N1754 | data_masked[5532];
  assign N1754 = N1753 | data_masked[5660];
  assign N1753 = N1752 | data_masked[5788];
  assign N1752 = N1751 | data_masked[5916];
  assign N1751 = N1750 | data_masked[6044];
  assign N1750 = N1749 | data_masked[6172];
  assign N1749 = N1748 | data_masked[6300];
  assign N1748 = N1747 | data_masked[6428];
  assign N1747 = N1746 | data_masked[6556];
  assign N1746 = N1745 | data_masked[6684];
  assign N1745 = N1744 | data_masked[6812];
  assign N1744 = N1743 | data_masked[6940];
  assign N1743 = N1742 | data_masked[7068];
  assign N1742 = N1741 | data_masked[7196];
  assign N1741 = N1740 | data_masked[7324];
  assign N1740 = N1739 | data_masked[7452];
  assign N1739 = N1738 | data_masked[7580];
  assign N1738 = N1737 | data_masked[7708];
  assign N1737 = N1736 | data_masked[7836];
  assign N1736 = data_masked[8092] | data_masked[7964];
  assign data_o[29] = N1859 | data_masked[29];
  assign N1859 = N1858 | data_masked[157];
  assign N1858 = N1857 | data_masked[285];
  assign N1857 = N1856 | data_masked[413];
  assign N1856 = N1855 | data_masked[541];
  assign N1855 = N1854 | data_masked[669];
  assign N1854 = N1853 | data_masked[797];
  assign N1853 = N1852 | data_masked[925];
  assign N1852 = N1851 | data_masked[1053];
  assign N1851 = N1850 | data_masked[1181];
  assign N1850 = N1849 | data_masked[1309];
  assign N1849 = N1848 | data_masked[1437];
  assign N1848 = N1847 | data_masked[1565];
  assign N1847 = N1846 | data_masked[1693];
  assign N1846 = N1845 | data_masked[1821];
  assign N1845 = N1844 | data_masked[1949];
  assign N1844 = N1843 | data_masked[2077];
  assign N1843 = N1842 | data_masked[2205];
  assign N1842 = N1841 | data_masked[2333];
  assign N1841 = N1840 | data_masked[2461];
  assign N1840 = N1839 | data_masked[2589];
  assign N1839 = N1838 | data_masked[2717];
  assign N1838 = N1837 | data_masked[2845];
  assign N1837 = N1836 | data_masked[2973];
  assign N1836 = N1835 | data_masked[3101];
  assign N1835 = N1834 | data_masked[3229];
  assign N1834 = N1833 | data_masked[3357];
  assign N1833 = N1832 | data_masked[3485];
  assign N1832 = N1831 | data_masked[3613];
  assign N1831 = N1830 | data_masked[3741];
  assign N1830 = N1829 | data_masked[3869];
  assign N1829 = N1828 | data_masked[3997];
  assign N1828 = N1827 | data_masked[4125];
  assign N1827 = N1826 | data_masked[4253];
  assign N1826 = N1825 | data_masked[4381];
  assign N1825 = N1824 | data_masked[4509];
  assign N1824 = N1823 | data_masked[4637];
  assign N1823 = N1822 | data_masked[4765];
  assign N1822 = N1821 | data_masked[4893];
  assign N1821 = N1820 | data_masked[5021];
  assign N1820 = N1819 | data_masked[5149];
  assign N1819 = N1818 | data_masked[5277];
  assign N1818 = N1817 | data_masked[5405];
  assign N1817 = N1816 | data_masked[5533];
  assign N1816 = N1815 | data_masked[5661];
  assign N1815 = N1814 | data_masked[5789];
  assign N1814 = N1813 | data_masked[5917];
  assign N1813 = N1812 | data_masked[6045];
  assign N1812 = N1811 | data_masked[6173];
  assign N1811 = N1810 | data_masked[6301];
  assign N1810 = N1809 | data_masked[6429];
  assign N1809 = N1808 | data_masked[6557];
  assign N1808 = N1807 | data_masked[6685];
  assign N1807 = N1806 | data_masked[6813];
  assign N1806 = N1805 | data_masked[6941];
  assign N1805 = N1804 | data_masked[7069];
  assign N1804 = N1803 | data_masked[7197];
  assign N1803 = N1802 | data_masked[7325];
  assign N1802 = N1801 | data_masked[7453];
  assign N1801 = N1800 | data_masked[7581];
  assign N1800 = N1799 | data_masked[7709];
  assign N1799 = N1798 | data_masked[7837];
  assign N1798 = data_masked[8093] | data_masked[7965];
  assign data_o[30] = N1921 | data_masked[30];
  assign N1921 = N1920 | data_masked[158];
  assign N1920 = N1919 | data_masked[286];
  assign N1919 = N1918 | data_masked[414];
  assign N1918 = N1917 | data_masked[542];
  assign N1917 = N1916 | data_masked[670];
  assign N1916 = N1915 | data_masked[798];
  assign N1915 = N1914 | data_masked[926];
  assign N1914 = N1913 | data_masked[1054];
  assign N1913 = N1912 | data_masked[1182];
  assign N1912 = N1911 | data_masked[1310];
  assign N1911 = N1910 | data_masked[1438];
  assign N1910 = N1909 | data_masked[1566];
  assign N1909 = N1908 | data_masked[1694];
  assign N1908 = N1907 | data_masked[1822];
  assign N1907 = N1906 | data_masked[1950];
  assign N1906 = N1905 | data_masked[2078];
  assign N1905 = N1904 | data_masked[2206];
  assign N1904 = N1903 | data_masked[2334];
  assign N1903 = N1902 | data_masked[2462];
  assign N1902 = N1901 | data_masked[2590];
  assign N1901 = N1900 | data_masked[2718];
  assign N1900 = N1899 | data_masked[2846];
  assign N1899 = N1898 | data_masked[2974];
  assign N1898 = N1897 | data_masked[3102];
  assign N1897 = N1896 | data_masked[3230];
  assign N1896 = N1895 | data_masked[3358];
  assign N1895 = N1894 | data_masked[3486];
  assign N1894 = N1893 | data_masked[3614];
  assign N1893 = N1892 | data_masked[3742];
  assign N1892 = N1891 | data_masked[3870];
  assign N1891 = N1890 | data_masked[3998];
  assign N1890 = N1889 | data_masked[4126];
  assign N1889 = N1888 | data_masked[4254];
  assign N1888 = N1887 | data_masked[4382];
  assign N1887 = N1886 | data_masked[4510];
  assign N1886 = N1885 | data_masked[4638];
  assign N1885 = N1884 | data_masked[4766];
  assign N1884 = N1883 | data_masked[4894];
  assign N1883 = N1882 | data_masked[5022];
  assign N1882 = N1881 | data_masked[5150];
  assign N1881 = N1880 | data_masked[5278];
  assign N1880 = N1879 | data_masked[5406];
  assign N1879 = N1878 | data_masked[5534];
  assign N1878 = N1877 | data_masked[5662];
  assign N1877 = N1876 | data_masked[5790];
  assign N1876 = N1875 | data_masked[5918];
  assign N1875 = N1874 | data_masked[6046];
  assign N1874 = N1873 | data_masked[6174];
  assign N1873 = N1872 | data_masked[6302];
  assign N1872 = N1871 | data_masked[6430];
  assign N1871 = N1870 | data_masked[6558];
  assign N1870 = N1869 | data_masked[6686];
  assign N1869 = N1868 | data_masked[6814];
  assign N1868 = N1867 | data_masked[6942];
  assign N1867 = N1866 | data_masked[7070];
  assign N1866 = N1865 | data_masked[7198];
  assign N1865 = N1864 | data_masked[7326];
  assign N1864 = N1863 | data_masked[7454];
  assign N1863 = N1862 | data_masked[7582];
  assign N1862 = N1861 | data_masked[7710];
  assign N1861 = N1860 | data_masked[7838];
  assign N1860 = data_masked[8094] | data_masked[7966];
  assign data_o[31] = N1983 | data_masked[31];
  assign N1983 = N1982 | data_masked[159];
  assign N1982 = N1981 | data_masked[287];
  assign N1981 = N1980 | data_masked[415];
  assign N1980 = N1979 | data_masked[543];
  assign N1979 = N1978 | data_masked[671];
  assign N1978 = N1977 | data_masked[799];
  assign N1977 = N1976 | data_masked[927];
  assign N1976 = N1975 | data_masked[1055];
  assign N1975 = N1974 | data_masked[1183];
  assign N1974 = N1973 | data_masked[1311];
  assign N1973 = N1972 | data_masked[1439];
  assign N1972 = N1971 | data_masked[1567];
  assign N1971 = N1970 | data_masked[1695];
  assign N1970 = N1969 | data_masked[1823];
  assign N1969 = N1968 | data_masked[1951];
  assign N1968 = N1967 | data_masked[2079];
  assign N1967 = N1966 | data_masked[2207];
  assign N1966 = N1965 | data_masked[2335];
  assign N1965 = N1964 | data_masked[2463];
  assign N1964 = N1963 | data_masked[2591];
  assign N1963 = N1962 | data_masked[2719];
  assign N1962 = N1961 | data_masked[2847];
  assign N1961 = N1960 | data_masked[2975];
  assign N1960 = N1959 | data_masked[3103];
  assign N1959 = N1958 | data_masked[3231];
  assign N1958 = N1957 | data_masked[3359];
  assign N1957 = N1956 | data_masked[3487];
  assign N1956 = N1955 | data_masked[3615];
  assign N1955 = N1954 | data_masked[3743];
  assign N1954 = N1953 | data_masked[3871];
  assign N1953 = N1952 | data_masked[3999];
  assign N1952 = N1951 | data_masked[4127];
  assign N1951 = N1950 | data_masked[4255];
  assign N1950 = N1949 | data_masked[4383];
  assign N1949 = N1948 | data_masked[4511];
  assign N1948 = N1947 | data_masked[4639];
  assign N1947 = N1946 | data_masked[4767];
  assign N1946 = N1945 | data_masked[4895];
  assign N1945 = N1944 | data_masked[5023];
  assign N1944 = N1943 | data_masked[5151];
  assign N1943 = N1942 | data_masked[5279];
  assign N1942 = N1941 | data_masked[5407];
  assign N1941 = N1940 | data_masked[5535];
  assign N1940 = N1939 | data_masked[5663];
  assign N1939 = N1938 | data_masked[5791];
  assign N1938 = N1937 | data_masked[5919];
  assign N1937 = N1936 | data_masked[6047];
  assign N1936 = N1935 | data_masked[6175];
  assign N1935 = N1934 | data_masked[6303];
  assign N1934 = N1933 | data_masked[6431];
  assign N1933 = N1932 | data_masked[6559];
  assign N1932 = N1931 | data_masked[6687];
  assign N1931 = N1930 | data_masked[6815];
  assign N1930 = N1929 | data_masked[6943];
  assign N1929 = N1928 | data_masked[7071];
  assign N1928 = N1927 | data_masked[7199];
  assign N1927 = N1926 | data_masked[7327];
  assign N1926 = N1925 | data_masked[7455];
  assign N1925 = N1924 | data_masked[7583];
  assign N1924 = N1923 | data_masked[7711];
  assign N1923 = N1922 | data_masked[7839];
  assign N1922 = data_masked[8095] | data_masked[7967];
  assign data_o[32] = N2045 | data_masked[32];
  assign N2045 = N2044 | data_masked[160];
  assign N2044 = N2043 | data_masked[288];
  assign N2043 = N2042 | data_masked[416];
  assign N2042 = N2041 | data_masked[544];
  assign N2041 = N2040 | data_masked[672];
  assign N2040 = N2039 | data_masked[800];
  assign N2039 = N2038 | data_masked[928];
  assign N2038 = N2037 | data_masked[1056];
  assign N2037 = N2036 | data_masked[1184];
  assign N2036 = N2035 | data_masked[1312];
  assign N2035 = N2034 | data_masked[1440];
  assign N2034 = N2033 | data_masked[1568];
  assign N2033 = N2032 | data_masked[1696];
  assign N2032 = N2031 | data_masked[1824];
  assign N2031 = N2030 | data_masked[1952];
  assign N2030 = N2029 | data_masked[2080];
  assign N2029 = N2028 | data_masked[2208];
  assign N2028 = N2027 | data_masked[2336];
  assign N2027 = N2026 | data_masked[2464];
  assign N2026 = N2025 | data_masked[2592];
  assign N2025 = N2024 | data_masked[2720];
  assign N2024 = N2023 | data_masked[2848];
  assign N2023 = N2022 | data_masked[2976];
  assign N2022 = N2021 | data_masked[3104];
  assign N2021 = N2020 | data_masked[3232];
  assign N2020 = N2019 | data_masked[3360];
  assign N2019 = N2018 | data_masked[3488];
  assign N2018 = N2017 | data_masked[3616];
  assign N2017 = N2016 | data_masked[3744];
  assign N2016 = N2015 | data_masked[3872];
  assign N2015 = N2014 | data_masked[4000];
  assign N2014 = N2013 | data_masked[4128];
  assign N2013 = N2012 | data_masked[4256];
  assign N2012 = N2011 | data_masked[4384];
  assign N2011 = N2010 | data_masked[4512];
  assign N2010 = N2009 | data_masked[4640];
  assign N2009 = N2008 | data_masked[4768];
  assign N2008 = N2007 | data_masked[4896];
  assign N2007 = N2006 | data_masked[5024];
  assign N2006 = N2005 | data_masked[5152];
  assign N2005 = N2004 | data_masked[5280];
  assign N2004 = N2003 | data_masked[5408];
  assign N2003 = N2002 | data_masked[5536];
  assign N2002 = N2001 | data_masked[5664];
  assign N2001 = N2000 | data_masked[5792];
  assign N2000 = N1999 | data_masked[5920];
  assign N1999 = N1998 | data_masked[6048];
  assign N1998 = N1997 | data_masked[6176];
  assign N1997 = N1996 | data_masked[6304];
  assign N1996 = N1995 | data_masked[6432];
  assign N1995 = N1994 | data_masked[6560];
  assign N1994 = N1993 | data_masked[6688];
  assign N1993 = N1992 | data_masked[6816];
  assign N1992 = N1991 | data_masked[6944];
  assign N1991 = N1990 | data_masked[7072];
  assign N1990 = N1989 | data_masked[7200];
  assign N1989 = N1988 | data_masked[7328];
  assign N1988 = N1987 | data_masked[7456];
  assign N1987 = N1986 | data_masked[7584];
  assign N1986 = N1985 | data_masked[7712];
  assign N1985 = N1984 | data_masked[7840];
  assign N1984 = data_masked[8096] | data_masked[7968];
  assign data_o[33] = N2107 | data_masked[33];
  assign N2107 = N2106 | data_masked[161];
  assign N2106 = N2105 | data_masked[289];
  assign N2105 = N2104 | data_masked[417];
  assign N2104 = N2103 | data_masked[545];
  assign N2103 = N2102 | data_masked[673];
  assign N2102 = N2101 | data_masked[801];
  assign N2101 = N2100 | data_masked[929];
  assign N2100 = N2099 | data_masked[1057];
  assign N2099 = N2098 | data_masked[1185];
  assign N2098 = N2097 | data_masked[1313];
  assign N2097 = N2096 | data_masked[1441];
  assign N2096 = N2095 | data_masked[1569];
  assign N2095 = N2094 | data_masked[1697];
  assign N2094 = N2093 | data_masked[1825];
  assign N2093 = N2092 | data_masked[1953];
  assign N2092 = N2091 | data_masked[2081];
  assign N2091 = N2090 | data_masked[2209];
  assign N2090 = N2089 | data_masked[2337];
  assign N2089 = N2088 | data_masked[2465];
  assign N2088 = N2087 | data_masked[2593];
  assign N2087 = N2086 | data_masked[2721];
  assign N2086 = N2085 | data_masked[2849];
  assign N2085 = N2084 | data_masked[2977];
  assign N2084 = N2083 | data_masked[3105];
  assign N2083 = N2082 | data_masked[3233];
  assign N2082 = N2081 | data_masked[3361];
  assign N2081 = N2080 | data_masked[3489];
  assign N2080 = N2079 | data_masked[3617];
  assign N2079 = N2078 | data_masked[3745];
  assign N2078 = N2077 | data_masked[3873];
  assign N2077 = N2076 | data_masked[4001];
  assign N2076 = N2075 | data_masked[4129];
  assign N2075 = N2074 | data_masked[4257];
  assign N2074 = N2073 | data_masked[4385];
  assign N2073 = N2072 | data_masked[4513];
  assign N2072 = N2071 | data_masked[4641];
  assign N2071 = N2070 | data_masked[4769];
  assign N2070 = N2069 | data_masked[4897];
  assign N2069 = N2068 | data_masked[5025];
  assign N2068 = N2067 | data_masked[5153];
  assign N2067 = N2066 | data_masked[5281];
  assign N2066 = N2065 | data_masked[5409];
  assign N2065 = N2064 | data_masked[5537];
  assign N2064 = N2063 | data_masked[5665];
  assign N2063 = N2062 | data_masked[5793];
  assign N2062 = N2061 | data_masked[5921];
  assign N2061 = N2060 | data_masked[6049];
  assign N2060 = N2059 | data_masked[6177];
  assign N2059 = N2058 | data_masked[6305];
  assign N2058 = N2057 | data_masked[6433];
  assign N2057 = N2056 | data_masked[6561];
  assign N2056 = N2055 | data_masked[6689];
  assign N2055 = N2054 | data_masked[6817];
  assign N2054 = N2053 | data_masked[6945];
  assign N2053 = N2052 | data_masked[7073];
  assign N2052 = N2051 | data_masked[7201];
  assign N2051 = N2050 | data_masked[7329];
  assign N2050 = N2049 | data_masked[7457];
  assign N2049 = N2048 | data_masked[7585];
  assign N2048 = N2047 | data_masked[7713];
  assign N2047 = N2046 | data_masked[7841];
  assign N2046 = data_masked[8097] | data_masked[7969];
  assign data_o[34] = N2169 | data_masked[34];
  assign N2169 = N2168 | data_masked[162];
  assign N2168 = N2167 | data_masked[290];
  assign N2167 = N2166 | data_masked[418];
  assign N2166 = N2165 | data_masked[546];
  assign N2165 = N2164 | data_masked[674];
  assign N2164 = N2163 | data_masked[802];
  assign N2163 = N2162 | data_masked[930];
  assign N2162 = N2161 | data_masked[1058];
  assign N2161 = N2160 | data_masked[1186];
  assign N2160 = N2159 | data_masked[1314];
  assign N2159 = N2158 | data_masked[1442];
  assign N2158 = N2157 | data_masked[1570];
  assign N2157 = N2156 | data_masked[1698];
  assign N2156 = N2155 | data_masked[1826];
  assign N2155 = N2154 | data_masked[1954];
  assign N2154 = N2153 | data_masked[2082];
  assign N2153 = N2152 | data_masked[2210];
  assign N2152 = N2151 | data_masked[2338];
  assign N2151 = N2150 | data_masked[2466];
  assign N2150 = N2149 | data_masked[2594];
  assign N2149 = N2148 | data_masked[2722];
  assign N2148 = N2147 | data_masked[2850];
  assign N2147 = N2146 | data_masked[2978];
  assign N2146 = N2145 | data_masked[3106];
  assign N2145 = N2144 | data_masked[3234];
  assign N2144 = N2143 | data_masked[3362];
  assign N2143 = N2142 | data_masked[3490];
  assign N2142 = N2141 | data_masked[3618];
  assign N2141 = N2140 | data_masked[3746];
  assign N2140 = N2139 | data_masked[3874];
  assign N2139 = N2138 | data_masked[4002];
  assign N2138 = N2137 | data_masked[4130];
  assign N2137 = N2136 | data_masked[4258];
  assign N2136 = N2135 | data_masked[4386];
  assign N2135 = N2134 | data_masked[4514];
  assign N2134 = N2133 | data_masked[4642];
  assign N2133 = N2132 | data_masked[4770];
  assign N2132 = N2131 | data_masked[4898];
  assign N2131 = N2130 | data_masked[5026];
  assign N2130 = N2129 | data_masked[5154];
  assign N2129 = N2128 | data_masked[5282];
  assign N2128 = N2127 | data_masked[5410];
  assign N2127 = N2126 | data_masked[5538];
  assign N2126 = N2125 | data_masked[5666];
  assign N2125 = N2124 | data_masked[5794];
  assign N2124 = N2123 | data_masked[5922];
  assign N2123 = N2122 | data_masked[6050];
  assign N2122 = N2121 | data_masked[6178];
  assign N2121 = N2120 | data_masked[6306];
  assign N2120 = N2119 | data_masked[6434];
  assign N2119 = N2118 | data_masked[6562];
  assign N2118 = N2117 | data_masked[6690];
  assign N2117 = N2116 | data_masked[6818];
  assign N2116 = N2115 | data_masked[6946];
  assign N2115 = N2114 | data_masked[7074];
  assign N2114 = N2113 | data_masked[7202];
  assign N2113 = N2112 | data_masked[7330];
  assign N2112 = N2111 | data_masked[7458];
  assign N2111 = N2110 | data_masked[7586];
  assign N2110 = N2109 | data_masked[7714];
  assign N2109 = N2108 | data_masked[7842];
  assign N2108 = data_masked[8098] | data_masked[7970];
  assign data_o[35] = N2231 | data_masked[35];
  assign N2231 = N2230 | data_masked[163];
  assign N2230 = N2229 | data_masked[291];
  assign N2229 = N2228 | data_masked[419];
  assign N2228 = N2227 | data_masked[547];
  assign N2227 = N2226 | data_masked[675];
  assign N2226 = N2225 | data_masked[803];
  assign N2225 = N2224 | data_masked[931];
  assign N2224 = N2223 | data_masked[1059];
  assign N2223 = N2222 | data_masked[1187];
  assign N2222 = N2221 | data_masked[1315];
  assign N2221 = N2220 | data_masked[1443];
  assign N2220 = N2219 | data_masked[1571];
  assign N2219 = N2218 | data_masked[1699];
  assign N2218 = N2217 | data_masked[1827];
  assign N2217 = N2216 | data_masked[1955];
  assign N2216 = N2215 | data_masked[2083];
  assign N2215 = N2214 | data_masked[2211];
  assign N2214 = N2213 | data_masked[2339];
  assign N2213 = N2212 | data_masked[2467];
  assign N2212 = N2211 | data_masked[2595];
  assign N2211 = N2210 | data_masked[2723];
  assign N2210 = N2209 | data_masked[2851];
  assign N2209 = N2208 | data_masked[2979];
  assign N2208 = N2207 | data_masked[3107];
  assign N2207 = N2206 | data_masked[3235];
  assign N2206 = N2205 | data_masked[3363];
  assign N2205 = N2204 | data_masked[3491];
  assign N2204 = N2203 | data_masked[3619];
  assign N2203 = N2202 | data_masked[3747];
  assign N2202 = N2201 | data_masked[3875];
  assign N2201 = N2200 | data_masked[4003];
  assign N2200 = N2199 | data_masked[4131];
  assign N2199 = N2198 | data_masked[4259];
  assign N2198 = N2197 | data_masked[4387];
  assign N2197 = N2196 | data_masked[4515];
  assign N2196 = N2195 | data_masked[4643];
  assign N2195 = N2194 | data_masked[4771];
  assign N2194 = N2193 | data_masked[4899];
  assign N2193 = N2192 | data_masked[5027];
  assign N2192 = N2191 | data_masked[5155];
  assign N2191 = N2190 | data_masked[5283];
  assign N2190 = N2189 | data_masked[5411];
  assign N2189 = N2188 | data_masked[5539];
  assign N2188 = N2187 | data_masked[5667];
  assign N2187 = N2186 | data_masked[5795];
  assign N2186 = N2185 | data_masked[5923];
  assign N2185 = N2184 | data_masked[6051];
  assign N2184 = N2183 | data_masked[6179];
  assign N2183 = N2182 | data_masked[6307];
  assign N2182 = N2181 | data_masked[6435];
  assign N2181 = N2180 | data_masked[6563];
  assign N2180 = N2179 | data_masked[6691];
  assign N2179 = N2178 | data_masked[6819];
  assign N2178 = N2177 | data_masked[6947];
  assign N2177 = N2176 | data_masked[7075];
  assign N2176 = N2175 | data_masked[7203];
  assign N2175 = N2174 | data_masked[7331];
  assign N2174 = N2173 | data_masked[7459];
  assign N2173 = N2172 | data_masked[7587];
  assign N2172 = N2171 | data_masked[7715];
  assign N2171 = N2170 | data_masked[7843];
  assign N2170 = data_masked[8099] | data_masked[7971];
  assign data_o[36] = N2293 | data_masked[36];
  assign N2293 = N2292 | data_masked[164];
  assign N2292 = N2291 | data_masked[292];
  assign N2291 = N2290 | data_masked[420];
  assign N2290 = N2289 | data_masked[548];
  assign N2289 = N2288 | data_masked[676];
  assign N2288 = N2287 | data_masked[804];
  assign N2287 = N2286 | data_masked[932];
  assign N2286 = N2285 | data_masked[1060];
  assign N2285 = N2284 | data_masked[1188];
  assign N2284 = N2283 | data_masked[1316];
  assign N2283 = N2282 | data_masked[1444];
  assign N2282 = N2281 | data_masked[1572];
  assign N2281 = N2280 | data_masked[1700];
  assign N2280 = N2279 | data_masked[1828];
  assign N2279 = N2278 | data_masked[1956];
  assign N2278 = N2277 | data_masked[2084];
  assign N2277 = N2276 | data_masked[2212];
  assign N2276 = N2275 | data_masked[2340];
  assign N2275 = N2274 | data_masked[2468];
  assign N2274 = N2273 | data_masked[2596];
  assign N2273 = N2272 | data_masked[2724];
  assign N2272 = N2271 | data_masked[2852];
  assign N2271 = N2270 | data_masked[2980];
  assign N2270 = N2269 | data_masked[3108];
  assign N2269 = N2268 | data_masked[3236];
  assign N2268 = N2267 | data_masked[3364];
  assign N2267 = N2266 | data_masked[3492];
  assign N2266 = N2265 | data_masked[3620];
  assign N2265 = N2264 | data_masked[3748];
  assign N2264 = N2263 | data_masked[3876];
  assign N2263 = N2262 | data_masked[4004];
  assign N2262 = N2261 | data_masked[4132];
  assign N2261 = N2260 | data_masked[4260];
  assign N2260 = N2259 | data_masked[4388];
  assign N2259 = N2258 | data_masked[4516];
  assign N2258 = N2257 | data_masked[4644];
  assign N2257 = N2256 | data_masked[4772];
  assign N2256 = N2255 | data_masked[4900];
  assign N2255 = N2254 | data_masked[5028];
  assign N2254 = N2253 | data_masked[5156];
  assign N2253 = N2252 | data_masked[5284];
  assign N2252 = N2251 | data_masked[5412];
  assign N2251 = N2250 | data_masked[5540];
  assign N2250 = N2249 | data_masked[5668];
  assign N2249 = N2248 | data_masked[5796];
  assign N2248 = N2247 | data_masked[5924];
  assign N2247 = N2246 | data_masked[6052];
  assign N2246 = N2245 | data_masked[6180];
  assign N2245 = N2244 | data_masked[6308];
  assign N2244 = N2243 | data_masked[6436];
  assign N2243 = N2242 | data_masked[6564];
  assign N2242 = N2241 | data_masked[6692];
  assign N2241 = N2240 | data_masked[6820];
  assign N2240 = N2239 | data_masked[6948];
  assign N2239 = N2238 | data_masked[7076];
  assign N2238 = N2237 | data_masked[7204];
  assign N2237 = N2236 | data_masked[7332];
  assign N2236 = N2235 | data_masked[7460];
  assign N2235 = N2234 | data_masked[7588];
  assign N2234 = N2233 | data_masked[7716];
  assign N2233 = N2232 | data_masked[7844];
  assign N2232 = data_masked[8100] | data_masked[7972];
  assign data_o[37] = N2355 | data_masked[37];
  assign N2355 = N2354 | data_masked[165];
  assign N2354 = N2353 | data_masked[293];
  assign N2353 = N2352 | data_masked[421];
  assign N2352 = N2351 | data_masked[549];
  assign N2351 = N2350 | data_masked[677];
  assign N2350 = N2349 | data_masked[805];
  assign N2349 = N2348 | data_masked[933];
  assign N2348 = N2347 | data_masked[1061];
  assign N2347 = N2346 | data_masked[1189];
  assign N2346 = N2345 | data_masked[1317];
  assign N2345 = N2344 | data_masked[1445];
  assign N2344 = N2343 | data_masked[1573];
  assign N2343 = N2342 | data_masked[1701];
  assign N2342 = N2341 | data_masked[1829];
  assign N2341 = N2340 | data_masked[1957];
  assign N2340 = N2339 | data_masked[2085];
  assign N2339 = N2338 | data_masked[2213];
  assign N2338 = N2337 | data_masked[2341];
  assign N2337 = N2336 | data_masked[2469];
  assign N2336 = N2335 | data_masked[2597];
  assign N2335 = N2334 | data_masked[2725];
  assign N2334 = N2333 | data_masked[2853];
  assign N2333 = N2332 | data_masked[2981];
  assign N2332 = N2331 | data_masked[3109];
  assign N2331 = N2330 | data_masked[3237];
  assign N2330 = N2329 | data_masked[3365];
  assign N2329 = N2328 | data_masked[3493];
  assign N2328 = N2327 | data_masked[3621];
  assign N2327 = N2326 | data_masked[3749];
  assign N2326 = N2325 | data_masked[3877];
  assign N2325 = N2324 | data_masked[4005];
  assign N2324 = N2323 | data_masked[4133];
  assign N2323 = N2322 | data_masked[4261];
  assign N2322 = N2321 | data_masked[4389];
  assign N2321 = N2320 | data_masked[4517];
  assign N2320 = N2319 | data_masked[4645];
  assign N2319 = N2318 | data_masked[4773];
  assign N2318 = N2317 | data_masked[4901];
  assign N2317 = N2316 | data_masked[5029];
  assign N2316 = N2315 | data_masked[5157];
  assign N2315 = N2314 | data_masked[5285];
  assign N2314 = N2313 | data_masked[5413];
  assign N2313 = N2312 | data_masked[5541];
  assign N2312 = N2311 | data_masked[5669];
  assign N2311 = N2310 | data_masked[5797];
  assign N2310 = N2309 | data_masked[5925];
  assign N2309 = N2308 | data_masked[6053];
  assign N2308 = N2307 | data_masked[6181];
  assign N2307 = N2306 | data_masked[6309];
  assign N2306 = N2305 | data_masked[6437];
  assign N2305 = N2304 | data_masked[6565];
  assign N2304 = N2303 | data_masked[6693];
  assign N2303 = N2302 | data_masked[6821];
  assign N2302 = N2301 | data_masked[6949];
  assign N2301 = N2300 | data_masked[7077];
  assign N2300 = N2299 | data_masked[7205];
  assign N2299 = N2298 | data_masked[7333];
  assign N2298 = N2297 | data_masked[7461];
  assign N2297 = N2296 | data_masked[7589];
  assign N2296 = N2295 | data_masked[7717];
  assign N2295 = N2294 | data_masked[7845];
  assign N2294 = data_masked[8101] | data_masked[7973];
  assign data_o[38] = N2417 | data_masked[38];
  assign N2417 = N2416 | data_masked[166];
  assign N2416 = N2415 | data_masked[294];
  assign N2415 = N2414 | data_masked[422];
  assign N2414 = N2413 | data_masked[550];
  assign N2413 = N2412 | data_masked[678];
  assign N2412 = N2411 | data_masked[806];
  assign N2411 = N2410 | data_masked[934];
  assign N2410 = N2409 | data_masked[1062];
  assign N2409 = N2408 | data_masked[1190];
  assign N2408 = N2407 | data_masked[1318];
  assign N2407 = N2406 | data_masked[1446];
  assign N2406 = N2405 | data_masked[1574];
  assign N2405 = N2404 | data_masked[1702];
  assign N2404 = N2403 | data_masked[1830];
  assign N2403 = N2402 | data_masked[1958];
  assign N2402 = N2401 | data_masked[2086];
  assign N2401 = N2400 | data_masked[2214];
  assign N2400 = N2399 | data_masked[2342];
  assign N2399 = N2398 | data_masked[2470];
  assign N2398 = N2397 | data_masked[2598];
  assign N2397 = N2396 | data_masked[2726];
  assign N2396 = N2395 | data_masked[2854];
  assign N2395 = N2394 | data_masked[2982];
  assign N2394 = N2393 | data_masked[3110];
  assign N2393 = N2392 | data_masked[3238];
  assign N2392 = N2391 | data_masked[3366];
  assign N2391 = N2390 | data_masked[3494];
  assign N2390 = N2389 | data_masked[3622];
  assign N2389 = N2388 | data_masked[3750];
  assign N2388 = N2387 | data_masked[3878];
  assign N2387 = N2386 | data_masked[4006];
  assign N2386 = N2385 | data_masked[4134];
  assign N2385 = N2384 | data_masked[4262];
  assign N2384 = N2383 | data_masked[4390];
  assign N2383 = N2382 | data_masked[4518];
  assign N2382 = N2381 | data_masked[4646];
  assign N2381 = N2380 | data_masked[4774];
  assign N2380 = N2379 | data_masked[4902];
  assign N2379 = N2378 | data_masked[5030];
  assign N2378 = N2377 | data_masked[5158];
  assign N2377 = N2376 | data_masked[5286];
  assign N2376 = N2375 | data_masked[5414];
  assign N2375 = N2374 | data_masked[5542];
  assign N2374 = N2373 | data_masked[5670];
  assign N2373 = N2372 | data_masked[5798];
  assign N2372 = N2371 | data_masked[5926];
  assign N2371 = N2370 | data_masked[6054];
  assign N2370 = N2369 | data_masked[6182];
  assign N2369 = N2368 | data_masked[6310];
  assign N2368 = N2367 | data_masked[6438];
  assign N2367 = N2366 | data_masked[6566];
  assign N2366 = N2365 | data_masked[6694];
  assign N2365 = N2364 | data_masked[6822];
  assign N2364 = N2363 | data_masked[6950];
  assign N2363 = N2362 | data_masked[7078];
  assign N2362 = N2361 | data_masked[7206];
  assign N2361 = N2360 | data_masked[7334];
  assign N2360 = N2359 | data_masked[7462];
  assign N2359 = N2358 | data_masked[7590];
  assign N2358 = N2357 | data_masked[7718];
  assign N2357 = N2356 | data_masked[7846];
  assign N2356 = data_masked[8102] | data_masked[7974];
  assign data_o[39] = N2479 | data_masked[39];
  assign N2479 = N2478 | data_masked[167];
  assign N2478 = N2477 | data_masked[295];
  assign N2477 = N2476 | data_masked[423];
  assign N2476 = N2475 | data_masked[551];
  assign N2475 = N2474 | data_masked[679];
  assign N2474 = N2473 | data_masked[807];
  assign N2473 = N2472 | data_masked[935];
  assign N2472 = N2471 | data_masked[1063];
  assign N2471 = N2470 | data_masked[1191];
  assign N2470 = N2469 | data_masked[1319];
  assign N2469 = N2468 | data_masked[1447];
  assign N2468 = N2467 | data_masked[1575];
  assign N2467 = N2466 | data_masked[1703];
  assign N2466 = N2465 | data_masked[1831];
  assign N2465 = N2464 | data_masked[1959];
  assign N2464 = N2463 | data_masked[2087];
  assign N2463 = N2462 | data_masked[2215];
  assign N2462 = N2461 | data_masked[2343];
  assign N2461 = N2460 | data_masked[2471];
  assign N2460 = N2459 | data_masked[2599];
  assign N2459 = N2458 | data_masked[2727];
  assign N2458 = N2457 | data_masked[2855];
  assign N2457 = N2456 | data_masked[2983];
  assign N2456 = N2455 | data_masked[3111];
  assign N2455 = N2454 | data_masked[3239];
  assign N2454 = N2453 | data_masked[3367];
  assign N2453 = N2452 | data_masked[3495];
  assign N2452 = N2451 | data_masked[3623];
  assign N2451 = N2450 | data_masked[3751];
  assign N2450 = N2449 | data_masked[3879];
  assign N2449 = N2448 | data_masked[4007];
  assign N2448 = N2447 | data_masked[4135];
  assign N2447 = N2446 | data_masked[4263];
  assign N2446 = N2445 | data_masked[4391];
  assign N2445 = N2444 | data_masked[4519];
  assign N2444 = N2443 | data_masked[4647];
  assign N2443 = N2442 | data_masked[4775];
  assign N2442 = N2441 | data_masked[4903];
  assign N2441 = N2440 | data_masked[5031];
  assign N2440 = N2439 | data_masked[5159];
  assign N2439 = N2438 | data_masked[5287];
  assign N2438 = N2437 | data_masked[5415];
  assign N2437 = N2436 | data_masked[5543];
  assign N2436 = N2435 | data_masked[5671];
  assign N2435 = N2434 | data_masked[5799];
  assign N2434 = N2433 | data_masked[5927];
  assign N2433 = N2432 | data_masked[6055];
  assign N2432 = N2431 | data_masked[6183];
  assign N2431 = N2430 | data_masked[6311];
  assign N2430 = N2429 | data_masked[6439];
  assign N2429 = N2428 | data_masked[6567];
  assign N2428 = N2427 | data_masked[6695];
  assign N2427 = N2426 | data_masked[6823];
  assign N2426 = N2425 | data_masked[6951];
  assign N2425 = N2424 | data_masked[7079];
  assign N2424 = N2423 | data_masked[7207];
  assign N2423 = N2422 | data_masked[7335];
  assign N2422 = N2421 | data_masked[7463];
  assign N2421 = N2420 | data_masked[7591];
  assign N2420 = N2419 | data_masked[7719];
  assign N2419 = N2418 | data_masked[7847];
  assign N2418 = data_masked[8103] | data_masked[7975];
  assign data_o[40] = N2541 | data_masked[40];
  assign N2541 = N2540 | data_masked[168];
  assign N2540 = N2539 | data_masked[296];
  assign N2539 = N2538 | data_masked[424];
  assign N2538 = N2537 | data_masked[552];
  assign N2537 = N2536 | data_masked[680];
  assign N2536 = N2535 | data_masked[808];
  assign N2535 = N2534 | data_masked[936];
  assign N2534 = N2533 | data_masked[1064];
  assign N2533 = N2532 | data_masked[1192];
  assign N2532 = N2531 | data_masked[1320];
  assign N2531 = N2530 | data_masked[1448];
  assign N2530 = N2529 | data_masked[1576];
  assign N2529 = N2528 | data_masked[1704];
  assign N2528 = N2527 | data_masked[1832];
  assign N2527 = N2526 | data_masked[1960];
  assign N2526 = N2525 | data_masked[2088];
  assign N2525 = N2524 | data_masked[2216];
  assign N2524 = N2523 | data_masked[2344];
  assign N2523 = N2522 | data_masked[2472];
  assign N2522 = N2521 | data_masked[2600];
  assign N2521 = N2520 | data_masked[2728];
  assign N2520 = N2519 | data_masked[2856];
  assign N2519 = N2518 | data_masked[2984];
  assign N2518 = N2517 | data_masked[3112];
  assign N2517 = N2516 | data_masked[3240];
  assign N2516 = N2515 | data_masked[3368];
  assign N2515 = N2514 | data_masked[3496];
  assign N2514 = N2513 | data_masked[3624];
  assign N2513 = N2512 | data_masked[3752];
  assign N2512 = N2511 | data_masked[3880];
  assign N2511 = N2510 | data_masked[4008];
  assign N2510 = N2509 | data_masked[4136];
  assign N2509 = N2508 | data_masked[4264];
  assign N2508 = N2507 | data_masked[4392];
  assign N2507 = N2506 | data_masked[4520];
  assign N2506 = N2505 | data_masked[4648];
  assign N2505 = N2504 | data_masked[4776];
  assign N2504 = N2503 | data_masked[4904];
  assign N2503 = N2502 | data_masked[5032];
  assign N2502 = N2501 | data_masked[5160];
  assign N2501 = N2500 | data_masked[5288];
  assign N2500 = N2499 | data_masked[5416];
  assign N2499 = N2498 | data_masked[5544];
  assign N2498 = N2497 | data_masked[5672];
  assign N2497 = N2496 | data_masked[5800];
  assign N2496 = N2495 | data_masked[5928];
  assign N2495 = N2494 | data_masked[6056];
  assign N2494 = N2493 | data_masked[6184];
  assign N2493 = N2492 | data_masked[6312];
  assign N2492 = N2491 | data_masked[6440];
  assign N2491 = N2490 | data_masked[6568];
  assign N2490 = N2489 | data_masked[6696];
  assign N2489 = N2488 | data_masked[6824];
  assign N2488 = N2487 | data_masked[6952];
  assign N2487 = N2486 | data_masked[7080];
  assign N2486 = N2485 | data_masked[7208];
  assign N2485 = N2484 | data_masked[7336];
  assign N2484 = N2483 | data_masked[7464];
  assign N2483 = N2482 | data_masked[7592];
  assign N2482 = N2481 | data_masked[7720];
  assign N2481 = N2480 | data_masked[7848];
  assign N2480 = data_masked[8104] | data_masked[7976];
  assign data_o[41] = N2603 | data_masked[41];
  assign N2603 = N2602 | data_masked[169];
  assign N2602 = N2601 | data_masked[297];
  assign N2601 = N2600 | data_masked[425];
  assign N2600 = N2599 | data_masked[553];
  assign N2599 = N2598 | data_masked[681];
  assign N2598 = N2597 | data_masked[809];
  assign N2597 = N2596 | data_masked[937];
  assign N2596 = N2595 | data_masked[1065];
  assign N2595 = N2594 | data_masked[1193];
  assign N2594 = N2593 | data_masked[1321];
  assign N2593 = N2592 | data_masked[1449];
  assign N2592 = N2591 | data_masked[1577];
  assign N2591 = N2590 | data_masked[1705];
  assign N2590 = N2589 | data_masked[1833];
  assign N2589 = N2588 | data_masked[1961];
  assign N2588 = N2587 | data_masked[2089];
  assign N2587 = N2586 | data_masked[2217];
  assign N2586 = N2585 | data_masked[2345];
  assign N2585 = N2584 | data_masked[2473];
  assign N2584 = N2583 | data_masked[2601];
  assign N2583 = N2582 | data_masked[2729];
  assign N2582 = N2581 | data_masked[2857];
  assign N2581 = N2580 | data_masked[2985];
  assign N2580 = N2579 | data_masked[3113];
  assign N2579 = N2578 | data_masked[3241];
  assign N2578 = N2577 | data_masked[3369];
  assign N2577 = N2576 | data_masked[3497];
  assign N2576 = N2575 | data_masked[3625];
  assign N2575 = N2574 | data_masked[3753];
  assign N2574 = N2573 | data_masked[3881];
  assign N2573 = N2572 | data_masked[4009];
  assign N2572 = N2571 | data_masked[4137];
  assign N2571 = N2570 | data_masked[4265];
  assign N2570 = N2569 | data_masked[4393];
  assign N2569 = N2568 | data_masked[4521];
  assign N2568 = N2567 | data_masked[4649];
  assign N2567 = N2566 | data_masked[4777];
  assign N2566 = N2565 | data_masked[4905];
  assign N2565 = N2564 | data_masked[5033];
  assign N2564 = N2563 | data_masked[5161];
  assign N2563 = N2562 | data_masked[5289];
  assign N2562 = N2561 | data_masked[5417];
  assign N2561 = N2560 | data_masked[5545];
  assign N2560 = N2559 | data_masked[5673];
  assign N2559 = N2558 | data_masked[5801];
  assign N2558 = N2557 | data_masked[5929];
  assign N2557 = N2556 | data_masked[6057];
  assign N2556 = N2555 | data_masked[6185];
  assign N2555 = N2554 | data_masked[6313];
  assign N2554 = N2553 | data_masked[6441];
  assign N2553 = N2552 | data_masked[6569];
  assign N2552 = N2551 | data_masked[6697];
  assign N2551 = N2550 | data_masked[6825];
  assign N2550 = N2549 | data_masked[6953];
  assign N2549 = N2548 | data_masked[7081];
  assign N2548 = N2547 | data_masked[7209];
  assign N2547 = N2546 | data_masked[7337];
  assign N2546 = N2545 | data_masked[7465];
  assign N2545 = N2544 | data_masked[7593];
  assign N2544 = N2543 | data_masked[7721];
  assign N2543 = N2542 | data_masked[7849];
  assign N2542 = data_masked[8105] | data_masked[7977];
  assign data_o[42] = N2665 | data_masked[42];
  assign N2665 = N2664 | data_masked[170];
  assign N2664 = N2663 | data_masked[298];
  assign N2663 = N2662 | data_masked[426];
  assign N2662 = N2661 | data_masked[554];
  assign N2661 = N2660 | data_masked[682];
  assign N2660 = N2659 | data_masked[810];
  assign N2659 = N2658 | data_masked[938];
  assign N2658 = N2657 | data_masked[1066];
  assign N2657 = N2656 | data_masked[1194];
  assign N2656 = N2655 | data_masked[1322];
  assign N2655 = N2654 | data_masked[1450];
  assign N2654 = N2653 | data_masked[1578];
  assign N2653 = N2652 | data_masked[1706];
  assign N2652 = N2651 | data_masked[1834];
  assign N2651 = N2650 | data_masked[1962];
  assign N2650 = N2649 | data_masked[2090];
  assign N2649 = N2648 | data_masked[2218];
  assign N2648 = N2647 | data_masked[2346];
  assign N2647 = N2646 | data_masked[2474];
  assign N2646 = N2645 | data_masked[2602];
  assign N2645 = N2644 | data_masked[2730];
  assign N2644 = N2643 | data_masked[2858];
  assign N2643 = N2642 | data_masked[2986];
  assign N2642 = N2641 | data_masked[3114];
  assign N2641 = N2640 | data_masked[3242];
  assign N2640 = N2639 | data_masked[3370];
  assign N2639 = N2638 | data_masked[3498];
  assign N2638 = N2637 | data_masked[3626];
  assign N2637 = N2636 | data_masked[3754];
  assign N2636 = N2635 | data_masked[3882];
  assign N2635 = N2634 | data_masked[4010];
  assign N2634 = N2633 | data_masked[4138];
  assign N2633 = N2632 | data_masked[4266];
  assign N2632 = N2631 | data_masked[4394];
  assign N2631 = N2630 | data_masked[4522];
  assign N2630 = N2629 | data_masked[4650];
  assign N2629 = N2628 | data_masked[4778];
  assign N2628 = N2627 | data_masked[4906];
  assign N2627 = N2626 | data_masked[5034];
  assign N2626 = N2625 | data_masked[5162];
  assign N2625 = N2624 | data_masked[5290];
  assign N2624 = N2623 | data_masked[5418];
  assign N2623 = N2622 | data_masked[5546];
  assign N2622 = N2621 | data_masked[5674];
  assign N2621 = N2620 | data_masked[5802];
  assign N2620 = N2619 | data_masked[5930];
  assign N2619 = N2618 | data_masked[6058];
  assign N2618 = N2617 | data_masked[6186];
  assign N2617 = N2616 | data_masked[6314];
  assign N2616 = N2615 | data_masked[6442];
  assign N2615 = N2614 | data_masked[6570];
  assign N2614 = N2613 | data_masked[6698];
  assign N2613 = N2612 | data_masked[6826];
  assign N2612 = N2611 | data_masked[6954];
  assign N2611 = N2610 | data_masked[7082];
  assign N2610 = N2609 | data_masked[7210];
  assign N2609 = N2608 | data_masked[7338];
  assign N2608 = N2607 | data_masked[7466];
  assign N2607 = N2606 | data_masked[7594];
  assign N2606 = N2605 | data_masked[7722];
  assign N2605 = N2604 | data_masked[7850];
  assign N2604 = data_masked[8106] | data_masked[7978];
  assign data_o[43] = N2727 | data_masked[43];
  assign N2727 = N2726 | data_masked[171];
  assign N2726 = N2725 | data_masked[299];
  assign N2725 = N2724 | data_masked[427];
  assign N2724 = N2723 | data_masked[555];
  assign N2723 = N2722 | data_masked[683];
  assign N2722 = N2721 | data_masked[811];
  assign N2721 = N2720 | data_masked[939];
  assign N2720 = N2719 | data_masked[1067];
  assign N2719 = N2718 | data_masked[1195];
  assign N2718 = N2717 | data_masked[1323];
  assign N2717 = N2716 | data_masked[1451];
  assign N2716 = N2715 | data_masked[1579];
  assign N2715 = N2714 | data_masked[1707];
  assign N2714 = N2713 | data_masked[1835];
  assign N2713 = N2712 | data_masked[1963];
  assign N2712 = N2711 | data_masked[2091];
  assign N2711 = N2710 | data_masked[2219];
  assign N2710 = N2709 | data_masked[2347];
  assign N2709 = N2708 | data_masked[2475];
  assign N2708 = N2707 | data_masked[2603];
  assign N2707 = N2706 | data_masked[2731];
  assign N2706 = N2705 | data_masked[2859];
  assign N2705 = N2704 | data_masked[2987];
  assign N2704 = N2703 | data_masked[3115];
  assign N2703 = N2702 | data_masked[3243];
  assign N2702 = N2701 | data_masked[3371];
  assign N2701 = N2700 | data_masked[3499];
  assign N2700 = N2699 | data_masked[3627];
  assign N2699 = N2698 | data_masked[3755];
  assign N2698 = N2697 | data_masked[3883];
  assign N2697 = N2696 | data_masked[4011];
  assign N2696 = N2695 | data_masked[4139];
  assign N2695 = N2694 | data_masked[4267];
  assign N2694 = N2693 | data_masked[4395];
  assign N2693 = N2692 | data_masked[4523];
  assign N2692 = N2691 | data_masked[4651];
  assign N2691 = N2690 | data_masked[4779];
  assign N2690 = N2689 | data_masked[4907];
  assign N2689 = N2688 | data_masked[5035];
  assign N2688 = N2687 | data_masked[5163];
  assign N2687 = N2686 | data_masked[5291];
  assign N2686 = N2685 | data_masked[5419];
  assign N2685 = N2684 | data_masked[5547];
  assign N2684 = N2683 | data_masked[5675];
  assign N2683 = N2682 | data_masked[5803];
  assign N2682 = N2681 | data_masked[5931];
  assign N2681 = N2680 | data_masked[6059];
  assign N2680 = N2679 | data_masked[6187];
  assign N2679 = N2678 | data_masked[6315];
  assign N2678 = N2677 | data_masked[6443];
  assign N2677 = N2676 | data_masked[6571];
  assign N2676 = N2675 | data_masked[6699];
  assign N2675 = N2674 | data_masked[6827];
  assign N2674 = N2673 | data_masked[6955];
  assign N2673 = N2672 | data_masked[7083];
  assign N2672 = N2671 | data_masked[7211];
  assign N2671 = N2670 | data_masked[7339];
  assign N2670 = N2669 | data_masked[7467];
  assign N2669 = N2668 | data_masked[7595];
  assign N2668 = N2667 | data_masked[7723];
  assign N2667 = N2666 | data_masked[7851];
  assign N2666 = data_masked[8107] | data_masked[7979];
  assign data_o[44] = N2789 | data_masked[44];
  assign N2789 = N2788 | data_masked[172];
  assign N2788 = N2787 | data_masked[300];
  assign N2787 = N2786 | data_masked[428];
  assign N2786 = N2785 | data_masked[556];
  assign N2785 = N2784 | data_masked[684];
  assign N2784 = N2783 | data_masked[812];
  assign N2783 = N2782 | data_masked[940];
  assign N2782 = N2781 | data_masked[1068];
  assign N2781 = N2780 | data_masked[1196];
  assign N2780 = N2779 | data_masked[1324];
  assign N2779 = N2778 | data_masked[1452];
  assign N2778 = N2777 | data_masked[1580];
  assign N2777 = N2776 | data_masked[1708];
  assign N2776 = N2775 | data_masked[1836];
  assign N2775 = N2774 | data_masked[1964];
  assign N2774 = N2773 | data_masked[2092];
  assign N2773 = N2772 | data_masked[2220];
  assign N2772 = N2771 | data_masked[2348];
  assign N2771 = N2770 | data_masked[2476];
  assign N2770 = N2769 | data_masked[2604];
  assign N2769 = N2768 | data_masked[2732];
  assign N2768 = N2767 | data_masked[2860];
  assign N2767 = N2766 | data_masked[2988];
  assign N2766 = N2765 | data_masked[3116];
  assign N2765 = N2764 | data_masked[3244];
  assign N2764 = N2763 | data_masked[3372];
  assign N2763 = N2762 | data_masked[3500];
  assign N2762 = N2761 | data_masked[3628];
  assign N2761 = N2760 | data_masked[3756];
  assign N2760 = N2759 | data_masked[3884];
  assign N2759 = N2758 | data_masked[4012];
  assign N2758 = N2757 | data_masked[4140];
  assign N2757 = N2756 | data_masked[4268];
  assign N2756 = N2755 | data_masked[4396];
  assign N2755 = N2754 | data_masked[4524];
  assign N2754 = N2753 | data_masked[4652];
  assign N2753 = N2752 | data_masked[4780];
  assign N2752 = N2751 | data_masked[4908];
  assign N2751 = N2750 | data_masked[5036];
  assign N2750 = N2749 | data_masked[5164];
  assign N2749 = N2748 | data_masked[5292];
  assign N2748 = N2747 | data_masked[5420];
  assign N2747 = N2746 | data_masked[5548];
  assign N2746 = N2745 | data_masked[5676];
  assign N2745 = N2744 | data_masked[5804];
  assign N2744 = N2743 | data_masked[5932];
  assign N2743 = N2742 | data_masked[6060];
  assign N2742 = N2741 | data_masked[6188];
  assign N2741 = N2740 | data_masked[6316];
  assign N2740 = N2739 | data_masked[6444];
  assign N2739 = N2738 | data_masked[6572];
  assign N2738 = N2737 | data_masked[6700];
  assign N2737 = N2736 | data_masked[6828];
  assign N2736 = N2735 | data_masked[6956];
  assign N2735 = N2734 | data_masked[7084];
  assign N2734 = N2733 | data_masked[7212];
  assign N2733 = N2732 | data_masked[7340];
  assign N2732 = N2731 | data_masked[7468];
  assign N2731 = N2730 | data_masked[7596];
  assign N2730 = N2729 | data_masked[7724];
  assign N2729 = N2728 | data_masked[7852];
  assign N2728 = data_masked[8108] | data_masked[7980];
  assign data_o[45] = N2851 | data_masked[45];
  assign N2851 = N2850 | data_masked[173];
  assign N2850 = N2849 | data_masked[301];
  assign N2849 = N2848 | data_masked[429];
  assign N2848 = N2847 | data_masked[557];
  assign N2847 = N2846 | data_masked[685];
  assign N2846 = N2845 | data_masked[813];
  assign N2845 = N2844 | data_masked[941];
  assign N2844 = N2843 | data_masked[1069];
  assign N2843 = N2842 | data_masked[1197];
  assign N2842 = N2841 | data_masked[1325];
  assign N2841 = N2840 | data_masked[1453];
  assign N2840 = N2839 | data_masked[1581];
  assign N2839 = N2838 | data_masked[1709];
  assign N2838 = N2837 | data_masked[1837];
  assign N2837 = N2836 | data_masked[1965];
  assign N2836 = N2835 | data_masked[2093];
  assign N2835 = N2834 | data_masked[2221];
  assign N2834 = N2833 | data_masked[2349];
  assign N2833 = N2832 | data_masked[2477];
  assign N2832 = N2831 | data_masked[2605];
  assign N2831 = N2830 | data_masked[2733];
  assign N2830 = N2829 | data_masked[2861];
  assign N2829 = N2828 | data_masked[2989];
  assign N2828 = N2827 | data_masked[3117];
  assign N2827 = N2826 | data_masked[3245];
  assign N2826 = N2825 | data_masked[3373];
  assign N2825 = N2824 | data_masked[3501];
  assign N2824 = N2823 | data_masked[3629];
  assign N2823 = N2822 | data_masked[3757];
  assign N2822 = N2821 | data_masked[3885];
  assign N2821 = N2820 | data_masked[4013];
  assign N2820 = N2819 | data_masked[4141];
  assign N2819 = N2818 | data_masked[4269];
  assign N2818 = N2817 | data_masked[4397];
  assign N2817 = N2816 | data_masked[4525];
  assign N2816 = N2815 | data_masked[4653];
  assign N2815 = N2814 | data_masked[4781];
  assign N2814 = N2813 | data_masked[4909];
  assign N2813 = N2812 | data_masked[5037];
  assign N2812 = N2811 | data_masked[5165];
  assign N2811 = N2810 | data_masked[5293];
  assign N2810 = N2809 | data_masked[5421];
  assign N2809 = N2808 | data_masked[5549];
  assign N2808 = N2807 | data_masked[5677];
  assign N2807 = N2806 | data_masked[5805];
  assign N2806 = N2805 | data_masked[5933];
  assign N2805 = N2804 | data_masked[6061];
  assign N2804 = N2803 | data_masked[6189];
  assign N2803 = N2802 | data_masked[6317];
  assign N2802 = N2801 | data_masked[6445];
  assign N2801 = N2800 | data_masked[6573];
  assign N2800 = N2799 | data_masked[6701];
  assign N2799 = N2798 | data_masked[6829];
  assign N2798 = N2797 | data_masked[6957];
  assign N2797 = N2796 | data_masked[7085];
  assign N2796 = N2795 | data_masked[7213];
  assign N2795 = N2794 | data_masked[7341];
  assign N2794 = N2793 | data_masked[7469];
  assign N2793 = N2792 | data_masked[7597];
  assign N2792 = N2791 | data_masked[7725];
  assign N2791 = N2790 | data_masked[7853];
  assign N2790 = data_masked[8109] | data_masked[7981];
  assign data_o[46] = N2913 | data_masked[46];
  assign N2913 = N2912 | data_masked[174];
  assign N2912 = N2911 | data_masked[302];
  assign N2911 = N2910 | data_masked[430];
  assign N2910 = N2909 | data_masked[558];
  assign N2909 = N2908 | data_masked[686];
  assign N2908 = N2907 | data_masked[814];
  assign N2907 = N2906 | data_masked[942];
  assign N2906 = N2905 | data_masked[1070];
  assign N2905 = N2904 | data_masked[1198];
  assign N2904 = N2903 | data_masked[1326];
  assign N2903 = N2902 | data_masked[1454];
  assign N2902 = N2901 | data_masked[1582];
  assign N2901 = N2900 | data_masked[1710];
  assign N2900 = N2899 | data_masked[1838];
  assign N2899 = N2898 | data_masked[1966];
  assign N2898 = N2897 | data_masked[2094];
  assign N2897 = N2896 | data_masked[2222];
  assign N2896 = N2895 | data_masked[2350];
  assign N2895 = N2894 | data_masked[2478];
  assign N2894 = N2893 | data_masked[2606];
  assign N2893 = N2892 | data_masked[2734];
  assign N2892 = N2891 | data_masked[2862];
  assign N2891 = N2890 | data_masked[2990];
  assign N2890 = N2889 | data_masked[3118];
  assign N2889 = N2888 | data_masked[3246];
  assign N2888 = N2887 | data_masked[3374];
  assign N2887 = N2886 | data_masked[3502];
  assign N2886 = N2885 | data_masked[3630];
  assign N2885 = N2884 | data_masked[3758];
  assign N2884 = N2883 | data_masked[3886];
  assign N2883 = N2882 | data_masked[4014];
  assign N2882 = N2881 | data_masked[4142];
  assign N2881 = N2880 | data_masked[4270];
  assign N2880 = N2879 | data_masked[4398];
  assign N2879 = N2878 | data_masked[4526];
  assign N2878 = N2877 | data_masked[4654];
  assign N2877 = N2876 | data_masked[4782];
  assign N2876 = N2875 | data_masked[4910];
  assign N2875 = N2874 | data_masked[5038];
  assign N2874 = N2873 | data_masked[5166];
  assign N2873 = N2872 | data_masked[5294];
  assign N2872 = N2871 | data_masked[5422];
  assign N2871 = N2870 | data_masked[5550];
  assign N2870 = N2869 | data_masked[5678];
  assign N2869 = N2868 | data_masked[5806];
  assign N2868 = N2867 | data_masked[5934];
  assign N2867 = N2866 | data_masked[6062];
  assign N2866 = N2865 | data_masked[6190];
  assign N2865 = N2864 | data_masked[6318];
  assign N2864 = N2863 | data_masked[6446];
  assign N2863 = N2862 | data_masked[6574];
  assign N2862 = N2861 | data_masked[6702];
  assign N2861 = N2860 | data_masked[6830];
  assign N2860 = N2859 | data_masked[6958];
  assign N2859 = N2858 | data_masked[7086];
  assign N2858 = N2857 | data_masked[7214];
  assign N2857 = N2856 | data_masked[7342];
  assign N2856 = N2855 | data_masked[7470];
  assign N2855 = N2854 | data_masked[7598];
  assign N2854 = N2853 | data_masked[7726];
  assign N2853 = N2852 | data_masked[7854];
  assign N2852 = data_masked[8110] | data_masked[7982];
  assign data_o[47] = N2975 | data_masked[47];
  assign N2975 = N2974 | data_masked[175];
  assign N2974 = N2973 | data_masked[303];
  assign N2973 = N2972 | data_masked[431];
  assign N2972 = N2971 | data_masked[559];
  assign N2971 = N2970 | data_masked[687];
  assign N2970 = N2969 | data_masked[815];
  assign N2969 = N2968 | data_masked[943];
  assign N2968 = N2967 | data_masked[1071];
  assign N2967 = N2966 | data_masked[1199];
  assign N2966 = N2965 | data_masked[1327];
  assign N2965 = N2964 | data_masked[1455];
  assign N2964 = N2963 | data_masked[1583];
  assign N2963 = N2962 | data_masked[1711];
  assign N2962 = N2961 | data_masked[1839];
  assign N2961 = N2960 | data_masked[1967];
  assign N2960 = N2959 | data_masked[2095];
  assign N2959 = N2958 | data_masked[2223];
  assign N2958 = N2957 | data_masked[2351];
  assign N2957 = N2956 | data_masked[2479];
  assign N2956 = N2955 | data_masked[2607];
  assign N2955 = N2954 | data_masked[2735];
  assign N2954 = N2953 | data_masked[2863];
  assign N2953 = N2952 | data_masked[2991];
  assign N2952 = N2951 | data_masked[3119];
  assign N2951 = N2950 | data_masked[3247];
  assign N2950 = N2949 | data_masked[3375];
  assign N2949 = N2948 | data_masked[3503];
  assign N2948 = N2947 | data_masked[3631];
  assign N2947 = N2946 | data_masked[3759];
  assign N2946 = N2945 | data_masked[3887];
  assign N2945 = N2944 | data_masked[4015];
  assign N2944 = N2943 | data_masked[4143];
  assign N2943 = N2942 | data_masked[4271];
  assign N2942 = N2941 | data_masked[4399];
  assign N2941 = N2940 | data_masked[4527];
  assign N2940 = N2939 | data_masked[4655];
  assign N2939 = N2938 | data_masked[4783];
  assign N2938 = N2937 | data_masked[4911];
  assign N2937 = N2936 | data_masked[5039];
  assign N2936 = N2935 | data_masked[5167];
  assign N2935 = N2934 | data_masked[5295];
  assign N2934 = N2933 | data_masked[5423];
  assign N2933 = N2932 | data_masked[5551];
  assign N2932 = N2931 | data_masked[5679];
  assign N2931 = N2930 | data_masked[5807];
  assign N2930 = N2929 | data_masked[5935];
  assign N2929 = N2928 | data_masked[6063];
  assign N2928 = N2927 | data_masked[6191];
  assign N2927 = N2926 | data_masked[6319];
  assign N2926 = N2925 | data_masked[6447];
  assign N2925 = N2924 | data_masked[6575];
  assign N2924 = N2923 | data_masked[6703];
  assign N2923 = N2922 | data_masked[6831];
  assign N2922 = N2921 | data_masked[6959];
  assign N2921 = N2920 | data_masked[7087];
  assign N2920 = N2919 | data_masked[7215];
  assign N2919 = N2918 | data_masked[7343];
  assign N2918 = N2917 | data_masked[7471];
  assign N2917 = N2916 | data_masked[7599];
  assign N2916 = N2915 | data_masked[7727];
  assign N2915 = N2914 | data_masked[7855];
  assign N2914 = data_masked[8111] | data_masked[7983];
  assign data_o[48] = N3037 | data_masked[48];
  assign N3037 = N3036 | data_masked[176];
  assign N3036 = N3035 | data_masked[304];
  assign N3035 = N3034 | data_masked[432];
  assign N3034 = N3033 | data_masked[560];
  assign N3033 = N3032 | data_masked[688];
  assign N3032 = N3031 | data_masked[816];
  assign N3031 = N3030 | data_masked[944];
  assign N3030 = N3029 | data_masked[1072];
  assign N3029 = N3028 | data_masked[1200];
  assign N3028 = N3027 | data_masked[1328];
  assign N3027 = N3026 | data_masked[1456];
  assign N3026 = N3025 | data_masked[1584];
  assign N3025 = N3024 | data_masked[1712];
  assign N3024 = N3023 | data_masked[1840];
  assign N3023 = N3022 | data_masked[1968];
  assign N3022 = N3021 | data_masked[2096];
  assign N3021 = N3020 | data_masked[2224];
  assign N3020 = N3019 | data_masked[2352];
  assign N3019 = N3018 | data_masked[2480];
  assign N3018 = N3017 | data_masked[2608];
  assign N3017 = N3016 | data_masked[2736];
  assign N3016 = N3015 | data_masked[2864];
  assign N3015 = N3014 | data_masked[2992];
  assign N3014 = N3013 | data_masked[3120];
  assign N3013 = N3012 | data_masked[3248];
  assign N3012 = N3011 | data_masked[3376];
  assign N3011 = N3010 | data_masked[3504];
  assign N3010 = N3009 | data_masked[3632];
  assign N3009 = N3008 | data_masked[3760];
  assign N3008 = N3007 | data_masked[3888];
  assign N3007 = N3006 | data_masked[4016];
  assign N3006 = N3005 | data_masked[4144];
  assign N3005 = N3004 | data_masked[4272];
  assign N3004 = N3003 | data_masked[4400];
  assign N3003 = N3002 | data_masked[4528];
  assign N3002 = N3001 | data_masked[4656];
  assign N3001 = N3000 | data_masked[4784];
  assign N3000 = N2999 | data_masked[4912];
  assign N2999 = N2998 | data_masked[5040];
  assign N2998 = N2997 | data_masked[5168];
  assign N2997 = N2996 | data_masked[5296];
  assign N2996 = N2995 | data_masked[5424];
  assign N2995 = N2994 | data_masked[5552];
  assign N2994 = N2993 | data_masked[5680];
  assign N2993 = N2992 | data_masked[5808];
  assign N2992 = N2991 | data_masked[5936];
  assign N2991 = N2990 | data_masked[6064];
  assign N2990 = N2989 | data_masked[6192];
  assign N2989 = N2988 | data_masked[6320];
  assign N2988 = N2987 | data_masked[6448];
  assign N2987 = N2986 | data_masked[6576];
  assign N2986 = N2985 | data_masked[6704];
  assign N2985 = N2984 | data_masked[6832];
  assign N2984 = N2983 | data_masked[6960];
  assign N2983 = N2982 | data_masked[7088];
  assign N2982 = N2981 | data_masked[7216];
  assign N2981 = N2980 | data_masked[7344];
  assign N2980 = N2979 | data_masked[7472];
  assign N2979 = N2978 | data_masked[7600];
  assign N2978 = N2977 | data_masked[7728];
  assign N2977 = N2976 | data_masked[7856];
  assign N2976 = data_masked[8112] | data_masked[7984];
  assign data_o[49] = N3099 | data_masked[49];
  assign N3099 = N3098 | data_masked[177];
  assign N3098 = N3097 | data_masked[305];
  assign N3097 = N3096 | data_masked[433];
  assign N3096 = N3095 | data_masked[561];
  assign N3095 = N3094 | data_masked[689];
  assign N3094 = N3093 | data_masked[817];
  assign N3093 = N3092 | data_masked[945];
  assign N3092 = N3091 | data_masked[1073];
  assign N3091 = N3090 | data_masked[1201];
  assign N3090 = N3089 | data_masked[1329];
  assign N3089 = N3088 | data_masked[1457];
  assign N3088 = N3087 | data_masked[1585];
  assign N3087 = N3086 | data_masked[1713];
  assign N3086 = N3085 | data_masked[1841];
  assign N3085 = N3084 | data_masked[1969];
  assign N3084 = N3083 | data_masked[2097];
  assign N3083 = N3082 | data_masked[2225];
  assign N3082 = N3081 | data_masked[2353];
  assign N3081 = N3080 | data_masked[2481];
  assign N3080 = N3079 | data_masked[2609];
  assign N3079 = N3078 | data_masked[2737];
  assign N3078 = N3077 | data_masked[2865];
  assign N3077 = N3076 | data_masked[2993];
  assign N3076 = N3075 | data_masked[3121];
  assign N3075 = N3074 | data_masked[3249];
  assign N3074 = N3073 | data_masked[3377];
  assign N3073 = N3072 | data_masked[3505];
  assign N3072 = N3071 | data_masked[3633];
  assign N3071 = N3070 | data_masked[3761];
  assign N3070 = N3069 | data_masked[3889];
  assign N3069 = N3068 | data_masked[4017];
  assign N3068 = N3067 | data_masked[4145];
  assign N3067 = N3066 | data_masked[4273];
  assign N3066 = N3065 | data_masked[4401];
  assign N3065 = N3064 | data_masked[4529];
  assign N3064 = N3063 | data_masked[4657];
  assign N3063 = N3062 | data_masked[4785];
  assign N3062 = N3061 | data_masked[4913];
  assign N3061 = N3060 | data_masked[5041];
  assign N3060 = N3059 | data_masked[5169];
  assign N3059 = N3058 | data_masked[5297];
  assign N3058 = N3057 | data_masked[5425];
  assign N3057 = N3056 | data_masked[5553];
  assign N3056 = N3055 | data_masked[5681];
  assign N3055 = N3054 | data_masked[5809];
  assign N3054 = N3053 | data_masked[5937];
  assign N3053 = N3052 | data_masked[6065];
  assign N3052 = N3051 | data_masked[6193];
  assign N3051 = N3050 | data_masked[6321];
  assign N3050 = N3049 | data_masked[6449];
  assign N3049 = N3048 | data_masked[6577];
  assign N3048 = N3047 | data_masked[6705];
  assign N3047 = N3046 | data_masked[6833];
  assign N3046 = N3045 | data_masked[6961];
  assign N3045 = N3044 | data_masked[7089];
  assign N3044 = N3043 | data_masked[7217];
  assign N3043 = N3042 | data_masked[7345];
  assign N3042 = N3041 | data_masked[7473];
  assign N3041 = N3040 | data_masked[7601];
  assign N3040 = N3039 | data_masked[7729];
  assign N3039 = N3038 | data_masked[7857];
  assign N3038 = data_masked[8113] | data_masked[7985];
  assign data_o[50] = N3161 | data_masked[50];
  assign N3161 = N3160 | data_masked[178];
  assign N3160 = N3159 | data_masked[306];
  assign N3159 = N3158 | data_masked[434];
  assign N3158 = N3157 | data_masked[562];
  assign N3157 = N3156 | data_masked[690];
  assign N3156 = N3155 | data_masked[818];
  assign N3155 = N3154 | data_masked[946];
  assign N3154 = N3153 | data_masked[1074];
  assign N3153 = N3152 | data_masked[1202];
  assign N3152 = N3151 | data_masked[1330];
  assign N3151 = N3150 | data_masked[1458];
  assign N3150 = N3149 | data_masked[1586];
  assign N3149 = N3148 | data_masked[1714];
  assign N3148 = N3147 | data_masked[1842];
  assign N3147 = N3146 | data_masked[1970];
  assign N3146 = N3145 | data_masked[2098];
  assign N3145 = N3144 | data_masked[2226];
  assign N3144 = N3143 | data_masked[2354];
  assign N3143 = N3142 | data_masked[2482];
  assign N3142 = N3141 | data_masked[2610];
  assign N3141 = N3140 | data_masked[2738];
  assign N3140 = N3139 | data_masked[2866];
  assign N3139 = N3138 | data_masked[2994];
  assign N3138 = N3137 | data_masked[3122];
  assign N3137 = N3136 | data_masked[3250];
  assign N3136 = N3135 | data_masked[3378];
  assign N3135 = N3134 | data_masked[3506];
  assign N3134 = N3133 | data_masked[3634];
  assign N3133 = N3132 | data_masked[3762];
  assign N3132 = N3131 | data_masked[3890];
  assign N3131 = N3130 | data_masked[4018];
  assign N3130 = N3129 | data_masked[4146];
  assign N3129 = N3128 | data_masked[4274];
  assign N3128 = N3127 | data_masked[4402];
  assign N3127 = N3126 | data_masked[4530];
  assign N3126 = N3125 | data_masked[4658];
  assign N3125 = N3124 | data_masked[4786];
  assign N3124 = N3123 | data_masked[4914];
  assign N3123 = N3122 | data_masked[5042];
  assign N3122 = N3121 | data_masked[5170];
  assign N3121 = N3120 | data_masked[5298];
  assign N3120 = N3119 | data_masked[5426];
  assign N3119 = N3118 | data_masked[5554];
  assign N3118 = N3117 | data_masked[5682];
  assign N3117 = N3116 | data_masked[5810];
  assign N3116 = N3115 | data_masked[5938];
  assign N3115 = N3114 | data_masked[6066];
  assign N3114 = N3113 | data_masked[6194];
  assign N3113 = N3112 | data_masked[6322];
  assign N3112 = N3111 | data_masked[6450];
  assign N3111 = N3110 | data_masked[6578];
  assign N3110 = N3109 | data_masked[6706];
  assign N3109 = N3108 | data_masked[6834];
  assign N3108 = N3107 | data_masked[6962];
  assign N3107 = N3106 | data_masked[7090];
  assign N3106 = N3105 | data_masked[7218];
  assign N3105 = N3104 | data_masked[7346];
  assign N3104 = N3103 | data_masked[7474];
  assign N3103 = N3102 | data_masked[7602];
  assign N3102 = N3101 | data_masked[7730];
  assign N3101 = N3100 | data_masked[7858];
  assign N3100 = data_masked[8114] | data_masked[7986];
  assign data_o[51] = N3223 | data_masked[51];
  assign N3223 = N3222 | data_masked[179];
  assign N3222 = N3221 | data_masked[307];
  assign N3221 = N3220 | data_masked[435];
  assign N3220 = N3219 | data_masked[563];
  assign N3219 = N3218 | data_masked[691];
  assign N3218 = N3217 | data_masked[819];
  assign N3217 = N3216 | data_masked[947];
  assign N3216 = N3215 | data_masked[1075];
  assign N3215 = N3214 | data_masked[1203];
  assign N3214 = N3213 | data_masked[1331];
  assign N3213 = N3212 | data_masked[1459];
  assign N3212 = N3211 | data_masked[1587];
  assign N3211 = N3210 | data_masked[1715];
  assign N3210 = N3209 | data_masked[1843];
  assign N3209 = N3208 | data_masked[1971];
  assign N3208 = N3207 | data_masked[2099];
  assign N3207 = N3206 | data_masked[2227];
  assign N3206 = N3205 | data_masked[2355];
  assign N3205 = N3204 | data_masked[2483];
  assign N3204 = N3203 | data_masked[2611];
  assign N3203 = N3202 | data_masked[2739];
  assign N3202 = N3201 | data_masked[2867];
  assign N3201 = N3200 | data_masked[2995];
  assign N3200 = N3199 | data_masked[3123];
  assign N3199 = N3198 | data_masked[3251];
  assign N3198 = N3197 | data_masked[3379];
  assign N3197 = N3196 | data_masked[3507];
  assign N3196 = N3195 | data_masked[3635];
  assign N3195 = N3194 | data_masked[3763];
  assign N3194 = N3193 | data_masked[3891];
  assign N3193 = N3192 | data_masked[4019];
  assign N3192 = N3191 | data_masked[4147];
  assign N3191 = N3190 | data_masked[4275];
  assign N3190 = N3189 | data_masked[4403];
  assign N3189 = N3188 | data_masked[4531];
  assign N3188 = N3187 | data_masked[4659];
  assign N3187 = N3186 | data_masked[4787];
  assign N3186 = N3185 | data_masked[4915];
  assign N3185 = N3184 | data_masked[5043];
  assign N3184 = N3183 | data_masked[5171];
  assign N3183 = N3182 | data_masked[5299];
  assign N3182 = N3181 | data_masked[5427];
  assign N3181 = N3180 | data_masked[5555];
  assign N3180 = N3179 | data_masked[5683];
  assign N3179 = N3178 | data_masked[5811];
  assign N3178 = N3177 | data_masked[5939];
  assign N3177 = N3176 | data_masked[6067];
  assign N3176 = N3175 | data_masked[6195];
  assign N3175 = N3174 | data_masked[6323];
  assign N3174 = N3173 | data_masked[6451];
  assign N3173 = N3172 | data_masked[6579];
  assign N3172 = N3171 | data_masked[6707];
  assign N3171 = N3170 | data_masked[6835];
  assign N3170 = N3169 | data_masked[6963];
  assign N3169 = N3168 | data_masked[7091];
  assign N3168 = N3167 | data_masked[7219];
  assign N3167 = N3166 | data_masked[7347];
  assign N3166 = N3165 | data_masked[7475];
  assign N3165 = N3164 | data_masked[7603];
  assign N3164 = N3163 | data_masked[7731];
  assign N3163 = N3162 | data_masked[7859];
  assign N3162 = data_masked[8115] | data_masked[7987];
  assign data_o[52] = N3285 | data_masked[52];
  assign N3285 = N3284 | data_masked[180];
  assign N3284 = N3283 | data_masked[308];
  assign N3283 = N3282 | data_masked[436];
  assign N3282 = N3281 | data_masked[564];
  assign N3281 = N3280 | data_masked[692];
  assign N3280 = N3279 | data_masked[820];
  assign N3279 = N3278 | data_masked[948];
  assign N3278 = N3277 | data_masked[1076];
  assign N3277 = N3276 | data_masked[1204];
  assign N3276 = N3275 | data_masked[1332];
  assign N3275 = N3274 | data_masked[1460];
  assign N3274 = N3273 | data_masked[1588];
  assign N3273 = N3272 | data_masked[1716];
  assign N3272 = N3271 | data_masked[1844];
  assign N3271 = N3270 | data_masked[1972];
  assign N3270 = N3269 | data_masked[2100];
  assign N3269 = N3268 | data_masked[2228];
  assign N3268 = N3267 | data_masked[2356];
  assign N3267 = N3266 | data_masked[2484];
  assign N3266 = N3265 | data_masked[2612];
  assign N3265 = N3264 | data_masked[2740];
  assign N3264 = N3263 | data_masked[2868];
  assign N3263 = N3262 | data_masked[2996];
  assign N3262 = N3261 | data_masked[3124];
  assign N3261 = N3260 | data_masked[3252];
  assign N3260 = N3259 | data_masked[3380];
  assign N3259 = N3258 | data_masked[3508];
  assign N3258 = N3257 | data_masked[3636];
  assign N3257 = N3256 | data_masked[3764];
  assign N3256 = N3255 | data_masked[3892];
  assign N3255 = N3254 | data_masked[4020];
  assign N3254 = N3253 | data_masked[4148];
  assign N3253 = N3252 | data_masked[4276];
  assign N3252 = N3251 | data_masked[4404];
  assign N3251 = N3250 | data_masked[4532];
  assign N3250 = N3249 | data_masked[4660];
  assign N3249 = N3248 | data_masked[4788];
  assign N3248 = N3247 | data_masked[4916];
  assign N3247 = N3246 | data_masked[5044];
  assign N3246 = N3245 | data_masked[5172];
  assign N3245 = N3244 | data_masked[5300];
  assign N3244 = N3243 | data_masked[5428];
  assign N3243 = N3242 | data_masked[5556];
  assign N3242 = N3241 | data_masked[5684];
  assign N3241 = N3240 | data_masked[5812];
  assign N3240 = N3239 | data_masked[5940];
  assign N3239 = N3238 | data_masked[6068];
  assign N3238 = N3237 | data_masked[6196];
  assign N3237 = N3236 | data_masked[6324];
  assign N3236 = N3235 | data_masked[6452];
  assign N3235 = N3234 | data_masked[6580];
  assign N3234 = N3233 | data_masked[6708];
  assign N3233 = N3232 | data_masked[6836];
  assign N3232 = N3231 | data_masked[6964];
  assign N3231 = N3230 | data_masked[7092];
  assign N3230 = N3229 | data_masked[7220];
  assign N3229 = N3228 | data_masked[7348];
  assign N3228 = N3227 | data_masked[7476];
  assign N3227 = N3226 | data_masked[7604];
  assign N3226 = N3225 | data_masked[7732];
  assign N3225 = N3224 | data_masked[7860];
  assign N3224 = data_masked[8116] | data_masked[7988];
  assign data_o[53] = N3347 | data_masked[53];
  assign N3347 = N3346 | data_masked[181];
  assign N3346 = N3345 | data_masked[309];
  assign N3345 = N3344 | data_masked[437];
  assign N3344 = N3343 | data_masked[565];
  assign N3343 = N3342 | data_masked[693];
  assign N3342 = N3341 | data_masked[821];
  assign N3341 = N3340 | data_masked[949];
  assign N3340 = N3339 | data_masked[1077];
  assign N3339 = N3338 | data_masked[1205];
  assign N3338 = N3337 | data_masked[1333];
  assign N3337 = N3336 | data_masked[1461];
  assign N3336 = N3335 | data_masked[1589];
  assign N3335 = N3334 | data_masked[1717];
  assign N3334 = N3333 | data_masked[1845];
  assign N3333 = N3332 | data_masked[1973];
  assign N3332 = N3331 | data_masked[2101];
  assign N3331 = N3330 | data_masked[2229];
  assign N3330 = N3329 | data_masked[2357];
  assign N3329 = N3328 | data_masked[2485];
  assign N3328 = N3327 | data_masked[2613];
  assign N3327 = N3326 | data_masked[2741];
  assign N3326 = N3325 | data_masked[2869];
  assign N3325 = N3324 | data_masked[2997];
  assign N3324 = N3323 | data_masked[3125];
  assign N3323 = N3322 | data_masked[3253];
  assign N3322 = N3321 | data_masked[3381];
  assign N3321 = N3320 | data_masked[3509];
  assign N3320 = N3319 | data_masked[3637];
  assign N3319 = N3318 | data_masked[3765];
  assign N3318 = N3317 | data_masked[3893];
  assign N3317 = N3316 | data_masked[4021];
  assign N3316 = N3315 | data_masked[4149];
  assign N3315 = N3314 | data_masked[4277];
  assign N3314 = N3313 | data_masked[4405];
  assign N3313 = N3312 | data_masked[4533];
  assign N3312 = N3311 | data_masked[4661];
  assign N3311 = N3310 | data_masked[4789];
  assign N3310 = N3309 | data_masked[4917];
  assign N3309 = N3308 | data_masked[5045];
  assign N3308 = N3307 | data_masked[5173];
  assign N3307 = N3306 | data_masked[5301];
  assign N3306 = N3305 | data_masked[5429];
  assign N3305 = N3304 | data_masked[5557];
  assign N3304 = N3303 | data_masked[5685];
  assign N3303 = N3302 | data_masked[5813];
  assign N3302 = N3301 | data_masked[5941];
  assign N3301 = N3300 | data_masked[6069];
  assign N3300 = N3299 | data_masked[6197];
  assign N3299 = N3298 | data_masked[6325];
  assign N3298 = N3297 | data_masked[6453];
  assign N3297 = N3296 | data_masked[6581];
  assign N3296 = N3295 | data_masked[6709];
  assign N3295 = N3294 | data_masked[6837];
  assign N3294 = N3293 | data_masked[6965];
  assign N3293 = N3292 | data_masked[7093];
  assign N3292 = N3291 | data_masked[7221];
  assign N3291 = N3290 | data_masked[7349];
  assign N3290 = N3289 | data_masked[7477];
  assign N3289 = N3288 | data_masked[7605];
  assign N3288 = N3287 | data_masked[7733];
  assign N3287 = N3286 | data_masked[7861];
  assign N3286 = data_masked[8117] | data_masked[7989];
  assign data_o[54] = N3409 | data_masked[54];
  assign N3409 = N3408 | data_masked[182];
  assign N3408 = N3407 | data_masked[310];
  assign N3407 = N3406 | data_masked[438];
  assign N3406 = N3405 | data_masked[566];
  assign N3405 = N3404 | data_masked[694];
  assign N3404 = N3403 | data_masked[822];
  assign N3403 = N3402 | data_masked[950];
  assign N3402 = N3401 | data_masked[1078];
  assign N3401 = N3400 | data_masked[1206];
  assign N3400 = N3399 | data_masked[1334];
  assign N3399 = N3398 | data_masked[1462];
  assign N3398 = N3397 | data_masked[1590];
  assign N3397 = N3396 | data_masked[1718];
  assign N3396 = N3395 | data_masked[1846];
  assign N3395 = N3394 | data_masked[1974];
  assign N3394 = N3393 | data_masked[2102];
  assign N3393 = N3392 | data_masked[2230];
  assign N3392 = N3391 | data_masked[2358];
  assign N3391 = N3390 | data_masked[2486];
  assign N3390 = N3389 | data_masked[2614];
  assign N3389 = N3388 | data_masked[2742];
  assign N3388 = N3387 | data_masked[2870];
  assign N3387 = N3386 | data_masked[2998];
  assign N3386 = N3385 | data_masked[3126];
  assign N3385 = N3384 | data_masked[3254];
  assign N3384 = N3383 | data_masked[3382];
  assign N3383 = N3382 | data_masked[3510];
  assign N3382 = N3381 | data_masked[3638];
  assign N3381 = N3380 | data_masked[3766];
  assign N3380 = N3379 | data_masked[3894];
  assign N3379 = N3378 | data_masked[4022];
  assign N3378 = N3377 | data_masked[4150];
  assign N3377 = N3376 | data_masked[4278];
  assign N3376 = N3375 | data_masked[4406];
  assign N3375 = N3374 | data_masked[4534];
  assign N3374 = N3373 | data_masked[4662];
  assign N3373 = N3372 | data_masked[4790];
  assign N3372 = N3371 | data_masked[4918];
  assign N3371 = N3370 | data_masked[5046];
  assign N3370 = N3369 | data_masked[5174];
  assign N3369 = N3368 | data_masked[5302];
  assign N3368 = N3367 | data_masked[5430];
  assign N3367 = N3366 | data_masked[5558];
  assign N3366 = N3365 | data_masked[5686];
  assign N3365 = N3364 | data_masked[5814];
  assign N3364 = N3363 | data_masked[5942];
  assign N3363 = N3362 | data_masked[6070];
  assign N3362 = N3361 | data_masked[6198];
  assign N3361 = N3360 | data_masked[6326];
  assign N3360 = N3359 | data_masked[6454];
  assign N3359 = N3358 | data_masked[6582];
  assign N3358 = N3357 | data_masked[6710];
  assign N3357 = N3356 | data_masked[6838];
  assign N3356 = N3355 | data_masked[6966];
  assign N3355 = N3354 | data_masked[7094];
  assign N3354 = N3353 | data_masked[7222];
  assign N3353 = N3352 | data_masked[7350];
  assign N3352 = N3351 | data_masked[7478];
  assign N3351 = N3350 | data_masked[7606];
  assign N3350 = N3349 | data_masked[7734];
  assign N3349 = N3348 | data_masked[7862];
  assign N3348 = data_masked[8118] | data_masked[7990];
  assign data_o[55] = N3471 | data_masked[55];
  assign N3471 = N3470 | data_masked[183];
  assign N3470 = N3469 | data_masked[311];
  assign N3469 = N3468 | data_masked[439];
  assign N3468 = N3467 | data_masked[567];
  assign N3467 = N3466 | data_masked[695];
  assign N3466 = N3465 | data_masked[823];
  assign N3465 = N3464 | data_masked[951];
  assign N3464 = N3463 | data_masked[1079];
  assign N3463 = N3462 | data_masked[1207];
  assign N3462 = N3461 | data_masked[1335];
  assign N3461 = N3460 | data_masked[1463];
  assign N3460 = N3459 | data_masked[1591];
  assign N3459 = N3458 | data_masked[1719];
  assign N3458 = N3457 | data_masked[1847];
  assign N3457 = N3456 | data_masked[1975];
  assign N3456 = N3455 | data_masked[2103];
  assign N3455 = N3454 | data_masked[2231];
  assign N3454 = N3453 | data_masked[2359];
  assign N3453 = N3452 | data_masked[2487];
  assign N3452 = N3451 | data_masked[2615];
  assign N3451 = N3450 | data_masked[2743];
  assign N3450 = N3449 | data_masked[2871];
  assign N3449 = N3448 | data_masked[2999];
  assign N3448 = N3447 | data_masked[3127];
  assign N3447 = N3446 | data_masked[3255];
  assign N3446 = N3445 | data_masked[3383];
  assign N3445 = N3444 | data_masked[3511];
  assign N3444 = N3443 | data_masked[3639];
  assign N3443 = N3442 | data_masked[3767];
  assign N3442 = N3441 | data_masked[3895];
  assign N3441 = N3440 | data_masked[4023];
  assign N3440 = N3439 | data_masked[4151];
  assign N3439 = N3438 | data_masked[4279];
  assign N3438 = N3437 | data_masked[4407];
  assign N3437 = N3436 | data_masked[4535];
  assign N3436 = N3435 | data_masked[4663];
  assign N3435 = N3434 | data_masked[4791];
  assign N3434 = N3433 | data_masked[4919];
  assign N3433 = N3432 | data_masked[5047];
  assign N3432 = N3431 | data_masked[5175];
  assign N3431 = N3430 | data_masked[5303];
  assign N3430 = N3429 | data_masked[5431];
  assign N3429 = N3428 | data_masked[5559];
  assign N3428 = N3427 | data_masked[5687];
  assign N3427 = N3426 | data_masked[5815];
  assign N3426 = N3425 | data_masked[5943];
  assign N3425 = N3424 | data_masked[6071];
  assign N3424 = N3423 | data_masked[6199];
  assign N3423 = N3422 | data_masked[6327];
  assign N3422 = N3421 | data_masked[6455];
  assign N3421 = N3420 | data_masked[6583];
  assign N3420 = N3419 | data_masked[6711];
  assign N3419 = N3418 | data_masked[6839];
  assign N3418 = N3417 | data_masked[6967];
  assign N3417 = N3416 | data_masked[7095];
  assign N3416 = N3415 | data_masked[7223];
  assign N3415 = N3414 | data_masked[7351];
  assign N3414 = N3413 | data_masked[7479];
  assign N3413 = N3412 | data_masked[7607];
  assign N3412 = N3411 | data_masked[7735];
  assign N3411 = N3410 | data_masked[7863];
  assign N3410 = data_masked[8119] | data_masked[7991];
  assign data_o[56] = N3533 | data_masked[56];
  assign N3533 = N3532 | data_masked[184];
  assign N3532 = N3531 | data_masked[312];
  assign N3531 = N3530 | data_masked[440];
  assign N3530 = N3529 | data_masked[568];
  assign N3529 = N3528 | data_masked[696];
  assign N3528 = N3527 | data_masked[824];
  assign N3527 = N3526 | data_masked[952];
  assign N3526 = N3525 | data_masked[1080];
  assign N3525 = N3524 | data_masked[1208];
  assign N3524 = N3523 | data_masked[1336];
  assign N3523 = N3522 | data_masked[1464];
  assign N3522 = N3521 | data_masked[1592];
  assign N3521 = N3520 | data_masked[1720];
  assign N3520 = N3519 | data_masked[1848];
  assign N3519 = N3518 | data_masked[1976];
  assign N3518 = N3517 | data_masked[2104];
  assign N3517 = N3516 | data_masked[2232];
  assign N3516 = N3515 | data_masked[2360];
  assign N3515 = N3514 | data_masked[2488];
  assign N3514 = N3513 | data_masked[2616];
  assign N3513 = N3512 | data_masked[2744];
  assign N3512 = N3511 | data_masked[2872];
  assign N3511 = N3510 | data_masked[3000];
  assign N3510 = N3509 | data_masked[3128];
  assign N3509 = N3508 | data_masked[3256];
  assign N3508 = N3507 | data_masked[3384];
  assign N3507 = N3506 | data_masked[3512];
  assign N3506 = N3505 | data_masked[3640];
  assign N3505 = N3504 | data_masked[3768];
  assign N3504 = N3503 | data_masked[3896];
  assign N3503 = N3502 | data_masked[4024];
  assign N3502 = N3501 | data_masked[4152];
  assign N3501 = N3500 | data_masked[4280];
  assign N3500 = N3499 | data_masked[4408];
  assign N3499 = N3498 | data_masked[4536];
  assign N3498 = N3497 | data_masked[4664];
  assign N3497 = N3496 | data_masked[4792];
  assign N3496 = N3495 | data_masked[4920];
  assign N3495 = N3494 | data_masked[5048];
  assign N3494 = N3493 | data_masked[5176];
  assign N3493 = N3492 | data_masked[5304];
  assign N3492 = N3491 | data_masked[5432];
  assign N3491 = N3490 | data_masked[5560];
  assign N3490 = N3489 | data_masked[5688];
  assign N3489 = N3488 | data_masked[5816];
  assign N3488 = N3487 | data_masked[5944];
  assign N3487 = N3486 | data_masked[6072];
  assign N3486 = N3485 | data_masked[6200];
  assign N3485 = N3484 | data_masked[6328];
  assign N3484 = N3483 | data_masked[6456];
  assign N3483 = N3482 | data_masked[6584];
  assign N3482 = N3481 | data_masked[6712];
  assign N3481 = N3480 | data_masked[6840];
  assign N3480 = N3479 | data_masked[6968];
  assign N3479 = N3478 | data_masked[7096];
  assign N3478 = N3477 | data_masked[7224];
  assign N3477 = N3476 | data_masked[7352];
  assign N3476 = N3475 | data_masked[7480];
  assign N3475 = N3474 | data_masked[7608];
  assign N3474 = N3473 | data_masked[7736];
  assign N3473 = N3472 | data_masked[7864];
  assign N3472 = data_masked[8120] | data_masked[7992];
  assign data_o[57] = N3595 | data_masked[57];
  assign N3595 = N3594 | data_masked[185];
  assign N3594 = N3593 | data_masked[313];
  assign N3593 = N3592 | data_masked[441];
  assign N3592 = N3591 | data_masked[569];
  assign N3591 = N3590 | data_masked[697];
  assign N3590 = N3589 | data_masked[825];
  assign N3589 = N3588 | data_masked[953];
  assign N3588 = N3587 | data_masked[1081];
  assign N3587 = N3586 | data_masked[1209];
  assign N3586 = N3585 | data_masked[1337];
  assign N3585 = N3584 | data_masked[1465];
  assign N3584 = N3583 | data_masked[1593];
  assign N3583 = N3582 | data_masked[1721];
  assign N3582 = N3581 | data_masked[1849];
  assign N3581 = N3580 | data_masked[1977];
  assign N3580 = N3579 | data_masked[2105];
  assign N3579 = N3578 | data_masked[2233];
  assign N3578 = N3577 | data_masked[2361];
  assign N3577 = N3576 | data_masked[2489];
  assign N3576 = N3575 | data_masked[2617];
  assign N3575 = N3574 | data_masked[2745];
  assign N3574 = N3573 | data_masked[2873];
  assign N3573 = N3572 | data_masked[3001];
  assign N3572 = N3571 | data_masked[3129];
  assign N3571 = N3570 | data_masked[3257];
  assign N3570 = N3569 | data_masked[3385];
  assign N3569 = N3568 | data_masked[3513];
  assign N3568 = N3567 | data_masked[3641];
  assign N3567 = N3566 | data_masked[3769];
  assign N3566 = N3565 | data_masked[3897];
  assign N3565 = N3564 | data_masked[4025];
  assign N3564 = N3563 | data_masked[4153];
  assign N3563 = N3562 | data_masked[4281];
  assign N3562 = N3561 | data_masked[4409];
  assign N3561 = N3560 | data_masked[4537];
  assign N3560 = N3559 | data_masked[4665];
  assign N3559 = N3558 | data_masked[4793];
  assign N3558 = N3557 | data_masked[4921];
  assign N3557 = N3556 | data_masked[5049];
  assign N3556 = N3555 | data_masked[5177];
  assign N3555 = N3554 | data_masked[5305];
  assign N3554 = N3553 | data_masked[5433];
  assign N3553 = N3552 | data_masked[5561];
  assign N3552 = N3551 | data_masked[5689];
  assign N3551 = N3550 | data_masked[5817];
  assign N3550 = N3549 | data_masked[5945];
  assign N3549 = N3548 | data_masked[6073];
  assign N3548 = N3547 | data_masked[6201];
  assign N3547 = N3546 | data_masked[6329];
  assign N3546 = N3545 | data_masked[6457];
  assign N3545 = N3544 | data_masked[6585];
  assign N3544 = N3543 | data_masked[6713];
  assign N3543 = N3542 | data_masked[6841];
  assign N3542 = N3541 | data_masked[6969];
  assign N3541 = N3540 | data_masked[7097];
  assign N3540 = N3539 | data_masked[7225];
  assign N3539 = N3538 | data_masked[7353];
  assign N3538 = N3537 | data_masked[7481];
  assign N3537 = N3536 | data_masked[7609];
  assign N3536 = N3535 | data_masked[7737];
  assign N3535 = N3534 | data_masked[7865];
  assign N3534 = data_masked[8121] | data_masked[7993];
  assign data_o[58] = N3657 | data_masked[58];
  assign N3657 = N3656 | data_masked[186];
  assign N3656 = N3655 | data_masked[314];
  assign N3655 = N3654 | data_masked[442];
  assign N3654 = N3653 | data_masked[570];
  assign N3653 = N3652 | data_masked[698];
  assign N3652 = N3651 | data_masked[826];
  assign N3651 = N3650 | data_masked[954];
  assign N3650 = N3649 | data_masked[1082];
  assign N3649 = N3648 | data_masked[1210];
  assign N3648 = N3647 | data_masked[1338];
  assign N3647 = N3646 | data_masked[1466];
  assign N3646 = N3645 | data_masked[1594];
  assign N3645 = N3644 | data_masked[1722];
  assign N3644 = N3643 | data_masked[1850];
  assign N3643 = N3642 | data_masked[1978];
  assign N3642 = N3641 | data_masked[2106];
  assign N3641 = N3640 | data_masked[2234];
  assign N3640 = N3639 | data_masked[2362];
  assign N3639 = N3638 | data_masked[2490];
  assign N3638 = N3637 | data_masked[2618];
  assign N3637 = N3636 | data_masked[2746];
  assign N3636 = N3635 | data_masked[2874];
  assign N3635 = N3634 | data_masked[3002];
  assign N3634 = N3633 | data_masked[3130];
  assign N3633 = N3632 | data_masked[3258];
  assign N3632 = N3631 | data_masked[3386];
  assign N3631 = N3630 | data_masked[3514];
  assign N3630 = N3629 | data_masked[3642];
  assign N3629 = N3628 | data_masked[3770];
  assign N3628 = N3627 | data_masked[3898];
  assign N3627 = N3626 | data_masked[4026];
  assign N3626 = N3625 | data_masked[4154];
  assign N3625 = N3624 | data_masked[4282];
  assign N3624 = N3623 | data_masked[4410];
  assign N3623 = N3622 | data_masked[4538];
  assign N3622 = N3621 | data_masked[4666];
  assign N3621 = N3620 | data_masked[4794];
  assign N3620 = N3619 | data_masked[4922];
  assign N3619 = N3618 | data_masked[5050];
  assign N3618 = N3617 | data_masked[5178];
  assign N3617 = N3616 | data_masked[5306];
  assign N3616 = N3615 | data_masked[5434];
  assign N3615 = N3614 | data_masked[5562];
  assign N3614 = N3613 | data_masked[5690];
  assign N3613 = N3612 | data_masked[5818];
  assign N3612 = N3611 | data_masked[5946];
  assign N3611 = N3610 | data_masked[6074];
  assign N3610 = N3609 | data_masked[6202];
  assign N3609 = N3608 | data_masked[6330];
  assign N3608 = N3607 | data_masked[6458];
  assign N3607 = N3606 | data_masked[6586];
  assign N3606 = N3605 | data_masked[6714];
  assign N3605 = N3604 | data_masked[6842];
  assign N3604 = N3603 | data_masked[6970];
  assign N3603 = N3602 | data_masked[7098];
  assign N3602 = N3601 | data_masked[7226];
  assign N3601 = N3600 | data_masked[7354];
  assign N3600 = N3599 | data_masked[7482];
  assign N3599 = N3598 | data_masked[7610];
  assign N3598 = N3597 | data_masked[7738];
  assign N3597 = N3596 | data_masked[7866];
  assign N3596 = data_masked[8122] | data_masked[7994];
  assign data_o[59] = N3719 | data_masked[59];
  assign N3719 = N3718 | data_masked[187];
  assign N3718 = N3717 | data_masked[315];
  assign N3717 = N3716 | data_masked[443];
  assign N3716 = N3715 | data_masked[571];
  assign N3715 = N3714 | data_masked[699];
  assign N3714 = N3713 | data_masked[827];
  assign N3713 = N3712 | data_masked[955];
  assign N3712 = N3711 | data_masked[1083];
  assign N3711 = N3710 | data_masked[1211];
  assign N3710 = N3709 | data_masked[1339];
  assign N3709 = N3708 | data_masked[1467];
  assign N3708 = N3707 | data_masked[1595];
  assign N3707 = N3706 | data_masked[1723];
  assign N3706 = N3705 | data_masked[1851];
  assign N3705 = N3704 | data_masked[1979];
  assign N3704 = N3703 | data_masked[2107];
  assign N3703 = N3702 | data_masked[2235];
  assign N3702 = N3701 | data_masked[2363];
  assign N3701 = N3700 | data_masked[2491];
  assign N3700 = N3699 | data_masked[2619];
  assign N3699 = N3698 | data_masked[2747];
  assign N3698 = N3697 | data_masked[2875];
  assign N3697 = N3696 | data_masked[3003];
  assign N3696 = N3695 | data_masked[3131];
  assign N3695 = N3694 | data_masked[3259];
  assign N3694 = N3693 | data_masked[3387];
  assign N3693 = N3692 | data_masked[3515];
  assign N3692 = N3691 | data_masked[3643];
  assign N3691 = N3690 | data_masked[3771];
  assign N3690 = N3689 | data_masked[3899];
  assign N3689 = N3688 | data_masked[4027];
  assign N3688 = N3687 | data_masked[4155];
  assign N3687 = N3686 | data_masked[4283];
  assign N3686 = N3685 | data_masked[4411];
  assign N3685 = N3684 | data_masked[4539];
  assign N3684 = N3683 | data_masked[4667];
  assign N3683 = N3682 | data_masked[4795];
  assign N3682 = N3681 | data_masked[4923];
  assign N3681 = N3680 | data_masked[5051];
  assign N3680 = N3679 | data_masked[5179];
  assign N3679 = N3678 | data_masked[5307];
  assign N3678 = N3677 | data_masked[5435];
  assign N3677 = N3676 | data_masked[5563];
  assign N3676 = N3675 | data_masked[5691];
  assign N3675 = N3674 | data_masked[5819];
  assign N3674 = N3673 | data_masked[5947];
  assign N3673 = N3672 | data_masked[6075];
  assign N3672 = N3671 | data_masked[6203];
  assign N3671 = N3670 | data_masked[6331];
  assign N3670 = N3669 | data_masked[6459];
  assign N3669 = N3668 | data_masked[6587];
  assign N3668 = N3667 | data_masked[6715];
  assign N3667 = N3666 | data_masked[6843];
  assign N3666 = N3665 | data_masked[6971];
  assign N3665 = N3664 | data_masked[7099];
  assign N3664 = N3663 | data_masked[7227];
  assign N3663 = N3662 | data_masked[7355];
  assign N3662 = N3661 | data_masked[7483];
  assign N3661 = N3660 | data_masked[7611];
  assign N3660 = N3659 | data_masked[7739];
  assign N3659 = N3658 | data_masked[7867];
  assign N3658 = data_masked[8123] | data_masked[7995];
  assign data_o[60] = N3781 | data_masked[60];
  assign N3781 = N3780 | data_masked[188];
  assign N3780 = N3779 | data_masked[316];
  assign N3779 = N3778 | data_masked[444];
  assign N3778 = N3777 | data_masked[572];
  assign N3777 = N3776 | data_masked[700];
  assign N3776 = N3775 | data_masked[828];
  assign N3775 = N3774 | data_masked[956];
  assign N3774 = N3773 | data_masked[1084];
  assign N3773 = N3772 | data_masked[1212];
  assign N3772 = N3771 | data_masked[1340];
  assign N3771 = N3770 | data_masked[1468];
  assign N3770 = N3769 | data_masked[1596];
  assign N3769 = N3768 | data_masked[1724];
  assign N3768 = N3767 | data_masked[1852];
  assign N3767 = N3766 | data_masked[1980];
  assign N3766 = N3765 | data_masked[2108];
  assign N3765 = N3764 | data_masked[2236];
  assign N3764 = N3763 | data_masked[2364];
  assign N3763 = N3762 | data_masked[2492];
  assign N3762 = N3761 | data_masked[2620];
  assign N3761 = N3760 | data_masked[2748];
  assign N3760 = N3759 | data_masked[2876];
  assign N3759 = N3758 | data_masked[3004];
  assign N3758 = N3757 | data_masked[3132];
  assign N3757 = N3756 | data_masked[3260];
  assign N3756 = N3755 | data_masked[3388];
  assign N3755 = N3754 | data_masked[3516];
  assign N3754 = N3753 | data_masked[3644];
  assign N3753 = N3752 | data_masked[3772];
  assign N3752 = N3751 | data_masked[3900];
  assign N3751 = N3750 | data_masked[4028];
  assign N3750 = N3749 | data_masked[4156];
  assign N3749 = N3748 | data_masked[4284];
  assign N3748 = N3747 | data_masked[4412];
  assign N3747 = N3746 | data_masked[4540];
  assign N3746 = N3745 | data_masked[4668];
  assign N3745 = N3744 | data_masked[4796];
  assign N3744 = N3743 | data_masked[4924];
  assign N3743 = N3742 | data_masked[5052];
  assign N3742 = N3741 | data_masked[5180];
  assign N3741 = N3740 | data_masked[5308];
  assign N3740 = N3739 | data_masked[5436];
  assign N3739 = N3738 | data_masked[5564];
  assign N3738 = N3737 | data_masked[5692];
  assign N3737 = N3736 | data_masked[5820];
  assign N3736 = N3735 | data_masked[5948];
  assign N3735 = N3734 | data_masked[6076];
  assign N3734 = N3733 | data_masked[6204];
  assign N3733 = N3732 | data_masked[6332];
  assign N3732 = N3731 | data_masked[6460];
  assign N3731 = N3730 | data_masked[6588];
  assign N3730 = N3729 | data_masked[6716];
  assign N3729 = N3728 | data_masked[6844];
  assign N3728 = N3727 | data_masked[6972];
  assign N3727 = N3726 | data_masked[7100];
  assign N3726 = N3725 | data_masked[7228];
  assign N3725 = N3724 | data_masked[7356];
  assign N3724 = N3723 | data_masked[7484];
  assign N3723 = N3722 | data_masked[7612];
  assign N3722 = N3721 | data_masked[7740];
  assign N3721 = N3720 | data_masked[7868];
  assign N3720 = data_masked[8124] | data_masked[7996];
  assign data_o[61] = N3843 | data_masked[61];
  assign N3843 = N3842 | data_masked[189];
  assign N3842 = N3841 | data_masked[317];
  assign N3841 = N3840 | data_masked[445];
  assign N3840 = N3839 | data_masked[573];
  assign N3839 = N3838 | data_masked[701];
  assign N3838 = N3837 | data_masked[829];
  assign N3837 = N3836 | data_masked[957];
  assign N3836 = N3835 | data_masked[1085];
  assign N3835 = N3834 | data_masked[1213];
  assign N3834 = N3833 | data_masked[1341];
  assign N3833 = N3832 | data_masked[1469];
  assign N3832 = N3831 | data_masked[1597];
  assign N3831 = N3830 | data_masked[1725];
  assign N3830 = N3829 | data_masked[1853];
  assign N3829 = N3828 | data_masked[1981];
  assign N3828 = N3827 | data_masked[2109];
  assign N3827 = N3826 | data_masked[2237];
  assign N3826 = N3825 | data_masked[2365];
  assign N3825 = N3824 | data_masked[2493];
  assign N3824 = N3823 | data_masked[2621];
  assign N3823 = N3822 | data_masked[2749];
  assign N3822 = N3821 | data_masked[2877];
  assign N3821 = N3820 | data_masked[3005];
  assign N3820 = N3819 | data_masked[3133];
  assign N3819 = N3818 | data_masked[3261];
  assign N3818 = N3817 | data_masked[3389];
  assign N3817 = N3816 | data_masked[3517];
  assign N3816 = N3815 | data_masked[3645];
  assign N3815 = N3814 | data_masked[3773];
  assign N3814 = N3813 | data_masked[3901];
  assign N3813 = N3812 | data_masked[4029];
  assign N3812 = N3811 | data_masked[4157];
  assign N3811 = N3810 | data_masked[4285];
  assign N3810 = N3809 | data_masked[4413];
  assign N3809 = N3808 | data_masked[4541];
  assign N3808 = N3807 | data_masked[4669];
  assign N3807 = N3806 | data_masked[4797];
  assign N3806 = N3805 | data_masked[4925];
  assign N3805 = N3804 | data_masked[5053];
  assign N3804 = N3803 | data_masked[5181];
  assign N3803 = N3802 | data_masked[5309];
  assign N3802 = N3801 | data_masked[5437];
  assign N3801 = N3800 | data_masked[5565];
  assign N3800 = N3799 | data_masked[5693];
  assign N3799 = N3798 | data_masked[5821];
  assign N3798 = N3797 | data_masked[5949];
  assign N3797 = N3796 | data_masked[6077];
  assign N3796 = N3795 | data_masked[6205];
  assign N3795 = N3794 | data_masked[6333];
  assign N3794 = N3793 | data_masked[6461];
  assign N3793 = N3792 | data_masked[6589];
  assign N3792 = N3791 | data_masked[6717];
  assign N3791 = N3790 | data_masked[6845];
  assign N3790 = N3789 | data_masked[6973];
  assign N3789 = N3788 | data_masked[7101];
  assign N3788 = N3787 | data_masked[7229];
  assign N3787 = N3786 | data_masked[7357];
  assign N3786 = N3785 | data_masked[7485];
  assign N3785 = N3784 | data_masked[7613];
  assign N3784 = N3783 | data_masked[7741];
  assign N3783 = N3782 | data_masked[7869];
  assign N3782 = data_masked[8125] | data_masked[7997];
  assign data_o[62] = N3905 | data_masked[62];
  assign N3905 = N3904 | data_masked[190];
  assign N3904 = N3903 | data_masked[318];
  assign N3903 = N3902 | data_masked[446];
  assign N3902 = N3901 | data_masked[574];
  assign N3901 = N3900 | data_masked[702];
  assign N3900 = N3899 | data_masked[830];
  assign N3899 = N3898 | data_masked[958];
  assign N3898 = N3897 | data_masked[1086];
  assign N3897 = N3896 | data_masked[1214];
  assign N3896 = N3895 | data_masked[1342];
  assign N3895 = N3894 | data_masked[1470];
  assign N3894 = N3893 | data_masked[1598];
  assign N3893 = N3892 | data_masked[1726];
  assign N3892 = N3891 | data_masked[1854];
  assign N3891 = N3890 | data_masked[1982];
  assign N3890 = N3889 | data_masked[2110];
  assign N3889 = N3888 | data_masked[2238];
  assign N3888 = N3887 | data_masked[2366];
  assign N3887 = N3886 | data_masked[2494];
  assign N3886 = N3885 | data_masked[2622];
  assign N3885 = N3884 | data_masked[2750];
  assign N3884 = N3883 | data_masked[2878];
  assign N3883 = N3882 | data_masked[3006];
  assign N3882 = N3881 | data_masked[3134];
  assign N3881 = N3880 | data_masked[3262];
  assign N3880 = N3879 | data_masked[3390];
  assign N3879 = N3878 | data_masked[3518];
  assign N3878 = N3877 | data_masked[3646];
  assign N3877 = N3876 | data_masked[3774];
  assign N3876 = N3875 | data_masked[3902];
  assign N3875 = N3874 | data_masked[4030];
  assign N3874 = N3873 | data_masked[4158];
  assign N3873 = N3872 | data_masked[4286];
  assign N3872 = N3871 | data_masked[4414];
  assign N3871 = N3870 | data_masked[4542];
  assign N3870 = N3869 | data_masked[4670];
  assign N3869 = N3868 | data_masked[4798];
  assign N3868 = N3867 | data_masked[4926];
  assign N3867 = N3866 | data_masked[5054];
  assign N3866 = N3865 | data_masked[5182];
  assign N3865 = N3864 | data_masked[5310];
  assign N3864 = N3863 | data_masked[5438];
  assign N3863 = N3862 | data_masked[5566];
  assign N3862 = N3861 | data_masked[5694];
  assign N3861 = N3860 | data_masked[5822];
  assign N3860 = N3859 | data_masked[5950];
  assign N3859 = N3858 | data_masked[6078];
  assign N3858 = N3857 | data_masked[6206];
  assign N3857 = N3856 | data_masked[6334];
  assign N3856 = N3855 | data_masked[6462];
  assign N3855 = N3854 | data_masked[6590];
  assign N3854 = N3853 | data_masked[6718];
  assign N3853 = N3852 | data_masked[6846];
  assign N3852 = N3851 | data_masked[6974];
  assign N3851 = N3850 | data_masked[7102];
  assign N3850 = N3849 | data_masked[7230];
  assign N3849 = N3848 | data_masked[7358];
  assign N3848 = N3847 | data_masked[7486];
  assign N3847 = N3846 | data_masked[7614];
  assign N3846 = N3845 | data_masked[7742];
  assign N3845 = N3844 | data_masked[7870];
  assign N3844 = data_masked[8126] | data_masked[7998];
  assign data_o[63] = N3967 | data_masked[63];
  assign N3967 = N3966 | data_masked[191];
  assign N3966 = N3965 | data_masked[319];
  assign N3965 = N3964 | data_masked[447];
  assign N3964 = N3963 | data_masked[575];
  assign N3963 = N3962 | data_masked[703];
  assign N3962 = N3961 | data_masked[831];
  assign N3961 = N3960 | data_masked[959];
  assign N3960 = N3959 | data_masked[1087];
  assign N3959 = N3958 | data_masked[1215];
  assign N3958 = N3957 | data_masked[1343];
  assign N3957 = N3956 | data_masked[1471];
  assign N3956 = N3955 | data_masked[1599];
  assign N3955 = N3954 | data_masked[1727];
  assign N3954 = N3953 | data_masked[1855];
  assign N3953 = N3952 | data_masked[1983];
  assign N3952 = N3951 | data_masked[2111];
  assign N3951 = N3950 | data_masked[2239];
  assign N3950 = N3949 | data_masked[2367];
  assign N3949 = N3948 | data_masked[2495];
  assign N3948 = N3947 | data_masked[2623];
  assign N3947 = N3946 | data_masked[2751];
  assign N3946 = N3945 | data_masked[2879];
  assign N3945 = N3944 | data_masked[3007];
  assign N3944 = N3943 | data_masked[3135];
  assign N3943 = N3942 | data_masked[3263];
  assign N3942 = N3941 | data_masked[3391];
  assign N3941 = N3940 | data_masked[3519];
  assign N3940 = N3939 | data_masked[3647];
  assign N3939 = N3938 | data_masked[3775];
  assign N3938 = N3937 | data_masked[3903];
  assign N3937 = N3936 | data_masked[4031];
  assign N3936 = N3935 | data_masked[4159];
  assign N3935 = N3934 | data_masked[4287];
  assign N3934 = N3933 | data_masked[4415];
  assign N3933 = N3932 | data_masked[4543];
  assign N3932 = N3931 | data_masked[4671];
  assign N3931 = N3930 | data_masked[4799];
  assign N3930 = N3929 | data_masked[4927];
  assign N3929 = N3928 | data_masked[5055];
  assign N3928 = N3927 | data_masked[5183];
  assign N3927 = N3926 | data_masked[5311];
  assign N3926 = N3925 | data_masked[5439];
  assign N3925 = N3924 | data_masked[5567];
  assign N3924 = N3923 | data_masked[5695];
  assign N3923 = N3922 | data_masked[5823];
  assign N3922 = N3921 | data_masked[5951];
  assign N3921 = N3920 | data_masked[6079];
  assign N3920 = N3919 | data_masked[6207];
  assign N3919 = N3918 | data_masked[6335];
  assign N3918 = N3917 | data_masked[6463];
  assign N3917 = N3916 | data_masked[6591];
  assign N3916 = N3915 | data_masked[6719];
  assign N3915 = N3914 | data_masked[6847];
  assign N3914 = N3913 | data_masked[6975];
  assign N3913 = N3912 | data_masked[7103];
  assign N3912 = N3911 | data_masked[7231];
  assign N3911 = N3910 | data_masked[7359];
  assign N3910 = N3909 | data_masked[7487];
  assign N3909 = N3908 | data_masked[7615];
  assign N3908 = N3907 | data_masked[7743];
  assign N3907 = N3906 | data_masked[7871];
  assign N3906 = data_masked[8127] | data_masked[7999];
  assign data_o[64] = N4029 | data_masked[64];
  assign N4029 = N4028 | data_masked[192];
  assign N4028 = N4027 | data_masked[320];
  assign N4027 = N4026 | data_masked[448];
  assign N4026 = N4025 | data_masked[576];
  assign N4025 = N4024 | data_masked[704];
  assign N4024 = N4023 | data_masked[832];
  assign N4023 = N4022 | data_masked[960];
  assign N4022 = N4021 | data_masked[1088];
  assign N4021 = N4020 | data_masked[1216];
  assign N4020 = N4019 | data_masked[1344];
  assign N4019 = N4018 | data_masked[1472];
  assign N4018 = N4017 | data_masked[1600];
  assign N4017 = N4016 | data_masked[1728];
  assign N4016 = N4015 | data_masked[1856];
  assign N4015 = N4014 | data_masked[1984];
  assign N4014 = N4013 | data_masked[2112];
  assign N4013 = N4012 | data_masked[2240];
  assign N4012 = N4011 | data_masked[2368];
  assign N4011 = N4010 | data_masked[2496];
  assign N4010 = N4009 | data_masked[2624];
  assign N4009 = N4008 | data_masked[2752];
  assign N4008 = N4007 | data_masked[2880];
  assign N4007 = N4006 | data_masked[3008];
  assign N4006 = N4005 | data_masked[3136];
  assign N4005 = N4004 | data_masked[3264];
  assign N4004 = N4003 | data_masked[3392];
  assign N4003 = N4002 | data_masked[3520];
  assign N4002 = N4001 | data_masked[3648];
  assign N4001 = N4000 | data_masked[3776];
  assign N4000 = N3999 | data_masked[3904];
  assign N3999 = N3998 | data_masked[4032];
  assign N3998 = N3997 | data_masked[4160];
  assign N3997 = N3996 | data_masked[4288];
  assign N3996 = N3995 | data_masked[4416];
  assign N3995 = N3994 | data_masked[4544];
  assign N3994 = N3993 | data_masked[4672];
  assign N3993 = N3992 | data_masked[4800];
  assign N3992 = N3991 | data_masked[4928];
  assign N3991 = N3990 | data_masked[5056];
  assign N3990 = N3989 | data_masked[5184];
  assign N3989 = N3988 | data_masked[5312];
  assign N3988 = N3987 | data_masked[5440];
  assign N3987 = N3986 | data_masked[5568];
  assign N3986 = N3985 | data_masked[5696];
  assign N3985 = N3984 | data_masked[5824];
  assign N3984 = N3983 | data_masked[5952];
  assign N3983 = N3982 | data_masked[6080];
  assign N3982 = N3981 | data_masked[6208];
  assign N3981 = N3980 | data_masked[6336];
  assign N3980 = N3979 | data_masked[6464];
  assign N3979 = N3978 | data_masked[6592];
  assign N3978 = N3977 | data_masked[6720];
  assign N3977 = N3976 | data_masked[6848];
  assign N3976 = N3975 | data_masked[6976];
  assign N3975 = N3974 | data_masked[7104];
  assign N3974 = N3973 | data_masked[7232];
  assign N3973 = N3972 | data_masked[7360];
  assign N3972 = N3971 | data_masked[7488];
  assign N3971 = N3970 | data_masked[7616];
  assign N3970 = N3969 | data_masked[7744];
  assign N3969 = N3968 | data_masked[7872];
  assign N3968 = data_masked[8128] | data_masked[8000];
  assign data_o[65] = N4091 | data_masked[65];
  assign N4091 = N4090 | data_masked[193];
  assign N4090 = N4089 | data_masked[321];
  assign N4089 = N4088 | data_masked[449];
  assign N4088 = N4087 | data_masked[577];
  assign N4087 = N4086 | data_masked[705];
  assign N4086 = N4085 | data_masked[833];
  assign N4085 = N4084 | data_masked[961];
  assign N4084 = N4083 | data_masked[1089];
  assign N4083 = N4082 | data_masked[1217];
  assign N4082 = N4081 | data_masked[1345];
  assign N4081 = N4080 | data_masked[1473];
  assign N4080 = N4079 | data_masked[1601];
  assign N4079 = N4078 | data_masked[1729];
  assign N4078 = N4077 | data_masked[1857];
  assign N4077 = N4076 | data_masked[1985];
  assign N4076 = N4075 | data_masked[2113];
  assign N4075 = N4074 | data_masked[2241];
  assign N4074 = N4073 | data_masked[2369];
  assign N4073 = N4072 | data_masked[2497];
  assign N4072 = N4071 | data_masked[2625];
  assign N4071 = N4070 | data_masked[2753];
  assign N4070 = N4069 | data_masked[2881];
  assign N4069 = N4068 | data_masked[3009];
  assign N4068 = N4067 | data_masked[3137];
  assign N4067 = N4066 | data_masked[3265];
  assign N4066 = N4065 | data_masked[3393];
  assign N4065 = N4064 | data_masked[3521];
  assign N4064 = N4063 | data_masked[3649];
  assign N4063 = N4062 | data_masked[3777];
  assign N4062 = N4061 | data_masked[3905];
  assign N4061 = N4060 | data_masked[4033];
  assign N4060 = N4059 | data_masked[4161];
  assign N4059 = N4058 | data_masked[4289];
  assign N4058 = N4057 | data_masked[4417];
  assign N4057 = N4056 | data_masked[4545];
  assign N4056 = N4055 | data_masked[4673];
  assign N4055 = N4054 | data_masked[4801];
  assign N4054 = N4053 | data_masked[4929];
  assign N4053 = N4052 | data_masked[5057];
  assign N4052 = N4051 | data_masked[5185];
  assign N4051 = N4050 | data_masked[5313];
  assign N4050 = N4049 | data_masked[5441];
  assign N4049 = N4048 | data_masked[5569];
  assign N4048 = N4047 | data_masked[5697];
  assign N4047 = N4046 | data_masked[5825];
  assign N4046 = N4045 | data_masked[5953];
  assign N4045 = N4044 | data_masked[6081];
  assign N4044 = N4043 | data_masked[6209];
  assign N4043 = N4042 | data_masked[6337];
  assign N4042 = N4041 | data_masked[6465];
  assign N4041 = N4040 | data_masked[6593];
  assign N4040 = N4039 | data_masked[6721];
  assign N4039 = N4038 | data_masked[6849];
  assign N4038 = N4037 | data_masked[6977];
  assign N4037 = N4036 | data_masked[7105];
  assign N4036 = N4035 | data_masked[7233];
  assign N4035 = N4034 | data_masked[7361];
  assign N4034 = N4033 | data_masked[7489];
  assign N4033 = N4032 | data_masked[7617];
  assign N4032 = N4031 | data_masked[7745];
  assign N4031 = N4030 | data_masked[7873];
  assign N4030 = data_masked[8129] | data_masked[8001];
  assign data_o[66] = N4153 | data_masked[66];
  assign N4153 = N4152 | data_masked[194];
  assign N4152 = N4151 | data_masked[322];
  assign N4151 = N4150 | data_masked[450];
  assign N4150 = N4149 | data_masked[578];
  assign N4149 = N4148 | data_masked[706];
  assign N4148 = N4147 | data_masked[834];
  assign N4147 = N4146 | data_masked[962];
  assign N4146 = N4145 | data_masked[1090];
  assign N4145 = N4144 | data_masked[1218];
  assign N4144 = N4143 | data_masked[1346];
  assign N4143 = N4142 | data_masked[1474];
  assign N4142 = N4141 | data_masked[1602];
  assign N4141 = N4140 | data_masked[1730];
  assign N4140 = N4139 | data_masked[1858];
  assign N4139 = N4138 | data_masked[1986];
  assign N4138 = N4137 | data_masked[2114];
  assign N4137 = N4136 | data_masked[2242];
  assign N4136 = N4135 | data_masked[2370];
  assign N4135 = N4134 | data_masked[2498];
  assign N4134 = N4133 | data_masked[2626];
  assign N4133 = N4132 | data_masked[2754];
  assign N4132 = N4131 | data_masked[2882];
  assign N4131 = N4130 | data_masked[3010];
  assign N4130 = N4129 | data_masked[3138];
  assign N4129 = N4128 | data_masked[3266];
  assign N4128 = N4127 | data_masked[3394];
  assign N4127 = N4126 | data_masked[3522];
  assign N4126 = N4125 | data_masked[3650];
  assign N4125 = N4124 | data_masked[3778];
  assign N4124 = N4123 | data_masked[3906];
  assign N4123 = N4122 | data_masked[4034];
  assign N4122 = N4121 | data_masked[4162];
  assign N4121 = N4120 | data_masked[4290];
  assign N4120 = N4119 | data_masked[4418];
  assign N4119 = N4118 | data_masked[4546];
  assign N4118 = N4117 | data_masked[4674];
  assign N4117 = N4116 | data_masked[4802];
  assign N4116 = N4115 | data_masked[4930];
  assign N4115 = N4114 | data_masked[5058];
  assign N4114 = N4113 | data_masked[5186];
  assign N4113 = N4112 | data_masked[5314];
  assign N4112 = N4111 | data_masked[5442];
  assign N4111 = N4110 | data_masked[5570];
  assign N4110 = N4109 | data_masked[5698];
  assign N4109 = N4108 | data_masked[5826];
  assign N4108 = N4107 | data_masked[5954];
  assign N4107 = N4106 | data_masked[6082];
  assign N4106 = N4105 | data_masked[6210];
  assign N4105 = N4104 | data_masked[6338];
  assign N4104 = N4103 | data_masked[6466];
  assign N4103 = N4102 | data_masked[6594];
  assign N4102 = N4101 | data_masked[6722];
  assign N4101 = N4100 | data_masked[6850];
  assign N4100 = N4099 | data_masked[6978];
  assign N4099 = N4098 | data_masked[7106];
  assign N4098 = N4097 | data_masked[7234];
  assign N4097 = N4096 | data_masked[7362];
  assign N4096 = N4095 | data_masked[7490];
  assign N4095 = N4094 | data_masked[7618];
  assign N4094 = N4093 | data_masked[7746];
  assign N4093 = N4092 | data_masked[7874];
  assign N4092 = data_masked[8130] | data_masked[8002];
  assign data_o[67] = N4215 | data_masked[67];
  assign N4215 = N4214 | data_masked[195];
  assign N4214 = N4213 | data_masked[323];
  assign N4213 = N4212 | data_masked[451];
  assign N4212 = N4211 | data_masked[579];
  assign N4211 = N4210 | data_masked[707];
  assign N4210 = N4209 | data_masked[835];
  assign N4209 = N4208 | data_masked[963];
  assign N4208 = N4207 | data_masked[1091];
  assign N4207 = N4206 | data_masked[1219];
  assign N4206 = N4205 | data_masked[1347];
  assign N4205 = N4204 | data_masked[1475];
  assign N4204 = N4203 | data_masked[1603];
  assign N4203 = N4202 | data_masked[1731];
  assign N4202 = N4201 | data_masked[1859];
  assign N4201 = N4200 | data_masked[1987];
  assign N4200 = N4199 | data_masked[2115];
  assign N4199 = N4198 | data_masked[2243];
  assign N4198 = N4197 | data_masked[2371];
  assign N4197 = N4196 | data_masked[2499];
  assign N4196 = N4195 | data_masked[2627];
  assign N4195 = N4194 | data_masked[2755];
  assign N4194 = N4193 | data_masked[2883];
  assign N4193 = N4192 | data_masked[3011];
  assign N4192 = N4191 | data_masked[3139];
  assign N4191 = N4190 | data_masked[3267];
  assign N4190 = N4189 | data_masked[3395];
  assign N4189 = N4188 | data_masked[3523];
  assign N4188 = N4187 | data_masked[3651];
  assign N4187 = N4186 | data_masked[3779];
  assign N4186 = N4185 | data_masked[3907];
  assign N4185 = N4184 | data_masked[4035];
  assign N4184 = N4183 | data_masked[4163];
  assign N4183 = N4182 | data_masked[4291];
  assign N4182 = N4181 | data_masked[4419];
  assign N4181 = N4180 | data_masked[4547];
  assign N4180 = N4179 | data_masked[4675];
  assign N4179 = N4178 | data_masked[4803];
  assign N4178 = N4177 | data_masked[4931];
  assign N4177 = N4176 | data_masked[5059];
  assign N4176 = N4175 | data_masked[5187];
  assign N4175 = N4174 | data_masked[5315];
  assign N4174 = N4173 | data_masked[5443];
  assign N4173 = N4172 | data_masked[5571];
  assign N4172 = N4171 | data_masked[5699];
  assign N4171 = N4170 | data_masked[5827];
  assign N4170 = N4169 | data_masked[5955];
  assign N4169 = N4168 | data_masked[6083];
  assign N4168 = N4167 | data_masked[6211];
  assign N4167 = N4166 | data_masked[6339];
  assign N4166 = N4165 | data_masked[6467];
  assign N4165 = N4164 | data_masked[6595];
  assign N4164 = N4163 | data_masked[6723];
  assign N4163 = N4162 | data_masked[6851];
  assign N4162 = N4161 | data_masked[6979];
  assign N4161 = N4160 | data_masked[7107];
  assign N4160 = N4159 | data_masked[7235];
  assign N4159 = N4158 | data_masked[7363];
  assign N4158 = N4157 | data_masked[7491];
  assign N4157 = N4156 | data_masked[7619];
  assign N4156 = N4155 | data_masked[7747];
  assign N4155 = N4154 | data_masked[7875];
  assign N4154 = data_masked[8131] | data_masked[8003];
  assign data_o[68] = N4277 | data_masked[68];
  assign N4277 = N4276 | data_masked[196];
  assign N4276 = N4275 | data_masked[324];
  assign N4275 = N4274 | data_masked[452];
  assign N4274 = N4273 | data_masked[580];
  assign N4273 = N4272 | data_masked[708];
  assign N4272 = N4271 | data_masked[836];
  assign N4271 = N4270 | data_masked[964];
  assign N4270 = N4269 | data_masked[1092];
  assign N4269 = N4268 | data_masked[1220];
  assign N4268 = N4267 | data_masked[1348];
  assign N4267 = N4266 | data_masked[1476];
  assign N4266 = N4265 | data_masked[1604];
  assign N4265 = N4264 | data_masked[1732];
  assign N4264 = N4263 | data_masked[1860];
  assign N4263 = N4262 | data_masked[1988];
  assign N4262 = N4261 | data_masked[2116];
  assign N4261 = N4260 | data_masked[2244];
  assign N4260 = N4259 | data_masked[2372];
  assign N4259 = N4258 | data_masked[2500];
  assign N4258 = N4257 | data_masked[2628];
  assign N4257 = N4256 | data_masked[2756];
  assign N4256 = N4255 | data_masked[2884];
  assign N4255 = N4254 | data_masked[3012];
  assign N4254 = N4253 | data_masked[3140];
  assign N4253 = N4252 | data_masked[3268];
  assign N4252 = N4251 | data_masked[3396];
  assign N4251 = N4250 | data_masked[3524];
  assign N4250 = N4249 | data_masked[3652];
  assign N4249 = N4248 | data_masked[3780];
  assign N4248 = N4247 | data_masked[3908];
  assign N4247 = N4246 | data_masked[4036];
  assign N4246 = N4245 | data_masked[4164];
  assign N4245 = N4244 | data_masked[4292];
  assign N4244 = N4243 | data_masked[4420];
  assign N4243 = N4242 | data_masked[4548];
  assign N4242 = N4241 | data_masked[4676];
  assign N4241 = N4240 | data_masked[4804];
  assign N4240 = N4239 | data_masked[4932];
  assign N4239 = N4238 | data_masked[5060];
  assign N4238 = N4237 | data_masked[5188];
  assign N4237 = N4236 | data_masked[5316];
  assign N4236 = N4235 | data_masked[5444];
  assign N4235 = N4234 | data_masked[5572];
  assign N4234 = N4233 | data_masked[5700];
  assign N4233 = N4232 | data_masked[5828];
  assign N4232 = N4231 | data_masked[5956];
  assign N4231 = N4230 | data_masked[6084];
  assign N4230 = N4229 | data_masked[6212];
  assign N4229 = N4228 | data_masked[6340];
  assign N4228 = N4227 | data_masked[6468];
  assign N4227 = N4226 | data_masked[6596];
  assign N4226 = N4225 | data_masked[6724];
  assign N4225 = N4224 | data_masked[6852];
  assign N4224 = N4223 | data_masked[6980];
  assign N4223 = N4222 | data_masked[7108];
  assign N4222 = N4221 | data_masked[7236];
  assign N4221 = N4220 | data_masked[7364];
  assign N4220 = N4219 | data_masked[7492];
  assign N4219 = N4218 | data_masked[7620];
  assign N4218 = N4217 | data_masked[7748];
  assign N4217 = N4216 | data_masked[7876];
  assign N4216 = data_masked[8132] | data_masked[8004];
  assign data_o[69] = N4339 | data_masked[69];
  assign N4339 = N4338 | data_masked[197];
  assign N4338 = N4337 | data_masked[325];
  assign N4337 = N4336 | data_masked[453];
  assign N4336 = N4335 | data_masked[581];
  assign N4335 = N4334 | data_masked[709];
  assign N4334 = N4333 | data_masked[837];
  assign N4333 = N4332 | data_masked[965];
  assign N4332 = N4331 | data_masked[1093];
  assign N4331 = N4330 | data_masked[1221];
  assign N4330 = N4329 | data_masked[1349];
  assign N4329 = N4328 | data_masked[1477];
  assign N4328 = N4327 | data_masked[1605];
  assign N4327 = N4326 | data_masked[1733];
  assign N4326 = N4325 | data_masked[1861];
  assign N4325 = N4324 | data_masked[1989];
  assign N4324 = N4323 | data_masked[2117];
  assign N4323 = N4322 | data_masked[2245];
  assign N4322 = N4321 | data_masked[2373];
  assign N4321 = N4320 | data_masked[2501];
  assign N4320 = N4319 | data_masked[2629];
  assign N4319 = N4318 | data_masked[2757];
  assign N4318 = N4317 | data_masked[2885];
  assign N4317 = N4316 | data_masked[3013];
  assign N4316 = N4315 | data_masked[3141];
  assign N4315 = N4314 | data_masked[3269];
  assign N4314 = N4313 | data_masked[3397];
  assign N4313 = N4312 | data_masked[3525];
  assign N4312 = N4311 | data_masked[3653];
  assign N4311 = N4310 | data_masked[3781];
  assign N4310 = N4309 | data_masked[3909];
  assign N4309 = N4308 | data_masked[4037];
  assign N4308 = N4307 | data_masked[4165];
  assign N4307 = N4306 | data_masked[4293];
  assign N4306 = N4305 | data_masked[4421];
  assign N4305 = N4304 | data_masked[4549];
  assign N4304 = N4303 | data_masked[4677];
  assign N4303 = N4302 | data_masked[4805];
  assign N4302 = N4301 | data_masked[4933];
  assign N4301 = N4300 | data_masked[5061];
  assign N4300 = N4299 | data_masked[5189];
  assign N4299 = N4298 | data_masked[5317];
  assign N4298 = N4297 | data_masked[5445];
  assign N4297 = N4296 | data_masked[5573];
  assign N4296 = N4295 | data_masked[5701];
  assign N4295 = N4294 | data_masked[5829];
  assign N4294 = N4293 | data_masked[5957];
  assign N4293 = N4292 | data_masked[6085];
  assign N4292 = N4291 | data_masked[6213];
  assign N4291 = N4290 | data_masked[6341];
  assign N4290 = N4289 | data_masked[6469];
  assign N4289 = N4288 | data_masked[6597];
  assign N4288 = N4287 | data_masked[6725];
  assign N4287 = N4286 | data_masked[6853];
  assign N4286 = N4285 | data_masked[6981];
  assign N4285 = N4284 | data_masked[7109];
  assign N4284 = N4283 | data_masked[7237];
  assign N4283 = N4282 | data_masked[7365];
  assign N4282 = N4281 | data_masked[7493];
  assign N4281 = N4280 | data_masked[7621];
  assign N4280 = N4279 | data_masked[7749];
  assign N4279 = N4278 | data_masked[7877];
  assign N4278 = data_masked[8133] | data_masked[8005];
  assign data_o[70] = N4401 | data_masked[70];
  assign N4401 = N4400 | data_masked[198];
  assign N4400 = N4399 | data_masked[326];
  assign N4399 = N4398 | data_masked[454];
  assign N4398 = N4397 | data_masked[582];
  assign N4397 = N4396 | data_masked[710];
  assign N4396 = N4395 | data_masked[838];
  assign N4395 = N4394 | data_masked[966];
  assign N4394 = N4393 | data_masked[1094];
  assign N4393 = N4392 | data_masked[1222];
  assign N4392 = N4391 | data_masked[1350];
  assign N4391 = N4390 | data_masked[1478];
  assign N4390 = N4389 | data_masked[1606];
  assign N4389 = N4388 | data_masked[1734];
  assign N4388 = N4387 | data_masked[1862];
  assign N4387 = N4386 | data_masked[1990];
  assign N4386 = N4385 | data_masked[2118];
  assign N4385 = N4384 | data_masked[2246];
  assign N4384 = N4383 | data_masked[2374];
  assign N4383 = N4382 | data_masked[2502];
  assign N4382 = N4381 | data_masked[2630];
  assign N4381 = N4380 | data_masked[2758];
  assign N4380 = N4379 | data_masked[2886];
  assign N4379 = N4378 | data_masked[3014];
  assign N4378 = N4377 | data_masked[3142];
  assign N4377 = N4376 | data_masked[3270];
  assign N4376 = N4375 | data_masked[3398];
  assign N4375 = N4374 | data_masked[3526];
  assign N4374 = N4373 | data_masked[3654];
  assign N4373 = N4372 | data_masked[3782];
  assign N4372 = N4371 | data_masked[3910];
  assign N4371 = N4370 | data_masked[4038];
  assign N4370 = N4369 | data_masked[4166];
  assign N4369 = N4368 | data_masked[4294];
  assign N4368 = N4367 | data_masked[4422];
  assign N4367 = N4366 | data_masked[4550];
  assign N4366 = N4365 | data_masked[4678];
  assign N4365 = N4364 | data_masked[4806];
  assign N4364 = N4363 | data_masked[4934];
  assign N4363 = N4362 | data_masked[5062];
  assign N4362 = N4361 | data_masked[5190];
  assign N4361 = N4360 | data_masked[5318];
  assign N4360 = N4359 | data_masked[5446];
  assign N4359 = N4358 | data_masked[5574];
  assign N4358 = N4357 | data_masked[5702];
  assign N4357 = N4356 | data_masked[5830];
  assign N4356 = N4355 | data_masked[5958];
  assign N4355 = N4354 | data_masked[6086];
  assign N4354 = N4353 | data_masked[6214];
  assign N4353 = N4352 | data_masked[6342];
  assign N4352 = N4351 | data_masked[6470];
  assign N4351 = N4350 | data_masked[6598];
  assign N4350 = N4349 | data_masked[6726];
  assign N4349 = N4348 | data_masked[6854];
  assign N4348 = N4347 | data_masked[6982];
  assign N4347 = N4346 | data_masked[7110];
  assign N4346 = N4345 | data_masked[7238];
  assign N4345 = N4344 | data_masked[7366];
  assign N4344 = N4343 | data_masked[7494];
  assign N4343 = N4342 | data_masked[7622];
  assign N4342 = N4341 | data_masked[7750];
  assign N4341 = N4340 | data_masked[7878];
  assign N4340 = data_masked[8134] | data_masked[8006];
  assign data_o[71] = N4463 | data_masked[71];
  assign N4463 = N4462 | data_masked[199];
  assign N4462 = N4461 | data_masked[327];
  assign N4461 = N4460 | data_masked[455];
  assign N4460 = N4459 | data_masked[583];
  assign N4459 = N4458 | data_masked[711];
  assign N4458 = N4457 | data_masked[839];
  assign N4457 = N4456 | data_masked[967];
  assign N4456 = N4455 | data_masked[1095];
  assign N4455 = N4454 | data_masked[1223];
  assign N4454 = N4453 | data_masked[1351];
  assign N4453 = N4452 | data_masked[1479];
  assign N4452 = N4451 | data_masked[1607];
  assign N4451 = N4450 | data_masked[1735];
  assign N4450 = N4449 | data_masked[1863];
  assign N4449 = N4448 | data_masked[1991];
  assign N4448 = N4447 | data_masked[2119];
  assign N4447 = N4446 | data_masked[2247];
  assign N4446 = N4445 | data_masked[2375];
  assign N4445 = N4444 | data_masked[2503];
  assign N4444 = N4443 | data_masked[2631];
  assign N4443 = N4442 | data_masked[2759];
  assign N4442 = N4441 | data_masked[2887];
  assign N4441 = N4440 | data_masked[3015];
  assign N4440 = N4439 | data_masked[3143];
  assign N4439 = N4438 | data_masked[3271];
  assign N4438 = N4437 | data_masked[3399];
  assign N4437 = N4436 | data_masked[3527];
  assign N4436 = N4435 | data_masked[3655];
  assign N4435 = N4434 | data_masked[3783];
  assign N4434 = N4433 | data_masked[3911];
  assign N4433 = N4432 | data_masked[4039];
  assign N4432 = N4431 | data_masked[4167];
  assign N4431 = N4430 | data_masked[4295];
  assign N4430 = N4429 | data_masked[4423];
  assign N4429 = N4428 | data_masked[4551];
  assign N4428 = N4427 | data_masked[4679];
  assign N4427 = N4426 | data_masked[4807];
  assign N4426 = N4425 | data_masked[4935];
  assign N4425 = N4424 | data_masked[5063];
  assign N4424 = N4423 | data_masked[5191];
  assign N4423 = N4422 | data_masked[5319];
  assign N4422 = N4421 | data_masked[5447];
  assign N4421 = N4420 | data_masked[5575];
  assign N4420 = N4419 | data_masked[5703];
  assign N4419 = N4418 | data_masked[5831];
  assign N4418 = N4417 | data_masked[5959];
  assign N4417 = N4416 | data_masked[6087];
  assign N4416 = N4415 | data_masked[6215];
  assign N4415 = N4414 | data_masked[6343];
  assign N4414 = N4413 | data_masked[6471];
  assign N4413 = N4412 | data_masked[6599];
  assign N4412 = N4411 | data_masked[6727];
  assign N4411 = N4410 | data_masked[6855];
  assign N4410 = N4409 | data_masked[6983];
  assign N4409 = N4408 | data_masked[7111];
  assign N4408 = N4407 | data_masked[7239];
  assign N4407 = N4406 | data_masked[7367];
  assign N4406 = N4405 | data_masked[7495];
  assign N4405 = N4404 | data_masked[7623];
  assign N4404 = N4403 | data_masked[7751];
  assign N4403 = N4402 | data_masked[7879];
  assign N4402 = data_masked[8135] | data_masked[8007];
  assign data_o[72] = N4525 | data_masked[72];
  assign N4525 = N4524 | data_masked[200];
  assign N4524 = N4523 | data_masked[328];
  assign N4523 = N4522 | data_masked[456];
  assign N4522 = N4521 | data_masked[584];
  assign N4521 = N4520 | data_masked[712];
  assign N4520 = N4519 | data_masked[840];
  assign N4519 = N4518 | data_masked[968];
  assign N4518 = N4517 | data_masked[1096];
  assign N4517 = N4516 | data_masked[1224];
  assign N4516 = N4515 | data_masked[1352];
  assign N4515 = N4514 | data_masked[1480];
  assign N4514 = N4513 | data_masked[1608];
  assign N4513 = N4512 | data_masked[1736];
  assign N4512 = N4511 | data_masked[1864];
  assign N4511 = N4510 | data_masked[1992];
  assign N4510 = N4509 | data_masked[2120];
  assign N4509 = N4508 | data_masked[2248];
  assign N4508 = N4507 | data_masked[2376];
  assign N4507 = N4506 | data_masked[2504];
  assign N4506 = N4505 | data_masked[2632];
  assign N4505 = N4504 | data_masked[2760];
  assign N4504 = N4503 | data_masked[2888];
  assign N4503 = N4502 | data_masked[3016];
  assign N4502 = N4501 | data_masked[3144];
  assign N4501 = N4500 | data_masked[3272];
  assign N4500 = N4499 | data_masked[3400];
  assign N4499 = N4498 | data_masked[3528];
  assign N4498 = N4497 | data_masked[3656];
  assign N4497 = N4496 | data_masked[3784];
  assign N4496 = N4495 | data_masked[3912];
  assign N4495 = N4494 | data_masked[4040];
  assign N4494 = N4493 | data_masked[4168];
  assign N4493 = N4492 | data_masked[4296];
  assign N4492 = N4491 | data_masked[4424];
  assign N4491 = N4490 | data_masked[4552];
  assign N4490 = N4489 | data_masked[4680];
  assign N4489 = N4488 | data_masked[4808];
  assign N4488 = N4487 | data_masked[4936];
  assign N4487 = N4486 | data_masked[5064];
  assign N4486 = N4485 | data_masked[5192];
  assign N4485 = N4484 | data_masked[5320];
  assign N4484 = N4483 | data_masked[5448];
  assign N4483 = N4482 | data_masked[5576];
  assign N4482 = N4481 | data_masked[5704];
  assign N4481 = N4480 | data_masked[5832];
  assign N4480 = N4479 | data_masked[5960];
  assign N4479 = N4478 | data_masked[6088];
  assign N4478 = N4477 | data_masked[6216];
  assign N4477 = N4476 | data_masked[6344];
  assign N4476 = N4475 | data_masked[6472];
  assign N4475 = N4474 | data_masked[6600];
  assign N4474 = N4473 | data_masked[6728];
  assign N4473 = N4472 | data_masked[6856];
  assign N4472 = N4471 | data_masked[6984];
  assign N4471 = N4470 | data_masked[7112];
  assign N4470 = N4469 | data_masked[7240];
  assign N4469 = N4468 | data_masked[7368];
  assign N4468 = N4467 | data_masked[7496];
  assign N4467 = N4466 | data_masked[7624];
  assign N4466 = N4465 | data_masked[7752];
  assign N4465 = N4464 | data_masked[7880];
  assign N4464 = data_masked[8136] | data_masked[8008];
  assign data_o[73] = N4587 | data_masked[73];
  assign N4587 = N4586 | data_masked[201];
  assign N4586 = N4585 | data_masked[329];
  assign N4585 = N4584 | data_masked[457];
  assign N4584 = N4583 | data_masked[585];
  assign N4583 = N4582 | data_masked[713];
  assign N4582 = N4581 | data_masked[841];
  assign N4581 = N4580 | data_masked[969];
  assign N4580 = N4579 | data_masked[1097];
  assign N4579 = N4578 | data_masked[1225];
  assign N4578 = N4577 | data_masked[1353];
  assign N4577 = N4576 | data_masked[1481];
  assign N4576 = N4575 | data_masked[1609];
  assign N4575 = N4574 | data_masked[1737];
  assign N4574 = N4573 | data_masked[1865];
  assign N4573 = N4572 | data_masked[1993];
  assign N4572 = N4571 | data_masked[2121];
  assign N4571 = N4570 | data_masked[2249];
  assign N4570 = N4569 | data_masked[2377];
  assign N4569 = N4568 | data_masked[2505];
  assign N4568 = N4567 | data_masked[2633];
  assign N4567 = N4566 | data_masked[2761];
  assign N4566 = N4565 | data_masked[2889];
  assign N4565 = N4564 | data_masked[3017];
  assign N4564 = N4563 | data_masked[3145];
  assign N4563 = N4562 | data_masked[3273];
  assign N4562 = N4561 | data_masked[3401];
  assign N4561 = N4560 | data_masked[3529];
  assign N4560 = N4559 | data_masked[3657];
  assign N4559 = N4558 | data_masked[3785];
  assign N4558 = N4557 | data_masked[3913];
  assign N4557 = N4556 | data_masked[4041];
  assign N4556 = N4555 | data_masked[4169];
  assign N4555 = N4554 | data_masked[4297];
  assign N4554 = N4553 | data_masked[4425];
  assign N4553 = N4552 | data_masked[4553];
  assign N4552 = N4551 | data_masked[4681];
  assign N4551 = N4550 | data_masked[4809];
  assign N4550 = N4549 | data_masked[4937];
  assign N4549 = N4548 | data_masked[5065];
  assign N4548 = N4547 | data_masked[5193];
  assign N4547 = N4546 | data_masked[5321];
  assign N4546 = N4545 | data_masked[5449];
  assign N4545 = N4544 | data_masked[5577];
  assign N4544 = N4543 | data_masked[5705];
  assign N4543 = N4542 | data_masked[5833];
  assign N4542 = N4541 | data_masked[5961];
  assign N4541 = N4540 | data_masked[6089];
  assign N4540 = N4539 | data_masked[6217];
  assign N4539 = N4538 | data_masked[6345];
  assign N4538 = N4537 | data_masked[6473];
  assign N4537 = N4536 | data_masked[6601];
  assign N4536 = N4535 | data_masked[6729];
  assign N4535 = N4534 | data_masked[6857];
  assign N4534 = N4533 | data_masked[6985];
  assign N4533 = N4532 | data_masked[7113];
  assign N4532 = N4531 | data_masked[7241];
  assign N4531 = N4530 | data_masked[7369];
  assign N4530 = N4529 | data_masked[7497];
  assign N4529 = N4528 | data_masked[7625];
  assign N4528 = N4527 | data_masked[7753];
  assign N4527 = N4526 | data_masked[7881];
  assign N4526 = data_masked[8137] | data_masked[8009];
  assign data_o[74] = N4649 | data_masked[74];
  assign N4649 = N4648 | data_masked[202];
  assign N4648 = N4647 | data_masked[330];
  assign N4647 = N4646 | data_masked[458];
  assign N4646 = N4645 | data_masked[586];
  assign N4645 = N4644 | data_masked[714];
  assign N4644 = N4643 | data_masked[842];
  assign N4643 = N4642 | data_masked[970];
  assign N4642 = N4641 | data_masked[1098];
  assign N4641 = N4640 | data_masked[1226];
  assign N4640 = N4639 | data_masked[1354];
  assign N4639 = N4638 | data_masked[1482];
  assign N4638 = N4637 | data_masked[1610];
  assign N4637 = N4636 | data_masked[1738];
  assign N4636 = N4635 | data_masked[1866];
  assign N4635 = N4634 | data_masked[1994];
  assign N4634 = N4633 | data_masked[2122];
  assign N4633 = N4632 | data_masked[2250];
  assign N4632 = N4631 | data_masked[2378];
  assign N4631 = N4630 | data_masked[2506];
  assign N4630 = N4629 | data_masked[2634];
  assign N4629 = N4628 | data_masked[2762];
  assign N4628 = N4627 | data_masked[2890];
  assign N4627 = N4626 | data_masked[3018];
  assign N4626 = N4625 | data_masked[3146];
  assign N4625 = N4624 | data_masked[3274];
  assign N4624 = N4623 | data_masked[3402];
  assign N4623 = N4622 | data_masked[3530];
  assign N4622 = N4621 | data_masked[3658];
  assign N4621 = N4620 | data_masked[3786];
  assign N4620 = N4619 | data_masked[3914];
  assign N4619 = N4618 | data_masked[4042];
  assign N4618 = N4617 | data_masked[4170];
  assign N4617 = N4616 | data_masked[4298];
  assign N4616 = N4615 | data_masked[4426];
  assign N4615 = N4614 | data_masked[4554];
  assign N4614 = N4613 | data_masked[4682];
  assign N4613 = N4612 | data_masked[4810];
  assign N4612 = N4611 | data_masked[4938];
  assign N4611 = N4610 | data_masked[5066];
  assign N4610 = N4609 | data_masked[5194];
  assign N4609 = N4608 | data_masked[5322];
  assign N4608 = N4607 | data_masked[5450];
  assign N4607 = N4606 | data_masked[5578];
  assign N4606 = N4605 | data_masked[5706];
  assign N4605 = N4604 | data_masked[5834];
  assign N4604 = N4603 | data_masked[5962];
  assign N4603 = N4602 | data_masked[6090];
  assign N4602 = N4601 | data_masked[6218];
  assign N4601 = N4600 | data_masked[6346];
  assign N4600 = N4599 | data_masked[6474];
  assign N4599 = N4598 | data_masked[6602];
  assign N4598 = N4597 | data_masked[6730];
  assign N4597 = N4596 | data_masked[6858];
  assign N4596 = N4595 | data_masked[6986];
  assign N4595 = N4594 | data_masked[7114];
  assign N4594 = N4593 | data_masked[7242];
  assign N4593 = N4592 | data_masked[7370];
  assign N4592 = N4591 | data_masked[7498];
  assign N4591 = N4590 | data_masked[7626];
  assign N4590 = N4589 | data_masked[7754];
  assign N4589 = N4588 | data_masked[7882];
  assign N4588 = data_masked[8138] | data_masked[8010];
  assign data_o[75] = N4711 | data_masked[75];
  assign N4711 = N4710 | data_masked[203];
  assign N4710 = N4709 | data_masked[331];
  assign N4709 = N4708 | data_masked[459];
  assign N4708 = N4707 | data_masked[587];
  assign N4707 = N4706 | data_masked[715];
  assign N4706 = N4705 | data_masked[843];
  assign N4705 = N4704 | data_masked[971];
  assign N4704 = N4703 | data_masked[1099];
  assign N4703 = N4702 | data_masked[1227];
  assign N4702 = N4701 | data_masked[1355];
  assign N4701 = N4700 | data_masked[1483];
  assign N4700 = N4699 | data_masked[1611];
  assign N4699 = N4698 | data_masked[1739];
  assign N4698 = N4697 | data_masked[1867];
  assign N4697 = N4696 | data_masked[1995];
  assign N4696 = N4695 | data_masked[2123];
  assign N4695 = N4694 | data_masked[2251];
  assign N4694 = N4693 | data_masked[2379];
  assign N4693 = N4692 | data_masked[2507];
  assign N4692 = N4691 | data_masked[2635];
  assign N4691 = N4690 | data_masked[2763];
  assign N4690 = N4689 | data_masked[2891];
  assign N4689 = N4688 | data_masked[3019];
  assign N4688 = N4687 | data_masked[3147];
  assign N4687 = N4686 | data_masked[3275];
  assign N4686 = N4685 | data_masked[3403];
  assign N4685 = N4684 | data_masked[3531];
  assign N4684 = N4683 | data_masked[3659];
  assign N4683 = N4682 | data_masked[3787];
  assign N4682 = N4681 | data_masked[3915];
  assign N4681 = N4680 | data_masked[4043];
  assign N4680 = N4679 | data_masked[4171];
  assign N4679 = N4678 | data_masked[4299];
  assign N4678 = N4677 | data_masked[4427];
  assign N4677 = N4676 | data_masked[4555];
  assign N4676 = N4675 | data_masked[4683];
  assign N4675 = N4674 | data_masked[4811];
  assign N4674 = N4673 | data_masked[4939];
  assign N4673 = N4672 | data_masked[5067];
  assign N4672 = N4671 | data_masked[5195];
  assign N4671 = N4670 | data_masked[5323];
  assign N4670 = N4669 | data_masked[5451];
  assign N4669 = N4668 | data_masked[5579];
  assign N4668 = N4667 | data_masked[5707];
  assign N4667 = N4666 | data_masked[5835];
  assign N4666 = N4665 | data_masked[5963];
  assign N4665 = N4664 | data_masked[6091];
  assign N4664 = N4663 | data_masked[6219];
  assign N4663 = N4662 | data_masked[6347];
  assign N4662 = N4661 | data_masked[6475];
  assign N4661 = N4660 | data_masked[6603];
  assign N4660 = N4659 | data_masked[6731];
  assign N4659 = N4658 | data_masked[6859];
  assign N4658 = N4657 | data_masked[6987];
  assign N4657 = N4656 | data_masked[7115];
  assign N4656 = N4655 | data_masked[7243];
  assign N4655 = N4654 | data_masked[7371];
  assign N4654 = N4653 | data_masked[7499];
  assign N4653 = N4652 | data_masked[7627];
  assign N4652 = N4651 | data_masked[7755];
  assign N4651 = N4650 | data_masked[7883];
  assign N4650 = data_masked[8139] | data_masked[8011];
  assign data_o[76] = N4773 | data_masked[76];
  assign N4773 = N4772 | data_masked[204];
  assign N4772 = N4771 | data_masked[332];
  assign N4771 = N4770 | data_masked[460];
  assign N4770 = N4769 | data_masked[588];
  assign N4769 = N4768 | data_masked[716];
  assign N4768 = N4767 | data_masked[844];
  assign N4767 = N4766 | data_masked[972];
  assign N4766 = N4765 | data_masked[1100];
  assign N4765 = N4764 | data_masked[1228];
  assign N4764 = N4763 | data_masked[1356];
  assign N4763 = N4762 | data_masked[1484];
  assign N4762 = N4761 | data_masked[1612];
  assign N4761 = N4760 | data_masked[1740];
  assign N4760 = N4759 | data_masked[1868];
  assign N4759 = N4758 | data_masked[1996];
  assign N4758 = N4757 | data_masked[2124];
  assign N4757 = N4756 | data_masked[2252];
  assign N4756 = N4755 | data_masked[2380];
  assign N4755 = N4754 | data_masked[2508];
  assign N4754 = N4753 | data_masked[2636];
  assign N4753 = N4752 | data_masked[2764];
  assign N4752 = N4751 | data_masked[2892];
  assign N4751 = N4750 | data_masked[3020];
  assign N4750 = N4749 | data_masked[3148];
  assign N4749 = N4748 | data_masked[3276];
  assign N4748 = N4747 | data_masked[3404];
  assign N4747 = N4746 | data_masked[3532];
  assign N4746 = N4745 | data_masked[3660];
  assign N4745 = N4744 | data_masked[3788];
  assign N4744 = N4743 | data_masked[3916];
  assign N4743 = N4742 | data_masked[4044];
  assign N4742 = N4741 | data_masked[4172];
  assign N4741 = N4740 | data_masked[4300];
  assign N4740 = N4739 | data_masked[4428];
  assign N4739 = N4738 | data_masked[4556];
  assign N4738 = N4737 | data_masked[4684];
  assign N4737 = N4736 | data_masked[4812];
  assign N4736 = N4735 | data_masked[4940];
  assign N4735 = N4734 | data_masked[5068];
  assign N4734 = N4733 | data_masked[5196];
  assign N4733 = N4732 | data_masked[5324];
  assign N4732 = N4731 | data_masked[5452];
  assign N4731 = N4730 | data_masked[5580];
  assign N4730 = N4729 | data_masked[5708];
  assign N4729 = N4728 | data_masked[5836];
  assign N4728 = N4727 | data_masked[5964];
  assign N4727 = N4726 | data_masked[6092];
  assign N4726 = N4725 | data_masked[6220];
  assign N4725 = N4724 | data_masked[6348];
  assign N4724 = N4723 | data_masked[6476];
  assign N4723 = N4722 | data_masked[6604];
  assign N4722 = N4721 | data_masked[6732];
  assign N4721 = N4720 | data_masked[6860];
  assign N4720 = N4719 | data_masked[6988];
  assign N4719 = N4718 | data_masked[7116];
  assign N4718 = N4717 | data_masked[7244];
  assign N4717 = N4716 | data_masked[7372];
  assign N4716 = N4715 | data_masked[7500];
  assign N4715 = N4714 | data_masked[7628];
  assign N4714 = N4713 | data_masked[7756];
  assign N4713 = N4712 | data_masked[7884];
  assign N4712 = data_masked[8140] | data_masked[8012];
  assign data_o[77] = N4835 | data_masked[77];
  assign N4835 = N4834 | data_masked[205];
  assign N4834 = N4833 | data_masked[333];
  assign N4833 = N4832 | data_masked[461];
  assign N4832 = N4831 | data_masked[589];
  assign N4831 = N4830 | data_masked[717];
  assign N4830 = N4829 | data_masked[845];
  assign N4829 = N4828 | data_masked[973];
  assign N4828 = N4827 | data_masked[1101];
  assign N4827 = N4826 | data_masked[1229];
  assign N4826 = N4825 | data_masked[1357];
  assign N4825 = N4824 | data_masked[1485];
  assign N4824 = N4823 | data_masked[1613];
  assign N4823 = N4822 | data_masked[1741];
  assign N4822 = N4821 | data_masked[1869];
  assign N4821 = N4820 | data_masked[1997];
  assign N4820 = N4819 | data_masked[2125];
  assign N4819 = N4818 | data_masked[2253];
  assign N4818 = N4817 | data_masked[2381];
  assign N4817 = N4816 | data_masked[2509];
  assign N4816 = N4815 | data_masked[2637];
  assign N4815 = N4814 | data_masked[2765];
  assign N4814 = N4813 | data_masked[2893];
  assign N4813 = N4812 | data_masked[3021];
  assign N4812 = N4811 | data_masked[3149];
  assign N4811 = N4810 | data_masked[3277];
  assign N4810 = N4809 | data_masked[3405];
  assign N4809 = N4808 | data_masked[3533];
  assign N4808 = N4807 | data_masked[3661];
  assign N4807 = N4806 | data_masked[3789];
  assign N4806 = N4805 | data_masked[3917];
  assign N4805 = N4804 | data_masked[4045];
  assign N4804 = N4803 | data_masked[4173];
  assign N4803 = N4802 | data_masked[4301];
  assign N4802 = N4801 | data_masked[4429];
  assign N4801 = N4800 | data_masked[4557];
  assign N4800 = N4799 | data_masked[4685];
  assign N4799 = N4798 | data_masked[4813];
  assign N4798 = N4797 | data_masked[4941];
  assign N4797 = N4796 | data_masked[5069];
  assign N4796 = N4795 | data_masked[5197];
  assign N4795 = N4794 | data_masked[5325];
  assign N4794 = N4793 | data_masked[5453];
  assign N4793 = N4792 | data_masked[5581];
  assign N4792 = N4791 | data_masked[5709];
  assign N4791 = N4790 | data_masked[5837];
  assign N4790 = N4789 | data_masked[5965];
  assign N4789 = N4788 | data_masked[6093];
  assign N4788 = N4787 | data_masked[6221];
  assign N4787 = N4786 | data_masked[6349];
  assign N4786 = N4785 | data_masked[6477];
  assign N4785 = N4784 | data_masked[6605];
  assign N4784 = N4783 | data_masked[6733];
  assign N4783 = N4782 | data_masked[6861];
  assign N4782 = N4781 | data_masked[6989];
  assign N4781 = N4780 | data_masked[7117];
  assign N4780 = N4779 | data_masked[7245];
  assign N4779 = N4778 | data_masked[7373];
  assign N4778 = N4777 | data_masked[7501];
  assign N4777 = N4776 | data_masked[7629];
  assign N4776 = N4775 | data_masked[7757];
  assign N4775 = N4774 | data_masked[7885];
  assign N4774 = data_masked[8141] | data_masked[8013];
  assign data_o[78] = N4897 | data_masked[78];
  assign N4897 = N4896 | data_masked[206];
  assign N4896 = N4895 | data_masked[334];
  assign N4895 = N4894 | data_masked[462];
  assign N4894 = N4893 | data_masked[590];
  assign N4893 = N4892 | data_masked[718];
  assign N4892 = N4891 | data_masked[846];
  assign N4891 = N4890 | data_masked[974];
  assign N4890 = N4889 | data_masked[1102];
  assign N4889 = N4888 | data_masked[1230];
  assign N4888 = N4887 | data_masked[1358];
  assign N4887 = N4886 | data_masked[1486];
  assign N4886 = N4885 | data_masked[1614];
  assign N4885 = N4884 | data_masked[1742];
  assign N4884 = N4883 | data_masked[1870];
  assign N4883 = N4882 | data_masked[1998];
  assign N4882 = N4881 | data_masked[2126];
  assign N4881 = N4880 | data_masked[2254];
  assign N4880 = N4879 | data_masked[2382];
  assign N4879 = N4878 | data_masked[2510];
  assign N4878 = N4877 | data_masked[2638];
  assign N4877 = N4876 | data_masked[2766];
  assign N4876 = N4875 | data_masked[2894];
  assign N4875 = N4874 | data_masked[3022];
  assign N4874 = N4873 | data_masked[3150];
  assign N4873 = N4872 | data_masked[3278];
  assign N4872 = N4871 | data_masked[3406];
  assign N4871 = N4870 | data_masked[3534];
  assign N4870 = N4869 | data_masked[3662];
  assign N4869 = N4868 | data_masked[3790];
  assign N4868 = N4867 | data_masked[3918];
  assign N4867 = N4866 | data_masked[4046];
  assign N4866 = N4865 | data_masked[4174];
  assign N4865 = N4864 | data_masked[4302];
  assign N4864 = N4863 | data_masked[4430];
  assign N4863 = N4862 | data_masked[4558];
  assign N4862 = N4861 | data_masked[4686];
  assign N4861 = N4860 | data_masked[4814];
  assign N4860 = N4859 | data_masked[4942];
  assign N4859 = N4858 | data_masked[5070];
  assign N4858 = N4857 | data_masked[5198];
  assign N4857 = N4856 | data_masked[5326];
  assign N4856 = N4855 | data_masked[5454];
  assign N4855 = N4854 | data_masked[5582];
  assign N4854 = N4853 | data_masked[5710];
  assign N4853 = N4852 | data_masked[5838];
  assign N4852 = N4851 | data_masked[5966];
  assign N4851 = N4850 | data_masked[6094];
  assign N4850 = N4849 | data_masked[6222];
  assign N4849 = N4848 | data_masked[6350];
  assign N4848 = N4847 | data_masked[6478];
  assign N4847 = N4846 | data_masked[6606];
  assign N4846 = N4845 | data_masked[6734];
  assign N4845 = N4844 | data_masked[6862];
  assign N4844 = N4843 | data_masked[6990];
  assign N4843 = N4842 | data_masked[7118];
  assign N4842 = N4841 | data_masked[7246];
  assign N4841 = N4840 | data_masked[7374];
  assign N4840 = N4839 | data_masked[7502];
  assign N4839 = N4838 | data_masked[7630];
  assign N4838 = N4837 | data_masked[7758];
  assign N4837 = N4836 | data_masked[7886];
  assign N4836 = data_masked[8142] | data_masked[8014];
  assign data_o[79] = N4959 | data_masked[79];
  assign N4959 = N4958 | data_masked[207];
  assign N4958 = N4957 | data_masked[335];
  assign N4957 = N4956 | data_masked[463];
  assign N4956 = N4955 | data_masked[591];
  assign N4955 = N4954 | data_masked[719];
  assign N4954 = N4953 | data_masked[847];
  assign N4953 = N4952 | data_masked[975];
  assign N4952 = N4951 | data_masked[1103];
  assign N4951 = N4950 | data_masked[1231];
  assign N4950 = N4949 | data_masked[1359];
  assign N4949 = N4948 | data_masked[1487];
  assign N4948 = N4947 | data_masked[1615];
  assign N4947 = N4946 | data_masked[1743];
  assign N4946 = N4945 | data_masked[1871];
  assign N4945 = N4944 | data_masked[1999];
  assign N4944 = N4943 | data_masked[2127];
  assign N4943 = N4942 | data_masked[2255];
  assign N4942 = N4941 | data_masked[2383];
  assign N4941 = N4940 | data_masked[2511];
  assign N4940 = N4939 | data_masked[2639];
  assign N4939 = N4938 | data_masked[2767];
  assign N4938 = N4937 | data_masked[2895];
  assign N4937 = N4936 | data_masked[3023];
  assign N4936 = N4935 | data_masked[3151];
  assign N4935 = N4934 | data_masked[3279];
  assign N4934 = N4933 | data_masked[3407];
  assign N4933 = N4932 | data_masked[3535];
  assign N4932 = N4931 | data_masked[3663];
  assign N4931 = N4930 | data_masked[3791];
  assign N4930 = N4929 | data_masked[3919];
  assign N4929 = N4928 | data_masked[4047];
  assign N4928 = N4927 | data_masked[4175];
  assign N4927 = N4926 | data_masked[4303];
  assign N4926 = N4925 | data_masked[4431];
  assign N4925 = N4924 | data_masked[4559];
  assign N4924 = N4923 | data_masked[4687];
  assign N4923 = N4922 | data_masked[4815];
  assign N4922 = N4921 | data_masked[4943];
  assign N4921 = N4920 | data_masked[5071];
  assign N4920 = N4919 | data_masked[5199];
  assign N4919 = N4918 | data_masked[5327];
  assign N4918 = N4917 | data_masked[5455];
  assign N4917 = N4916 | data_masked[5583];
  assign N4916 = N4915 | data_masked[5711];
  assign N4915 = N4914 | data_masked[5839];
  assign N4914 = N4913 | data_masked[5967];
  assign N4913 = N4912 | data_masked[6095];
  assign N4912 = N4911 | data_masked[6223];
  assign N4911 = N4910 | data_masked[6351];
  assign N4910 = N4909 | data_masked[6479];
  assign N4909 = N4908 | data_masked[6607];
  assign N4908 = N4907 | data_masked[6735];
  assign N4907 = N4906 | data_masked[6863];
  assign N4906 = N4905 | data_masked[6991];
  assign N4905 = N4904 | data_masked[7119];
  assign N4904 = N4903 | data_masked[7247];
  assign N4903 = N4902 | data_masked[7375];
  assign N4902 = N4901 | data_masked[7503];
  assign N4901 = N4900 | data_masked[7631];
  assign N4900 = N4899 | data_masked[7759];
  assign N4899 = N4898 | data_masked[7887];
  assign N4898 = data_masked[8143] | data_masked[8015];
  assign data_o[80] = N5021 | data_masked[80];
  assign N5021 = N5020 | data_masked[208];
  assign N5020 = N5019 | data_masked[336];
  assign N5019 = N5018 | data_masked[464];
  assign N5018 = N5017 | data_masked[592];
  assign N5017 = N5016 | data_masked[720];
  assign N5016 = N5015 | data_masked[848];
  assign N5015 = N5014 | data_masked[976];
  assign N5014 = N5013 | data_masked[1104];
  assign N5013 = N5012 | data_masked[1232];
  assign N5012 = N5011 | data_masked[1360];
  assign N5011 = N5010 | data_masked[1488];
  assign N5010 = N5009 | data_masked[1616];
  assign N5009 = N5008 | data_masked[1744];
  assign N5008 = N5007 | data_masked[1872];
  assign N5007 = N5006 | data_masked[2000];
  assign N5006 = N5005 | data_masked[2128];
  assign N5005 = N5004 | data_masked[2256];
  assign N5004 = N5003 | data_masked[2384];
  assign N5003 = N5002 | data_masked[2512];
  assign N5002 = N5001 | data_masked[2640];
  assign N5001 = N5000 | data_masked[2768];
  assign N5000 = N4999 | data_masked[2896];
  assign N4999 = N4998 | data_masked[3024];
  assign N4998 = N4997 | data_masked[3152];
  assign N4997 = N4996 | data_masked[3280];
  assign N4996 = N4995 | data_masked[3408];
  assign N4995 = N4994 | data_masked[3536];
  assign N4994 = N4993 | data_masked[3664];
  assign N4993 = N4992 | data_masked[3792];
  assign N4992 = N4991 | data_masked[3920];
  assign N4991 = N4990 | data_masked[4048];
  assign N4990 = N4989 | data_masked[4176];
  assign N4989 = N4988 | data_masked[4304];
  assign N4988 = N4987 | data_masked[4432];
  assign N4987 = N4986 | data_masked[4560];
  assign N4986 = N4985 | data_masked[4688];
  assign N4985 = N4984 | data_masked[4816];
  assign N4984 = N4983 | data_masked[4944];
  assign N4983 = N4982 | data_masked[5072];
  assign N4982 = N4981 | data_masked[5200];
  assign N4981 = N4980 | data_masked[5328];
  assign N4980 = N4979 | data_masked[5456];
  assign N4979 = N4978 | data_masked[5584];
  assign N4978 = N4977 | data_masked[5712];
  assign N4977 = N4976 | data_masked[5840];
  assign N4976 = N4975 | data_masked[5968];
  assign N4975 = N4974 | data_masked[6096];
  assign N4974 = N4973 | data_masked[6224];
  assign N4973 = N4972 | data_masked[6352];
  assign N4972 = N4971 | data_masked[6480];
  assign N4971 = N4970 | data_masked[6608];
  assign N4970 = N4969 | data_masked[6736];
  assign N4969 = N4968 | data_masked[6864];
  assign N4968 = N4967 | data_masked[6992];
  assign N4967 = N4966 | data_masked[7120];
  assign N4966 = N4965 | data_masked[7248];
  assign N4965 = N4964 | data_masked[7376];
  assign N4964 = N4963 | data_masked[7504];
  assign N4963 = N4962 | data_masked[7632];
  assign N4962 = N4961 | data_masked[7760];
  assign N4961 = N4960 | data_masked[7888];
  assign N4960 = data_masked[8144] | data_masked[8016];
  assign data_o[81] = N5083 | data_masked[81];
  assign N5083 = N5082 | data_masked[209];
  assign N5082 = N5081 | data_masked[337];
  assign N5081 = N5080 | data_masked[465];
  assign N5080 = N5079 | data_masked[593];
  assign N5079 = N5078 | data_masked[721];
  assign N5078 = N5077 | data_masked[849];
  assign N5077 = N5076 | data_masked[977];
  assign N5076 = N5075 | data_masked[1105];
  assign N5075 = N5074 | data_masked[1233];
  assign N5074 = N5073 | data_masked[1361];
  assign N5073 = N5072 | data_masked[1489];
  assign N5072 = N5071 | data_masked[1617];
  assign N5071 = N5070 | data_masked[1745];
  assign N5070 = N5069 | data_masked[1873];
  assign N5069 = N5068 | data_masked[2001];
  assign N5068 = N5067 | data_masked[2129];
  assign N5067 = N5066 | data_masked[2257];
  assign N5066 = N5065 | data_masked[2385];
  assign N5065 = N5064 | data_masked[2513];
  assign N5064 = N5063 | data_masked[2641];
  assign N5063 = N5062 | data_masked[2769];
  assign N5062 = N5061 | data_masked[2897];
  assign N5061 = N5060 | data_masked[3025];
  assign N5060 = N5059 | data_masked[3153];
  assign N5059 = N5058 | data_masked[3281];
  assign N5058 = N5057 | data_masked[3409];
  assign N5057 = N5056 | data_masked[3537];
  assign N5056 = N5055 | data_masked[3665];
  assign N5055 = N5054 | data_masked[3793];
  assign N5054 = N5053 | data_masked[3921];
  assign N5053 = N5052 | data_masked[4049];
  assign N5052 = N5051 | data_masked[4177];
  assign N5051 = N5050 | data_masked[4305];
  assign N5050 = N5049 | data_masked[4433];
  assign N5049 = N5048 | data_masked[4561];
  assign N5048 = N5047 | data_masked[4689];
  assign N5047 = N5046 | data_masked[4817];
  assign N5046 = N5045 | data_masked[4945];
  assign N5045 = N5044 | data_masked[5073];
  assign N5044 = N5043 | data_masked[5201];
  assign N5043 = N5042 | data_masked[5329];
  assign N5042 = N5041 | data_masked[5457];
  assign N5041 = N5040 | data_masked[5585];
  assign N5040 = N5039 | data_masked[5713];
  assign N5039 = N5038 | data_masked[5841];
  assign N5038 = N5037 | data_masked[5969];
  assign N5037 = N5036 | data_masked[6097];
  assign N5036 = N5035 | data_masked[6225];
  assign N5035 = N5034 | data_masked[6353];
  assign N5034 = N5033 | data_masked[6481];
  assign N5033 = N5032 | data_masked[6609];
  assign N5032 = N5031 | data_masked[6737];
  assign N5031 = N5030 | data_masked[6865];
  assign N5030 = N5029 | data_masked[6993];
  assign N5029 = N5028 | data_masked[7121];
  assign N5028 = N5027 | data_masked[7249];
  assign N5027 = N5026 | data_masked[7377];
  assign N5026 = N5025 | data_masked[7505];
  assign N5025 = N5024 | data_masked[7633];
  assign N5024 = N5023 | data_masked[7761];
  assign N5023 = N5022 | data_masked[7889];
  assign N5022 = data_masked[8145] | data_masked[8017];
  assign data_o[82] = N5145 | data_masked[82];
  assign N5145 = N5144 | data_masked[210];
  assign N5144 = N5143 | data_masked[338];
  assign N5143 = N5142 | data_masked[466];
  assign N5142 = N5141 | data_masked[594];
  assign N5141 = N5140 | data_masked[722];
  assign N5140 = N5139 | data_masked[850];
  assign N5139 = N5138 | data_masked[978];
  assign N5138 = N5137 | data_masked[1106];
  assign N5137 = N5136 | data_masked[1234];
  assign N5136 = N5135 | data_masked[1362];
  assign N5135 = N5134 | data_masked[1490];
  assign N5134 = N5133 | data_masked[1618];
  assign N5133 = N5132 | data_masked[1746];
  assign N5132 = N5131 | data_masked[1874];
  assign N5131 = N5130 | data_masked[2002];
  assign N5130 = N5129 | data_masked[2130];
  assign N5129 = N5128 | data_masked[2258];
  assign N5128 = N5127 | data_masked[2386];
  assign N5127 = N5126 | data_masked[2514];
  assign N5126 = N5125 | data_masked[2642];
  assign N5125 = N5124 | data_masked[2770];
  assign N5124 = N5123 | data_masked[2898];
  assign N5123 = N5122 | data_masked[3026];
  assign N5122 = N5121 | data_masked[3154];
  assign N5121 = N5120 | data_masked[3282];
  assign N5120 = N5119 | data_masked[3410];
  assign N5119 = N5118 | data_masked[3538];
  assign N5118 = N5117 | data_masked[3666];
  assign N5117 = N5116 | data_masked[3794];
  assign N5116 = N5115 | data_masked[3922];
  assign N5115 = N5114 | data_masked[4050];
  assign N5114 = N5113 | data_masked[4178];
  assign N5113 = N5112 | data_masked[4306];
  assign N5112 = N5111 | data_masked[4434];
  assign N5111 = N5110 | data_masked[4562];
  assign N5110 = N5109 | data_masked[4690];
  assign N5109 = N5108 | data_masked[4818];
  assign N5108 = N5107 | data_masked[4946];
  assign N5107 = N5106 | data_masked[5074];
  assign N5106 = N5105 | data_masked[5202];
  assign N5105 = N5104 | data_masked[5330];
  assign N5104 = N5103 | data_masked[5458];
  assign N5103 = N5102 | data_masked[5586];
  assign N5102 = N5101 | data_masked[5714];
  assign N5101 = N5100 | data_masked[5842];
  assign N5100 = N5099 | data_masked[5970];
  assign N5099 = N5098 | data_masked[6098];
  assign N5098 = N5097 | data_masked[6226];
  assign N5097 = N5096 | data_masked[6354];
  assign N5096 = N5095 | data_masked[6482];
  assign N5095 = N5094 | data_masked[6610];
  assign N5094 = N5093 | data_masked[6738];
  assign N5093 = N5092 | data_masked[6866];
  assign N5092 = N5091 | data_masked[6994];
  assign N5091 = N5090 | data_masked[7122];
  assign N5090 = N5089 | data_masked[7250];
  assign N5089 = N5088 | data_masked[7378];
  assign N5088 = N5087 | data_masked[7506];
  assign N5087 = N5086 | data_masked[7634];
  assign N5086 = N5085 | data_masked[7762];
  assign N5085 = N5084 | data_masked[7890];
  assign N5084 = data_masked[8146] | data_masked[8018];
  assign data_o[83] = N5207 | data_masked[83];
  assign N5207 = N5206 | data_masked[211];
  assign N5206 = N5205 | data_masked[339];
  assign N5205 = N5204 | data_masked[467];
  assign N5204 = N5203 | data_masked[595];
  assign N5203 = N5202 | data_masked[723];
  assign N5202 = N5201 | data_masked[851];
  assign N5201 = N5200 | data_masked[979];
  assign N5200 = N5199 | data_masked[1107];
  assign N5199 = N5198 | data_masked[1235];
  assign N5198 = N5197 | data_masked[1363];
  assign N5197 = N5196 | data_masked[1491];
  assign N5196 = N5195 | data_masked[1619];
  assign N5195 = N5194 | data_masked[1747];
  assign N5194 = N5193 | data_masked[1875];
  assign N5193 = N5192 | data_masked[2003];
  assign N5192 = N5191 | data_masked[2131];
  assign N5191 = N5190 | data_masked[2259];
  assign N5190 = N5189 | data_masked[2387];
  assign N5189 = N5188 | data_masked[2515];
  assign N5188 = N5187 | data_masked[2643];
  assign N5187 = N5186 | data_masked[2771];
  assign N5186 = N5185 | data_masked[2899];
  assign N5185 = N5184 | data_masked[3027];
  assign N5184 = N5183 | data_masked[3155];
  assign N5183 = N5182 | data_masked[3283];
  assign N5182 = N5181 | data_masked[3411];
  assign N5181 = N5180 | data_masked[3539];
  assign N5180 = N5179 | data_masked[3667];
  assign N5179 = N5178 | data_masked[3795];
  assign N5178 = N5177 | data_masked[3923];
  assign N5177 = N5176 | data_masked[4051];
  assign N5176 = N5175 | data_masked[4179];
  assign N5175 = N5174 | data_masked[4307];
  assign N5174 = N5173 | data_masked[4435];
  assign N5173 = N5172 | data_masked[4563];
  assign N5172 = N5171 | data_masked[4691];
  assign N5171 = N5170 | data_masked[4819];
  assign N5170 = N5169 | data_masked[4947];
  assign N5169 = N5168 | data_masked[5075];
  assign N5168 = N5167 | data_masked[5203];
  assign N5167 = N5166 | data_masked[5331];
  assign N5166 = N5165 | data_masked[5459];
  assign N5165 = N5164 | data_masked[5587];
  assign N5164 = N5163 | data_masked[5715];
  assign N5163 = N5162 | data_masked[5843];
  assign N5162 = N5161 | data_masked[5971];
  assign N5161 = N5160 | data_masked[6099];
  assign N5160 = N5159 | data_masked[6227];
  assign N5159 = N5158 | data_masked[6355];
  assign N5158 = N5157 | data_masked[6483];
  assign N5157 = N5156 | data_masked[6611];
  assign N5156 = N5155 | data_masked[6739];
  assign N5155 = N5154 | data_masked[6867];
  assign N5154 = N5153 | data_masked[6995];
  assign N5153 = N5152 | data_masked[7123];
  assign N5152 = N5151 | data_masked[7251];
  assign N5151 = N5150 | data_masked[7379];
  assign N5150 = N5149 | data_masked[7507];
  assign N5149 = N5148 | data_masked[7635];
  assign N5148 = N5147 | data_masked[7763];
  assign N5147 = N5146 | data_masked[7891];
  assign N5146 = data_masked[8147] | data_masked[8019];
  assign data_o[84] = N5269 | data_masked[84];
  assign N5269 = N5268 | data_masked[212];
  assign N5268 = N5267 | data_masked[340];
  assign N5267 = N5266 | data_masked[468];
  assign N5266 = N5265 | data_masked[596];
  assign N5265 = N5264 | data_masked[724];
  assign N5264 = N5263 | data_masked[852];
  assign N5263 = N5262 | data_masked[980];
  assign N5262 = N5261 | data_masked[1108];
  assign N5261 = N5260 | data_masked[1236];
  assign N5260 = N5259 | data_masked[1364];
  assign N5259 = N5258 | data_masked[1492];
  assign N5258 = N5257 | data_masked[1620];
  assign N5257 = N5256 | data_masked[1748];
  assign N5256 = N5255 | data_masked[1876];
  assign N5255 = N5254 | data_masked[2004];
  assign N5254 = N5253 | data_masked[2132];
  assign N5253 = N5252 | data_masked[2260];
  assign N5252 = N5251 | data_masked[2388];
  assign N5251 = N5250 | data_masked[2516];
  assign N5250 = N5249 | data_masked[2644];
  assign N5249 = N5248 | data_masked[2772];
  assign N5248 = N5247 | data_masked[2900];
  assign N5247 = N5246 | data_masked[3028];
  assign N5246 = N5245 | data_masked[3156];
  assign N5245 = N5244 | data_masked[3284];
  assign N5244 = N5243 | data_masked[3412];
  assign N5243 = N5242 | data_masked[3540];
  assign N5242 = N5241 | data_masked[3668];
  assign N5241 = N5240 | data_masked[3796];
  assign N5240 = N5239 | data_masked[3924];
  assign N5239 = N5238 | data_masked[4052];
  assign N5238 = N5237 | data_masked[4180];
  assign N5237 = N5236 | data_masked[4308];
  assign N5236 = N5235 | data_masked[4436];
  assign N5235 = N5234 | data_masked[4564];
  assign N5234 = N5233 | data_masked[4692];
  assign N5233 = N5232 | data_masked[4820];
  assign N5232 = N5231 | data_masked[4948];
  assign N5231 = N5230 | data_masked[5076];
  assign N5230 = N5229 | data_masked[5204];
  assign N5229 = N5228 | data_masked[5332];
  assign N5228 = N5227 | data_masked[5460];
  assign N5227 = N5226 | data_masked[5588];
  assign N5226 = N5225 | data_masked[5716];
  assign N5225 = N5224 | data_masked[5844];
  assign N5224 = N5223 | data_masked[5972];
  assign N5223 = N5222 | data_masked[6100];
  assign N5222 = N5221 | data_masked[6228];
  assign N5221 = N5220 | data_masked[6356];
  assign N5220 = N5219 | data_masked[6484];
  assign N5219 = N5218 | data_masked[6612];
  assign N5218 = N5217 | data_masked[6740];
  assign N5217 = N5216 | data_masked[6868];
  assign N5216 = N5215 | data_masked[6996];
  assign N5215 = N5214 | data_masked[7124];
  assign N5214 = N5213 | data_masked[7252];
  assign N5213 = N5212 | data_masked[7380];
  assign N5212 = N5211 | data_masked[7508];
  assign N5211 = N5210 | data_masked[7636];
  assign N5210 = N5209 | data_masked[7764];
  assign N5209 = N5208 | data_masked[7892];
  assign N5208 = data_masked[8148] | data_masked[8020];
  assign data_o[85] = N5331 | data_masked[85];
  assign N5331 = N5330 | data_masked[213];
  assign N5330 = N5329 | data_masked[341];
  assign N5329 = N5328 | data_masked[469];
  assign N5328 = N5327 | data_masked[597];
  assign N5327 = N5326 | data_masked[725];
  assign N5326 = N5325 | data_masked[853];
  assign N5325 = N5324 | data_masked[981];
  assign N5324 = N5323 | data_masked[1109];
  assign N5323 = N5322 | data_masked[1237];
  assign N5322 = N5321 | data_masked[1365];
  assign N5321 = N5320 | data_masked[1493];
  assign N5320 = N5319 | data_masked[1621];
  assign N5319 = N5318 | data_masked[1749];
  assign N5318 = N5317 | data_masked[1877];
  assign N5317 = N5316 | data_masked[2005];
  assign N5316 = N5315 | data_masked[2133];
  assign N5315 = N5314 | data_masked[2261];
  assign N5314 = N5313 | data_masked[2389];
  assign N5313 = N5312 | data_masked[2517];
  assign N5312 = N5311 | data_masked[2645];
  assign N5311 = N5310 | data_masked[2773];
  assign N5310 = N5309 | data_masked[2901];
  assign N5309 = N5308 | data_masked[3029];
  assign N5308 = N5307 | data_masked[3157];
  assign N5307 = N5306 | data_masked[3285];
  assign N5306 = N5305 | data_masked[3413];
  assign N5305 = N5304 | data_masked[3541];
  assign N5304 = N5303 | data_masked[3669];
  assign N5303 = N5302 | data_masked[3797];
  assign N5302 = N5301 | data_masked[3925];
  assign N5301 = N5300 | data_masked[4053];
  assign N5300 = N5299 | data_masked[4181];
  assign N5299 = N5298 | data_masked[4309];
  assign N5298 = N5297 | data_masked[4437];
  assign N5297 = N5296 | data_masked[4565];
  assign N5296 = N5295 | data_masked[4693];
  assign N5295 = N5294 | data_masked[4821];
  assign N5294 = N5293 | data_masked[4949];
  assign N5293 = N5292 | data_masked[5077];
  assign N5292 = N5291 | data_masked[5205];
  assign N5291 = N5290 | data_masked[5333];
  assign N5290 = N5289 | data_masked[5461];
  assign N5289 = N5288 | data_masked[5589];
  assign N5288 = N5287 | data_masked[5717];
  assign N5287 = N5286 | data_masked[5845];
  assign N5286 = N5285 | data_masked[5973];
  assign N5285 = N5284 | data_masked[6101];
  assign N5284 = N5283 | data_masked[6229];
  assign N5283 = N5282 | data_masked[6357];
  assign N5282 = N5281 | data_masked[6485];
  assign N5281 = N5280 | data_masked[6613];
  assign N5280 = N5279 | data_masked[6741];
  assign N5279 = N5278 | data_masked[6869];
  assign N5278 = N5277 | data_masked[6997];
  assign N5277 = N5276 | data_masked[7125];
  assign N5276 = N5275 | data_masked[7253];
  assign N5275 = N5274 | data_masked[7381];
  assign N5274 = N5273 | data_masked[7509];
  assign N5273 = N5272 | data_masked[7637];
  assign N5272 = N5271 | data_masked[7765];
  assign N5271 = N5270 | data_masked[7893];
  assign N5270 = data_masked[8149] | data_masked[8021];
  assign data_o[86] = N5393 | data_masked[86];
  assign N5393 = N5392 | data_masked[214];
  assign N5392 = N5391 | data_masked[342];
  assign N5391 = N5390 | data_masked[470];
  assign N5390 = N5389 | data_masked[598];
  assign N5389 = N5388 | data_masked[726];
  assign N5388 = N5387 | data_masked[854];
  assign N5387 = N5386 | data_masked[982];
  assign N5386 = N5385 | data_masked[1110];
  assign N5385 = N5384 | data_masked[1238];
  assign N5384 = N5383 | data_masked[1366];
  assign N5383 = N5382 | data_masked[1494];
  assign N5382 = N5381 | data_masked[1622];
  assign N5381 = N5380 | data_masked[1750];
  assign N5380 = N5379 | data_masked[1878];
  assign N5379 = N5378 | data_masked[2006];
  assign N5378 = N5377 | data_masked[2134];
  assign N5377 = N5376 | data_masked[2262];
  assign N5376 = N5375 | data_masked[2390];
  assign N5375 = N5374 | data_masked[2518];
  assign N5374 = N5373 | data_masked[2646];
  assign N5373 = N5372 | data_masked[2774];
  assign N5372 = N5371 | data_masked[2902];
  assign N5371 = N5370 | data_masked[3030];
  assign N5370 = N5369 | data_masked[3158];
  assign N5369 = N5368 | data_masked[3286];
  assign N5368 = N5367 | data_masked[3414];
  assign N5367 = N5366 | data_masked[3542];
  assign N5366 = N5365 | data_masked[3670];
  assign N5365 = N5364 | data_masked[3798];
  assign N5364 = N5363 | data_masked[3926];
  assign N5363 = N5362 | data_masked[4054];
  assign N5362 = N5361 | data_masked[4182];
  assign N5361 = N5360 | data_masked[4310];
  assign N5360 = N5359 | data_masked[4438];
  assign N5359 = N5358 | data_masked[4566];
  assign N5358 = N5357 | data_masked[4694];
  assign N5357 = N5356 | data_masked[4822];
  assign N5356 = N5355 | data_masked[4950];
  assign N5355 = N5354 | data_masked[5078];
  assign N5354 = N5353 | data_masked[5206];
  assign N5353 = N5352 | data_masked[5334];
  assign N5352 = N5351 | data_masked[5462];
  assign N5351 = N5350 | data_masked[5590];
  assign N5350 = N5349 | data_masked[5718];
  assign N5349 = N5348 | data_masked[5846];
  assign N5348 = N5347 | data_masked[5974];
  assign N5347 = N5346 | data_masked[6102];
  assign N5346 = N5345 | data_masked[6230];
  assign N5345 = N5344 | data_masked[6358];
  assign N5344 = N5343 | data_masked[6486];
  assign N5343 = N5342 | data_masked[6614];
  assign N5342 = N5341 | data_masked[6742];
  assign N5341 = N5340 | data_masked[6870];
  assign N5340 = N5339 | data_masked[6998];
  assign N5339 = N5338 | data_masked[7126];
  assign N5338 = N5337 | data_masked[7254];
  assign N5337 = N5336 | data_masked[7382];
  assign N5336 = N5335 | data_masked[7510];
  assign N5335 = N5334 | data_masked[7638];
  assign N5334 = N5333 | data_masked[7766];
  assign N5333 = N5332 | data_masked[7894];
  assign N5332 = data_masked[8150] | data_masked[8022];
  assign data_o[87] = N5455 | data_masked[87];
  assign N5455 = N5454 | data_masked[215];
  assign N5454 = N5453 | data_masked[343];
  assign N5453 = N5452 | data_masked[471];
  assign N5452 = N5451 | data_masked[599];
  assign N5451 = N5450 | data_masked[727];
  assign N5450 = N5449 | data_masked[855];
  assign N5449 = N5448 | data_masked[983];
  assign N5448 = N5447 | data_masked[1111];
  assign N5447 = N5446 | data_masked[1239];
  assign N5446 = N5445 | data_masked[1367];
  assign N5445 = N5444 | data_masked[1495];
  assign N5444 = N5443 | data_masked[1623];
  assign N5443 = N5442 | data_masked[1751];
  assign N5442 = N5441 | data_masked[1879];
  assign N5441 = N5440 | data_masked[2007];
  assign N5440 = N5439 | data_masked[2135];
  assign N5439 = N5438 | data_masked[2263];
  assign N5438 = N5437 | data_masked[2391];
  assign N5437 = N5436 | data_masked[2519];
  assign N5436 = N5435 | data_masked[2647];
  assign N5435 = N5434 | data_masked[2775];
  assign N5434 = N5433 | data_masked[2903];
  assign N5433 = N5432 | data_masked[3031];
  assign N5432 = N5431 | data_masked[3159];
  assign N5431 = N5430 | data_masked[3287];
  assign N5430 = N5429 | data_masked[3415];
  assign N5429 = N5428 | data_masked[3543];
  assign N5428 = N5427 | data_masked[3671];
  assign N5427 = N5426 | data_masked[3799];
  assign N5426 = N5425 | data_masked[3927];
  assign N5425 = N5424 | data_masked[4055];
  assign N5424 = N5423 | data_masked[4183];
  assign N5423 = N5422 | data_masked[4311];
  assign N5422 = N5421 | data_masked[4439];
  assign N5421 = N5420 | data_masked[4567];
  assign N5420 = N5419 | data_masked[4695];
  assign N5419 = N5418 | data_masked[4823];
  assign N5418 = N5417 | data_masked[4951];
  assign N5417 = N5416 | data_masked[5079];
  assign N5416 = N5415 | data_masked[5207];
  assign N5415 = N5414 | data_masked[5335];
  assign N5414 = N5413 | data_masked[5463];
  assign N5413 = N5412 | data_masked[5591];
  assign N5412 = N5411 | data_masked[5719];
  assign N5411 = N5410 | data_masked[5847];
  assign N5410 = N5409 | data_masked[5975];
  assign N5409 = N5408 | data_masked[6103];
  assign N5408 = N5407 | data_masked[6231];
  assign N5407 = N5406 | data_masked[6359];
  assign N5406 = N5405 | data_masked[6487];
  assign N5405 = N5404 | data_masked[6615];
  assign N5404 = N5403 | data_masked[6743];
  assign N5403 = N5402 | data_masked[6871];
  assign N5402 = N5401 | data_masked[6999];
  assign N5401 = N5400 | data_masked[7127];
  assign N5400 = N5399 | data_masked[7255];
  assign N5399 = N5398 | data_masked[7383];
  assign N5398 = N5397 | data_masked[7511];
  assign N5397 = N5396 | data_masked[7639];
  assign N5396 = N5395 | data_masked[7767];
  assign N5395 = N5394 | data_masked[7895];
  assign N5394 = data_masked[8151] | data_masked[8023];
  assign data_o[88] = N5517 | data_masked[88];
  assign N5517 = N5516 | data_masked[216];
  assign N5516 = N5515 | data_masked[344];
  assign N5515 = N5514 | data_masked[472];
  assign N5514 = N5513 | data_masked[600];
  assign N5513 = N5512 | data_masked[728];
  assign N5512 = N5511 | data_masked[856];
  assign N5511 = N5510 | data_masked[984];
  assign N5510 = N5509 | data_masked[1112];
  assign N5509 = N5508 | data_masked[1240];
  assign N5508 = N5507 | data_masked[1368];
  assign N5507 = N5506 | data_masked[1496];
  assign N5506 = N5505 | data_masked[1624];
  assign N5505 = N5504 | data_masked[1752];
  assign N5504 = N5503 | data_masked[1880];
  assign N5503 = N5502 | data_masked[2008];
  assign N5502 = N5501 | data_masked[2136];
  assign N5501 = N5500 | data_masked[2264];
  assign N5500 = N5499 | data_masked[2392];
  assign N5499 = N5498 | data_masked[2520];
  assign N5498 = N5497 | data_masked[2648];
  assign N5497 = N5496 | data_masked[2776];
  assign N5496 = N5495 | data_masked[2904];
  assign N5495 = N5494 | data_masked[3032];
  assign N5494 = N5493 | data_masked[3160];
  assign N5493 = N5492 | data_masked[3288];
  assign N5492 = N5491 | data_masked[3416];
  assign N5491 = N5490 | data_masked[3544];
  assign N5490 = N5489 | data_masked[3672];
  assign N5489 = N5488 | data_masked[3800];
  assign N5488 = N5487 | data_masked[3928];
  assign N5487 = N5486 | data_masked[4056];
  assign N5486 = N5485 | data_masked[4184];
  assign N5485 = N5484 | data_masked[4312];
  assign N5484 = N5483 | data_masked[4440];
  assign N5483 = N5482 | data_masked[4568];
  assign N5482 = N5481 | data_masked[4696];
  assign N5481 = N5480 | data_masked[4824];
  assign N5480 = N5479 | data_masked[4952];
  assign N5479 = N5478 | data_masked[5080];
  assign N5478 = N5477 | data_masked[5208];
  assign N5477 = N5476 | data_masked[5336];
  assign N5476 = N5475 | data_masked[5464];
  assign N5475 = N5474 | data_masked[5592];
  assign N5474 = N5473 | data_masked[5720];
  assign N5473 = N5472 | data_masked[5848];
  assign N5472 = N5471 | data_masked[5976];
  assign N5471 = N5470 | data_masked[6104];
  assign N5470 = N5469 | data_masked[6232];
  assign N5469 = N5468 | data_masked[6360];
  assign N5468 = N5467 | data_masked[6488];
  assign N5467 = N5466 | data_masked[6616];
  assign N5466 = N5465 | data_masked[6744];
  assign N5465 = N5464 | data_masked[6872];
  assign N5464 = N5463 | data_masked[7000];
  assign N5463 = N5462 | data_masked[7128];
  assign N5462 = N5461 | data_masked[7256];
  assign N5461 = N5460 | data_masked[7384];
  assign N5460 = N5459 | data_masked[7512];
  assign N5459 = N5458 | data_masked[7640];
  assign N5458 = N5457 | data_masked[7768];
  assign N5457 = N5456 | data_masked[7896];
  assign N5456 = data_masked[8152] | data_masked[8024];
  assign data_o[89] = N5579 | data_masked[89];
  assign N5579 = N5578 | data_masked[217];
  assign N5578 = N5577 | data_masked[345];
  assign N5577 = N5576 | data_masked[473];
  assign N5576 = N5575 | data_masked[601];
  assign N5575 = N5574 | data_masked[729];
  assign N5574 = N5573 | data_masked[857];
  assign N5573 = N5572 | data_masked[985];
  assign N5572 = N5571 | data_masked[1113];
  assign N5571 = N5570 | data_masked[1241];
  assign N5570 = N5569 | data_masked[1369];
  assign N5569 = N5568 | data_masked[1497];
  assign N5568 = N5567 | data_masked[1625];
  assign N5567 = N5566 | data_masked[1753];
  assign N5566 = N5565 | data_masked[1881];
  assign N5565 = N5564 | data_masked[2009];
  assign N5564 = N5563 | data_masked[2137];
  assign N5563 = N5562 | data_masked[2265];
  assign N5562 = N5561 | data_masked[2393];
  assign N5561 = N5560 | data_masked[2521];
  assign N5560 = N5559 | data_masked[2649];
  assign N5559 = N5558 | data_masked[2777];
  assign N5558 = N5557 | data_masked[2905];
  assign N5557 = N5556 | data_masked[3033];
  assign N5556 = N5555 | data_masked[3161];
  assign N5555 = N5554 | data_masked[3289];
  assign N5554 = N5553 | data_masked[3417];
  assign N5553 = N5552 | data_masked[3545];
  assign N5552 = N5551 | data_masked[3673];
  assign N5551 = N5550 | data_masked[3801];
  assign N5550 = N5549 | data_masked[3929];
  assign N5549 = N5548 | data_masked[4057];
  assign N5548 = N5547 | data_masked[4185];
  assign N5547 = N5546 | data_masked[4313];
  assign N5546 = N5545 | data_masked[4441];
  assign N5545 = N5544 | data_masked[4569];
  assign N5544 = N5543 | data_masked[4697];
  assign N5543 = N5542 | data_masked[4825];
  assign N5542 = N5541 | data_masked[4953];
  assign N5541 = N5540 | data_masked[5081];
  assign N5540 = N5539 | data_masked[5209];
  assign N5539 = N5538 | data_masked[5337];
  assign N5538 = N5537 | data_masked[5465];
  assign N5537 = N5536 | data_masked[5593];
  assign N5536 = N5535 | data_masked[5721];
  assign N5535 = N5534 | data_masked[5849];
  assign N5534 = N5533 | data_masked[5977];
  assign N5533 = N5532 | data_masked[6105];
  assign N5532 = N5531 | data_masked[6233];
  assign N5531 = N5530 | data_masked[6361];
  assign N5530 = N5529 | data_masked[6489];
  assign N5529 = N5528 | data_masked[6617];
  assign N5528 = N5527 | data_masked[6745];
  assign N5527 = N5526 | data_masked[6873];
  assign N5526 = N5525 | data_masked[7001];
  assign N5525 = N5524 | data_masked[7129];
  assign N5524 = N5523 | data_masked[7257];
  assign N5523 = N5522 | data_masked[7385];
  assign N5522 = N5521 | data_masked[7513];
  assign N5521 = N5520 | data_masked[7641];
  assign N5520 = N5519 | data_masked[7769];
  assign N5519 = N5518 | data_masked[7897];
  assign N5518 = data_masked[8153] | data_masked[8025];
  assign data_o[90] = N5641 | data_masked[90];
  assign N5641 = N5640 | data_masked[218];
  assign N5640 = N5639 | data_masked[346];
  assign N5639 = N5638 | data_masked[474];
  assign N5638 = N5637 | data_masked[602];
  assign N5637 = N5636 | data_masked[730];
  assign N5636 = N5635 | data_masked[858];
  assign N5635 = N5634 | data_masked[986];
  assign N5634 = N5633 | data_masked[1114];
  assign N5633 = N5632 | data_masked[1242];
  assign N5632 = N5631 | data_masked[1370];
  assign N5631 = N5630 | data_masked[1498];
  assign N5630 = N5629 | data_masked[1626];
  assign N5629 = N5628 | data_masked[1754];
  assign N5628 = N5627 | data_masked[1882];
  assign N5627 = N5626 | data_masked[2010];
  assign N5626 = N5625 | data_masked[2138];
  assign N5625 = N5624 | data_masked[2266];
  assign N5624 = N5623 | data_masked[2394];
  assign N5623 = N5622 | data_masked[2522];
  assign N5622 = N5621 | data_masked[2650];
  assign N5621 = N5620 | data_masked[2778];
  assign N5620 = N5619 | data_masked[2906];
  assign N5619 = N5618 | data_masked[3034];
  assign N5618 = N5617 | data_masked[3162];
  assign N5617 = N5616 | data_masked[3290];
  assign N5616 = N5615 | data_masked[3418];
  assign N5615 = N5614 | data_masked[3546];
  assign N5614 = N5613 | data_masked[3674];
  assign N5613 = N5612 | data_masked[3802];
  assign N5612 = N5611 | data_masked[3930];
  assign N5611 = N5610 | data_masked[4058];
  assign N5610 = N5609 | data_masked[4186];
  assign N5609 = N5608 | data_masked[4314];
  assign N5608 = N5607 | data_masked[4442];
  assign N5607 = N5606 | data_masked[4570];
  assign N5606 = N5605 | data_masked[4698];
  assign N5605 = N5604 | data_masked[4826];
  assign N5604 = N5603 | data_masked[4954];
  assign N5603 = N5602 | data_masked[5082];
  assign N5602 = N5601 | data_masked[5210];
  assign N5601 = N5600 | data_masked[5338];
  assign N5600 = N5599 | data_masked[5466];
  assign N5599 = N5598 | data_masked[5594];
  assign N5598 = N5597 | data_masked[5722];
  assign N5597 = N5596 | data_masked[5850];
  assign N5596 = N5595 | data_masked[5978];
  assign N5595 = N5594 | data_masked[6106];
  assign N5594 = N5593 | data_masked[6234];
  assign N5593 = N5592 | data_masked[6362];
  assign N5592 = N5591 | data_masked[6490];
  assign N5591 = N5590 | data_masked[6618];
  assign N5590 = N5589 | data_masked[6746];
  assign N5589 = N5588 | data_masked[6874];
  assign N5588 = N5587 | data_masked[7002];
  assign N5587 = N5586 | data_masked[7130];
  assign N5586 = N5585 | data_masked[7258];
  assign N5585 = N5584 | data_masked[7386];
  assign N5584 = N5583 | data_masked[7514];
  assign N5583 = N5582 | data_masked[7642];
  assign N5582 = N5581 | data_masked[7770];
  assign N5581 = N5580 | data_masked[7898];
  assign N5580 = data_masked[8154] | data_masked[8026];
  assign data_o[91] = N5703 | data_masked[91];
  assign N5703 = N5702 | data_masked[219];
  assign N5702 = N5701 | data_masked[347];
  assign N5701 = N5700 | data_masked[475];
  assign N5700 = N5699 | data_masked[603];
  assign N5699 = N5698 | data_masked[731];
  assign N5698 = N5697 | data_masked[859];
  assign N5697 = N5696 | data_masked[987];
  assign N5696 = N5695 | data_masked[1115];
  assign N5695 = N5694 | data_masked[1243];
  assign N5694 = N5693 | data_masked[1371];
  assign N5693 = N5692 | data_masked[1499];
  assign N5692 = N5691 | data_masked[1627];
  assign N5691 = N5690 | data_masked[1755];
  assign N5690 = N5689 | data_masked[1883];
  assign N5689 = N5688 | data_masked[2011];
  assign N5688 = N5687 | data_masked[2139];
  assign N5687 = N5686 | data_masked[2267];
  assign N5686 = N5685 | data_masked[2395];
  assign N5685 = N5684 | data_masked[2523];
  assign N5684 = N5683 | data_masked[2651];
  assign N5683 = N5682 | data_masked[2779];
  assign N5682 = N5681 | data_masked[2907];
  assign N5681 = N5680 | data_masked[3035];
  assign N5680 = N5679 | data_masked[3163];
  assign N5679 = N5678 | data_masked[3291];
  assign N5678 = N5677 | data_masked[3419];
  assign N5677 = N5676 | data_masked[3547];
  assign N5676 = N5675 | data_masked[3675];
  assign N5675 = N5674 | data_masked[3803];
  assign N5674 = N5673 | data_masked[3931];
  assign N5673 = N5672 | data_masked[4059];
  assign N5672 = N5671 | data_masked[4187];
  assign N5671 = N5670 | data_masked[4315];
  assign N5670 = N5669 | data_masked[4443];
  assign N5669 = N5668 | data_masked[4571];
  assign N5668 = N5667 | data_masked[4699];
  assign N5667 = N5666 | data_masked[4827];
  assign N5666 = N5665 | data_masked[4955];
  assign N5665 = N5664 | data_masked[5083];
  assign N5664 = N5663 | data_masked[5211];
  assign N5663 = N5662 | data_masked[5339];
  assign N5662 = N5661 | data_masked[5467];
  assign N5661 = N5660 | data_masked[5595];
  assign N5660 = N5659 | data_masked[5723];
  assign N5659 = N5658 | data_masked[5851];
  assign N5658 = N5657 | data_masked[5979];
  assign N5657 = N5656 | data_masked[6107];
  assign N5656 = N5655 | data_masked[6235];
  assign N5655 = N5654 | data_masked[6363];
  assign N5654 = N5653 | data_masked[6491];
  assign N5653 = N5652 | data_masked[6619];
  assign N5652 = N5651 | data_masked[6747];
  assign N5651 = N5650 | data_masked[6875];
  assign N5650 = N5649 | data_masked[7003];
  assign N5649 = N5648 | data_masked[7131];
  assign N5648 = N5647 | data_masked[7259];
  assign N5647 = N5646 | data_masked[7387];
  assign N5646 = N5645 | data_masked[7515];
  assign N5645 = N5644 | data_masked[7643];
  assign N5644 = N5643 | data_masked[7771];
  assign N5643 = N5642 | data_masked[7899];
  assign N5642 = data_masked[8155] | data_masked[8027];
  assign data_o[92] = N5765 | data_masked[92];
  assign N5765 = N5764 | data_masked[220];
  assign N5764 = N5763 | data_masked[348];
  assign N5763 = N5762 | data_masked[476];
  assign N5762 = N5761 | data_masked[604];
  assign N5761 = N5760 | data_masked[732];
  assign N5760 = N5759 | data_masked[860];
  assign N5759 = N5758 | data_masked[988];
  assign N5758 = N5757 | data_masked[1116];
  assign N5757 = N5756 | data_masked[1244];
  assign N5756 = N5755 | data_masked[1372];
  assign N5755 = N5754 | data_masked[1500];
  assign N5754 = N5753 | data_masked[1628];
  assign N5753 = N5752 | data_masked[1756];
  assign N5752 = N5751 | data_masked[1884];
  assign N5751 = N5750 | data_masked[2012];
  assign N5750 = N5749 | data_masked[2140];
  assign N5749 = N5748 | data_masked[2268];
  assign N5748 = N5747 | data_masked[2396];
  assign N5747 = N5746 | data_masked[2524];
  assign N5746 = N5745 | data_masked[2652];
  assign N5745 = N5744 | data_masked[2780];
  assign N5744 = N5743 | data_masked[2908];
  assign N5743 = N5742 | data_masked[3036];
  assign N5742 = N5741 | data_masked[3164];
  assign N5741 = N5740 | data_masked[3292];
  assign N5740 = N5739 | data_masked[3420];
  assign N5739 = N5738 | data_masked[3548];
  assign N5738 = N5737 | data_masked[3676];
  assign N5737 = N5736 | data_masked[3804];
  assign N5736 = N5735 | data_masked[3932];
  assign N5735 = N5734 | data_masked[4060];
  assign N5734 = N5733 | data_masked[4188];
  assign N5733 = N5732 | data_masked[4316];
  assign N5732 = N5731 | data_masked[4444];
  assign N5731 = N5730 | data_masked[4572];
  assign N5730 = N5729 | data_masked[4700];
  assign N5729 = N5728 | data_masked[4828];
  assign N5728 = N5727 | data_masked[4956];
  assign N5727 = N5726 | data_masked[5084];
  assign N5726 = N5725 | data_masked[5212];
  assign N5725 = N5724 | data_masked[5340];
  assign N5724 = N5723 | data_masked[5468];
  assign N5723 = N5722 | data_masked[5596];
  assign N5722 = N5721 | data_masked[5724];
  assign N5721 = N5720 | data_masked[5852];
  assign N5720 = N5719 | data_masked[5980];
  assign N5719 = N5718 | data_masked[6108];
  assign N5718 = N5717 | data_masked[6236];
  assign N5717 = N5716 | data_masked[6364];
  assign N5716 = N5715 | data_masked[6492];
  assign N5715 = N5714 | data_masked[6620];
  assign N5714 = N5713 | data_masked[6748];
  assign N5713 = N5712 | data_masked[6876];
  assign N5712 = N5711 | data_masked[7004];
  assign N5711 = N5710 | data_masked[7132];
  assign N5710 = N5709 | data_masked[7260];
  assign N5709 = N5708 | data_masked[7388];
  assign N5708 = N5707 | data_masked[7516];
  assign N5707 = N5706 | data_masked[7644];
  assign N5706 = N5705 | data_masked[7772];
  assign N5705 = N5704 | data_masked[7900];
  assign N5704 = data_masked[8156] | data_masked[8028];
  assign data_o[93] = N5827 | data_masked[93];
  assign N5827 = N5826 | data_masked[221];
  assign N5826 = N5825 | data_masked[349];
  assign N5825 = N5824 | data_masked[477];
  assign N5824 = N5823 | data_masked[605];
  assign N5823 = N5822 | data_masked[733];
  assign N5822 = N5821 | data_masked[861];
  assign N5821 = N5820 | data_masked[989];
  assign N5820 = N5819 | data_masked[1117];
  assign N5819 = N5818 | data_masked[1245];
  assign N5818 = N5817 | data_masked[1373];
  assign N5817 = N5816 | data_masked[1501];
  assign N5816 = N5815 | data_masked[1629];
  assign N5815 = N5814 | data_masked[1757];
  assign N5814 = N5813 | data_masked[1885];
  assign N5813 = N5812 | data_masked[2013];
  assign N5812 = N5811 | data_masked[2141];
  assign N5811 = N5810 | data_masked[2269];
  assign N5810 = N5809 | data_masked[2397];
  assign N5809 = N5808 | data_masked[2525];
  assign N5808 = N5807 | data_masked[2653];
  assign N5807 = N5806 | data_masked[2781];
  assign N5806 = N5805 | data_masked[2909];
  assign N5805 = N5804 | data_masked[3037];
  assign N5804 = N5803 | data_masked[3165];
  assign N5803 = N5802 | data_masked[3293];
  assign N5802 = N5801 | data_masked[3421];
  assign N5801 = N5800 | data_masked[3549];
  assign N5800 = N5799 | data_masked[3677];
  assign N5799 = N5798 | data_masked[3805];
  assign N5798 = N5797 | data_masked[3933];
  assign N5797 = N5796 | data_masked[4061];
  assign N5796 = N5795 | data_masked[4189];
  assign N5795 = N5794 | data_masked[4317];
  assign N5794 = N5793 | data_masked[4445];
  assign N5793 = N5792 | data_masked[4573];
  assign N5792 = N5791 | data_masked[4701];
  assign N5791 = N5790 | data_masked[4829];
  assign N5790 = N5789 | data_masked[4957];
  assign N5789 = N5788 | data_masked[5085];
  assign N5788 = N5787 | data_masked[5213];
  assign N5787 = N5786 | data_masked[5341];
  assign N5786 = N5785 | data_masked[5469];
  assign N5785 = N5784 | data_masked[5597];
  assign N5784 = N5783 | data_masked[5725];
  assign N5783 = N5782 | data_masked[5853];
  assign N5782 = N5781 | data_masked[5981];
  assign N5781 = N5780 | data_masked[6109];
  assign N5780 = N5779 | data_masked[6237];
  assign N5779 = N5778 | data_masked[6365];
  assign N5778 = N5777 | data_masked[6493];
  assign N5777 = N5776 | data_masked[6621];
  assign N5776 = N5775 | data_masked[6749];
  assign N5775 = N5774 | data_masked[6877];
  assign N5774 = N5773 | data_masked[7005];
  assign N5773 = N5772 | data_masked[7133];
  assign N5772 = N5771 | data_masked[7261];
  assign N5771 = N5770 | data_masked[7389];
  assign N5770 = N5769 | data_masked[7517];
  assign N5769 = N5768 | data_masked[7645];
  assign N5768 = N5767 | data_masked[7773];
  assign N5767 = N5766 | data_masked[7901];
  assign N5766 = data_masked[8157] | data_masked[8029];
  assign data_o[94] = N5889 | data_masked[94];
  assign N5889 = N5888 | data_masked[222];
  assign N5888 = N5887 | data_masked[350];
  assign N5887 = N5886 | data_masked[478];
  assign N5886 = N5885 | data_masked[606];
  assign N5885 = N5884 | data_masked[734];
  assign N5884 = N5883 | data_masked[862];
  assign N5883 = N5882 | data_masked[990];
  assign N5882 = N5881 | data_masked[1118];
  assign N5881 = N5880 | data_masked[1246];
  assign N5880 = N5879 | data_masked[1374];
  assign N5879 = N5878 | data_masked[1502];
  assign N5878 = N5877 | data_masked[1630];
  assign N5877 = N5876 | data_masked[1758];
  assign N5876 = N5875 | data_masked[1886];
  assign N5875 = N5874 | data_masked[2014];
  assign N5874 = N5873 | data_masked[2142];
  assign N5873 = N5872 | data_masked[2270];
  assign N5872 = N5871 | data_masked[2398];
  assign N5871 = N5870 | data_masked[2526];
  assign N5870 = N5869 | data_masked[2654];
  assign N5869 = N5868 | data_masked[2782];
  assign N5868 = N5867 | data_masked[2910];
  assign N5867 = N5866 | data_masked[3038];
  assign N5866 = N5865 | data_masked[3166];
  assign N5865 = N5864 | data_masked[3294];
  assign N5864 = N5863 | data_masked[3422];
  assign N5863 = N5862 | data_masked[3550];
  assign N5862 = N5861 | data_masked[3678];
  assign N5861 = N5860 | data_masked[3806];
  assign N5860 = N5859 | data_masked[3934];
  assign N5859 = N5858 | data_masked[4062];
  assign N5858 = N5857 | data_masked[4190];
  assign N5857 = N5856 | data_masked[4318];
  assign N5856 = N5855 | data_masked[4446];
  assign N5855 = N5854 | data_masked[4574];
  assign N5854 = N5853 | data_masked[4702];
  assign N5853 = N5852 | data_masked[4830];
  assign N5852 = N5851 | data_masked[4958];
  assign N5851 = N5850 | data_masked[5086];
  assign N5850 = N5849 | data_masked[5214];
  assign N5849 = N5848 | data_masked[5342];
  assign N5848 = N5847 | data_masked[5470];
  assign N5847 = N5846 | data_masked[5598];
  assign N5846 = N5845 | data_masked[5726];
  assign N5845 = N5844 | data_masked[5854];
  assign N5844 = N5843 | data_masked[5982];
  assign N5843 = N5842 | data_masked[6110];
  assign N5842 = N5841 | data_masked[6238];
  assign N5841 = N5840 | data_masked[6366];
  assign N5840 = N5839 | data_masked[6494];
  assign N5839 = N5838 | data_masked[6622];
  assign N5838 = N5837 | data_masked[6750];
  assign N5837 = N5836 | data_masked[6878];
  assign N5836 = N5835 | data_masked[7006];
  assign N5835 = N5834 | data_masked[7134];
  assign N5834 = N5833 | data_masked[7262];
  assign N5833 = N5832 | data_masked[7390];
  assign N5832 = N5831 | data_masked[7518];
  assign N5831 = N5830 | data_masked[7646];
  assign N5830 = N5829 | data_masked[7774];
  assign N5829 = N5828 | data_masked[7902];
  assign N5828 = data_masked[8158] | data_masked[8030];
  assign data_o[95] = N5951 | data_masked[95];
  assign N5951 = N5950 | data_masked[223];
  assign N5950 = N5949 | data_masked[351];
  assign N5949 = N5948 | data_masked[479];
  assign N5948 = N5947 | data_masked[607];
  assign N5947 = N5946 | data_masked[735];
  assign N5946 = N5945 | data_masked[863];
  assign N5945 = N5944 | data_masked[991];
  assign N5944 = N5943 | data_masked[1119];
  assign N5943 = N5942 | data_masked[1247];
  assign N5942 = N5941 | data_masked[1375];
  assign N5941 = N5940 | data_masked[1503];
  assign N5940 = N5939 | data_masked[1631];
  assign N5939 = N5938 | data_masked[1759];
  assign N5938 = N5937 | data_masked[1887];
  assign N5937 = N5936 | data_masked[2015];
  assign N5936 = N5935 | data_masked[2143];
  assign N5935 = N5934 | data_masked[2271];
  assign N5934 = N5933 | data_masked[2399];
  assign N5933 = N5932 | data_masked[2527];
  assign N5932 = N5931 | data_masked[2655];
  assign N5931 = N5930 | data_masked[2783];
  assign N5930 = N5929 | data_masked[2911];
  assign N5929 = N5928 | data_masked[3039];
  assign N5928 = N5927 | data_masked[3167];
  assign N5927 = N5926 | data_masked[3295];
  assign N5926 = N5925 | data_masked[3423];
  assign N5925 = N5924 | data_masked[3551];
  assign N5924 = N5923 | data_masked[3679];
  assign N5923 = N5922 | data_masked[3807];
  assign N5922 = N5921 | data_masked[3935];
  assign N5921 = N5920 | data_masked[4063];
  assign N5920 = N5919 | data_masked[4191];
  assign N5919 = N5918 | data_masked[4319];
  assign N5918 = N5917 | data_masked[4447];
  assign N5917 = N5916 | data_masked[4575];
  assign N5916 = N5915 | data_masked[4703];
  assign N5915 = N5914 | data_masked[4831];
  assign N5914 = N5913 | data_masked[4959];
  assign N5913 = N5912 | data_masked[5087];
  assign N5912 = N5911 | data_masked[5215];
  assign N5911 = N5910 | data_masked[5343];
  assign N5910 = N5909 | data_masked[5471];
  assign N5909 = N5908 | data_masked[5599];
  assign N5908 = N5907 | data_masked[5727];
  assign N5907 = N5906 | data_masked[5855];
  assign N5906 = N5905 | data_masked[5983];
  assign N5905 = N5904 | data_masked[6111];
  assign N5904 = N5903 | data_masked[6239];
  assign N5903 = N5902 | data_masked[6367];
  assign N5902 = N5901 | data_masked[6495];
  assign N5901 = N5900 | data_masked[6623];
  assign N5900 = N5899 | data_masked[6751];
  assign N5899 = N5898 | data_masked[6879];
  assign N5898 = N5897 | data_masked[7007];
  assign N5897 = N5896 | data_masked[7135];
  assign N5896 = N5895 | data_masked[7263];
  assign N5895 = N5894 | data_masked[7391];
  assign N5894 = N5893 | data_masked[7519];
  assign N5893 = N5892 | data_masked[7647];
  assign N5892 = N5891 | data_masked[7775];
  assign N5891 = N5890 | data_masked[7903];
  assign N5890 = data_masked[8159] | data_masked[8031];
  assign data_o[96] = N6013 | data_masked[96];
  assign N6013 = N6012 | data_masked[224];
  assign N6012 = N6011 | data_masked[352];
  assign N6011 = N6010 | data_masked[480];
  assign N6010 = N6009 | data_masked[608];
  assign N6009 = N6008 | data_masked[736];
  assign N6008 = N6007 | data_masked[864];
  assign N6007 = N6006 | data_masked[992];
  assign N6006 = N6005 | data_masked[1120];
  assign N6005 = N6004 | data_masked[1248];
  assign N6004 = N6003 | data_masked[1376];
  assign N6003 = N6002 | data_masked[1504];
  assign N6002 = N6001 | data_masked[1632];
  assign N6001 = N6000 | data_masked[1760];
  assign N6000 = N5999 | data_masked[1888];
  assign N5999 = N5998 | data_masked[2016];
  assign N5998 = N5997 | data_masked[2144];
  assign N5997 = N5996 | data_masked[2272];
  assign N5996 = N5995 | data_masked[2400];
  assign N5995 = N5994 | data_masked[2528];
  assign N5994 = N5993 | data_masked[2656];
  assign N5993 = N5992 | data_masked[2784];
  assign N5992 = N5991 | data_masked[2912];
  assign N5991 = N5990 | data_masked[3040];
  assign N5990 = N5989 | data_masked[3168];
  assign N5989 = N5988 | data_masked[3296];
  assign N5988 = N5987 | data_masked[3424];
  assign N5987 = N5986 | data_masked[3552];
  assign N5986 = N5985 | data_masked[3680];
  assign N5985 = N5984 | data_masked[3808];
  assign N5984 = N5983 | data_masked[3936];
  assign N5983 = N5982 | data_masked[4064];
  assign N5982 = N5981 | data_masked[4192];
  assign N5981 = N5980 | data_masked[4320];
  assign N5980 = N5979 | data_masked[4448];
  assign N5979 = N5978 | data_masked[4576];
  assign N5978 = N5977 | data_masked[4704];
  assign N5977 = N5976 | data_masked[4832];
  assign N5976 = N5975 | data_masked[4960];
  assign N5975 = N5974 | data_masked[5088];
  assign N5974 = N5973 | data_masked[5216];
  assign N5973 = N5972 | data_masked[5344];
  assign N5972 = N5971 | data_masked[5472];
  assign N5971 = N5970 | data_masked[5600];
  assign N5970 = N5969 | data_masked[5728];
  assign N5969 = N5968 | data_masked[5856];
  assign N5968 = N5967 | data_masked[5984];
  assign N5967 = N5966 | data_masked[6112];
  assign N5966 = N5965 | data_masked[6240];
  assign N5965 = N5964 | data_masked[6368];
  assign N5964 = N5963 | data_masked[6496];
  assign N5963 = N5962 | data_masked[6624];
  assign N5962 = N5961 | data_masked[6752];
  assign N5961 = N5960 | data_masked[6880];
  assign N5960 = N5959 | data_masked[7008];
  assign N5959 = N5958 | data_masked[7136];
  assign N5958 = N5957 | data_masked[7264];
  assign N5957 = N5956 | data_masked[7392];
  assign N5956 = N5955 | data_masked[7520];
  assign N5955 = N5954 | data_masked[7648];
  assign N5954 = N5953 | data_masked[7776];
  assign N5953 = N5952 | data_masked[7904];
  assign N5952 = data_masked[8160] | data_masked[8032];
  assign data_o[97] = N6075 | data_masked[97];
  assign N6075 = N6074 | data_masked[225];
  assign N6074 = N6073 | data_masked[353];
  assign N6073 = N6072 | data_masked[481];
  assign N6072 = N6071 | data_masked[609];
  assign N6071 = N6070 | data_masked[737];
  assign N6070 = N6069 | data_masked[865];
  assign N6069 = N6068 | data_masked[993];
  assign N6068 = N6067 | data_masked[1121];
  assign N6067 = N6066 | data_masked[1249];
  assign N6066 = N6065 | data_masked[1377];
  assign N6065 = N6064 | data_masked[1505];
  assign N6064 = N6063 | data_masked[1633];
  assign N6063 = N6062 | data_masked[1761];
  assign N6062 = N6061 | data_masked[1889];
  assign N6061 = N6060 | data_masked[2017];
  assign N6060 = N6059 | data_masked[2145];
  assign N6059 = N6058 | data_masked[2273];
  assign N6058 = N6057 | data_masked[2401];
  assign N6057 = N6056 | data_masked[2529];
  assign N6056 = N6055 | data_masked[2657];
  assign N6055 = N6054 | data_masked[2785];
  assign N6054 = N6053 | data_masked[2913];
  assign N6053 = N6052 | data_masked[3041];
  assign N6052 = N6051 | data_masked[3169];
  assign N6051 = N6050 | data_masked[3297];
  assign N6050 = N6049 | data_masked[3425];
  assign N6049 = N6048 | data_masked[3553];
  assign N6048 = N6047 | data_masked[3681];
  assign N6047 = N6046 | data_masked[3809];
  assign N6046 = N6045 | data_masked[3937];
  assign N6045 = N6044 | data_masked[4065];
  assign N6044 = N6043 | data_masked[4193];
  assign N6043 = N6042 | data_masked[4321];
  assign N6042 = N6041 | data_masked[4449];
  assign N6041 = N6040 | data_masked[4577];
  assign N6040 = N6039 | data_masked[4705];
  assign N6039 = N6038 | data_masked[4833];
  assign N6038 = N6037 | data_masked[4961];
  assign N6037 = N6036 | data_masked[5089];
  assign N6036 = N6035 | data_masked[5217];
  assign N6035 = N6034 | data_masked[5345];
  assign N6034 = N6033 | data_masked[5473];
  assign N6033 = N6032 | data_masked[5601];
  assign N6032 = N6031 | data_masked[5729];
  assign N6031 = N6030 | data_masked[5857];
  assign N6030 = N6029 | data_masked[5985];
  assign N6029 = N6028 | data_masked[6113];
  assign N6028 = N6027 | data_masked[6241];
  assign N6027 = N6026 | data_masked[6369];
  assign N6026 = N6025 | data_masked[6497];
  assign N6025 = N6024 | data_masked[6625];
  assign N6024 = N6023 | data_masked[6753];
  assign N6023 = N6022 | data_masked[6881];
  assign N6022 = N6021 | data_masked[7009];
  assign N6021 = N6020 | data_masked[7137];
  assign N6020 = N6019 | data_masked[7265];
  assign N6019 = N6018 | data_masked[7393];
  assign N6018 = N6017 | data_masked[7521];
  assign N6017 = N6016 | data_masked[7649];
  assign N6016 = N6015 | data_masked[7777];
  assign N6015 = N6014 | data_masked[7905];
  assign N6014 = data_masked[8161] | data_masked[8033];
  assign data_o[98] = N6137 | data_masked[98];
  assign N6137 = N6136 | data_masked[226];
  assign N6136 = N6135 | data_masked[354];
  assign N6135 = N6134 | data_masked[482];
  assign N6134 = N6133 | data_masked[610];
  assign N6133 = N6132 | data_masked[738];
  assign N6132 = N6131 | data_masked[866];
  assign N6131 = N6130 | data_masked[994];
  assign N6130 = N6129 | data_masked[1122];
  assign N6129 = N6128 | data_masked[1250];
  assign N6128 = N6127 | data_masked[1378];
  assign N6127 = N6126 | data_masked[1506];
  assign N6126 = N6125 | data_masked[1634];
  assign N6125 = N6124 | data_masked[1762];
  assign N6124 = N6123 | data_masked[1890];
  assign N6123 = N6122 | data_masked[2018];
  assign N6122 = N6121 | data_masked[2146];
  assign N6121 = N6120 | data_masked[2274];
  assign N6120 = N6119 | data_masked[2402];
  assign N6119 = N6118 | data_masked[2530];
  assign N6118 = N6117 | data_masked[2658];
  assign N6117 = N6116 | data_masked[2786];
  assign N6116 = N6115 | data_masked[2914];
  assign N6115 = N6114 | data_masked[3042];
  assign N6114 = N6113 | data_masked[3170];
  assign N6113 = N6112 | data_masked[3298];
  assign N6112 = N6111 | data_masked[3426];
  assign N6111 = N6110 | data_masked[3554];
  assign N6110 = N6109 | data_masked[3682];
  assign N6109 = N6108 | data_masked[3810];
  assign N6108 = N6107 | data_masked[3938];
  assign N6107 = N6106 | data_masked[4066];
  assign N6106 = N6105 | data_masked[4194];
  assign N6105 = N6104 | data_masked[4322];
  assign N6104 = N6103 | data_masked[4450];
  assign N6103 = N6102 | data_masked[4578];
  assign N6102 = N6101 | data_masked[4706];
  assign N6101 = N6100 | data_masked[4834];
  assign N6100 = N6099 | data_masked[4962];
  assign N6099 = N6098 | data_masked[5090];
  assign N6098 = N6097 | data_masked[5218];
  assign N6097 = N6096 | data_masked[5346];
  assign N6096 = N6095 | data_masked[5474];
  assign N6095 = N6094 | data_masked[5602];
  assign N6094 = N6093 | data_masked[5730];
  assign N6093 = N6092 | data_masked[5858];
  assign N6092 = N6091 | data_masked[5986];
  assign N6091 = N6090 | data_masked[6114];
  assign N6090 = N6089 | data_masked[6242];
  assign N6089 = N6088 | data_masked[6370];
  assign N6088 = N6087 | data_masked[6498];
  assign N6087 = N6086 | data_masked[6626];
  assign N6086 = N6085 | data_masked[6754];
  assign N6085 = N6084 | data_masked[6882];
  assign N6084 = N6083 | data_masked[7010];
  assign N6083 = N6082 | data_masked[7138];
  assign N6082 = N6081 | data_masked[7266];
  assign N6081 = N6080 | data_masked[7394];
  assign N6080 = N6079 | data_masked[7522];
  assign N6079 = N6078 | data_masked[7650];
  assign N6078 = N6077 | data_masked[7778];
  assign N6077 = N6076 | data_masked[7906];
  assign N6076 = data_masked[8162] | data_masked[8034];
  assign data_o[99] = N6199 | data_masked[99];
  assign N6199 = N6198 | data_masked[227];
  assign N6198 = N6197 | data_masked[355];
  assign N6197 = N6196 | data_masked[483];
  assign N6196 = N6195 | data_masked[611];
  assign N6195 = N6194 | data_masked[739];
  assign N6194 = N6193 | data_masked[867];
  assign N6193 = N6192 | data_masked[995];
  assign N6192 = N6191 | data_masked[1123];
  assign N6191 = N6190 | data_masked[1251];
  assign N6190 = N6189 | data_masked[1379];
  assign N6189 = N6188 | data_masked[1507];
  assign N6188 = N6187 | data_masked[1635];
  assign N6187 = N6186 | data_masked[1763];
  assign N6186 = N6185 | data_masked[1891];
  assign N6185 = N6184 | data_masked[2019];
  assign N6184 = N6183 | data_masked[2147];
  assign N6183 = N6182 | data_masked[2275];
  assign N6182 = N6181 | data_masked[2403];
  assign N6181 = N6180 | data_masked[2531];
  assign N6180 = N6179 | data_masked[2659];
  assign N6179 = N6178 | data_masked[2787];
  assign N6178 = N6177 | data_masked[2915];
  assign N6177 = N6176 | data_masked[3043];
  assign N6176 = N6175 | data_masked[3171];
  assign N6175 = N6174 | data_masked[3299];
  assign N6174 = N6173 | data_masked[3427];
  assign N6173 = N6172 | data_masked[3555];
  assign N6172 = N6171 | data_masked[3683];
  assign N6171 = N6170 | data_masked[3811];
  assign N6170 = N6169 | data_masked[3939];
  assign N6169 = N6168 | data_masked[4067];
  assign N6168 = N6167 | data_masked[4195];
  assign N6167 = N6166 | data_masked[4323];
  assign N6166 = N6165 | data_masked[4451];
  assign N6165 = N6164 | data_masked[4579];
  assign N6164 = N6163 | data_masked[4707];
  assign N6163 = N6162 | data_masked[4835];
  assign N6162 = N6161 | data_masked[4963];
  assign N6161 = N6160 | data_masked[5091];
  assign N6160 = N6159 | data_masked[5219];
  assign N6159 = N6158 | data_masked[5347];
  assign N6158 = N6157 | data_masked[5475];
  assign N6157 = N6156 | data_masked[5603];
  assign N6156 = N6155 | data_masked[5731];
  assign N6155 = N6154 | data_masked[5859];
  assign N6154 = N6153 | data_masked[5987];
  assign N6153 = N6152 | data_masked[6115];
  assign N6152 = N6151 | data_masked[6243];
  assign N6151 = N6150 | data_masked[6371];
  assign N6150 = N6149 | data_masked[6499];
  assign N6149 = N6148 | data_masked[6627];
  assign N6148 = N6147 | data_masked[6755];
  assign N6147 = N6146 | data_masked[6883];
  assign N6146 = N6145 | data_masked[7011];
  assign N6145 = N6144 | data_masked[7139];
  assign N6144 = N6143 | data_masked[7267];
  assign N6143 = N6142 | data_masked[7395];
  assign N6142 = N6141 | data_masked[7523];
  assign N6141 = N6140 | data_masked[7651];
  assign N6140 = N6139 | data_masked[7779];
  assign N6139 = N6138 | data_masked[7907];
  assign N6138 = data_masked[8163] | data_masked[8035];
  assign data_o[100] = N6261 | data_masked[100];
  assign N6261 = N6260 | data_masked[228];
  assign N6260 = N6259 | data_masked[356];
  assign N6259 = N6258 | data_masked[484];
  assign N6258 = N6257 | data_masked[612];
  assign N6257 = N6256 | data_masked[740];
  assign N6256 = N6255 | data_masked[868];
  assign N6255 = N6254 | data_masked[996];
  assign N6254 = N6253 | data_masked[1124];
  assign N6253 = N6252 | data_masked[1252];
  assign N6252 = N6251 | data_masked[1380];
  assign N6251 = N6250 | data_masked[1508];
  assign N6250 = N6249 | data_masked[1636];
  assign N6249 = N6248 | data_masked[1764];
  assign N6248 = N6247 | data_masked[1892];
  assign N6247 = N6246 | data_masked[2020];
  assign N6246 = N6245 | data_masked[2148];
  assign N6245 = N6244 | data_masked[2276];
  assign N6244 = N6243 | data_masked[2404];
  assign N6243 = N6242 | data_masked[2532];
  assign N6242 = N6241 | data_masked[2660];
  assign N6241 = N6240 | data_masked[2788];
  assign N6240 = N6239 | data_masked[2916];
  assign N6239 = N6238 | data_masked[3044];
  assign N6238 = N6237 | data_masked[3172];
  assign N6237 = N6236 | data_masked[3300];
  assign N6236 = N6235 | data_masked[3428];
  assign N6235 = N6234 | data_masked[3556];
  assign N6234 = N6233 | data_masked[3684];
  assign N6233 = N6232 | data_masked[3812];
  assign N6232 = N6231 | data_masked[3940];
  assign N6231 = N6230 | data_masked[4068];
  assign N6230 = N6229 | data_masked[4196];
  assign N6229 = N6228 | data_masked[4324];
  assign N6228 = N6227 | data_masked[4452];
  assign N6227 = N6226 | data_masked[4580];
  assign N6226 = N6225 | data_masked[4708];
  assign N6225 = N6224 | data_masked[4836];
  assign N6224 = N6223 | data_masked[4964];
  assign N6223 = N6222 | data_masked[5092];
  assign N6222 = N6221 | data_masked[5220];
  assign N6221 = N6220 | data_masked[5348];
  assign N6220 = N6219 | data_masked[5476];
  assign N6219 = N6218 | data_masked[5604];
  assign N6218 = N6217 | data_masked[5732];
  assign N6217 = N6216 | data_masked[5860];
  assign N6216 = N6215 | data_masked[5988];
  assign N6215 = N6214 | data_masked[6116];
  assign N6214 = N6213 | data_masked[6244];
  assign N6213 = N6212 | data_masked[6372];
  assign N6212 = N6211 | data_masked[6500];
  assign N6211 = N6210 | data_masked[6628];
  assign N6210 = N6209 | data_masked[6756];
  assign N6209 = N6208 | data_masked[6884];
  assign N6208 = N6207 | data_masked[7012];
  assign N6207 = N6206 | data_masked[7140];
  assign N6206 = N6205 | data_masked[7268];
  assign N6205 = N6204 | data_masked[7396];
  assign N6204 = N6203 | data_masked[7524];
  assign N6203 = N6202 | data_masked[7652];
  assign N6202 = N6201 | data_masked[7780];
  assign N6201 = N6200 | data_masked[7908];
  assign N6200 = data_masked[8164] | data_masked[8036];
  assign data_o[101] = N6323 | data_masked[101];
  assign N6323 = N6322 | data_masked[229];
  assign N6322 = N6321 | data_masked[357];
  assign N6321 = N6320 | data_masked[485];
  assign N6320 = N6319 | data_masked[613];
  assign N6319 = N6318 | data_masked[741];
  assign N6318 = N6317 | data_masked[869];
  assign N6317 = N6316 | data_masked[997];
  assign N6316 = N6315 | data_masked[1125];
  assign N6315 = N6314 | data_masked[1253];
  assign N6314 = N6313 | data_masked[1381];
  assign N6313 = N6312 | data_masked[1509];
  assign N6312 = N6311 | data_masked[1637];
  assign N6311 = N6310 | data_masked[1765];
  assign N6310 = N6309 | data_masked[1893];
  assign N6309 = N6308 | data_masked[2021];
  assign N6308 = N6307 | data_masked[2149];
  assign N6307 = N6306 | data_masked[2277];
  assign N6306 = N6305 | data_masked[2405];
  assign N6305 = N6304 | data_masked[2533];
  assign N6304 = N6303 | data_masked[2661];
  assign N6303 = N6302 | data_masked[2789];
  assign N6302 = N6301 | data_masked[2917];
  assign N6301 = N6300 | data_masked[3045];
  assign N6300 = N6299 | data_masked[3173];
  assign N6299 = N6298 | data_masked[3301];
  assign N6298 = N6297 | data_masked[3429];
  assign N6297 = N6296 | data_masked[3557];
  assign N6296 = N6295 | data_masked[3685];
  assign N6295 = N6294 | data_masked[3813];
  assign N6294 = N6293 | data_masked[3941];
  assign N6293 = N6292 | data_masked[4069];
  assign N6292 = N6291 | data_masked[4197];
  assign N6291 = N6290 | data_masked[4325];
  assign N6290 = N6289 | data_masked[4453];
  assign N6289 = N6288 | data_masked[4581];
  assign N6288 = N6287 | data_masked[4709];
  assign N6287 = N6286 | data_masked[4837];
  assign N6286 = N6285 | data_masked[4965];
  assign N6285 = N6284 | data_masked[5093];
  assign N6284 = N6283 | data_masked[5221];
  assign N6283 = N6282 | data_masked[5349];
  assign N6282 = N6281 | data_masked[5477];
  assign N6281 = N6280 | data_masked[5605];
  assign N6280 = N6279 | data_masked[5733];
  assign N6279 = N6278 | data_masked[5861];
  assign N6278 = N6277 | data_masked[5989];
  assign N6277 = N6276 | data_masked[6117];
  assign N6276 = N6275 | data_masked[6245];
  assign N6275 = N6274 | data_masked[6373];
  assign N6274 = N6273 | data_masked[6501];
  assign N6273 = N6272 | data_masked[6629];
  assign N6272 = N6271 | data_masked[6757];
  assign N6271 = N6270 | data_masked[6885];
  assign N6270 = N6269 | data_masked[7013];
  assign N6269 = N6268 | data_masked[7141];
  assign N6268 = N6267 | data_masked[7269];
  assign N6267 = N6266 | data_masked[7397];
  assign N6266 = N6265 | data_masked[7525];
  assign N6265 = N6264 | data_masked[7653];
  assign N6264 = N6263 | data_masked[7781];
  assign N6263 = N6262 | data_masked[7909];
  assign N6262 = data_masked[8165] | data_masked[8037];
  assign data_o[102] = N6385 | data_masked[102];
  assign N6385 = N6384 | data_masked[230];
  assign N6384 = N6383 | data_masked[358];
  assign N6383 = N6382 | data_masked[486];
  assign N6382 = N6381 | data_masked[614];
  assign N6381 = N6380 | data_masked[742];
  assign N6380 = N6379 | data_masked[870];
  assign N6379 = N6378 | data_masked[998];
  assign N6378 = N6377 | data_masked[1126];
  assign N6377 = N6376 | data_masked[1254];
  assign N6376 = N6375 | data_masked[1382];
  assign N6375 = N6374 | data_masked[1510];
  assign N6374 = N6373 | data_masked[1638];
  assign N6373 = N6372 | data_masked[1766];
  assign N6372 = N6371 | data_masked[1894];
  assign N6371 = N6370 | data_masked[2022];
  assign N6370 = N6369 | data_masked[2150];
  assign N6369 = N6368 | data_masked[2278];
  assign N6368 = N6367 | data_masked[2406];
  assign N6367 = N6366 | data_masked[2534];
  assign N6366 = N6365 | data_masked[2662];
  assign N6365 = N6364 | data_masked[2790];
  assign N6364 = N6363 | data_masked[2918];
  assign N6363 = N6362 | data_masked[3046];
  assign N6362 = N6361 | data_masked[3174];
  assign N6361 = N6360 | data_masked[3302];
  assign N6360 = N6359 | data_masked[3430];
  assign N6359 = N6358 | data_masked[3558];
  assign N6358 = N6357 | data_masked[3686];
  assign N6357 = N6356 | data_masked[3814];
  assign N6356 = N6355 | data_masked[3942];
  assign N6355 = N6354 | data_masked[4070];
  assign N6354 = N6353 | data_masked[4198];
  assign N6353 = N6352 | data_masked[4326];
  assign N6352 = N6351 | data_masked[4454];
  assign N6351 = N6350 | data_masked[4582];
  assign N6350 = N6349 | data_masked[4710];
  assign N6349 = N6348 | data_masked[4838];
  assign N6348 = N6347 | data_masked[4966];
  assign N6347 = N6346 | data_masked[5094];
  assign N6346 = N6345 | data_masked[5222];
  assign N6345 = N6344 | data_masked[5350];
  assign N6344 = N6343 | data_masked[5478];
  assign N6343 = N6342 | data_masked[5606];
  assign N6342 = N6341 | data_masked[5734];
  assign N6341 = N6340 | data_masked[5862];
  assign N6340 = N6339 | data_masked[5990];
  assign N6339 = N6338 | data_masked[6118];
  assign N6338 = N6337 | data_masked[6246];
  assign N6337 = N6336 | data_masked[6374];
  assign N6336 = N6335 | data_masked[6502];
  assign N6335 = N6334 | data_masked[6630];
  assign N6334 = N6333 | data_masked[6758];
  assign N6333 = N6332 | data_masked[6886];
  assign N6332 = N6331 | data_masked[7014];
  assign N6331 = N6330 | data_masked[7142];
  assign N6330 = N6329 | data_masked[7270];
  assign N6329 = N6328 | data_masked[7398];
  assign N6328 = N6327 | data_masked[7526];
  assign N6327 = N6326 | data_masked[7654];
  assign N6326 = N6325 | data_masked[7782];
  assign N6325 = N6324 | data_masked[7910];
  assign N6324 = data_masked[8166] | data_masked[8038];
  assign data_o[103] = N6447 | data_masked[103];
  assign N6447 = N6446 | data_masked[231];
  assign N6446 = N6445 | data_masked[359];
  assign N6445 = N6444 | data_masked[487];
  assign N6444 = N6443 | data_masked[615];
  assign N6443 = N6442 | data_masked[743];
  assign N6442 = N6441 | data_masked[871];
  assign N6441 = N6440 | data_masked[999];
  assign N6440 = N6439 | data_masked[1127];
  assign N6439 = N6438 | data_masked[1255];
  assign N6438 = N6437 | data_masked[1383];
  assign N6437 = N6436 | data_masked[1511];
  assign N6436 = N6435 | data_masked[1639];
  assign N6435 = N6434 | data_masked[1767];
  assign N6434 = N6433 | data_masked[1895];
  assign N6433 = N6432 | data_masked[2023];
  assign N6432 = N6431 | data_masked[2151];
  assign N6431 = N6430 | data_masked[2279];
  assign N6430 = N6429 | data_masked[2407];
  assign N6429 = N6428 | data_masked[2535];
  assign N6428 = N6427 | data_masked[2663];
  assign N6427 = N6426 | data_masked[2791];
  assign N6426 = N6425 | data_masked[2919];
  assign N6425 = N6424 | data_masked[3047];
  assign N6424 = N6423 | data_masked[3175];
  assign N6423 = N6422 | data_masked[3303];
  assign N6422 = N6421 | data_masked[3431];
  assign N6421 = N6420 | data_masked[3559];
  assign N6420 = N6419 | data_masked[3687];
  assign N6419 = N6418 | data_masked[3815];
  assign N6418 = N6417 | data_masked[3943];
  assign N6417 = N6416 | data_masked[4071];
  assign N6416 = N6415 | data_masked[4199];
  assign N6415 = N6414 | data_masked[4327];
  assign N6414 = N6413 | data_masked[4455];
  assign N6413 = N6412 | data_masked[4583];
  assign N6412 = N6411 | data_masked[4711];
  assign N6411 = N6410 | data_masked[4839];
  assign N6410 = N6409 | data_masked[4967];
  assign N6409 = N6408 | data_masked[5095];
  assign N6408 = N6407 | data_masked[5223];
  assign N6407 = N6406 | data_masked[5351];
  assign N6406 = N6405 | data_masked[5479];
  assign N6405 = N6404 | data_masked[5607];
  assign N6404 = N6403 | data_masked[5735];
  assign N6403 = N6402 | data_masked[5863];
  assign N6402 = N6401 | data_masked[5991];
  assign N6401 = N6400 | data_masked[6119];
  assign N6400 = N6399 | data_masked[6247];
  assign N6399 = N6398 | data_masked[6375];
  assign N6398 = N6397 | data_masked[6503];
  assign N6397 = N6396 | data_masked[6631];
  assign N6396 = N6395 | data_masked[6759];
  assign N6395 = N6394 | data_masked[6887];
  assign N6394 = N6393 | data_masked[7015];
  assign N6393 = N6392 | data_masked[7143];
  assign N6392 = N6391 | data_masked[7271];
  assign N6391 = N6390 | data_masked[7399];
  assign N6390 = N6389 | data_masked[7527];
  assign N6389 = N6388 | data_masked[7655];
  assign N6388 = N6387 | data_masked[7783];
  assign N6387 = N6386 | data_masked[7911];
  assign N6386 = data_masked[8167] | data_masked[8039];
  assign data_o[104] = N6509 | data_masked[104];
  assign N6509 = N6508 | data_masked[232];
  assign N6508 = N6507 | data_masked[360];
  assign N6507 = N6506 | data_masked[488];
  assign N6506 = N6505 | data_masked[616];
  assign N6505 = N6504 | data_masked[744];
  assign N6504 = N6503 | data_masked[872];
  assign N6503 = N6502 | data_masked[1000];
  assign N6502 = N6501 | data_masked[1128];
  assign N6501 = N6500 | data_masked[1256];
  assign N6500 = N6499 | data_masked[1384];
  assign N6499 = N6498 | data_masked[1512];
  assign N6498 = N6497 | data_masked[1640];
  assign N6497 = N6496 | data_masked[1768];
  assign N6496 = N6495 | data_masked[1896];
  assign N6495 = N6494 | data_masked[2024];
  assign N6494 = N6493 | data_masked[2152];
  assign N6493 = N6492 | data_masked[2280];
  assign N6492 = N6491 | data_masked[2408];
  assign N6491 = N6490 | data_masked[2536];
  assign N6490 = N6489 | data_masked[2664];
  assign N6489 = N6488 | data_masked[2792];
  assign N6488 = N6487 | data_masked[2920];
  assign N6487 = N6486 | data_masked[3048];
  assign N6486 = N6485 | data_masked[3176];
  assign N6485 = N6484 | data_masked[3304];
  assign N6484 = N6483 | data_masked[3432];
  assign N6483 = N6482 | data_masked[3560];
  assign N6482 = N6481 | data_masked[3688];
  assign N6481 = N6480 | data_masked[3816];
  assign N6480 = N6479 | data_masked[3944];
  assign N6479 = N6478 | data_masked[4072];
  assign N6478 = N6477 | data_masked[4200];
  assign N6477 = N6476 | data_masked[4328];
  assign N6476 = N6475 | data_masked[4456];
  assign N6475 = N6474 | data_masked[4584];
  assign N6474 = N6473 | data_masked[4712];
  assign N6473 = N6472 | data_masked[4840];
  assign N6472 = N6471 | data_masked[4968];
  assign N6471 = N6470 | data_masked[5096];
  assign N6470 = N6469 | data_masked[5224];
  assign N6469 = N6468 | data_masked[5352];
  assign N6468 = N6467 | data_masked[5480];
  assign N6467 = N6466 | data_masked[5608];
  assign N6466 = N6465 | data_masked[5736];
  assign N6465 = N6464 | data_masked[5864];
  assign N6464 = N6463 | data_masked[5992];
  assign N6463 = N6462 | data_masked[6120];
  assign N6462 = N6461 | data_masked[6248];
  assign N6461 = N6460 | data_masked[6376];
  assign N6460 = N6459 | data_masked[6504];
  assign N6459 = N6458 | data_masked[6632];
  assign N6458 = N6457 | data_masked[6760];
  assign N6457 = N6456 | data_masked[6888];
  assign N6456 = N6455 | data_masked[7016];
  assign N6455 = N6454 | data_masked[7144];
  assign N6454 = N6453 | data_masked[7272];
  assign N6453 = N6452 | data_masked[7400];
  assign N6452 = N6451 | data_masked[7528];
  assign N6451 = N6450 | data_masked[7656];
  assign N6450 = N6449 | data_masked[7784];
  assign N6449 = N6448 | data_masked[7912];
  assign N6448 = data_masked[8168] | data_masked[8040];
  assign data_o[105] = N6571 | data_masked[105];
  assign N6571 = N6570 | data_masked[233];
  assign N6570 = N6569 | data_masked[361];
  assign N6569 = N6568 | data_masked[489];
  assign N6568 = N6567 | data_masked[617];
  assign N6567 = N6566 | data_masked[745];
  assign N6566 = N6565 | data_masked[873];
  assign N6565 = N6564 | data_masked[1001];
  assign N6564 = N6563 | data_masked[1129];
  assign N6563 = N6562 | data_masked[1257];
  assign N6562 = N6561 | data_masked[1385];
  assign N6561 = N6560 | data_masked[1513];
  assign N6560 = N6559 | data_masked[1641];
  assign N6559 = N6558 | data_masked[1769];
  assign N6558 = N6557 | data_masked[1897];
  assign N6557 = N6556 | data_masked[2025];
  assign N6556 = N6555 | data_masked[2153];
  assign N6555 = N6554 | data_masked[2281];
  assign N6554 = N6553 | data_masked[2409];
  assign N6553 = N6552 | data_masked[2537];
  assign N6552 = N6551 | data_masked[2665];
  assign N6551 = N6550 | data_masked[2793];
  assign N6550 = N6549 | data_masked[2921];
  assign N6549 = N6548 | data_masked[3049];
  assign N6548 = N6547 | data_masked[3177];
  assign N6547 = N6546 | data_masked[3305];
  assign N6546 = N6545 | data_masked[3433];
  assign N6545 = N6544 | data_masked[3561];
  assign N6544 = N6543 | data_masked[3689];
  assign N6543 = N6542 | data_masked[3817];
  assign N6542 = N6541 | data_masked[3945];
  assign N6541 = N6540 | data_masked[4073];
  assign N6540 = N6539 | data_masked[4201];
  assign N6539 = N6538 | data_masked[4329];
  assign N6538 = N6537 | data_masked[4457];
  assign N6537 = N6536 | data_masked[4585];
  assign N6536 = N6535 | data_masked[4713];
  assign N6535 = N6534 | data_masked[4841];
  assign N6534 = N6533 | data_masked[4969];
  assign N6533 = N6532 | data_masked[5097];
  assign N6532 = N6531 | data_masked[5225];
  assign N6531 = N6530 | data_masked[5353];
  assign N6530 = N6529 | data_masked[5481];
  assign N6529 = N6528 | data_masked[5609];
  assign N6528 = N6527 | data_masked[5737];
  assign N6527 = N6526 | data_masked[5865];
  assign N6526 = N6525 | data_masked[5993];
  assign N6525 = N6524 | data_masked[6121];
  assign N6524 = N6523 | data_masked[6249];
  assign N6523 = N6522 | data_masked[6377];
  assign N6522 = N6521 | data_masked[6505];
  assign N6521 = N6520 | data_masked[6633];
  assign N6520 = N6519 | data_masked[6761];
  assign N6519 = N6518 | data_masked[6889];
  assign N6518 = N6517 | data_masked[7017];
  assign N6517 = N6516 | data_masked[7145];
  assign N6516 = N6515 | data_masked[7273];
  assign N6515 = N6514 | data_masked[7401];
  assign N6514 = N6513 | data_masked[7529];
  assign N6513 = N6512 | data_masked[7657];
  assign N6512 = N6511 | data_masked[7785];
  assign N6511 = N6510 | data_masked[7913];
  assign N6510 = data_masked[8169] | data_masked[8041];
  assign data_o[106] = N6633 | data_masked[106];
  assign N6633 = N6632 | data_masked[234];
  assign N6632 = N6631 | data_masked[362];
  assign N6631 = N6630 | data_masked[490];
  assign N6630 = N6629 | data_masked[618];
  assign N6629 = N6628 | data_masked[746];
  assign N6628 = N6627 | data_masked[874];
  assign N6627 = N6626 | data_masked[1002];
  assign N6626 = N6625 | data_masked[1130];
  assign N6625 = N6624 | data_masked[1258];
  assign N6624 = N6623 | data_masked[1386];
  assign N6623 = N6622 | data_masked[1514];
  assign N6622 = N6621 | data_masked[1642];
  assign N6621 = N6620 | data_masked[1770];
  assign N6620 = N6619 | data_masked[1898];
  assign N6619 = N6618 | data_masked[2026];
  assign N6618 = N6617 | data_masked[2154];
  assign N6617 = N6616 | data_masked[2282];
  assign N6616 = N6615 | data_masked[2410];
  assign N6615 = N6614 | data_masked[2538];
  assign N6614 = N6613 | data_masked[2666];
  assign N6613 = N6612 | data_masked[2794];
  assign N6612 = N6611 | data_masked[2922];
  assign N6611 = N6610 | data_masked[3050];
  assign N6610 = N6609 | data_masked[3178];
  assign N6609 = N6608 | data_masked[3306];
  assign N6608 = N6607 | data_masked[3434];
  assign N6607 = N6606 | data_masked[3562];
  assign N6606 = N6605 | data_masked[3690];
  assign N6605 = N6604 | data_masked[3818];
  assign N6604 = N6603 | data_masked[3946];
  assign N6603 = N6602 | data_masked[4074];
  assign N6602 = N6601 | data_masked[4202];
  assign N6601 = N6600 | data_masked[4330];
  assign N6600 = N6599 | data_masked[4458];
  assign N6599 = N6598 | data_masked[4586];
  assign N6598 = N6597 | data_masked[4714];
  assign N6597 = N6596 | data_masked[4842];
  assign N6596 = N6595 | data_masked[4970];
  assign N6595 = N6594 | data_masked[5098];
  assign N6594 = N6593 | data_masked[5226];
  assign N6593 = N6592 | data_masked[5354];
  assign N6592 = N6591 | data_masked[5482];
  assign N6591 = N6590 | data_masked[5610];
  assign N6590 = N6589 | data_masked[5738];
  assign N6589 = N6588 | data_masked[5866];
  assign N6588 = N6587 | data_masked[5994];
  assign N6587 = N6586 | data_masked[6122];
  assign N6586 = N6585 | data_masked[6250];
  assign N6585 = N6584 | data_masked[6378];
  assign N6584 = N6583 | data_masked[6506];
  assign N6583 = N6582 | data_masked[6634];
  assign N6582 = N6581 | data_masked[6762];
  assign N6581 = N6580 | data_masked[6890];
  assign N6580 = N6579 | data_masked[7018];
  assign N6579 = N6578 | data_masked[7146];
  assign N6578 = N6577 | data_masked[7274];
  assign N6577 = N6576 | data_masked[7402];
  assign N6576 = N6575 | data_masked[7530];
  assign N6575 = N6574 | data_masked[7658];
  assign N6574 = N6573 | data_masked[7786];
  assign N6573 = N6572 | data_masked[7914];
  assign N6572 = data_masked[8170] | data_masked[8042];
  assign data_o[107] = N6695 | data_masked[107];
  assign N6695 = N6694 | data_masked[235];
  assign N6694 = N6693 | data_masked[363];
  assign N6693 = N6692 | data_masked[491];
  assign N6692 = N6691 | data_masked[619];
  assign N6691 = N6690 | data_masked[747];
  assign N6690 = N6689 | data_masked[875];
  assign N6689 = N6688 | data_masked[1003];
  assign N6688 = N6687 | data_masked[1131];
  assign N6687 = N6686 | data_masked[1259];
  assign N6686 = N6685 | data_masked[1387];
  assign N6685 = N6684 | data_masked[1515];
  assign N6684 = N6683 | data_masked[1643];
  assign N6683 = N6682 | data_masked[1771];
  assign N6682 = N6681 | data_masked[1899];
  assign N6681 = N6680 | data_masked[2027];
  assign N6680 = N6679 | data_masked[2155];
  assign N6679 = N6678 | data_masked[2283];
  assign N6678 = N6677 | data_masked[2411];
  assign N6677 = N6676 | data_masked[2539];
  assign N6676 = N6675 | data_masked[2667];
  assign N6675 = N6674 | data_masked[2795];
  assign N6674 = N6673 | data_masked[2923];
  assign N6673 = N6672 | data_masked[3051];
  assign N6672 = N6671 | data_masked[3179];
  assign N6671 = N6670 | data_masked[3307];
  assign N6670 = N6669 | data_masked[3435];
  assign N6669 = N6668 | data_masked[3563];
  assign N6668 = N6667 | data_masked[3691];
  assign N6667 = N6666 | data_masked[3819];
  assign N6666 = N6665 | data_masked[3947];
  assign N6665 = N6664 | data_masked[4075];
  assign N6664 = N6663 | data_masked[4203];
  assign N6663 = N6662 | data_masked[4331];
  assign N6662 = N6661 | data_masked[4459];
  assign N6661 = N6660 | data_masked[4587];
  assign N6660 = N6659 | data_masked[4715];
  assign N6659 = N6658 | data_masked[4843];
  assign N6658 = N6657 | data_masked[4971];
  assign N6657 = N6656 | data_masked[5099];
  assign N6656 = N6655 | data_masked[5227];
  assign N6655 = N6654 | data_masked[5355];
  assign N6654 = N6653 | data_masked[5483];
  assign N6653 = N6652 | data_masked[5611];
  assign N6652 = N6651 | data_masked[5739];
  assign N6651 = N6650 | data_masked[5867];
  assign N6650 = N6649 | data_masked[5995];
  assign N6649 = N6648 | data_masked[6123];
  assign N6648 = N6647 | data_masked[6251];
  assign N6647 = N6646 | data_masked[6379];
  assign N6646 = N6645 | data_masked[6507];
  assign N6645 = N6644 | data_masked[6635];
  assign N6644 = N6643 | data_masked[6763];
  assign N6643 = N6642 | data_masked[6891];
  assign N6642 = N6641 | data_masked[7019];
  assign N6641 = N6640 | data_masked[7147];
  assign N6640 = N6639 | data_masked[7275];
  assign N6639 = N6638 | data_masked[7403];
  assign N6638 = N6637 | data_masked[7531];
  assign N6637 = N6636 | data_masked[7659];
  assign N6636 = N6635 | data_masked[7787];
  assign N6635 = N6634 | data_masked[7915];
  assign N6634 = data_masked[8171] | data_masked[8043];
  assign data_o[108] = N6757 | data_masked[108];
  assign N6757 = N6756 | data_masked[236];
  assign N6756 = N6755 | data_masked[364];
  assign N6755 = N6754 | data_masked[492];
  assign N6754 = N6753 | data_masked[620];
  assign N6753 = N6752 | data_masked[748];
  assign N6752 = N6751 | data_masked[876];
  assign N6751 = N6750 | data_masked[1004];
  assign N6750 = N6749 | data_masked[1132];
  assign N6749 = N6748 | data_masked[1260];
  assign N6748 = N6747 | data_masked[1388];
  assign N6747 = N6746 | data_masked[1516];
  assign N6746 = N6745 | data_masked[1644];
  assign N6745 = N6744 | data_masked[1772];
  assign N6744 = N6743 | data_masked[1900];
  assign N6743 = N6742 | data_masked[2028];
  assign N6742 = N6741 | data_masked[2156];
  assign N6741 = N6740 | data_masked[2284];
  assign N6740 = N6739 | data_masked[2412];
  assign N6739 = N6738 | data_masked[2540];
  assign N6738 = N6737 | data_masked[2668];
  assign N6737 = N6736 | data_masked[2796];
  assign N6736 = N6735 | data_masked[2924];
  assign N6735 = N6734 | data_masked[3052];
  assign N6734 = N6733 | data_masked[3180];
  assign N6733 = N6732 | data_masked[3308];
  assign N6732 = N6731 | data_masked[3436];
  assign N6731 = N6730 | data_masked[3564];
  assign N6730 = N6729 | data_masked[3692];
  assign N6729 = N6728 | data_masked[3820];
  assign N6728 = N6727 | data_masked[3948];
  assign N6727 = N6726 | data_masked[4076];
  assign N6726 = N6725 | data_masked[4204];
  assign N6725 = N6724 | data_masked[4332];
  assign N6724 = N6723 | data_masked[4460];
  assign N6723 = N6722 | data_masked[4588];
  assign N6722 = N6721 | data_masked[4716];
  assign N6721 = N6720 | data_masked[4844];
  assign N6720 = N6719 | data_masked[4972];
  assign N6719 = N6718 | data_masked[5100];
  assign N6718 = N6717 | data_masked[5228];
  assign N6717 = N6716 | data_masked[5356];
  assign N6716 = N6715 | data_masked[5484];
  assign N6715 = N6714 | data_masked[5612];
  assign N6714 = N6713 | data_masked[5740];
  assign N6713 = N6712 | data_masked[5868];
  assign N6712 = N6711 | data_masked[5996];
  assign N6711 = N6710 | data_masked[6124];
  assign N6710 = N6709 | data_masked[6252];
  assign N6709 = N6708 | data_masked[6380];
  assign N6708 = N6707 | data_masked[6508];
  assign N6707 = N6706 | data_masked[6636];
  assign N6706 = N6705 | data_masked[6764];
  assign N6705 = N6704 | data_masked[6892];
  assign N6704 = N6703 | data_masked[7020];
  assign N6703 = N6702 | data_masked[7148];
  assign N6702 = N6701 | data_masked[7276];
  assign N6701 = N6700 | data_masked[7404];
  assign N6700 = N6699 | data_masked[7532];
  assign N6699 = N6698 | data_masked[7660];
  assign N6698 = N6697 | data_masked[7788];
  assign N6697 = N6696 | data_masked[7916];
  assign N6696 = data_masked[8172] | data_masked[8044];
  assign data_o[109] = N6819 | data_masked[109];
  assign N6819 = N6818 | data_masked[237];
  assign N6818 = N6817 | data_masked[365];
  assign N6817 = N6816 | data_masked[493];
  assign N6816 = N6815 | data_masked[621];
  assign N6815 = N6814 | data_masked[749];
  assign N6814 = N6813 | data_masked[877];
  assign N6813 = N6812 | data_masked[1005];
  assign N6812 = N6811 | data_masked[1133];
  assign N6811 = N6810 | data_masked[1261];
  assign N6810 = N6809 | data_masked[1389];
  assign N6809 = N6808 | data_masked[1517];
  assign N6808 = N6807 | data_masked[1645];
  assign N6807 = N6806 | data_masked[1773];
  assign N6806 = N6805 | data_masked[1901];
  assign N6805 = N6804 | data_masked[2029];
  assign N6804 = N6803 | data_masked[2157];
  assign N6803 = N6802 | data_masked[2285];
  assign N6802 = N6801 | data_masked[2413];
  assign N6801 = N6800 | data_masked[2541];
  assign N6800 = N6799 | data_masked[2669];
  assign N6799 = N6798 | data_masked[2797];
  assign N6798 = N6797 | data_masked[2925];
  assign N6797 = N6796 | data_masked[3053];
  assign N6796 = N6795 | data_masked[3181];
  assign N6795 = N6794 | data_masked[3309];
  assign N6794 = N6793 | data_masked[3437];
  assign N6793 = N6792 | data_masked[3565];
  assign N6792 = N6791 | data_masked[3693];
  assign N6791 = N6790 | data_masked[3821];
  assign N6790 = N6789 | data_masked[3949];
  assign N6789 = N6788 | data_masked[4077];
  assign N6788 = N6787 | data_masked[4205];
  assign N6787 = N6786 | data_masked[4333];
  assign N6786 = N6785 | data_masked[4461];
  assign N6785 = N6784 | data_masked[4589];
  assign N6784 = N6783 | data_masked[4717];
  assign N6783 = N6782 | data_masked[4845];
  assign N6782 = N6781 | data_masked[4973];
  assign N6781 = N6780 | data_masked[5101];
  assign N6780 = N6779 | data_masked[5229];
  assign N6779 = N6778 | data_masked[5357];
  assign N6778 = N6777 | data_masked[5485];
  assign N6777 = N6776 | data_masked[5613];
  assign N6776 = N6775 | data_masked[5741];
  assign N6775 = N6774 | data_masked[5869];
  assign N6774 = N6773 | data_masked[5997];
  assign N6773 = N6772 | data_masked[6125];
  assign N6772 = N6771 | data_masked[6253];
  assign N6771 = N6770 | data_masked[6381];
  assign N6770 = N6769 | data_masked[6509];
  assign N6769 = N6768 | data_masked[6637];
  assign N6768 = N6767 | data_masked[6765];
  assign N6767 = N6766 | data_masked[6893];
  assign N6766 = N6765 | data_masked[7021];
  assign N6765 = N6764 | data_masked[7149];
  assign N6764 = N6763 | data_masked[7277];
  assign N6763 = N6762 | data_masked[7405];
  assign N6762 = N6761 | data_masked[7533];
  assign N6761 = N6760 | data_masked[7661];
  assign N6760 = N6759 | data_masked[7789];
  assign N6759 = N6758 | data_masked[7917];
  assign N6758 = data_masked[8173] | data_masked[8045];
  assign data_o[110] = N6881 | data_masked[110];
  assign N6881 = N6880 | data_masked[238];
  assign N6880 = N6879 | data_masked[366];
  assign N6879 = N6878 | data_masked[494];
  assign N6878 = N6877 | data_masked[622];
  assign N6877 = N6876 | data_masked[750];
  assign N6876 = N6875 | data_masked[878];
  assign N6875 = N6874 | data_masked[1006];
  assign N6874 = N6873 | data_masked[1134];
  assign N6873 = N6872 | data_masked[1262];
  assign N6872 = N6871 | data_masked[1390];
  assign N6871 = N6870 | data_masked[1518];
  assign N6870 = N6869 | data_masked[1646];
  assign N6869 = N6868 | data_masked[1774];
  assign N6868 = N6867 | data_masked[1902];
  assign N6867 = N6866 | data_masked[2030];
  assign N6866 = N6865 | data_masked[2158];
  assign N6865 = N6864 | data_masked[2286];
  assign N6864 = N6863 | data_masked[2414];
  assign N6863 = N6862 | data_masked[2542];
  assign N6862 = N6861 | data_masked[2670];
  assign N6861 = N6860 | data_masked[2798];
  assign N6860 = N6859 | data_masked[2926];
  assign N6859 = N6858 | data_masked[3054];
  assign N6858 = N6857 | data_masked[3182];
  assign N6857 = N6856 | data_masked[3310];
  assign N6856 = N6855 | data_masked[3438];
  assign N6855 = N6854 | data_masked[3566];
  assign N6854 = N6853 | data_masked[3694];
  assign N6853 = N6852 | data_masked[3822];
  assign N6852 = N6851 | data_masked[3950];
  assign N6851 = N6850 | data_masked[4078];
  assign N6850 = N6849 | data_masked[4206];
  assign N6849 = N6848 | data_masked[4334];
  assign N6848 = N6847 | data_masked[4462];
  assign N6847 = N6846 | data_masked[4590];
  assign N6846 = N6845 | data_masked[4718];
  assign N6845 = N6844 | data_masked[4846];
  assign N6844 = N6843 | data_masked[4974];
  assign N6843 = N6842 | data_masked[5102];
  assign N6842 = N6841 | data_masked[5230];
  assign N6841 = N6840 | data_masked[5358];
  assign N6840 = N6839 | data_masked[5486];
  assign N6839 = N6838 | data_masked[5614];
  assign N6838 = N6837 | data_masked[5742];
  assign N6837 = N6836 | data_masked[5870];
  assign N6836 = N6835 | data_masked[5998];
  assign N6835 = N6834 | data_masked[6126];
  assign N6834 = N6833 | data_masked[6254];
  assign N6833 = N6832 | data_masked[6382];
  assign N6832 = N6831 | data_masked[6510];
  assign N6831 = N6830 | data_masked[6638];
  assign N6830 = N6829 | data_masked[6766];
  assign N6829 = N6828 | data_masked[6894];
  assign N6828 = N6827 | data_masked[7022];
  assign N6827 = N6826 | data_masked[7150];
  assign N6826 = N6825 | data_masked[7278];
  assign N6825 = N6824 | data_masked[7406];
  assign N6824 = N6823 | data_masked[7534];
  assign N6823 = N6822 | data_masked[7662];
  assign N6822 = N6821 | data_masked[7790];
  assign N6821 = N6820 | data_masked[7918];
  assign N6820 = data_masked[8174] | data_masked[8046];
  assign data_o[111] = N6943 | data_masked[111];
  assign N6943 = N6942 | data_masked[239];
  assign N6942 = N6941 | data_masked[367];
  assign N6941 = N6940 | data_masked[495];
  assign N6940 = N6939 | data_masked[623];
  assign N6939 = N6938 | data_masked[751];
  assign N6938 = N6937 | data_masked[879];
  assign N6937 = N6936 | data_masked[1007];
  assign N6936 = N6935 | data_masked[1135];
  assign N6935 = N6934 | data_masked[1263];
  assign N6934 = N6933 | data_masked[1391];
  assign N6933 = N6932 | data_masked[1519];
  assign N6932 = N6931 | data_masked[1647];
  assign N6931 = N6930 | data_masked[1775];
  assign N6930 = N6929 | data_masked[1903];
  assign N6929 = N6928 | data_masked[2031];
  assign N6928 = N6927 | data_masked[2159];
  assign N6927 = N6926 | data_masked[2287];
  assign N6926 = N6925 | data_masked[2415];
  assign N6925 = N6924 | data_masked[2543];
  assign N6924 = N6923 | data_masked[2671];
  assign N6923 = N6922 | data_masked[2799];
  assign N6922 = N6921 | data_masked[2927];
  assign N6921 = N6920 | data_masked[3055];
  assign N6920 = N6919 | data_masked[3183];
  assign N6919 = N6918 | data_masked[3311];
  assign N6918 = N6917 | data_masked[3439];
  assign N6917 = N6916 | data_masked[3567];
  assign N6916 = N6915 | data_masked[3695];
  assign N6915 = N6914 | data_masked[3823];
  assign N6914 = N6913 | data_masked[3951];
  assign N6913 = N6912 | data_masked[4079];
  assign N6912 = N6911 | data_masked[4207];
  assign N6911 = N6910 | data_masked[4335];
  assign N6910 = N6909 | data_masked[4463];
  assign N6909 = N6908 | data_masked[4591];
  assign N6908 = N6907 | data_masked[4719];
  assign N6907 = N6906 | data_masked[4847];
  assign N6906 = N6905 | data_masked[4975];
  assign N6905 = N6904 | data_masked[5103];
  assign N6904 = N6903 | data_masked[5231];
  assign N6903 = N6902 | data_masked[5359];
  assign N6902 = N6901 | data_masked[5487];
  assign N6901 = N6900 | data_masked[5615];
  assign N6900 = N6899 | data_masked[5743];
  assign N6899 = N6898 | data_masked[5871];
  assign N6898 = N6897 | data_masked[5999];
  assign N6897 = N6896 | data_masked[6127];
  assign N6896 = N6895 | data_masked[6255];
  assign N6895 = N6894 | data_masked[6383];
  assign N6894 = N6893 | data_masked[6511];
  assign N6893 = N6892 | data_masked[6639];
  assign N6892 = N6891 | data_masked[6767];
  assign N6891 = N6890 | data_masked[6895];
  assign N6890 = N6889 | data_masked[7023];
  assign N6889 = N6888 | data_masked[7151];
  assign N6888 = N6887 | data_masked[7279];
  assign N6887 = N6886 | data_masked[7407];
  assign N6886 = N6885 | data_masked[7535];
  assign N6885 = N6884 | data_masked[7663];
  assign N6884 = N6883 | data_masked[7791];
  assign N6883 = N6882 | data_masked[7919];
  assign N6882 = data_masked[8175] | data_masked[8047];
  assign data_o[112] = N7005 | data_masked[112];
  assign N7005 = N7004 | data_masked[240];
  assign N7004 = N7003 | data_masked[368];
  assign N7003 = N7002 | data_masked[496];
  assign N7002 = N7001 | data_masked[624];
  assign N7001 = N7000 | data_masked[752];
  assign N7000 = N6999 | data_masked[880];
  assign N6999 = N6998 | data_masked[1008];
  assign N6998 = N6997 | data_masked[1136];
  assign N6997 = N6996 | data_masked[1264];
  assign N6996 = N6995 | data_masked[1392];
  assign N6995 = N6994 | data_masked[1520];
  assign N6994 = N6993 | data_masked[1648];
  assign N6993 = N6992 | data_masked[1776];
  assign N6992 = N6991 | data_masked[1904];
  assign N6991 = N6990 | data_masked[2032];
  assign N6990 = N6989 | data_masked[2160];
  assign N6989 = N6988 | data_masked[2288];
  assign N6988 = N6987 | data_masked[2416];
  assign N6987 = N6986 | data_masked[2544];
  assign N6986 = N6985 | data_masked[2672];
  assign N6985 = N6984 | data_masked[2800];
  assign N6984 = N6983 | data_masked[2928];
  assign N6983 = N6982 | data_masked[3056];
  assign N6982 = N6981 | data_masked[3184];
  assign N6981 = N6980 | data_masked[3312];
  assign N6980 = N6979 | data_masked[3440];
  assign N6979 = N6978 | data_masked[3568];
  assign N6978 = N6977 | data_masked[3696];
  assign N6977 = N6976 | data_masked[3824];
  assign N6976 = N6975 | data_masked[3952];
  assign N6975 = N6974 | data_masked[4080];
  assign N6974 = N6973 | data_masked[4208];
  assign N6973 = N6972 | data_masked[4336];
  assign N6972 = N6971 | data_masked[4464];
  assign N6971 = N6970 | data_masked[4592];
  assign N6970 = N6969 | data_masked[4720];
  assign N6969 = N6968 | data_masked[4848];
  assign N6968 = N6967 | data_masked[4976];
  assign N6967 = N6966 | data_masked[5104];
  assign N6966 = N6965 | data_masked[5232];
  assign N6965 = N6964 | data_masked[5360];
  assign N6964 = N6963 | data_masked[5488];
  assign N6963 = N6962 | data_masked[5616];
  assign N6962 = N6961 | data_masked[5744];
  assign N6961 = N6960 | data_masked[5872];
  assign N6960 = N6959 | data_masked[6000];
  assign N6959 = N6958 | data_masked[6128];
  assign N6958 = N6957 | data_masked[6256];
  assign N6957 = N6956 | data_masked[6384];
  assign N6956 = N6955 | data_masked[6512];
  assign N6955 = N6954 | data_masked[6640];
  assign N6954 = N6953 | data_masked[6768];
  assign N6953 = N6952 | data_masked[6896];
  assign N6952 = N6951 | data_masked[7024];
  assign N6951 = N6950 | data_masked[7152];
  assign N6950 = N6949 | data_masked[7280];
  assign N6949 = N6948 | data_masked[7408];
  assign N6948 = N6947 | data_masked[7536];
  assign N6947 = N6946 | data_masked[7664];
  assign N6946 = N6945 | data_masked[7792];
  assign N6945 = N6944 | data_masked[7920];
  assign N6944 = data_masked[8176] | data_masked[8048];
  assign data_o[113] = N7067 | data_masked[113];
  assign N7067 = N7066 | data_masked[241];
  assign N7066 = N7065 | data_masked[369];
  assign N7065 = N7064 | data_masked[497];
  assign N7064 = N7063 | data_masked[625];
  assign N7063 = N7062 | data_masked[753];
  assign N7062 = N7061 | data_masked[881];
  assign N7061 = N7060 | data_masked[1009];
  assign N7060 = N7059 | data_masked[1137];
  assign N7059 = N7058 | data_masked[1265];
  assign N7058 = N7057 | data_masked[1393];
  assign N7057 = N7056 | data_masked[1521];
  assign N7056 = N7055 | data_masked[1649];
  assign N7055 = N7054 | data_masked[1777];
  assign N7054 = N7053 | data_masked[1905];
  assign N7053 = N7052 | data_masked[2033];
  assign N7052 = N7051 | data_masked[2161];
  assign N7051 = N7050 | data_masked[2289];
  assign N7050 = N7049 | data_masked[2417];
  assign N7049 = N7048 | data_masked[2545];
  assign N7048 = N7047 | data_masked[2673];
  assign N7047 = N7046 | data_masked[2801];
  assign N7046 = N7045 | data_masked[2929];
  assign N7045 = N7044 | data_masked[3057];
  assign N7044 = N7043 | data_masked[3185];
  assign N7043 = N7042 | data_masked[3313];
  assign N7042 = N7041 | data_masked[3441];
  assign N7041 = N7040 | data_masked[3569];
  assign N7040 = N7039 | data_masked[3697];
  assign N7039 = N7038 | data_masked[3825];
  assign N7038 = N7037 | data_masked[3953];
  assign N7037 = N7036 | data_masked[4081];
  assign N7036 = N7035 | data_masked[4209];
  assign N7035 = N7034 | data_masked[4337];
  assign N7034 = N7033 | data_masked[4465];
  assign N7033 = N7032 | data_masked[4593];
  assign N7032 = N7031 | data_masked[4721];
  assign N7031 = N7030 | data_masked[4849];
  assign N7030 = N7029 | data_masked[4977];
  assign N7029 = N7028 | data_masked[5105];
  assign N7028 = N7027 | data_masked[5233];
  assign N7027 = N7026 | data_masked[5361];
  assign N7026 = N7025 | data_masked[5489];
  assign N7025 = N7024 | data_masked[5617];
  assign N7024 = N7023 | data_masked[5745];
  assign N7023 = N7022 | data_masked[5873];
  assign N7022 = N7021 | data_masked[6001];
  assign N7021 = N7020 | data_masked[6129];
  assign N7020 = N7019 | data_masked[6257];
  assign N7019 = N7018 | data_masked[6385];
  assign N7018 = N7017 | data_masked[6513];
  assign N7017 = N7016 | data_masked[6641];
  assign N7016 = N7015 | data_masked[6769];
  assign N7015 = N7014 | data_masked[6897];
  assign N7014 = N7013 | data_masked[7025];
  assign N7013 = N7012 | data_masked[7153];
  assign N7012 = N7011 | data_masked[7281];
  assign N7011 = N7010 | data_masked[7409];
  assign N7010 = N7009 | data_masked[7537];
  assign N7009 = N7008 | data_masked[7665];
  assign N7008 = N7007 | data_masked[7793];
  assign N7007 = N7006 | data_masked[7921];
  assign N7006 = data_masked[8177] | data_masked[8049];
  assign data_o[114] = N7129 | data_masked[114];
  assign N7129 = N7128 | data_masked[242];
  assign N7128 = N7127 | data_masked[370];
  assign N7127 = N7126 | data_masked[498];
  assign N7126 = N7125 | data_masked[626];
  assign N7125 = N7124 | data_masked[754];
  assign N7124 = N7123 | data_masked[882];
  assign N7123 = N7122 | data_masked[1010];
  assign N7122 = N7121 | data_masked[1138];
  assign N7121 = N7120 | data_masked[1266];
  assign N7120 = N7119 | data_masked[1394];
  assign N7119 = N7118 | data_masked[1522];
  assign N7118 = N7117 | data_masked[1650];
  assign N7117 = N7116 | data_masked[1778];
  assign N7116 = N7115 | data_masked[1906];
  assign N7115 = N7114 | data_masked[2034];
  assign N7114 = N7113 | data_masked[2162];
  assign N7113 = N7112 | data_masked[2290];
  assign N7112 = N7111 | data_masked[2418];
  assign N7111 = N7110 | data_masked[2546];
  assign N7110 = N7109 | data_masked[2674];
  assign N7109 = N7108 | data_masked[2802];
  assign N7108 = N7107 | data_masked[2930];
  assign N7107 = N7106 | data_masked[3058];
  assign N7106 = N7105 | data_masked[3186];
  assign N7105 = N7104 | data_masked[3314];
  assign N7104 = N7103 | data_masked[3442];
  assign N7103 = N7102 | data_masked[3570];
  assign N7102 = N7101 | data_masked[3698];
  assign N7101 = N7100 | data_masked[3826];
  assign N7100 = N7099 | data_masked[3954];
  assign N7099 = N7098 | data_masked[4082];
  assign N7098 = N7097 | data_masked[4210];
  assign N7097 = N7096 | data_masked[4338];
  assign N7096 = N7095 | data_masked[4466];
  assign N7095 = N7094 | data_masked[4594];
  assign N7094 = N7093 | data_masked[4722];
  assign N7093 = N7092 | data_masked[4850];
  assign N7092 = N7091 | data_masked[4978];
  assign N7091 = N7090 | data_masked[5106];
  assign N7090 = N7089 | data_masked[5234];
  assign N7089 = N7088 | data_masked[5362];
  assign N7088 = N7087 | data_masked[5490];
  assign N7087 = N7086 | data_masked[5618];
  assign N7086 = N7085 | data_masked[5746];
  assign N7085 = N7084 | data_masked[5874];
  assign N7084 = N7083 | data_masked[6002];
  assign N7083 = N7082 | data_masked[6130];
  assign N7082 = N7081 | data_masked[6258];
  assign N7081 = N7080 | data_masked[6386];
  assign N7080 = N7079 | data_masked[6514];
  assign N7079 = N7078 | data_masked[6642];
  assign N7078 = N7077 | data_masked[6770];
  assign N7077 = N7076 | data_masked[6898];
  assign N7076 = N7075 | data_masked[7026];
  assign N7075 = N7074 | data_masked[7154];
  assign N7074 = N7073 | data_masked[7282];
  assign N7073 = N7072 | data_masked[7410];
  assign N7072 = N7071 | data_masked[7538];
  assign N7071 = N7070 | data_masked[7666];
  assign N7070 = N7069 | data_masked[7794];
  assign N7069 = N7068 | data_masked[7922];
  assign N7068 = data_masked[8178] | data_masked[8050];
  assign data_o[115] = N7191 | data_masked[115];
  assign N7191 = N7190 | data_masked[243];
  assign N7190 = N7189 | data_masked[371];
  assign N7189 = N7188 | data_masked[499];
  assign N7188 = N7187 | data_masked[627];
  assign N7187 = N7186 | data_masked[755];
  assign N7186 = N7185 | data_masked[883];
  assign N7185 = N7184 | data_masked[1011];
  assign N7184 = N7183 | data_masked[1139];
  assign N7183 = N7182 | data_masked[1267];
  assign N7182 = N7181 | data_masked[1395];
  assign N7181 = N7180 | data_masked[1523];
  assign N7180 = N7179 | data_masked[1651];
  assign N7179 = N7178 | data_masked[1779];
  assign N7178 = N7177 | data_masked[1907];
  assign N7177 = N7176 | data_masked[2035];
  assign N7176 = N7175 | data_masked[2163];
  assign N7175 = N7174 | data_masked[2291];
  assign N7174 = N7173 | data_masked[2419];
  assign N7173 = N7172 | data_masked[2547];
  assign N7172 = N7171 | data_masked[2675];
  assign N7171 = N7170 | data_masked[2803];
  assign N7170 = N7169 | data_masked[2931];
  assign N7169 = N7168 | data_masked[3059];
  assign N7168 = N7167 | data_masked[3187];
  assign N7167 = N7166 | data_masked[3315];
  assign N7166 = N7165 | data_masked[3443];
  assign N7165 = N7164 | data_masked[3571];
  assign N7164 = N7163 | data_masked[3699];
  assign N7163 = N7162 | data_masked[3827];
  assign N7162 = N7161 | data_masked[3955];
  assign N7161 = N7160 | data_masked[4083];
  assign N7160 = N7159 | data_masked[4211];
  assign N7159 = N7158 | data_masked[4339];
  assign N7158 = N7157 | data_masked[4467];
  assign N7157 = N7156 | data_masked[4595];
  assign N7156 = N7155 | data_masked[4723];
  assign N7155 = N7154 | data_masked[4851];
  assign N7154 = N7153 | data_masked[4979];
  assign N7153 = N7152 | data_masked[5107];
  assign N7152 = N7151 | data_masked[5235];
  assign N7151 = N7150 | data_masked[5363];
  assign N7150 = N7149 | data_masked[5491];
  assign N7149 = N7148 | data_masked[5619];
  assign N7148 = N7147 | data_masked[5747];
  assign N7147 = N7146 | data_masked[5875];
  assign N7146 = N7145 | data_masked[6003];
  assign N7145 = N7144 | data_masked[6131];
  assign N7144 = N7143 | data_masked[6259];
  assign N7143 = N7142 | data_masked[6387];
  assign N7142 = N7141 | data_masked[6515];
  assign N7141 = N7140 | data_masked[6643];
  assign N7140 = N7139 | data_masked[6771];
  assign N7139 = N7138 | data_masked[6899];
  assign N7138 = N7137 | data_masked[7027];
  assign N7137 = N7136 | data_masked[7155];
  assign N7136 = N7135 | data_masked[7283];
  assign N7135 = N7134 | data_masked[7411];
  assign N7134 = N7133 | data_masked[7539];
  assign N7133 = N7132 | data_masked[7667];
  assign N7132 = N7131 | data_masked[7795];
  assign N7131 = N7130 | data_masked[7923];
  assign N7130 = data_masked[8179] | data_masked[8051];
  assign data_o[116] = N7253 | data_masked[116];
  assign N7253 = N7252 | data_masked[244];
  assign N7252 = N7251 | data_masked[372];
  assign N7251 = N7250 | data_masked[500];
  assign N7250 = N7249 | data_masked[628];
  assign N7249 = N7248 | data_masked[756];
  assign N7248 = N7247 | data_masked[884];
  assign N7247 = N7246 | data_masked[1012];
  assign N7246 = N7245 | data_masked[1140];
  assign N7245 = N7244 | data_masked[1268];
  assign N7244 = N7243 | data_masked[1396];
  assign N7243 = N7242 | data_masked[1524];
  assign N7242 = N7241 | data_masked[1652];
  assign N7241 = N7240 | data_masked[1780];
  assign N7240 = N7239 | data_masked[1908];
  assign N7239 = N7238 | data_masked[2036];
  assign N7238 = N7237 | data_masked[2164];
  assign N7237 = N7236 | data_masked[2292];
  assign N7236 = N7235 | data_masked[2420];
  assign N7235 = N7234 | data_masked[2548];
  assign N7234 = N7233 | data_masked[2676];
  assign N7233 = N7232 | data_masked[2804];
  assign N7232 = N7231 | data_masked[2932];
  assign N7231 = N7230 | data_masked[3060];
  assign N7230 = N7229 | data_masked[3188];
  assign N7229 = N7228 | data_masked[3316];
  assign N7228 = N7227 | data_masked[3444];
  assign N7227 = N7226 | data_masked[3572];
  assign N7226 = N7225 | data_masked[3700];
  assign N7225 = N7224 | data_masked[3828];
  assign N7224 = N7223 | data_masked[3956];
  assign N7223 = N7222 | data_masked[4084];
  assign N7222 = N7221 | data_masked[4212];
  assign N7221 = N7220 | data_masked[4340];
  assign N7220 = N7219 | data_masked[4468];
  assign N7219 = N7218 | data_masked[4596];
  assign N7218 = N7217 | data_masked[4724];
  assign N7217 = N7216 | data_masked[4852];
  assign N7216 = N7215 | data_masked[4980];
  assign N7215 = N7214 | data_masked[5108];
  assign N7214 = N7213 | data_masked[5236];
  assign N7213 = N7212 | data_masked[5364];
  assign N7212 = N7211 | data_masked[5492];
  assign N7211 = N7210 | data_masked[5620];
  assign N7210 = N7209 | data_masked[5748];
  assign N7209 = N7208 | data_masked[5876];
  assign N7208 = N7207 | data_masked[6004];
  assign N7207 = N7206 | data_masked[6132];
  assign N7206 = N7205 | data_masked[6260];
  assign N7205 = N7204 | data_masked[6388];
  assign N7204 = N7203 | data_masked[6516];
  assign N7203 = N7202 | data_masked[6644];
  assign N7202 = N7201 | data_masked[6772];
  assign N7201 = N7200 | data_masked[6900];
  assign N7200 = N7199 | data_masked[7028];
  assign N7199 = N7198 | data_masked[7156];
  assign N7198 = N7197 | data_masked[7284];
  assign N7197 = N7196 | data_masked[7412];
  assign N7196 = N7195 | data_masked[7540];
  assign N7195 = N7194 | data_masked[7668];
  assign N7194 = N7193 | data_masked[7796];
  assign N7193 = N7192 | data_masked[7924];
  assign N7192 = data_masked[8180] | data_masked[8052];
  assign data_o[117] = N7315 | data_masked[117];
  assign N7315 = N7314 | data_masked[245];
  assign N7314 = N7313 | data_masked[373];
  assign N7313 = N7312 | data_masked[501];
  assign N7312 = N7311 | data_masked[629];
  assign N7311 = N7310 | data_masked[757];
  assign N7310 = N7309 | data_masked[885];
  assign N7309 = N7308 | data_masked[1013];
  assign N7308 = N7307 | data_masked[1141];
  assign N7307 = N7306 | data_masked[1269];
  assign N7306 = N7305 | data_masked[1397];
  assign N7305 = N7304 | data_masked[1525];
  assign N7304 = N7303 | data_masked[1653];
  assign N7303 = N7302 | data_masked[1781];
  assign N7302 = N7301 | data_masked[1909];
  assign N7301 = N7300 | data_masked[2037];
  assign N7300 = N7299 | data_masked[2165];
  assign N7299 = N7298 | data_masked[2293];
  assign N7298 = N7297 | data_masked[2421];
  assign N7297 = N7296 | data_masked[2549];
  assign N7296 = N7295 | data_masked[2677];
  assign N7295 = N7294 | data_masked[2805];
  assign N7294 = N7293 | data_masked[2933];
  assign N7293 = N7292 | data_masked[3061];
  assign N7292 = N7291 | data_masked[3189];
  assign N7291 = N7290 | data_masked[3317];
  assign N7290 = N7289 | data_masked[3445];
  assign N7289 = N7288 | data_masked[3573];
  assign N7288 = N7287 | data_masked[3701];
  assign N7287 = N7286 | data_masked[3829];
  assign N7286 = N7285 | data_masked[3957];
  assign N7285 = N7284 | data_masked[4085];
  assign N7284 = N7283 | data_masked[4213];
  assign N7283 = N7282 | data_masked[4341];
  assign N7282 = N7281 | data_masked[4469];
  assign N7281 = N7280 | data_masked[4597];
  assign N7280 = N7279 | data_masked[4725];
  assign N7279 = N7278 | data_masked[4853];
  assign N7278 = N7277 | data_masked[4981];
  assign N7277 = N7276 | data_masked[5109];
  assign N7276 = N7275 | data_masked[5237];
  assign N7275 = N7274 | data_masked[5365];
  assign N7274 = N7273 | data_masked[5493];
  assign N7273 = N7272 | data_masked[5621];
  assign N7272 = N7271 | data_masked[5749];
  assign N7271 = N7270 | data_masked[5877];
  assign N7270 = N7269 | data_masked[6005];
  assign N7269 = N7268 | data_masked[6133];
  assign N7268 = N7267 | data_masked[6261];
  assign N7267 = N7266 | data_masked[6389];
  assign N7266 = N7265 | data_masked[6517];
  assign N7265 = N7264 | data_masked[6645];
  assign N7264 = N7263 | data_masked[6773];
  assign N7263 = N7262 | data_masked[6901];
  assign N7262 = N7261 | data_masked[7029];
  assign N7261 = N7260 | data_masked[7157];
  assign N7260 = N7259 | data_masked[7285];
  assign N7259 = N7258 | data_masked[7413];
  assign N7258 = N7257 | data_masked[7541];
  assign N7257 = N7256 | data_masked[7669];
  assign N7256 = N7255 | data_masked[7797];
  assign N7255 = N7254 | data_masked[7925];
  assign N7254 = data_masked[8181] | data_masked[8053];
  assign data_o[118] = N7377 | data_masked[118];
  assign N7377 = N7376 | data_masked[246];
  assign N7376 = N7375 | data_masked[374];
  assign N7375 = N7374 | data_masked[502];
  assign N7374 = N7373 | data_masked[630];
  assign N7373 = N7372 | data_masked[758];
  assign N7372 = N7371 | data_masked[886];
  assign N7371 = N7370 | data_masked[1014];
  assign N7370 = N7369 | data_masked[1142];
  assign N7369 = N7368 | data_masked[1270];
  assign N7368 = N7367 | data_masked[1398];
  assign N7367 = N7366 | data_masked[1526];
  assign N7366 = N7365 | data_masked[1654];
  assign N7365 = N7364 | data_masked[1782];
  assign N7364 = N7363 | data_masked[1910];
  assign N7363 = N7362 | data_masked[2038];
  assign N7362 = N7361 | data_masked[2166];
  assign N7361 = N7360 | data_masked[2294];
  assign N7360 = N7359 | data_masked[2422];
  assign N7359 = N7358 | data_masked[2550];
  assign N7358 = N7357 | data_masked[2678];
  assign N7357 = N7356 | data_masked[2806];
  assign N7356 = N7355 | data_masked[2934];
  assign N7355 = N7354 | data_masked[3062];
  assign N7354 = N7353 | data_masked[3190];
  assign N7353 = N7352 | data_masked[3318];
  assign N7352 = N7351 | data_masked[3446];
  assign N7351 = N7350 | data_masked[3574];
  assign N7350 = N7349 | data_masked[3702];
  assign N7349 = N7348 | data_masked[3830];
  assign N7348 = N7347 | data_masked[3958];
  assign N7347 = N7346 | data_masked[4086];
  assign N7346 = N7345 | data_masked[4214];
  assign N7345 = N7344 | data_masked[4342];
  assign N7344 = N7343 | data_masked[4470];
  assign N7343 = N7342 | data_masked[4598];
  assign N7342 = N7341 | data_masked[4726];
  assign N7341 = N7340 | data_masked[4854];
  assign N7340 = N7339 | data_masked[4982];
  assign N7339 = N7338 | data_masked[5110];
  assign N7338 = N7337 | data_masked[5238];
  assign N7337 = N7336 | data_masked[5366];
  assign N7336 = N7335 | data_masked[5494];
  assign N7335 = N7334 | data_masked[5622];
  assign N7334 = N7333 | data_masked[5750];
  assign N7333 = N7332 | data_masked[5878];
  assign N7332 = N7331 | data_masked[6006];
  assign N7331 = N7330 | data_masked[6134];
  assign N7330 = N7329 | data_masked[6262];
  assign N7329 = N7328 | data_masked[6390];
  assign N7328 = N7327 | data_masked[6518];
  assign N7327 = N7326 | data_masked[6646];
  assign N7326 = N7325 | data_masked[6774];
  assign N7325 = N7324 | data_masked[6902];
  assign N7324 = N7323 | data_masked[7030];
  assign N7323 = N7322 | data_masked[7158];
  assign N7322 = N7321 | data_masked[7286];
  assign N7321 = N7320 | data_masked[7414];
  assign N7320 = N7319 | data_masked[7542];
  assign N7319 = N7318 | data_masked[7670];
  assign N7318 = N7317 | data_masked[7798];
  assign N7317 = N7316 | data_masked[7926];
  assign N7316 = data_masked[8182] | data_masked[8054];
  assign data_o[119] = N7439 | data_masked[119];
  assign N7439 = N7438 | data_masked[247];
  assign N7438 = N7437 | data_masked[375];
  assign N7437 = N7436 | data_masked[503];
  assign N7436 = N7435 | data_masked[631];
  assign N7435 = N7434 | data_masked[759];
  assign N7434 = N7433 | data_masked[887];
  assign N7433 = N7432 | data_masked[1015];
  assign N7432 = N7431 | data_masked[1143];
  assign N7431 = N7430 | data_masked[1271];
  assign N7430 = N7429 | data_masked[1399];
  assign N7429 = N7428 | data_masked[1527];
  assign N7428 = N7427 | data_masked[1655];
  assign N7427 = N7426 | data_masked[1783];
  assign N7426 = N7425 | data_masked[1911];
  assign N7425 = N7424 | data_masked[2039];
  assign N7424 = N7423 | data_masked[2167];
  assign N7423 = N7422 | data_masked[2295];
  assign N7422 = N7421 | data_masked[2423];
  assign N7421 = N7420 | data_masked[2551];
  assign N7420 = N7419 | data_masked[2679];
  assign N7419 = N7418 | data_masked[2807];
  assign N7418 = N7417 | data_masked[2935];
  assign N7417 = N7416 | data_masked[3063];
  assign N7416 = N7415 | data_masked[3191];
  assign N7415 = N7414 | data_masked[3319];
  assign N7414 = N7413 | data_masked[3447];
  assign N7413 = N7412 | data_masked[3575];
  assign N7412 = N7411 | data_masked[3703];
  assign N7411 = N7410 | data_masked[3831];
  assign N7410 = N7409 | data_masked[3959];
  assign N7409 = N7408 | data_masked[4087];
  assign N7408 = N7407 | data_masked[4215];
  assign N7407 = N7406 | data_masked[4343];
  assign N7406 = N7405 | data_masked[4471];
  assign N7405 = N7404 | data_masked[4599];
  assign N7404 = N7403 | data_masked[4727];
  assign N7403 = N7402 | data_masked[4855];
  assign N7402 = N7401 | data_masked[4983];
  assign N7401 = N7400 | data_masked[5111];
  assign N7400 = N7399 | data_masked[5239];
  assign N7399 = N7398 | data_masked[5367];
  assign N7398 = N7397 | data_masked[5495];
  assign N7397 = N7396 | data_masked[5623];
  assign N7396 = N7395 | data_masked[5751];
  assign N7395 = N7394 | data_masked[5879];
  assign N7394 = N7393 | data_masked[6007];
  assign N7393 = N7392 | data_masked[6135];
  assign N7392 = N7391 | data_masked[6263];
  assign N7391 = N7390 | data_masked[6391];
  assign N7390 = N7389 | data_masked[6519];
  assign N7389 = N7388 | data_masked[6647];
  assign N7388 = N7387 | data_masked[6775];
  assign N7387 = N7386 | data_masked[6903];
  assign N7386 = N7385 | data_masked[7031];
  assign N7385 = N7384 | data_masked[7159];
  assign N7384 = N7383 | data_masked[7287];
  assign N7383 = N7382 | data_masked[7415];
  assign N7382 = N7381 | data_masked[7543];
  assign N7381 = N7380 | data_masked[7671];
  assign N7380 = N7379 | data_masked[7799];
  assign N7379 = N7378 | data_masked[7927];
  assign N7378 = data_masked[8183] | data_masked[8055];
  assign data_o[120] = N7501 | data_masked[120];
  assign N7501 = N7500 | data_masked[248];
  assign N7500 = N7499 | data_masked[376];
  assign N7499 = N7498 | data_masked[504];
  assign N7498 = N7497 | data_masked[632];
  assign N7497 = N7496 | data_masked[760];
  assign N7496 = N7495 | data_masked[888];
  assign N7495 = N7494 | data_masked[1016];
  assign N7494 = N7493 | data_masked[1144];
  assign N7493 = N7492 | data_masked[1272];
  assign N7492 = N7491 | data_masked[1400];
  assign N7491 = N7490 | data_masked[1528];
  assign N7490 = N7489 | data_masked[1656];
  assign N7489 = N7488 | data_masked[1784];
  assign N7488 = N7487 | data_masked[1912];
  assign N7487 = N7486 | data_masked[2040];
  assign N7486 = N7485 | data_masked[2168];
  assign N7485 = N7484 | data_masked[2296];
  assign N7484 = N7483 | data_masked[2424];
  assign N7483 = N7482 | data_masked[2552];
  assign N7482 = N7481 | data_masked[2680];
  assign N7481 = N7480 | data_masked[2808];
  assign N7480 = N7479 | data_masked[2936];
  assign N7479 = N7478 | data_masked[3064];
  assign N7478 = N7477 | data_masked[3192];
  assign N7477 = N7476 | data_masked[3320];
  assign N7476 = N7475 | data_masked[3448];
  assign N7475 = N7474 | data_masked[3576];
  assign N7474 = N7473 | data_masked[3704];
  assign N7473 = N7472 | data_masked[3832];
  assign N7472 = N7471 | data_masked[3960];
  assign N7471 = N7470 | data_masked[4088];
  assign N7470 = N7469 | data_masked[4216];
  assign N7469 = N7468 | data_masked[4344];
  assign N7468 = N7467 | data_masked[4472];
  assign N7467 = N7466 | data_masked[4600];
  assign N7466 = N7465 | data_masked[4728];
  assign N7465 = N7464 | data_masked[4856];
  assign N7464 = N7463 | data_masked[4984];
  assign N7463 = N7462 | data_masked[5112];
  assign N7462 = N7461 | data_masked[5240];
  assign N7461 = N7460 | data_masked[5368];
  assign N7460 = N7459 | data_masked[5496];
  assign N7459 = N7458 | data_masked[5624];
  assign N7458 = N7457 | data_masked[5752];
  assign N7457 = N7456 | data_masked[5880];
  assign N7456 = N7455 | data_masked[6008];
  assign N7455 = N7454 | data_masked[6136];
  assign N7454 = N7453 | data_masked[6264];
  assign N7453 = N7452 | data_masked[6392];
  assign N7452 = N7451 | data_masked[6520];
  assign N7451 = N7450 | data_masked[6648];
  assign N7450 = N7449 | data_masked[6776];
  assign N7449 = N7448 | data_masked[6904];
  assign N7448 = N7447 | data_masked[7032];
  assign N7447 = N7446 | data_masked[7160];
  assign N7446 = N7445 | data_masked[7288];
  assign N7445 = N7444 | data_masked[7416];
  assign N7444 = N7443 | data_masked[7544];
  assign N7443 = N7442 | data_masked[7672];
  assign N7442 = N7441 | data_masked[7800];
  assign N7441 = N7440 | data_masked[7928];
  assign N7440 = data_masked[8184] | data_masked[8056];
  assign data_o[121] = N7563 | data_masked[121];
  assign N7563 = N7562 | data_masked[249];
  assign N7562 = N7561 | data_masked[377];
  assign N7561 = N7560 | data_masked[505];
  assign N7560 = N7559 | data_masked[633];
  assign N7559 = N7558 | data_masked[761];
  assign N7558 = N7557 | data_masked[889];
  assign N7557 = N7556 | data_masked[1017];
  assign N7556 = N7555 | data_masked[1145];
  assign N7555 = N7554 | data_masked[1273];
  assign N7554 = N7553 | data_masked[1401];
  assign N7553 = N7552 | data_masked[1529];
  assign N7552 = N7551 | data_masked[1657];
  assign N7551 = N7550 | data_masked[1785];
  assign N7550 = N7549 | data_masked[1913];
  assign N7549 = N7548 | data_masked[2041];
  assign N7548 = N7547 | data_masked[2169];
  assign N7547 = N7546 | data_masked[2297];
  assign N7546 = N7545 | data_masked[2425];
  assign N7545 = N7544 | data_masked[2553];
  assign N7544 = N7543 | data_masked[2681];
  assign N7543 = N7542 | data_masked[2809];
  assign N7542 = N7541 | data_masked[2937];
  assign N7541 = N7540 | data_masked[3065];
  assign N7540 = N7539 | data_masked[3193];
  assign N7539 = N7538 | data_masked[3321];
  assign N7538 = N7537 | data_masked[3449];
  assign N7537 = N7536 | data_masked[3577];
  assign N7536 = N7535 | data_masked[3705];
  assign N7535 = N7534 | data_masked[3833];
  assign N7534 = N7533 | data_masked[3961];
  assign N7533 = N7532 | data_masked[4089];
  assign N7532 = N7531 | data_masked[4217];
  assign N7531 = N7530 | data_masked[4345];
  assign N7530 = N7529 | data_masked[4473];
  assign N7529 = N7528 | data_masked[4601];
  assign N7528 = N7527 | data_masked[4729];
  assign N7527 = N7526 | data_masked[4857];
  assign N7526 = N7525 | data_masked[4985];
  assign N7525 = N7524 | data_masked[5113];
  assign N7524 = N7523 | data_masked[5241];
  assign N7523 = N7522 | data_masked[5369];
  assign N7522 = N7521 | data_masked[5497];
  assign N7521 = N7520 | data_masked[5625];
  assign N7520 = N7519 | data_masked[5753];
  assign N7519 = N7518 | data_masked[5881];
  assign N7518 = N7517 | data_masked[6009];
  assign N7517 = N7516 | data_masked[6137];
  assign N7516 = N7515 | data_masked[6265];
  assign N7515 = N7514 | data_masked[6393];
  assign N7514 = N7513 | data_masked[6521];
  assign N7513 = N7512 | data_masked[6649];
  assign N7512 = N7511 | data_masked[6777];
  assign N7511 = N7510 | data_masked[6905];
  assign N7510 = N7509 | data_masked[7033];
  assign N7509 = N7508 | data_masked[7161];
  assign N7508 = N7507 | data_masked[7289];
  assign N7507 = N7506 | data_masked[7417];
  assign N7506 = N7505 | data_masked[7545];
  assign N7505 = N7504 | data_masked[7673];
  assign N7504 = N7503 | data_masked[7801];
  assign N7503 = N7502 | data_masked[7929];
  assign N7502 = data_masked[8185] | data_masked[8057];
  assign data_o[122] = N7625 | data_masked[122];
  assign N7625 = N7624 | data_masked[250];
  assign N7624 = N7623 | data_masked[378];
  assign N7623 = N7622 | data_masked[506];
  assign N7622 = N7621 | data_masked[634];
  assign N7621 = N7620 | data_masked[762];
  assign N7620 = N7619 | data_masked[890];
  assign N7619 = N7618 | data_masked[1018];
  assign N7618 = N7617 | data_masked[1146];
  assign N7617 = N7616 | data_masked[1274];
  assign N7616 = N7615 | data_masked[1402];
  assign N7615 = N7614 | data_masked[1530];
  assign N7614 = N7613 | data_masked[1658];
  assign N7613 = N7612 | data_masked[1786];
  assign N7612 = N7611 | data_masked[1914];
  assign N7611 = N7610 | data_masked[2042];
  assign N7610 = N7609 | data_masked[2170];
  assign N7609 = N7608 | data_masked[2298];
  assign N7608 = N7607 | data_masked[2426];
  assign N7607 = N7606 | data_masked[2554];
  assign N7606 = N7605 | data_masked[2682];
  assign N7605 = N7604 | data_masked[2810];
  assign N7604 = N7603 | data_masked[2938];
  assign N7603 = N7602 | data_masked[3066];
  assign N7602 = N7601 | data_masked[3194];
  assign N7601 = N7600 | data_masked[3322];
  assign N7600 = N7599 | data_masked[3450];
  assign N7599 = N7598 | data_masked[3578];
  assign N7598 = N7597 | data_masked[3706];
  assign N7597 = N7596 | data_masked[3834];
  assign N7596 = N7595 | data_masked[3962];
  assign N7595 = N7594 | data_masked[4090];
  assign N7594 = N7593 | data_masked[4218];
  assign N7593 = N7592 | data_masked[4346];
  assign N7592 = N7591 | data_masked[4474];
  assign N7591 = N7590 | data_masked[4602];
  assign N7590 = N7589 | data_masked[4730];
  assign N7589 = N7588 | data_masked[4858];
  assign N7588 = N7587 | data_masked[4986];
  assign N7587 = N7586 | data_masked[5114];
  assign N7586 = N7585 | data_masked[5242];
  assign N7585 = N7584 | data_masked[5370];
  assign N7584 = N7583 | data_masked[5498];
  assign N7583 = N7582 | data_masked[5626];
  assign N7582 = N7581 | data_masked[5754];
  assign N7581 = N7580 | data_masked[5882];
  assign N7580 = N7579 | data_masked[6010];
  assign N7579 = N7578 | data_masked[6138];
  assign N7578 = N7577 | data_masked[6266];
  assign N7577 = N7576 | data_masked[6394];
  assign N7576 = N7575 | data_masked[6522];
  assign N7575 = N7574 | data_masked[6650];
  assign N7574 = N7573 | data_masked[6778];
  assign N7573 = N7572 | data_masked[6906];
  assign N7572 = N7571 | data_masked[7034];
  assign N7571 = N7570 | data_masked[7162];
  assign N7570 = N7569 | data_masked[7290];
  assign N7569 = N7568 | data_masked[7418];
  assign N7568 = N7567 | data_masked[7546];
  assign N7567 = N7566 | data_masked[7674];
  assign N7566 = N7565 | data_masked[7802];
  assign N7565 = N7564 | data_masked[7930];
  assign N7564 = data_masked[8186] | data_masked[8058];
  assign data_o[123] = N7687 | data_masked[123];
  assign N7687 = N7686 | data_masked[251];
  assign N7686 = N7685 | data_masked[379];
  assign N7685 = N7684 | data_masked[507];
  assign N7684 = N7683 | data_masked[635];
  assign N7683 = N7682 | data_masked[763];
  assign N7682 = N7681 | data_masked[891];
  assign N7681 = N7680 | data_masked[1019];
  assign N7680 = N7679 | data_masked[1147];
  assign N7679 = N7678 | data_masked[1275];
  assign N7678 = N7677 | data_masked[1403];
  assign N7677 = N7676 | data_masked[1531];
  assign N7676 = N7675 | data_masked[1659];
  assign N7675 = N7674 | data_masked[1787];
  assign N7674 = N7673 | data_masked[1915];
  assign N7673 = N7672 | data_masked[2043];
  assign N7672 = N7671 | data_masked[2171];
  assign N7671 = N7670 | data_masked[2299];
  assign N7670 = N7669 | data_masked[2427];
  assign N7669 = N7668 | data_masked[2555];
  assign N7668 = N7667 | data_masked[2683];
  assign N7667 = N7666 | data_masked[2811];
  assign N7666 = N7665 | data_masked[2939];
  assign N7665 = N7664 | data_masked[3067];
  assign N7664 = N7663 | data_masked[3195];
  assign N7663 = N7662 | data_masked[3323];
  assign N7662 = N7661 | data_masked[3451];
  assign N7661 = N7660 | data_masked[3579];
  assign N7660 = N7659 | data_masked[3707];
  assign N7659 = N7658 | data_masked[3835];
  assign N7658 = N7657 | data_masked[3963];
  assign N7657 = N7656 | data_masked[4091];
  assign N7656 = N7655 | data_masked[4219];
  assign N7655 = N7654 | data_masked[4347];
  assign N7654 = N7653 | data_masked[4475];
  assign N7653 = N7652 | data_masked[4603];
  assign N7652 = N7651 | data_masked[4731];
  assign N7651 = N7650 | data_masked[4859];
  assign N7650 = N7649 | data_masked[4987];
  assign N7649 = N7648 | data_masked[5115];
  assign N7648 = N7647 | data_masked[5243];
  assign N7647 = N7646 | data_masked[5371];
  assign N7646 = N7645 | data_masked[5499];
  assign N7645 = N7644 | data_masked[5627];
  assign N7644 = N7643 | data_masked[5755];
  assign N7643 = N7642 | data_masked[5883];
  assign N7642 = N7641 | data_masked[6011];
  assign N7641 = N7640 | data_masked[6139];
  assign N7640 = N7639 | data_masked[6267];
  assign N7639 = N7638 | data_masked[6395];
  assign N7638 = N7637 | data_masked[6523];
  assign N7637 = N7636 | data_masked[6651];
  assign N7636 = N7635 | data_masked[6779];
  assign N7635 = N7634 | data_masked[6907];
  assign N7634 = N7633 | data_masked[7035];
  assign N7633 = N7632 | data_masked[7163];
  assign N7632 = N7631 | data_masked[7291];
  assign N7631 = N7630 | data_masked[7419];
  assign N7630 = N7629 | data_masked[7547];
  assign N7629 = N7628 | data_masked[7675];
  assign N7628 = N7627 | data_masked[7803];
  assign N7627 = N7626 | data_masked[7931];
  assign N7626 = data_masked[8187] | data_masked[8059];
  assign data_o[124] = N7749 | data_masked[124];
  assign N7749 = N7748 | data_masked[252];
  assign N7748 = N7747 | data_masked[380];
  assign N7747 = N7746 | data_masked[508];
  assign N7746 = N7745 | data_masked[636];
  assign N7745 = N7744 | data_masked[764];
  assign N7744 = N7743 | data_masked[892];
  assign N7743 = N7742 | data_masked[1020];
  assign N7742 = N7741 | data_masked[1148];
  assign N7741 = N7740 | data_masked[1276];
  assign N7740 = N7739 | data_masked[1404];
  assign N7739 = N7738 | data_masked[1532];
  assign N7738 = N7737 | data_masked[1660];
  assign N7737 = N7736 | data_masked[1788];
  assign N7736 = N7735 | data_masked[1916];
  assign N7735 = N7734 | data_masked[2044];
  assign N7734 = N7733 | data_masked[2172];
  assign N7733 = N7732 | data_masked[2300];
  assign N7732 = N7731 | data_masked[2428];
  assign N7731 = N7730 | data_masked[2556];
  assign N7730 = N7729 | data_masked[2684];
  assign N7729 = N7728 | data_masked[2812];
  assign N7728 = N7727 | data_masked[2940];
  assign N7727 = N7726 | data_masked[3068];
  assign N7726 = N7725 | data_masked[3196];
  assign N7725 = N7724 | data_masked[3324];
  assign N7724 = N7723 | data_masked[3452];
  assign N7723 = N7722 | data_masked[3580];
  assign N7722 = N7721 | data_masked[3708];
  assign N7721 = N7720 | data_masked[3836];
  assign N7720 = N7719 | data_masked[3964];
  assign N7719 = N7718 | data_masked[4092];
  assign N7718 = N7717 | data_masked[4220];
  assign N7717 = N7716 | data_masked[4348];
  assign N7716 = N7715 | data_masked[4476];
  assign N7715 = N7714 | data_masked[4604];
  assign N7714 = N7713 | data_masked[4732];
  assign N7713 = N7712 | data_masked[4860];
  assign N7712 = N7711 | data_masked[4988];
  assign N7711 = N7710 | data_masked[5116];
  assign N7710 = N7709 | data_masked[5244];
  assign N7709 = N7708 | data_masked[5372];
  assign N7708 = N7707 | data_masked[5500];
  assign N7707 = N7706 | data_masked[5628];
  assign N7706 = N7705 | data_masked[5756];
  assign N7705 = N7704 | data_masked[5884];
  assign N7704 = N7703 | data_masked[6012];
  assign N7703 = N7702 | data_masked[6140];
  assign N7702 = N7701 | data_masked[6268];
  assign N7701 = N7700 | data_masked[6396];
  assign N7700 = N7699 | data_masked[6524];
  assign N7699 = N7698 | data_masked[6652];
  assign N7698 = N7697 | data_masked[6780];
  assign N7697 = N7696 | data_masked[6908];
  assign N7696 = N7695 | data_masked[7036];
  assign N7695 = N7694 | data_masked[7164];
  assign N7694 = N7693 | data_masked[7292];
  assign N7693 = N7692 | data_masked[7420];
  assign N7692 = N7691 | data_masked[7548];
  assign N7691 = N7690 | data_masked[7676];
  assign N7690 = N7689 | data_masked[7804];
  assign N7689 = N7688 | data_masked[7932];
  assign N7688 = data_masked[8188] | data_masked[8060];
  assign data_o[125] = N7811 | data_masked[125];
  assign N7811 = N7810 | data_masked[253];
  assign N7810 = N7809 | data_masked[381];
  assign N7809 = N7808 | data_masked[509];
  assign N7808 = N7807 | data_masked[637];
  assign N7807 = N7806 | data_masked[765];
  assign N7806 = N7805 | data_masked[893];
  assign N7805 = N7804 | data_masked[1021];
  assign N7804 = N7803 | data_masked[1149];
  assign N7803 = N7802 | data_masked[1277];
  assign N7802 = N7801 | data_masked[1405];
  assign N7801 = N7800 | data_masked[1533];
  assign N7800 = N7799 | data_masked[1661];
  assign N7799 = N7798 | data_masked[1789];
  assign N7798 = N7797 | data_masked[1917];
  assign N7797 = N7796 | data_masked[2045];
  assign N7796 = N7795 | data_masked[2173];
  assign N7795 = N7794 | data_masked[2301];
  assign N7794 = N7793 | data_masked[2429];
  assign N7793 = N7792 | data_masked[2557];
  assign N7792 = N7791 | data_masked[2685];
  assign N7791 = N7790 | data_masked[2813];
  assign N7790 = N7789 | data_masked[2941];
  assign N7789 = N7788 | data_masked[3069];
  assign N7788 = N7787 | data_masked[3197];
  assign N7787 = N7786 | data_masked[3325];
  assign N7786 = N7785 | data_masked[3453];
  assign N7785 = N7784 | data_masked[3581];
  assign N7784 = N7783 | data_masked[3709];
  assign N7783 = N7782 | data_masked[3837];
  assign N7782 = N7781 | data_masked[3965];
  assign N7781 = N7780 | data_masked[4093];
  assign N7780 = N7779 | data_masked[4221];
  assign N7779 = N7778 | data_masked[4349];
  assign N7778 = N7777 | data_masked[4477];
  assign N7777 = N7776 | data_masked[4605];
  assign N7776 = N7775 | data_masked[4733];
  assign N7775 = N7774 | data_masked[4861];
  assign N7774 = N7773 | data_masked[4989];
  assign N7773 = N7772 | data_masked[5117];
  assign N7772 = N7771 | data_masked[5245];
  assign N7771 = N7770 | data_masked[5373];
  assign N7770 = N7769 | data_masked[5501];
  assign N7769 = N7768 | data_masked[5629];
  assign N7768 = N7767 | data_masked[5757];
  assign N7767 = N7766 | data_masked[5885];
  assign N7766 = N7765 | data_masked[6013];
  assign N7765 = N7764 | data_masked[6141];
  assign N7764 = N7763 | data_masked[6269];
  assign N7763 = N7762 | data_masked[6397];
  assign N7762 = N7761 | data_masked[6525];
  assign N7761 = N7760 | data_masked[6653];
  assign N7760 = N7759 | data_masked[6781];
  assign N7759 = N7758 | data_masked[6909];
  assign N7758 = N7757 | data_masked[7037];
  assign N7757 = N7756 | data_masked[7165];
  assign N7756 = N7755 | data_masked[7293];
  assign N7755 = N7754 | data_masked[7421];
  assign N7754 = N7753 | data_masked[7549];
  assign N7753 = N7752 | data_masked[7677];
  assign N7752 = N7751 | data_masked[7805];
  assign N7751 = N7750 | data_masked[7933];
  assign N7750 = data_masked[8189] | data_masked[8061];
  assign data_o[126] = N7873 | data_masked[126];
  assign N7873 = N7872 | data_masked[254];
  assign N7872 = N7871 | data_masked[382];
  assign N7871 = N7870 | data_masked[510];
  assign N7870 = N7869 | data_masked[638];
  assign N7869 = N7868 | data_masked[766];
  assign N7868 = N7867 | data_masked[894];
  assign N7867 = N7866 | data_masked[1022];
  assign N7866 = N7865 | data_masked[1150];
  assign N7865 = N7864 | data_masked[1278];
  assign N7864 = N7863 | data_masked[1406];
  assign N7863 = N7862 | data_masked[1534];
  assign N7862 = N7861 | data_masked[1662];
  assign N7861 = N7860 | data_masked[1790];
  assign N7860 = N7859 | data_masked[1918];
  assign N7859 = N7858 | data_masked[2046];
  assign N7858 = N7857 | data_masked[2174];
  assign N7857 = N7856 | data_masked[2302];
  assign N7856 = N7855 | data_masked[2430];
  assign N7855 = N7854 | data_masked[2558];
  assign N7854 = N7853 | data_masked[2686];
  assign N7853 = N7852 | data_masked[2814];
  assign N7852 = N7851 | data_masked[2942];
  assign N7851 = N7850 | data_masked[3070];
  assign N7850 = N7849 | data_masked[3198];
  assign N7849 = N7848 | data_masked[3326];
  assign N7848 = N7847 | data_masked[3454];
  assign N7847 = N7846 | data_masked[3582];
  assign N7846 = N7845 | data_masked[3710];
  assign N7845 = N7844 | data_masked[3838];
  assign N7844 = N7843 | data_masked[3966];
  assign N7843 = N7842 | data_masked[4094];
  assign N7842 = N7841 | data_masked[4222];
  assign N7841 = N7840 | data_masked[4350];
  assign N7840 = N7839 | data_masked[4478];
  assign N7839 = N7838 | data_masked[4606];
  assign N7838 = N7837 | data_masked[4734];
  assign N7837 = N7836 | data_masked[4862];
  assign N7836 = N7835 | data_masked[4990];
  assign N7835 = N7834 | data_masked[5118];
  assign N7834 = N7833 | data_masked[5246];
  assign N7833 = N7832 | data_masked[5374];
  assign N7832 = N7831 | data_masked[5502];
  assign N7831 = N7830 | data_masked[5630];
  assign N7830 = N7829 | data_masked[5758];
  assign N7829 = N7828 | data_masked[5886];
  assign N7828 = N7827 | data_masked[6014];
  assign N7827 = N7826 | data_masked[6142];
  assign N7826 = N7825 | data_masked[6270];
  assign N7825 = N7824 | data_masked[6398];
  assign N7824 = N7823 | data_masked[6526];
  assign N7823 = N7822 | data_masked[6654];
  assign N7822 = N7821 | data_masked[6782];
  assign N7821 = N7820 | data_masked[6910];
  assign N7820 = N7819 | data_masked[7038];
  assign N7819 = N7818 | data_masked[7166];
  assign N7818 = N7817 | data_masked[7294];
  assign N7817 = N7816 | data_masked[7422];
  assign N7816 = N7815 | data_masked[7550];
  assign N7815 = N7814 | data_masked[7678];
  assign N7814 = N7813 | data_masked[7806];
  assign N7813 = N7812 | data_masked[7934];
  assign N7812 = data_masked[8190] | data_masked[8062];
  assign data_o[127] = N7935 | data_masked[127];
  assign N7935 = N7934 | data_masked[255];
  assign N7934 = N7933 | data_masked[383];
  assign N7933 = N7932 | data_masked[511];
  assign N7932 = N7931 | data_masked[639];
  assign N7931 = N7930 | data_masked[767];
  assign N7930 = N7929 | data_masked[895];
  assign N7929 = N7928 | data_masked[1023];
  assign N7928 = N7927 | data_masked[1151];
  assign N7927 = N7926 | data_masked[1279];
  assign N7926 = N7925 | data_masked[1407];
  assign N7925 = N7924 | data_masked[1535];
  assign N7924 = N7923 | data_masked[1663];
  assign N7923 = N7922 | data_masked[1791];
  assign N7922 = N7921 | data_masked[1919];
  assign N7921 = N7920 | data_masked[2047];
  assign N7920 = N7919 | data_masked[2175];
  assign N7919 = N7918 | data_masked[2303];
  assign N7918 = N7917 | data_masked[2431];
  assign N7917 = N7916 | data_masked[2559];
  assign N7916 = N7915 | data_masked[2687];
  assign N7915 = N7914 | data_masked[2815];
  assign N7914 = N7913 | data_masked[2943];
  assign N7913 = N7912 | data_masked[3071];
  assign N7912 = N7911 | data_masked[3199];
  assign N7911 = N7910 | data_masked[3327];
  assign N7910 = N7909 | data_masked[3455];
  assign N7909 = N7908 | data_masked[3583];
  assign N7908 = N7907 | data_masked[3711];
  assign N7907 = N7906 | data_masked[3839];
  assign N7906 = N7905 | data_masked[3967];
  assign N7905 = N7904 | data_masked[4095];
  assign N7904 = N7903 | data_masked[4223];
  assign N7903 = N7902 | data_masked[4351];
  assign N7902 = N7901 | data_masked[4479];
  assign N7901 = N7900 | data_masked[4607];
  assign N7900 = N7899 | data_masked[4735];
  assign N7899 = N7898 | data_masked[4863];
  assign N7898 = N7897 | data_masked[4991];
  assign N7897 = N7896 | data_masked[5119];
  assign N7896 = N7895 | data_masked[5247];
  assign N7895 = N7894 | data_masked[5375];
  assign N7894 = N7893 | data_masked[5503];
  assign N7893 = N7892 | data_masked[5631];
  assign N7892 = N7891 | data_masked[5759];
  assign N7891 = N7890 | data_masked[5887];
  assign N7890 = N7889 | data_masked[6015];
  assign N7889 = N7888 | data_masked[6143];
  assign N7888 = N7887 | data_masked[6271];
  assign N7887 = N7886 | data_masked[6399];
  assign N7886 = N7885 | data_masked[6527];
  assign N7885 = N7884 | data_masked[6655];
  assign N7884 = N7883 | data_masked[6783];
  assign N7883 = N7882 | data_masked[6911];
  assign N7882 = N7881 | data_masked[7039];
  assign N7881 = N7880 | data_masked[7167];
  assign N7880 = N7879 | data_masked[7295];
  assign N7879 = N7878 | data_masked[7423];
  assign N7878 = N7877 | data_masked[7551];
  assign N7877 = N7876 | data_masked[7679];
  assign N7876 = N7875 | data_masked[7807];
  assign N7875 = N7874 | data_masked[7935];
  assign N7874 = data_masked[8191] | data_masked[8063];

endmodule

