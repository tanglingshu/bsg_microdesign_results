

module top
(
  clk_i,
  reset_i,
  v_i,
  tag_i,
  data_i,
  yumi_o,
  v_o,
  yumi_i,
  data_o
);

  input [7:0] tag_i;
  input [7:0] data_i;
  output [255:0] v_o;
  input [255:0] yumi_i;
  output [2047:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  output yumi_o;

  bsg_1_to_n_tagged_fifo
  wrapper
  (
    .tag_i(tag_i),
    .data_i(data_i),
    .v_o(v_o),
    .yumi_i(yumi_i),
    .data_o(data_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .yumi_o(yumi_o)
  );


endmodule



module bsg_decode_num_out_p256
(
  i,
  o
);

  input [7:0] i;
  output [255:0] o;
  wire [255:0] o;
  assign o = { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1 } << i;

endmodule



module bsg_decode_with_v_num_out_p256
(
  i,
  v_i,
  o
);

  input [7:0] i;
  output [255:0] o;
  input v_i;
  wire [255:0] o,lo;

  bsg_decode_num_out_p256
  bd
  (
    .i(i),
    .o(lo)
  );

  assign o[255] = v_i & lo[255];
  assign o[254] = v_i & lo[254];
  assign o[253] = v_i & lo[253];
  assign o[252] = v_i & lo[252];
  assign o[251] = v_i & lo[251];
  assign o[250] = v_i & lo[250];
  assign o[249] = v_i & lo[249];
  assign o[248] = v_i & lo[248];
  assign o[247] = v_i & lo[247];
  assign o[246] = v_i & lo[246];
  assign o[245] = v_i & lo[245];
  assign o[244] = v_i & lo[244];
  assign o[243] = v_i & lo[243];
  assign o[242] = v_i & lo[242];
  assign o[241] = v_i & lo[241];
  assign o[240] = v_i & lo[240];
  assign o[239] = v_i & lo[239];
  assign o[238] = v_i & lo[238];
  assign o[237] = v_i & lo[237];
  assign o[236] = v_i & lo[236];
  assign o[235] = v_i & lo[235];
  assign o[234] = v_i & lo[234];
  assign o[233] = v_i & lo[233];
  assign o[232] = v_i & lo[232];
  assign o[231] = v_i & lo[231];
  assign o[230] = v_i & lo[230];
  assign o[229] = v_i & lo[229];
  assign o[228] = v_i & lo[228];
  assign o[227] = v_i & lo[227];
  assign o[226] = v_i & lo[226];
  assign o[225] = v_i & lo[225];
  assign o[224] = v_i & lo[224];
  assign o[223] = v_i & lo[223];
  assign o[222] = v_i & lo[222];
  assign o[221] = v_i & lo[221];
  assign o[220] = v_i & lo[220];
  assign o[219] = v_i & lo[219];
  assign o[218] = v_i & lo[218];
  assign o[217] = v_i & lo[217];
  assign o[216] = v_i & lo[216];
  assign o[215] = v_i & lo[215];
  assign o[214] = v_i & lo[214];
  assign o[213] = v_i & lo[213];
  assign o[212] = v_i & lo[212];
  assign o[211] = v_i & lo[211];
  assign o[210] = v_i & lo[210];
  assign o[209] = v_i & lo[209];
  assign o[208] = v_i & lo[208];
  assign o[207] = v_i & lo[207];
  assign o[206] = v_i & lo[206];
  assign o[205] = v_i & lo[205];
  assign o[204] = v_i & lo[204];
  assign o[203] = v_i & lo[203];
  assign o[202] = v_i & lo[202];
  assign o[201] = v_i & lo[201];
  assign o[200] = v_i & lo[200];
  assign o[199] = v_i & lo[199];
  assign o[198] = v_i & lo[198];
  assign o[197] = v_i & lo[197];
  assign o[196] = v_i & lo[196];
  assign o[195] = v_i & lo[195];
  assign o[194] = v_i & lo[194];
  assign o[193] = v_i & lo[193];
  assign o[192] = v_i & lo[192];
  assign o[191] = v_i & lo[191];
  assign o[190] = v_i & lo[190];
  assign o[189] = v_i & lo[189];
  assign o[188] = v_i & lo[188];
  assign o[187] = v_i & lo[187];
  assign o[186] = v_i & lo[186];
  assign o[185] = v_i & lo[185];
  assign o[184] = v_i & lo[184];
  assign o[183] = v_i & lo[183];
  assign o[182] = v_i & lo[182];
  assign o[181] = v_i & lo[181];
  assign o[180] = v_i & lo[180];
  assign o[179] = v_i & lo[179];
  assign o[178] = v_i & lo[178];
  assign o[177] = v_i & lo[177];
  assign o[176] = v_i & lo[176];
  assign o[175] = v_i & lo[175];
  assign o[174] = v_i & lo[174];
  assign o[173] = v_i & lo[173];
  assign o[172] = v_i & lo[172];
  assign o[171] = v_i & lo[171];
  assign o[170] = v_i & lo[170];
  assign o[169] = v_i & lo[169];
  assign o[168] = v_i & lo[168];
  assign o[167] = v_i & lo[167];
  assign o[166] = v_i & lo[166];
  assign o[165] = v_i & lo[165];
  assign o[164] = v_i & lo[164];
  assign o[163] = v_i & lo[163];
  assign o[162] = v_i & lo[162];
  assign o[161] = v_i & lo[161];
  assign o[160] = v_i & lo[160];
  assign o[159] = v_i & lo[159];
  assign o[158] = v_i & lo[158];
  assign o[157] = v_i & lo[157];
  assign o[156] = v_i & lo[156];
  assign o[155] = v_i & lo[155];
  assign o[154] = v_i & lo[154];
  assign o[153] = v_i & lo[153];
  assign o[152] = v_i & lo[152];
  assign o[151] = v_i & lo[151];
  assign o[150] = v_i & lo[150];
  assign o[149] = v_i & lo[149];
  assign o[148] = v_i & lo[148];
  assign o[147] = v_i & lo[147];
  assign o[146] = v_i & lo[146];
  assign o[145] = v_i & lo[145];
  assign o[144] = v_i & lo[144];
  assign o[143] = v_i & lo[143];
  assign o[142] = v_i & lo[142];
  assign o[141] = v_i & lo[141];
  assign o[140] = v_i & lo[140];
  assign o[139] = v_i & lo[139];
  assign o[138] = v_i & lo[138];
  assign o[137] = v_i & lo[137];
  assign o[136] = v_i & lo[136];
  assign o[135] = v_i & lo[135];
  assign o[134] = v_i & lo[134];
  assign o[133] = v_i & lo[133];
  assign o[132] = v_i & lo[132];
  assign o[131] = v_i & lo[131];
  assign o[130] = v_i & lo[130];
  assign o[129] = v_i & lo[129];
  assign o[128] = v_i & lo[128];
  assign o[127] = v_i & lo[127];
  assign o[126] = v_i & lo[126];
  assign o[125] = v_i & lo[125];
  assign o[124] = v_i & lo[124];
  assign o[123] = v_i & lo[123];
  assign o[122] = v_i & lo[122];
  assign o[121] = v_i & lo[121];
  assign o[120] = v_i & lo[120];
  assign o[119] = v_i & lo[119];
  assign o[118] = v_i & lo[118];
  assign o[117] = v_i & lo[117];
  assign o[116] = v_i & lo[116];
  assign o[115] = v_i & lo[115];
  assign o[114] = v_i & lo[114];
  assign o[113] = v_i & lo[113];
  assign o[112] = v_i & lo[112];
  assign o[111] = v_i & lo[111];
  assign o[110] = v_i & lo[110];
  assign o[109] = v_i & lo[109];
  assign o[108] = v_i & lo[108];
  assign o[107] = v_i & lo[107];
  assign o[106] = v_i & lo[106];
  assign o[105] = v_i & lo[105];
  assign o[104] = v_i & lo[104];
  assign o[103] = v_i & lo[103];
  assign o[102] = v_i & lo[102];
  assign o[101] = v_i & lo[101];
  assign o[100] = v_i & lo[100];
  assign o[99] = v_i & lo[99];
  assign o[98] = v_i & lo[98];
  assign o[97] = v_i & lo[97];
  assign o[96] = v_i & lo[96];
  assign o[95] = v_i & lo[95];
  assign o[94] = v_i & lo[94];
  assign o[93] = v_i & lo[93];
  assign o[92] = v_i & lo[92];
  assign o[91] = v_i & lo[91];
  assign o[90] = v_i & lo[90];
  assign o[89] = v_i & lo[89];
  assign o[88] = v_i & lo[88];
  assign o[87] = v_i & lo[87];
  assign o[86] = v_i & lo[86];
  assign o[85] = v_i & lo[85];
  assign o[84] = v_i & lo[84];
  assign o[83] = v_i & lo[83];
  assign o[82] = v_i & lo[82];
  assign o[81] = v_i & lo[81];
  assign o[80] = v_i & lo[80];
  assign o[79] = v_i & lo[79];
  assign o[78] = v_i & lo[78];
  assign o[77] = v_i & lo[77];
  assign o[76] = v_i & lo[76];
  assign o[75] = v_i & lo[75];
  assign o[74] = v_i & lo[74];
  assign o[73] = v_i & lo[73];
  assign o[72] = v_i & lo[72];
  assign o[71] = v_i & lo[71];
  assign o[70] = v_i & lo[70];
  assign o[69] = v_i & lo[69];
  assign o[68] = v_i & lo[68];
  assign o[67] = v_i & lo[67];
  assign o[66] = v_i & lo[66];
  assign o[65] = v_i & lo[65];
  assign o[64] = v_i & lo[64];
  assign o[63] = v_i & lo[63];
  assign o[62] = v_i & lo[62];
  assign o[61] = v_i & lo[61];
  assign o[60] = v_i & lo[60];
  assign o[59] = v_i & lo[59];
  assign o[58] = v_i & lo[58];
  assign o[57] = v_i & lo[57];
  assign o[56] = v_i & lo[56];
  assign o[55] = v_i & lo[55];
  assign o[54] = v_i & lo[54];
  assign o[53] = v_i & lo[53];
  assign o[52] = v_i & lo[52];
  assign o[51] = v_i & lo[51];
  assign o[50] = v_i & lo[50];
  assign o[49] = v_i & lo[49];
  assign o[48] = v_i & lo[48];
  assign o[47] = v_i & lo[47];
  assign o[46] = v_i & lo[46];
  assign o[45] = v_i & lo[45];
  assign o[44] = v_i & lo[44];
  assign o[43] = v_i & lo[43];
  assign o[42] = v_i & lo[42];
  assign o[41] = v_i & lo[41];
  assign o[40] = v_i & lo[40];
  assign o[39] = v_i & lo[39];
  assign o[38] = v_i & lo[38];
  assign o[37] = v_i & lo[37];
  assign o[36] = v_i & lo[36];
  assign o[35] = v_i & lo[35];
  assign o[34] = v_i & lo[34];
  assign o[33] = v_i & lo[33];
  assign o[32] = v_i & lo[32];
  assign o[31] = v_i & lo[31];
  assign o[30] = v_i & lo[30];
  assign o[29] = v_i & lo[29];
  assign o[28] = v_i & lo[28];
  assign o[27] = v_i & lo[27];
  assign o[26] = v_i & lo[26];
  assign o[25] = v_i & lo[25];
  assign o[24] = v_i & lo[24];
  assign o[23] = v_i & lo[23];
  assign o[22] = v_i & lo[22];
  assign o[21] = v_i & lo[21];
  assign o[20] = v_i & lo[20];
  assign o[19] = v_i & lo[19];
  assign o[18] = v_i & lo[18];
  assign o[17] = v_i & lo[17];
  assign o[16] = v_i & lo[16];
  assign o[15] = v_i & lo[15];
  assign o[14] = v_i & lo[14];
  assign o[13] = v_i & lo[13];
  assign o[12] = v_i & lo[12];
  assign o[11] = v_i & lo[11];
  assign o[10] = v_i & lo[10];
  assign o[9] = v_i & lo[9];
  assign o[8] = v_i & lo[8];
  assign o[7] = v_i & lo[7];
  assign o[6] = v_i & lo[6];
  assign o[5] = v_i & lo[5];
  assign o[4] = v_i & lo[4];
  assign o[3] = v_i & lo[3];
  assign o[2] = v_i & lo[2];
  assign o[1] = v_i & lo[1];
  assign o[0] = v_i & lo[0];

endmodule



module bsg_1_to_n_tagged_num_out_p256
(
  clk_i,
  reset_i,
  v_i,
  tag_i,
  yumi_o,
  v_o,
  ready_i
);

  input [7:0] tag_i;
  output [255:0] v_o;
  input [255:0] ready_i;
  input clk_i;
  input reset_i;
  input v_i;
  output yumi_o;
  wire [255:0] v_o;
  wire yumi_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,
  N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,
  N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,
  N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,
  N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,
  N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,
  N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,
  N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,
  N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,
  N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,
  N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,
  N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,
  N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,
  N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,
  N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
  N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,
  N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,
  N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,
  N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,
  N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,
  N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,
  N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,
  N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,
  N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,
  N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,
  N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,
  N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,
  N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,
  N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,
  N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,
  N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,
  N516;

  bsg_decode_with_v_num_out_p256
  many_bdv
  (
    .i(tag_i),
    .v_i(v_i),
    .o(v_o)
  );

  assign N516 = (N260)? ready_i[0] : 
                (N262)? ready_i[1] : 
                (N264)? ready_i[2] : 
                (N266)? ready_i[3] : 
                (N268)? ready_i[4] : 
                (N270)? ready_i[5] : 
                (N272)? ready_i[6] : 
                (N274)? ready_i[7] : 
                (N276)? ready_i[8] : 
                (N278)? ready_i[9] : 
                (N280)? ready_i[10] : 
                (N282)? ready_i[11] : 
                (N284)? ready_i[12] : 
                (N286)? ready_i[13] : 
                (N288)? ready_i[14] : 
                (N290)? ready_i[15] : 
                (N292)? ready_i[16] : 
                (N294)? ready_i[17] : 
                (N296)? ready_i[18] : 
                (N298)? ready_i[19] : 
                (N300)? ready_i[20] : 
                (N302)? ready_i[21] : 
                (N304)? ready_i[22] : 
                (N306)? ready_i[23] : 
                (N308)? ready_i[24] : 
                (N310)? ready_i[25] : 
                (N312)? ready_i[26] : 
                (N314)? ready_i[27] : 
                (N316)? ready_i[28] : 
                (N318)? ready_i[29] : 
                (N320)? ready_i[30] : 
                (N322)? ready_i[31] : 
                (N324)? ready_i[32] : 
                (N326)? ready_i[33] : 
                (N328)? ready_i[34] : 
                (N330)? ready_i[35] : 
                (N332)? ready_i[36] : 
                (N334)? ready_i[37] : 
                (N336)? ready_i[38] : 
                (N338)? ready_i[39] : 
                (N340)? ready_i[40] : 
                (N342)? ready_i[41] : 
                (N344)? ready_i[42] : 
                (N346)? ready_i[43] : 
                (N348)? ready_i[44] : 
                (N350)? ready_i[45] : 
                (N352)? ready_i[46] : 
                (N354)? ready_i[47] : 
                (N356)? ready_i[48] : 
                (N358)? ready_i[49] : 
                (N360)? ready_i[50] : 
                (N362)? ready_i[51] : 
                (N364)? ready_i[52] : 
                (N366)? ready_i[53] : 
                (N368)? ready_i[54] : 
                (N370)? ready_i[55] : 
                (N372)? ready_i[56] : 
                (N374)? ready_i[57] : 
                (N376)? ready_i[58] : 
                (N378)? ready_i[59] : 
                (N380)? ready_i[60] : 
                (N382)? ready_i[61] : 
                (N384)? ready_i[62] : 
                (N386)? ready_i[63] : 
                (N388)? ready_i[64] : 
                (N390)? ready_i[65] : 
                (N392)? ready_i[66] : 
                (N394)? ready_i[67] : 
                (N396)? ready_i[68] : 
                (N398)? ready_i[69] : 
                (N400)? ready_i[70] : 
                (N402)? ready_i[71] : 
                (N404)? ready_i[72] : 
                (N406)? ready_i[73] : 
                (N408)? ready_i[74] : 
                (N410)? ready_i[75] : 
                (N412)? ready_i[76] : 
                (N414)? ready_i[77] : 
                (N416)? ready_i[78] : 
                (N418)? ready_i[79] : 
                (N420)? ready_i[80] : 
                (N422)? ready_i[81] : 
                (N424)? ready_i[82] : 
                (N426)? ready_i[83] : 
                (N428)? ready_i[84] : 
                (N430)? ready_i[85] : 
                (N432)? ready_i[86] : 
                (N434)? ready_i[87] : 
                (N436)? ready_i[88] : 
                (N438)? ready_i[89] : 
                (N440)? ready_i[90] : 
                (N442)? ready_i[91] : 
                (N444)? ready_i[92] : 
                (N446)? ready_i[93] : 
                (N448)? ready_i[94] : 
                (N450)? ready_i[95] : 
                (N452)? ready_i[96] : 
                (N454)? ready_i[97] : 
                (N456)? ready_i[98] : 
                (N458)? ready_i[99] : 
                (N460)? ready_i[100] : 
                (N462)? ready_i[101] : 
                (N464)? ready_i[102] : 
                (N466)? ready_i[103] : 
                (N468)? ready_i[104] : 
                (N470)? ready_i[105] : 
                (N472)? ready_i[106] : 
                (N474)? ready_i[107] : 
                (N476)? ready_i[108] : 
                (N478)? ready_i[109] : 
                (N480)? ready_i[110] : 
                (N482)? ready_i[111] : 
                (N484)? ready_i[112] : 
                (N486)? ready_i[113] : 
                (N488)? ready_i[114] : 
                (N490)? ready_i[115] : 
                (N492)? ready_i[116] : 
                (N494)? ready_i[117] : 
                (N496)? ready_i[118] : 
                (N498)? ready_i[119] : 
                (N500)? ready_i[120] : 
                (N502)? ready_i[121] : 
                (N504)? ready_i[122] : 
                (N506)? ready_i[123] : 
                (N508)? ready_i[124] : 
                (N510)? ready_i[125] : 
                (N512)? ready_i[126] : 
                (N514)? ready_i[127] : 
                (N261)? ready_i[128] : 
                (N263)? ready_i[129] : 
                (N265)? ready_i[130] : 
                (N267)? ready_i[131] : 
                (N269)? ready_i[132] : 
                (N271)? ready_i[133] : 
                (N273)? ready_i[134] : 
                (N275)? ready_i[135] : 
                (N277)? ready_i[136] : 
                (N279)? ready_i[137] : 
                (N281)? ready_i[138] : 
                (N283)? ready_i[139] : 
                (N285)? ready_i[140] : 
                (N287)? ready_i[141] : 
                (N289)? ready_i[142] : 
                (N291)? ready_i[143] : 
                (N293)? ready_i[144] : 
                (N295)? ready_i[145] : 
                (N297)? ready_i[146] : 
                (N299)? ready_i[147] : 
                (N301)? ready_i[148] : 
                (N303)? ready_i[149] : 
                (N305)? ready_i[150] : 
                (N307)? ready_i[151] : 
                (N309)? ready_i[152] : 
                (N311)? ready_i[153] : 
                (N313)? ready_i[154] : 
                (N315)? ready_i[155] : 
                (N317)? ready_i[156] : 
                (N319)? ready_i[157] : 
                (N321)? ready_i[158] : 
                (N323)? ready_i[159] : 
                (N325)? ready_i[160] : 
                (N327)? ready_i[161] : 
                (N329)? ready_i[162] : 
                (N331)? ready_i[163] : 
                (N333)? ready_i[164] : 
                (N335)? ready_i[165] : 
                (N337)? ready_i[166] : 
                (N339)? ready_i[167] : 
                (N341)? ready_i[168] : 
                (N343)? ready_i[169] : 
                (N345)? ready_i[170] : 
                (N347)? ready_i[171] : 
                (N349)? ready_i[172] : 
                (N351)? ready_i[173] : 
                (N353)? ready_i[174] : 
                (N355)? ready_i[175] : 
                (N357)? ready_i[176] : 
                (N359)? ready_i[177] : 
                (N361)? ready_i[178] : 
                (N363)? ready_i[179] : 
                (N365)? ready_i[180] : 
                (N367)? ready_i[181] : 
                (N369)? ready_i[182] : 
                (N371)? ready_i[183] : 
                (N373)? ready_i[184] : 
                (N375)? ready_i[185] : 
                (N377)? ready_i[186] : 
                (N379)? ready_i[187] : 
                (N381)? ready_i[188] : 
                (N383)? ready_i[189] : 
                (N385)? ready_i[190] : 
                (N387)? ready_i[191] : 
                (N389)? ready_i[192] : 
                (N391)? ready_i[193] : 
                (N393)? ready_i[194] : 
                (N395)? ready_i[195] : 
                (N397)? ready_i[196] : 
                (N399)? ready_i[197] : 
                (N401)? ready_i[198] : 
                (N403)? ready_i[199] : 
                (N405)? ready_i[200] : 
                (N407)? ready_i[201] : 
                (N409)? ready_i[202] : 
                (N411)? ready_i[203] : 
                (N413)? ready_i[204] : 
                (N415)? ready_i[205] : 
                (N417)? ready_i[206] : 
                (N419)? ready_i[207] : 
                (N421)? ready_i[208] : 
                (N423)? ready_i[209] : 
                (N425)? ready_i[210] : 
                (N427)? ready_i[211] : 
                (N429)? ready_i[212] : 
                (N431)? ready_i[213] : 
                (N433)? ready_i[214] : 
                (N435)? ready_i[215] : 
                (N437)? ready_i[216] : 
                (N439)? ready_i[217] : 
                (N441)? ready_i[218] : 
                (N443)? ready_i[219] : 
                (N445)? ready_i[220] : 
                (N447)? ready_i[221] : 
                (N449)? ready_i[222] : 
                (N451)? ready_i[223] : 
                (N453)? ready_i[224] : 
                (N455)? ready_i[225] : 
                (N457)? ready_i[226] : 
                (N459)? ready_i[227] : 
                (N461)? ready_i[228] : 
                (N463)? ready_i[229] : 
                (N465)? ready_i[230] : 
                (N467)? ready_i[231] : 
                (N469)? ready_i[232] : 
                (N471)? ready_i[233] : 
                (N473)? ready_i[234] : 
                (N475)? ready_i[235] : 
                (N477)? ready_i[236] : 
                (N479)? ready_i[237] : 
                (N481)? ready_i[238] : 
                (N483)? ready_i[239] : 
                (N485)? ready_i[240] : 
                (N487)? ready_i[241] : 
                (N489)? ready_i[242] : 
                (N491)? ready_i[243] : 
                (N493)? ready_i[244] : 
                (N495)? ready_i[245] : 
                (N497)? ready_i[246] : 
                (N499)? ready_i[247] : 
                (N501)? ready_i[248] : 
                (N503)? ready_i[249] : 
                (N505)? ready_i[250] : 
                (N507)? ready_i[251] : 
                (N509)? ready_i[252] : 
                (N511)? ready_i[253] : 
                (N513)? ready_i[254] : 
                (N515)? ready_i[255] : 1'b0;
  assign N0 = ~tag_i[0];
  assign N1 = ~tag_i[1];
  assign N2 = N0 & N1;
  assign N3 = N0 & tag_i[1];
  assign N4 = tag_i[0] & N1;
  assign N5 = tag_i[0] & tag_i[1];
  assign N6 = ~tag_i[2];
  assign N7 = N2 & N6;
  assign N8 = N2 & tag_i[2];
  assign N9 = N4 & N6;
  assign N10 = N4 & tag_i[2];
  assign N11 = N3 & N6;
  assign N12 = N3 & tag_i[2];
  assign N13 = N5 & N6;
  assign N14 = N5 & tag_i[2];
  assign N15 = ~tag_i[3];
  assign N16 = N7 & N15;
  assign N17 = N7 & tag_i[3];
  assign N18 = N9 & N15;
  assign N19 = N9 & tag_i[3];
  assign N20 = N11 & N15;
  assign N21 = N11 & tag_i[3];
  assign N22 = N13 & N15;
  assign N23 = N13 & tag_i[3];
  assign N24 = N8 & N15;
  assign N25 = N8 & tag_i[3];
  assign N26 = N10 & N15;
  assign N27 = N10 & tag_i[3];
  assign N28 = N12 & N15;
  assign N29 = N12 & tag_i[3];
  assign N30 = N14 & N15;
  assign N31 = N14 & tag_i[3];
  assign N32 = ~tag_i[4];
  assign N33 = N16 & N32;
  assign N34 = N16 & tag_i[4];
  assign N35 = N18 & N32;
  assign N36 = N18 & tag_i[4];
  assign N37 = N20 & N32;
  assign N38 = N20 & tag_i[4];
  assign N39 = N22 & N32;
  assign N40 = N22 & tag_i[4];
  assign N41 = N24 & N32;
  assign N42 = N24 & tag_i[4];
  assign N43 = N26 & N32;
  assign N44 = N26 & tag_i[4];
  assign N45 = N28 & N32;
  assign N46 = N28 & tag_i[4];
  assign N47 = N30 & N32;
  assign N48 = N30 & tag_i[4];
  assign N49 = N17 & N32;
  assign N50 = N17 & tag_i[4];
  assign N51 = N19 & N32;
  assign N52 = N19 & tag_i[4];
  assign N53 = N21 & N32;
  assign N54 = N21 & tag_i[4];
  assign N55 = N23 & N32;
  assign N56 = N23 & tag_i[4];
  assign N57 = N25 & N32;
  assign N58 = N25 & tag_i[4];
  assign N59 = N27 & N32;
  assign N60 = N27 & tag_i[4];
  assign N61 = N29 & N32;
  assign N62 = N29 & tag_i[4];
  assign N63 = N31 & N32;
  assign N64 = N31 & tag_i[4];
  assign N65 = ~tag_i[5];
  assign N66 = N33 & N65;
  assign N67 = N33 & tag_i[5];
  assign N68 = N35 & N65;
  assign N69 = N35 & tag_i[5];
  assign N70 = N37 & N65;
  assign N71 = N37 & tag_i[5];
  assign N72 = N39 & N65;
  assign N73 = N39 & tag_i[5];
  assign N74 = N41 & N65;
  assign N75 = N41 & tag_i[5];
  assign N76 = N43 & N65;
  assign N77 = N43 & tag_i[5];
  assign N78 = N45 & N65;
  assign N79 = N45 & tag_i[5];
  assign N80 = N47 & N65;
  assign N81 = N47 & tag_i[5];
  assign N82 = N49 & N65;
  assign N83 = N49 & tag_i[5];
  assign N84 = N51 & N65;
  assign N85 = N51 & tag_i[5];
  assign N86 = N53 & N65;
  assign N87 = N53 & tag_i[5];
  assign N88 = N55 & N65;
  assign N89 = N55 & tag_i[5];
  assign N90 = N57 & N65;
  assign N91 = N57 & tag_i[5];
  assign N92 = N59 & N65;
  assign N93 = N59 & tag_i[5];
  assign N94 = N61 & N65;
  assign N95 = N61 & tag_i[5];
  assign N96 = N63 & N65;
  assign N97 = N63 & tag_i[5];
  assign N98 = N34 & N65;
  assign N99 = N34 & tag_i[5];
  assign N100 = N36 & N65;
  assign N101 = N36 & tag_i[5];
  assign N102 = N38 & N65;
  assign N103 = N38 & tag_i[5];
  assign N104 = N40 & N65;
  assign N105 = N40 & tag_i[5];
  assign N106 = N42 & N65;
  assign N107 = N42 & tag_i[5];
  assign N108 = N44 & N65;
  assign N109 = N44 & tag_i[5];
  assign N110 = N46 & N65;
  assign N111 = N46 & tag_i[5];
  assign N112 = N48 & N65;
  assign N113 = N48 & tag_i[5];
  assign N114 = N50 & N65;
  assign N115 = N50 & tag_i[5];
  assign N116 = N52 & N65;
  assign N117 = N52 & tag_i[5];
  assign N118 = N54 & N65;
  assign N119 = N54 & tag_i[5];
  assign N120 = N56 & N65;
  assign N121 = N56 & tag_i[5];
  assign N122 = N58 & N65;
  assign N123 = N58 & tag_i[5];
  assign N124 = N60 & N65;
  assign N125 = N60 & tag_i[5];
  assign N126 = N62 & N65;
  assign N127 = N62 & tag_i[5];
  assign N128 = N64 & N65;
  assign N129 = N64 & tag_i[5];
  assign N130 = ~tag_i[6];
  assign N131 = N66 & N130;
  assign N132 = N66 & tag_i[6];
  assign N133 = N68 & N130;
  assign N134 = N68 & tag_i[6];
  assign N135 = N70 & N130;
  assign N136 = N70 & tag_i[6];
  assign N137 = N72 & N130;
  assign N138 = N72 & tag_i[6];
  assign N139 = N74 & N130;
  assign N140 = N74 & tag_i[6];
  assign N141 = N76 & N130;
  assign N142 = N76 & tag_i[6];
  assign N143 = N78 & N130;
  assign N144 = N78 & tag_i[6];
  assign N145 = N80 & N130;
  assign N146 = N80 & tag_i[6];
  assign N147 = N82 & N130;
  assign N148 = N82 & tag_i[6];
  assign N149 = N84 & N130;
  assign N150 = N84 & tag_i[6];
  assign N151 = N86 & N130;
  assign N152 = N86 & tag_i[6];
  assign N153 = N88 & N130;
  assign N154 = N88 & tag_i[6];
  assign N155 = N90 & N130;
  assign N156 = N90 & tag_i[6];
  assign N157 = N92 & N130;
  assign N158 = N92 & tag_i[6];
  assign N159 = N94 & N130;
  assign N160 = N94 & tag_i[6];
  assign N161 = N96 & N130;
  assign N162 = N96 & tag_i[6];
  assign N163 = N98 & N130;
  assign N164 = N98 & tag_i[6];
  assign N165 = N100 & N130;
  assign N166 = N100 & tag_i[6];
  assign N167 = N102 & N130;
  assign N168 = N102 & tag_i[6];
  assign N169 = N104 & N130;
  assign N170 = N104 & tag_i[6];
  assign N171 = N106 & N130;
  assign N172 = N106 & tag_i[6];
  assign N173 = N108 & N130;
  assign N174 = N108 & tag_i[6];
  assign N175 = N110 & N130;
  assign N176 = N110 & tag_i[6];
  assign N177 = N112 & N130;
  assign N178 = N112 & tag_i[6];
  assign N179 = N114 & N130;
  assign N180 = N114 & tag_i[6];
  assign N181 = N116 & N130;
  assign N182 = N116 & tag_i[6];
  assign N183 = N118 & N130;
  assign N184 = N118 & tag_i[6];
  assign N185 = N120 & N130;
  assign N186 = N120 & tag_i[6];
  assign N187 = N122 & N130;
  assign N188 = N122 & tag_i[6];
  assign N189 = N124 & N130;
  assign N190 = N124 & tag_i[6];
  assign N191 = N126 & N130;
  assign N192 = N126 & tag_i[6];
  assign N193 = N128 & N130;
  assign N194 = N128 & tag_i[6];
  assign N195 = N67 & N130;
  assign N196 = N67 & tag_i[6];
  assign N197 = N69 & N130;
  assign N198 = N69 & tag_i[6];
  assign N199 = N71 & N130;
  assign N200 = N71 & tag_i[6];
  assign N201 = N73 & N130;
  assign N202 = N73 & tag_i[6];
  assign N203 = N75 & N130;
  assign N204 = N75 & tag_i[6];
  assign N205 = N77 & N130;
  assign N206 = N77 & tag_i[6];
  assign N207 = N79 & N130;
  assign N208 = N79 & tag_i[6];
  assign N209 = N81 & N130;
  assign N210 = N81 & tag_i[6];
  assign N211 = N83 & N130;
  assign N212 = N83 & tag_i[6];
  assign N213 = N85 & N130;
  assign N214 = N85 & tag_i[6];
  assign N215 = N87 & N130;
  assign N216 = N87 & tag_i[6];
  assign N217 = N89 & N130;
  assign N218 = N89 & tag_i[6];
  assign N219 = N91 & N130;
  assign N220 = N91 & tag_i[6];
  assign N221 = N93 & N130;
  assign N222 = N93 & tag_i[6];
  assign N223 = N95 & N130;
  assign N224 = N95 & tag_i[6];
  assign N225 = N97 & N130;
  assign N226 = N97 & tag_i[6];
  assign N227 = N99 & N130;
  assign N228 = N99 & tag_i[6];
  assign N229 = N101 & N130;
  assign N230 = N101 & tag_i[6];
  assign N231 = N103 & N130;
  assign N232 = N103 & tag_i[6];
  assign N233 = N105 & N130;
  assign N234 = N105 & tag_i[6];
  assign N235 = N107 & N130;
  assign N236 = N107 & tag_i[6];
  assign N237 = N109 & N130;
  assign N238 = N109 & tag_i[6];
  assign N239 = N111 & N130;
  assign N240 = N111 & tag_i[6];
  assign N241 = N113 & N130;
  assign N242 = N113 & tag_i[6];
  assign N243 = N115 & N130;
  assign N244 = N115 & tag_i[6];
  assign N245 = N117 & N130;
  assign N246 = N117 & tag_i[6];
  assign N247 = N119 & N130;
  assign N248 = N119 & tag_i[6];
  assign N249 = N121 & N130;
  assign N250 = N121 & tag_i[6];
  assign N251 = N123 & N130;
  assign N252 = N123 & tag_i[6];
  assign N253 = N125 & N130;
  assign N254 = N125 & tag_i[6];
  assign N255 = N127 & N130;
  assign N256 = N127 & tag_i[6];
  assign N257 = N129 & N130;
  assign N258 = N129 & tag_i[6];
  assign N259 = ~tag_i[7];
  assign N260 = N131 & N259;
  assign N261 = N131 & tag_i[7];
  assign N262 = N133 & N259;
  assign N263 = N133 & tag_i[7];
  assign N264 = N135 & N259;
  assign N265 = N135 & tag_i[7];
  assign N266 = N137 & N259;
  assign N267 = N137 & tag_i[7];
  assign N268 = N139 & N259;
  assign N269 = N139 & tag_i[7];
  assign N270 = N141 & N259;
  assign N271 = N141 & tag_i[7];
  assign N272 = N143 & N259;
  assign N273 = N143 & tag_i[7];
  assign N274 = N145 & N259;
  assign N275 = N145 & tag_i[7];
  assign N276 = N147 & N259;
  assign N277 = N147 & tag_i[7];
  assign N278 = N149 & N259;
  assign N279 = N149 & tag_i[7];
  assign N280 = N151 & N259;
  assign N281 = N151 & tag_i[7];
  assign N282 = N153 & N259;
  assign N283 = N153 & tag_i[7];
  assign N284 = N155 & N259;
  assign N285 = N155 & tag_i[7];
  assign N286 = N157 & N259;
  assign N287 = N157 & tag_i[7];
  assign N288 = N159 & N259;
  assign N289 = N159 & tag_i[7];
  assign N290 = N161 & N259;
  assign N291 = N161 & tag_i[7];
  assign N292 = N163 & N259;
  assign N293 = N163 & tag_i[7];
  assign N294 = N165 & N259;
  assign N295 = N165 & tag_i[7];
  assign N296 = N167 & N259;
  assign N297 = N167 & tag_i[7];
  assign N298 = N169 & N259;
  assign N299 = N169 & tag_i[7];
  assign N300 = N171 & N259;
  assign N301 = N171 & tag_i[7];
  assign N302 = N173 & N259;
  assign N303 = N173 & tag_i[7];
  assign N304 = N175 & N259;
  assign N305 = N175 & tag_i[7];
  assign N306 = N177 & N259;
  assign N307 = N177 & tag_i[7];
  assign N308 = N179 & N259;
  assign N309 = N179 & tag_i[7];
  assign N310 = N181 & N259;
  assign N311 = N181 & tag_i[7];
  assign N312 = N183 & N259;
  assign N313 = N183 & tag_i[7];
  assign N314 = N185 & N259;
  assign N315 = N185 & tag_i[7];
  assign N316 = N187 & N259;
  assign N317 = N187 & tag_i[7];
  assign N318 = N189 & N259;
  assign N319 = N189 & tag_i[7];
  assign N320 = N191 & N259;
  assign N321 = N191 & tag_i[7];
  assign N322 = N193 & N259;
  assign N323 = N193 & tag_i[7];
  assign N324 = N195 & N259;
  assign N325 = N195 & tag_i[7];
  assign N326 = N197 & N259;
  assign N327 = N197 & tag_i[7];
  assign N328 = N199 & N259;
  assign N329 = N199 & tag_i[7];
  assign N330 = N201 & N259;
  assign N331 = N201 & tag_i[7];
  assign N332 = N203 & N259;
  assign N333 = N203 & tag_i[7];
  assign N334 = N205 & N259;
  assign N335 = N205 & tag_i[7];
  assign N336 = N207 & N259;
  assign N337 = N207 & tag_i[7];
  assign N338 = N209 & N259;
  assign N339 = N209 & tag_i[7];
  assign N340 = N211 & N259;
  assign N341 = N211 & tag_i[7];
  assign N342 = N213 & N259;
  assign N343 = N213 & tag_i[7];
  assign N344 = N215 & N259;
  assign N345 = N215 & tag_i[7];
  assign N346 = N217 & N259;
  assign N347 = N217 & tag_i[7];
  assign N348 = N219 & N259;
  assign N349 = N219 & tag_i[7];
  assign N350 = N221 & N259;
  assign N351 = N221 & tag_i[7];
  assign N352 = N223 & N259;
  assign N353 = N223 & tag_i[7];
  assign N354 = N225 & N259;
  assign N355 = N225 & tag_i[7];
  assign N356 = N227 & N259;
  assign N357 = N227 & tag_i[7];
  assign N358 = N229 & N259;
  assign N359 = N229 & tag_i[7];
  assign N360 = N231 & N259;
  assign N361 = N231 & tag_i[7];
  assign N362 = N233 & N259;
  assign N363 = N233 & tag_i[7];
  assign N364 = N235 & N259;
  assign N365 = N235 & tag_i[7];
  assign N366 = N237 & N259;
  assign N367 = N237 & tag_i[7];
  assign N368 = N239 & N259;
  assign N369 = N239 & tag_i[7];
  assign N370 = N241 & N259;
  assign N371 = N241 & tag_i[7];
  assign N372 = N243 & N259;
  assign N373 = N243 & tag_i[7];
  assign N374 = N245 & N259;
  assign N375 = N245 & tag_i[7];
  assign N376 = N247 & N259;
  assign N377 = N247 & tag_i[7];
  assign N378 = N249 & N259;
  assign N379 = N249 & tag_i[7];
  assign N380 = N251 & N259;
  assign N381 = N251 & tag_i[7];
  assign N382 = N253 & N259;
  assign N383 = N253 & tag_i[7];
  assign N384 = N255 & N259;
  assign N385 = N255 & tag_i[7];
  assign N386 = N257 & N259;
  assign N387 = N257 & tag_i[7];
  assign N388 = N132 & N259;
  assign N389 = N132 & tag_i[7];
  assign N390 = N134 & N259;
  assign N391 = N134 & tag_i[7];
  assign N392 = N136 & N259;
  assign N393 = N136 & tag_i[7];
  assign N394 = N138 & N259;
  assign N395 = N138 & tag_i[7];
  assign N396 = N140 & N259;
  assign N397 = N140 & tag_i[7];
  assign N398 = N142 & N259;
  assign N399 = N142 & tag_i[7];
  assign N400 = N144 & N259;
  assign N401 = N144 & tag_i[7];
  assign N402 = N146 & N259;
  assign N403 = N146 & tag_i[7];
  assign N404 = N148 & N259;
  assign N405 = N148 & tag_i[7];
  assign N406 = N150 & N259;
  assign N407 = N150 & tag_i[7];
  assign N408 = N152 & N259;
  assign N409 = N152 & tag_i[7];
  assign N410 = N154 & N259;
  assign N411 = N154 & tag_i[7];
  assign N412 = N156 & N259;
  assign N413 = N156 & tag_i[7];
  assign N414 = N158 & N259;
  assign N415 = N158 & tag_i[7];
  assign N416 = N160 & N259;
  assign N417 = N160 & tag_i[7];
  assign N418 = N162 & N259;
  assign N419 = N162 & tag_i[7];
  assign N420 = N164 & N259;
  assign N421 = N164 & tag_i[7];
  assign N422 = N166 & N259;
  assign N423 = N166 & tag_i[7];
  assign N424 = N168 & N259;
  assign N425 = N168 & tag_i[7];
  assign N426 = N170 & N259;
  assign N427 = N170 & tag_i[7];
  assign N428 = N172 & N259;
  assign N429 = N172 & tag_i[7];
  assign N430 = N174 & N259;
  assign N431 = N174 & tag_i[7];
  assign N432 = N176 & N259;
  assign N433 = N176 & tag_i[7];
  assign N434 = N178 & N259;
  assign N435 = N178 & tag_i[7];
  assign N436 = N180 & N259;
  assign N437 = N180 & tag_i[7];
  assign N438 = N182 & N259;
  assign N439 = N182 & tag_i[7];
  assign N440 = N184 & N259;
  assign N441 = N184 & tag_i[7];
  assign N442 = N186 & N259;
  assign N443 = N186 & tag_i[7];
  assign N444 = N188 & N259;
  assign N445 = N188 & tag_i[7];
  assign N446 = N190 & N259;
  assign N447 = N190 & tag_i[7];
  assign N448 = N192 & N259;
  assign N449 = N192 & tag_i[7];
  assign N450 = N194 & N259;
  assign N451 = N194 & tag_i[7];
  assign N452 = N196 & N259;
  assign N453 = N196 & tag_i[7];
  assign N454 = N198 & N259;
  assign N455 = N198 & tag_i[7];
  assign N456 = N200 & N259;
  assign N457 = N200 & tag_i[7];
  assign N458 = N202 & N259;
  assign N459 = N202 & tag_i[7];
  assign N460 = N204 & N259;
  assign N461 = N204 & tag_i[7];
  assign N462 = N206 & N259;
  assign N463 = N206 & tag_i[7];
  assign N464 = N208 & N259;
  assign N465 = N208 & tag_i[7];
  assign N466 = N210 & N259;
  assign N467 = N210 & tag_i[7];
  assign N468 = N212 & N259;
  assign N469 = N212 & tag_i[7];
  assign N470 = N214 & N259;
  assign N471 = N214 & tag_i[7];
  assign N472 = N216 & N259;
  assign N473 = N216 & tag_i[7];
  assign N474 = N218 & N259;
  assign N475 = N218 & tag_i[7];
  assign N476 = N220 & N259;
  assign N477 = N220 & tag_i[7];
  assign N478 = N222 & N259;
  assign N479 = N222 & tag_i[7];
  assign N480 = N224 & N259;
  assign N481 = N224 & tag_i[7];
  assign N482 = N226 & N259;
  assign N483 = N226 & tag_i[7];
  assign N484 = N228 & N259;
  assign N485 = N228 & tag_i[7];
  assign N486 = N230 & N259;
  assign N487 = N230 & tag_i[7];
  assign N488 = N232 & N259;
  assign N489 = N232 & tag_i[7];
  assign N490 = N234 & N259;
  assign N491 = N234 & tag_i[7];
  assign N492 = N236 & N259;
  assign N493 = N236 & tag_i[7];
  assign N494 = N238 & N259;
  assign N495 = N238 & tag_i[7];
  assign N496 = N240 & N259;
  assign N497 = N240 & tag_i[7];
  assign N498 = N242 & N259;
  assign N499 = N242 & tag_i[7];
  assign N500 = N244 & N259;
  assign N501 = N244 & tag_i[7];
  assign N502 = N246 & N259;
  assign N503 = N246 & tag_i[7];
  assign N504 = N248 & N259;
  assign N505 = N248 & tag_i[7];
  assign N506 = N250 & N259;
  assign N507 = N250 & tag_i[7];
  assign N508 = N252 & N259;
  assign N509 = N252 & tag_i[7];
  assign N510 = N254 & N259;
  assign N511 = N254 & tag_i[7];
  assign N512 = N256 & N259;
  assign N513 = N256 & tag_i[7];
  assign N514 = N258 & N259;
  assign N515 = N258 & tag_i[7];
  assign yumi_o = N516 & v_i;

endmodule



module bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
(
  clk_i,
  reset_i,
  data_i,
  v_i,
  ready_o,
  v_o,
  data_o,
  yumi_i
);

  input [7:0] data_i;
  output [7:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  input yumi_i;
  output ready_o;
  output v_o;
  wire [7:0] data_o,little_data,big_data_lo;
  wire ready_o,v_o,N0,N1,N2,N3,little_ready_lo,little_will_have_space,N4,N5,big_deq,N6,
  big_full_lo,big_empty_lo,N7,N8,little_valid,big_enq,N9,N10,N11,N12,N13,
  big_valid,N14,N15,N16,N17,N18,N19,N20,N21,N22,N23;
  reg big_deq_r;

  bsg_fifo_1rw_large
  big1p
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(big_valid),
    .enq_not_deq_i(big_enq),
    .full_o(big_full_lo),
    .empty_o(big_empty_lo),
    .data_o(big_data_lo)
  );


  bsg_two_fifo
  little2p
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .ready_o(little_ready_lo),
    .data_i(little_data),
    .v_i(little_valid),
    .v_o(v_o),
    .data_o(data_o),
    .yumi_i(yumi_i)
  );

  assign N6 = (N0)? 1'b0 : 
              (N1)? big_deq : 1'b0;
  assign N0 = N5;
  assign N1 = N4;
  assign little_valid = (N2)? 1'b1 : 
                        (N15)? N10 : 
                        (N8)? 1'b0 : 1'b0;
  assign N2 = big_deq_r;
  assign big_enq = (N2)? v_i : 
                   (N15)? N11 : 
                   (N8)? N12 : 1'b0;
  assign big_deq = (N2)? N9 : 
                   (N15)? 1'b0 : 
                   (N8)? N13 : 1'b0;
  assign little_data = (N2)? big_data_lo : 
                       (N3)? data_i : 1'b0;
  assign N3 = N16;
  assign little_will_have_space = little_ready_lo | yumi_i;
  assign N4 = ~reset_i;
  assign N5 = reset_i;
  assign ready_o = ~big_full_lo;
  assign N7 = big_empty_lo | big_deq_r;
  assign N8 = ~N7;
  assign N9 = N19 & N20;
  assign N19 = N17 & N18;
  assign N17 = ~big_empty_lo;
  assign N18 = ~v_i;
  assign N20 = ~v_o;
  assign N10 = v_i & little_will_have_space;
  assign N11 = v_i & N21;
  assign N21 = ~little_will_have_space;
  assign N12 = v_i & N22;
  assign N22 = ~big_full_lo;
  assign N13 = N23 & little_will_have_space;
  assign N23 = ~N12;
  assign big_valid = big_enq | big_deq;
  assign N14 = ~big_deq_r;
  assign N15 = big_empty_lo & N14;
  assign N16 = ~big_deq_r;

  always @(posedge clk_i) begin
    if(1'b1) begin
      big_deq_r <= N6;
    end 
  end


endmodule



module bsg_1_to_n_tagged_fifo
(
  clk_i,
  reset_i,
  v_i,
  tag_i,
  data_i,
  yumi_o,
  v_o,
  yumi_i,
  data_o
);

  input [7:0] tag_i;
  input [7:0] data_i;
  output [255:0] v_o;
  input [255:0] yumi_i;
  output [2047:0] data_o;
  input clk_i;
  input reset_i;
  input v_i;
  output yumi_o;
  wire [255:0] v_o,valid_lo,ready_li;
  wire [2047:0] data_o;
  wire yumi_o;

  bsg_1_to_n_tagged_num_out_p256
  u_1_to_n
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .v_i(v_i),
    .tag_i(tag_i),
    .yumi_o(yumi_o),
    .v_o(valid_lo),
    .ready_i(ready_li)
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_0__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[0]),
    .ready_o(ready_li[0]),
    .v_o(v_o[0]),
    .data_o(data_o[7:0]),
    .yumi_i(yumi_i[0])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_1__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[1]),
    .ready_o(ready_li[1]),
    .v_o(v_o[1]),
    .data_o(data_o[15:8]),
    .yumi_i(yumi_i[1])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_2__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[2]),
    .ready_o(ready_li[2]),
    .v_o(v_o[2]),
    .data_o(data_o[23:16]),
    .yumi_i(yumi_i[2])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_3__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[3]),
    .ready_o(ready_li[3]),
    .v_o(v_o[3]),
    .data_o(data_o[31:24]),
    .yumi_i(yumi_i[3])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_4__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[4]),
    .ready_o(ready_li[4]),
    .v_o(v_o[4]),
    .data_o(data_o[39:32]),
    .yumi_i(yumi_i[4])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_5__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[5]),
    .ready_o(ready_li[5]),
    .v_o(v_o[5]),
    .data_o(data_o[47:40]),
    .yumi_i(yumi_i[5])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_6__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[6]),
    .ready_o(ready_li[6]),
    .v_o(v_o[6]),
    .data_o(data_o[55:48]),
    .yumi_i(yumi_i[6])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_7__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[7]),
    .ready_o(ready_li[7]),
    .v_o(v_o[7]),
    .data_o(data_o[63:56]),
    .yumi_i(yumi_i[7])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_8__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[8]),
    .ready_o(ready_li[8]),
    .v_o(v_o[8]),
    .data_o(data_o[71:64]),
    .yumi_i(yumi_i[8])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_9__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[9]),
    .ready_o(ready_li[9]),
    .v_o(v_o[9]),
    .data_o(data_o[79:72]),
    .yumi_i(yumi_i[9])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_10__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[10]),
    .ready_o(ready_li[10]),
    .v_o(v_o[10]),
    .data_o(data_o[87:80]),
    .yumi_i(yumi_i[10])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_11__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[11]),
    .ready_o(ready_li[11]),
    .v_o(v_o[11]),
    .data_o(data_o[95:88]),
    .yumi_i(yumi_i[11])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_12__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[12]),
    .ready_o(ready_li[12]),
    .v_o(v_o[12]),
    .data_o(data_o[103:96]),
    .yumi_i(yumi_i[12])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_13__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[13]),
    .ready_o(ready_li[13]),
    .v_o(v_o[13]),
    .data_o(data_o[111:104]),
    .yumi_i(yumi_i[13])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_14__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[14]),
    .ready_o(ready_li[14]),
    .v_o(v_o[14]),
    .data_o(data_o[119:112]),
    .yumi_i(yumi_i[14])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_15__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[15]),
    .ready_o(ready_li[15]),
    .v_o(v_o[15]),
    .data_o(data_o[127:120]),
    .yumi_i(yumi_i[15])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_16__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[16]),
    .ready_o(ready_li[16]),
    .v_o(v_o[16]),
    .data_o(data_o[135:128]),
    .yumi_i(yumi_i[16])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_17__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[17]),
    .ready_o(ready_li[17]),
    .v_o(v_o[17]),
    .data_o(data_o[143:136]),
    .yumi_i(yumi_i[17])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_18__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[18]),
    .ready_o(ready_li[18]),
    .v_o(v_o[18]),
    .data_o(data_o[151:144]),
    .yumi_i(yumi_i[18])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_19__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[19]),
    .ready_o(ready_li[19]),
    .v_o(v_o[19]),
    .data_o(data_o[159:152]),
    .yumi_i(yumi_i[19])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_20__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[20]),
    .ready_o(ready_li[20]),
    .v_o(v_o[20]),
    .data_o(data_o[167:160]),
    .yumi_i(yumi_i[20])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_21__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[21]),
    .ready_o(ready_li[21]),
    .v_o(v_o[21]),
    .data_o(data_o[175:168]),
    .yumi_i(yumi_i[21])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_22__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[22]),
    .ready_o(ready_li[22]),
    .v_o(v_o[22]),
    .data_o(data_o[183:176]),
    .yumi_i(yumi_i[22])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_23__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[23]),
    .ready_o(ready_li[23]),
    .v_o(v_o[23]),
    .data_o(data_o[191:184]),
    .yumi_i(yumi_i[23])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_24__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[24]),
    .ready_o(ready_li[24]),
    .v_o(v_o[24]),
    .data_o(data_o[199:192]),
    .yumi_i(yumi_i[24])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_25__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[25]),
    .ready_o(ready_li[25]),
    .v_o(v_o[25]),
    .data_o(data_o[207:200]),
    .yumi_i(yumi_i[25])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_26__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[26]),
    .ready_o(ready_li[26]),
    .v_o(v_o[26]),
    .data_o(data_o[215:208]),
    .yumi_i(yumi_i[26])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_27__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[27]),
    .ready_o(ready_li[27]),
    .v_o(v_o[27]),
    .data_o(data_o[223:216]),
    .yumi_i(yumi_i[27])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_28__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[28]),
    .ready_o(ready_li[28]),
    .v_o(v_o[28]),
    .data_o(data_o[231:224]),
    .yumi_i(yumi_i[28])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_29__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[29]),
    .ready_o(ready_li[29]),
    .v_o(v_o[29]),
    .data_o(data_o[239:232]),
    .yumi_i(yumi_i[29])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_30__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[30]),
    .ready_o(ready_li[30]),
    .v_o(v_o[30]),
    .data_o(data_o[247:240]),
    .yumi_i(yumi_i[30])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_31__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[31]),
    .ready_o(ready_li[31]),
    .v_o(v_o[31]),
    .data_o(data_o[255:248]),
    .yumi_i(yumi_i[31])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_32__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[32]),
    .ready_o(ready_li[32]),
    .v_o(v_o[32]),
    .data_o(data_o[263:256]),
    .yumi_i(yumi_i[32])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_33__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[33]),
    .ready_o(ready_li[33]),
    .v_o(v_o[33]),
    .data_o(data_o[271:264]),
    .yumi_i(yumi_i[33])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_34__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[34]),
    .ready_o(ready_li[34]),
    .v_o(v_o[34]),
    .data_o(data_o[279:272]),
    .yumi_i(yumi_i[34])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_35__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[35]),
    .ready_o(ready_li[35]),
    .v_o(v_o[35]),
    .data_o(data_o[287:280]),
    .yumi_i(yumi_i[35])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_36__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[36]),
    .ready_o(ready_li[36]),
    .v_o(v_o[36]),
    .data_o(data_o[295:288]),
    .yumi_i(yumi_i[36])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_37__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[37]),
    .ready_o(ready_li[37]),
    .v_o(v_o[37]),
    .data_o(data_o[303:296]),
    .yumi_i(yumi_i[37])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_38__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[38]),
    .ready_o(ready_li[38]),
    .v_o(v_o[38]),
    .data_o(data_o[311:304]),
    .yumi_i(yumi_i[38])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_39__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[39]),
    .ready_o(ready_li[39]),
    .v_o(v_o[39]),
    .data_o(data_o[319:312]),
    .yumi_i(yumi_i[39])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_40__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[40]),
    .ready_o(ready_li[40]),
    .v_o(v_o[40]),
    .data_o(data_o[327:320]),
    .yumi_i(yumi_i[40])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_41__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[41]),
    .ready_o(ready_li[41]),
    .v_o(v_o[41]),
    .data_o(data_o[335:328]),
    .yumi_i(yumi_i[41])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_42__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[42]),
    .ready_o(ready_li[42]),
    .v_o(v_o[42]),
    .data_o(data_o[343:336]),
    .yumi_i(yumi_i[42])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_43__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[43]),
    .ready_o(ready_li[43]),
    .v_o(v_o[43]),
    .data_o(data_o[351:344]),
    .yumi_i(yumi_i[43])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_44__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[44]),
    .ready_o(ready_li[44]),
    .v_o(v_o[44]),
    .data_o(data_o[359:352]),
    .yumi_i(yumi_i[44])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_45__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[45]),
    .ready_o(ready_li[45]),
    .v_o(v_o[45]),
    .data_o(data_o[367:360]),
    .yumi_i(yumi_i[45])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_46__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[46]),
    .ready_o(ready_li[46]),
    .v_o(v_o[46]),
    .data_o(data_o[375:368]),
    .yumi_i(yumi_i[46])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_47__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[47]),
    .ready_o(ready_li[47]),
    .v_o(v_o[47]),
    .data_o(data_o[383:376]),
    .yumi_i(yumi_i[47])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_48__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[48]),
    .ready_o(ready_li[48]),
    .v_o(v_o[48]),
    .data_o(data_o[391:384]),
    .yumi_i(yumi_i[48])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_49__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[49]),
    .ready_o(ready_li[49]),
    .v_o(v_o[49]),
    .data_o(data_o[399:392]),
    .yumi_i(yumi_i[49])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_50__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[50]),
    .ready_o(ready_li[50]),
    .v_o(v_o[50]),
    .data_o(data_o[407:400]),
    .yumi_i(yumi_i[50])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_51__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[51]),
    .ready_o(ready_li[51]),
    .v_o(v_o[51]),
    .data_o(data_o[415:408]),
    .yumi_i(yumi_i[51])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_52__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[52]),
    .ready_o(ready_li[52]),
    .v_o(v_o[52]),
    .data_o(data_o[423:416]),
    .yumi_i(yumi_i[52])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_53__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[53]),
    .ready_o(ready_li[53]),
    .v_o(v_o[53]),
    .data_o(data_o[431:424]),
    .yumi_i(yumi_i[53])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_54__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[54]),
    .ready_o(ready_li[54]),
    .v_o(v_o[54]),
    .data_o(data_o[439:432]),
    .yumi_i(yumi_i[54])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_55__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[55]),
    .ready_o(ready_li[55]),
    .v_o(v_o[55]),
    .data_o(data_o[447:440]),
    .yumi_i(yumi_i[55])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_56__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[56]),
    .ready_o(ready_li[56]),
    .v_o(v_o[56]),
    .data_o(data_o[455:448]),
    .yumi_i(yumi_i[56])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_57__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[57]),
    .ready_o(ready_li[57]),
    .v_o(v_o[57]),
    .data_o(data_o[463:456]),
    .yumi_i(yumi_i[57])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_58__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[58]),
    .ready_o(ready_li[58]),
    .v_o(v_o[58]),
    .data_o(data_o[471:464]),
    .yumi_i(yumi_i[58])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_59__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[59]),
    .ready_o(ready_li[59]),
    .v_o(v_o[59]),
    .data_o(data_o[479:472]),
    .yumi_i(yumi_i[59])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_60__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[60]),
    .ready_o(ready_li[60]),
    .v_o(v_o[60]),
    .data_o(data_o[487:480]),
    .yumi_i(yumi_i[60])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_61__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[61]),
    .ready_o(ready_li[61]),
    .v_o(v_o[61]),
    .data_o(data_o[495:488]),
    .yumi_i(yumi_i[61])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_62__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[62]),
    .ready_o(ready_li[62]),
    .v_o(v_o[62]),
    .data_o(data_o[503:496]),
    .yumi_i(yumi_i[62])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_63__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[63]),
    .ready_o(ready_li[63]),
    .v_o(v_o[63]),
    .data_o(data_o[511:504]),
    .yumi_i(yumi_i[63])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_64__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[64]),
    .ready_o(ready_li[64]),
    .v_o(v_o[64]),
    .data_o(data_o[519:512]),
    .yumi_i(yumi_i[64])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_65__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[65]),
    .ready_o(ready_li[65]),
    .v_o(v_o[65]),
    .data_o(data_o[527:520]),
    .yumi_i(yumi_i[65])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_66__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[66]),
    .ready_o(ready_li[66]),
    .v_o(v_o[66]),
    .data_o(data_o[535:528]),
    .yumi_i(yumi_i[66])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_67__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[67]),
    .ready_o(ready_li[67]),
    .v_o(v_o[67]),
    .data_o(data_o[543:536]),
    .yumi_i(yumi_i[67])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_68__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[68]),
    .ready_o(ready_li[68]),
    .v_o(v_o[68]),
    .data_o(data_o[551:544]),
    .yumi_i(yumi_i[68])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_69__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[69]),
    .ready_o(ready_li[69]),
    .v_o(v_o[69]),
    .data_o(data_o[559:552]),
    .yumi_i(yumi_i[69])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_70__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[70]),
    .ready_o(ready_li[70]),
    .v_o(v_o[70]),
    .data_o(data_o[567:560]),
    .yumi_i(yumi_i[70])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_71__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[71]),
    .ready_o(ready_li[71]),
    .v_o(v_o[71]),
    .data_o(data_o[575:568]),
    .yumi_i(yumi_i[71])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_72__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[72]),
    .ready_o(ready_li[72]),
    .v_o(v_o[72]),
    .data_o(data_o[583:576]),
    .yumi_i(yumi_i[72])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_73__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[73]),
    .ready_o(ready_li[73]),
    .v_o(v_o[73]),
    .data_o(data_o[591:584]),
    .yumi_i(yumi_i[73])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_74__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[74]),
    .ready_o(ready_li[74]),
    .v_o(v_o[74]),
    .data_o(data_o[599:592]),
    .yumi_i(yumi_i[74])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_75__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[75]),
    .ready_o(ready_li[75]),
    .v_o(v_o[75]),
    .data_o(data_o[607:600]),
    .yumi_i(yumi_i[75])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_76__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[76]),
    .ready_o(ready_li[76]),
    .v_o(v_o[76]),
    .data_o(data_o[615:608]),
    .yumi_i(yumi_i[76])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_77__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[77]),
    .ready_o(ready_li[77]),
    .v_o(v_o[77]),
    .data_o(data_o[623:616]),
    .yumi_i(yumi_i[77])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_78__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[78]),
    .ready_o(ready_li[78]),
    .v_o(v_o[78]),
    .data_o(data_o[631:624]),
    .yumi_i(yumi_i[78])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_79__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[79]),
    .ready_o(ready_li[79]),
    .v_o(v_o[79]),
    .data_o(data_o[639:632]),
    .yumi_i(yumi_i[79])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_80__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[80]),
    .ready_o(ready_li[80]),
    .v_o(v_o[80]),
    .data_o(data_o[647:640]),
    .yumi_i(yumi_i[80])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_81__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[81]),
    .ready_o(ready_li[81]),
    .v_o(v_o[81]),
    .data_o(data_o[655:648]),
    .yumi_i(yumi_i[81])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_82__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[82]),
    .ready_o(ready_li[82]),
    .v_o(v_o[82]),
    .data_o(data_o[663:656]),
    .yumi_i(yumi_i[82])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_83__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[83]),
    .ready_o(ready_li[83]),
    .v_o(v_o[83]),
    .data_o(data_o[671:664]),
    .yumi_i(yumi_i[83])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_84__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[84]),
    .ready_o(ready_li[84]),
    .v_o(v_o[84]),
    .data_o(data_o[679:672]),
    .yumi_i(yumi_i[84])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_85__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[85]),
    .ready_o(ready_li[85]),
    .v_o(v_o[85]),
    .data_o(data_o[687:680]),
    .yumi_i(yumi_i[85])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_86__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[86]),
    .ready_o(ready_li[86]),
    .v_o(v_o[86]),
    .data_o(data_o[695:688]),
    .yumi_i(yumi_i[86])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_87__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[87]),
    .ready_o(ready_li[87]),
    .v_o(v_o[87]),
    .data_o(data_o[703:696]),
    .yumi_i(yumi_i[87])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_88__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[88]),
    .ready_o(ready_li[88]),
    .v_o(v_o[88]),
    .data_o(data_o[711:704]),
    .yumi_i(yumi_i[88])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_89__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[89]),
    .ready_o(ready_li[89]),
    .v_o(v_o[89]),
    .data_o(data_o[719:712]),
    .yumi_i(yumi_i[89])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_90__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[90]),
    .ready_o(ready_li[90]),
    .v_o(v_o[90]),
    .data_o(data_o[727:720]),
    .yumi_i(yumi_i[90])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_91__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[91]),
    .ready_o(ready_li[91]),
    .v_o(v_o[91]),
    .data_o(data_o[735:728]),
    .yumi_i(yumi_i[91])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_92__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[92]),
    .ready_o(ready_li[92]),
    .v_o(v_o[92]),
    .data_o(data_o[743:736]),
    .yumi_i(yumi_i[92])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_93__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[93]),
    .ready_o(ready_li[93]),
    .v_o(v_o[93]),
    .data_o(data_o[751:744]),
    .yumi_i(yumi_i[93])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_94__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[94]),
    .ready_o(ready_li[94]),
    .v_o(v_o[94]),
    .data_o(data_o[759:752]),
    .yumi_i(yumi_i[94])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_95__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[95]),
    .ready_o(ready_li[95]),
    .v_o(v_o[95]),
    .data_o(data_o[767:760]),
    .yumi_i(yumi_i[95])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_96__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[96]),
    .ready_o(ready_li[96]),
    .v_o(v_o[96]),
    .data_o(data_o[775:768]),
    .yumi_i(yumi_i[96])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_97__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[97]),
    .ready_o(ready_li[97]),
    .v_o(v_o[97]),
    .data_o(data_o[783:776]),
    .yumi_i(yumi_i[97])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_98__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[98]),
    .ready_o(ready_li[98]),
    .v_o(v_o[98]),
    .data_o(data_o[791:784]),
    .yumi_i(yumi_i[98])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_99__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[99]),
    .ready_o(ready_li[99]),
    .v_o(v_o[99]),
    .data_o(data_o[799:792]),
    .yumi_i(yumi_i[99])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_100__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[100]),
    .ready_o(ready_li[100]),
    .v_o(v_o[100]),
    .data_o(data_o[807:800]),
    .yumi_i(yumi_i[100])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_101__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[101]),
    .ready_o(ready_li[101]),
    .v_o(v_o[101]),
    .data_o(data_o[815:808]),
    .yumi_i(yumi_i[101])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_102__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[102]),
    .ready_o(ready_li[102]),
    .v_o(v_o[102]),
    .data_o(data_o[823:816]),
    .yumi_i(yumi_i[102])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_103__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[103]),
    .ready_o(ready_li[103]),
    .v_o(v_o[103]),
    .data_o(data_o[831:824]),
    .yumi_i(yumi_i[103])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_104__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[104]),
    .ready_o(ready_li[104]),
    .v_o(v_o[104]),
    .data_o(data_o[839:832]),
    .yumi_i(yumi_i[104])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_105__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[105]),
    .ready_o(ready_li[105]),
    .v_o(v_o[105]),
    .data_o(data_o[847:840]),
    .yumi_i(yumi_i[105])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_106__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[106]),
    .ready_o(ready_li[106]),
    .v_o(v_o[106]),
    .data_o(data_o[855:848]),
    .yumi_i(yumi_i[106])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_107__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[107]),
    .ready_o(ready_li[107]),
    .v_o(v_o[107]),
    .data_o(data_o[863:856]),
    .yumi_i(yumi_i[107])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_108__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[108]),
    .ready_o(ready_li[108]),
    .v_o(v_o[108]),
    .data_o(data_o[871:864]),
    .yumi_i(yumi_i[108])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_109__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[109]),
    .ready_o(ready_li[109]),
    .v_o(v_o[109]),
    .data_o(data_o[879:872]),
    .yumi_i(yumi_i[109])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_110__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[110]),
    .ready_o(ready_li[110]),
    .v_o(v_o[110]),
    .data_o(data_o[887:880]),
    .yumi_i(yumi_i[110])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_111__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[111]),
    .ready_o(ready_li[111]),
    .v_o(v_o[111]),
    .data_o(data_o[895:888]),
    .yumi_i(yumi_i[111])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_112__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[112]),
    .ready_o(ready_li[112]),
    .v_o(v_o[112]),
    .data_o(data_o[903:896]),
    .yumi_i(yumi_i[112])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_113__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[113]),
    .ready_o(ready_li[113]),
    .v_o(v_o[113]),
    .data_o(data_o[911:904]),
    .yumi_i(yumi_i[113])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_114__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[114]),
    .ready_o(ready_li[114]),
    .v_o(v_o[114]),
    .data_o(data_o[919:912]),
    .yumi_i(yumi_i[114])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_115__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[115]),
    .ready_o(ready_li[115]),
    .v_o(v_o[115]),
    .data_o(data_o[927:920]),
    .yumi_i(yumi_i[115])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_116__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[116]),
    .ready_o(ready_li[116]),
    .v_o(v_o[116]),
    .data_o(data_o[935:928]),
    .yumi_i(yumi_i[116])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_117__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[117]),
    .ready_o(ready_li[117]),
    .v_o(v_o[117]),
    .data_o(data_o[943:936]),
    .yumi_i(yumi_i[117])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_118__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[118]),
    .ready_o(ready_li[118]),
    .v_o(v_o[118]),
    .data_o(data_o[951:944]),
    .yumi_i(yumi_i[118])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_119__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[119]),
    .ready_o(ready_li[119]),
    .v_o(v_o[119]),
    .data_o(data_o[959:952]),
    .yumi_i(yumi_i[119])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_120__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[120]),
    .ready_o(ready_li[120]),
    .v_o(v_o[120]),
    .data_o(data_o[967:960]),
    .yumi_i(yumi_i[120])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_121__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[121]),
    .ready_o(ready_li[121]),
    .v_o(v_o[121]),
    .data_o(data_o[975:968]),
    .yumi_i(yumi_i[121])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_122__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[122]),
    .ready_o(ready_li[122]),
    .v_o(v_o[122]),
    .data_o(data_o[983:976]),
    .yumi_i(yumi_i[122])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_123__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[123]),
    .ready_o(ready_li[123]),
    .v_o(v_o[123]),
    .data_o(data_o[991:984]),
    .yumi_i(yumi_i[123])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_124__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[124]),
    .ready_o(ready_li[124]),
    .v_o(v_o[124]),
    .data_o(data_o[999:992]),
    .yumi_i(yumi_i[124])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_125__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[125]),
    .ready_o(ready_li[125]),
    .v_o(v_o[125]),
    .data_o(data_o[1007:1000]),
    .yumi_i(yumi_i[125])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_126__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[126]),
    .ready_o(ready_li[126]),
    .v_o(v_o[126]),
    .data_o(data_o[1015:1008]),
    .yumi_i(yumi_i[126])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_127__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[127]),
    .ready_o(ready_li[127]),
    .v_o(v_o[127]),
    .data_o(data_o[1023:1016]),
    .yumi_i(yumi_i[127])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_128__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[128]),
    .ready_o(ready_li[128]),
    .v_o(v_o[128]),
    .data_o(data_o[1031:1024]),
    .yumi_i(yumi_i[128])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_129__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[129]),
    .ready_o(ready_li[129]),
    .v_o(v_o[129]),
    .data_o(data_o[1039:1032]),
    .yumi_i(yumi_i[129])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_130__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[130]),
    .ready_o(ready_li[130]),
    .v_o(v_o[130]),
    .data_o(data_o[1047:1040]),
    .yumi_i(yumi_i[130])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_131__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[131]),
    .ready_o(ready_li[131]),
    .v_o(v_o[131]),
    .data_o(data_o[1055:1048]),
    .yumi_i(yumi_i[131])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_132__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[132]),
    .ready_o(ready_li[132]),
    .v_o(v_o[132]),
    .data_o(data_o[1063:1056]),
    .yumi_i(yumi_i[132])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_133__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[133]),
    .ready_o(ready_li[133]),
    .v_o(v_o[133]),
    .data_o(data_o[1071:1064]),
    .yumi_i(yumi_i[133])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_134__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[134]),
    .ready_o(ready_li[134]),
    .v_o(v_o[134]),
    .data_o(data_o[1079:1072]),
    .yumi_i(yumi_i[134])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_135__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[135]),
    .ready_o(ready_li[135]),
    .v_o(v_o[135]),
    .data_o(data_o[1087:1080]),
    .yumi_i(yumi_i[135])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_136__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[136]),
    .ready_o(ready_li[136]),
    .v_o(v_o[136]),
    .data_o(data_o[1095:1088]),
    .yumi_i(yumi_i[136])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_137__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[137]),
    .ready_o(ready_li[137]),
    .v_o(v_o[137]),
    .data_o(data_o[1103:1096]),
    .yumi_i(yumi_i[137])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_138__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[138]),
    .ready_o(ready_li[138]),
    .v_o(v_o[138]),
    .data_o(data_o[1111:1104]),
    .yumi_i(yumi_i[138])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_139__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[139]),
    .ready_o(ready_li[139]),
    .v_o(v_o[139]),
    .data_o(data_o[1119:1112]),
    .yumi_i(yumi_i[139])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_140__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[140]),
    .ready_o(ready_li[140]),
    .v_o(v_o[140]),
    .data_o(data_o[1127:1120]),
    .yumi_i(yumi_i[140])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_141__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[141]),
    .ready_o(ready_li[141]),
    .v_o(v_o[141]),
    .data_o(data_o[1135:1128]),
    .yumi_i(yumi_i[141])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_142__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[142]),
    .ready_o(ready_li[142]),
    .v_o(v_o[142]),
    .data_o(data_o[1143:1136]),
    .yumi_i(yumi_i[142])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_143__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[143]),
    .ready_o(ready_li[143]),
    .v_o(v_o[143]),
    .data_o(data_o[1151:1144]),
    .yumi_i(yumi_i[143])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_144__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[144]),
    .ready_o(ready_li[144]),
    .v_o(v_o[144]),
    .data_o(data_o[1159:1152]),
    .yumi_i(yumi_i[144])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_145__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[145]),
    .ready_o(ready_li[145]),
    .v_o(v_o[145]),
    .data_o(data_o[1167:1160]),
    .yumi_i(yumi_i[145])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_146__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[146]),
    .ready_o(ready_li[146]),
    .v_o(v_o[146]),
    .data_o(data_o[1175:1168]),
    .yumi_i(yumi_i[146])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_147__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[147]),
    .ready_o(ready_li[147]),
    .v_o(v_o[147]),
    .data_o(data_o[1183:1176]),
    .yumi_i(yumi_i[147])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_148__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[148]),
    .ready_o(ready_li[148]),
    .v_o(v_o[148]),
    .data_o(data_o[1191:1184]),
    .yumi_i(yumi_i[148])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_149__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[149]),
    .ready_o(ready_li[149]),
    .v_o(v_o[149]),
    .data_o(data_o[1199:1192]),
    .yumi_i(yumi_i[149])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_150__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[150]),
    .ready_o(ready_li[150]),
    .v_o(v_o[150]),
    .data_o(data_o[1207:1200]),
    .yumi_i(yumi_i[150])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_151__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[151]),
    .ready_o(ready_li[151]),
    .v_o(v_o[151]),
    .data_o(data_o[1215:1208]),
    .yumi_i(yumi_i[151])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_152__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[152]),
    .ready_o(ready_li[152]),
    .v_o(v_o[152]),
    .data_o(data_o[1223:1216]),
    .yumi_i(yumi_i[152])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_153__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[153]),
    .ready_o(ready_li[153]),
    .v_o(v_o[153]),
    .data_o(data_o[1231:1224]),
    .yumi_i(yumi_i[153])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_154__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[154]),
    .ready_o(ready_li[154]),
    .v_o(v_o[154]),
    .data_o(data_o[1239:1232]),
    .yumi_i(yumi_i[154])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_155__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[155]),
    .ready_o(ready_li[155]),
    .v_o(v_o[155]),
    .data_o(data_o[1247:1240]),
    .yumi_i(yumi_i[155])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_156__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[156]),
    .ready_o(ready_li[156]),
    .v_o(v_o[156]),
    .data_o(data_o[1255:1248]),
    .yumi_i(yumi_i[156])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_157__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[157]),
    .ready_o(ready_li[157]),
    .v_o(v_o[157]),
    .data_o(data_o[1263:1256]),
    .yumi_i(yumi_i[157])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_158__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[158]),
    .ready_o(ready_li[158]),
    .v_o(v_o[158]),
    .data_o(data_o[1271:1264]),
    .yumi_i(yumi_i[158])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_159__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[159]),
    .ready_o(ready_li[159]),
    .v_o(v_o[159]),
    .data_o(data_o[1279:1272]),
    .yumi_i(yumi_i[159])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_160__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[160]),
    .ready_o(ready_li[160]),
    .v_o(v_o[160]),
    .data_o(data_o[1287:1280]),
    .yumi_i(yumi_i[160])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_161__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[161]),
    .ready_o(ready_li[161]),
    .v_o(v_o[161]),
    .data_o(data_o[1295:1288]),
    .yumi_i(yumi_i[161])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_162__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[162]),
    .ready_o(ready_li[162]),
    .v_o(v_o[162]),
    .data_o(data_o[1303:1296]),
    .yumi_i(yumi_i[162])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_163__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[163]),
    .ready_o(ready_li[163]),
    .v_o(v_o[163]),
    .data_o(data_o[1311:1304]),
    .yumi_i(yumi_i[163])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_164__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[164]),
    .ready_o(ready_li[164]),
    .v_o(v_o[164]),
    .data_o(data_o[1319:1312]),
    .yumi_i(yumi_i[164])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_165__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[165]),
    .ready_o(ready_li[165]),
    .v_o(v_o[165]),
    .data_o(data_o[1327:1320]),
    .yumi_i(yumi_i[165])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_166__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[166]),
    .ready_o(ready_li[166]),
    .v_o(v_o[166]),
    .data_o(data_o[1335:1328]),
    .yumi_i(yumi_i[166])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_167__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[167]),
    .ready_o(ready_li[167]),
    .v_o(v_o[167]),
    .data_o(data_o[1343:1336]),
    .yumi_i(yumi_i[167])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_168__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[168]),
    .ready_o(ready_li[168]),
    .v_o(v_o[168]),
    .data_o(data_o[1351:1344]),
    .yumi_i(yumi_i[168])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_169__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[169]),
    .ready_o(ready_li[169]),
    .v_o(v_o[169]),
    .data_o(data_o[1359:1352]),
    .yumi_i(yumi_i[169])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_170__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[170]),
    .ready_o(ready_li[170]),
    .v_o(v_o[170]),
    .data_o(data_o[1367:1360]),
    .yumi_i(yumi_i[170])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_171__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[171]),
    .ready_o(ready_li[171]),
    .v_o(v_o[171]),
    .data_o(data_o[1375:1368]),
    .yumi_i(yumi_i[171])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_172__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[172]),
    .ready_o(ready_li[172]),
    .v_o(v_o[172]),
    .data_o(data_o[1383:1376]),
    .yumi_i(yumi_i[172])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_173__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[173]),
    .ready_o(ready_li[173]),
    .v_o(v_o[173]),
    .data_o(data_o[1391:1384]),
    .yumi_i(yumi_i[173])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_174__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[174]),
    .ready_o(ready_li[174]),
    .v_o(v_o[174]),
    .data_o(data_o[1399:1392]),
    .yumi_i(yumi_i[174])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_175__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[175]),
    .ready_o(ready_li[175]),
    .v_o(v_o[175]),
    .data_o(data_o[1407:1400]),
    .yumi_i(yumi_i[175])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_176__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[176]),
    .ready_o(ready_li[176]),
    .v_o(v_o[176]),
    .data_o(data_o[1415:1408]),
    .yumi_i(yumi_i[176])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_177__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[177]),
    .ready_o(ready_li[177]),
    .v_o(v_o[177]),
    .data_o(data_o[1423:1416]),
    .yumi_i(yumi_i[177])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_178__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[178]),
    .ready_o(ready_li[178]),
    .v_o(v_o[178]),
    .data_o(data_o[1431:1424]),
    .yumi_i(yumi_i[178])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_179__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[179]),
    .ready_o(ready_li[179]),
    .v_o(v_o[179]),
    .data_o(data_o[1439:1432]),
    .yumi_i(yumi_i[179])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_180__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[180]),
    .ready_o(ready_li[180]),
    .v_o(v_o[180]),
    .data_o(data_o[1447:1440]),
    .yumi_i(yumi_i[180])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_181__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[181]),
    .ready_o(ready_li[181]),
    .v_o(v_o[181]),
    .data_o(data_o[1455:1448]),
    .yumi_i(yumi_i[181])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_182__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[182]),
    .ready_o(ready_li[182]),
    .v_o(v_o[182]),
    .data_o(data_o[1463:1456]),
    .yumi_i(yumi_i[182])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_183__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[183]),
    .ready_o(ready_li[183]),
    .v_o(v_o[183]),
    .data_o(data_o[1471:1464]),
    .yumi_i(yumi_i[183])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_184__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[184]),
    .ready_o(ready_li[184]),
    .v_o(v_o[184]),
    .data_o(data_o[1479:1472]),
    .yumi_i(yumi_i[184])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_185__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[185]),
    .ready_o(ready_li[185]),
    .v_o(v_o[185]),
    .data_o(data_o[1487:1480]),
    .yumi_i(yumi_i[185])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_186__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[186]),
    .ready_o(ready_li[186]),
    .v_o(v_o[186]),
    .data_o(data_o[1495:1488]),
    .yumi_i(yumi_i[186])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_187__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[187]),
    .ready_o(ready_li[187]),
    .v_o(v_o[187]),
    .data_o(data_o[1503:1496]),
    .yumi_i(yumi_i[187])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_188__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[188]),
    .ready_o(ready_li[188]),
    .v_o(v_o[188]),
    .data_o(data_o[1511:1504]),
    .yumi_i(yumi_i[188])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_189__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[189]),
    .ready_o(ready_li[189]),
    .v_o(v_o[189]),
    .data_o(data_o[1519:1512]),
    .yumi_i(yumi_i[189])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_190__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[190]),
    .ready_o(ready_li[190]),
    .v_o(v_o[190]),
    .data_o(data_o[1527:1520]),
    .yumi_i(yumi_i[190])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_191__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[191]),
    .ready_o(ready_li[191]),
    .v_o(v_o[191]),
    .data_o(data_o[1535:1528]),
    .yumi_i(yumi_i[191])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_192__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[192]),
    .ready_o(ready_li[192]),
    .v_o(v_o[192]),
    .data_o(data_o[1543:1536]),
    .yumi_i(yumi_i[192])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_193__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[193]),
    .ready_o(ready_li[193]),
    .v_o(v_o[193]),
    .data_o(data_o[1551:1544]),
    .yumi_i(yumi_i[193])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_194__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[194]),
    .ready_o(ready_li[194]),
    .v_o(v_o[194]),
    .data_o(data_o[1559:1552]),
    .yumi_i(yumi_i[194])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_195__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[195]),
    .ready_o(ready_li[195]),
    .v_o(v_o[195]),
    .data_o(data_o[1567:1560]),
    .yumi_i(yumi_i[195])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_196__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[196]),
    .ready_o(ready_li[196]),
    .v_o(v_o[196]),
    .data_o(data_o[1575:1568]),
    .yumi_i(yumi_i[196])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_197__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[197]),
    .ready_o(ready_li[197]),
    .v_o(v_o[197]),
    .data_o(data_o[1583:1576]),
    .yumi_i(yumi_i[197])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_198__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[198]),
    .ready_o(ready_li[198]),
    .v_o(v_o[198]),
    .data_o(data_o[1591:1584]),
    .yumi_i(yumi_i[198])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_199__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[199]),
    .ready_o(ready_li[199]),
    .v_o(v_o[199]),
    .data_o(data_o[1599:1592]),
    .yumi_i(yumi_i[199])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_200__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[200]),
    .ready_o(ready_li[200]),
    .v_o(v_o[200]),
    .data_o(data_o[1607:1600]),
    .yumi_i(yumi_i[200])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_201__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[201]),
    .ready_o(ready_li[201]),
    .v_o(v_o[201]),
    .data_o(data_o[1615:1608]),
    .yumi_i(yumi_i[201])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_202__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[202]),
    .ready_o(ready_li[202]),
    .v_o(v_o[202]),
    .data_o(data_o[1623:1616]),
    .yumi_i(yumi_i[202])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_203__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[203]),
    .ready_o(ready_li[203]),
    .v_o(v_o[203]),
    .data_o(data_o[1631:1624]),
    .yumi_i(yumi_i[203])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_204__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[204]),
    .ready_o(ready_li[204]),
    .v_o(v_o[204]),
    .data_o(data_o[1639:1632]),
    .yumi_i(yumi_i[204])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_205__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[205]),
    .ready_o(ready_li[205]),
    .v_o(v_o[205]),
    .data_o(data_o[1647:1640]),
    .yumi_i(yumi_i[205])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_206__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[206]),
    .ready_o(ready_li[206]),
    .v_o(v_o[206]),
    .data_o(data_o[1655:1648]),
    .yumi_i(yumi_i[206])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_207__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[207]),
    .ready_o(ready_li[207]),
    .v_o(v_o[207]),
    .data_o(data_o[1663:1656]),
    .yumi_i(yumi_i[207])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_208__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[208]),
    .ready_o(ready_li[208]),
    .v_o(v_o[208]),
    .data_o(data_o[1671:1664]),
    .yumi_i(yumi_i[208])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_209__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[209]),
    .ready_o(ready_li[209]),
    .v_o(v_o[209]),
    .data_o(data_o[1679:1672]),
    .yumi_i(yumi_i[209])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_210__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[210]),
    .ready_o(ready_li[210]),
    .v_o(v_o[210]),
    .data_o(data_o[1687:1680]),
    .yumi_i(yumi_i[210])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_211__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[211]),
    .ready_o(ready_li[211]),
    .v_o(v_o[211]),
    .data_o(data_o[1695:1688]),
    .yumi_i(yumi_i[211])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_212__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[212]),
    .ready_o(ready_li[212]),
    .v_o(v_o[212]),
    .data_o(data_o[1703:1696]),
    .yumi_i(yumi_i[212])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_213__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[213]),
    .ready_o(ready_li[213]),
    .v_o(v_o[213]),
    .data_o(data_o[1711:1704]),
    .yumi_i(yumi_i[213])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_214__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[214]),
    .ready_o(ready_li[214]),
    .v_o(v_o[214]),
    .data_o(data_o[1719:1712]),
    .yumi_i(yumi_i[214])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_215__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[215]),
    .ready_o(ready_li[215]),
    .v_o(v_o[215]),
    .data_o(data_o[1727:1720]),
    .yumi_i(yumi_i[215])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_216__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[216]),
    .ready_o(ready_li[216]),
    .v_o(v_o[216]),
    .data_o(data_o[1735:1728]),
    .yumi_i(yumi_i[216])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_217__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[217]),
    .ready_o(ready_li[217]),
    .v_o(v_o[217]),
    .data_o(data_o[1743:1736]),
    .yumi_i(yumi_i[217])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_218__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[218]),
    .ready_o(ready_li[218]),
    .v_o(v_o[218]),
    .data_o(data_o[1751:1744]),
    .yumi_i(yumi_i[218])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_219__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[219]),
    .ready_o(ready_li[219]),
    .v_o(v_o[219]),
    .data_o(data_o[1759:1752]),
    .yumi_i(yumi_i[219])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_220__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[220]),
    .ready_o(ready_li[220]),
    .v_o(v_o[220]),
    .data_o(data_o[1767:1760]),
    .yumi_i(yumi_i[220])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_221__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[221]),
    .ready_o(ready_li[221]),
    .v_o(v_o[221]),
    .data_o(data_o[1775:1768]),
    .yumi_i(yumi_i[221])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_222__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[222]),
    .ready_o(ready_li[222]),
    .v_o(v_o[222]),
    .data_o(data_o[1783:1776]),
    .yumi_i(yumi_i[222])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_223__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[223]),
    .ready_o(ready_li[223]),
    .v_o(v_o[223]),
    .data_o(data_o[1791:1784]),
    .yumi_i(yumi_i[223])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_224__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[224]),
    .ready_o(ready_li[224]),
    .v_o(v_o[224]),
    .data_o(data_o[1799:1792]),
    .yumi_i(yumi_i[224])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_225__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[225]),
    .ready_o(ready_li[225]),
    .v_o(v_o[225]),
    .data_o(data_o[1807:1800]),
    .yumi_i(yumi_i[225])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_226__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[226]),
    .ready_o(ready_li[226]),
    .v_o(v_o[226]),
    .data_o(data_o[1815:1808]),
    .yumi_i(yumi_i[226])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_227__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[227]),
    .ready_o(ready_li[227]),
    .v_o(v_o[227]),
    .data_o(data_o[1823:1816]),
    .yumi_i(yumi_i[227])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_228__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[228]),
    .ready_o(ready_li[228]),
    .v_o(v_o[228]),
    .data_o(data_o[1831:1824]),
    .yumi_i(yumi_i[228])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_229__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[229]),
    .ready_o(ready_li[229]),
    .v_o(v_o[229]),
    .data_o(data_o[1839:1832]),
    .yumi_i(yumi_i[229])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_230__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[230]),
    .ready_o(ready_li[230]),
    .v_o(v_o[230]),
    .data_o(data_o[1847:1840]),
    .yumi_i(yumi_i[230])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_231__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[231]),
    .ready_o(ready_li[231]),
    .v_o(v_o[231]),
    .data_o(data_o[1855:1848]),
    .yumi_i(yumi_i[231])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_232__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[232]),
    .ready_o(ready_li[232]),
    .v_o(v_o[232]),
    .data_o(data_o[1863:1856]),
    .yumi_i(yumi_i[232])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_233__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[233]),
    .ready_o(ready_li[233]),
    .v_o(v_o[233]),
    .data_o(data_o[1871:1864]),
    .yumi_i(yumi_i[233])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_234__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[234]),
    .ready_o(ready_li[234]),
    .v_o(v_o[234]),
    .data_o(data_o[1879:1872]),
    .yumi_i(yumi_i[234])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_235__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[235]),
    .ready_o(ready_li[235]),
    .v_o(v_o[235]),
    .data_o(data_o[1887:1880]),
    .yumi_i(yumi_i[235])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_236__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[236]),
    .ready_o(ready_li[236]),
    .v_o(v_o[236]),
    .data_o(data_o[1895:1888]),
    .yumi_i(yumi_i[236])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_237__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[237]),
    .ready_o(ready_li[237]),
    .v_o(v_o[237]),
    .data_o(data_o[1903:1896]),
    .yumi_i(yumi_i[237])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_238__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[238]),
    .ready_o(ready_li[238]),
    .v_o(v_o[238]),
    .data_o(data_o[1911:1904]),
    .yumi_i(yumi_i[238])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_239__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[239]),
    .ready_o(ready_li[239]),
    .v_o(v_o[239]),
    .data_o(data_o[1919:1912]),
    .yumi_i(yumi_i[239])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_240__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[240]),
    .ready_o(ready_li[240]),
    .v_o(v_o[240]),
    .data_o(data_o[1927:1920]),
    .yumi_i(yumi_i[240])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_241__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[241]),
    .ready_o(ready_li[241]),
    .v_o(v_o[241]),
    .data_o(data_o[1935:1928]),
    .yumi_i(yumi_i[241])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_242__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[242]),
    .ready_o(ready_li[242]),
    .v_o(v_o[242]),
    .data_o(data_o[1943:1936]),
    .yumi_i(yumi_i[242])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_243__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[243]),
    .ready_o(ready_li[243]),
    .v_o(v_o[243]),
    .data_o(data_o[1951:1944]),
    .yumi_i(yumi_i[243])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_244__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[244]),
    .ready_o(ready_li[244]),
    .v_o(v_o[244]),
    .data_o(data_o[1959:1952]),
    .yumi_i(yumi_i[244])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_245__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[245]),
    .ready_o(ready_li[245]),
    .v_o(v_o[245]),
    .data_o(data_o[1967:1960]),
    .yumi_i(yumi_i[245])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_246__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[246]),
    .ready_o(ready_li[246]),
    .v_o(v_o[246]),
    .data_o(data_o[1975:1968]),
    .yumi_i(yumi_i[246])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_247__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[247]),
    .ready_o(ready_li[247]),
    .v_o(v_o[247]),
    .data_o(data_o[1983:1976]),
    .yumi_i(yumi_i[247])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_248__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[248]),
    .ready_o(ready_li[248]),
    .v_o(v_o[248]),
    .data_o(data_o[1991:1984]),
    .yumi_i(yumi_i[248])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_249__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[249]),
    .ready_o(ready_li[249]),
    .v_o(v_o[249]),
    .data_o(data_o[1999:1992]),
    .yumi_i(yumi_i[249])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_250__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[250]),
    .ready_o(ready_li[250]),
    .v_o(v_o[250]),
    .data_o(data_o[2007:2000]),
    .yumi_i(yumi_i[250])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_251__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[251]),
    .ready_o(ready_li[251]),
    .v_o(v_o[251]),
    .data_o(data_o[2015:2008]),
    .yumi_i(yumi_i[251])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_252__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[252]),
    .ready_o(ready_li[252]),
    .v_o(v_o[252]),
    .data_o(data_o[2023:2016]),
    .yumi_i(yumi_i[252])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_253__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[253]),
    .ready_o(ready_li[253]),
    .v_o(v_o[253]),
    .data_o(data_o[2031:2024]),
    .yumi_i(yumi_i[253])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_254__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[254]),
    .ready_o(ready_li[254]),
    .v_o(v_o[254]),
    .data_o(data_o[2039:2032]),
    .yumi_i(yumi_i[254])
  );


  bsg_fifo_1r1w_pseudo_large_width_p8_els_p8
  rof_255__psdlrg_fifo
  (
    .clk_i(clk_i),
    .reset_i(reset_i),
    .data_i(data_i),
    .v_i(valid_lo[255]),
    .ready_o(ready_li[255]),
    .v_o(v_o[255]),
    .data_o(data_o[2047:2040]),
    .yumi_i(yumi_i[255])
  );


endmodule

