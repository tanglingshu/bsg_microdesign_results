

module top
(
  gray_i,
  binary_o
);

  input [127:0] gray_i;
  output [127:0] binary_o;

  bsg_gray_to_binary
  wrapper
  (
    .gray_i(gray_i),
    .binary_o(binary_o)
  );


endmodule



module bsg_scan_width_p128_xor_p1
(
  i,
  o
);

  input [127:0] i;
  output [127:0] o;
  wire [127:0] o;
  wire t_3__127_,t_3__126_,t_3__125_,t_3__124_,t_3__123_,t_3__122_,t_3__121_,t_3__120_,
  t_3__119_,t_3__118_,t_3__117_,t_3__116_,t_3__115_,t_3__114_,t_3__113_,t_3__112_,
  t_3__111_,t_3__110_,t_3__109_,t_3__108_,t_3__107_,t_3__106_,t_3__105_,t_3__104_,
  t_3__103_,t_3__102_,t_3__101_,t_3__100_,t_3__99_,t_3__98_,t_3__97_,t_3__96_,
  t_3__95_,t_3__94_,t_3__93_,t_3__92_,t_3__91_,t_3__90_,t_3__89_,t_3__88_,t_3__87_,
  t_3__86_,t_3__85_,t_3__84_,t_3__83_,t_3__82_,t_3__81_,t_3__80_,t_3__79_,t_3__78_,
  t_3__77_,t_3__76_,t_3__75_,t_3__74_,t_3__73_,t_3__72_,t_3__71_,t_3__70_,t_3__69_,
  t_3__68_,t_3__67_,t_3__66_,t_3__65_,t_3__64_,t_3__63_,t_3__62_,t_3__61_,t_3__60_,
  t_3__59_,t_3__58_,t_3__57_,t_3__56_,t_3__55_,t_3__54_,t_3__53_,t_3__52_,
  t_3__51_,t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,t_3__45_,t_3__44_,t_3__43_,
  t_3__42_,t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,t_3__36_,t_3__35_,t_3__34_,
  t_3__33_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,t_3__26_,t_3__25_,
  t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,t_3__17_,t_3__16_,
  t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,t_3__7_,
  t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_2__127_,t_2__126_,t_2__125_,
  t_2__124_,t_2__123_,t_2__122_,t_2__121_,t_2__120_,t_2__119_,t_2__118_,t_2__117_,
  t_2__116_,t_2__115_,t_2__114_,t_2__113_,t_2__112_,t_2__111_,t_2__110_,t_2__109_,
  t_2__108_,t_2__107_,t_2__106_,t_2__105_,t_2__104_,t_2__103_,t_2__102_,t_2__101_,
  t_2__100_,t_2__99_,t_2__98_,t_2__97_,t_2__96_,t_2__95_,t_2__94_,t_2__93_,
  t_2__92_,t_2__91_,t_2__90_,t_2__89_,t_2__88_,t_2__87_,t_2__86_,t_2__85_,t_2__84_,
  t_2__83_,t_2__82_,t_2__81_,t_2__80_,t_2__79_,t_2__78_,t_2__77_,t_2__76_,t_2__75_,
  t_2__74_,t_2__73_,t_2__72_,t_2__71_,t_2__70_,t_2__69_,t_2__68_,t_2__67_,t_2__66_,
  t_2__65_,t_2__64_,t_2__63_,t_2__62_,t_2__61_,t_2__60_,t_2__59_,t_2__58_,t_2__57_,
  t_2__56_,t_2__55_,t_2__54_,t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,t_2__48_,
  t_2__47_,t_2__46_,t_2__45_,t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,t_2__39_,
  t_2__38_,t_2__37_,t_2__36_,t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,t_2__30_,
  t_2__29_,t_2__28_,t_2__27_,t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,
  t_2__21_,t_2__20_,t_2__19_,t_2__18_,t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,
  t_2__12_,t_2__11_,t_2__10_,t_2__9_,t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,
  t_2__2_,t_2__1_,t_2__0_,t_1__127_,t_1__126_,t_1__125_,t_1__124_,t_1__123_,t_1__122_,
  t_1__121_,t_1__120_,t_1__119_,t_1__118_,t_1__117_,t_1__116_,t_1__115_,t_1__114_,
  t_1__113_,t_1__112_,t_1__111_,t_1__110_,t_1__109_,t_1__108_,t_1__107_,t_1__106_,
  t_1__105_,t_1__104_,t_1__103_,t_1__102_,t_1__101_,t_1__100_,t_1__99_,t_1__98_,
  t_1__97_,t_1__96_,t_1__95_,t_1__94_,t_1__93_,t_1__92_,t_1__91_,t_1__90_,t_1__89_,
  t_1__88_,t_1__87_,t_1__86_,t_1__85_,t_1__84_,t_1__83_,t_1__82_,t_1__81_,t_1__80_,
  t_1__79_,t_1__78_,t_1__77_,t_1__76_,t_1__75_,t_1__74_,t_1__73_,t_1__72_,
  t_1__71_,t_1__70_,t_1__69_,t_1__68_,t_1__67_,t_1__66_,t_1__65_,t_1__64_,t_1__63_,
  t_1__62_,t_1__61_,t_1__60_,t_1__59_,t_1__58_,t_1__57_,t_1__56_,t_1__55_,t_1__54_,
  t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,t_1__48_,t_1__47_,t_1__46_,t_1__45_,
  t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,t_1__39_,t_1__38_,t_1__37_,t_1__36_,
  t_1__35_,t_1__34_,t_1__33_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,t_1__27_,
  t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,t_1__18_,
  t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,t_1__9_,
  t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_,t_6__127_,
  t_6__126_,t_6__125_,t_6__124_,t_6__123_,t_6__122_,t_6__121_,t_6__120_,t_6__119_,
  t_6__118_,t_6__117_,t_6__116_,t_6__115_,t_6__114_,t_6__113_,t_6__112_,t_6__111_,
  t_6__110_,t_6__109_,t_6__108_,t_6__107_,t_6__106_,t_6__105_,t_6__104_,t_6__103_,
  t_6__102_,t_6__101_,t_6__100_,t_6__99_,t_6__98_,t_6__97_,t_6__96_,t_6__95_,
  t_6__94_,t_6__93_,t_6__92_,t_6__91_,t_6__90_,t_6__89_,t_6__88_,t_6__87_,t_6__86_,
  t_6__85_,t_6__84_,t_6__83_,t_6__82_,t_6__81_,t_6__80_,t_6__79_,t_6__78_,t_6__77_,
  t_6__76_,t_6__75_,t_6__74_,t_6__73_,t_6__72_,t_6__71_,t_6__70_,t_6__69_,t_6__68_,
  t_6__67_,t_6__66_,t_6__65_,t_6__64_,t_6__63_,t_6__62_,t_6__61_,t_6__60_,t_6__59_,
  t_6__58_,t_6__57_,t_6__56_,t_6__55_,t_6__54_,t_6__53_,t_6__52_,t_6__51_,t_6__50_,
  t_6__49_,t_6__48_,t_6__47_,t_6__46_,t_6__45_,t_6__44_,t_6__43_,t_6__42_,
  t_6__41_,t_6__40_,t_6__39_,t_6__38_,t_6__37_,t_6__36_,t_6__35_,t_6__34_,t_6__33_,
  t_6__32_,t_6__31_,t_6__30_,t_6__29_,t_6__28_,t_6__27_,t_6__26_,t_6__25_,t_6__24_,
  t_6__23_,t_6__22_,t_6__21_,t_6__20_,t_6__19_,t_6__18_,t_6__17_,t_6__16_,t_6__15_,
  t_6__14_,t_6__13_,t_6__12_,t_6__11_,t_6__10_,t_6__9_,t_6__8_,t_6__7_,t_6__6_,t_6__5_,
  t_6__4_,t_6__3_,t_6__2_,t_6__1_,t_6__0_,t_5__127_,t_5__126_,t_5__125_,t_5__124_,
  t_5__123_,t_5__122_,t_5__121_,t_5__120_,t_5__119_,t_5__118_,t_5__117_,t_5__116_,
  t_5__115_,t_5__114_,t_5__113_,t_5__112_,t_5__111_,t_5__110_,t_5__109_,t_5__108_,
  t_5__107_,t_5__106_,t_5__105_,t_5__104_,t_5__103_,t_5__102_,t_5__101_,t_5__100_,
  t_5__99_,t_5__98_,t_5__97_,t_5__96_,t_5__95_,t_5__94_,t_5__93_,t_5__92_,
  t_5__91_,t_5__90_,t_5__89_,t_5__88_,t_5__87_,t_5__86_,t_5__85_,t_5__84_,t_5__83_,
  t_5__82_,t_5__81_,t_5__80_,t_5__79_,t_5__78_,t_5__77_,t_5__76_,t_5__75_,t_5__74_,
  t_5__73_,t_5__72_,t_5__71_,t_5__70_,t_5__69_,t_5__68_,t_5__67_,t_5__66_,t_5__65_,
  t_5__64_,t_5__63_,t_5__62_,t_5__61_,t_5__60_,t_5__59_,t_5__58_,t_5__57_,t_5__56_,
  t_5__55_,t_5__54_,t_5__53_,t_5__52_,t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,
  t_5__46_,t_5__45_,t_5__44_,t_5__43_,t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,
  t_5__37_,t_5__36_,t_5__35_,t_5__34_,t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,
  t_5__28_,t_5__27_,t_5__26_,t_5__25_,t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,
  t_5__19_,t_5__18_,t_5__17_,t_5__16_,t_5__15_,t_5__14_,t_5__13_,t_5__12_,
  t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,
  t_5__1_,t_5__0_,t_4__127_,t_4__126_,t_4__125_,t_4__124_,t_4__123_,t_4__122_,t_4__121_,
  t_4__120_,t_4__119_,t_4__118_,t_4__117_,t_4__116_,t_4__115_,t_4__114_,t_4__113_,
  t_4__112_,t_4__111_,t_4__110_,t_4__109_,t_4__108_,t_4__107_,t_4__106_,t_4__105_,
  t_4__104_,t_4__103_,t_4__102_,t_4__101_,t_4__100_,t_4__99_,t_4__98_,t_4__97_,
  t_4__96_,t_4__95_,t_4__94_,t_4__93_,t_4__92_,t_4__91_,t_4__90_,t_4__89_,t_4__88_,
  t_4__87_,t_4__86_,t_4__85_,t_4__84_,t_4__83_,t_4__82_,t_4__81_,t_4__80_,t_4__79_,
  t_4__78_,t_4__77_,t_4__76_,t_4__75_,t_4__74_,t_4__73_,t_4__72_,t_4__71_,t_4__70_,
  t_4__69_,t_4__68_,t_4__67_,t_4__66_,t_4__65_,t_4__64_,t_4__63_,t_4__62_,
  t_4__61_,t_4__60_,t_4__59_,t_4__58_,t_4__57_,t_4__56_,t_4__55_,t_4__54_,t_4__53_,
  t_4__52_,t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,
  t_4__43_,t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,
  t_4__34_,t_4__33_,t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,
  t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,
  t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,
  t_4__7_,t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_;
  assign t_1__127_ = i[127] ^ 1'b0;
  assign t_1__126_ = i[126] ^ i[127];
  assign t_1__125_ = i[125] ^ i[126];
  assign t_1__124_ = i[124] ^ i[125];
  assign t_1__123_ = i[123] ^ i[124];
  assign t_1__122_ = i[122] ^ i[123];
  assign t_1__121_ = i[121] ^ i[122];
  assign t_1__120_ = i[120] ^ i[121];
  assign t_1__119_ = i[119] ^ i[120];
  assign t_1__118_ = i[118] ^ i[119];
  assign t_1__117_ = i[117] ^ i[118];
  assign t_1__116_ = i[116] ^ i[117];
  assign t_1__115_ = i[115] ^ i[116];
  assign t_1__114_ = i[114] ^ i[115];
  assign t_1__113_ = i[113] ^ i[114];
  assign t_1__112_ = i[112] ^ i[113];
  assign t_1__111_ = i[111] ^ i[112];
  assign t_1__110_ = i[110] ^ i[111];
  assign t_1__109_ = i[109] ^ i[110];
  assign t_1__108_ = i[108] ^ i[109];
  assign t_1__107_ = i[107] ^ i[108];
  assign t_1__106_ = i[106] ^ i[107];
  assign t_1__105_ = i[105] ^ i[106];
  assign t_1__104_ = i[104] ^ i[105];
  assign t_1__103_ = i[103] ^ i[104];
  assign t_1__102_ = i[102] ^ i[103];
  assign t_1__101_ = i[101] ^ i[102];
  assign t_1__100_ = i[100] ^ i[101];
  assign t_1__99_ = i[99] ^ i[100];
  assign t_1__98_ = i[98] ^ i[99];
  assign t_1__97_ = i[97] ^ i[98];
  assign t_1__96_ = i[96] ^ i[97];
  assign t_1__95_ = i[95] ^ i[96];
  assign t_1__94_ = i[94] ^ i[95];
  assign t_1__93_ = i[93] ^ i[94];
  assign t_1__92_ = i[92] ^ i[93];
  assign t_1__91_ = i[91] ^ i[92];
  assign t_1__90_ = i[90] ^ i[91];
  assign t_1__89_ = i[89] ^ i[90];
  assign t_1__88_ = i[88] ^ i[89];
  assign t_1__87_ = i[87] ^ i[88];
  assign t_1__86_ = i[86] ^ i[87];
  assign t_1__85_ = i[85] ^ i[86];
  assign t_1__84_ = i[84] ^ i[85];
  assign t_1__83_ = i[83] ^ i[84];
  assign t_1__82_ = i[82] ^ i[83];
  assign t_1__81_ = i[81] ^ i[82];
  assign t_1__80_ = i[80] ^ i[81];
  assign t_1__79_ = i[79] ^ i[80];
  assign t_1__78_ = i[78] ^ i[79];
  assign t_1__77_ = i[77] ^ i[78];
  assign t_1__76_ = i[76] ^ i[77];
  assign t_1__75_ = i[75] ^ i[76];
  assign t_1__74_ = i[74] ^ i[75];
  assign t_1__73_ = i[73] ^ i[74];
  assign t_1__72_ = i[72] ^ i[73];
  assign t_1__71_ = i[71] ^ i[72];
  assign t_1__70_ = i[70] ^ i[71];
  assign t_1__69_ = i[69] ^ i[70];
  assign t_1__68_ = i[68] ^ i[69];
  assign t_1__67_ = i[67] ^ i[68];
  assign t_1__66_ = i[66] ^ i[67];
  assign t_1__65_ = i[65] ^ i[66];
  assign t_1__64_ = i[64] ^ i[65];
  assign t_1__63_ = i[63] ^ i[64];
  assign t_1__62_ = i[62] ^ i[63];
  assign t_1__61_ = i[61] ^ i[62];
  assign t_1__60_ = i[60] ^ i[61];
  assign t_1__59_ = i[59] ^ i[60];
  assign t_1__58_ = i[58] ^ i[59];
  assign t_1__57_ = i[57] ^ i[58];
  assign t_1__56_ = i[56] ^ i[57];
  assign t_1__55_ = i[55] ^ i[56];
  assign t_1__54_ = i[54] ^ i[55];
  assign t_1__53_ = i[53] ^ i[54];
  assign t_1__52_ = i[52] ^ i[53];
  assign t_1__51_ = i[51] ^ i[52];
  assign t_1__50_ = i[50] ^ i[51];
  assign t_1__49_ = i[49] ^ i[50];
  assign t_1__48_ = i[48] ^ i[49];
  assign t_1__47_ = i[47] ^ i[48];
  assign t_1__46_ = i[46] ^ i[47];
  assign t_1__45_ = i[45] ^ i[46];
  assign t_1__44_ = i[44] ^ i[45];
  assign t_1__43_ = i[43] ^ i[44];
  assign t_1__42_ = i[42] ^ i[43];
  assign t_1__41_ = i[41] ^ i[42];
  assign t_1__40_ = i[40] ^ i[41];
  assign t_1__39_ = i[39] ^ i[40];
  assign t_1__38_ = i[38] ^ i[39];
  assign t_1__37_ = i[37] ^ i[38];
  assign t_1__36_ = i[36] ^ i[37];
  assign t_1__35_ = i[35] ^ i[36];
  assign t_1__34_ = i[34] ^ i[35];
  assign t_1__33_ = i[33] ^ i[34];
  assign t_1__32_ = i[32] ^ i[33];
  assign t_1__31_ = i[31] ^ i[32];
  assign t_1__30_ = i[30] ^ i[31];
  assign t_1__29_ = i[29] ^ i[30];
  assign t_1__28_ = i[28] ^ i[29];
  assign t_1__27_ = i[27] ^ i[28];
  assign t_1__26_ = i[26] ^ i[27];
  assign t_1__25_ = i[25] ^ i[26];
  assign t_1__24_ = i[24] ^ i[25];
  assign t_1__23_ = i[23] ^ i[24];
  assign t_1__22_ = i[22] ^ i[23];
  assign t_1__21_ = i[21] ^ i[22];
  assign t_1__20_ = i[20] ^ i[21];
  assign t_1__19_ = i[19] ^ i[20];
  assign t_1__18_ = i[18] ^ i[19];
  assign t_1__17_ = i[17] ^ i[18];
  assign t_1__16_ = i[16] ^ i[17];
  assign t_1__15_ = i[15] ^ i[16];
  assign t_1__14_ = i[14] ^ i[15];
  assign t_1__13_ = i[13] ^ i[14];
  assign t_1__12_ = i[12] ^ i[13];
  assign t_1__11_ = i[11] ^ i[12];
  assign t_1__10_ = i[10] ^ i[11];
  assign t_1__9_ = i[9] ^ i[10];
  assign t_1__8_ = i[8] ^ i[9];
  assign t_1__7_ = i[7] ^ i[8];
  assign t_1__6_ = i[6] ^ i[7];
  assign t_1__5_ = i[5] ^ i[6];
  assign t_1__4_ = i[4] ^ i[5];
  assign t_1__3_ = i[3] ^ i[4];
  assign t_1__2_ = i[2] ^ i[3];
  assign t_1__1_ = i[1] ^ i[2];
  assign t_1__0_ = i[0] ^ i[1];
  assign t_2__127_ = t_1__127_ ^ 1'b0;
  assign t_2__126_ = t_1__126_ ^ 1'b0;
  assign t_2__125_ = t_1__125_ ^ t_1__127_;
  assign t_2__124_ = t_1__124_ ^ t_1__126_;
  assign t_2__123_ = t_1__123_ ^ t_1__125_;
  assign t_2__122_ = t_1__122_ ^ t_1__124_;
  assign t_2__121_ = t_1__121_ ^ t_1__123_;
  assign t_2__120_ = t_1__120_ ^ t_1__122_;
  assign t_2__119_ = t_1__119_ ^ t_1__121_;
  assign t_2__118_ = t_1__118_ ^ t_1__120_;
  assign t_2__117_ = t_1__117_ ^ t_1__119_;
  assign t_2__116_ = t_1__116_ ^ t_1__118_;
  assign t_2__115_ = t_1__115_ ^ t_1__117_;
  assign t_2__114_ = t_1__114_ ^ t_1__116_;
  assign t_2__113_ = t_1__113_ ^ t_1__115_;
  assign t_2__112_ = t_1__112_ ^ t_1__114_;
  assign t_2__111_ = t_1__111_ ^ t_1__113_;
  assign t_2__110_ = t_1__110_ ^ t_1__112_;
  assign t_2__109_ = t_1__109_ ^ t_1__111_;
  assign t_2__108_ = t_1__108_ ^ t_1__110_;
  assign t_2__107_ = t_1__107_ ^ t_1__109_;
  assign t_2__106_ = t_1__106_ ^ t_1__108_;
  assign t_2__105_ = t_1__105_ ^ t_1__107_;
  assign t_2__104_ = t_1__104_ ^ t_1__106_;
  assign t_2__103_ = t_1__103_ ^ t_1__105_;
  assign t_2__102_ = t_1__102_ ^ t_1__104_;
  assign t_2__101_ = t_1__101_ ^ t_1__103_;
  assign t_2__100_ = t_1__100_ ^ t_1__102_;
  assign t_2__99_ = t_1__99_ ^ t_1__101_;
  assign t_2__98_ = t_1__98_ ^ t_1__100_;
  assign t_2__97_ = t_1__97_ ^ t_1__99_;
  assign t_2__96_ = t_1__96_ ^ t_1__98_;
  assign t_2__95_ = t_1__95_ ^ t_1__97_;
  assign t_2__94_ = t_1__94_ ^ t_1__96_;
  assign t_2__93_ = t_1__93_ ^ t_1__95_;
  assign t_2__92_ = t_1__92_ ^ t_1__94_;
  assign t_2__91_ = t_1__91_ ^ t_1__93_;
  assign t_2__90_ = t_1__90_ ^ t_1__92_;
  assign t_2__89_ = t_1__89_ ^ t_1__91_;
  assign t_2__88_ = t_1__88_ ^ t_1__90_;
  assign t_2__87_ = t_1__87_ ^ t_1__89_;
  assign t_2__86_ = t_1__86_ ^ t_1__88_;
  assign t_2__85_ = t_1__85_ ^ t_1__87_;
  assign t_2__84_ = t_1__84_ ^ t_1__86_;
  assign t_2__83_ = t_1__83_ ^ t_1__85_;
  assign t_2__82_ = t_1__82_ ^ t_1__84_;
  assign t_2__81_ = t_1__81_ ^ t_1__83_;
  assign t_2__80_ = t_1__80_ ^ t_1__82_;
  assign t_2__79_ = t_1__79_ ^ t_1__81_;
  assign t_2__78_ = t_1__78_ ^ t_1__80_;
  assign t_2__77_ = t_1__77_ ^ t_1__79_;
  assign t_2__76_ = t_1__76_ ^ t_1__78_;
  assign t_2__75_ = t_1__75_ ^ t_1__77_;
  assign t_2__74_ = t_1__74_ ^ t_1__76_;
  assign t_2__73_ = t_1__73_ ^ t_1__75_;
  assign t_2__72_ = t_1__72_ ^ t_1__74_;
  assign t_2__71_ = t_1__71_ ^ t_1__73_;
  assign t_2__70_ = t_1__70_ ^ t_1__72_;
  assign t_2__69_ = t_1__69_ ^ t_1__71_;
  assign t_2__68_ = t_1__68_ ^ t_1__70_;
  assign t_2__67_ = t_1__67_ ^ t_1__69_;
  assign t_2__66_ = t_1__66_ ^ t_1__68_;
  assign t_2__65_ = t_1__65_ ^ t_1__67_;
  assign t_2__64_ = t_1__64_ ^ t_1__66_;
  assign t_2__63_ = t_1__63_ ^ t_1__65_;
  assign t_2__62_ = t_1__62_ ^ t_1__64_;
  assign t_2__61_ = t_1__61_ ^ t_1__63_;
  assign t_2__60_ = t_1__60_ ^ t_1__62_;
  assign t_2__59_ = t_1__59_ ^ t_1__61_;
  assign t_2__58_ = t_1__58_ ^ t_1__60_;
  assign t_2__57_ = t_1__57_ ^ t_1__59_;
  assign t_2__56_ = t_1__56_ ^ t_1__58_;
  assign t_2__55_ = t_1__55_ ^ t_1__57_;
  assign t_2__54_ = t_1__54_ ^ t_1__56_;
  assign t_2__53_ = t_1__53_ ^ t_1__55_;
  assign t_2__52_ = t_1__52_ ^ t_1__54_;
  assign t_2__51_ = t_1__51_ ^ t_1__53_;
  assign t_2__50_ = t_1__50_ ^ t_1__52_;
  assign t_2__49_ = t_1__49_ ^ t_1__51_;
  assign t_2__48_ = t_1__48_ ^ t_1__50_;
  assign t_2__47_ = t_1__47_ ^ t_1__49_;
  assign t_2__46_ = t_1__46_ ^ t_1__48_;
  assign t_2__45_ = t_1__45_ ^ t_1__47_;
  assign t_2__44_ = t_1__44_ ^ t_1__46_;
  assign t_2__43_ = t_1__43_ ^ t_1__45_;
  assign t_2__42_ = t_1__42_ ^ t_1__44_;
  assign t_2__41_ = t_1__41_ ^ t_1__43_;
  assign t_2__40_ = t_1__40_ ^ t_1__42_;
  assign t_2__39_ = t_1__39_ ^ t_1__41_;
  assign t_2__38_ = t_1__38_ ^ t_1__40_;
  assign t_2__37_ = t_1__37_ ^ t_1__39_;
  assign t_2__36_ = t_1__36_ ^ t_1__38_;
  assign t_2__35_ = t_1__35_ ^ t_1__37_;
  assign t_2__34_ = t_1__34_ ^ t_1__36_;
  assign t_2__33_ = t_1__33_ ^ t_1__35_;
  assign t_2__32_ = t_1__32_ ^ t_1__34_;
  assign t_2__31_ = t_1__31_ ^ t_1__33_;
  assign t_2__30_ = t_1__30_ ^ t_1__32_;
  assign t_2__29_ = t_1__29_ ^ t_1__31_;
  assign t_2__28_ = t_1__28_ ^ t_1__30_;
  assign t_2__27_ = t_1__27_ ^ t_1__29_;
  assign t_2__26_ = t_1__26_ ^ t_1__28_;
  assign t_2__25_ = t_1__25_ ^ t_1__27_;
  assign t_2__24_ = t_1__24_ ^ t_1__26_;
  assign t_2__23_ = t_1__23_ ^ t_1__25_;
  assign t_2__22_ = t_1__22_ ^ t_1__24_;
  assign t_2__21_ = t_1__21_ ^ t_1__23_;
  assign t_2__20_ = t_1__20_ ^ t_1__22_;
  assign t_2__19_ = t_1__19_ ^ t_1__21_;
  assign t_2__18_ = t_1__18_ ^ t_1__20_;
  assign t_2__17_ = t_1__17_ ^ t_1__19_;
  assign t_2__16_ = t_1__16_ ^ t_1__18_;
  assign t_2__15_ = t_1__15_ ^ t_1__17_;
  assign t_2__14_ = t_1__14_ ^ t_1__16_;
  assign t_2__13_ = t_1__13_ ^ t_1__15_;
  assign t_2__12_ = t_1__12_ ^ t_1__14_;
  assign t_2__11_ = t_1__11_ ^ t_1__13_;
  assign t_2__10_ = t_1__10_ ^ t_1__12_;
  assign t_2__9_ = t_1__9_ ^ t_1__11_;
  assign t_2__8_ = t_1__8_ ^ t_1__10_;
  assign t_2__7_ = t_1__7_ ^ t_1__9_;
  assign t_2__6_ = t_1__6_ ^ t_1__8_;
  assign t_2__5_ = t_1__5_ ^ t_1__7_;
  assign t_2__4_ = t_1__4_ ^ t_1__6_;
  assign t_2__3_ = t_1__3_ ^ t_1__5_;
  assign t_2__2_ = t_1__2_ ^ t_1__4_;
  assign t_2__1_ = t_1__1_ ^ t_1__3_;
  assign t_2__0_ = t_1__0_ ^ t_1__2_;
  assign t_3__127_ = t_2__127_ ^ 1'b0;
  assign t_3__126_ = t_2__126_ ^ 1'b0;
  assign t_3__125_ = t_2__125_ ^ 1'b0;
  assign t_3__124_ = t_2__124_ ^ 1'b0;
  assign t_3__123_ = t_2__123_ ^ t_2__127_;
  assign t_3__122_ = t_2__122_ ^ t_2__126_;
  assign t_3__121_ = t_2__121_ ^ t_2__125_;
  assign t_3__120_ = t_2__120_ ^ t_2__124_;
  assign t_3__119_ = t_2__119_ ^ t_2__123_;
  assign t_3__118_ = t_2__118_ ^ t_2__122_;
  assign t_3__117_ = t_2__117_ ^ t_2__121_;
  assign t_3__116_ = t_2__116_ ^ t_2__120_;
  assign t_3__115_ = t_2__115_ ^ t_2__119_;
  assign t_3__114_ = t_2__114_ ^ t_2__118_;
  assign t_3__113_ = t_2__113_ ^ t_2__117_;
  assign t_3__112_ = t_2__112_ ^ t_2__116_;
  assign t_3__111_ = t_2__111_ ^ t_2__115_;
  assign t_3__110_ = t_2__110_ ^ t_2__114_;
  assign t_3__109_ = t_2__109_ ^ t_2__113_;
  assign t_3__108_ = t_2__108_ ^ t_2__112_;
  assign t_3__107_ = t_2__107_ ^ t_2__111_;
  assign t_3__106_ = t_2__106_ ^ t_2__110_;
  assign t_3__105_ = t_2__105_ ^ t_2__109_;
  assign t_3__104_ = t_2__104_ ^ t_2__108_;
  assign t_3__103_ = t_2__103_ ^ t_2__107_;
  assign t_3__102_ = t_2__102_ ^ t_2__106_;
  assign t_3__101_ = t_2__101_ ^ t_2__105_;
  assign t_3__100_ = t_2__100_ ^ t_2__104_;
  assign t_3__99_ = t_2__99_ ^ t_2__103_;
  assign t_3__98_ = t_2__98_ ^ t_2__102_;
  assign t_3__97_ = t_2__97_ ^ t_2__101_;
  assign t_3__96_ = t_2__96_ ^ t_2__100_;
  assign t_3__95_ = t_2__95_ ^ t_2__99_;
  assign t_3__94_ = t_2__94_ ^ t_2__98_;
  assign t_3__93_ = t_2__93_ ^ t_2__97_;
  assign t_3__92_ = t_2__92_ ^ t_2__96_;
  assign t_3__91_ = t_2__91_ ^ t_2__95_;
  assign t_3__90_ = t_2__90_ ^ t_2__94_;
  assign t_3__89_ = t_2__89_ ^ t_2__93_;
  assign t_3__88_ = t_2__88_ ^ t_2__92_;
  assign t_3__87_ = t_2__87_ ^ t_2__91_;
  assign t_3__86_ = t_2__86_ ^ t_2__90_;
  assign t_3__85_ = t_2__85_ ^ t_2__89_;
  assign t_3__84_ = t_2__84_ ^ t_2__88_;
  assign t_3__83_ = t_2__83_ ^ t_2__87_;
  assign t_3__82_ = t_2__82_ ^ t_2__86_;
  assign t_3__81_ = t_2__81_ ^ t_2__85_;
  assign t_3__80_ = t_2__80_ ^ t_2__84_;
  assign t_3__79_ = t_2__79_ ^ t_2__83_;
  assign t_3__78_ = t_2__78_ ^ t_2__82_;
  assign t_3__77_ = t_2__77_ ^ t_2__81_;
  assign t_3__76_ = t_2__76_ ^ t_2__80_;
  assign t_3__75_ = t_2__75_ ^ t_2__79_;
  assign t_3__74_ = t_2__74_ ^ t_2__78_;
  assign t_3__73_ = t_2__73_ ^ t_2__77_;
  assign t_3__72_ = t_2__72_ ^ t_2__76_;
  assign t_3__71_ = t_2__71_ ^ t_2__75_;
  assign t_3__70_ = t_2__70_ ^ t_2__74_;
  assign t_3__69_ = t_2__69_ ^ t_2__73_;
  assign t_3__68_ = t_2__68_ ^ t_2__72_;
  assign t_3__67_ = t_2__67_ ^ t_2__71_;
  assign t_3__66_ = t_2__66_ ^ t_2__70_;
  assign t_3__65_ = t_2__65_ ^ t_2__69_;
  assign t_3__64_ = t_2__64_ ^ t_2__68_;
  assign t_3__63_ = t_2__63_ ^ t_2__67_;
  assign t_3__62_ = t_2__62_ ^ t_2__66_;
  assign t_3__61_ = t_2__61_ ^ t_2__65_;
  assign t_3__60_ = t_2__60_ ^ t_2__64_;
  assign t_3__59_ = t_2__59_ ^ t_2__63_;
  assign t_3__58_ = t_2__58_ ^ t_2__62_;
  assign t_3__57_ = t_2__57_ ^ t_2__61_;
  assign t_3__56_ = t_2__56_ ^ t_2__60_;
  assign t_3__55_ = t_2__55_ ^ t_2__59_;
  assign t_3__54_ = t_2__54_ ^ t_2__58_;
  assign t_3__53_ = t_2__53_ ^ t_2__57_;
  assign t_3__52_ = t_2__52_ ^ t_2__56_;
  assign t_3__51_ = t_2__51_ ^ t_2__55_;
  assign t_3__50_ = t_2__50_ ^ t_2__54_;
  assign t_3__49_ = t_2__49_ ^ t_2__53_;
  assign t_3__48_ = t_2__48_ ^ t_2__52_;
  assign t_3__47_ = t_2__47_ ^ t_2__51_;
  assign t_3__46_ = t_2__46_ ^ t_2__50_;
  assign t_3__45_ = t_2__45_ ^ t_2__49_;
  assign t_3__44_ = t_2__44_ ^ t_2__48_;
  assign t_3__43_ = t_2__43_ ^ t_2__47_;
  assign t_3__42_ = t_2__42_ ^ t_2__46_;
  assign t_3__41_ = t_2__41_ ^ t_2__45_;
  assign t_3__40_ = t_2__40_ ^ t_2__44_;
  assign t_3__39_ = t_2__39_ ^ t_2__43_;
  assign t_3__38_ = t_2__38_ ^ t_2__42_;
  assign t_3__37_ = t_2__37_ ^ t_2__41_;
  assign t_3__36_ = t_2__36_ ^ t_2__40_;
  assign t_3__35_ = t_2__35_ ^ t_2__39_;
  assign t_3__34_ = t_2__34_ ^ t_2__38_;
  assign t_3__33_ = t_2__33_ ^ t_2__37_;
  assign t_3__32_ = t_2__32_ ^ t_2__36_;
  assign t_3__31_ = t_2__31_ ^ t_2__35_;
  assign t_3__30_ = t_2__30_ ^ t_2__34_;
  assign t_3__29_ = t_2__29_ ^ t_2__33_;
  assign t_3__28_ = t_2__28_ ^ t_2__32_;
  assign t_3__27_ = t_2__27_ ^ t_2__31_;
  assign t_3__26_ = t_2__26_ ^ t_2__30_;
  assign t_3__25_ = t_2__25_ ^ t_2__29_;
  assign t_3__24_ = t_2__24_ ^ t_2__28_;
  assign t_3__23_ = t_2__23_ ^ t_2__27_;
  assign t_3__22_ = t_2__22_ ^ t_2__26_;
  assign t_3__21_ = t_2__21_ ^ t_2__25_;
  assign t_3__20_ = t_2__20_ ^ t_2__24_;
  assign t_3__19_ = t_2__19_ ^ t_2__23_;
  assign t_3__18_ = t_2__18_ ^ t_2__22_;
  assign t_3__17_ = t_2__17_ ^ t_2__21_;
  assign t_3__16_ = t_2__16_ ^ t_2__20_;
  assign t_3__15_ = t_2__15_ ^ t_2__19_;
  assign t_3__14_ = t_2__14_ ^ t_2__18_;
  assign t_3__13_ = t_2__13_ ^ t_2__17_;
  assign t_3__12_ = t_2__12_ ^ t_2__16_;
  assign t_3__11_ = t_2__11_ ^ t_2__15_;
  assign t_3__10_ = t_2__10_ ^ t_2__14_;
  assign t_3__9_ = t_2__9_ ^ t_2__13_;
  assign t_3__8_ = t_2__8_ ^ t_2__12_;
  assign t_3__7_ = t_2__7_ ^ t_2__11_;
  assign t_3__6_ = t_2__6_ ^ t_2__10_;
  assign t_3__5_ = t_2__5_ ^ t_2__9_;
  assign t_3__4_ = t_2__4_ ^ t_2__8_;
  assign t_3__3_ = t_2__3_ ^ t_2__7_;
  assign t_3__2_ = t_2__2_ ^ t_2__6_;
  assign t_3__1_ = t_2__1_ ^ t_2__5_;
  assign t_3__0_ = t_2__0_ ^ t_2__4_;
  assign t_4__127_ = t_3__127_ ^ 1'b0;
  assign t_4__126_ = t_3__126_ ^ 1'b0;
  assign t_4__125_ = t_3__125_ ^ 1'b0;
  assign t_4__124_ = t_3__124_ ^ 1'b0;
  assign t_4__123_ = t_3__123_ ^ 1'b0;
  assign t_4__122_ = t_3__122_ ^ 1'b0;
  assign t_4__121_ = t_3__121_ ^ 1'b0;
  assign t_4__120_ = t_3__120_ ^ 1'b0;
  assign t_4__119_ = t_3__119_ ^ t_3__127_;
  assign t_4__118_ = t_3__118_ ^ t_3__126_;
  assign t_4__117_ = t_3__117_ ^ t_3__125_;
  assign t_4__116_ = t_3__116_ ^ t_3__124_;
  assign t_4__115_ = t_3__115_ ^ t_3__123_;
  assign t_4__114_ = t_3__114_ ^ t_3__122_;
  assign t_4__113_ = t_3__113_ ^ t_3__121_;
  assign t_4__112_ = t_3__112_ ^ t_3__120_;
  assign t_4__111_ = t_3__111_ ^ t_3__119_;
  assign t_4__110_ = t_3__110_ ^ t_3__118_;
  assign t_4__109_ = t_3__109_ ^ t_3__117_;
  assign t_4__108_ = t_3__108_ ^ t_3__116_;
  assign t_4__107_ = t_3__107_ ^ t_3__115_;
  assign t_4__106_ = t_3__106_ ^ t_3__114_;
  assign t_4__105_ = t_3__105_ ^ t_3__113_;
  assign t_4__104_ = t_3__104_ ^ t_3__112_;
  assign t_4__103_ = t_3__103_ ^ t_3__111_;
  assign t_4__102_ = t_3__102_ ^ t_3__110_;
  assign t_4__101_ = t_3__101_ ^ t_3__109_;
  assign t_4__100_ = t_3__100_ ^ t_3__108_;
  assign t_4__99_ = t_3__99_ ^ t_3__107_;
  assign t_4__98_ = t_3__98_ ^ t_3__106_;
  assign t_4__97_ = t_3__97_ ^ t_3__105_;
  assign t_4__96_ = t_3__96_ ^ t_3__104_;
  assign t_4__95_ = t_3__95_ ^ t_3__103_;
  assign t_4__94_ = t_3__94_ ^ t_3__102_;
  assign t_4__93_ = t_3__93_ ^ t_3__101_;
  assign t_4__92_ = t_3__92_ ^ t_3__100_;
  assign t_4__91_ = t_3__91_ ^ t_3__99_;
  assign t_4__90_ = t_3__90_ ^ t_3__98_;
  assign t_4__89_ = t_3__89_ ^ t_3__97_;
  assign t_4__88_ = t_3__88_ ^ t_3__96_;
  assign t_4__87_ = t_3__87_ ^ t_3__95_;
  assign t_4__86_ = t_3__86_ ^ t_3__94_;
  assign t_4__85_ = t_3__85_ ^ t_3__93_;
  assign t_4__84_ = t_3__84_ ^ t_3__92_;
  assign t_4__83_ = t_3__83_ ^ t_3__91_;
  assign t_4__82_ = t_3__82_ ^ t_3__90_;
  assign t_4__81_ = t_3__81_ ^ t_3__89_;
  assign t_4__80_ = t_3__80_ ^ t_3__88_;
  assign t_4__79_ = t_3__79_ ^ t_3__87_;
  assign t_4__78_ = t_3__78_ ^ t_3__86_;
  assign t_4__77_ = t_3__77_ ^ t_3__85_;
  assign t_4__76_ = t_3__76_ ^ t_3__84_;
  assign t_4__75_ = t_3__75_ ^ t_3__83_;
  assign t_4__74_ = t_3__74_ ^ t_3__82_;
  assign t_4__73_ = t_3__73_ ^ t_3__81_;
  assign t_4__72_ = t_3__72_ ^ t_3__80_;
  assign t_4__71_ = t_3__71_ ^ t_3__79_;
  assign t_4__70_ = t_3__70_ ^ t_3__78_;
  assign t_4__69_ = t_3__69_ ^ t_3__77_;
  assign t_4__68_ = t_3__68_ ^ t_3__76_;
  assign t_4__67_ = t_3__67_ ^ t_3__75_;
  assign t_4__66_ = t_3__66_ ^ t_3__74_;
  assign t_4__65_ = t_3__65_ ^ t_3__73_;
  assign t_4__64_ = t_3__64_ ^ t_3__72_;
  assign t_4__63_ = t_3__63_ ^ t_3__71_;
  assign t_4__62_ = t_3__62_ ^ t_3__70_;
  assign t_4__61_ = t_3__61_ ^ t_3__69_;
  assign t_4__60_ = t_3__60_ ^ t_3__68_;
  assign t_4__59_ = t_3__59_ ^ t_3__67_;
  assign t_4__58_ = t_3__58_ ^ t_3__66_;
  assign t_4__57_ = t_3__57_ ^ t_3__65_;
  assign t_4__56_ = t_3__56_ ^ t_3__64_;
  assign t_4__55_ = t_3__55_ ^ t_3__63_;
  assign t_4__54_ = t_3__54_ ^ t_3__62_;
  assign t_4__53_ = t_3__53_ ^ t_3__61_;
  assign t_4__52_ = t_3__52_ ^ t_3__60_;
  assign t_4__51_ = t_3__51_ ^ t_3__59_;
  assign t_4__50_ = t_3__50_ ^ t_3__58_;
  assign t_4__49_ = t_3__49_ ^ t_3__57_;
  assign t_4__48_ = t_3__48_ ^ t_3__56_;
  assign t_4__47_ = t_3__47_ ^ t_3__55_;
  assign t_4__46_ = t_3__46_ ^ t_3__54_;
  assign t_4__45_ = t_3__45_ ^ t_3__53_;
  assign t_4__44_ = t_3__44_ ^ t_3__52_;
  assign t_4__43_ = t_3__43_ ^ t_3__51_;
  assign t_4__42_ = t_3__42_ ^ t_3__50_;
  assign t_4__41_ = t_3__41_ ^ t_3__49_;
  assign t_4__40_ = t_3__40_ ^ t_3__48_;
  assign t_4__39_ = t_3__39_ ^ t_3__47_;
  assign t_4__38_ = t_3__38_ ^ t_3__46_;
  assign t_4__37_ = t_3__37_ ^ t_3__45_;
  assign t_4__36_ = t_3__36_ ^ t_3__44_;
  assign t_4__35_ = t_3__35_ ^ t_3__43_;
  assign t_4__34_ = t_3__34_ ^ t_3__42_;
  assign t_4__33_ = t_3__33_ ^ t_3__41_;
  assign t_4__32_ = t_3__32_ ^ t_3__40_;
  assign t_4__31_ = t_3__31_ ^ t_3__39_;
  assign t_4__30_ = t_3__30_ ^ t_3__38_;
  assign t_4__29_ = t_3__29_ ^ t_3__37_;
  assign t_4__28_ = t_3__28_ ^ t_3__36_;
  assign t_4__27_ = t_3__27_ ^ t_3__35_;
  assign t_4__26_ = t_3__26_ ^ t_3__34_;
  assign t_4__25_ = t_3__25_ ^ t_3__33_;
  assign t_4__24_ = t_3__24_ ^ t_3__32_;
  assign t_4__23_ = t_3__23_ ^ t_3__31_;
  assign t_4__22_ = t_3__22_ ^ t_3__30_;
  assign t_4__21_ = t_3__21_ ^ t_3__29_;
  assign t_4__20_ = t_3__20_ ^ t_3__28_;
  assign t_4__19_ = t_3__19_ ^ t_3__27_;
  assign t_4__18_ = t_3__18_ ^ t_3__26_;
  assign t_4__17_ = t_3__17_ ^ t_3__25_;
  assign t_4__16_ = t_3__16_ ^ t_3__24_;
  assign t_4__15_ = t_3__15_ ^ t_3__23_;
  assign t_4__14_ = t_3__14_ ^ t_3__22_;
  assign t_4__13_ = t_3__13_ ^ t_3__21_;
  assign t_4__12_ = t_3__12_ ^ t_3__20_;
  assign t_4__11_ = t_3__11_ ^ t_3__19_;
  assign t_4__10_ = t_3__10_ ^ t_3__18_;
  assign t_4__9_ = t_3__9_ ^ t_3__17_;
  assign t_4__8_ = t_3__8_ ^ t_3__16_;
  assign t_4__7_ = t_3__7_ ^ t_3__15_;
  assign t_4__6_ = t_3__6_ ^ t_3__14_;
  assign t_4__5_ = t_3__5_ ^ t_3__13_;
  assign t_4__4_ = t_3__4_ ^ t_3__12_;
  assign t_4__3_ = t_3__3_ ^ t_3__11_;
  assign t_4__2_ = t_3__2_ ^ t_3__10_;
  assign t_4__1_ = t_3__1_ ^ t_3__9_;
  assign t_4__0_ = t_3__0_ ^ t_3__8_;
  assign t_5__127_ = t_4__127_ ^ 1'b0;
  assign t_5__126_ = t_4__126_ ^ 1'b0;
  assign t_5__125_ = t_4__125_ ^ 1'b0;
  assign t_5__124_ = t_4__124_ ^ 1'b0;
  assign t_5__123_ = t_4__123_ ^ 1'b0;
  assign t_5__122_ = t_4__122_ ^ 1'b0;
  assign t_5__121_ = t_4__121_ ^ 1'b0;
  assign t_5__120_ = t_4__120_ ^ 1'b0;
  assign t_5__119_ = t_4__119_ ^ 1'b0;
  assign t_5__118_ = t_4__118_ ^ 1'b0;
  assign t_5__117_ = t_4__117_ ^ 1'b0;
  assign t_5__116_ = t_4__116_ ^ 1'b0;
  assign t_5__115_ = t_4__115_ ^ 1'b0;
  assign t_5__114_ = t_4__114_ ^ 1'b0;
  assign t_5__113_ = t_4__113_ ^ 1'b0;
  assign t_5__112_ = t_4__112_ ^ 1'b0;
  assign t_5__111_ = t_4__111_ ^ t_4__127_;
  assign t_5__110_ = t_4__110_ ^ t_4__126_;
  assign t_5__109_ = t_4__109_ ^ t_4__125_;
  assign t_5__108_ = t_4__108_ ^ t_4__124_;
  assign t_5__107_ = t_4__107_ ^ t_4__123_;
  assign t_5__106_ = t_4__106_ ^ t_4__122_;
  assign t_5__105_ = t_4__105_ ^ t_4__121_;
  assign t_5__104_ = t_4__104_ ^ t_4__120_;
  assign t_5__103_ = t_4__103_ ^ t_4__119_;
  assign t_5__102_ = t_4__102_ ^ t_4__118_;
  assign t_5__101_ = t_4__101_ ^ t_4__117_;
  assign t_5__100_ = t_4__100_ ^ t_4__116_;
  assign t_5__99_ = t_4__99_ ^ t_4__115_;
  assign t_5__98_ = t_4__98_ ^ t_4__114_;
  assign t_5__97_ = t_4__97_ ^ t_4__113_;
  assign t_5__96_ = t_4__96_ ^ t_4__112_;
  assign t_5__95_ = t_4__95_ ^ t_4__111_;
  assign t_5__94_ = t_4__94_ ^ t_4__110_;
  assign t_5__93_ = t_4__93_ ^ t_4__109_;
  assign t_5__92_ = t_4__92_ ^ t_4__108_;
  assign t_5__91_ = t_4__91_ ^ t_4__107_;
  assign t_5__90_ = t_4__90_ ^ t_4__106_;
  assign t_5__89_ = t_4__89_ ^ t_4__105_;
  assign t_5__88_ = t_4__88_ ^ t_4__104_;
  assign t_5__87_ = t_4__87_ ^ t_4__103_;
  assign t_5__86_ = t_4__86_ ^ t_4__102_;
  assign t_5__85_ = t_4__85_ ^ t_4__101_;
  assign t_5__84_ = t_4__84_ ^ t_4__100_;
  assign t_5__83_ = t_4__83_ ^ t_4__99_;
  assign t_5__82_ = t_4__82_ ^ t_4__98_;
  assign t_5__81_ = t_4__81_ ^ t_4__97_;
  assign t_5__80_ = t_4__80_ ^ t_4__96_;
  assign t_5__79_ = t_4__79_ ^ t_4__95_;
  assign t_5__78_ = t_4__78_ ^ t_4__94_;
  assign t_5__77_ = t_4__77_ ^ t_4__93_;
  assign t_5__76_ = t_4__76_ ^ t_4__92_;
  assign t_5__75_ = t_4__75_ ^ t_4__91_;
  assign t_5__74_ = t_4__74_ ^ t_4__90_;
  assign t_5__73_ = t_4__73_ ^ t_4__89_;
  assign t_5__72_ = t_4__72_ ^ t_4__88_;
  assign t_5__71_ = t_4__71_ ^ t_4__87_;
  assign t_5__70_ = t_4__70_ ^ t_4__86_;
  assign t_5__69_ = t_4__69_ ^ t_4__85_;
  assign t_5__68_ = t_4__68_ ^ t_4__84_;
  assign t_5__67_ = t_4__67_ ^ t_4__83_;
  assign t_5__66_ = t_4__66_ ^ t_4__82_;
  assign t_5__65_ = t_4__65_ ^ t_4__81_;
  assign t_5__64_ = t_4__64_ ^ t_4__80_;
  assign t_5__63_ = t_4__63_ ^ t_4__79_;
  assign t_5__62_ = t_4__62_ ^ t_4__78_;
  assign t_5__61_ = t_4__61_ ^ t_4__77_;
  assign t_5__60_ = t_4__60_ ^ t_4__76_;
  assign t_5__59_ = t_4__59_ ^ t_4__75_;
  assign t_5__58_ = t_4__58_ ^ t_4__74_;
  assign t_5__57_ = t_4__57_ ^ t_4__73_;
  assign t_5__56_ = t_4__56_ ^ t_4__72_;
  assign t_5__55_ = t_4__55_ ^ t_4__71_;
  assign t_5__54_ = t_4__54_ ^ t_4__70_;
  assign t_5__53_ = t_4__53_ ^ t_4__69_;
  assign t_5__52_ = t_4__52_ ^ t_4__68_;
  assign t_5__51_ = t_4__51_ ^ t_4__67_;
  assign t_5__50_ = t_4__50_ ^ t_4__66_;
  assign t_5__49_ = t_4__49_ ^ t_4__65_;
  assign t_5__48_ = t_4__48_ ^ t_4__64_;
  assign t_5__47_ = t_4__47_ ^ t_4__63_;
  assign t_5__46_ = t_4__46_ ^ t_4__62_;
  assign t_5__45_ = t_4__45_ ^ t_4__61_;
  assign t_5__44_ = t_4__44_ ^ t_4__60_;
  assign t_5__43_ = t_4__43_ ^ t_4__59_;
  assign t_5__42_ = t_4__42_ ^ t_4__58_;
  assign t_5__41_ = t_4__41_ ^ t_4__57_;
  assign t_5__40_ = t_4__40_ ^ t_4__56_;
  assign t_5__39_ = t_4__39_ ^ t_4__55_;
  assign t_5__38_ = t_4__38_ ^ t_4__54_;
  assign t_5__37_ = t_4__37_ ^ t_4__53_;
  assign t_5__36_ = t_4__36_ ^ t_4__52_;
  assign t_5__35_ = t_4__35_ ^ t_4__51_;
  assign t_5__34_ = t_4__34_ ^ t_4__50_;
  assign t_5__33_ = t_4__33_ ^ t_4__49_;
  assign t_5__32_ = t_4__32_ ^ t_4__48_;
  assign t_5__31_ = t_4__31_ ^ t_4__47_;
  assign t_5__30_ = t_4__30_ ^ t_4__46_;
  assign t_5__29_ = t_4__29_ ^ t_4__45_;
  assign t_5__28_ = t_4__28_ ^ t_4__44_;
  assign t_5__27_ = t_4__27_ ^ t_4__43_;
  assign t_5__26_ = t_4__26_ ^ t_4__42_;
  assign t_5__25_ = t_4__25_ ^ t_4__41_;
  assign t_5__24_ = t_4__24_ ^ t_4__40_;
  assign t_5__23_ = t_4__23_ ^ t_4__39_;
  assign t_5__22_ = t_4__22_ ^ t_4__38_;
  assign t_5__21_ = t_4__21_ ^ t_4__37_;
  assign t_5__20_ = t_4__20_ ^ t_4__36_;
  assign t_5__19_ = t_4__19_ ^ t_4__35_;
  assign t_5__18_ = t_4__18_ ^ t_4__34_;
  assign t_5__17_ = t_4__17_ ^ t_4__33_;
  assign t_5__16_ = t_4__16_ ^ t_4__32_;
  assign t_5__15_ = t_4__15_ ^ t_4__31_;
  assign t_5__14_ = t_4__14_ ^ t_4__30_;
  assign t_5__13_ = t_4__13_ ^ t_4__29_;
  assign t_5__12_ = t_4__12_ ^ t_4__28_;
  assign t_5__11_ = t_4__11_ ^ t_4__27_;
  assign t_5__10_ = t_4__10_ ^ t_4__26_;
  assign t_5__9_ = t_4__9_ ^ t_4__25_;
  assign t_5__8_ = t_4__8_ ^ t_4__24_;
  assign t_5__7_ = t_4__7_ ^ t_4__23_;
  assign t_5__6_ = t_4__6_ ^ t_4__22_;
  assign t_5__5_ = t_4__5_ ^ t_4__21_;
  assign t_5__4_ = t_4__4_ ^ t_4__20_;
  assign t_5__3_ = t_4__3_ ^ t_4__19_;
  assign t_5__2_ = t_4__2_ ^ t_4__18_;
  assign t_5__1_ = t_4__1_ ^ t_4__17_;
  assign t_5__0_ = t_4__0_ ^ t_4__16_;
  assign t_6__127_ = t_5__127_ ^ 1'b0;
  assign t_6__126_ = t_5__126_ ^ 1'b0;
  assign t_6__125_ = t_5__125_ ^ 1'b0;
  assign t_6__124_ = t_5__124_ ^ 1'b0;
  assign t_6__123_ = t_5__123_ ^ 1'b0;
  assign t_6__122_ = t_5__122_ ^ 1'b0;
  assign t_6__121_ = t_5__121_ ^ 1'b0;
  assign t_6__120_ = t_5__120_ ^ 1'b0;
  assign t_6__119_ = t_5__119_ ^ 1'b0;
  assign t_6__118_ = t_5__118_ ^ 1'b0;
  assign t_6__117_ = t_5__117_ ^ 1'b0;
  assign t_6__116_ = t_5__116_ ^ 1'b0;
  assign t_6__115_ = t_5__115_ ^ 1'b0;
  assign t_6__114_ = t_5__114_ ^ 1'b0;
  assign t_6__113_ = t_5__113_ ^ 1'b0;
  assign t_6__112_ = t_5__112_ ^ 1'b0;
  assign t_6__111_ = t_5__111_ ^ 1'b0;
  assign t_6__110_ = t_5__110_ ^ 1'b0;
  assign t_6__109_ = t_5__109_ ^ 1'b0;
  assign t_6__108_ = t_5__108_ ^ 1'b0;
  assign t_6__107_ = t_5__107_ ^ 1'b0;
  assign t_6__106_ = t_5__106_ ^ 1'b0;
  assign t_6__105_ = t_5__105_ ^ 1'b0;
  assign t_6__104_ = t_5__104_ ^ 1'b0;
  assign t_6__103_ = t_5__103_ ^ 1'b0;
  assign t_6__102_ = t_5__102_ ^ 1'b0;
  assign t_6__101_ = t_5__101_ ^ 1'b0;
  assign t_6__100_ = t_5__100_ ^ 1'b0;
  assign t_6__99_ = t_5__99_ ^ 1'b0;
  assign t_6__98_ = t_5__98_ ^ 1'b0;
  assign t_6__97_ = t_5__97_ ^ 1'b0;
  assign t_6__96_ = t_5__96_ ^ 1'b0;
  assign t_6__95_ = t_5__95_ ^ t_5__127_;
  assign t_6__94_ = t_5__94_ ^ t_5__126_;
  assign t_6__93_ = t_5__93_ ^ t_5__125_;
  assign t_6__92_ = t_5__92_ ^ t_5__124_;
  assign t_6__91_ = t_5__91_ ^ t_5__123_;
  assign t_6__90_ = t_5__90_ ^ t_5__122_;
  assign t_6__89_ = t_5__89_ ^ t_5__121_;
  assign t_6__88_ = t_5__88_ ^ t_5__120_;
  assign t_6__87_ = t_5__87_ ^ t_5__119_;
  assign t_6__86_ = t_5__86_ ^ t_5__118_;
  assign t_6__85_ = t_5__85_ ^ t_5__117_;
  assign t_6__84_ = t_5__84_ ^ t_5__116_;
  assign t_6__83_ = t_5__83_ ^ t_5__115_;
  assign t_6__82_ = t_5__82_ ^ t_5__114_;
  assign t_6__81_ = t_5__81_ ^ t_5__113_;
  assign t_6__80_ = t_5__80_ ^ t_5__112_;
  assign t_6__79_ = t_5__79_ ^ t_5__111_;
  assign t_6__78_ = t_5__78_ ^ t_5__110_;
  assign t_6__77_ = t_5__77_ ^ t_5__109_;
  assign t_6__76_ = t_5__76_ ^ t_5__108_;
  assign t_6__75_ = t_5__75_ ^ t_5__107_;
  assign t_6__74_ = t_5__74_ ^ t_5__106_;
  assign t_6__73_ = t_5__73_ ^ t_5__105_;
  assign t_6__72_ = t_5__72_ ^ t_5__104_;
  assign t_6__71_ = t_5__71_ ^ t_5__103_;
  assign t_6__70_ = t_5__70_ ^ t_5__102_;
  assign t_6__69_ = t_5__69_ ^ t_5__101_;
  assign t_6__68_ = t_5__68_ ^ t_5__100_;
  assign t_6__67_ = t_5__67_ ^ t_5__99_;
  assign t_6__66_ = t_5__66_ ^ t_5__98_;
  assign t_6__65_ = t_5__65_ ^ t_5__97_;
  assign t_6__64_ = t_5__64_ ^ t_5__96_;
  assign t_6__63_ = t_5__63_ ^ t_5__95_;
  assign t_6__62_ = t_5__62_ ^ t_5__94_;
  assign t_6__61_ = t_5__61_ ^ t_5__93_;
  assign t_6__60_ = t_5__60_ ^ t_5__92_;
  assign t_6__59_ = t_5__59_ ^ t_5__91_;
  assign t_6__58_ = t_5__58_ ^ t_5__90_;
  assign t_6__57_ = t_5__57_ ^ t_5__89_;
  assign t_6__56_ = t_5__56_ ^ t_5__88_;
  assign t_6__55_ = t_5__55_ ^ t_5__87_;
  assign t_6__54_ = t_5__54_ ^ t_5__86_;
  assign t_6__53_ = t_5__53_ ^ t_5__85_;
  assign t_6__52_ = t_5__52_ ^ t_5__84_;
  assign t_6__51_ = t_5__51_ ^ t_5__83_;
  assign t_6__50_ = t_5__50_ ^ t_5__82_;
  assign t_6__49_ = t_5__49_ ^ t_5__81_;
  assign t_6__48_ = t_5__48_ ^ t_5__80_;
  assign t_6__47_ = t_5__47_ ^ t_5__79_;
  assign t_6__46_ = t_5__46_ ^ t_5__78_;
  assign t_6__45_ = t_5__45_ ^ t_5__77_;
  assign t_6__44_ = t_5__44_ ^ t_5__76_;
  assign t_6__43_ = t_5__43_ ^ t_5__75_;
  assign t_6__42_ = t_5__42_ ^ t_5__74_;
  assign t_6__41_ = t_5__41_ ^ t_5__73_;
  assign t_6__40_ = t_5__40_ ^ t_5__72_;
  assign t_6__39_ = t_5__39_ ^ t_5__71_;
  assign t_6__38_ = t_5__38_ ^ t_5__70_;
  assign t_6__37_ = t_5__37_ ^ t_5__69_;
  assign t_6__36_ = t_5__36_ ^ t_5__68_;
  assign t_6__35_ = t_5__35_ ^ t_5__67_;
  assign t_6__34_ = t_5__34_ ^ t_5__66_;
  assign t_6__33_ = t_5__33_ ^ t_5__65_;
  assign t_6__32_ = t_5__32_ ^ t_5__64_;
  assign t_6__31_ = t_5__31_ ^ t_5__63_;
  assign t_6__30_ = t_5__30_ ^ t_5__62_;
  assign t_6__29_ = t_5__29_ ^ t_5__61_;
  assign t_6__28_ = t_5__28_ ^ t_5__60_;
  assign t_6__27_ = t_5__27_ ^ t_5__59_;
  assign t_6__26_ = t_5__26_ ^ t_5__58_;
  assign t_6__25_ = t_5__25_ ^ t_5__57_;
  assign t_6__24_ = t_5__24_ ^ t_5__56_;
  assign t_6__23_ = t_5__23_ ^ t_5__55_;
  assign t_6__22_ = t_5__22_ ^ t_5__54_;
  assign t_6__21_ = t_5__21_ ^ t_5__53_;
  assign t_6__20_ = t_5__20_ ^ t_5__52_;
  assign t_6__19_ = t_5__19_ ^ t_5__51_;
  assign t_6__18_ = t_5__18_ ^ t_5__50_;
  assign t_6__17_ = t_5__17_ ^ t_5__49_;
  assign t_6__16_ = t_5__16_ ^ t_5__48_;
  assign t_6__15_ = t_5__15_ ^ t_5__47_;
  assign t_6__14_ = t_5__14_ ^ t_5__46_;
  assign t_6__13_ = t_5__13_ ^ t_5__45_;
  assign t_6__12_ = t_5__12_ ^ t_5__44_;
  assign t_6__11_ = t_5__11_ ^ t_5__43_;
  assign t_6__10_ = t_5__10_ ^ t_5__42_;
  assign t_6__9_ = t_5__9_ ^ t_5__41_;
  assign t_6__8_ = t_5__8_ ^ t_5__40_;
  assign t_6__7_ = t_5__7_ ^ t_5__39_;
  assign t_6__6_ = t_5__6_ ^ t_5__38_;
  assign t_6__5_ = t_5__5_ ^ t_5__37_;
  assign t_6__4_ = t_5__4_ ^ t_5__36_;
  assign t_6__3_ = t_5__3_ ^ t_5__35_;
  assign t_6__2_ = t_5__2_ ^ t_5__34_;
  assign t_6__1_ = t_5__1_ ^ t_5__33_;
  assign t_6__0_ = t_5__0_ ^ t_5__32_;
  assign o[127] = t_6__127_ ^ 1'b0;
  assign o[126] = t_6__126_ ^ 1'b0;
  assign o[125] = t_6__125_ ^ 1'b0;
  assign o[124] = t_6__124_ ^ 1'b0;
  assign o[123] = t_6__123_ ^ 1'b0;
  assign o[122] = t_6__122_ ^ 1'b0;
  assign o[121] = t_6__121_ ^ 1'b0;
  assign o[120] = t_6__120_ ^ 1'b0;
  assign o[119] = t_6__119_ ^ 1'b0;
  assign o[118] = t_6__118_ ^ 1'b0;
  assign o[117] = t_6__117_ ^ 1'b0;
  assign o[116] = t_6__116_ ^ 1'b0;
  assign o[115] = t_6__115_ ^ 1'b0;
  assign o[114] = t_6__114_ ^ 1'b0;
  assign o[113] = t_6__113_ ^ 1'b0;
  assign o[112] = t_6__112_ ^ 1'b0;
  assign o[111] = t_6__111_ ^ 1'b0;
  assign o[110] = t_6__110_ ^ 1'b0;
  assign o[109] = t_6__109_ ^ 1'b0;
  assign o[108] = t_6__108_ ^ 1'b0;
  assign o[107] = t_6__107_ ^ 1'b0;
  assign o[106] = t_6__106_ ^ 1'b0;
  assign o[105] = t_6__105_ ^ 1'b0;
  assign o[104] = t_6__104_ ^ 1'b0;
  assign o[103] = t_6__103_ ^ 1'b0;
  assign o[102] = t_6__102_ ^ 1'b0;
  assign o[101] = t_6__101_ ^ 1'b0;
  assign o[100] = t_6__100_ ^ 1'b0;
  assign o[99] = t_6__99_ ^ 1'b0;
  assign o[98] = t_6__98_ ^ 1'b0;
  assign o[97] = t_6__97_ ^ 1'b0;
  assign o[96] = t_6__96_ ^ 1'b0;
  assign o[95] = t_6__95_ ^ 1'b0;
  assign o[94] = t_6__94_ ^ 1'b0;
  assign o[93] = t_6__93_ ^ 1'b0;
  assign o[92] = t_6__92_ ^ 1'b0;
  assign o[91] = t_6__91_ ^ 1'b0;
  assign o[90] = t_6__90_ ^ 1'b0;
  assign o[89] = t_6__89_ ^ 1'b0;
  assign o[88] = t_6__88_ ^ 1'b0;
  assign o[87] = t_6__87_ ^ 1'b0;
  assign o[86] = t_6__86_ ^ 1'b0;
  assign o[85] = t_6__85_ ^ 1'b0;
  assign o[84] = t_6__84_ ^ 1'b0;
  assign o[83] = t_6__83_ ^ 1'b0;
  assign o[82] = t_6__82_ ^ 1'b0;
  assign o[81] = t_6__81_ ^ 1'b0;
  assign o[80] = t_6__80_ ^ 1'b0;
  assign o[79] = t_6__79_ ^ 1'b0;
  assign o[78] = t_6__78_ ^ 1'b0;
  assign o[77] = t_6__77_ ^ 1'b0;
  assign o[76] = t_6__76_ ^ 1'b0;
  assign o[75] = t_6__75_ ^ 1'b0;
  assign o[74] = t_6__74_ ^ 1'b0;
  assign o[73] = t_6__73_ ^ 1'b0;
  assign o[72] = t_6__72_ ^ 1'b0;
  assign o[71] = t_6__71_ ^ 1'b0;
  assign o[70] = t_6__70_ ^ 1'b0;
  assign o[69] = t_6__69_ ^ 1'b0;
  assign o[68] = t_6__68_ ^ 1'b0;
  assign o[67] = t_6__67_ ^ 1'b0;
  assign o[66] = t_6__66_ ^ 1'b0;
  assign o[65] = t_6__65_ ^ 1'b0;
  assign o[64] = t_6__64_ ^ 1'b0;
  assign o[63] = t_6__63_ ^ t_6__127_;
  assign o[62] = t_6__62_ ^ t_6__126_;
  assign o[61] = t_6__61_ ^ t_6__125_;
  assign o[60] = t_6__60_ ^ t_6__124_;
  assign o[59] = t_6__59_ ^ t_6__123_;
  assign o[58] = t_6__58_ ^ t_6__122_;
  assign o[57] = t_6__57_ ^ t_6__121_;
  assign o[56] = t_6__56_ ^ t_6__120_;
  assign o[55] = t_6__55_ ^ t_6__119_;
  assign o[54] = t_6__54_ ^ t_6__118_;
  assign o[53] = t_6__53_ ^ t_6__117_;
  assign o[52] = t_6__52_ ^ t_6__116_;
  assign o[51] = t_6__51_ ^ t_6__115_;
  assign o[50] = t_6__50_ ^ t_6__114_;
  assign o[49] = t_6__49_ ^ t_6__113_;
  assign o[48] = t_6__48_ ^ t_6__112_;
  assign o[47] = t_6__47_ ^ t_6__111_;
  assign o[46] = t_6__46_ ^ t_6__110_;
  assign o[45] = t_6__45_ ^ t_6__109_;
  assign o[44] = t_6__44_ ^ t_6__108_;
  assign o[43] = t_6__43_ ^ t_6__107_;
  assign o[42] = t_6__42_ ^ t_6__106_;
  assign o[41] = t_6__41_ ^ t_6__105_;
  assign o[40] = t_6__40_ ^ t_6__104_;
  assign o[39] = t_6__39_ ^ t_6__103_;
  assign o[38] = t_6__38_ ^ t_6__102_;
  assign o[37] = t_6__37_ ^ t_6__101_;
  assign o[36] = t_6__36_ ^ t_6__100_;
  assign o[35] = t_6__35_ ^ t_6__99_;
  assign o[34] = t_6__34_ ^ t_6__98_;
  assign o[33] = t_6__33_ ^ t_6__97_;
  assign o[32] = t_6__32_ ^ t_6__96_;
  assign o[31] = t_6__31_ ^ t_6__95_;
  assign o[30] = t_6__30_ ^ t_6__94_;
  assign o[29] = t_6__29_ ^ t_6__93_;
  assign o[28] = t_6__28_ ^ t_6__92_;
  assign o[27] = t_6__27_ ^ t_6__91_;
  assign o[26] = t_6__26_ ^ t_6__90_;
  assign o[25] = t_6__25_ ^ t_6__89_;
  assign o[24] = t_6__24_ ^ t_6__88_;
  assign o[23] = t_6__23_ ^ t_6__87_;
  assign o[22] = t_6__22_ ^ t_6__86_;
  assign o[21] = t_6__21_ ^ t_6__85_;
  assign o[20] = t_6__20_ ^ t_6__84_;
  assign o[19] = t_6__19_ ^ t_6__83_;
  assign o[18] = t_6__18_ ^ t_6__82_;
  assign o[17] = t_6__17_ ^ t_6__81_;
  assign o[16] = t_6__16_ ^ t_6__80_;
  assign o[15] = t_6__15_ ^ t_6__79_;
  assign o[14] = t_6__14_ ^ t_6__78_;
  assign o[13] = t_6__13_ ^ t_6__77_;
  assign o[12] = t_6__12_ ^ t_6__76_;
  assign o[11] = t_6__11_ ^ t_6__75_;
  assign o[10] = t_6__10_ ^ t_6__74_;
  assign o[9] = t_6__9_ ^ t_6__73_;
  assign o[8] = t_6__8_ ^ t_6__72_;
  assign o[7] = t_6__7_ ^ t_6__71_;
  assign o[6] = t_6__6_ ^ t_6__70_;
  assign o[5] = t_6__5_ ^ t_6__69_;
  assign o[4] = t_6__4_ ^ t_6__68_;
  assign o[3] = t_6__3_ ^ t_6__67_;
  assign o[2] = t_6__2_ ^ t_6__66_;
  assign o[1] = t_6__1_ ^ t_6__65_;
  assign o[0] = t_6__0_ ^ t_6__64_;

endmodule



module bsg_gray_to_binary
(
  gray_i,
  binary_o
);

  input [127:0] gray_i;
  output [127:0] binary_o;
  wire [127:0] binary_o;

  bsg_scan_width_p128_xor_p1
  scan_xor
  (
    .i(gray_i),
    .o(binary_o)
  );


endmodule

