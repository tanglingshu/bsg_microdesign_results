

module top
(
  clk_i,
  reset_i,
  en_i,
  w_v_i,
  w_set_not_clear_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_data_i,
  r_v_o,
  r_addr_o,
  empty_v_o,
  empty_addr_o
);

  input [9:0] w_addr_i;
  input [31:0] w_data_i;
  input [31:0] r_data_i;
  output [9:0] r_addr_o;
  output [9:0] empty_addr_o;
  input clk_i;
  input reset_i;
  input en_i;
  input w_v_i;
  input w_set_not_clear_i;
  input r_v_i;
  output r_v_o;
  output empty_v_o;

  bsg_cam_1r1w
  wrapper
  (
    .w_addr_i(w_addr_i),
    .w_data_i(w_data_i),
    .r_data_i(r_data_i),
    .r_addr_o(r_addr_o),
    .empty_addr_o(empty_addr_o),
    .clk_i(clk_i),
    .reset_i(reset_i),
    .en_i(en_i),
    .w_v_i(w_v_i),
    .w_set_not_clear_i(w_set_not_clear_i),
    .r_v_i(r_v_i),
    .r_v_o(r_v_o),
    .empty_v_o(empty_v_o)
  );


endmodule



module bsg_scan_width_p1024_or_p1_lo_to_hi_p1
(
  i,
  o
);

  input [1023:0] i;
  output [1023:0] o;
  wire [1023:0] o;
  wire t_1__1023_,t_1__1022_,t_1__1021_,t_1__1020_,t_1__1019_,t_1__1018_,t_1__1017_,
  t_1__1016_,t_1__1015_,t_1__1014_,t_1__1013_,t_1__1012_,t_1__1011_,t_1__1010_,
  t_1__1009_,t_1__1008_,t_1__1007_,t_1__1006_,t_1__1005_,t_1__1004_,t_1__1003_,
  t_1__1002_,t_1__1001_,t_1__1000_,t_1__999_,t_1__998_,t_1__997_,t_1__996_,t_1__995_,
  t_1__994_,t_1__993_,t_1__992_,t_1__991_,t_1__990_,t_1__989_,t_1__988_,t_1__987_,
  t_1__986_,t_1__985_,t_1__984_,t_1__983_,t_1__982_,t_1__981_,t_1__980_,t_1__979_,
  t_1__978_,t_1__977_,t_1__976_,t_1__975_,t_1__974_,t_1__973_,t_1__972_,t_1__971_,
  t_1__970_,t_1__969_,t_1__968_,t_1__967_,t_1__966_,t_1__965_,t_1__964_,t_1__963_,
  t_1__962_,t_1__961_,t_1__960_,t_1__959_,t_1__958_,t_1__957_,t_1__956_,t_1__955_,
  t_1__954_,t_1__953_,t_1__952_,t_1__951_,t_1__950_,t_1__949_,t_1__948_,t_1__947_,
  t_1__946_,t_1__945_,t_1__944_,t_1__943_,t_1__942_,t_1__941_,t_1__940_,t_1__939_,
  t_1__938_,t_1__937_,t_1__936_,t_1__935_,t_1__934_,t_1__933_,t_1__932_,t_1__931_,
  t_1__930_,t_1__929_,t_1__928_,t_1__927_,t_1__926_,t_1__925_,t_1__924_,t_1__923_,
  t_1__922_,t_1__921_,t_1__920_,t_1__919_,t_1__918_,t_1__917_,t_1__916_,t_1__915_,
  t_1__914_,t_1__913_,t_1__912_,t_1__911_,t_1__910_,t_1__909_,t_1__908_,t_1__907_,
  t_1__906_,t_1__905_,t_1__904_,t_1__903_,t_1__902_,t_1__901_,t_1__900_,t_1__899_,
  t_1__898_,t_1__897_,t_1__896_,t_1__895_,t_1__894_,t_1__893_,t_1__892_,t_1__891_,
  t_1__890_,t_1__889_,t_1__888_,t_1__887_,t_1__886_,t_1__885_,t_1__884_,t_1__883_,
  t_1__882_,t_1__881_,t_1__880_,t_1__879_,t_1__878_,t_1__877_,t_1__876_,t_1__875_,
  t_1__874_,t_1__873_,t_1__872_,t_1__871_,t_1__870_,t_1__869_,t_1__868_,t_1__867_,
  t_1__866_,t_1__865_,t_1__864_,t_1__863_,t_1__862_,t_1__861_,t_1__860_,t_1__859_,
  t_1__858_,t_1__857_,t_1__856_,t_1__855_,t_1__854_,t_1__853_,t_1__852_,t_1__851_,
  t_1__850_,t_1__849_,t_1__848_,t_1__847_,t_1__846_,t_1__845_,t_1__844_,t_1__843_,
  t_1__842_,t_1__841_,t_1__840_,t_1__839_,t_1__838_,t_1__837_,t_1__836_,t_1__835_,
  t_1__834_,t_1__833_,t_1__832_,t_1__831_,t_1__830_,t_1__829_,t_1__828_,t_1__827_,
  t_1__826_,t_1__825_,t_1__824_,t_1__823_,t_1__822_,t_1__821_,t_1__820_,t_1__819_,
  t_1__818_,t_1__817_,t_1__816_,t_1__815_,t_1__814_,t_1__813_,t_1__812_,t_1__811_,
  t_1__810_,t_1__809_,t_1__808_,t_1__807_,t_1__806_,t_1__805_,t_1__804_,t_1__803_,
  t_1__802_,t_1__801_,t_1__800_,t_1__799_,t_1__798_,t_1__797_,t_1__796_,t_1__795_,
  t_1__794_,t_1__793_,t_1__792_,t_1__791_,t_1__790_,t_1__789_,t_1__788_,t_1__787_,
  t_1__786_,t_1__785_,t_1__784_,t_1__783_,t_1__782_,t_1__781_,t_1__780_,t_1__779_,
  t_1__778_,t_1__777_,t_1__776_,t_1__775_,t_1__774_,t_1__773_,t_1__772_,t_1__771_,
  t_1__770_,t_1__769_,t_1__768_,t_1__767_,t_1__766_,t_1__765_,t_1__764_,t_1__763_,
  t_1__762_,t_1__761_,t_1__760_,t_1__759_,t_1__758_,t_1__757_,t_1__756_,t_1__755_,
  t_1__754_,t_1__753_,t_1__752_,t_1__751_,t_1__750_,t_1__749_,t_1__748_,t_1__747_,
  t_1__746_,t_1__745_,t_1__744_,t_1__743_,t_1__742_,t_1__741_,t_1__740_,t_1__739_,
  t_1__738_,t_1__737_,t_1__736_,t_1__735_,t_1__734_,t_1__733_,t_1__732_,t_1__731_,
  t_1__730_,t_1__729_,t_1__728_,t_1__727_,t_1__726_,t_1__725_,t_1__724_,t_1__723_,
  t_1__722_,t_1__721_,t_1__720_,t_1__719_,t_1__718_,t_1__717_,t_1__716_,t_1__715_,
  t_1__714_,t_1__713_,t_1__712_,t_1__711_,t_1__710_,t_1__709_,t_1__708_,t_1__707_,
  t_1__706_,t_1__705_,t_1__704_,t_1__703_,t_1__702_,t_1__701_,t_1__700_,t_1__699_,
  t_1__698_,t_1__697_,t_1__696_,t_1__695_,t_1__694_,t_1__693_,t_1__692_,t_1__691_,
  t_1__690_,t_1__689_,t_1__688_,t_1__687_,t_1__686_,t_1__685_,t_1__684_,t_1__683_,
  t_1__682_,t_1__681_,t_1__680_,t_1__679_,t_1__678_,t_1__677_,t_1__676_,t_1__675_,
  t_1__674_,t_1__673_,t_1__672_,t_1__671_,t_1__670_,t_1__669_,t_1__668_,t_1__667_,
  t_1__666_,t_1__665_,t_1__664_,t_1__663_,t_1__662_,t_1__661_,t_1__660_,t_1__659_,
  t_1__658_,t_1__657_,t_1__656_,t_1__655_,t_1__654_,t_1__653_,t_1__652_,t_1__651_,
  t_1__650_,t_1__649_,t_1__648_,t_1__647_,t_1__646_,t_1__645_,t_1__644_,t_1__643_,
  t_1__642_,t_1__641_,t_1__640_,t_1__639_,t_1__638_,t_1__637_,t_1__636_,t_1__635_,
  t_1__634_,t_1__633_,t_1__632_,t_1__631_,t_1__630_,t_1__629_,t_1__628_,t_1__627_,
  t_1__626_,t_1__625_,t_1__624_,t_1__623_,t_1__622_,t_1__621_,t_1__620_,t_1__619_,
  t_1__618_,t_1__617_,t_1__616_,t_1__615_,t_1__614_,t_1__613_,t_1__612_,t_1__611_,
  t_1__610_,t_1__609_,t_1__608_,t_1__607_,t_1__606_,t_1__605_,t_1__604_,t_1__603_,
  t_1__602_,t_1__601_,t_1__600_,t_1__599_,t_1__598_,t_1__597_,t_1__596_,t_1__595_,
  t_1__594_,t_1__593_,t_1__592_,t_1__591_,t_1__590_,t_1__589_,t_1__588_,t_1__587_,
  t_1__586_,t_1__585_,t_1__584_,t_1__583_,t_1__582_,t_1__581_,t_1__580_,t_1__579_,
  t_1__578_,t_1__577_,t_1__576_,t_1__575_,t_1__574_,t_1__573_,t_1__572_,t_1__571_,
  t_1__570_,t_1__569_,t_1__568_,t_1__567_,t_1__566_,t_1__565_,t_1__564_,t_1__563_,
  t_1__562_,t_1__561_,t_1__560_,t_1__559_,t_1__558_,t_1__557_,t_1__556_,t_1__555_,
  t_1__554_,t_1__553_,t_1__552_,t_1__551_,t_1__550_,t_1__549_,t_1__548_,t_1__547_,
  t_1__546_,t_1__545_,t_1__544_,t_1__543_,t_1__542_,t_1__541_,t_1__540_,t_1__539_,
  t_1__538_,t_1__537_,t_1__536_,t_1__535_,t_1__534_,t_1__533_,t_1__532_,t_1__531_,
  t_1__530_,t_1__529_,t_1__528_,t_1__527_,t_1__526_,t_1__525_,t_1__524_,t_1__523_,
  t_1__522_,t_1__521_,t_1__520_,t_1__519_,t_1__518_,t_1__517_,t_1__516_,t_1__515_,
  t_1__514_,t_1__513_,t_1__512_,t_1__511_,t_1__510_,t_1__509_,t_1__508_,t_1__507_,
  t_1__506_,t_1__505_,t_1__504_,t_1__503_,t_1__502_,t_1__501_,t_1__500_,t_1__499_,
  t_1__498_,t_1__497_,t_1__496_,t_1__495_,t_1__494_,t_1__493_,t_1__492_,t_1__491_,
  t_1__490_,t_1__489_,t_1__488_,t_1__487_,t_1__486_,t_1__485_,t_1__484_,t_1__483_,
  t_1__482_,t_1__481_,t_1__480_,t_1__479_,t_1__478_,t_1__477_,t_1__476_,t_1__475_,
  t_1__474_,t_1__473_,t_1__472_,t_1__471_,t_1__470_,t_1__469_,t_1__468_,t_1__467_,
  t_1__466_,t_1__465_,t_1__464_,t_1__463_,t_1__462_,t_1__461_,t_1__460_,t_1__459_,
  t_1__458_,t_1__457_,t_1__456_,t_1__455_,t_1__454_,t_1__453_,t_1__452_,t_1__451_,
  t_1__450_,t_1__449_,t_1__448_,t_1__447_,t_1__446_,t_1__445_,t_1__444_,t_1__443_,
  t_1__442_,t_1__441_,t_1__440_,t_1__439_,t_1__438_,t_1__437_,t_1__436_,t_1__435_,
  t_1__434_,t_1__433_,t_1__432_,t_1__431_,t_1__430_,t_1__429_,t_1__428_,t_1__427_,
  t_1__426_,t_1__425_,t_1__424_,t_1__423_,t_1__422_,t_1__421_,t_1__420_,t_1__419_,
  t_1__418_,t_1__417_,t_1__416_,t_1__415_,t_1__414_,t_1__413_,t_1__412_,t_1__411_,
  t_1__410_,t_1__409_,t_1__408_,t_1__407_,t_1__406_,t_1__405_,t_1__404_,t_1__403_,
  t_1__402_,t_1__401_,t_1__400_,t_1__399_,t_1__398_,t_1__397_,t_1__396_,t_1__395_,
  t_1__394_,t_1__393_,t_1__392_,t_1__391_,t_1__390_,t_1__389_,t_1__388_,t_1__387_,
  t_1__386_,t_1__385_,t_1__384_,t_1__383_,t_1__382_,t_1__381_,t_1__380_,t_1__379_,
  t_1__378_,t_1__377_,t_1__376_,t_1__375_,t_1__374_,t_1__373_,t_1__372_,t_1__371_,
  t_1__370_,t_1__369_,t_1__368_,t_1__367_,t_1__366_,t_1__365_,t_1__364_,t_1__363_,
  t_1__362_,t_1__361_,t_1__360_,t_1__359_,t_1__358_,t_1__357_,t_1__356_,t_1__355_,
  t_1__354_,t_1__353_,t_1__352_,t_1__351_,t_1__350_,t_1__349_,t_1__348_,t_1__347_,
  t_1__346_,t_1__345_,t_1__344_,t_1__343_,t_1__342_,t_1__341_,t_1__340_,t_1__339_,
  t_1__338_,t_1__337_,t_1__336_,t_1__335_,t_1__334_,t_1__333_,t_1__332_,t_1__331_,
  t_1__330_,t_1__329_,t_1__328_,t_1__327_,t_1__326_,t_1__325_,t_1__324_,t_1__323_,
  t_1__322_,t_1__321_,t_1__320_,t_1__319_,t_1__318_,t_1__317_,t_1__316_,t_1__315_,
  t_1__314_,t_1__313_,t_1__312_,t_1__311_,t_1__310_,t_1__309_,t_1__308_,t_1__307_,
  t_1__306_,t_1__305_,t_1__304_,t_1__303_,t_1__302_,t_1__301_,t_1__300_,t_1__299_,
  t_1__298_,t_1__297_,t_1__296_,t_1__295_,t_1__294_,t_1__293_,t_1__292_,t_1__291_,
  t_1__290_,t_1__289_,t_1__288_,t_1__287_,t_1__286_,t_1__285_,t_1__284_,t_1__283_,
  t_1__282_,t_1__281_,t_1__280_,t_1__279_,t_1__278_,t_1__277_,t_1__276_,t_1__275_,
  t_1__274_,t_1__273_,t_1__272_,t_1__271_,t_1__270_,t_1__269_,t_1__268_,t_1__267_,
  t_1__266_,t_1__265_,t_1__264_,t_1__263_,t_1__262_,t_1__261_,t_1__260_,t_1__259_,
  t_1__258_,t_1__257_,t_1__256_,t_1__255_,t_1__254_,t_1__253_,t_1__252_,t_1__251_,
  t_1__250_,t_1__249_,t_1__248_,t_1__247_,t_1__246_,t_1__245_,t_1__244_,t_1__243_,
  t_1__242_,t_1__241_,t_1__240_,t_1__239_,t_1__238_,t_1__237_,t_1__236_,t_1__235_,
  t_1__234_,t_1__233_,t_1__232_,t_1__231_,t_1__230_,t_1__229_,t_1__228_,t_1__227_,
  t_1__226_,t_1__225_,t_1__224_,t_1__223_,t_1__222_,t_1__221_,t_1__220_,t_1__219_,
  t_1__218_,t_1__217_,t_1__216_,t_1__215_,t_1__214_,t_1__213_,t_1__212_,t_1__211_,
  t_1__210_,t_1__209_,t_1__208_,t_1__207_,t_1__206_,t_1__205_,t_1__204_,t_1__203_,
  t_1__202_,t_1__201_,t_1__200_,t_1__199_,t_1__198_,t_1__197_,t_1__196_,t_1__195_,
  t_1__194_,t_1__193_,t_1__192_,t_1__191_,t_1__190_,t_1__189_,t_1__188_,t_1__187_,
  t_1__186_,t_1__185_,t_1__184_,t_1__183_,t_1__182_,t_1__181_,t_1__180_,t_1__179_,
  t_1__178_,t_1__177_,t_1__176_,t_1__175_,t_1__174_,t_1__173_,t_1__172_,t_1__171_,
  t_1__170_,t_1__169_,t_1__168_,t_1__167_,t_1__166_,t_1__165_,t_1__164_,t_1__163_,
  t_1__162_,t_1__161_,t_1__160_,t_1__159_,t_1__158_,t_1__157_,t_1__156_,t_1__155_,
  t_1__154_,t_1__153_,t_1__152_,t_1__151_,t_1__150_,t_1__149_,t_1__148_,t_1__147_,
  t_1__146_,t_1__145_,t_1__144_,t_1__143_,t_1__142_,t_1__141_,t_1__140_,t_1__139_,
  t_1__138_,t_1__137_,t_1__136_,t_1__135_,t_1__134_,t_1__133_,t_1__132_,t_1__131_,
  t_1__130_,t_1__129_,t_1__128_,t_1__127_,t_1__126_,t_1__125_,t_1__124_,t_1__123_,
  t_1__122_,t_1__121_,t_1__120_,t_1__119_,t_1__118_,t_1__117_,t_1__116_,t_1__115_,
  t_1__114_,t_1__113_,t_1__112_,t_1__111_,t_1__110_,t_1__109_,t_1__108_,t_1__107_,
  t_1__106_,t_1__105_,t_1__104_,t_1__103_,t_1__102_,t_1__101_,t_1__100_,t_1__99_,
  t_1__98_,t_1__97_,t_1__96_,t_1__95_,t_1__94_,t_1__93_,t_1__92_,t_1__91_,t_1__90_,
  t_1__89_,t_1__88_,t_1__87_,t_1__86_,t_1__85_,t_1__84_,t_1__83_,t_1__82_,t_1__81_,
  t_1__80_,t_1__79_,t_1__78_,t_1__77_,t_1__76_,t_1__75_,t_1__74_,t_1__73_,t_1__72_,
  t_1__71_,t_1__70_,t_1__69_,t_1__68_,t_1__67_,t_1__66_,t_1__65_,t_1__64_,t_1__63_,
  t_1__62_,t_1__61_,t_1__60_,t_1__59_,t_1__58_,t_1__57_,t_1__56_,t_1__55_,t_1__54_,
  t_1__53_,t_1__52_,t_1__51_,t_1__50_,t_1__49_,t_1__48_,t_1__47_,t_1__46_,t_1__45_,
  t_1__44_,t_1__43_,t_1__42_,t_1__41_,t_1__40_,t_1__39_,t_1__38_,t_1__37_,t_1__36_,
  t_1__35_,t_1__34_,t_1__33_,t_1__32_,t_1__31_,t_1__30_,t_1__29_,t_1__28_,
  t_1__27_,t_1__26_,t_1__25_,t_1__24_,t_1__23_,t_1__22_,t_1__21_,t_1__20_,t_1__19_,
  t_1__18_,t_1__17_,t_1__16_,t_1__15_,t_1__14_,t_1__13_,t_1__12_,t_1__11_,t_1__10_,
  t_1__9_,t_1__8_,t_1__7_,t_1__6_,t_1__5_,t_1__4_,t_1__3_,t_1__2_,t_1__1_,t_1__0_,
  t_2__1023_,t_2__1022_,t_2__1021_,t_2__1020_,t_2__1019_,t_2__1018_,t_2__1017_,
  t_2__1016_,t_2__1015_,t_2__1014_,t_2__1013_,t_2__1012_,t_2__1011_,t_2__1010_,t_2__1009_,
  t_2__1008_,t_2__1007_,t_2__1006_,t_2__1005_,t_2__1004_,t_2__1003_,t_2__1002_,
  t_2__1001_,t_2__1000_,t_2__999_,t_2__998_,t_2__997_,t_2__996_,t_2__995_,t_2__994_,
  t_2__993_,t_2__992_,t_2__991_,t_2__990_,t_2__989_,t_2__988_,t_2__987_,t_2__986_,
  t_2__985_,t_2__984_,t_2__983_,t_2__982_,t_2__981_,t_2__980_,t_2__979_,t_2__978_,
  t_2__977_,t_2__976_,t_2__975_,t_2__974_,t_2__973_,t_2__972_,t_2__971_,t_2__970_,
  t_2__969_,t_2__968_,t_2__967_,t_2__966_,t_2__965_,t_2__964_,t_2__963_,t_2__962_,
  t_2__961_,t_2__960_,t_2__959_,t_2__958_,t_2__957_,t_2__956_,t_2__955_,t_2__954_,
  t_2__953_,t_2__952_,t_2__951_,t_2__950_,t_2__949_,t_2__948_,t_2__947_,t_2__946_,
  t_2__945_,t_2__944_,t_2__943_,t_2__942_,t_2__941_,t_2__940_,t_2__939_,t_2__938_,
  t_2__937_,t_2__936_,t_2__935_,t_2__934_,t_2__933_,t_2__932_,t_2__931_,t_2__930_,
  t_2__929_,t_2__928_,t_2__927_,t_2__926_,t_2__925_,t_2__924_,t_2__923_,t_2__922_,
  t_2__921_,t_2__920_,t_2__919_,t_2__918_,t_2__917_,t_2__916_,t_2__915_,t_2__914_,
  t_2__913_,t_2__912_,t_2__911_,t_2__910_,t_2__909_,t_2__908_,t_2__907_,t_2__906_,
  t_2__905_,t_2__904_,t_2__903_,t_2__902_,t_2__901_,t_2__900_,t_2__899_,t_2__898_,
  t_2__897_,t_2__896_,t_2__895_,t_2__894_,t_2__893_,t_2__892_,t_2__891_,t_2__890_,
  t_2__889_,t_2__888_,t_2__887_,t_2__886_,t_2__885_,t_2__884_,t_2__883_,t_2__882_,
  t_2__881_,t_2__880_,t_2__879_,t_2__878_,t_2__877_,t_2__876_,t_2__875_,t_2__874_,
  t_2__873_,t_2__872_,t_2__871_,t_2__870_,t_2__869_,t_2__868_,t_2__867_,t_2__866_,
  t_2__865_,t_2__864_,t_2__863_,t_2__862_,t_2__861_,t_2__860_,t_2__859_,t_2__858_,
  t_2__857_,t_2__856_,t_2__855_,t_2__854_,t_2__853_,t_2__852_,t_2__851_,t_2__850_,
  t_2__849_,t_2__848_,t_2__847_,t_2__846_,t_2__845_,t_2__844_,t_2__843_,t_2__842_,
  t_2__841_,t_2__840_,t_2__839_,t_2__838_,t_2__837_,t_2__836_,t_2__835_,t_2__834_,
  t_2__833_,t_2__832_,t_2__831_,t_2__830_,t_2__829_,t_2__828_,t_2__827_,t_2__826_,
  t_2__825_,t_2__824_,t_2__823_,t_2__822_,t_2__821_,t_2__820_,t_2__819_,t_2__818_,
  t_2__817_,t_2__816_,t_2__815_,t_2__814_,t_2__813_,t_2__812_,t_2__811_,t_2__810_,
  t_2__809_,t_2__808_,t_2__807_,t_2__806_,t_2__805_,t_2__804_,t_2__803_,t_2__802_,
  t_2__801_,t_2__800_,t_2__799_,t_2__798_,t_2__797_,t_2__796_,t_2__795_,t_2__794_,
  t_2__793_,t_2__792_,t_2__791_,t_2__790_,t_2__789_,t_2__788_,t_2__787_,t_2__786_,
  t_2__785_,t_2__784_,t_2__783_,t_2__782_,t_2__781_,t_2__780_,t_2__779_,t_2__778_,
  t_2__777_,t_2__776_,t_2__775_,t_2__774_,t_2__773_,t_2__772_,t_2__771_,t_2__770_,
  t_2__769_,t_2__768_,t_2__767_,t_2__766_,t_2__765_,t_2__764_,t_2__763_,t_2__762_,
  t_2__761_,t_2__760_,t_2__759_,t_2__758_,t_2__757_,t_2__756_,t_2__755_,t_2__754_,
  t_2__753_,t_2__752_,t_2__751_,t_2__750_,t_2__749_,t_2__748_,t_2__747_,t_2__746_,
  t_2__745_,t_2__744_,t_2__743_,t_2__742_,t_2__741_,t_2__740_,t_2__739_,t_2__738_,
  t_2__737_,t_2__736_,t_2__735_,t_2__734_,t_2__733_,t_2__732_,t_2__731_,t_2__730_,
  t_2__729_,t_2__728_,t_2__727_,t_2__726_,t_2__725_,t_2__724_,t_2__723_,t_2__722_,
  t_2__721_,t_2__720_,t_2__719_,t_2__718_,t_2__717_,t_2__716_,t_2__715_,t_2__714_,
  t_2__713_,t_2__712_,t_2__711_,t_2__710_,t_2__709_,t_2__708_,t_2__707_,t_2__706_,
  t_2__705_,t_2__704_,t_2__703_,t_2__702_,t_2__701_,t_2__700_,t_2__699_,t_2__698_,
  t_2__697_,t_2__696_,t_2__695_,t_2__694_,t_2__693_,t_2__692_,t_2__691_,t_2__690_,
  t_2__689_,t_2__688_,t_2__687_,t_2__686_,t_2__685_,t_2__684_,t_2__683_,t_2__682_,
  t_2__681_,t_2__680_,t_2__679_,t_2__678_,t_2__677_,t_2__676_,t_2__675_,t_2__674_,
  t_2__673_,t_2__672_,t_2__671_,t_2__670_,t_2__669_,t_2__668_,t_2__667_,t_2__666_,
  t_2__665_,t_2__664_,t_2__663_,t_2__662_,t_2__661_,t_2__660_,t_2__659_,t_2__658_,
  t_2__657_,t_2__656_,t_2__655_,t_2__654_,t_2__653_,t_2__652_,t_2__651_,t_2__650_,
  t_2__649_,t_2__648_,t_2__647_,t_2__646_,t_2__645_,t_2__644_,t_2__643_,t_2__642_,
  t_2__641_,t_2__640_,t_2__639_,t_2__638_,t_2__637_,t_2__636_,t_2__635_,t_2__634_,
  t_2__633_,t_2__632_,t_2__631_,t_2__630_,t_2__629_,t_2__628_,t_2__627_,t_2__626_,
  t_2__625_,t_2__624_,t_2__623_,t_2__622_,t_2__621_,t_2__620_,t_2__619_,t_2__618_,
  t_2__617_,t_2__616_,t_2__615_,t_2__614_,t_2__613_,t_2__612_,t_2__611_,t_2__610_,
  t_2__609_,t_2__608_,t_2__607_,t_2__606_,t_2__605_,t_2__604_,t_2__603_,t_2__602_,
  t_2__601_,t_2__600_,t_2__599_,t_2__598_,t_2__597_,t_2__596_,t_2__595_,t_2__594_,
  t_2__593_,t_2__592_,t_2__591_,t_2__590_,t_2__589_,t_2__588_,t_2__587_,t_2__586_,
  t_2__585_,t_2__584_,t_2__583_,t_2__582_,t_2__581_,t_2__580_,t_2__579_,t_2__578_,
  t_2__577_,t_2__576_,t_2__575_,t_2__574_,t_2__573_,t_2__572_,t_2__571_,t_2__570_,
  t_2__569_,t_2__568_,t_2__567_,t_2__566_,t_2__565_,t_2__564_,t_2__563_,t_2__562_,
  t_2__561_,t_2__560_,t_2__559_,t_2__558_,t_2__557_,t_2__556_,t_2__555_,t_2__554_,
  t_2__553_,t_2__552_,t_2__551_,t_2__550_,t_2__549_,t_2__548_,t_2__547_,t_2__546_,
  t_2__545_,t_2__544_,t_2__543_,t_2__542_,t_2__541_,t_2__540_,t_2__539_,t_2__538_,
  t_2__537_,t_2__536_,t_2__535_,t_2__534_,t_2__533_,t_2__532_,t_2__531_,t_2__530_,
  t_2__529_,t_2__528_,t_2__527_,t_2__526_,t_2__525_,t_2__524_,t_2__523_,t_2__522_,
  t_2__521_,t_2__520_,t_2__519_,t_2__518_,t_2__517_,t_2__516_,t_2__515_,t_2__514_,
  t_2__513_,t_2__512_,t_2__511_,t_2__510_,t_2__509_,t_2__508_,t_2__507_,t_2__506_,
  t_2__505_,t_2__504_,t_2__503_,t_2__502_,t_2__501_,t_2__500_,t_2__499_,t_2__498_,
  t_2__497_,t_2__496_,t_2__495_,t_2__494_,t_2__493_,t_2__492_,t_2__491_,t_2__490_,
  t_2__489_,t_2__488_,t_2__487_,t_2__486_,t_2__485_,t_2__484_,t_2__483_,t_2__482_,
  t_2__481_,t_2__480_,t_2__479_,t_2__478_,t_2__477_,t_2__476_,t_2__475_,t_2__474_,
  t_2__473_,t_2__472_,t_2__471_,t_2__470_,t_2__469_,t_2__468_,t_2__467_,t_2__466_,
  t_2__465_,t_2__464_,t_2__463_,t_2__462_,t_2__461_,t_2__460_,t_2__459_,t_2__458_,
  t_2__457_,t_2__456_,t_2__455_,t_2__454_,t_2__453_,t_2__452_,t_2__451_,t_2__450_,
  t_2__449_,t_2__448_,t_2__447_,t_2__446_,t_2__445_,t_2__444_,t_2__443_,t_2__442_,
  t_2__441_,t_2__440_,t_2__439_,t_2__438_,t_2__437_,t_2__436_,t_2__435_,t_2__434_,
  t_2__433_,t_2__432_,t_2__431_,t_2__430_,t_2__429_,t_2__428_,t_2__427_,t_2__426_,
  t_2__425_,t_2__424_,t_2__423_,t_2__422_,t_2__421_,t_2__420_,t_2__419_,t_2__418_,
  t_2__417_,t_2__416_,t_2__415_,t_2__414_,t_2__413_,t_2__412_,t_2__411_,t_2__410_,
  t_2__409_,t_2__408_,t_2__407_,t_2__406_,t_2__405_,t_2__404_,t_2__403_,t_2__402_,
  t_2__401_,t_2__400_,t_2__399_,t_2__398_,t_2__397_,t_2__396_,t_2__395_,t_2__394_,
  t_2__393_,t_2__392_,t_2__391_,t_2__390_,t_2__389_,t_2__388_,t_2__387_,t_2__386_,
  t_2__385_,t_2__384_,t_2__383_,t_2__382_,t_2__381_,t_2__380_,t_2__379_,t_2__378_,
  t_2__377_,t_2__376_,t_2__375_,t_2__374_,t_2__373_,t_2__372_,t_2__371_,t_2__370_,
  t_2__369_,t_2__368_,t_2__367_,t_2__366_,t_2__365_,t_2__364_,t_2__363_,t_2__362_,
  t_2__361_,t_2__360_,t_2__359_,t_2__358_,t_2__357_,t_2__356_,t_2__355_,t_2__354_,
  t_2__353_,t_2__352_,t_2__351_,t_2__350_,t_2__349_,t_2__348_,t_2__347_,t_2__346_,
  t_2__345_,t_2__344_,t_2__343_,t_2__342_,t_2__341_,t_2__340_,t_2__339_,t_2__338_,
  t_2__337_,t_2__336_,t_2__335_,t_2__334_,t_2__333_,t_2__332_,t_2__331_,t_2__330_,
  t_2__329_,t_2__328_,t_2__327_,t_2__326_,t_2__325_,t_2__324_,t_2__323_,t_2__322_,
  t_2__321_,t_2__320_,t_2__319_,t_2__318_,t_2__317_,t_2__316_,t_2__315_,t_2__314_,
  t_2__313_,t_2__312_,t_2__311_,t_2__310_,t_2__309_,t_2__308_,t_2__307_,t_2__306_,
  t_2__305_,t_2__304_,t_2__303_,t_2__302_,t_2__301_,t_2__300_,t_2__299_,t_2__298_,
  t_2__297_,t_2__296_,t_2__295_,t_2__294_,t_2__293_,t_2__292_,t_2__291_,t_2__290_,
  t_2__289_,t_2__288_,t_2__287_,t_2__286_,t_2__285_,t_2__284_,t_2__283_,t_2__282_,
  t_2__281_,t_2__280_,t_2__279_,t_2__278_,t_2__277_,t_2__276_,t_2__275_,t_2__274_,
  t_2__273_,t_2__272_,t_2__271_,t_2__270_,t_2__269_,t_2__268_,t_2__267_,t_2__266_,
  t_2__265_,t_2__264_,t_2__263_,t_2__262_,t_2__261_,t_2__260_,t_2__259_,t_2__258_,
  t_2__257_,t_2__256_,t_2__255_,t_2__254_,t_2__253_,t_2__252_,t_2__251_,t_2__250_,
  t_2__249_,t_2__248_,t_2__247_,t_2__246_,t_2__245_,t_2__244_,t_2__243_,t_2__242_,
  t_2__241_,t_2__240_,t_2__239_,t_2__238_,t_2__237_,t_2__236_,t_2__235_,t_2__234_,
  t_2__233_,t_2__232_,t_2__231_,t_2__230_,t_2__229_,t_2__228_,t_2__227_,t_2__226_,
  t_2__225_,t_2__224_,t_2__223_,t_2__222_,t_2__221_,t_2__220_,t_2__219_,t_2__218_,
  t_2__217_,t_2__216_,t_2__215_,t_2__214_,t_2__213_,t_2__212_,t_2__211_,t_2__210_,
  t_2__209_,t_2__208_,t_2__207_,t_2__206_,t_2__205_,t_2__204_,t_2__203_,t_2__202_,
  t_2__201_,t_2__200_,t_2__199_,t_2__198_,t_2__197_,t_2__196_,t_2__195_,t_2__194_,
  t_2__193_,t_2__192_,t_2__191_,t_2__190_,t_2__189_,t_2__188_,t_2__187_,t_2__186_,
  t_2__185_,t_2__184_,t_2__183_,t_2__182_,t_2__181_,t_2__180_,t_2__179_,t_2__178_,
  t_2__177_,t_2__176_,t_2__175_,t_2__174_,t_2__173_,t_2__172_,t_2__171_,t_2__170_,
  t_2__169_,t_2__168_,t_2__167_,t_2__166_,t_2__165_,t_2__164_,t_2__163_,t_2__162_,
  t_2__161_,t_2__160_,t_2__159_,t_2__158_,t_2__157_,t_2__156_,t_2__155_,t_2__154_,
  t_2__153_,t_2__152_,t_2__151_,t_2__150_,t_2__149_,t_2__148_,t_2__147_,t_2__146_,
  t_2__145_,t_2__144_,t_2__143_,t_2__142_,t_2__141_,t_2__140_,t_2__139_,t_2__138_,
  t_2__137_,t_2__136_,t_2__135_,t_2__134_,t_2__133_,t_2__132_,t_2__131_,t_2__130_,
  t_2__129_,t_2__128_,t_2__127_,t_2__126_,t_2__125_,t_2__124_,t_2__123_,t_2__122_,
  t_2__121_,t_2__120_,t_2__119_,t_2__118_,t_2__117_,t_2__116_,t_2__115_,t_2__114_,
  t_2__113_,t_2__112_,t_2__111_,t_2__110_,t_2__109_,t_2__108_,t_2__107_,t_2__106_,
  t_2__105_,t_2__104_,t_2__103_,t_2__102_,t_2__101_,t_2__100_,t_2__99_,t_2__98_,
  t_2__97_,t_2__96_,t_2__95_,t_2__94_,t_2__93_,t_2__92_,t_2__91_,t_2__90_,t_2__89_,
  t_2__88_,t_2__87_,t_2__86_,t_2__85_,t_2__84_,t_2__83_,t_2__82_,t_2__81_,t_2__80_,
  t_2__79_,t_2__78_,t_2__77_,t_2__76_,t_2__75_,t_2__74_,t_2__73_,t_2__72_,t_2__71_,
  t_2__70_,t_2__69_,t_2__68_,t_2__67_,t_2__66_,t_2__65_,t_2__64_,t_2__63_,t_2__62_,
  t_2__61_,t_2__60_,t_2__59_,t_2__58_,t_2__57_,t_2__56_,t_2__55_,t_2__54_,
  t_2__53_,t_2__52_,t_2__51_,t_2__50_,t_2__49_,t_2__48_,t_2__47_,t_2__46_,t_2__45_,
  t_2__44_,t_2__43_,t_2__42_,t_2__41_,t_2__40_,t_2__39_,t_2__38_,t_2__37_,t_2__36_,
  t_2__35_,t_2__34_,t_2__33_,t_2__32_,t_2__31_,t_2__30_,t_2__29_,t_2__28_,t_2__27_,
  t_2__26_,t_2__25_,t_2__24_,t_2__23_,t_2__22_,t_2__21_,t_2__20_,t_2__19_,t_2__18_,
  t_2__17_,t_2__16_,t_2__15_,t_2__14_,t_2__13_,t_2__12_,t_2__11_,t_2__10_,t_2__9_,
  t_2__8_,t_2__7_,t_2__6_,t_2__5_,t_2__4_,t_2__3_,t_2__2_,t_2__1_,t_2__0_,t_3__1023_,
  t_3__1022_,t_3__1021_,t_3__1020_,t_3__1019_,t_3__1018_,t_3__1017_,t_3__1016_,
  t_3__1015_,t_3__1014_,t_3__1013_,t_3__1012_,t_3__1011_,t_3__1010_,t_3__1009_,
  t_3__1008_,t_3__1007_,t_3__1006_,t_3__1005_,t_3__1004_,t_3__1003_,t_3__1002_,
  t_3__1001_,t_3__1000_,t_3__999_,t_3__998_,t_3__997_,t_3__996_,t_3__995_,t_3__994_,
  t_3__993_,t_3__992_,t_3__991_,t_3__990_,t_3__989_,t_3__988_,t_3__987_,t_3__986_,
  t_3__985_,t_3__984_,t_3__983_,t_3__982_,t_3__981_,t_3__980_,t_3__979_,t_3__978_,
  t_3__977_,t_3__976_,t_3__975_,t_3__974_,t_3__973_,t_3__972_,t_3__971_,t_3__970_,
  t_3__969_,t_3__968_,t_3__967_,t_3__966_,t_3__965_,t_3__964_,t_3__963_,t_3__962_,
  t_3__961_,t_3__960_,t_3__959_,t_3__958_,t_3__957_,t_3__956_,t_3__955_,t_3__954_,
  t_3__953_,t_3__952_,t_3__951_,t_3__950_,t_3__949_,t_3__948_,t_3__947_,t_3__946_,
  t_3__945_,t_3__944_,t_3__943_,t_3__942_,t_3__941_,t_3__940_,t_3__939_,t_3__938_,
  t_3__937_,t_3__936_,t_3__935_,t_3__934_,t_3__933_,t_3__932_,t_3__931_,t_3__930_,
  t_3__929_,t_3__928_,t_3__927_,t_3__926_,t_3__925_,t_3__924_,t_3__923_,t_3__922_,
  t_3__921_,t_3__920_,t_3__919_,t_3__918_,t_3__917_,t_3__916_,t_3__915_,t_3__914_,
  t_3__913_,t_3__912_,t_3__911_,t_3__910_,t_3__909_,t_3__908_,t_3__907_,t_3__906_,
  t_3__905_,t_3__904_,t_3__903_,t_3__902_,t_3__901_,t_3__900_,t_3__899_,t_3__898_,
  t_3__897_,t_3__896_,t_3__895_,t_3__894_,t_3__893_,t_3__892_,t_3__891_,t_3__890_,
  t_3__889_,t_3__888_,t_3__887_,t_3__886_,t_3__885_,t_3__884_,t_3__883_,t_3__882_,
  t_3__881_,t_3__880_,t_3__879_,t_3__878_,t_3__877_,t_3__876_,t_3__875_,t_3__874_,
  t_3__873_,t_3__872_,t_3__871_,t_3__870_,t_3__869_,t_3__868_,t_3__867_,t_3__866_,
  t_3__865_,t_3__864_,t_3__863_,t_3__862_,t_3__861_,t_3__860_,t_3__859_,t_3__858_,
  t_3__857_,t_3__856_,t_3__855_,t_3__854_,t_3__853_,t_3__852_,t_3__851_,t_3__850_,
  t_3__849_,t_3__848_,t_3__847_,t_3__846_,t_3__845_,t_3__844_,t_3__843_,t_3__842_,
  t_3__841_,t_3__840_,t_3__839_,t_3__838_,t_3__837_,t_3__836_,t_3__835_,t_3__834_,
  t_3__833_,t_3__832_,t_3__831_,t_3__830_,t_3__829_,t_3__828_,t_3__827_,t_3__826_,
  t_3__825_,t_3__824_,t_3__823_,t_3__822_,t_3__821_,t_3__820_,t_3__819_,t_3__818_,
  t_3__817_,t_3__816_,t_3__815_,t_3__814_,t_3__813_,t_3__812_,t_3__811_,t_3__810_,
  t_3__809_,t_3__808_,t_3__807_,t_3__806_,t_3__805_,t_3__804_,t_3__803_,t_3__802_,
  t_3__801_,t_3__800_,t_3__799_,t_3__798_,t_3__797_,t_3__796_,t_3__795_,t_3__794_,
  t_3__793_,t_3__792_,t_3__791_,t_3__790_,t_3__789_,t_3__788_,t_3__787_,t_3__786_,
  t_3__785_,t_3__784_,t_3__783_,t_3__782_,t_3__781_,t_3__780_,t_3__779_,t_3__778_,
  t_3__777_,t_3__776_,t_3__775_,t_3__774_,t_3__773_,t_3__772_,t_3__771_,t_3__770_,
  t_3__769_,t_3__768_,t_3__767_,t_3__766_,t_3__765_,t_3__764_,t_3__763_,t_3__762_,
  t_3__761_,t_3__760_,t_3__759_,t_3__758_,t_3__757_,t_3__756_,t_3__755_,t_3__754_,
  t_3__753_,t_3__752_,t_3__751_,t_3__750_,t_3__749_,t_3__748_,t_3__747_,t_3__746_,
  t_3__745_,t_3__744_,t_3__743_,t_3__742_,t_3__741_,t_3__740_,t_3__739_,t_3__738_,
  t_3__737_,t_3__736_,t_3__735_,t_3__734_,t_3__733_,t_3__732_,t_3__731_,t_3__730_,
  t_3__729_,t_3__728_,t_3__727_,t_3__726_,t_3__725_,t_3__724_,t_3__723_,t_3__722_,
  t_3__721_,t_3__720_,t_3__719_,t_3__718_,t_3__717_,t_3__716_,t_3__715_,t_3__714_,
  t_3__713_,t_3__712_,t_3__711_,t_3__710_,t_3__709_,t_3__708_,t_3__707_,t_3__706_,
  t_3__705_,t_3__704_,t_3__703_,t_3__702_,t_3__701_,t_3__700_,t_3__699_,t_3__698_,
  t_3__697_,t_3__696_,t_3__695_,t_3__694_,t_3__693_,t_3__692_,t_3__691_,t_3__690_,
  t_3__689_,t_3__688_,t_3__687_,t_3__686_,t_3__685_,t_3__684_,t_3__683_,t_3__682_,
  t_3__681_,t_3__680_,t_3__679_,t_3__678_,t_3__677_,t_3__676_,t_3__675_,t_3__674_,
  t_3__673_,t_3__672_,t_3__671_,t_3__670_,t_3__669_,t_3__668_,t_3__667_,t_3__666_,
  t_3__665_,t_3__664_,t_3__663_,t_3__662_,t_3__661_,t_3__660_,t_3__659_,t_3__658_,
  t_3__657_,t_3__656_,t_3__655_,t_3__654_,t_3__653_,t_3__652_,t_3__651_,t_3__650_,
  t_3__649_,t_3__648_,t_3__647_,t_3__646_,t_3__645_,t_3__644_,t_3__643_,t_3__642_,
  t_3__641_,t_3__640_,t_3__639_,t_3__638_,t_3__637_,t_3__636_,t_3__635_,t_3__634_,
  t_3__633_,t_3__632_,t_3__631_,t_3__630_,t_3__629_,t_3__628_,t_3__627_,t_3__626_,
  t_3__625_,t_3__624_,t_3__623_,t_3__622_,t_3__621_,t_3__620_,t_3__619_,t_3__618_,
  t_3__617_,t_3__616_,t_3__615_,t_3__614_,t_3__613_,t_3__612_,t_3__611_,t_3__610_,
  t_3__609_,t_3__608_,t_3__607_,t_3__606_,t_3__605_,t_3__604_,t_3__603_,t_3__602_,
  t_3__601_,t_3__600_,t_3__599_,t_3__598_,t_3__597_,t_3__596_,t_3__595_,t_3__594_,
  t_3__593_,t_3__592_,t_3__591_,t_3__590_,t_3__589_,t_3__588_,t_3__587_,t_3__586_,
  t_3__585_,t_3__584_,t_3__583_,t_3__582_,t_3__581_,t_3__580_,t_3__579_,t_3__578_,
  t_3__577_,t_3__576_,t_3__575_,t_3__574_,t_3__573_,t_3__572_,t_3__571_,t_3__570_,
  t_3__569_,t_3__568_,t_3__567_,t_3__566_,t_3__565_,t_3__564_,t_3__563_,t_3__562_,
  t_3__561_,t_3__560_,t_3__559_,t_3__558_,t_3__557_,t_3__556_,t_3__555_,t_3__554_,
  t_3__553_,t_3__552_,t_3__551_,t_3__550_,t_3__549_,t_3__548_,t_3__547_,t_3__546_,
  t_3__545_,t_3__544_,t_3__543_,t_3__542_,t_3__541_,t_3__540_,t_3__539_,t_3__538_,
  t_3__537_,t_3__536_,t_3__535_,t_3__534_,t_3__533_,t_3__532_,t_3__531_,t_3__530_,
  t_3__529_,t_3__528_,t_3__527_,t_3__526_,t_3__525_,t_3__524_,t_3__523_,t_3__522_,
  t_3__521_,t_3__520_,t_3__519_,t_3__518_,t_3__517_,t_3__516_,t_3__515_,t_3__514_,
  t_3__513_,t_3__512_,t_3__511_,t_3__510_,t_3__509_,t_3__508_,t_3__507_,t_3__506_,
  t_3__505_,t_3__504_,t_3__503_,t_3__502_,t_3__501_,t_3__500_,t_3__499_,t_3__498_,
  t_3__497_,t_3__496_,t_3__495_,t_3__494_,t_3__493_,t_3__492_,t_3__491_,t_3__490_,
  t_3__489_,t_3__488_,t_3__487_,t_3__486_,t_3__485_,t_3__484_,t_3__483_,t_3__482_,
  t_3__481_,t_3__480_,t_3__479_,t_3__478_,t_3__477_,t_3__476_,t_3__475_,t_3__474_,
  t_3__473_,t_3__472_,t_3__471_,t_3__470_,t_3__469_,t_3__468_,t_3__467_,t_3__466_,
  t_3__465_,t_3__464_,t_3__463_,t_3__462_,t_3__461_,t_3__460_,t_3__459_,t_3__458_,
  t_3__457_,t_3__456_,t_3__455_,t_3__454_,t_3__453_,t_3__452_,t_3__451_,t_3__450_,
  t_3__449_,t_3__448_,t_3__447_,t_3__446_,t_3__445_,t_3__444_,t_3__443_,t_3__442_,
  t_3__441_,t_3__440_,t_3__439_,t_3__438_,t_3__437_,t_3__436_,t_3__435_,t_3__434_,
  t_3__433_,t_3__432_,t_3__431_,t_3__430_,t_3__429_,t_3__428_,t_3__427_,t_3__426_,
  t_3__425_,t_3__424_,t_3__423_,t_3__422_,t_3__421_,t_3__420_,t_3__419_,t_3__418_,
  t_3__417_,t_3__416_,t_3__415_,t_3__414_,t_3__413_,t_3__412_,t_3__411_,t_3__410_,
  t_3__409_,t_3__408_,t_3__407_,t_3__406_,t_3__405_,t_3__404_,t_3__403_,t_3__402_,
  t_3__401_,t_3__400_,t_3__399_,t_3__398_,t_3__397_,t_3__396_,t_3__395_,t_3__394_,
  t_3__393_,t_3__392_,t_3__391_,t_3__390_,t_3__389_,t_3__388_,t_3__387_,t_3__386_,
  t_3__385_,t_3__384_,t_3__383_,t_3__382_,t_3__381_,t_3__380_,t_3__379_,t_3__378_,
  t_3__377_,t_3__376_,t_3__375_,t_3__374_,t_3__373_,t_3__372_,t_3__371_,t_3__370_,
  t_3__369_,t_3__368_,t_3__367_,t_3__366_,t_3__365_,t_3__364_,t_3__363_,t_3__362_,
  t_3__361_,t_3__360_,t_3__359_,t_3__358_,t_3__357_,t_3__356_,t_3__355_,t_3__354_,
  t_3__353_,t_3__352_,t_3__351_,t_3__350_,t_3__349_,t_3__348_,t_3__347_,t_3__346_,
  t_3__345_,t_3__344_,t_3__343_,t_3__342_,t_3__341_,t_3__340_,t_3__339_,t_3__338_,
  t_3__337_,t_3__336_,t_3__335_,t_3__334_,t_3__333_,t_3__332_,t_3__331_,t_3__330_,
  t_3__329_,t_3__328_,t_3__327_,t_3__326_,t_3__325_,t_3__324_,t_3__323_,t_3__322_,
  t_3__321_,t_3__320_,t_3__319_,t_3__318_,t_3__317_,t_3__316_,t_3__315_,t_3__314_,
  t_3__313_,t_3__312_,t_3__311_,t_3__310_,t_3__309_,t_3__308_,t_3__307_,t_3__306_,
  t_3__305_,t_3__304_,t_3__303_,t_3__302_,t_3__301_,t_3__300_,t_3__299_,t_3__298_,
  t_3__297_,t_3__296_,t_3__295_,t_3__294_,t_3__293_,t_3__292_,t_3__291_,t_3__290_,
  t_3__289_,t_3__288_,t_3__287_,t_3__286_,t_3__285_,t_3__284_,t_3__283_,t_3__282_,
  t_3__281_,t_3__280_,t_3__279_,t_3__278_,t_3__277_,t_3__276_,t_3__275_,t_3__274_,
  t_3__273_,t_3__272_,t_3__271_,t_3__270_,t_3__269_,t_3__268_,t_3__267_,t_3__266_,
  t_3__265_,t_3__264_,t_3__263_,t_3__262_,t_3__261_,t_3__260_,t_3__259_,t_3__258_,
  t_3__257_,t_3__256_,t_3__255_,t_3__254_,t_3__253_,t_3__252_,t_3__251_,t_3__250_,
  t_3__249_,t_3__248_,t_3__247_,t_3__246_,t_3__245_,t_3__244_,t_3__243_,t_3__242_,
  t_3__241_,t_3__240_,t_3__239_,t_3__238_,t_3__237_,t_3__236_,t_3__235_,t_3__234_,
  t_3__233_,t_3__232_,t_3__231_,t_3__230_,t_3__229_,t_3__228_,t_3__227_,t_3__226_,
  t_3__225_,t_3__224_,t_3__223_,t_3__222_,t_3__221_,t_3__220_,t_3__219_,t_3__218_,
  t_3__217_,t_3__216_,t_3__215_,t_3__214_,t_3__213_,t_3__212_,t_3__211_,t_3__210_,
  t_3__209_,t_3__208_,t_3__207_,t_3__206_,t_3__205_,t_3__204_,t_3__203_,t_3__202_,
  t_3__201_,t_3__200_,t_3__199_,t_3__198_,t_3__197_,t_3__196_,t_3__195_,t_3__194_,
  t_3__193_,t_3__192_,t_3__191_,t_3__190_,t_3__189_,t_3__188_,t_3__187_,t_3__186_,
  t_3__185_,t_3__184_,t_3__183_,t_3__182_,t_3__181_,t_3__180_,t_3__179_,t_3__178_,
  t_3__177_,t_3__176_,t_3__175_,t_3__174_,t_3__173_,t_3__172_,t_3__171_,t_3__170_,
  t_3__169_,t_3__168_,t_3__167_,t_3__166_,t_3__165_,t_3__164_,t_3__163_,t_3__162_,
  t_3__161_,t_3__160_,t_3__159_,t_3__158_,t_3__157_,t_3__156_,t_3__155_,t_3__154_,
  t_3__153_,t_3__152_,t_3__151_,t_3__150_,t_3__149_,t_3__148_,t_3__147_,t_3__146_,
  t_3__145_,t_3__144_,t_3__143_,t_3__142_,t_3__141_,t_3__140_,t_3__139_,t_3__138_,
  t_3__137_,t_3__136_,t_3__135_,t_3__134_,t_3__133_,t_3__132_,t_3__131_,t_3__130_,
  t_3__129_,t_3__128_,t_3__127_,t_3__126_,t_3__125_,t_3__124_,t_3__123_,t_3__122_,
  t_3__121_,t_3__120_,t_3__119_,t_3__118_,t_3__117_,t_3__116_,t_3__115_,t_3__114_,
  t_3__113_,t_3__112_,t_3__111_,t_3__110_,t_3__109_,t_3__108_,t_3__107_,t_3__106_,
  t_3__105_,t_3__104_,t_3__103_,t_3__102_,t_3__101_,t_3__100_,t_3__99_,t_3__98_,t_3__97_,
  t_3__96_,t_3__95_,t_3__94_,t_3__93_,t_3__92_,t_3__91_,t_3__90_,t_3__89_,t_3__88_,
  t_3__87_,t_3__86_,t_3__85_,t_3__84_,t_3__83_,t_3__82_,t_3__81_,t_3__80_,
  t_3__79_,t_3__78_,t_3__77_,t_3__76_,t_3__75_,t_3__74_,t_3__73_,t_3__72_,t_3__71_,
  t_3__70_,t_3__69_,t_3__68_,t_3__67_,t_3__66_,t_3__65_,t_3__64_,t_3__63_,t_3__62_,
  t_3__61_,t_3__60_,t_3__59_,t_3__58_,t_3__57_,t_3__56_,t_3__55_,t_3__54_,t_3__53_,
  t_3__52_,t_3__51_,t_3__50_,t_3__49_,t_3__48_,t_3__47_,t_3__46_,t_3__45_,t_3__44_,
  t_3__43_,t_3__42_,t_3__41_,t_3__40_,t_3__39_,t_3__38_,t_3__37_,t_3__36_,t_3__35_,
  t_3__34_,t_3__33_,t_3__32_,t_3__31_,t_3__30_,t_3__29_,t_3__28_,t_3__27_,t_3__26_,
  t_3__25_,t_3__24_,t_3__23_,t_3__22_,t_3__21_,t_3__20_,t_3__19_,t_3__18_,t_3__17_,
  t_3__16_,t_3__15_,t_3__14_,t_3__13_,t_3__12_,t_3__11_,t_3__10_,t_3__9_,t_3__8_,
  t_3__7_,t_3__6_,t_3__5_,t_3__4_,t_3__3_,t_3__2_,t_3__1_,t_3__0_,t_4__1023_,
  t_4__1022_,t_4__1021_,t_4__1020_,t_4__1019_,t_4__1018_,t_4__1017_,t_4__1016_,
  t_4__1015_,t_4__1014_,t_4__1013_,t_4__1012_,t_4__1011_,t_4__1010_,t_4__1009_,t_4__1008_,
  t_4__1007_,t_4__1006_,t_4__1005_,t_4__1004_,t_4__1003_,t_4__1002_,t_4__1001_,
  t_4__1000_,t_4__999_,t_4__998_,t_4__997_,t_4__996_,t_4__995_,t_4__994_,t_4__993_,
  t_4__992_,t_4__991_,t_4__990_,t_4__989_,t_4__988_,t_4__987_,t_4__986_,t_4__985_,
  t_4__984_,t_4__983_,t_4__982_,t_4__981_,t_4__980_,t_4__979_,t_4__978_,t_4__977_,
  t_4__976_,t_4__975_,t_4__974_,t_4__973_,t_4__972_,t_4__971_,t_4__970_,t_4__969_,
  t_4__968_,t_4__967_,t_4__966_,t_4__965_,t_4__964_,t_4__963_,t_4__962_,t_4__961_,
  t_4__960_,t_4__959_,t_4__958_,t_4__957_,t_4__956_,t_4__955_,t_4__954_,t_4__953_,
  t_4__952_,t_4__951_,t_4__950_,t_4__949_,t_4__948_,t_4__947_,t_4__946_,t_4__945_,
  t_4__944_,t_4__943_,t_4__942_,t_4__941_,t_4__940_,t_4__939_,t_4__938_,t_4__937_,
  t_4__936_,t_4__935_,t_4__934_,t_4__933_,t_4__932_,t_4__931_,t_4__930_,t_4__929_,
  t_4__928_,t_4__927_,t_4__926_,t_4__925_,t_4__924_,t_4__923_,t_4__922_,t_4__921_,
  t_4__920_,t_4__919_,t_4__918_,t_4__917_,t_4__916_,t_4__915_,t_4__914_,t_4__913_,
  t_4__912_,t_4__911_,t_4__910_,t_4__909_,t_4__908_,t_4__907_,t_4__906_,t_4__905_,
  t_4__904_,t_4__903_,t_4__902_,t_4__901_,t_4__900_,t_4__899_,t_4__898_,t_4__897_,
  t_4__896_,t_4__895_,t_4__894_,t_4__893_,t_4__892_,t_4__891_,t_4__890_,t_4__889_,
  t_4__888_,t_4__887_,t_4__886_,t_4__885_,t_4__884_,t_4__883_,t_4__882_,t_4__881_,
  t_4__880_,t_4__879_,t_4__878_,t_4__877_,t_4__876_,t_4__875_,t_4__874_,t_4__873_,
  t_4__872_,t_4__871_,t_4__870_,t_4__869_,t_4__868_,t_4__867_,t_4__866_,t_4__865_,
  t_4__864_,t_4__863_,t_4__862_,t_4__861_,t_4__860_,t_4__859_,t_4__858_,t_4__857_,
  t_4__856_,t_4__855_,t_4__854_,t_4__853_,t_4__852_,t_4__851_,t_4__850_,t_4__849_,
  t_4__848_,t_4__847_,t_4__846_,t_4__845_,t_4__844_,t_4__843_,t_4__842_,t_4__841_,
  t_4__840_,t_4__839_,t_4__838_,t_4__837_,t_4__836_,t_4__835_,t_4__834_,t_4__833_,
  t_4__832_,t_4__831_,t_4__830_,t_4__829_,t_4__828_,t_4__827_,t_4__826_,t_4__825_,
  t_4__824_,t_4__823_,t_4__822_,t_4__821_,t_4__820_,t_4__819_,t_4__818_,t_4__817_,
  t_4__816_,t_4__815_,t_4__814_,t_4__813_,t_4__812_,t_4__811_,t_4__810_,t_4__809_,
  t_4__808_,t_4__807_,t_4__806_,t_4__805_,t_4__804_,t_4__803_,t_4__802_,t_4__801_,
  t_4__800_,t_4__799_,t_4__798_,t_4__797_,t_4__796_,t_4__795_,t_4__794_,t_4__793_,
  t_4__792_,t_4__791_,t_4__790_,t_4__789_,t_4__788_,t_4__787_,t_4__786_,t_4__785_,
  t_4__784_,t_4__783_,t_4__782_,t_4__781_,t_4__780_,t_4__779_,t_4__778_,t_4__777_,
  t_4__776_,t_4__775_,t_4__774_,t_4__773_,t_4__772_,t_4__771_,t_4__770_,t_4__769_,
  t_4__768_,t_4__767_,t_4__766_,t_4__765_,t_4__764_,t_4__763_,t_4__762_,t_4__761_,
  t_4__760_,t_4__759_,t_4__758_,t_4__757_,t_4__756_,t_4__755_,t_4__754_,t_4__753_,
  t_4__752_,t_4__751_,t_4__750_,t_4__749_,t_4__748_,t_4__747_,t_4__746_,t_4__745_,
  t_4__744_,t_4__743_,t_4__742_,t_4__741_,t_4__740_,t_4__739_,t_4__738_,t_4__737_,
  t_4__736_,t_4__735_,t_4__734_,t_4__733_,t_4__732_,t_4__731_,t_4__730_,t_4__729_,
  t_4__728_,t_4__727_,t_4__726_,t_4__725_,t_4__724_,t_4__723_,t_4__722_,t_4__721_,
  t_4__720_,t_4__719_,t_4__718_,t_4__717_,t_4__716_,t_4__715_,t_4__714_,t_4__713_,
  t_4__712_,t_4__711_,t_4__710_,t_4__709_,t_4__708_,t_4__707_,t_4__706_,t_4__705_,
  t_4__704_,t_4__703_,t_4__702_,t_4__701_,t_4__700_,t_4__699_,t_4__698_,t_4__697_,
  t_4__696_,t_4__695_,t_4__694_,t_4__693_,t_4__692_,t_4__691_,t_4__690_,t_4__689_,
  t_4__688_,t_4__687_,t_4__686_,t_4__685_,t_4__684_,t_4__683_,t_4__682_,t_4__681_,
  t_4__680_,t_4__679_,t_4__678_,t_4__677_,t_4__676_,t_4__675_,t_4__674_,t_4__673_,
  t_4__672_,t_4__671_,t_4__670_,t_4__669_,t_4__668_,t_4__667_,t_4__666_,t_4__665_,
  t_4__664_,t_4__663_,t_4__662_,t_4__661_,t_4__660_,t_4__659_,t_4__658_,t_4__657_,
  t_4__656_,t_4__655_,t_4__654_,t_4__653_,t_4__652_,t_4__651_,t_4__650_,t_4__649_,
  t_4__648_,t_4__647_,t_4__646_,t_4__645_,t_4__644_,t_4__643_,t_4__642_,t_4__641_,
  t_4__640_,t_4__639_,t_4__638_,t_4__637_,t_4__636_,t_4__635_,t_4__634_,t_4__633_,
  t_4__632_,t_4__631_,t_4__630_,t_4__629_,t_4__628_,t_4__627_,t_4__626_,t_4__625_,
  t_4__624_,t_4__623_,t_4__622_,t_4__621_,t_4__620_,t_4__619_,t_4__618_,t_4__617_,
  t_4__616_,t_4__615_,t_4__614_,t_4__613_,t_4__612_,t_4__611_,t_4__610_,t_4__609_,
  t_4__608_,t_4__607_,t_4__606_,t_4__605_,t_4__604_,t_4__603_,t_4__602_,t_4__601_,
  t_4__600_,t_4__599_,t_4__598_,t_4__597_,t_4__596_,t_4__595_,t_4__594_,t_4__593_,
  t_4__592_,t_4__591_,t_4__590_,t_4__589_,t_4__588_,t_4__587_,t_4__586_,t_4__585_,
  t_4__584_,t_4__583_,t_4__582_,t_4__581_,t_4__580_,t_4__579_,t_4__578_,t_4__577_,
  t_4__576_,t_4__575_,t_4__574_,t_4__573_,t_4__572_,t_4__571_,t_4__570_,t_4__569_,
  t_4__568_,t_4__567_,t_4__566_,t_4__565_,t_4__564_,t_4__563_,t_4__562_,t_4__561_,
  t_4__560_,t_4__559_,t_4__558_,t_4__557_,t_4__556_,t_4__555_,t_4__554_,t_4__553_,
  t_4__552_,t_4__551_,t_4__550_,t_4__549_,t_4__548_,t_4__547_,t_4__546_,t_4__545_,
  t_4__544_,t_4__543_,t_4__542_,t_4__541_,t_4__540_,t_4__539_,t_4__538_,t_4__537_,
  t_4__536_,t_4__535_,t_4__534_,t_4__533_,t_4__532_,t_4__531_,t_4__530_,t_4__529_,
  t_4__528_,t_4__527_,t_4__526_,t_4__525_,t_4__524_,t_4__523_,t_4__522_,t_4__521_,
  t_4__520_,t_4__519_,t_4__518_,t_4__517_,t_4__516_,t_4__515_,t_4__514_,t_4__513_,
  t_4__512_,t_4__511_,t_4__510_,t_4__509_,t_4__508_,t_4__507_,t_4__506_,t_4__505_,
  t_4__504_,t_4__503_,t_4__502_,t_4__501_,t_4__500_,t_4__499_,t_4__498_,t_4__497_,
  t_4__496_,t_4__495_,t_4__494_,t_4__493_,t_4__492_,t_4__491_,t_4__490_,t_4__489_,
  t_4__488_,t_4__487_,t_4__486_,t_4__485_,t_4__484_,t_4__483_,t_4__482_,t_4__481_,
  t_4__480_,t_4__479_,t_4__478_,t_4__477_,t_4__476_,t_4__475_,t_4__474_,t_4__473_,
  t_4__472_,t_4__471_,t_4__470_,t_4__469_,t_4__468_,t_4__467_,t_4__466_,t_4__465_,
  t_4__464_,t_4__463_,t_4__462_,t_4__461_,t_4__460_,t_4__459_,t_4__458_,t_4__457_,
  t_4__456_,t_4__455_,t_4__454_,t_4__453_,t_4__452_,t_4__451_,t_4__450_,t_4__449_,
  t_4__448_,t_4__447_,t_4__446_,t_4__445_,t_4__444_,t_4__443_,t_4__442_,t_4__441_,
  t_4__440_,t_4__439_,t_4__438_,t_4__437_,t_4__436_,t_4__435_,t_4__434_,t_4__433_,
  t_4__432_,t_4__431_,t_4__430_,t_4__429_,t_4__428_,t_4__427_,t_4__426_,t_4__425_,
  t_4__424_,t_4__423_,t_4__422_,t_4__421_,t_4__420_,t_4__419_,t_4__418_,t_4__417_,
  t_4__416_,t_4__415_,t_4__414_,t_4__413_,t_4__412_,t_4__411_,t_4__410_,t_4__409_,
  t_4__408_,t_4__407_,t_4__406_,t_4__405_,t_4__404_,t_4__403_,t_4__402_,t_4__401_,
  t_4__400_,t_4__399_,t_4__398_,t_4__397_,t_4__396_,t_4__395_,t_4__394_,t_4__393_,
  t_4__392_,t_4__391_,t_4__390_,t_4__389_,t_4__388_,t_4__387_,t_4__386_,t_4__385_,
  t_4__384_,t_4__383_,t_4__382_,t_4__381_,t_4__380_,t_4__379_,t_4__378_,t_4__377_,
  t_4__376_,t_4__375_,t_4__374_,t_4__373_,t_4__372_,t_4__371_,t_4__370_,t_4__369_,
  t_4__368_,t_4__367_,t_4__366_,t_4__365_,t_4__364_,t_4__363_,t_4__362_,t_4__361_,
  t_4__360_,t_4__359_,t_4__358_,t_4__357_,t_4__356_,t_4__355_,t_4__354_,t_4__353_,
  t_4__352_,t_4__351_,t_4__350_,t_4__349_,t_4__348_,t_4__347_,t_4__346_,t_4__345_,
  t_4__344_,t_4__343_,t_4__342_,t_4__341_,t_4__340_,t_4__339_,t_4__338_,t_4__337_,
  t_4__336_,t_4__335_,t_4__334_,t_4__333_,t_4__332_,t_4__331_,t_4__330_,t_4__329_,
  t_4__328_,t_4__327_,t_4__326_,t_4__325_,t_4__324_,t_4__323_,t_4__322_,t_4__321_,
  t_4__320_,t_4__319_,t_4__318_,t_4__317_,t_4__316_,t_4__315_,t_4__314_,t_4__313_,
  t_4__312_,t_4__311_,t_4__310_,t_4__309_,t_4__308_,t_4__307_,t_4__306_,t_4__305_,
  t_4__304_,t_4__303_,t_4__302_,t_4__301_,t_4__300_,t_4__299_,t_4__298_,t_4__297_,
  t_4__296_,t_4__295_,t_4__294_,t_4__293_,t_4__292_,t_4__291_,t_4__290_,t_4__289_,
  t_4__288_,t_4__287_,t_4__286_,t_4__285_,t_4__284_,t_4__283_,t_4__282_,t_4__281_,
  t_4__280_,t_4__279_,t_4__278_,t_4__277_,t_4__276_,t_4__275_,t_4__274_,t_4__273_,
  t_4__272_,t_4__271_,t_4__270_,t_4__269_,t_4__268_,t_4__267_,t_4__266_,t_4__265_,
  t_4__264_,t_4__263_,t_4__262_,t_4__261_,t_4__260_,t_4__259_,t_4__258_,t_4__257_,
  t_4__256_,t_4__255_,t_4__254_,t_4__253_,t_4__252_,t_4__251_,t_4__250_,t_4__249_,
  t_4__248_,t_4__247_,t_4__246_,t_4__245_,t_4__244_,t_4__243_,t_4__242_,t_4__241_,
  t_4__240_,t_4__239_,t_4__238_,t_4__237_,t_4__236_,t_4__235_,t_4__234_,t_4__233_,
  t_4__232_,t_4__231_,t_4__230_,t_4__229_,t_4__228_,t_4__227_,t_4__226_,t_4__225_,
  t_4__224_,t_4__223_,t_4__222_,t_4__221_,t_4__220_,t_4__219_,t_4__218_,t_4__217_,
  t_4__216_,t_4__215_,t_4__214_,t_4__213_,t_4__212_,t_4__211_,t_4__210_,t_4__209_,
  t_4__208_,t_4__207_,t_4__206_,t_4__205_,t_4__204_,t_4__203_,t_4__202_,t_4__201_,
  t_4__200_,t_4__199_,t_4__198_,t_4__197_,t_4__196_,t_4__195_,t_4__194_,t_4__193_,
  t_4__192_,t_4__191_,t_4__190_,t_4__189_,t_4__188_,t_4__187_,t_4__186_,t_4__185_,
  t_4__184_,t_4__183_,t_4__182_,t_4__181_,t_4__180_,t_4__179_,t_4__178_,t_4__177_,
  t_4__176_,t_4__175_,t_4__174_,t_4__173_,t_4__172_,t_4__171_,t_4__170_,t_4__169_,
  t_4__168_,t_4__167_,t_4__166_,t_4__165_,t_4__164_,t_4__163_,t_4__162_,t_4__161_,
  t_4__160_,t_4__159_,t_4__158_,t_4__157_,t_4__156_,t_4__155_,t_4__154_,t_4__153_,
  t_4__152_,t_4__151_,t_4__150_,t_4__149_,t_4__148_,t_4__147_,t_4__146_,t_4__145_,
  t_4__144_,t_4__143_,t_4__142_,t_4__141_,t_4__140_,t_4__139_,t_4__138_,t_4__137_,
  t_4__136_,t_4__135_,t_4__134_,t_4__133_,t_4__132_,t_4__131_,t_4__130_,t_4__129_,
  t_4__128_,t_4__127_,t_4__126_,t_4__125_,t_4__124_,t_4__123_,t_4__122_,t_4__121_,
  t_4__120_,t_4__119_,t_4__118_,t_4__117_,t_4__116_,t_4__115_,t_4__114_,t_4__113_,
  t_4__112_,t_4__111_,t_4__110_,t_4__109_,t_4__108_,t_4__107_,t_4__106_,t_4__105_,
  t_4__104_,t_4__103_,t_4__102_,t_4__101_,t_4__100_,t_4__99_,t_4__98_,t_4__97_,
  t_4__96_,t_4__95_,t_4__94_,t_4__93_,t_4__92_,t_4__91_,t_4__90_,t_4__89_,t_4__88_,
  t_4__87_,t_4__86_,t_4__85_,t_4__84_,t_4__83_,t_4__82_,t_4__81_,t_4__80_,t_4__79_,
  t_4__78_,t_4__77_,t_4__76_,t_4__75_,t_4__74_,t_4__73_,t_4__72_,t_4__71_,t_4__70_,
  t_4__69_,t_4__68_,t_4__67_,t_4__66_,t_4__65_,t_4__64_,t_4__63_,t_4__62_,t_4__61_,
  t_4__60_,t_4__59_,t_4__58_,t_4__57_,t_4__56_,t_4__55_,t_4__54_,t_4__53_,t_4__52_,
  t_4__51_,t_4__50_,t_4__49_,t_4__48_,t_4__47_,t_4__46_,t_4__45_,t_4__44_,t_4__43_,
  t_4__42_,t_4__41_,t_4__40_,t_4__39_,t_4__38_,t_4__37_,t_4__36_,t_4__35_,t_4__34_,
  t_4__33_,t_4__32_,t_4__31_,t_4__30_,t_4__29_,t_4__28_,t_4__27_,t_4__26_,
  t_4__25_,t_4__24_,t_4__23_,t_4__22_,t_4__21_,t_4__20_,t_4__19_,t_4__18_,t_4__17_,
  t_4__16_,t_4__15_,t_4__14_,t_4__13_,t_4__12_,t_4__11_,t_4__10_,t_4__9_,t_4__8_,t_4__7_,
  t_4__6_,t_4__5_,t_4__4_,t_4__3_,t_4__2_,t_4__1_,t_4__0_,t_5__1023_,t_5__1022_,
  t_5__1021_,t_5__1020_,t_5__1019_,t_5__1018_,t_5__1017_,t_5__1016_,t_5__1015_,
  t_5__1014_,t_5__1013_,t_5__1012_,t_5__1011_,t_5__1010_,t_5__1009_,t_5__1008_,
  t_5__1007_,t_5__1006_,t_5__1005_,t_5__1004_,t_5__1003_,t_5__1002_,t_5__1001_,t_5__1000_,
  t_5__999_,t_5__998_,t_5__997_,t_5__996_,t_5__995_,t_5__994_,t_5__993_,t_5__992_,
  t_5__991_,t_5__990_,t_5__989_,t_5__988_,t_5__987_,t_5__986_,t_5__985_,t_5__984_,
  t_5__983_,t_5__982_,t_5__981_,t_5__980_,t_5__979_,t_5__978_,t_5__977_,t_5__976_,
  t_5__975_,t_5__974_,t_5__973_,t_5__972_,t_5__971_,t_5__970_,t_5__969_,t_5__968_,
  t_5__967_,t_5__966_,t_5__965_,t_5__964_,t_5__963_,t_5__962_,t_5__961_,t_5__960_,
  t_5__959_,t_5__958_,t_5__957_,t_5__956_,t_5__955_,t_5__954_,t_5__953_,t_5__952_,
  t_5__951_,t_5__950_,t_5__949_,t_5__948_,t_5__947_,t_5__946_,t_5__945_,t_5__944_,
  t_5__943_,t_5__942_,t_5__941_,t_5__940_,t_5__939_,t_5__938_,t_5__937_,t_5__936_,
  t_5__935_,t_5__934_,t_5__933_,t_5__932_,t_5__931_,t_5__930_,t_5__929_,t_5__928_,
  t_5__927_,t_5__926_,t_5__925_,t_5__924_,t_5__923_,t_5__922_,t_5__921_,t_5__920_,
  t_5__919_,t_5__918_,t_5__917_,t_5__916_,t_5__915_,t_5__914_,t_5__913_,t_5__912_,
  t_5__911_,t_5__910_,t_5__909_,t_5__908_,t_5__907_,t_5__906_,t_5__905_,t_5__904_,
  t_5__903_,t_5__902_,t_5__901_,t_5__900_,t_5__899_,t_5__898_,t_5__897_,t_5__896_,
  t_5__895_,t_5__894_,t_5__893_,t_5__892_,t_5__891_,t_5__890_,t_5__889_,t_5__888_,
  t_5__887_,t_5__886_,t_5__885_,t_5__884_,t_5__883_,t_5__882_,t_5__881_,t_5__880_,
  t_5__879_,t_5__878_,t_5__877_,t_5__876_,t_5__875_,t_5__874_,t_5__873_,t_5__872_,
  t_5__871_,t_5__870_,t_5__869_,t_5__868_,t_5__867_,t_5__866_,t_5__865_,t_5__864_,
  t_5__863_,t_5__862_,t_5__861_,t_5__860_,t_5__859_,t_5__858_,t_5__857_,t_5__856_,
  t_5__855_,t_5__854_,t_5__853_,t_5__852_,t_5__851_,t_5__850_,t_5__849_,t_5__848_,
  t_5__847_,t_5__846_,t_5__845_,t_5__844_,t_5__843_,t_5__842_,t_5__841_,t_5__840_,
  t_5__839_,t_5__838_,t_5__837_,t_5__836_,t_5__835_,t_5__834_,t_5__833_,t_5__832_,
  t_5__831_,t_5__830_,t_5__829_,t_5__828_,t_5__827_,t_5__826_,t_5__825_,t_5__824_,
  t_5__823_,t_5__822_,t_5__821_,t_5__820_,t_5__819_,t_5__818_,t_5__817_,t_5__816_,
  t_5__815_,t_5__814_,t_5__813_,t_5__812_,t_5__811_,t_5__810_,t_5__809_,t_5__808_,
  t_5__807_,t_5__806_,t_5__805_,t_5__804_,t_5__803_,t_5__802_,t_5__801_,t_5__800_,
  t_5__799_,t_5__798_,t_5__797_,t_5__796_,t_5__795_,t_5__794_,t_5__793_,t_5__792_,
  t_5__791_,t_5__790_,t_5__789_,t_5__788_,t_5__787_,t_5__786_,t_5__785_,t_5__784_,
  t_5__783_,t_5__782_,t_5__781_,t_5__780_,t_5__779_,t_5__778_,t_5__777_,t_5__776_,
  t_5__775_,t_5__774_,t_5__773_,t_5__772_,t_5__771_,t_5__770_,t_5__769_,t_5__768_,
  t_5__767_,t_5__766_,t_5__765_,t_5__764_,t_5__763_,t_5__762_,t_5__761_,t_5__760_,
  t_5__759_,t_5__758_,t_5__757_,t_5__756_,t_5__755_,t_5__754_,t_5__753_,t_5__752_,
  t_5__751_,t_5__750_,t_5__749_,t_5__748_,t_5__747_,t_5__746_,t_5__745_,t_5__744_,
  t_5__743_,t_5__742_,t_5__741_,t_5__740_,t_5__739_,t_5__738_,t_5__737_,t_5__736_,
  t_5__735_,t_5__734_,t_5__733_,t_5__732_,t_5__731_,t_5__730_,t_5__729_,t_5__728_,
  t_5__727_,t_5__726_,t_5__725_,t_5__724_,t_5__723_,t_5__722_,t_5__721_,t_5__720_,
  t_5__719_,t_5__718_,t_5__717_,t_5__716_,t_5__715_,t_5__714_,t_5__713_,t_5__712_,
  t_5__711_,t_5__710_,t_5__709_,t_5__708_,t_5__707_,t_5__706_,t_5__705_,t_5__704_,
  t_5__703_,t_5__702_,t_5__701_,t_5__700_,t_5__699_,t_5__698_,t_5__697_,t_5__696_,
  t_5__695_,t_5__694_,t_5__693_,t_5__692_,t_5__691_,t_5__690_,t_5__689_,t_5__688_,
  t_5__687_,t_5__686_,t_5__685_,t_5__684_,t_5__683_,t_5__682_,t_5__681_,t_5__680_,
  t_5__679_,t_5__678_,t_5__677_,t_5__676_,t_5__675_,t_5__674_,t_5__673_,t_5__672_,
  t_5__671_,t_5__670_,t_5__669_,t_5__668_,t_5__667_,t_5__666_,t_5__665_,t_5__664_,
  t_5__663_,t_5__662_,t_5__661_,t_5__660_,t_5__659_,t_5__658_,t_5__657_,t_5__656_,
  t_5__655_,t_5__654_,t_5__653_,t_5__652_,t_5__651_,t_5__650_,t_5__649_,t_5__648_,
  t_5__647_,t_5__646_,t_5__645_,t_5__644_,t_5__643_,t_5__642_,t_5__641_,t_5__640_,
  t_5__639_,t_5__638_,t_5__637_,t_5__636_,t_5__635_,t_5__634_,t_5__633_,t_5__632_,
  t_5__631_,t_5__630_,t_5__629_,t_5__628_,t_5__627_,t_5__626_,t_5__625_,t_5__624_,
  t_5__623_,t_5__622_,t_5__621_,t_5__620_,t_5__619_,t_5__618_,t_5__617_,t_5__616_,
  t_5__615_,t_5__614_,t_5__613_,t_5__612_,t_5__611_,t_5__610_,t_5__609_,t_5__608_,
  t_5__607_,t_5__606_,t_5__605_,t_5__604_,t_5__603_,t_5__602_,t_5__601_,t_5__600_,
  t_5__599_,t_5__598_,t_5__597_,t_5__596_,t_5__595_,t_5__594_,t_5__593_,t_5__592_,
  t_5__591_,t_5__590_,t_5__589_,t_5__588_,t_5__587_,t_5__586_,t_5__585_,t_5__584_,
  t_5__583_,t_5__582_,t_5__581_,t_5__580_,t_5__579_,t_5__578_,t_5__577_,t_5__576_,
  t_5__575_,t_5__574_,t_5__573_,t_5__572_,t_5__571_,t_5__570_,t_5__569_,t_5__568_,
  t_5__567_,t_5__566_,t_5__565_,t_5__564_,t_5__563_,t_5__562_,t_5__561_,t_5__560_,
  t_5__559_,t_5__558_,t_5__557_,t_5__556_,t_5__555_,t_5__554_,t_5__553_,t_5__552_,
  t_5__551_,t_5__550_,t_5__549_,t_5__548_,t_5__547_,t_5__546_,t_5__545_,t_5__544_,
  t_5__543_,t_5__542_,t_5__541_,t_5__540_,t_5__539_,t_5__538_,t_5__537_,t_5__536_,
  t_5__535_,t_5__534_,t_5__533_,t_5__532_,t_5__531_,t_5__530_,t_5__529_,t_5__528_,
  t_5__527_,t_5__526_,t_5__525_,t_5__524_,t_5__523_,t_5__522_,t_5__521_,t_5__520_,
  t_5__519_,t_5__518_,t_5__517_,t_5__516_,t_5__515_,t_5__514_,t_5__513_,t_5__512_,
  t_5__511_,t_5__510_,t_5__509_,t_5__508_,t_5__507_,t_5__506_,t_5__505_,t_5__504_,
  t_5__503_,t_5__502_,t_5__501_,t_5__500_,t_5__499_,t_5__498_,t_5__497_,t_5__496_,
  t_5__495_,t_5__494_,t_5__493_,t_5__492_,t_5__491_,t_5__490_,t_5__489_,t_5__488_,
  t_5__487_,t_5__486_,t_5__485_,t_5__484_,t_5__483_,t_5__482_,t_5__481_,t_5__480_,
  t_5__479_,t_5__478_,t_5__477_,t_5__476_,t_5__475_,t_5__474_,t_5__473_,t_5__472_,
  t_5__471_,t_5__470_,t_5__469_,t_5__468_,t_5__467_,t_5__466_,t_5__465_,t_5__464_,
  t_5__463_,t_5__462_,t_5__461_,t_5__460_,t_5__459_,t_5__458_,t_5__457_,t_5__456_,
  t_5__455_,t_5__454_,t_5__453_,t_5__452_,t_5__451_,t_5__450_,t_5__449_,t_5__448_,
  t_5__447_,t_5__446_,t_5__445_,t_5__444_,t_5__443_,t_5__442_,t_5__441_,t_5__440_,
  t_5__439_,t_5__438_,t_5__437_,t_5__436_,t_5__435_,t_5__434_,t_5__433_,t_5__432_,
  t_5__431_,t_5__430_,t_5__429_,t_5__428_,t_5__427_,t_5__426_,t_5__425_,t_5__424_,
  t_5__423_,t_5__422_,t_5__421_,t_5__420_,t_5__419_,t_5__418_,t_5__417_,t_5__416_,
  t_5__415_,t_5__414_,t_5__413_,t_5__412_,t_5__411_,t_5__410_,t_5__409_,t_5__408_,
  t_5__407_,t_5__406_,t_5__405_,t_5__404_,t_5__403_,t_5__402_,t_5__401_,t_5__400_,
  t_5__399_,t_5__398_,t_5__397_,t_5__396_,t_5__395_,t_5__394_,t_5__393_,t_5__392_,
  t_5__391_,t_5__390_,t_5__389_,t_5__388_,t_5__387_,t_5__386_,t_5__385_,t_5__384_,
  t_5__383_,t_5__382_,t_5__381_,t_5__380_,t_5__379_,t_5__378_,t_5__377_,t_5__376_,
  t_5__375_,t_5__374_,t_5__373_,t_5__372_,t_5__371_,t_5__370_,t_5__369_,t_5__368_,
  t_5__367_,t_5__366_,t_5__365_,t_5__364_,t_5__363_,t_5__362_,t_5__361_,t_5__360_,
  t_5__359_,t_5__358_,t_5__357_,t_5__356_,t_5__355_,t_5__354_,t_5__353_,t_5__352_,
  t_5__351_,t_5__350_,t_5__349_,t_5__348_,t_5__347_,t_5__346_,t_5__345_,t_5__344_,
  t_5__343_,t_5__342_,t_5__341_,t_5__340_,t_5__339_,t_5__338_,t_5__337_,t_5__336_,
  t_5__335_,t_5__334_,t_5__333_,t_5__332_,t_5__331_,t_5__330_,t_5__329_,t_5__328_,
  t_5__327_,t_5__326_,t_5__325_,t_5__324_,t_5__323_,t_5__322_,t_5__321_,t_5__320_,
  t_5__319_,t_5__318_,t_5__317_,t_5__316_,t_5__315_,t_5__314_,t_5__313_,t_5__312_,
  t_5__311_,t_5__310_,t_5__309_,t_5__308_,t_5__307_,t_5__306_,t_5__305_,t_5__304_,
  t_5__303_,t_5__302_,t_5__301_,t_5__300_,t_5__299_,t_5__298_,t_5__297_,t_5__296_,
  t_5__295_,t_5__294_,t_5__293_,t_5__292_,t_5__291_,t_5__290_,t_5__289_,t_5__288_,
  t_5__287_,t_5__286_,t_5__285_,t_5__284_,t_5__283_,t_5__282_,t_5__281_,t_5__280_,
  t_5__279_,t_5__278_,t_5__277_,t_5__276_,t_5__275_,t_5__274_,t_5__273_,t_5__272_,
  t_5__271_,t_5__270_,t_5__269_,t_5__268_,t_5__267_,t_5__266_,t_5__265_,t_5__264_,
  t_5__263_,t_5__262_,t_5__261_,t_5__260_,t_5__259_,t_5__258_,t_5__257_,t_5__256_,
  t_5__255_,t_5__254_,t_5__253_,t_5__252_,t_5__251_,t_5__250_,t_5__249_,t_5__248_,
  t_5__247_,t_5__246_,t_5__245_,t_5__244_,t_5__243_,t_5__242_,t_5__241_,t_5__240_,
  t_5__239_,t_5__238_,t_5__237_,t_5__236_,t_5__235_,t_5__234_,t_5__233_,t_5__232_,
  t_5__231_,t_5__230_,t_5__229_,t_5__228_,t_5__227_,t_5__226_,t_5__225_,t_5__224_,
  t_5__223_,t_5__222_,t_5__221_,t_5__220_,t_5__219_,t_5__218_,t_5__217_,t_5__216_,
  t_5__215_,t_5__214_,t_5__213_,t_5__212_,t_5__211_,t_5__210_,t_5__209_,t_5__208_,
  t_5__207_,t_5__206_,t_5__205_,t_5__204_,t_5__203_,t_5__202_,t_5__201_,t_5__200_,
  t_5__199_,t_5__198_,t_5__197_,t_5__196_,t_5__195_,t_5__194_,t_5__193_,t_5__192_,
  t_5__191_,t_5__190_,t_5__189_,t_5__188_,t_5__187_,t_5__186_,t_5__185_,t_5__184_,
  t_5__183_,t_5__182_,t_5__181_,t_5__180_,t_5__179_,t_5__178_,t_5__177_,t_5__176_,
  t_5__175_,t_5__174_,t_5__173_,t_5__172_,t_5__171_,t_5__170_,t_5__169_,t_5__168_,
  t_5__167_,t_5__166_,t_5__165_,t_5__164_,t_5__163_,t_5__162_,t_5__161_,t_5__160_,
  t_5__159_,t_5__158_,t_5__157_,t_5__156_,t_5__155_,t_5__154_,t_5__153_,t_5__152_,
  t_5__151_,t_5__150_,t_5__149_,t_5__148_,t_5__147_,t_5__146_,t_5__145_,t_5__144_,
  t_5__143_,t_5__142_,t_5__141_,t_5__140_,t_5__139_,t_5__138_,t_5__137_,t_5__136_,
  t_5__135_,t_5__134_,t_5__133_,t_5__132_,t_5__131_,t_5__130_,t_5__129_,t_5__128_,
  t_5__127_,t_5__126_,t_5__125_,t_5__124_,t_5__123_,t_5__122_,t_5__121_,t_5__120_,
  t_5__119_,t_5__118_,t_5__117_,t_5__116_,t_5__115_,t_5__114_,t_5__113_,t_5__112_,
  t_5__111_,t_5__110_,t_5__109_,t_5__108_,t_5__107_,t_5__106_,t_5__105_,t_5__104_,
  t_5__103_,t_5__102_,t_5__101_,t_5__100_,t_5__99_,t_5__98_,t_5__97_,t_5__96_,
  t_5__95_,t_5__94_,t_5__93_,t_5__92_,t_5__91_,t_5__90_,t_5__89_,t_5__88_,t_5__87_,
  t_5__86_,t_5__85_,t_5__84_,t_5__83_,t_5__82_,t_5__81_,t_5__80_,t_5__79_,t_5__78_,
  t_5__77_,t_5__76_,t_5__75_,t_5__74_,t_5__73_,t_5__72_,t_5__71_,t_5__70_,t_5__69_,
  t_5__68_,t_5__67_,t_5__66_,t_5__65_,t_5__64_,t_5__63_,t_5__62_,t_5__61_,t_5__60_,
  t_5__59_,t_5__58_,t_5__57_,t_5__56_,t_5__55_,t_5__54_,t_5__53_,t_5__52_,
  t_5__51_,t_5__50_,t_5__49_,t_5__48_,t_5__47_,t_5__46_,t_5__45_,t_5__44_,t_5__43_,
  t_5__42_,t_5__41_,t_5__40_,t_5__39_,t_5__38_,t_5__37_,t_5__36_,t_5__35_,t_5__34_,
  t_5__33_,t_5__32_,t_5__31_,t_5__30_,t_5__29_,t_5__28_,t_5__27_,t_5__26_,t_5__25_,
  t_5__24_,t_5__23_,t_5__22_,t_5__21_,t_5__20_,t_5__19_,t_5__18_,t_5__17_,t_5__16_,
  t_5__15_,t_5__14_,t_5__13_,t_5__12_,t_5__11_,t_5__10_,t_5__9_,t_5__8_,t_5__7_,
  t_5__6_,t_5__5_,t_5__4_,t_5__3_,t_5__2_,t_5__1_,t_5__0_,t_6__1023_,t_6__1022_,
  t_6__1021_,t_6__1020_,t_6__1019_,t_6__1018_,t_6__1017_,t_6__1016_,t_6__1015_,t_6__1014_,
  t_6__1013_,t_6__1012_,t_6__1011_,t_6__1010_,t_6__1009_,t_6__1008_,t_6__1007_,
  t_6__1006_,t_6__1005_,t_6__1004_,t_6__1003_,t_6__1002_,t_6__1001_,t_6__1000_,
  t_6__999_,t_6__998_,t_6__997_,t_6__996_,t_6__995_,t_6__994_,t_6__993_,t_6__992_,
  t_6__991_,t_6__990_,t_6__989_,t_6__988_,t_6__987_,t_6__986_,t_6__985_,t_6__984_,
  t_6__983_,t_6__982_,t_6__981_,t_6__980_,t_6__979_,t_6__978_,t_6__977_,t_6__976_,
  t_6__975_,t_6__974_,t_6__973_,t_6__972_,t_6__971_,t_6__970_,t_6__969_,t_6__968_,
  t_6__967_,t_6__966_,t_6__965_,t_6__964_,t_6__963_,t_6__962_,t_6__961_,t_6__960_,
  t_6__959_,t_6__958_,t_6__957_,t_6__956_,t_6__955_,t_6__954_,t_6__953_,t_6__952_,
  t_6__951_,t_6__950_,t_6__949_,t_6__948_,t_6__947_,t_6__946_,t_6__945_,t_6__944_,
  t_6__943_,t_6__942_,t_6__941_,t_6__940_,t_6__939_,t_6__938_,t_6__937_,t_6__936_,
  t_6__935_,t_6__934_,t_6__933_,t_6__932_,t_6__931_,t_6__930_,t_6__929_,t_6__928_,
  t_6__927_,t_6__926_,t_6__925_,t_6__924_,t_6__923_,t_6__922_,t_6__921_,t_6__920_,
  t_6__919_,t_6__918_,t_6__917_,t_6__916_,t_6__915_,t_6__914_,t_6__913_,t_6__912_,
  t_6__911_,t_6__910_,t_6__909_,t_6__908_,t_6__907_,t_6__906_,t_6__905_,t_6__904_,
  t_6__903_,t_6__902_,t_6__901_,t_6__900_,t_6__899_,t_6__898_,t_6__897_,t_6__896_,
  t_6__895_,t_6__894_,t_6__893_,t_6__892_,t_6__891_,t_6__890_,t_6__889_,t_6__888_,
  t_6__887_,t_6__886_,t_6__885_,t_6__884_,t_6__883_,t_6__882_,t_6__881_,t_6__880_,
  t_6__879_,t_6__878_,t_6__877_,t_6__876_,t_6__875_,t_6__874_,t_6__873_,t_6__872_,
  t_6__871_,t_6__870_,t_6__869_,t_6__868_,t_6__867_,t_6__866_,t_6__865_,t_6__864_,
  t_6__863_,t_6__862_,t_6__861_,t_6__860_,t_6__859_,t_6__858_,t_6__857_,t_6__856_,
  t_6__855_,t_6__854_,t_6__853_,t_6__852_,t_6__851_,t_6__850_,t_6__849_,t_6__848_,
  t_6__847_,t_6__846_,t_6__845_,t_6__844_,t_6__843_,t_6__842_,t_6__841_,t_6__840_,
  t_6__839_,t_6__838_,t_6__837_,t_6__836_,t_6__835_,t_6__834_,t_6__833_,t_6__832_,
  t_6__831_,t_6__830_,t_6__829_,t_6__828_,t_6__827_,t_6__826_,t_6__825_,t_6__824_,
  t_6__823_,t_6__822_,t_6__821_,t_6__820_,t_6__819_,t_6__818_,t_6__817_,t_6__816_,
  t_6__815_,t_6__814_,t_6__813_,t_6__812_,t_6__811_,t_6__810_,t_6__809_,t_6__808_,
  t_6__807_,t_6__806_,t_6__805_,t_6__804_,t_6__803_,t_6__802_,t_6__801_,t_6__800_,
  t_6__799_,t_6__798_,t_6__797_,t_6__796_,t_6__795_,t_6__794_,t_6__793_,t_6__792_,
  t_6__791_,t_6__790_,t_6__789_,t_6__788_,t_6__787_,t_6__786_,t_6__785_,t_6__784_,
  t_6__783_,t_6__782_,t_6__781_,t_6__780_,t_6__779_,t_6__778_,t_6__777_,t_6__776_,
  t_6__775_,t_6__774_,t_6__773_,t_6__772_,t_6__771_,t_6__770_,t_6__769_,t_6__768_,
  t_6__767_,t_6__766_,t_6__765_,t_6__764_,t_6__763_,t_6__762_,t_6__761_,t_6__760_,
  t_6__759_,t_6__758_,t_6__757_,t_6__756_,t_6__755_,t_6__754_,t_6__753_,t_6__752_,
  t_6__751_,t_6__750_,t_6__749_,t_6__748_,t_6__747_,t_6__746_,t_6__745_,t_6__744_,
  t_6__743_,t_6__742_,t_6__741_,t_6__740_,t_6__739_,t_6__738_,t_6__737_,t_6__736_,
  t_6__735_,t_6__734_,t_6__733_,t_6__732_,t_6__731_,t_6__730_,t_6__729_,t_6__728_,
  t_6__727_,t_6__726_,t_6__725_,t_6__724_,t_6__723_,t_6__722_,t_6__721_,t_6__720_,
  t_6__719_,t_6__718_,t_6__717_,t_6__716_,t_6__715_,t_6__714_,t_6__713_,t_6__712_,
  t_6__711_,t_6__710_,t_6__709_,t_6__708_,t_6__707_,t_6__706_,t_6__705_,t_6__704_,
  t_6__703_,t_6__702_,t_6__701_,t_6__700_,t_6__699_,t_6__698_,t_6__697_,t_6__696_,
  t_6__695_,t_6__694_,t_6__693_,t_6__692_,t_6__691_,t_6__690_,t_6__689_,t_6__688_,
  t_6__687_,t_6__686_,t_6__685_,t_6__684_,t_6__683_,t_6__682_,t_6__681_,t_6__680_,
  t_6__679_,t_6__678_,t_6__677_,t_6__676_,t_6__675_,t_6__674_,t_6__673_,t_6__672_,
  t_6__671_,t_6__670_,t_6__669_,t_6__668_,t_6__667_,t_6__666_,t_6__665_,t_6__664_,
  t_6__663_,t_6__662_,t_6__661_,t_6__660_,t_6__659_,t_6__658_,t_6__657_,t_6__656_,
  t_6__655_,t_6__654_,t_6__653_,t_6__652_,t_6__651_,t_6__650_,t_6__649_,t_6__648_,
  t_6__647_,t_6__646_,t_6__645_,t_6__644_,t_6__643_,t_6__642_,t_6__641_,t_6__640_,
  t_6__639_,t_6__638_,t_6__637_,t_6__636_,t_6__635_,t_6__634_,t_6__633_,t_6__632_,
  t_6__631_,t_6__630_,t_6__629_,t_6__628_,t_6__627_,t_6__626_,t_6__625_,t_6__624_,
  t_6__623_,t_6__622_,t_6__621_,t_6__620_,t_6__619_,t_6__618_,t_6__617_,t_6__616_,
  t_6__615_,t_6__614_,t_6__613_,t_6__612_,t_6__611_,t_6__610_,t_6__609_,t_6__608_,
  t_6__607_,t_6__606_,t_6__605_,t_6__604_,t_6__603_,t_6__602_,t_6__601_,t_6__600_,
  t_6__599_,t_6__598_,t_6__597_,t_6__596_,t_6__595_,t_6__594_,t_6__593_,t_6__592_,
  t_6__591_,t_6__590_,t_6__589_,t_6__588_,t_6__587_,t_6__586_,t_6__585_,t_6__584_,
  t_6__583_,t_6__582_,t_6__581_,t_6__580_,t_6__579_,t_6__578_,t_6__577_,t_6__576_,
  t_6__575_,t_6__574_,t_6__573_,t_6__572_,t_6__571_,t_6__570_,t_6__569_,t_6__568_,
  t_6__567_,t_6__566_,t_6__565_,t_6__564_,t_6__563_,t_6__562_,t_6__561_,t_6__560_,
  t_6__559_,t_6__558_,t_6__557_,t_6__556_,t_6__555_,t_6__554_,t_6__553_,t_6__552_,
  t_6__551_,t_6__550_,t_6__549_,t_6__548_,t_6__547_,t_6__546_,t_6__545_,t_6__544_,
  t_6__543_,t_6__542_,t_6__541_,t_6__540_,t_6__539_,t_6__538_,t_6__537_,t_6__536_,
  t_6__535_,t_6__534_,t_6__533_,t_6__532_,t_6__531_,t_6__530_,t_6__529_,t_6__528_,
  t_6__527_,t_6__526_,t_6__525_,t_6__524_,t_6__523_,t_6__522_,t_6__521_,t_6__520_,
  t_6__519_,t_6__518_,t_6__517_,t_6__516_,t_6__515_,t_6__514_,t_6__513_,t_6__512_,
  t_6__511_,t_6__510_,t_6__509_,t_6__508_,t_6__507_,t_6__506_,t_6__505_,t_6__504_,
  t_6__503_,t_6__502_,t_6__501_,t_6__500_,t_6__499_,t_6__498_,t_6__497_,t_6__496_,
  t_6__495_,t_6__494_,t_6__493_,t_6__492_,t_6__491_,t_6__490_,t_6__489_,t_6__488_,
  t_6__487_,t_6__486_,t_6__485_,t_6__484_,t_6__483_,t_6__482_,t_6__481_,t_6__480_,
  t_6__479_,t_6__478_,t_6__477_,t_6__476_,t_6__475_,t_6__474_,t_6__473_,t_6__472_,
  t_6__471_,t_6__470_,t_6__469_,t_6__468_,t_6__467_,t_6__466_,t_6__465_,t_6__464_,
  t_6__463_,t_6__462_,t_6__461_,t_6__460_,t_6__459_,t_6__458_,t_6__457_,t_6__456_,
  t_6__455_,t_6__454_,t_6__453_,t_6__452_,t_6__451_,t_6__450_,t_6__449_,t_6__448_,
  t_6__447_,t_6__446_,t_6__445_,t_6__444_,t_6__443_,t_6__442_,t_6__441_,t_6__440_,
  t_6__439_,t_6__438_,t_6__437_,t_6__436_,t_6__435_,t_6__434_,t_6__433_,t_6__432_,
  t_6__431_,t_6__430_,t_6__429_,t_6__428_,t_6__427_,t_6__426_,t_6__425_,t_6__424_,
  t_6__423_,t_6__422_,t_6__421_,t_6__420_,t_6__419_,t_6__418_,t_6__417_,t_6__416_,
  t_6__415_,t_6__414_,t_6__413_,t_6__412_,t_6__411_,t_6__410_,t_6__409_,t_6__408_,
  t_6__407_,t_6__406_,t_6__405_,t_6__404_,t_6__403_,t_6__402_,t_6__401_,t_6__400_,
  t_6__399_,t_6__398_,t_6__397_,t_6__396_,t_6__395_,t_6__394_,t_6__393_,t_6__392_,
  t_6__391_,t_6__390_,t_6__389_,t_6__388_,t_6__387_,t_6__386_,t_6__385_,t_6__384_,
  t_6__383_,t_6__382_,t_6__381_,t_6__380_,t_6__379_,t_6__378_,t_6__377_,t_6__376_,
  t_6__375_,t_6__374_,t_6__373_,t_6__372_,t_6__371_,t_6__370_,t_6__369_,t_6__368_,
  t_6__367_,t_6__366_,t_6__365_,t_6__364_,t_6__363_,t_6__362_,t_6__361_,t_6__360_,
  t_6__359_,t_6__358_,t_6__357_,t_6__356_,t_6__355_,t_6__354_,t_6__353_,t_6__352_,
  t_6__351_,t_6__350_,t_6__349_,t_6__348_,t_6__347_,t_6__346_,t_6__345_,t_6__344_,
  t_6__343_,t_6__342_,t_6__341_,t_6__340_,t_6__339_,t_6__338_,t_6__337_,t_6__336_,
  t_6__335_,t_6__334_,t_6__333_,t_6__332_,t_6__331_,t_6__330_,t_6__329_,t_6__328_,
  t_6__327_,t_6__326_,t_6__325_,t_6__324_,t_6__323_,t_6__322_,t_6__321_,t_6__320_,
  t_6__319_,t_6__318_,t_6__317_,t_6__316_,t_6__315_,t_6__314_,t_6__313_,t_6__312_,
  t_6__311_,t_6__310_,t_6__309_,t_6__308_,t_6__307_,t_6__306_,t_6__305_,t_6__304_,
  t_6__303_,t_6__302_,t_6__301_,t_6__300_,t_6__299_,t_6__298_,t_6__297_,t_6__296_,
  t_6__295_,t_6__294_,t_6__293_,t_6__292_,t_6__291_,t_6__290_,t_6__289_,t_6__288_,
  t_6__287_,t_6__286_,t_6__285_,t_6__284_,t_6__283_,t_6__282_,t_6__281_,t_6__280_,
  t_6__279_,t_6__278_,t_6__277_,t_6__276_,t_6__275_,t_6__274_,t_6__273_,t_6__272_,
  t_6__271_,t_6__270_,t_6__269_,t_6__268_,t_6__267_,t_6__266_,t_6__265_,t_6__264_,
  t_6__263_,t_6__262_,t_6__261_,t_6__260_,t_6__259_,t_6__258_,t_6__257_,t_6__256_,
  t_6__255_,t_6__254_,t_6__253_,t_6__252_,t_6__251_,t_6__250_,t_6__249_,t_6__248_,
  t_6__247_,t_6__246_,t_6__245_,t_6__244_,t_6__243_,t_6__242_,t_6__241_,t_6__240_,
  t_6__239_,t_6__238_,t_6__237_,t_6__236_,t_6__235_,t_6__234_,t_6__233_,t_6__232_,
  t_6__231_,t_6__230_,t_6__229_,t_6__228_,t_6__227_,t_6__226_,t_6__225_,t_6__224_,
  t_6__223_,t_6__222_,t_6__221_,t_6__220_,t_6__219_,t_6__218_,t_6__217_,t_6__216_,
  t_6__215_,t_6__214_,t_6__213_,t_6__212_,t_6__211_,t_6__210_,t_6__209_,t_6__208_,
  t_6__207_,t_6__206_,t_6__205_,t_6__204_,t_6__203_,t_6__202_,t_6__201_,t_6__200_,
  t_6__199_,t_6__198_,t_6__197_,t_6__196_,t_6__195_,t_6__194_,t_6__193_,t_6__192_,
  t_6__191_,t_6__190_,t_6__189_,t_6__188_,t_6__187_,t_6__186_,t_6__185_,t_6__184_,
  t_6__183_,t_6__182_,t_6__181_,t_6__180_,t_6__179_,t_6__178_,t_6__177_,t_6__176_,
  t_6__175_,t_6__174_,t_6__173_,t_6__172_,t_6__171_,t_6__170_,t_6__169_,t_6__168_,
  t_6__167_,t_6__166_,t_6__165_,t_6__164_,t_6__163_,t_6__162_,t_6__161_,t_6__160_,
  t_6__159_,t_6__158_,t_6__157_,t_6__156_,t_6__155_,t_6__154_,t_6__153_,t_6__152_,
  t_6__151_,t_6__150_,t_6__149_,t_6__148_,t_6__147_,t_6__146_,t_6__145_,t_6__144_,
  t_6__143_,t_6__142_,t_6__141_,t_6__140_,t_6__139_,t_6__138_,t_6__137_,t_6__136_,
  t_6__135_,t_6__134_,t_6__133_,t_6__132_,t_6__131_,t_6__130_,t_6__129_,t_6__128_,
  t_6__127_,t_6__126_,t_6__125_,t_6__124_,t_6__123_,t_6__122_,t_6__121_,t_6__120_,
  t_6__119_,t_6__118_,t_6__117_,t_6__116_,t_6__115_,t_6__114_,t_6__113_,t_6__112_,
  t_6__111_,t_6__110_,t_6__109_,t_6__108_,t_6__107_,t_6__106_,t_6__105_,t_6__104_,
  t_6__103_,t_6__102_,t_6__101_,t_6__100_,t_6__99_,t_6__98_,t_6__97_,t_6__96_,t_6__95_,
  t_6__94_,t_6__93_,t_6__92_,t_6__91_,t_6__90_,t_6__89_,t_6__88_,t_6__87_,t_6__86_,
  t_6__85_,t_6__84_,t_6__83_,t_6__82_,t_6__81_,t_6__80_,t_6__79_,t_6__78_,
  t_6__77_,t_6__76_,t_6__75_,t_6__74_,t_6__73_,t_6__72_,t_6__71_,t_6__70_,t_6__69_,
  t_6__68_,t_6__67_,t_6__66_,t_6__65_,t_6__64_,t_6__63_,t_6__62_,t_6__61_,t_6__60_,
  t_6__59_,t_6__58_,t_6__57_,t_6__56_,t_6__55_,t_6__54_,t_6__53_,t_6__52_,t_6__51_,
  t_6__50_,t_6__49_,t_6__48_,t_6__47_,t_6__46_,t_6__45_,t_6__44_,t_6__43_,t_6__42_,
  t_6__41_,t_6__40_,t_6__39_,t_6__38_,t_6__37_,t_6__36_,t_6__35_,t_6__34_,t_6__33_,
  t_6__32_,t_6__31_,t_6__30_,t_6__29_,t_6__28_,t_6__27_,t_6__26_,t_6__25_,t_6__24_,
  t_6__23_,t_6__22_,t_6__21_,t_6__20_,t_6__19_,t_6__18_,t_6__17_,t_6__16_,t_6__15_,
  t_6__14_,t_6__13_,t_6__12_,t_6__11_,t_6__10_,t_6__9_,t_6__8_,t_6__7_,t_6__6_,
  t_6__5_,t_6__4_,t_6__3_,t_6__2_,t_6__1_,t_6__0_,t_7__1023_,t_7__1022_,t_7__1021_,
  t_7__1020_,t_7__1019_,t_7__1018_,t_7__1017_,t_7__1016_,t_7__1015_,t_7__1014_,
  t_7__1013_,t_7__1012_,t_7__1011_,t_7__1010_,t_7__1009_,t_7__1008_,t_7__1007_,
  t_7__1006_,t_7__1005_,t_7__1004_,t_7__1003_,t_7__1002_,t_7__1001_,t_7__1000_,t_7__999_,
  t_7__998_,t_7__997_,t_7__996_,t_7__995_,t_7__994_,t_7__993_,t_7__992_,t_7__991_,
  t_7__990_,t_7__989_,t_7__988_,t_7__987_,t_7__986_,t_7__985_,t_7__984_,t_7__983_,
  t_7__982_,t_7__981_,t_7__980_,t_7__979_,t_7__978_,t_7__977_,t_7__976_,t_7__975_,
  t_7__974_,t_7__973_,t_7__972_,t_7__971_,t_7__970_,t_7__969_,t_7__968_,t_7__967_,
  t_7__966_,t_7__965_,t_7__964_,t_7__963_,t_7__962_,t_7__961_,t_7__960_,t_7__959_,
  t_7__958_,t_7__957_,t_7__956_,t_7__955_,t_7__954_,t_7__953_,t_7__952_,t_7__951_,
  t_7__950_,t_7__949_,t_7__948_,t_7__947_,t_7__946_,t_7__945_,t_7__944_,t_7__943_,
  t_7__942_,t_7__941_,t_7__940_,t_7__939_,t_7__938_,t_7__937_,t_7__936_,t_7__935_,
  t_7__934_,t_7__933_,t_7__932_,t_7__931_,t_7__930_,t_7__929_,t_7__928_,t_7__927_,
  t_7__926_,t_7__925_,t_7__924_,t_7__923_,t_7__922_,t_7__921_,t_7__920_,t_7__919_,
  t_7__918_,t_7__917_,t_7__916_,t_7__915_,t_7__914_,t_7__913_,t_7__912_,t_7__911_,
  t_7__910_,t_7__909_,t_7__908_,t_7__907_,t_7__906_,t_7__905_,t_7__904_,t_7__903_,
  t_7__902_,t_7__901_,t_7__900_,t_7__899_,t_7__898_,t_7__897_,t_7__896_,t_7__895_,
  t_7__894_,t_7__893_,t_7__892_,t_7__891_,t_7__890_,t_7__889_,t_7__888_,t_7__887_,
  t_7__886_,t_7__885_,t_7__884_,t_7__883_,t_7__882_,t_7__881_,t_7__880_,t_7__879_,
  t_7__878_,t_7__877_,t_7__876_,t_7__875_,t_7__874_,t_7__873_,t_7__872_,t_7__871_,
  t_7__870_,t_7__869_,t_7__868_,t_7__867_,t_7__866_,t_7__865_,t_7__864_,t_7__863_,
  t_7__862_,t_7__861_,t_7__860_,t_7__859_,t_7__858_,t_7__857_,t_7__856_,t_7__855_,
  t_7__854_,t_7__853_,t_7__852_,t_7__851_,t_7__850_,t_7__849_,t_7__848_,t_7__847_,
  t_7__846_,t_7__845_,t_7__844_,t_7__843_,t_7__842_,t_7__841_,t_7__840_,t_7__839_,
  t_7__838_,t_7__837_,t_7__836_,t_7__835_,t_7__834_,t_7__833_,t_7__832_,t_7__831_,
  t_7__830_,t_7__829_,t_7__828_,t_7__827_,t_7__826_,t_7__825_,t_7__824_,t_7__823_,
  t_7__822_,t_7__821_,t_7__820_,t_7__819_,t_7__818_,t_7__817_,t_7__816_,t_7__815_,
  t_7__814_,t_7__813_,t_7__812_,t_7__811_,t_7__810_,t_7__809_,t_7__808_,t_7__807_,
  t_7__806_,t_7__805_,t_7__804_,t_7__803_,t_7__802_,t_7__801_,t_7__800_,t_7__799_,
  t_7__798_,t_7__797_,t_7__796_,t_7__795_,t_7__794_,t_7__793_,t_7__792_,t_7__791_,
  t_7__790_,t_7__789_,t_7__788_,t_7__787_,t_7__786_,t_7__785_,t_7__784_,t_7__783_,
  t_7__782_,t_7__781_,t_7__780_,t_7__779_,t_7__778_,t_7__777_,t_7__776_,t_7__775_,
  t_7__774_,t_7__773_,t_7__772_,t_7__771_,t_7__770_,t_7__769_,t_7__768_,t_7__767_,
  t_7__766_,t_7__765_,t_7__764_,t_7__763_,t_7__762_,t_7__761_,t_7__760_,t_7__759_,
  t_7__758_,t_7__757_,t_7__756_,t_7__755_,t_7__754_,t_7__753_,t_7__752_,t_7__751_,
  t_7__750_,t_7__749_,t_7__748_,t_7__747_,t_7__746_,t_7__745_,t_7__744_,t_7__743_,
  t_7__742_,t_7__741_,t_7__740_,t_7__739_,t_7__738_,t_7__737_,t_7__736_,t_7__735_,
  t_7__734_,t_7__733_,t_7__732_,t_7__731_,t_7__730_,t_7__729_,t_7__728_,t_7__727_,
  t_7__726_,t_7__725_,t_7__724_,t_7__723_,t_7__722_,t_7__721_,t_7__720_,t_7__719_,
  t_7__718_,t_7__717_,t_7__716_,t_7__715_,t_7__714_,t_7__713_,t_7__712_,t_7__711_,
  t_7__710_,t_7__709_,t_7__708_,t_7__707_,t_7__706_,t_7__705_,t_7__704_,t_7__703_,
  t_7__702_,t_7__701_,t_7__700_,t_7__699_,t_7__698_,t_7__697_,t_7__696_,t_7__695_,
  t_7__694_,t_7__693_,t_7__692_,t_7__691_,t_7__690_,t_7__689_,t_7__688_,t_7__687_,
  t_7__686_,t_7__685_,t_7__684_,t_7__683_,t_7__682_,t_7__681_,t_7__680_,t_7__679_,
  t_7__678_,t_7__677_,t_7__676_,t_7__675_,t_7__674_,t_7__673_,t_7__672_,t_7__671_,
  t_7__670_,t_7__669_,t_7__668_,t_7__667_,t_7__666_,t_7__665_,t_7__664_,t_7__663_,
  t_7__662_,t_7__661_,t_7__660_,t_7__659_,t_7__658_,t_7__657_,t_7__656_,t_7__655_,
  t_7__654_,t_7__653_,t_7__652_,t_7__651_,t_7__650_,t_7__649_,t_7__648_,t_7__647_,
  t_7__646_,t_7__645_,t_7__644_,t_7__643_,t_7__642_,t_7__641_,t_7__640_,t_7__639_,
  t_7__638_,t_7__637_,t_7__636_,t_7__635_,t_7__634_,t_7__633_,t_7__632_,t_7__631_,
  t_7__630_,t_7__629_,t_7__628_,t_7__627_,t_7__626_,t_7__625_,t_7__624_,t_7__623_,
  t_7__622_,t_7__621_,t_7__620_,t_7__619_,t_7__618_,t_7__617_,t_7__616_,t_7__615_,
  t_7__614_,t_7__613_,t_7__612_,t_7__611_,t_7__610_,t_7__609_,t_7__608_,t_7__607_,
  t_7__606_,t_7__605_,t_7__604_,t_7__603_,t_7__602_,t_7__601_,t_7__600_,t_7__599_,
  t_7__598_,t_7__597_,t_7__596_,t_7__595_,t_7__594_,t_7__593_,t_7__592_,t_7__591_,
  t_7__590_,t_7__589_,t_7__588_,t_7__587_,t_7__586_,t_7__585_,t_7__584_,t_7__583_,
  t_7__582_,t_7__581_,t_7__580_,t_7__579_,t_7__578_,t_7__577_,t_7__576_,t_7__575_,
  t_7__574_,t_7__573_,t_7__572_,t_7__571_,t_7__570_,t_7__569_,t_7__568_,t_7__567_,
  t_7__566_,t_7__565_,t_7__564_,t_7__563_,t_7__562_,t_7__561_,t_7__560_,t_7__559_,
  t_7__558_,t_7__557_,t_7__556_,t_7__555_,t_7__554_,t_7__553_,t_7__552_,t_7__551_,
  t_7__550_,t_7__549_,t_7__548_,t_7__547_,t_7__546_,t_7__545_,t_7__544_,t_7__543_,
  t_7__542_,t_7__541_,t_7__540_,t_7__539_,t_7__538_,t_7__537_,t_7__536_,t_7__535_,
  t_7__534_,t_7__533_,t_7__532_,t_7__531_,t_7__530_,t_7__529_,t_7__528_,t_7__527_,
  t_7__526_,t_7__525_,t_7__524_,t_7__523_,t_7__522_,t_7__521_,t_7__520_,t_7__519_,
  t_7__518_,t_7__517_,t_7__516_,t_7__515_,t_7__514_,t_7__513_,t_7__512_,t_7__511_,
  t_7__510_,t_7__509_,t_7__508_,t_7__507_,t_7__506_,t_7__505_,t_7__504_,t_7__503_,
  t_7__502_,t_7__501_,t_7__500_,t_7__499_,t_7__498_,t_7__497_,t_7__496_,t_7__495_,
  t_7__494_,t_7__493_,t_7__492_,t_7__491_,t_7__490_,t_7__489_,t_7__488_,t_7__487_,
  t_7__486_,t_7__485_,t_7__484_,t_7__483_,t_7__482_,t_7__481_,t_7__480_,t_7__479_,
  t_7__478_,t_7__477_,t_7__476_,t_7__475_,t_7__474_,t_7__473_,t_7__472_,t_7__471_,
  t_7__470_,t_7__469_,t_7__468_,t_7__467_,t_7__466_,t_7__465_,t_7__464_,t_7__463_,
  t_7__462_,t_7__461_,t_7__460_,t_7__459_,t_7__458_,t_7__457_,t_7__456_,t_7__455_,
  t_7__454_,t_7__453_,t_7__452_,t_7__451_,t_7__450_,t_7__449_,t_7__448_,t_7__447_,
  t_7__446_,t_7__445_,t_7__444_,t_7__443_,t_7__442_,t_7__441_,t_7__440_,t_7__439_,
  t_7__438_,t_7__437_,t_7__436_,t_7__435_,t_7__434_,t_7__433_,t_7__432_,t_7__431_,
  t_7__430_,t_7__429_,t_7__428_,t_7__427_,t_7__426_,t_7__425_,t_7__424_,t_7__423_,
  t_7__422_,t_7__421_,t_7__420_,t_7__419_,t_7__418_,t_7__417_,t_7__416_,t_7__415_,
  t_7__414_,t_7__413_,t_7__412_,t_7__411_,t_7__410_,t_7__409_,t_7__408_,t_7__407_,
  t_7__406_,t_7__405_,t_7__404_,t_7__403_,t_7__402_,t_7__401_,t_7__400_,t_7__399_,
  t_7__398_,t_7__397_,t_7__396_,t_7__395_,t_7__394_,t_7__393_,t_7__392_,t_7__391_,
  t_7__390_,t_7__389_,t_7__388_,t_7__387_,t_7__386_,t_7__385_,t_7__384_,t_7__383_,
  t_7__382_,t_7__381_,t_7__380_,t_7__379_,t_7__378_,t_7__377_,t_7__376_,t_7__375_,
  t_7__374_,t_7__373_,t_7__372_,t_7__371_,t_7__370_,t_7__369_,t_7__368_,t_7__367_,
  t_7__366_,t_7__365_,t_7__364_,t_7__363_,t_7__362_,t_7__361_,t_7__360_,t_7__359_,
  t_7__358_,t_7__357_,t_7__356_,t_7__355_,t_7__354_,t_7__353_,t_7__352_,t_7__351_,
  t_7__350_,t_7__349_,t_7__348_,t_7__347_,t_7__346_,t_7__345_,t_7__344_,t_7__343_,
  t_7__342_,t_7__341_,t_7__340_,t_7__339_,t_7__338_,t_7__337_,t_7__336_,t_7__335_,
  t_7__334_,t_7__333_,t_7__332_,t_7__331_,t_7__330_,t_7__329_,t_7__328_,t_7__327_,
  t_7__326_,t_7__325_,t_7__324_,t_7__323_,t_7__322_,t_7__321_,t_7__320_,t_7__319_,
  t_7__318_,t_7__317_,t_7__316_,t_7__315_,t_7__314_,t_7__313_,t_7__312_,t_7__311_,
  t_7__310_,t_7__309_,t_7__308_,t_7__307_,t_7__306_,t_7__305_,t_7__304_,t_7__303_,
  t_7__302_,t_7__301_,t_7__300_,t_7__299_,t_7__298_,t_7__297_,t_7__296_,t_7__295_,
  t_7__294_,t_7__293_,t_7__292_,t_7__291_,t_7__290_,t_7__289_,t_7__288_,t_7__287_,
  t_7__286_,t_7__285_,t_7__284_,t_7__283_,t_7__282_,t_7__281_,t_7__280_,t_7__279_,
  t_7__278_,t_7__277_,t_7__276_,t_7__275_,t_7__274_,t_7__273_,t_7__272_,t_7__271_,
  t_7__270_,t_7__269_,t_7__268_,t_7__267_,t_7__266_,t_7__265_,t_7__264_,t_7__263_,
  t_7__262_,t_7__261_,t_7__260_,t_7__259_,t_7__258_,t_7__257_,t_7__256_,t_7__255_,
  t_7__254_,t_7__253_,t_7__252_,t_7__251_,t_7__250_,t_7__249_,t_7__248_,t_7__247_,
  t_7__246_,t_7__245_,t_7__244_,t_7__243_,t_7__242_,t_7__241_,t_7__240_,t_7__239_,
  t_7__238_,t_7__237_,t_7__236_,t_7__235_,t_7__234_,t_7__233_,t_7__232_,t_7__231_,
  t_7__230_,t_7__229_,t_7__228_,t_7__227_,t_7__226_,t_7__225_,t_7__224_,t_7__223_,
  t_7__222_,t_7__221_,t_7__220_,t_7__219_,t_7__218_,t_7__217_,t_7__216_,t_7__215_,
  t_7__214_,t_7__213_,t_7__212_,t_7__211_,t_7__210_,t_7__209_,t_7__208_,t_7__207_,
  t_7__206_,t_7__205_,t_7__204_,t_7__203_,t_7__202_,t_7__201_,t_7__200_,t_7__199_,
  t_7__198_,t_7__197_,t_7__196_,t_7__195_,t_7__194_,t_7__193_,t_7__192_,t_7__191_,
  t_7__190_,t_7__189_,t_7__188_,t_7__187_,t_7__186_,t_7__185_,t_7__184_,t_7__183_,
  t_7__182_,t_7__181_,t_7__180_,t_7__179_,t_7__178_,t_7__177_,t_7__176_,t_7__175_,
  t_7__174_,t_7__173_,t_7__172_,t_7__171_,t_7__170_,t_7__169_,t_7__168_,t_7__167_,
  t_7__166_,t_7__165_,t_7__164_,t_7__163_,t_7__162_,t_7__161_,t_7__160_,t_7__159_,
  t_7__158_,t_7__157_,t_7__156_,t_7__155_,t_7__154_,t_7__153_,t_7__152_,t_7__151_,
  t_7__150_,t_7__149_,t_7__148_,t_7__147_,t_7__146_,t_7__145_,t_7__144_,t_7__143_,
  t_7__142_,t_7__141_,t_7__140_,t_7__139_,t_7__138_,t_7__137_,t_7__136_,t_7__135_,
  t_7__134_,t_7__133_,t_7__132_,t_7__131_,t_7__130_,t_7__129_,t_7__128_,t_7__127_,
  t_7__126_,t_7__125_,t_7__124_,t_7__123_,t_7__122_,t_7__121_,t_7__120_,t_7__119_,
  t_7__118_,t_7__117_,t_7__116_,t_7__115_,t_7__114_,t_7__113_,t_7__112_,t_7__111_,
  t_7__110_,t_7__109_,t_7__108_,t_7__107_,t_7__106_,t_7__105_,t_7__104_,t_7__103_,
  t_7__102_,t_7__101_,t_7__100_,t_7__99_,t_7__98_,t_7__97_,t_7__96_,t_7__95_,
  t_7__94_,t_7__93_,t_7__92_,t_7__91_,t_7__90_,t_7__89_,t_7__88_,t_7__87_,t_7__86_,
  t_7__85_,t_7__84_,t_7__83_,t_7__82_,t_7__81_,t_7__80_,t_7__79_,t_7__78_,t_7__77_,
  t_7__76_,t_7__75_,t_7__74_,t_7__73_,t_7__72_,t_7__71_,t_7__70_,t_7__69_,t_7__68_,
  t_7__67_,t_7__66_,t_7__65_,t_7__64_,t_7__63_,t_7__62_,t_7__61_,t_7__60_,t_7__59_,
  t_7__58_,t_7__57_,t_7__56_,t_7__55_,t_7__54_,t_7__53_,t_7__52_,t_7__51_,t_7__50_,
  t_7__49_,t_7__48_,t_7__47_,t_7__46_,t_7__45_,t_7__44_,t_7__43_,t_7__42_,t_7__41_,
  t_7__40_,t_7__39_,t_7__38_,t_7__37_,t_7__36_,t_7__35_,t_7__34_,t_7__33_,t_7__32_,
  t_7__31_,t_7__30_,t_7__29_,t_7__28_,t_7__27_,t_7__26_,t_7__25_,t_7__24_,
  t_7__23_,t_7__22_,t_7__21_,t_7__20_,t_7__19_,t_7__18_,t_7__17_,t_7__16_,t_7__15_,
  t_7__14_,t_7__13_,t_7__12_,t_7__11_,t_7__10_,t_7__9_,t_7__8_,t_7__7_,t_7__6_,t_7__5_,
  t_7__4_,t_7__3_,t_7__2_,t_7__1_,t_7__0_,t_8__1023_,t_8__1022_,t_8__1021_,
  t_8__1020_,t_8__1019_,t_8__1018_,t_8__1017_,t_8__1016_,t_8__1015_,t_8__1014_,t_8__1013_,
  t_8__1012_,t_8__1011_,t_8__1010_,t_8__1009_,t_8__1008_,t_8__1007_,t_8__1006_,
  t_8__1005_,t_8__1004_,t_8__1003_,t_8__1002_,t_8__1001_,t_8__1000_,t_8__999_,
  t_8__998_,t_8__997_,t_8__996_,t_8__995_,t_8__994_,t_8__993_,t_8__992_,t_8__991_,
  t_8__990_,t_8__989_,t_8__988_,t_8__987_,t_8__986_,t_8__985_,t_8__984_,t_8__983_,
  t_8__982_,t_8__981_,t_8__980_,t_8__979_,t_8__978_,t_8__977_,t_8__976_,t_8__975_,
  t_8__974_,t_8__973_,t_8__972_,t_8__971_,t_8__970_,t_8__969_,t_8__968_,t_8__967_,
  t_8__966_,t_8__965_,t_8__964_,t_8__963_,t_8__962_,t_8__961_,t_8__960_,t_8__959_,
  t_8__958_,t_8__957_,t_8__956_,t_8__955_,t_8__954_,t_8__953_,t_8__952_,t_8__951_,
  t_8__950_,t_8__949_,t_8__948_,t_8__947_,t_8__946_,t_8__945_,t_8__944_,t_8__943_,
  t_8__942_,t_8__941_,t_8__940_,t_8__939_,t_8__938_,t_8__937_,t_8__936_,t_8__935_,
  t_8__934_,t_8__933_,t_8__932_,t_8__931_,t_8__930_,t_8__929_,t_8__928_,t_8__927_,
  t_8__926_,t_8__925_,t_8__924_,t_8__923_,t_8__922_,t_8__921_,t_8__920_,t_8__919_,
  t_8__918_,t_8__917_,t_8__916_,t_8__915_,t_8__914_,t_8__913_,t_8__912_,t_8__911_,
  t_8__910_,t_8__909_,t_8__908_,t_8__907_,t_8__906_,t_8__905_,t_8__904_,t_8__903_,
  t_8__902_,t_8__901_,t_8__900_,t_8__899_,t_8__898_,t_8__897_,t_8__896_,t_8__895_,
  t_8__894_,t_8__893_,t_8__892_,t_8__891_,t_8__890_,t_8__889_,t_8__888_,t_8__887_,
  t_8__886_,t_8__885_,t_8__884_,t_8__883_,t_8__882_,t_8__881_,t_8__880_,t_8__879_,
  t_8__878_,t_8__877_,t_8__876_,t_8__875_,t_8__874_,t_8__873_,t_8__872_,t_8__871_,
  t_8__870_,t_8__869_,t_8__868_,t_8__867_,t_8__866_,t_8__865_,t_8__864_,t_8__863_,
  t_8__862_,t_8__861_,t_8__860_,t_8__859_,t_8__858_,t_8__857_,t_8__856_,t_8__855_,
  t_8__854_,t_8__853_,t_8__852_,t_8__851_,t_8__850_,t_8__849_,t_8__848_,t_8__847_,
  t_8__846_,t_8__845_,t_8__844_,t_8__843_,t_8__842_,t_8__841_,t_8__840_,t_8__839_,
  t_8__838_,t_8__837_,t_8__836_,t_8__835_,t_8__834_,t_8__833_,t_8__832_,t_8__831_,
  t_8__830_,t_8__829_,t_8__828_,t_8__827_,t_8__826_,t_8__825_,t_8__824_,t_8__823_,
  t_8__822_,t_8__821_,t_8__820_,t_8__819_,t_8__818_,t_8__817_,t_8__816_,t_8__815_,
  t_8__814_,t_8__813_,t_8__812_,t_8__811_,t_8__810_,t_8__809_,t_8__808_,t_8__807_,
  t_8__806_,t_8__805_,t_8__804_,t_8__803_,t_8__802_,t_8__801_,t_8__800_,t_8__799_,
  t_8__798_,t_8__797_,t_8__796_,t_8__795_,t_8__794_,t_8__793_,t_8__792_,t_8__791_,
  t_8__790_,t_8__789_,t_8__788_,t_8__787_,t_8__786_,t_8__785_,t_8__784_,t_8__783_,
  t_8__782_,t_8__781_,t_8__780_,t_8__779_,t_8__778_,t_8__777_,t_8__776_,t_8__775_,
  t_8__774_,t_8__773_,t_8__772_,t_8__771_,t_8__770_,t_8__769_,t_8__768_,t_8__767_,
  t_8__766_,t_8__765_,t_8__764_,t_8__763_,t_8__762_,t_8__761_,t_8__760_,t_8__759_,
  t_8__758_,t_8__757_,t_8__756_,t_8__755_,t_8__754_,t_8__753_,t_8__752_,t_8__751_,
  t_8__750_,t_8__749_,t_8__748_,t_8__747_,t_8__746_,t_8__745_,t_8__744_,t_8__743_,
  t_8__742_,t_8__741_,t_8__740_,t_8__739_,t_8__738_,t_8__737_,t_8__736_,t_8__735_,
  t_8__734_,t_8__733_,t_8__732_,t_8__731_,t_8__730_,t_8__729_,t_8__728_,t_8__727_,
  t_8__726_,t_8__725_,t_8__724_,t_8__723_,t_8__722_,t_8__721_,t_8__720_,t_8__719_,
  t_8__718_,t_8__717_,t_8__716_,t_8__715_,t_8__714_,t_8__713_,t_8__712_,t_8__711_,
  t_8__710_,t_8__709_,t_8__708_,t_8__707_,t_8__706_,t_8__705_,t_8__704_,t_8__703_,
  t_8__702_,t_8__701_,t_8__700_,t_8__699_,t_8__698_,t_8__697_,t_8__696_,t_8__695_,
  t_8__694_,t_8__693_,t_8__692_,t_8__691_,t_8__690_,t_8__689_,t_8__688_,t_8__687_,
  t_8__686_,t_8__685_,t_8__684_,t_8__683_,t_8__682_,t_8__681_,t_8__680_,t_8__679_,
  t_8__678_,t_8__677_,t_8__676_,t_8__675_,t_8__674_,t_8__673_,t_8__672_,t_8__671_,
  t_8__670_,t_8__669_,t_8__668_,t_8__667_,t_8__666_,t_8__665_,t_8__664_,t_8__663_,
  t_8__662_,t_8__661_,t_8__660_,t_8__659_,t_8__658_,t_8__657_,t_8__656_,t_8__655_,
  t_8__654_,t_8__653_,t_8__652_,t_8__651_,t_8__650_,t_8__649_,t_8__648_,t_8__647_,
  t_8__646_,t_8__645_,t_8__644_,t_8__643_,t_8__642_,t_8__641_,t_8__640_,t_8__639_,
  t_8__638_,t_8__637_,t_8__636_,t_8__635_,t_8__634_,t_8__633_,t_8__632_,t_8__631_,
  t_8__630_,t_8__629_,t_8__628_,t_8__627_,t_8__626_,t_8__625_,t_8__624_,t_8__623_,
  t_8__622_,t_8__621_,t_8__620_,t_8__619_,t_8__618_,t_8__617_,t_8__616_,t_8__615_,
  t_8__614_,t_8__613_,t_8__612_,t_8__611_,t_8__610_,t_8__609_,t_8__608_,t_8__607_,
  t_8__606_,t_8__605_,t_8__604_,t_8__603_,t_8__602_,t_8__601_,t_8__600_,t_8__599_,
  t_8__598_,t_8__597_,t_8__596_,t_8__595_,t_8__594_,t_8__593_,t_8__592_,t_8__591_,
  t_8__590_,t_8__589_,t_8__588_,t_8__587_,t_8__586_,t_8__585_,t_8__584_,t_8__583_,
  t_8__582_,t_8__581_,t_8__580_,t_8__579_,t_8__578_,t_8__577_,t_8__576_,t_8__575_,
  t_8__574_,t_8__573_,t_8__572_,t_8__571_,t_8__570_,t_8__569_,t_8__568_,t_8__567_,
  t_8__566_,t_8__565_,t_8__564_,t_8__563_,t_8__562_,t_8__561_,t_8__560_,t_8__559_,
  t_8__558_,t_8__557_,t_8__556_,t_8__555_,t_8__554_,t_8__553_,t_8__552_,t_8__551_,
  t_8__550_,t_8__549_,t_8__548_,t_8__547_,t_8__546_,t_8__545_,t_8__544_,t_8__543_,
  t_8__542_,t_8__541_,t_8__540_,t_8__539_,t_8__538_,t_8__537_,t_8__536_,t_8__535_,
  t_8__534_,t_8__533_,t_8__532_,t_8__531_,t_8__530_,t_8__529_,t_8__528_,t_8__527_,
  t_8__526_,t_8__525_,t_8__524_,t_8__523_,t_8__522_,t_8__521_,t_8__520_,t_8__519_,
  t_8__518_,t_8__517_,t_8__516_,t_8__515_,t_8__514_,t_8__513_,t_8__512_,t_8__511_,
  t_8__510_,t_8__509_,t_8__508_,t_8__507_,t_8__506_,t_8__505_,t_8__504_,t_8__503_,
  t_8__502_,t_8__501_,t_8__500_,t_8__499_,t_8__498_,t_8__497_,t_8__496_,t_8__495_,
  t_8__494_,t_8__493_,t_8__492_,t_8__491_,t_8__490_,t_8__489_,t_8__488_,t_8__487_,
  t_8__486_,t_8__485_,t_8__484_,t_8__483_,t_8__482_,t_8__481_,t_8__480_,t_8__479_,
  t_8__478_,t_8__477_,t_8__476_,t_8__475_,t_8__474_,t_8__473_,t_8__472_,t_8__471_,
  t_8__470_,t_8__469_,t_8__468_,t_8__467_,t_8__466_,t_8__465_,t_8__464_,t_8__463_,
  t_8__462_,t_8__461_,t_8__460_,t_8__459_,t_8__458_,t_8__457_,t_8__456_,t_8__455_,
  t_8__454_,t_8__453_,t_8__452_,t_8__451_,t_8__450_,t_8__449_,t_8__448_,t_8__447_,
  t_8__446_,t_8__445_,t_8__444_,t_8__443_,t_8__442_,t_8__441_,t_8__440_,t_8__439_,
  t_8__438_,t_8__437_,t_8__436_,t_8__435_,t_8__434_,t_8__433_,t_8__432_,t_8__431_,
  t_8__430_,t_8__429_,t_8__428_,t_8__427_,t_8__426_,t_8__425_,t_8__424_,t_8__423_,
  t_8__422_,t_8__421_,t_8__420_,t_8__419_,t_8__418_,t_8__417_,t_8__416_,t_8__415_,
  t_8__414_,t_8__413_,t_8__412_,t_8__411_,t_8__410_,t_8__409_,t_8__408_,t_8__407_,
  t_8__406_,t_8__405_,t_8__404_,t_8__403_,t_8__402_,t_8__401_,t_8__400_,t_8__399_,
  t_8__398_,t_8__397_,t_8__396_,t_8__395_,t_8__394_,t_8__393_,t_8__392_,t_8__391_,
  t_8__390_,t_8__389_,t_8__388_,t_8__387_,t_8__386_,t_8__385_,t_8__384_,t_8__383_,
  t_8__382_,t_8__381_,t_8__380_,t_8__379_,t_8__378_,t_8__377_,t_8__376_,t_8__375_,
  t_8__374_,t_8__373_,t_8__372_,t_8__371_,t_8__370_,t_8__369_,t_8__368_,t_8__367_,
  t_8__366_,t_8__365_,t_8__364_,t_8__363_,t_8__362_,t_8__361_,t_8__360_,t_8__359_,
  t_8__358_,t_8__357_,t_8__356_,t_8__355_,t_8__354_,t_8__353_,t_8__352_,t_8__351_,
  t_8__350_,t_8__349_,t_8__348_,t_8__347_,t_8__346_,t_8__345_,t_8__344_,t_8__343_,
  t_8__342_,t_8__341_,t_8__340_,t_8__339_,t_8__338_,t_8__337_,t_8__336_,t_8__335_,
  t_8__334_,t_8__333_,t_8__332_,t_8__331_,t_8__330_,t_8__329_,t_8__328_,t_8__327_,
  t_8__326_,t_8__325_,t_8__324_,t_8__323_,t_8__322_,t_8__321_,t_8__320_,t_8__319_,
  t_8__318_,t_8__317_,t_8__316_,t_8__315_,t_8__314_,t_8__313_,t_8__312_,t_8__311_,
  t_8__310_,t_8__309_,t_8__308_,t_8__307_,t_8__306_,t_8__305_,t_8__304_,t_8__303_,
  t_8__302_,t_8__301_,t_8__300_,t_8__299_,t_8__298_,t_8__297_,t_8__296_,t_8__295_,
  t_8__294_,t_8__293_,t_8__292_,t_8__291_,t_8__290_,t_8__289_,t_8__288_,t_8__287_,
  t_8__286_,t_8__285_,t_8__284_,t_8__283_,t_8__282_,t_8__281_,t_8__280_,t_8__279_,
  t_8__278_,t_8__277_,t_8__276_,t_8__275_,t_8__274_,t_8__273_,t_8__272_,t_8__271_,
  t_8__270_,t_8__269_,t_8__268_,t_8__267_,t_8__266_,t_8__265_,t_8__264_,t_8__263_,
  t_8__262_,t_8__261_,t_8__260_,t_8__259_,t_8__258_,t_8__257_,t_8__256_,t_8__255_,
  t_8__254_,t_8__253_,t_8__252_,t_8__251_,t_8__250_,t_8__249_,t_8__248_,t_8__247_,
  t_8__246_,t_8__245_,t_8__244_,t_8__243_,t_8__242_,t_8__241_,t_8__240_,t_8__239_,
  t_8__238_,t_8__237_,t_8__236_,t_8__235_,t_8__234_,t_8__233_,t_8__232_,t_8__231_,
  t_8__230_,t_8__229_,t_8__228_,t_8__227_,t_8__226_,t_8__225_,t_8__224_,t_8__223_,
  t_8__222_,t_8__221_,t_8__220_,t_8__219_,t_8__218_,t_8__217_,t_8__216_,t_8__215_,
  t_8__214_,t_8__213_,t_8__212_,t_8__211_,t_8__210_,t_8__209_,t_8__208_,t_8__207_,
  t_8__206_,t_8__205_,t_8__204_,t_8__203_,t_8__202_,t_8__201_,t_8__200_,t_8__199_,
  t_8__198_,t_8__197_,t_8__196_,t_8__195_,t_8__194_,t_8__193_,t_8__192_,t_8__191_,
  t_8__190_,t_8__189_,t_8__188_,t_8__187_,t_8__186_,t_8__185_,t_8__184_,t_8__183_,
  t_8__182_,t_8__181_,t_8__180_,t_8__179_,t_8__178_,t_8__177_,t_8__176_,t_8__175_,
  t_8__174_,t_8__173_,t_8__172_,t_8__171_,t_8__170_,t_8__169_,t_8__168_,t_8__167_,
  t_8__166_,t_8__165_,t_8__164_,t_8__163_,t_8__162_,t_8__161_,t_8__160_,t_8__159_,
  t_8__158_,t_8__157_,t_8__156_,t_8__155_,t_8__154_,t_8__153_,t_8__152_,t_8__151_,
  t_8__150_,t_8__149_,t_8__148_,t_8__147_,t_8__146_,t_8__145_,t_8__144_,t_8__143_,
  t_8__142_,t_8__141_,t_8__140_,t_8__139_,t_8__138_,t_8__137_,t_8__136_,t_8__135_,
  t_8__134_,t_8__133_,t_8__132_,t_8__131_,t_8__130_,t_8__129_,t_8__128_,t_8__127_,
  t_8__126_,t_8__125_,t_8__124_,t_8__123_,t_8__122_,t_8__121_,t_8__120_,t_8__119_,
  t_8__118_,t_8__117_,t_8__116_,t_8__115_,t_8__114_,t_8__113_,t_8__112_,t_8__111_,
  t_8__110_,t_8__109_,t_8__108_,t_8__107_,t_8__106_,t_8__105_,t_8__104_,t_8__103_,
  t_8__102_,t_8__101_,t_8__100_,t_8__99_,t_8__98_,t_8__97_,t_8__96_,t_8__95_,t_8__94_,
  t_8__93_,t_8__92_,t_8__91_,t_8__90_,t_8__89_,t_8__88_,t_8__87_,t_8__86_,t_8__85_,
  t_8__84_,t_8__83_,t_8__82_,t_8__81_,t_8__80_,t_8__79_,t_8__78_,t_8__77_,t_8__76_,
  t_8__75_,t_8__74_,t_8__73_,t_8__72_,t_8__71_,t_8__70_,t_8__69_,t_8__68_,t_8__67_,
  t_8__66_,t_8__65_,t_8__64_,t_8__63_,t_8__62_,t_8__61_,t_8__60_,t_8__59_,t_8__58_,
  t_8__57_,t_8__56_,t_8__55_,t_8__54_,t_8__53_,t_8__52_,t_8__51_,t_8__50_,
  t_8__49_,t_8__48_,t_8__47_,t_8__46_,t_8__45_,t_8__44_,t_8__43_,t_8__42_,t_8__41_,
  t_8__40_,t_8__39_,t_8__38_,t_8__37_,t_8__36_,t_8__35_,t_8__34_,t_8__33_,t_8__32_,
  t_8__31_,t_8__30_,t_8__29_,t_8__28_,t_8__27_,t_8__26_,t_8__25_,t_8__24_,t_8__23_,
  t_8__22_,t_8__21_,t_8__20_,t_8__19_,t_8__18_,t_8__17_,t_8__16_,t_8__15_,t_8__14_,
  t_8__13_,t_8__12_,t_8__11_,t_8__10_,t_8__9_,t_8__8_,t_8__7_,t_8__6_,t_8__5_,t_8__4_,
  t_8__3_,t_8__2_,t_8__1_,t_8__0_,t_9__1023_,t_9__1022_,t_9__1021_,t_9__1020_,
  t_9__1019_,t_9__1018_,t_9__1017_,t_9__1016_,t_9__1015_,t_9__1014_,t_9__1013_,
  t_9__1012_,t_9__1011_,t_9__1010_,t_9__1009_,t_9__1008_,t_9__1007_,t_9__1006_,
  t_9__1005_,t_9__1004_,t_9__1003_,t_9__1002_,t_9__1001_,t_9__1000_,t_9__999_,t_9__998_,
  t_9__997_,t_9__996_,t_9__995_,t_9__994_,t_9__993_,t_9__992_,t_9__991_,t_9__990_,
  t_9__989_,t_9__988_,t_9__987_,t_9__986_,t_9__985_,t_9__984_,t_9__983_,t_9__982_,
  t_9__981_,t_9__980_,t_9__979_,t_9__978_,t_9__977_,t_9__976_,t_9__975_,t_9__974_,
  t_9__973_,t_9__972_,t_9__971_,t_9__970_,t_9__969_,t_9__968_,t_9__967_,t_9__966_,
  t_9__965_,t_9__964_,t_9__963_,t_9__962_,t_9__961_,t_9__960_,t_9__959_,t_9__958_,
  t_9__957_,t_9__956_,t_9__955_,t_9__954_,t_9__953_,t_9__952_,t_9__951_,t_9__950_,
  t_9__949_,t_9__948_,t_9__947_,t_9__946_,t_9__945_,t_9__944_,t_9__943_,t_9__942_,
  t_9__941_,t_9__940_,t_9__939_,t_9__938_,t_9__937_,t_9__936_,t_9__935_,t_9__934_,
  t_9__933_,t_9__932_,t_9__931_,t_9__930_,t_9__929_,t_9__928_,t_9__927_,t_9__926_,
  t_9__925_,t_9__924_,t_9__923_,t_9__922_,t_9__921_,t_9__920_,t_9__919_,t_9__918_,
  t_9__917_,t_9__916_,t_9__915_,t_9__914_,t_9__913_,t_9__912_,t_9__911_,t_9__910_,
  t_9__909_,t_9__908_,t_9__907_,t_9__906_,t_9__905_,t_9__904_,t_9__903_,t_9__902_,
  t_9__901_,t_9__900_,t_9__899_,t_9__898_,t_9__897_,t_9__896_,t_9__895_,t_9__894_,
  t_9__893_,t_9__892_,t_9__891_,t_9__890_,t_9__889_,t_9__888_,t_9__887_,t_9__886_,
  t_9__885_,t_9__884_,t_9__883_,t_9__882_,t_9__881_,t_9__880_,t_9__879_,t_9__878_,
  t_9__877_,t_9__876_,t_9__875_,t_9__874_,t_9__873_,t_9__872_,t_9__871_,t_9__870_,
  t_9__869_,t_9__868_,t_9__867_,t_9__866_,t_9__865_,t_9__864_,t_9__863_,t_9__862_,
  t_9__861_,t_9__860_,t_9__859_,t_9__858_,t_9__857_,t_9__856_,t_9__855_,t_9__854_,
  t_9__853_,t_9__852_,t_9__851_,t_9__850_,t_9__849_,t_9__848_,t_9__847_,t_9__846_,
  t_9__845_,t_9__844_,t_9__843_,t_9__842_,t_9__841_,t_9__840_,t_9__839_,t_9__838_,
  t_9__837_,t_9__836_,t_9__835_,t_9__834_,t_9__833_,t_9__832_,t_9__831_,t_9__830_,
  t_9__829_,t_9__828_,t_9__827_,t_9__826_,t_9__825_,t_9__824_,t_9__823_,t_9__822_,
  t_9__821_,t_9__820_,t_9__819_,t_9__818_,t_9__817_,t_9__816_,t_9__815_,t_9__814_,
  t_9__813_,t_9__812_,t_9__811_,t_9__810_,t_9__809_,t_9__808_,t_9__807_,t_9__806_,
  t_9__805_,t_9__804_,t_9__803_,t_9__802_,t_9__801_,t_9__800_,t_9__799_,t_9__798_,
  t_9__797_,t_9__796_,t_9__795_,t_9__794_,t_9__793_,t_9__792_,t_9__791_,t_9__790_,
  t_9__789_,t_9__788_,t_9__787_,t_9__786_,t_9__785_,t_9__784_,t_9__783_,t_9__782_,
  t_9__781_,t_9__780_,t_9__779_,t_9__778_,t_9__777_,t_9__776_,t_9__775_,t_9__774_,
  t_9__773_,t_9__772_,t_9__771_,t_9__770_,t_9__769_,t_9__768_,t_9__767_,t_9__766_,
  t_9__765_,t_9__764_,t_9__763_,t_9__762_,t_9__761_,t_9__760_,t_9__759_,t_9__758_,
  t_9__757_,t_9__756_,t_9__755_,t_9__754_,t_9__753_,t_9__752_,t_9__751_,t_9__750_,
  t_9__749_,t_9__748_,t_9__747_,t_9__746_,t_9__745_,t_9__744_,t_9__743_,t_9__742_,
  t_9__741_,t_9__740_,t_9__739_,t_9__738_,t_9__737_,t_9__736_,t_9__735_,t_9__734_,
  t_9__733_,t_9__732_,t_9__731_,t_9__730_,t_9__729_,t_9__728_,t_9__727_,t_9__726_,
  t_9__725_,t_9__724_,t_9__723_,t_9__722_,t_9__721_,t_9__720_,t_9__719_,t_9__718_,
  t_9__717_,t_9__716_,t_9__715_,t_9__714_,t_9__713_,t_9__712_,t_9__711_,t_9__710_,
  t_9__709_,t_9__708_,t_9__707_,t_9__706_,t_9__705_,t_9__704_,t_9__703_,t_9__702_,
  t_9__701_,t_9__700_,t_9__699_,t_9__698_,t_9__697_,t_9__696_,t_9__695_,t_9__694_,
  t_9__693_,t_9__692_,t_9__691_,t_9__690_,t_9__689_,t_9__688_,t_9__687_,t_9__686_,
  t_9__685_,t_9__684_,t_9__683_,t_9__682_,t_9__681_,t_9__680_,t_9__679_,t_9__678_,
  t_9__677_,t_9__676_,t_9__675_,t_9__674_,t_9__673_,t_9__672_,t_9__671_,t_9__670_,
  t_9__669_,t_9__668_,t_9__667_,t_9__666_,t_9__665_,t_9__664_,t_9__663_,t_9__662_,
  t_9__661_,t_9__660_,t_9__659_,t_9__658_,t_9__657_,t_9__656_,t_9__655_,t_9__654_,
  t_9__653_,t_9__652_,t_9__651_,t_9__650_,t_9__649_,t_9__648_,t_9__647_,t_9__646_,
  t_9__645_,t_9__644_,t_9__643_,t_9__642_,t_9__641_,t_9__640_,t_9__639_,t_9__638_,
  t_9__637_,t_9__636_,t_9__635_,t_9__634_,t_9__633_,t_9__632_,t_9__631_,t_9__630_,
  t_9__629_,t_9__628_,t_9__627_,t_9__626_,t_9__625_,t_9__624_,t_9__623_,t_9__622_,
  t_9__621_,t_9__620_,t_9__619_,t_9__618_,t_9__617_,t_9__616_,t_9__615_,t_9__614_,
  t_9__613_,t_9__612_,t_9__611_,t_9__610_,t_9__609_,t_9__608_,t_9__607_,t_9__606_,
  t_9__605_,t_9__604_,t_9__603_,t_9__602_,t_9__601_,t_9__600_,t_9__599_,t_9__598_,
  t_9__597_,t_9__596_,t_9__595_,t_9__594_,t_9__593_,t_9__592_,t_9__591_,t_9__590_,
  t_9__589_,t_9__588_,t_9__587_,t_9__586_,t_9__585_,t_9__584_,t_9__583_,t_9__582_,
  t_9__581_,t_9__580_,t_9__579_,t_9__578_,t_9__577_,t_9__576_,t_9__575_,t_9__574_,
  t_9__573_,t_9__572_,t_9__571_,t_9__570_,t_9__569_,t_9__568_,t_9__567_,t_9__566_,
  t_9__565_,t_9__564_,t_9__563_,t_9__562_,t_9__561_,t_9__560_,t_9__559_,t_9__558_,
  t_9__557_,t_9__556_,t_9__555_,t_9__554_,t_9__553_,t_9__552_,t_9__551_,t_9__550_,
  t_9__549_,t_9__548_,t_9__547_,t_9__546_,t_9__545_,t_9__544_,t_9__543_,t_9__542_,
  t_9__541_,t_9__540_,t_9__539_,t_9__538_,t_9__537_,t_9__536_,t_9__535_,t_9__534_,
  t_9__533_,t_9__532_,t_9__531_,t_9__530_,t_9__529_,t_9__528_,t_9__527_,t_9__526_,
  t_9__525_,t_9__524_,t_9__523_,t_9__522_,t_9__521_,t_9__520_,t_9__519_,t_9__518_,
  t_9__517_,t_9__516_,t_9__515_,t_9__514_,t_9__513_,t_9__512_,t_9__511_,t_9__510_,
  t_9__509_,t_9__508_,t_9__507_,t_9__506_,t_9__505_,t_9__504_,t_9__503_,t_9__502_,
  t_9__501_,t_9__500_,t_9__499_,t_9__498_,t_9__497_,t_9__496_,t_9__495_,t_9__494_,
  t_9__493_,t_9__492_,t_9__491_,t_9__490_,t_9__489_,t_9__488_,t_9__487_,t_9__486_,
  t_9__485_,t_9__484_,t_9__483_,t_9__482_,t_9__481_,t_9__480_,t_9__479_,t_9__478_,
  t_9__477_,t_9__476_,t_9__475_,t_9__474_,t_9__473_,t_9__472_,t_9__471_,t_9__470_,
  t_9__469_,t_9__468_,t_9__467_,t_9__466_,t_9__465_,t_9__464_,t_9__463_,t_9__462_,
  t_9__461_,t_9__460_,t_9__459_,t_9__458_,t_9__457_,t_9__456_,t_9__455_,t_9__454_,
  t_9__453_,t_9__452_,t_9__451_,t_9__450_,t_9__449_,t_9__448_,t_9__447_,t_9__446_,
  t_9__445_,t_9__444_,t_9__443_,t_9__442_,t_9__441_,t_9__440_,t_9__439_,t_9__438_,
  t_9__437_,t_9__436_,t_9__435_,t_9__434_,t_9__433_,t_9__432_,t_9__431_,t_9__430_,
  t_9__429_,t_9__428_,t_9__427_,t_9__426_,t_9__425_,t_9__424_,t_9__423_,t_9__422_,
  t_9__421_,t_9__420_,t_9__419_,t_9__418_,t_9__417_,t_9__416_,t_9__415_,t_9__414_,
  t_9__413_,t_9__412_,t_9__411_,t_9__410_,t_9__409_,t_9__408_,t_9__407_,t_9__406_,
  t_9__405_,t_9__404_,t_9__403_,t_9__402_,t_9__401_,t_9__400_,t_9__399_,t_9__398_,
  t_9__397_,t_9__396_,t_9__395_,t_9__394_,t_9__393_,t_9__392_,t_9__391_,t_9__390_,
  t_9__389_,t_9__388_,t_9__387_,t_9__386_,t_9__385_,t_9__384_,t_9__383_,t_9__382_,
  t_9__381_,t_9__380_,t_9__379_,t_9__378_,t_9__377_,t_9__376_,t_9__375_,t_9__374_,
  t_9__373_,t_9__372_,t_9__371_,t_9__370_,t_9__369_,t_9__368_,t_9__367_,t_9__366_,
  t_9__365_,t_9__364_,t_9__363_,t_9__362_,t_9__361_,t_9__360_,t_9__359_,t_9__358_,
  t_9__357_,t_9__356_,t_9__355_,t_9__354_,t_9__353_,t_9__352_,t_9__351_,t_9__350_,
  t_9__349_,t_9__348_,t_9__347_,t_9__346_,t_9__345_,t_9__344_,t_9__343_,t_9__342_,
  t_9__341_,t_9__340_,t_9__339_,t_9__338_,t_9__337_,t_9__336_,t_9__335_,t_9__334_,
  t_9__333_,t_9__332_,t_9__331_,t_9__330_,t_9__329_,t_9__328_,t_9__327_,t_9__326_,
  t_9__325_,t_9__324_,t_9__323_,t_9__322_,t_9__321_,t_9__320_,t_9__319_,t_9__318_,
  t_9__317_,t_9__316_,t_9__315_,t_9__314_,t_9__313_,t_9__312_,t_9__311_,t_9__310_,
  t_9__309_,t_9__308_,t_9__307_,t_9__306_,t_9__305_,t_9__304_,t_9__303_,t_9__302_,
  t_9__301_,t_9__300_,t_9__299_,t_9__298_,t_9__297_,t_9__296_,t_9__295_,t_9__294_,
  t_9__293_,t_9__292_,t_9__291_,t_9__290_,t_9__289_,t_9__288_,t_9__287_,t_9__286_,
  t_9__285_,t_9__284_,t_9__283_,t_9__282_,t_9__281_,t_9__280_,t_9__279_,t_9__278_,
  t_9__277_,t_9__276_,t_9__275_,t_9__274_,t_9__273_,t_9__272_,t_9__271_,t_9__270_,
  t_9__269_,t_9__268_,t_9__267_,t_9__266_,t_9__265_,t_9__264_,t_9__263_,t_9__262_,
  t_9__261_,t_9__260_,t_9__259_,t_9__258_,t_9__257_,t_9__256_,t_9__255_,t_9__254_,
  t_9__253_,t_9__252_,t_9__251_,t_9__250_,t_9__249_,t_9__248_,t_9__247_,t_9__246_,
  t_9__245_,t_9__244_,t_9__243_,t_9__242_,t_9__241_,t_9__240_,t_9__239_,t_9__238_,
  t_9__237_,t_9__236_,t_9__235_,t_9__234_,t_9__233_,t_9__232_,t_9__231_,t_9__230_,
  t_9__229_,t_9__228_,t_9__227_,t_9__226_,t_9__225_,t_9__224_,t_9__223_,t_9__222_,
  t_9__221_,t_9__220_,t_9__219_,t_9__218_,t_9__217_,t_9__216_,t_9__215_,t_9__214_,
  t_9__213_,t_9__212_,t_9__211_,t_9__210_,t_9__209_,t_9__208_,t_9__207_,t_9__206_,
  t_9__205_,t_9__204_,t_9__203_,t_9__202_,t_9__201_,t_9__200_,t_9__199_,t_9__198_,
  t_9__197_,t_9__196_,t_9__195_,t_9__194_,t_9__193_,t_9__192_,t_9__191_,t_9__190_,
  t_9__189_,t_9__188_,t_9__187_,t_9__186_,t_9__185_,t_9__184_,t_9__183_,t_9__182_,
  t_9__181_,t_9__180_,t_9__179_,t_9__178_,t_9__177_,t_9__176_,t_9__175_,t_9__174_,
  t_9__173_,t_9__172_,t_9__171_,t_9__170_,t_9__169_,t_9__168_,t_9__167_,t_9__166_,
  t_9__165_,t_9__164_,t_9__163_,t_9__162_,t_9__161_,t_9__160_,t_9__159_,t_9__158_,
  t_9__157_,t_9__156_,t_9__155_,t_9__154_,t_9__153_,t_9__152_,t_9__151_,t_9__150_,
  t_9__149_,t_9__148_,t_9__147_,t_9__146_,t_9__145_,t_9__144_,t_9__143_,t_9__142_,
  t_9__141_,t_9__140_,t_9__139_,t_9__138_,t_9__137_,t_9__136_,t_9__135_,t_9__134_,
  t_9__133_,t_9__132_,t_9__131_,t_9__130_,t_9__129_,t_9__128_,t_9__127_,t_9__126_,
  t_9__125_,t_9__124_,t_9__123_,t_9__122_,t_9__121_,t_9__120_,t_9__119_,t_9__118_,
  t_9__117_,t_9__116_,t_9__115_,t_9__114_,t_9__113_,t_9__112_,t_9__111_,t_9__110_,
  t_9__109_,t_9__108_,t_9__107_,t_9__106_,t_9__105_,t_9__104_,t_9__103_,t_9__102_,
  t_9__101_,t_9__100_,t_9__99_,t_9__98_,t_9__97_,t_9__96_,t_9__95_,t_9__94_,t_9__93_,
  t_9__92_,t_9__91_,t_9__90_,t_9__89_,t_9__88_,t_9__87_,t_9__86_,t_9__85_,t_9__84_,
  t_9__83_,t_9__82_,t_9__81_,t_9__80_,t_9__79_,t_9__78_,t_9__77_,t_9__76_,
  t_9__75_,t_9__74_,t_9__73_,t_9__72_,t_9__71_,t_9__70_,t_9__69_,t_9__68_,t_9__67_,
  t_9__66_,t_9__65_,t_9__64_,t_9__63_,t_9__62_,t_9__61_,t_9__60_,t_9__59_,t_9__58_,
  t_9__57_,t_9__56_,t_9__55_,t_9__54_,t_9__53_,t_9__52_,t_9__51_,t_9__50_,t_9__49_,
  t_9__48_,t_9__47_,t_9__46_,t_9__45_,t_9__44_,t_9__43_,t_9__42_,t_9__41_,t_9__40_,
  t_9__39_,t_9__38_,t_9__37_,t_9__36_,t_9__35_,t_9__34_,t_9__33_,t_9__32_,t_9__31_,
  t_9__30_,t_9__29_,t_9__28_,t_9__27_,t_9__26_,t_9__25_,t_9__24_,t_9__23_,t_9__22_,
  t_9__21_,t_9__20_,t_9__19_,t_9__18_,t_9__17_,t_9__16_,t_9__15_,t_9__14_,t_9__13_,
  t_9__12_,t_9__11_,t_9__10_,t_9__9_,t_9__8_,t_9__7_,t_9__6_,t_9__5_,t_9__4_,
  t_9__3_,t_9__2_,t_9__1_,t_9__0_;
  assign t_1__1023_ = i[0] | 1'b0;
  assign t_1__1022_ = i[1] | i[0];
  assign t_1__1021_ = i[2] | i[1];
  assign t_1__1020_ = i[3] | i[2];
  assign t_1__1019_ = i[4] | i[3];
  assign t_1__1018_ = i[5] | i[4];
  assign t_1__1017_ = i[6] | i[5];
  assign t_1__1016_ = i[7] | i[6];
  assign t_1__1015_ = i[8] | i[7];
  assign t_1__1014_ = i[9] | i[8];
  assign t_1__1013_ = i[10] | i[9];
  assign t_1__1012_ = i[11] | i[10];
  assign t_1__1011_ = i[12] | i[11];
  assign t_1__1010_ = i[13] | i[12];
  assign t_1__1009_ = i[14] | i[13];
  assign t_1__1008_ = i[15] | i[14];
  assign t_1__1007_ = i[16] | i[15];
  assign t_1__1006_ = i[17] | i[16];
  assign t_1__1005_ = i[18] | i[17];
  assign t_1__1004_ = i[19] | i[18];
  assign t_1__1003_ = i[20] | i[19];
  assign t_1__1002_ = i[21] | i[20];
  assign t_1__1001_ = i[22] | i[21];
  assign t_1__1000_ = i[23] | i[22];
  assign t_1__999_ = i[24] | i[23];
  assign t_1__998_ = i[25] | i[24];
  assign t_1__997_ = i[26] | i[25];
  assign t_1__996_ = i[27] | i[26];
  assign t_1__995_ = i[28] | i[27];
  assign t_1__994_ = i[29] | i[28];
  assign t_1__993_ = i[30] | i[29];
  assign t_1__992_ = i[31] | i[30];
  assign t_1__991_ = i[32] | i[31];
  assign t_1__990_ = i[33] | i[32];
  assign t_1__989_ = i[34] | i[33];
  assign t_1__988_ = i[35] | i[34];
  assign t_1__987_ = i[36] | i[35];
  assign t_1__986_ = i[37] | i[36];
  assign t_1__985_ = i[38] | i[37];
  assign t_1__984_ = i[39] | i[38];
  assign t_1__983_ = i[40] | i[39];
  assign t_1__982_ = i[41] | i[40];
  assign t_1__981_ = i[42] | i[41];
  assign t_1__980_ = i[43] | i[42];
  assign t_1__979_ = i[44] | i[43];
  assign t_1__978_ = i[45] | i[44];
  assign t_1__977_ = i[46] | i[45];
  assign t_1__976_ = i[47] | i[46];
  assign t_1__975_ = i[48] | i[47];
  assign t_1__974_ = i[49] | i[48];
  assign t_1__973_ = i[50] | i[49];
  assign t_1__972_ = i[51] | i[50];
  assign t_1__971_ = i[52] | i[51];
  assign t_1__970_ = i[53] | i[52];
  assign t_1__969_ = i[54] | i[53];
  assign t_1__968_ = i[55] | i[54];
  assign t_1__967_ = i[56] | i[55];
  assign t_1__966_ = i[57] | i[56];
  assign t_1__965_ = i[58] | i[57];
  assign t_1__964_ = i[59] | i[58];
  assign t_1__963_ = i[60] | i[59];
  assign t_1__962_ = i[61] | i[60];
  assign t_1__961_ = i[62] | i[61];
  assign t_1__960_ = i[63] | i[62];
  assign t_1__959_ = i[64] | i[63];
  assign t_1__958_ = i[65] | i[64];
  assign t_1__957_ = i[66] | i[65];
  assign t_1__956_ = i[67] | i[66];
  assign t_1__955_ = i[68] | i[67];
  assign t_1__954_ = i[69] | i[68];
  assign t_1__953_ = i[70] | i[69];
  assign t_1__952_ = i[71] | i[70];
  assign t_1__951_ = i[72] | i[71];
  assign t_1__950_ = i[73] | i[72];
  assign t_1__949_ = i[74] | i[73];
  assign t_1__948_ = i[75] | i[74];
  assign t_1__947_ = i[76] | i[75];
  assign t_1__946_ = i[77] | i[76];
  assign t_1__945_ = i[78] | i[77];
  assign t_1__944_ = i[79] | i[78];
  assign t_1__943_ = i[80] | i[79];
  assign t_1__942_ = i[81] | i[80];
  assign t_1__941_ = i[82] | i[81];
  assign t_1__940_ = i[83] | i[82];
  assign t_1__939_ = i[84] | i[83];
  assign t_1__938_ = i[85] | i[84];
  assign t_1__937_ = i[86] | i[85];
  assign t_1__936_ = i[87] | i[86];
  assign t_1__935_ = i[88] | i[87];
  assign t_1__934_ = i[89] | i[88];
  assign t_1__933_ = i[90] | i[89];
  assign t_1__932_ = i[91] | i[90];
  assign t_1__931_ = i[92] | i[91];
  assign t_1__930_ = i[93] | i[92];
  assign t_1__929_ = i[94] | i[93];
  assign t_1__928_ = i[95] | i[94];
  assign t_1__927_ = i[96] | i[95];
  assign t_1__926_ = i[97] | i[96];
  assign t_1__925_ = i[98] | i[97];
  assign t_1__924_ = i[99] | i[98];
  assign t_1__923_ = i[100] | i[99];
  assign t_1__922_ = i[101] | i[100];
  assign t_1__921_ = i[102] | i[101];
  assign t_1__920_ = i[103] | i[102];
  assign t_1__919_ = i[104] | i[103];
  assign t_1__918_ = i[105] | i[104];
  assign t_1__917_ = i[106] | i[105];
  assign t_1__916_ = i[107] | i[106];
  assign t_1__915_ = i[108] | i[107];
  assign t_1__914_ = i[109] | i[108];
  assign t_1__913_ = i[110] | i[109];
  assign t_1__912_ = i[111] | i[110];
  assign t_1__911_ = i[112] | i[111];
  assign t_1__910_ = i[113] | i[112];
  assign t_1__909_ = i[114] | i[113];
  assign t_1__908_ = i[115] | i[114];
  assign t_1__907_ = i[116] | i[115];
  assign t_1__906_ = i[117] | i[116];
  assign t_1__905_ = i[118] | i[117];
  assign t_1__904_ = i[119] | i[118];
  assign t_1__903_ = i[120] | i[119];
  assign t_1__902_ = i[121] | i[120];
  assign t_1__901_ = i[122] | i[121];
  assign t_1__900_ = i[123] | i[122];
  assign t_1__899_ = i[124] | i[123];
  assign t_1__898_ = i[125] | i[124];
  assign t_1__897_ = i[126] | i[125];
  assign t_1__896_ = i[127] | i[126];
  assign t_1__895_ = i[128] | i[127];
  assign t_1__894_ = i[129] | i[128];
  assign t_1__893_ = i[130] | i[129];
  assign t_1__892_ = i[131] | i[130];
  assign t_1__891_ = i[132] | i[131];
  assign t_1__890_ = i[133] | i[132];
  assign t_1__889_ = i[134] | i[133];
  assign t_1__888_ = i[135] | i[134];
  assign t_1__887_ = i[136] | i[135];
  assign t_1__886_ = i[137] | i[136];
  assign t_1__885_ = i[138] | i[137];
  assign t_1__884_ = i[139] | i[138];
  assign t_1__883_ = i[140] | i[139];
  assign t_1__882_ = i[141] | i[140];
  assign t_1__881_ = i[142] | i[141];
  assign t_1__880_ = i[143] | i[142];
  assign t_1__879_ = i[144] | i[143];
  assign t_1__878_ = i[145] | i[144];
  assign t_1__877_ = i[146] | i[145];
  assign t_1__876_ = i[147] | i[146];
  assign t_1__875_ = i[148] | i[147];
  assign t_1__874_ = i[149] | i[148];
  assign t_1__873_ = i[150] | i[149];
  assign t_1__872_ = i[151] | i[150];
  assign t_1__871_ = i[152] | i[151];
  assign t_1__870_ = i[153] | i[152];
  assign t_1__869_ = i[154] | i[153];
  assign t_1__868_ = i[155] | i[154];
  assign t_1__867_ = i[156] | i[155];
  assign t_1__866_ = i[157] | i[156];
  assign t_1__865_ = i[158] | i[157];
  assign t_1__864_ = i[159] | i[158];
  assign t_1__863_ = i[160] | i[159];
  assign t_1__862_ = i[161] | i[160];
  assign t_1__861_ = i[162] | i[161];
  assign t_1__860_ = i[163] | i[162];
  assign t_1__859_ = i[164] | i[163];
  assign t_1__858_ = i[165] | i[164];
  assign t_1__857_ = i[166] | i[165];
  assign t_1__856_ = i[167] | i[166];
  assign t_1__855_ = i[168] | i[167];
  assign t_1__854_ = i[169] | i[168];
  assign t_1__853_ = i[170] | i[169];
  assign t_1__852_ = i[171] | i[170];
  assign t_1__851_ = i[172] | i[171];
  assign t_1__850_ = i[173] | i[172];
  assign t_1__849_ = i[174] | i[173];
  assign t_1__848_ = i[175] | i[174];
  assign t_1__847_ = i[176] | i[175];
  assign t_1__846_ = i[177] | i[176];
  assign t_1__845_ = i[178] | i[177];
  assign t_1__844_ = i[179] | i[178];
  assign t_1__843_ = i[180] | i[179];
  assign t_1__842_ = i[181] | i[180];
  assign t_1__841_ = i[182] | i[181];
  assign t_1__840_ = i[183] | i[182];
  assign t_1__839_ = i[184] | i[183];
  assign t_1__838_ = i[185] | i[184];
  assign t_1__837_ = i[186] | i[185];
  assign t_1__836_ = i[187] | i[186];
  assign t_1__835_ = i[188] | i[187];
  assign t_1__834_ = i[189] | i[188];
  assign t_1__833_ = i[190] | i[189];
  assign t_1__832_ = i[191] | i[190];
  assign t_1__831_ = i[192] | i[191];
  assign t_1__830_ = i[193] | i[192];
  assign t_1__829_ = i[194] | i[193];
  assign t_1__828_ = i[195] | i[194];
  assign t_1__827_ = i[196] | i[195];
  assign t_1__826_ = i[197] | i[196];
  assign t_1__825_ = i[198] | i[197];
  assign t_1__824_ = i[199] | i[198];
  assign t_1__823_ = i[200] | i[199];
  assign t_1__822_ = i[201] | i[200];
  assign t_1__821_ = i[202] | i[201];
  assign t_1__820_ = i[203] | i[202];
  assign t_1__819_ = i[204] | i[203];
  assign t_1__818_ = i[205] | i[204];
  assign t_1__817_ = i[206] | i[205];
  assign t_1__816_ = i[207] | i[206];
  assign t_1__815_ = i[208] | i[207];
  assign t_1__814_ = i[209] | i[208];
  assign t_1__813_ = i[210] | i[209];
  assign t_1__812_ = i[211] | i[210];
  assign t_1__811_ = i[212] | i[211];
  assign t_1__810_ = i[213] | i[212];
  assign t_1__809_ = i[214] | i[213];
  assign t_1__808_ = i[215] | i[214];
  assign t_1__807_ = i[216] | i[215];
  assign t_1__806_ = i[217] | i[216];
  assign t_1__805_ = i[218] | i[217];
  assign t_1__804_ = i[219] | i[218];
  assign t_1__803_ = i[220] | i[219];
  assign t_1__802_ = i[221] | i[220];
  assign t_1__801_ = i[222] | i[221];
  assign t_1__800_ = i[223] | i[222];
  assign t_1__799_ = i[224] | i[223];
  assign t_1__798_ = i[225] | i[224];
  assign t_1__797_ = i[226] | i[225];
  assign t_1__796_ = i[227] | i[226];
  assign t_1__795_ = i[228] | i[227];
  assign t_1__794_ = i[229] | i[228];
  assign t_1__793_ = i[230] | i[229];
  assign t_1__792_ = i[231] | i[230];
  assign t_1__791_ = i[232] | i[231];
  assign t_1__790_ = i[233] | i[232];
  assign t_1__789_ = i[234] | i[233];
  assign t_1__788_ = i[235] | i[234];
  assign t_1__787_ = i[236] | i[235];
  assign t_1__786_ = i[237] | i[236];
  assign t_1__785_ = i[238] | i[237];
  assign t_1__784_ = i[239] | i[238];
  assign t_1__783_ = i[240] | i[239];
  assign t_1__782_ = i[241] | i[240];
  assign t_1__781_ = i[242] | i[241];
  assign t_1__780_ = i[243] | i[242];
  assign t_1__779_ = i[244] | i[243];
  assign t_1__778_ = i[245] | i[244];
  assign t_1__777_ = i[246] | i[245];
  assign t_1__776_ = i[247] | i[246];
  assign t_1__775_ = i[248] | i[247];
  assign t_1__774_ = i[249] | i[248];
  assign t_1__773_ = i[250] | i[249];
  assign t_1__772_ = i[251] | i[250];
  assign t_1__771_ = i[252] | i[251];
  assign t_1__770_ = i[253] | i[252];
  assign t_1__769_ = i[254] | i[253];
  assign t_1__768_ = i[255] | i[254];
  assign t_1__767_ = i[256] | i[255];
  assign t_1__766_ = i[257] | i[256];
  assign t_1__765_ = i[258] | i[257];
  assign t_1__764_ = i[259] | i[258];
  assign t_1__763_ = i[260] | i[259];
  assign t_1__762_ = i[261] | i[260];
  assign t_1__761_ = i[262] | i[261];
  assign t_1__760_ = i[263] | i[262];
  assign t_1__759_ = i[264] | i[263];
  assign t_1__758_ = i[265] | i[264];
  assign t_1__757_ = i[266] | i[265];
  assign t_1__756_ = i[267] | i[266];
  assign t_1__755_ = i[268] | i[267];
  assign t_1__754_ = i[269] | i[268];
  assign t_1__753_ = i[270] | i[269];
  assign t_1__752_ = i[271] | i[270];
  assign t_1__751_ = i[272] | i[271];
  assign t_1__750_ = i[273] | i[272];
  assign t_1__749_ = i[274] | i[273];
  assign t_1__748_ = i[275] | i[274];
  assign t_1__747_ = i[276] | i[275];
  assign t_1__746_ = i[277] | i[276];
  assign t_1__745_ = i[278] | i[277];
  assign t_1__744_ = i[279] | i[278];
  assign t_1__743_ = i[280] | i[279];
  assign t_1__742_ = i[281] | i[280];
  assign t_1__741_ = i[282] | i[281];
  assign t_1__740_ = i[283] | i[282];
  assign t_1__739_ = i[284] | i[283];
  assign t_1__738_ = i[285] | i[284];
  assign t_1__737_ = i[286] | i[285];
  assign t_1__736_ = i[287] | i[286];
  assign t_1__735_ = i[288] | i[287];
  assign t_1__734_ = i[289] | i[288];
  assign t_1__733_ = i[290] | i[289];
  assign t_1__732_ = i[291] | i[290];
  assign t_1__731_ = i[292] | i[291];
  assign t_1__730_ = i[293] | i[292];
  assign t_1__729_ = i[294] | i[293];
  assign t_1__728_ = i[295] | i[294];
  assign t_1__727_ = i[296] | i[295];
  assign t_1__726_ = i[297] | i[296];
  assign t_1__725_ = i[298] | i[297];
  assign t_1__724_ = i[299] | i[298];
  assign t_1__723_ = i[300] | i[299];
  assign t_1__722_ = i[301] | i[300];
  assign t_1__721_ = i[302] | i[301];
  assign t_1__720_ = i[303] | i[302];
  assign t_1__719_ = i[304] | i[303];
  assign t_1__718_ = i[305] | i[304];
  assign t_1__717_ = i[306] | i[305];
  assign t_1__716_ = i[307] | i[306];
  assign t_1__715_ = i[308] | i[307];
  assign t_1__714_ = i[309] | i[308];
  assign t_1__713_ = i[310] | i[309];
  assign t_1__712_ = i[311] | i[310];
  assign t_1__711_ = i[312] | i[311];
  assign t_1__710_ = i[313] | i[312];
  assign t_1__709_ = i[314] | i[313];
  assign t_1__708_ = i[315] | i[314];
  assign t_1__707_ = i[316] | i[315];
  assign t_1__706_ = i[317] | i[316];
  assign t_1__705_ = i[318] | i[317];
  assign t_1__704_ = i[319] | i[318];
  assign t_1__703_ = i[320] | i[319];
  assign t_1__702_ = i[321] | i[320];
  assign t_1__701_ = i[322] | i[321];
  assign t_1__700_ = i[323] | i[322];
  assign t_1__699_ = i[324] | i[323];
  assign t_1__698_ = i[325] | i[324];
  assign t_1__697_ = i[326] | i[325];
  assign t_1__696_ = i[327] | i[326];
  assign t_1__695_ = i[328] | i[327];
  assign t_1__694_ = i[329] | i[328];
  assign t_1__693_ = i[330] | i[329];
  assign t_1__692_ = i[331] | i[330];
  assign t_1__691_ = i[332] | i[331];
  assign t_1__690_ = i[333] | i[332];
  assign t_1__689_ = i[334] | i[333];
  assign t_1__688_ = i[335] | i[334];
  assign t_1__687_ = i[336] | i[335];
  assign t_1__686_ = i[337] | i[336];
  assign t_1__685_ = i[338] | i[337];
  assign t_1__684_ = i[339] | i[338];
  assign t_1__683_ = i[340] | i[339];
  assign t_1__682_ = i[341] | i[340];
  assign t_1__681_ = i[342] | i[341];
  assign t_1__680_ = i[343] | i[342];
  assign t_1__679_ = i[344] | i[343];
  assign t_1__678_ = i[345] | i[344];
  assign t_1__677_ = i[346] | i[345];
  assign t_1__676_ = i[347] | i[346];
  assign t_1__675_ = i[348] | i[347];
  assign t_1__674_ = i[349] | i[348];
  assign t_1__673_ = i[350] | i[349];
  assign t_1__672_ = i[351] | i[350];
  assign t_1__671_ = i[352] | i[351];
  assign t_1__670_ = i[353] | i[352];
  assign t_1__669_ = i[354] | i[353];
  assign t_1__668_ = i[355] | i[354];
  assign t_1__667_ = i[356] | i[355];
  assign t_1__666_ = i[357] | i[356];
  assign t_1__665_ = i[358] | i[357];
  assign t_1__664_ = i[359] | i[358];
  assign t_1__663_ = i[360] | i[359];
  assign t_1__662_ = i[361] | i[360];
  assign t_1__661_ = i[362] | i[361];
  assign t_1__660_ = i[363] | i[362];
  assign t_1__659_ = i[364] | i[363];
  assign t_1__658_ = i[365] | i[364];
  assign t_1__657_ = i[366] | i[365];
  assign t_1__656_ = i[367] | i[366];
  assign t_1__655_ = i[368] | i[367];
  assign t_1__654_ = i[369] | i[368];
  assign t_1__653_ = i[370] | i[369];
  assign t_1__652_ = i[371] | i[370];
  assign t_1__651_ = i[372] | i[371];
  assign t_1__650_ = i[373] | i[372];
  assign t_1__649_ = i[374] | i[373];
  assign t_1__648_ = i[375] | i[374];
  assign t_1__647_ = i[376] | i[375];
  assign t_1__646_ = i[377] | i[376];
  assign t_1__645_ = i[378] | i[377];
  assign t_1__644_ = i[379] | i[378];
  assign t_1__643_ = i[380] | i[379];
  assign t_1__642_ = i[381] | i[380];
  assign t_1__641_ = i[382] | i[381];
  assign t_1__640_ = i[383] | i[382];
  assign t_1__639_ = i[384] | i[383];
  assign t_1__638_ = i[385] | i[384];
  assign t_1__637_ = i[386] | i[385];
  assign t_1__636_ = i[387] | i[386];
  assign t_1__635_ = i[388] | i[387];
  assign t_1__634_ = i[389] | i[388];
  assign t_1__633_ = i[390] | i[389];
  assign t_1__632_ = i[391] | i[390];
  assign t_1__631_ = i[392] | i[391];
  assign t_1__630_ = i[393] | i[392];
  assign t_1__629_ = i[394] | i[393];
  assign t_1__628_ = i[395] | i[394];
  assign t_1__627_ = i[396] | i[395];
  assign t_1__626_ = i[397] | i[396];
  assign t_1__625_ = i[398] | i[397];
  assign t_1__624_ = i[399] | i[398];
  assign t_1__623_ = i[400] | i[399];
  assign t_1__622_ = i[401] | i[400];
  assign t_1__621_ = i[402] | i[401];
  assign t_1__620_ = i[403] | i[402];
  assign t_1__619_ = i[404] | i[403];
  assign t_1__618_ = i[405] | i[404];
  assign t_1__617_ = i[406] | i[405];
  assign t_1__616_ = i[407] | i[406];
  assign t_1__615_ = i[408] | i[407];
  assign t_1__614_ = i[409] | i[408];
  assign t_1__613_ = i[410] | i[409];
  assign t_1__612_ = i[411] | i[410];
  assign t_1__611_ = i[412] | i[411];
  assign t_1__610_ = i[413] | i[412];
  assign t_1__609_ = i[414] | i[413];
  assign t_1__608_ = i[415] | i[414];
  assign t_1__607_ = i[416] | i[415];
  assign t_1__606_ = i[417] | i[416];
  assign t_1__605_ = i[418] | i[417];
  assign t_1__604_ = i[419] | i[418];
  assign t_1__603_ = i[420] | i[419];
  assign t_1__602_ = i[421] | i[420];
  assign t_1__601_ = i[422] | i[421];
  assign t_1__600_ = i[423] | i[422];
  assign t_1__599_ = i[424] | i[423];
  assign t_1__598_ = i[425] | i[424];
  assign t_1__597_ = i[426] | i[425];
  assign t_1__596_ = i[427] | i[426];
  assign t_1__595_ = i[428] | i[427];
  assign t_1__594_ = i[429] | i[428];
  assign t_1__593_ = i[430] | i[429];
  assign t_1__592_ = i[431] | i[430];
  assign t_1__591_ = i[432] | i[431];
  assign t_1__590_ = i[433] | i[432];
  assign t_1__589_ = i[434] | i[433];
  assign t_1__588_ = i[435] | i[434];
  assign t_1__587_ = i[436] | i[435];
  assign t_1__586_ = i[437] | i[436];
  assign t_1__585_ = i[438] | i[437];
  assign t_1__584_ = i[439] | i[438];
  assign t_1__583_ = i[440] | i[439];
  assign t_1__582_ = i[441] | i[440];
  assign t_1__581_ = i[442] | i[441];
  assign t_1__580_ = i[443] | i[442];
  assign t_1__579_ = i[444] | i[443];
  assign t_1__578_ = i[445] | i[444];
  assign t_1__577_ = i[446] | i[445];
  assign t_1__576_ = i[447] | i[446];
  assign t_1__575_ = i[448] | i[447];
  assign t_1__574_ = i[449] | i[448];
  assign t_1__573_ = i[450] | i[449];
  assign t_1__572_ = i[451] | i[450];
  assign t_1__571_ = i[452] | i[451];
  assign t_1__570_ = i[453] | i[452];
  assign t_1__569_ = i[454] | i[453];
  assign t_1__568_ = i[455] | i[454];
  assign t_1__567_ = i[456] | i[455];
  assign t_1__566_ = i[457] | i[456];
  assign t_1__565_ = i[458] | i[457];
  assign t_1__564_ = i[459] | i[458];
  assign t_1__563_ = i[460] | i[459];
  assign t_1__562_ = i[461] | i[460];
  assign t_1__561_ = i[462] | i[461];
  assign t_1__560_ = i[463] | i[462];
  assign t_1__559_ = i[464] | i[463];
  assign t_1__558_ = i[465] | i[464];
  assign t_1__557_ = i[466] | i[465];
  assign t_1__556_ = i[467] | i[466];
  assign t_1__555_ = i[468] | i[467];
  assign t_1__554_ = i[469] | i[468];
  assign t_1__553_ = i[470] | i[469];
  assign t_1__552_ = i[471] | i[470];
  assign t_1__551_ = i[472] | i[471];
  assign t_1__550_ = i[473] | i[472];
  assign t_1__549_ = i[474] | i[473];
  assign t_1__548_ = i[475] | i[474];
  assign t_1__547_ = i[476] | i[475];
  assign t_1__546_ = i[477] | i[476];
  assign t_1__545_ = i[478] | i[477];
  assign t_1__544_ = i[479] | i[478];
  assign t_1__543_ = i[480] | i[479];
  assign t_1__542_ = i[481] | i[480];
  assign t_1__541_ = i[482] | i[481];
  assign t_1__540_ = i[483] | i[482];
  assign t_1__539_ = i[484] | i[483];
  assign t_1__538_ = i[485] | i[484];
  assign t_1__537_ = i[486] | i[485];
  assign t_1__536_ = i[487] | i[486];
  assign t_1__535_ = i[488] | i[487];
  assign t_1__534_ = i[489] | i[488];
  assign t_1__533_ = i[490] | i[489];
  assign t_1__532_ = i[491] | i[490];
  assign t_1__531_ = i[492] | i[491];
  assign t_1__530_ = i[493] | i[492];
  assign t_1__529_ = i[494] | i[493];
  assign t_1__528_ = i[495] | i[494];
  assign t_1__527_ = i[496] | i[495];
  assign t_1__526_ = i[497] | i[496];
  assign t_1__525_ = i[498] | i[497];
  assign t_1__524_ = i[499] | i[498];
  assign t_1__523_ = i[500] | i[499];
  assign t_1__522_ = i[501] | i[500];
  assign t_1__521_ = i[502] | i[501];
  assign t_1__520_ = i[503] | i[502];
  assign t_1__519_ = i[504] | i[503];
  assign t_1__518_ = i[505] | i[504];
  assign t_1__517_ = i[506] | i[505];
  assign t_1__516_ = i[507] | i[506];
  assign t_1__515_ = i[508] | i[507];
  assign t_1__514_ = i[509] | i[508];
  assign t_1__513_ = i[510] | i[509];
  assign t_1__512_ = i[511] | i[510];
  assign t_1__511_ = i[512] | i[511];
  assign t_1__510_ = i[513] | i[512];
  assign t_1__509_ = i[514] | i[513];
  assign t_1__508_ = i[515] | i[514];
  assign t_1__507_ = i[516] | i[515];
  assign t_1__506_ = i[517] | i[516];
  assign t_1__505_ = i[518] | i[517];
  assign t_1__504_ = i[519] | i[518];
  assign t_1__503_ = i[520] | i[519];
  assign t_1__502_ = i[521] | i[520];
  assign t_1__501_ = i[522] | i[521];
  assign t_1__500_ = i[523] | i[522];
  assign t_1__499_ = i[524] | i[523];
  assign t_1__498_ = i[525] | i[524];
  assign t_1__497_ = i[526] | i[525];
  assign t_1__496_ = i[527] | i[526];
  assign t_1__495_ = i[528] | i[527];
  assign t_1__494_ = i[529] | i[528];
  assign t_1__493_ = i[530] | i[529];
  assign t_1__492_ = i[531] | i[530];
  assign t_1__491_ = i[532] | i[531];
  assign t_1__490_ = i[533] | i[532];
  assign t_1__489_ = i[534] | i[533];
  assign t_1__488_ = i[535] | i[534];
  assign t_1__487_ = i[536] | i[535];
  assign t_1__486_ = i[537] | i[536];
  assign t_1__485_ = i[538] | i[537];
  assign t_1__484_ = i[539] | i[538];
  assign t_1__483_ = i[540] | i[539];
  assign t_1__482_ = i[541] | i[540];
  assign t_1__481_ = i[542] | i[541];
  assign t_1__480_ = i[543] | i[542];
  assign t_1__479_ = i[544] | i[543];
  assign t_1__478_ = i[545] | i[544];
  assign t_1__477_ = i[546] | i[545];
  assign t_1__476_ = i[547] | i[546];
  assign t_1__475_ = i[548] | i[547];
  assign t_1__474_ = i[549] | i[548];
  assign t_1__473_ = i[550] | i[549];
  assign t_1__472_ = i[551] | i[550];
  assign t_1__471_ = i[552] | i[551];
  assign t_1__470_ = i[553] | i[552];
  assign t_1__469_ = i[554] | i[553];
  assign t_1__468_ = i[555] | i[554];
  assign t_1__467_ = i[556] | i[555];
  assign t_1__466_ = i[557] | i[556];
  assign t_1__465_ = i[558] | i[557];
  assign t_1__464_ = i[559] | i[558];
  assign t_1__463_ = i[560] | i[559];
  assign t_1__462_ = i[561] | i[560];
  assign t_1__461_ = i[562] | i[561];
  assign t_1__460_ = i[563] | i[562];
  assign t_1__459_ = i[564] | i[563];
  assign t_1__458_ = i[565] | i[564];
  assign t_1__457_ = i[566] | i[565];
  assign t_1__456_ = i[567] | i[566];
  assign t_1__455_ = i[568] | i[567];
  assign t_1__454_ = i[569] | i[568];
  assign t_1__453_ = i[570] | i[569];
  assign t_1__452_ = i[571] | i[570];
  assign t_1__451_ = i[572] | i[571];
  assign t_1__450_ = i[573] | i[572];
  assign t_1__449_ = i[574] | i[573];
  assign t_1__448_ = i[575] | i[574];
  assign t_1__447_ = i[576] | i[575];
  assign t_1__446_ = i[577] | i[576];
  assign t_1__445_ = i[578] | i[577];
  assign t_1__444_ = i[579] | i[578];
  assign t_1__443_ = i[580] | i[579];
  assign t_1__442_ = i[581] | i[580];
  assign t_1__441_ = i[582] | i[581];
  assign t_1__440_ = i[583] | i[582];
  assign t_1__439_ = i[584] | i[583];
  assign t_1__438_ = i[585] | i[584];
  assign t_1__437_ = i[586] | i[585];
  assign t_1__436_ = i[587] | i[586];
  assign t_1__435_ = i[588] | i[587];
  assign t_1__434_ = i[589] | i[588];
  assign t_1__433_ = i[590] | i[589];
  assign t_1__432_ = i[591] | i[590];
  assign t_1__431_ = i[592] | i[591];
  assign t_1__430_ = i[593] | i[592];
  assign t_1__429_ = i[594] | i[593];
  assign t_1__428_ = i[595] | i[594];
  assign t_1__427_ = i[596] | i[595];
  assign t_1__426_ = i[597] | i[596];
  assign t_1__425_ = i[598] | i[597];
  assign t_1__424_ = i[599] | i[598];
  assign t_1__423_ = i[600] | i[599];
  assign t_1__422_ = i[601] | i[600];
  assign t_1__421_ = i[602] | i[601];
  assign t_1__420_ = i[603] | i[602];
  assign t_1__419_ = i[604] | i[603];
  assign t_1__418_ = i[605] | i[604];
  assign t_1__417_ = i[606] | i[605];
  assign t_1__416_ = i[607] | i[606];
  assign t_1__415_ = i[608] | i[607];
  assign t_1__414_ = i[609] | i[608];
  assign t_1__413_ = i[610] | i[609];
  assign t_1__412_ = i[611] | i[610];
  assign t_1__411_ = i[612] | i[611];
  assign t_1__410_ = i[613] | i[612];
  assign t_1__409_ = i[614] | i[613];
  assign t_1__408_ = i[615] | i[614];
  assign t_1__407_ = i[616] | i[615];
  assign t_1__406_ = i[617] | i[616];
  assign t_1__405_ = i[618] | i[617];
  assign t_1__404_ = i[619] | i[618];
  assign t_1__403_ = i[620] | i[619];
  assign t_1__402_ = i[621] | i[620];
  assign t_1__401_ = i[622] | i[621];
  assign t_1__400_ = i[623] | i[622];
  assign t_1__399_ = i[624] | i[623];
  assign t_1__398_ = i[625] | i[624];
  assign t_1__397_ = i[626] | i[625];
  assign t_1__396_ = i[627] | i[626];
  assign t_1__395_ = i[628] | i[627];
  assign t_1__394_ = i[629] | i[628];
  assign t_1__393_ = i[630] | i[629];
  assign t_1__392_ = i[631] | i[630];
  assign t_1__391_ = i[632] | i[631];
  assign t_1__390_ = i[633] | i[632];
  assign t_1__389_ = i[634] | i[633];
  assign t_1__388_ = i[635] | i[634];
  assign t_1__387_ = i[636] | i[635];
  assign t_1__386_ = i[637] | i[636];
  assign t_1__385_ = i[638] | i[637];
  assign t_1__384_ = i[639] | i[638];
  assign t_1__383_ = i[640] | i[639];
  assign t_1__382_ = i[641] | i[640];
  assign t_1__381_ = i[642] | i[641];
  assign t_1__380_ = i[643] | i[642];
  assign t_1__379_ = i[644] | i[643];
  assign t_1__378_ = i[645] | i[644];
  assign t_1__377_ = i[646] | i[645];
  assign t_1__376_ = i[647] | i[646];
  assign t_1__375_ = i[648] | i[647];
  assign t_1__374_ = i[649] | i[648];
  assign t_1__373_ = i[650] | i[649];
  assign t_1__372_ = i[651] | i[650];
  assign t_1__371_ = i[652] | i[651];
  assign t_1__370_ = i[653] | i[652];
  assign t_1__369_ = i[654] | i[653];
  assign t_1__368_ = i[655] | i[654];
  assign t_1__367_ = i[656] | i[655];
  assign t_1__366_ = i[657] | i[656];
  assign t_1__365_ = i[658] | i[657];
  assign t_1__364_ = i[659] | i[658];
  assign t_1__363_ = i[660] | i[659];
  assign t_1__362_ = i[661] | i[660];
  assign t_1__361_ = i[662] | i[661];
  assign t_1__360_ = i[663] | i[662];
  assign t_1__359_ = i[664] | i[663];
  assign t_1__358_ = i[665] | i[664];
  assign t_1__357_ = i[666] | i[665];
  assign t_1__356_ = i[667] | i[666];
  assign t_1__355_ = i[668] | i[667];
  assign t_1__354_ = i[669] | i[668];
  assign t_1__353_ = i[670] | i[669];
  assign t_1__352_ = i[671] | i[670];
  assign t_1__351_ = i[672] | i[671];
  assign t_1__350_ = i[673] | i[672];
  assign t_1__349_ = i[674] | i[673];
  assign t_1__348_ = i[675] | i[674];
  assign t_1__347_ = i[676] | i[675];
  assign t_1__346_ = i[677] | i[676];
  assign t_1__345_ = i[678] | i[677];
  assign t_1__344_ = i[679] | i[678];
  assign t_1__343_ = i[680] | i[679];
  assign t_1__342_ = i[681] | i[680];
  assign t_1__341_ = i[682] | i[681];
  assign t_1__340_ = i[683] | i[682];
  assign t_1__339_ = i[684] | i[683];
  assign t_1__338_ = i[685] | i[684];
  assign t_1__337_ = i[686] | i[685];
  assign t_1__336_ = i[687] | i[686];
  assign t_1__335_ = i[688] | i[687];
  assign t_1__334_ = i[689] | i[688];
  assign t_1__333_ = i[690] | i[689];
  assign t_1__332_ = i[691] | i[690];
  assign t_1__331_ = i[692] | i[691];
  assign t_1__330_ = i[693] | i[692];
  assign t_1__329_ = i[694] | i[693];
  assign t_1__328_ = i[695] | i[694];
  assign t_1__327_ = i[696] | i[695];
  assign t_1__326_ = i[697] | i[696];
  assign t_1__325_ = i[698] | i[697];
  assign t_1__324_ = i[699] | i[698];
  assign t_1__323_ = i[700] | i[699];
  assign t_1__322_ = i[701] | i[700];
  assign t_1__321_ = i[702] | i[701];
  assign t_1__320_ = i[703] | i[702];
  assign t_1__319_ = i[704] | i[703];
  assign t_1__318_ = i[705] | i[704];
  assign t_1__317_ = i[706] | i[705];
  assign t_1__316_ = i[707] | i[706];
  assign t_1__315_ = i[708] | i[707];
  assign t_1__314_ = i[709] | i[708];
  assign t_1__313_ = i[710] | i[709];
  assign t_1__312_ = i[711] | i[710];
  assign t_1__311_ = i[712] | i[711];
  assign t_1__310_ = i[713] | i[712];
  assign t_1__309_ = i[714] | i[713];
  assign t_1__308_ = i[715] | i[714];
  assign t_1__307_ = i[716] | i[715];
  assign t_1__306_ = i[717] | i[716];
  assign t_1__305_ = i[718] | i[717];
  assign t_1__304_ = i[719] | i[718];
  assign t_1__303_ = i[720] | i[719];
  assign t_1__302_ = i[721] | i[720];
  assign t_1__301_ = i[722] | i[721];
  assign t_1__300_ = i[723] | i[722];
  assign t_1__299_ = i[724] | i[723];
  assign t_1__298_ = i[725] | i[724];
  assign t_1__297_ = i[726] | i[725];
  assign t_1__296_ = i[727] | i[726];
  assign t_1__295_ = i[728] | i[727];
  assign t_1__294_ = i[729] | i[728];
  assign t_1__293_ = i[730] | i[729];
  assign t_1__292_ = i[731] | i[730];
  assign t_1__291_ = i[732] | i[731];
  assign t_1__290_ = i[733] | i[732];
  assign t_1__289_ = i[734] | i[733];
  assign t_1__288_ = i[735] | i[734];
  assign t_1__287_ = i[736] | i[735];
  assign t_1__286_ = i[737] | i[736];
  assign t_1__285_ = i[738] | i[737];
  assign t_1__284_ = i[739] | i[738];
  assign t_1__283_ = i[740] | i[739];
  assign t_1__282_ = i[741] | i[740];
  assign t_1__281_ = i[742] | i[741];
  assign t_1__280_ = i[743] | i[742];
  assign t_1__279_ = i[744] | i[743];
  assign t_1__278_ = i[745] | i[744];
  assign t_1__277_ = i[746] | i[745];
  assign t_1__276_ = i[747] | i[746];
  assign t_1__275_ = i[748] | i[747];
  assign t_1__274_ = i[749] | i[748];
  assign t_1__273_ = i[750] | i[749];
  assign t_1__272_ = i[751] | i[750];
  assign t_1__271_ = i[752] | i[751];
  assign t_1__270_ = i[753] | i[752];
  assign t_1__269_ = i[754] | i[753];
  assign t_1__268_ = i[755] | i[754];
  assign t_1__267_ = i[756] | i[755];
  assign t_1__266_ = i[757] | i[756];
  assign t_1__265_ = i[758] | i[757];
  assign t_1__264_ = i[759] | i[758];
  assign t_1__263_ = i[760] | i[759];
  assign t_1__262_ = i[761] | i[760];
  assign t_1__261_ = i[762] | i[761];
  assign t_1__260_ = i[763] | i[762];
  assign t_1__259_ = i[764] | i[763];
  assign t_1__258_ = i[765] | i[764];
  assign t_1__257_ = i[766] | i[765];
  assign t_1__256_ = i[767] | i[766];
  assign t_1__255_ = i[768] | i[767];
  assign t_1__254_ = i[769] | i[768];
  assign t_1__253_ = i[770] | i[769];
  assign t_1__252_ = i[771] | i[770];
  assign t_1__251_ = i[772] | i[771];
  assign t_1__250_ = i[773] | i[772];
  assign t_1__249_ = i[774] | i[773];
  assign t_1__248_ = i[775] | i[774];
  assign t_1__247_ = i[776] | i[775];
  assign t_1__246_ = i[777] | i[776];
  assign t_1__245_ = i[778] | i[777];
  assign t_1__244_ = i[779] | i[778];
  assign t_1__243_ = i[780] | i[779];
  assign t_1__242_ = i[781] | i[780];
  assign t_1__241_ = i[782] | i[781];
  assign t_1__240_ = i[783] | i[782];
  assign t_1__239_ = i[784] | i[783];
  assign t_1__238_ = i[785] | i[784];
  assign t_1__237_ = i[786] | i[785];
  assign t_1__236_ = i[787] | i[786];
  assign t_1__235_ = i[788] | i[787];
  assign t_1__234_ = i[789] | i[788];
  assign t_1__233_ = i[790] | i[789];
  assign t_1__232_ = i[791] | i[790];
  assign t_1__231_ = i[792] | i[791];
  assign t_1__230_ = i[793] | i[792];
  assign t_1__229_ = i[794] | i[793];
  assign t_1__228_ = i[795] | i[794];
  assign t_1__227_ = i[796] | i[795];
  assign t_1__226_ = i[797] | i[796];
  assign t_1__225_ = i[798] | i[797];
  assign t_1__224_ = i[799] | i[798];
  assign t_1__223_ = i[800] | i[799];
  assign t_1__222_ = i[801] | i[800];
  assign t_1__221_ = i[802] | i[801];
  assign t_1__220_ = i[803] | i[802];
  assign t_1__219_ = i[804] | i[803];
  assign t_1__218_ = i[805] | i[804];
  assign t_1__217_ = i[806] | i[805];
  assign t_1__216_ = i[807] | i[806];
  assign t_1__215_ = i[808] | i[807];
  assign t_1__214_ = i[809] | i[808];
  assign t_1__213_ = i[810] | i[809];
  assign t_1__212_ = i[811] | i[810];
  assign t_1__211_ = i[812] | i[811];
  assign t_1__210_ = i[813] | i[812];
  assign t_1__209_ = i[814] | i[813];
  assign t_1__208_ = i[815] | i[814];
  assign t_1__207_ = i[816] | i[815];
  assign t_1__206_ = i[817] | i[816];
  assign t_1__205_ = i[818] | i[817];
  assign t_1__204_ = i[819] | i[818];
  assign t_1__203_ = i[820] | i[819];
  assign t_1__202_ = i[821] | i[820];
  assign t_1__201_ = i[822] | i[821];
  assign t_1__200_ = i[823] | i[822];
  assign t_1__199_ = i[824] | i[823];
  assign t_1__198_ = i[825] | i[824];
  assign t_1__197_ = i[826] | i[825];
  assign t_1__196_ = i[827] | i[826];
  assign t_1__195_ = i[828] | i[827];
  assign t_1__194_ = i[829] | i[828];
  assign t_1__193_ = i[830] | i[829];
  assign t_1__192_ = i[831] | i[830];
  assign t_1__191_ = i[832] | i[831];
  assign t_1__190_ = i[833] | i[832];
  assign t_1__189_ = i[834] | i[833];
  assign t_1__188_ = i[835] | i[834];
  assign t_1__187_ = i[836] | i[835];
  assign t_1__186_ = i[837] | i[836];
  assign t_1__185_ = i[838] | i[837];
  assign t_1__184_ = i[839] | i[838];
  assign t_1__183_ = i[840] | i[839];
  assign t_1__182_ = i[841] | i[840];
  assign t_1__181_ = i[842] | i[841];
  assign t_1__180_ = i[843] | i[842];
  assign t_1__179_ = i[844] | i[843];
  assign t_1__178_ = i[845] | i[844];
  assign t_1__177_ = i[846] | i[845];
  assign t_1__176_ = i[847] | i[846];
  assign t_1__175_ = i[848] | i[847];
  assign t_1__174_ = i[849] | i[848];
  assign t_1__173_ = i[850] | i[849];
  assign t_1__172_ = i[851] | i[850];
  assign t_1__171_ = i[852] | i[851];
  assign t_1__170_ = i[853] | i[852];
  assign t_1__169_ = i[854] | i[853];
  assign t_1__168_ = i[855] | i[854];
  assign t_1__167_ = i[856] | i[855];
  assign t_1__166_ = i[857] | i[856];
  assign t_1__165_ = i[858] | i[857];
  assign t_1__164_ = i[859] | i[858];
  assign t_1__163_ = i[860] | i[859];
  assign t_1__162_ = i[861] | i[860];
  assign t_1__161_ = i[862] | i[861];
  assign t_1__160_ = i[863] | i[862];
  assign t_1__159_ = i[864] | i[863];
  assign t_1__158_ = i[865] | i[864];
  assign t_1__157_ = i[866] | i[865];
  assign t_1__156_ = i[867] | i[866];
  assign t_1__155_ = i[868] | i[867];
  assign t_1__154_ = i[869] | i[868];
  assign t_1__153_ = i[870] | i[869];
  assign t_1__152_ = i[871] | i[870];
  assign t_1__151_ = i[872] | i[871];
  assign t_1__150_ = i[873] | i[872];
  assign t_1__149_ = i[874] | i[873];
  assign t_1__148_ = i[875] | i[874];
  assign t_1__147_ = i[876] | i[875];
  assign t_1__146_ = i[877] | i[876];
  assign t_1__145_ = i[878] | i[877];
  assign t_1__144_ = i[879] | i[878];
  assign t_1__143_ = i[880] | i[879];
  assign t_1__142_ = i[881] | i[880];
  assign t_1__141_ = i[882] | i[881];
  assign t_1__140_ = i[883] | i[882];
  assign t_1__139_ = i[884] | i[883];
  assign t_1__138_ = i[885] | i[884];
  assign t_1__137_ = i[886] | i[885];
  assign t_1__136_ = i[887] | i[886];
  assign t_1__135_ = i[888] | i[887];
  assign t_1__134_ = i[889] | i[888];
  assign t_1__133_ = i[890] | i[889];
  assign t_1__132_ = i[891] | i[890];
  assign t_1__131_ = i[892] | i[891];
  assign t_1__130_ = i[893] | i[892];
  assign t_1__129_ = i[894] | i[893];
  assign t_1__128_ = i[895] | i[894];
  assign t_1__127_ = i[896] | i[895];
  assign t_1__126_ = i[897] | i[896];
  assign t_1__125_ = i[898] | i[897];
  assign t_1__124_ = i[899] | i[898];
  assign t_1__123_ = i[900] | i[899];
  assign t_1__122_ = i[901] | i[900];
  assign t_1__121_ = i[902] | i[901];
  assign t_1__120_ = i[903] | i[902];
  assign t_1__119_ = i[904] | i[903];
  assign t_1__118_ = i[905] | i[904];
  assign t_1__117_ = i[906] | i[905];
  assign t_1__116_ = i[907] | i[906];
  assign t_1__115_ = i[908] | i[907];
  assign t_1__114_ = i[909] | i[908];
  assign t_1__113_ = i[910] | i[909];
  assign t_1__112_ = i[911] | i[910];
  assign t_1__111_ = i[912] | i[911];
  assign t_1__110_ = i[913] | i[912];
  assign t_1__109_ = i[914] | i[913];
  assign t_1__108_ = i[915] | i[914];
  assign t_1__107_ = i[916] | i[915];
  assign t_1__106_ = i[917] | i[916];
  assign t_1__105_ = i[918] | i[917];
  assign t_1__104_ = i[919] | i[918];
  assign t_1__103_ = i[920] | i[919];
  assign t_1__102_ = i[921] | i[920];
  assign t_1__101_ = i[922] | i[921];
  assign t_1__100_ = i[923] | i[922];
  assign t_1__99_ = i[924] | i[923];
  assign t_1__98_ = i[925] | i[924];
  assign t_1__97_ = i[926] | i[925];
  assign t_1__96_ = i[927] | i[926];
  assign t_1__95_ = i[928] | i[927];
  assign t_1__94_ = i[929] | i[928];
  assign t_1__93_ = i[930] | i[929];
  assign t_1__92_ = i[931] | i[930];
  assign t_1__91_ = i[932] | i[931];
  assign t_1__90_ = i[933] | i[932];
  assign t_1__89_ = i[934] | i[933];
  assign t_1__88_ = i[935] | i[934];
  assign t_1__87_ = i[936] | i[935];
  assign t_1__86_ = i[937] | i[936];
  assign t_1__85_ = i[938] | i[937];
  assign t_1__84_ = i[939] | i[938];
  assign t_1__83_ = i[940] | i[939];
  assign t_1__82_ = i[941] | i[940];
  assign t_1__81_ = i[942] | i[941];
  assign t_1__80_ = i[943] | i[942];
  assign t_1__79_ = i[944] | i[943];
  assign t_1__78_ = i[945] | i[944];
  assign t_1__77_ = i[946] | i[945];
  assign t_1__76_ = i[947] | i[946];
  assign t_1__75_ = i[948] | i[947];
  assign t_1__74_ = i[949] | i[948];
  assign t_1__73_ = i[950] | i[949];
  assign t_1__72_ = i[951] | i[950];
  assign t_1__71_ = i[952] | i[951];
  assign t_1__70_ = i[953] | i[952];
  assign t_1__69_ = i[954] | i[953];
  assign t_1__68_ = i[955] | i[954];
  assign t_1__67_ = i[956] | i[955];
  assign t_1__66_ = i[957] | i[956];
  assign t_1__65_ = i[958] | i[957];
  assign t_1__64_ = i[959] | i[958];
  assign t_1__63_ = i[960] | i[959];
  assign t_1__62_ = i[961] | i[960];
  assign t_1__61_ = i[962] | i[961];
  assign t_1__60_ = i[963] | i[962];
  assign t_1__59_ = i[964] | i[963];
  assign t_1__58_ = i[965] | i[964];
  assign t_1__57_ = i[966] | i[965];
  assign t_1__56_ = i[967] | i[966];
  assign t_1__55_ = i[968] | i[967];
  assign t_1__54_ = i[969] | i[968];
  assign t_1__53_ = i[970] | i[969];
  assign t_1__52_ = i[971] | i[970];
  assign t_1__51_ = i[972] | i[971];
  assign t_1__50_ = i[973] | i[972];
  assign t_1__49_ = i[974] | i[973];
  assign t_1__48_ = i[975] | i[974];
  assign t_1__47_ = i[976] | i[975];
  assign t_1__46_ = i[977] | i[976];
  assign t_1__45_ = i[978] | i[977];
  assign t_1__44_ = i[979] | i[978];
  assign t_1__43_ = i[980] | i[979];
  assign t_1__42_ = i[981] | i[980];
  assign t_1__41_ = i[982] | i[981];
  assign t_1__40_ = i[983] | i[982];
  assign t_1__39_ = i[984] | i[983];
  assign t_1__38_ = i[985] | i[984];
  assign t_1__37_ = i[986] | i[985];
  assign t_1__36_ = i[987] | i[986];
  assign t_1__35_ = i[988] | i[987];
  assign t_1__34_ = i[989] | i[988];
  assign t_1__33_ = i[990] | i[989];
  assign t_1__32_ = i[991] | i[990];
  assign t_1__31_ = i[992] | i[991];
  assign t_1__30_ = i[993] | i[992];
  assign t_1__29_ = i[994] | i[993];
  assign t_1__28_ = i[995] | i[994];
  assign t_1__27_ = i[996] | i[995];
  assign t_1__26_ = i[997] | i[996];
  assign t_1__25_ = i[998] | i[997];
  assign t_1__24_ = i[999] | i[998];
  assign t_1__23_ = i[1000] | i[999];
  assign t_1__22_ = i[1001] | i[1000];
  assign t_1__21_ = i[1002] | i[1001];
  assign t_1__20_ = i[1003] | i[1002];
  assign t_1__19_ = i[1004] | i[1003];
  assign t_1__18_ = i[1005] | i[1004];
  assign t_1__17_ = i[1006] | i[1005];
  assign t_1__16_ = i[1007] | i[1006];
  assign t_1__15_ = i[1008] | i[1007];
  assign t_1__14_ = i[1009] | i[1008];
  assign t_1__13_ = i[1010] | i[1009];
  assign t_1__12_ = i[1011] | i[1010];
  assign t_1__11_ = i[1012] | i[1011];
  assign t_1__10_ = i[1013] | i[1012];
  assign t_1__9_ = i[1014] | i[1013];
  assign t_1__8_ = i[1015] | i[1014];
  assign t_1__7_ = i[1016] | i[1015];
  assign t_1__6_ = i[1017] | i[1016];
  assign t_1__5_ = i[1018] | i[1017];
  assign t_1__4_ = i[1019] | i[1018];
  assign t_1__3_ = i[1020] | i[1019];
  assign t_1__2_ = i[1021] | i[1020];
  assign t_1__1_ = i[1022] | i[1021];
  assign t_1__0_ = i[1023] | i[1022];
  assign t_2__1023_ = t_1__1023_ | 1'b0;
  assign t_2__1022_ = t_1__1022_ | 1'b0;
  assign t_2__1021_ = t_1__1021_ | t_1__1023_;
  assign t_2__1020_ = t_1__1020_ | t_1__1022_;
  assign t_2__1019_ = t_1__1019_ | t_1__1021_;
  assign t_2__1018_ = t_1__1018_ | t_1__1020_;
  assign t_2__1017_ = t_1__1017_ | t_1__1019_;
  assign t_2__1016_ = t_1__1016_ | t_1__1018_;
  assign t_2__1015_ = t_1__1015_ | t_1__1017_;
  assign t_2__1014_ = t_1__1014_ | t_1__1016_;
  assign t_2__1013_ = t_1__1013_ | t_1__1015_;
  assign t_2__1012_ = t_1__1012_ | t_1__1014_;
  assign t_2__1011_ = t_1__1011_ | t_1__1013_;
  assign t_2__1010_ = t_1__1010_ | t_1__1012_;
  assign t_2__1009_ = t_1__1009_ | t_1__1011_;
  assign t_2__1008_ = t_1__1008_ | t_1__1010_;
  assign t_2__1007_ = t_1__1007_ | t_1__1009_;
  assign t_2__1006_ = t_1__1006_ | t_1__1008_;
  assign t_2__1005_ = t_1__1005_ | t_1__1007_;
  assign t_2__1004_ = t_1__1004_ | t_1__1006_;
  assign t_2__1003_ = t_1__1003_ | t_1__1005_;
  assign t_2__1002_ = t_1__1002_ | t_1__1004_;
  assign t_2__1001_ = t_1__1001_ | t_1__1003_;
  assign t_2__1000_ = t_1__1000_ | t_1__1002_;
  assign t_2__999_ = t_1__999_ | t_1__1001_;
  assign t_2__998_ = t_1__998_ | t_1__1000_;
  assign t_2__997_ = t_1__997_ | t_1__999_;
  assign t_2__996_ = t_1__996_ | t_1__998_;
  assign t_2__995_ = t_1__995_ | t_1__997_;
  assign t_2__994_ = t_1__994_ | t_1__996_;
  assign t_2__993_ = t_1__993_ | t_1__995_;
  assign t_2__992_ = t_1__992_ | t_1__994_;
  assign t_2__991_ = t_1__991_ | t_1__993_;
  assign t_2__990_ = t_1__990_ | t_1__992_;
  assign t_2__989_ = t_1__989_ | t_1__991_;
  assign t_2__988_ = t_1__988_ | t_1__990_;
  assign t_2__987_ = t_1__987_ | t_1__989_;
  assign t_2__986_ = t_1__986_ | t_1__988_;
  assign t_2__985_ = t_1__985_ | t_1__987_;
  assign t_2__984_ = t_1__984_ | t_1__986_;
  assign t_2__983_ = t_1__983_ | t_1__985_;
  assign t_2__982_ = t_1__982_ | t_1__984_;
  assign t_2__981_ = t_1__981_ | t_1__983_;
  assign t_2__980_ = t_1__980_ | t_1__982_;
  assign t_2__979_ = t_1__979_ | t_1__981_;
  assign t_2__978_ = t_1__978_ | t_1__980_;
  assign t_2__977_ = t_1__977_ | t_1__979_;
  assign t_2__976_ = t_1__976_ | t_1__978_;
  assign t_2__975_ = t_1__975_ | t_1__977_;
  assign t_2__974_ = t_1__974_ | t_1__976_;
  assign t_2__973_ = t_1__973_ | t_1__975_;
  assign t_2__972_ = t_1__972_ | t_1__974_;
  assign t_2__971_ = t_1__971_ | t_1__973_;
  assign t_2__970_ = t_1__970_ | t_1__972_;
  assign t_2__969_ = t_1__969_ | t_1__971_;
  assign t_2__968_ = t_1__968_ | t_1__970_;
  assign t_2__967_ = t_1__967_ | t_1__969_;
  assign t_2__966_ = t_1__966_ | t_1__968_;
  assign t_2__965_ = t_1__965_ | t_1__967_;
  assign t_2__964_ = t_1__964_ | t_1__966_;
  assign t_2__963_ = t_1__963_ | t_1__965_;
  assign t_2__962_ = t_1__962_ | t_1__964_;
  assign t_2__961_ = t_1__961_ | t_1__963_;
  assign t_2__960_ = t_1__960_ | t_1__962_;
  assign t_2__959_ = t_1__959_ | t_1__961_;
  assign t_2__958_ = t_1__958_ | t_1__960_;
  assign t_2__957_ = t_1__957_ | t_1__959_;
  assign t_2__956_ = t_1__956_ | t_1__958_;
  assign t_2__955_ = t_1__955_ | t_1__957_;
  assign t_2__954_ = t_1__954_ | t_1__956_;
  assign t_2__953_ = t_1__953_ | t_1__955_;
  assign t_2__952_ = t_1__952_ | t_1__954_;
  assign t_2__951_ = t_1__951_ | t_1__953_;
  assign t_2__950_ = t_1__950_ | t_1__952_;
  assign t_2__949_ = t_1__949_ | t_1__951_;
  assign t_2__948_ = t_1__948_ | t_1__950_;
  assign t_2__947_ = t_1__947_ | t_1__949_;
  assign t_2__946_ = t_1__946_ | t_1__948_;
  assign t_2__945_ = t_1__945_ | t_1__947_;
  assign t_2__944_ = t_1__944_ | t_1__946_;
  assign t_2__943_ = t_1__943_ | t_1__945_;
  assign t_2__942_ = t_1__942_ | t_1__944_;
  assign t_2__941_ = t_1__941_ | t_1__943_;
  assign t_2__940_ = t_1__940_ | t_1__942_;
  assign t_2__939_ = t_1__939_ | t_1__941_;
  assign t_2__938_ = t_1__938_ | t_1__940_;
  assign t_2__937_ = t_1__937_ | t_1__939_;
  assign t_2__936_ = t_1__936_ | t_1__938_;
  assign t_2__935_ = t_1__935_ | t_1__937_;
  assign t_2__934_ = t_1__934_ | t_1__936_;
  assign t_2__933_ = t_1__933_ | t_1__935_;
  assign t_2__932_ = t_1__932_ | t_1__934_;
  assign t_2__931_ = t_1__931_ | t_1__933_;
  assign t_2__930_ = t_1__930_ | t_1__932_;
  assign t_2__929_ = t_1__929_ | t_1__931_;
  assign t_2__928_ = t_1__928_ | t_1__930_;
  assign t_2__927_ = t_1__927_ | t_1__929_;
  assign t_2__926_ = t_1__926_ | t_1__928_;
  assign t_2__925_ = t_1__925_ | t_1__927_;
  assign t_2__924_ = t_1__924_ | t_1__926_;
  assign t_2__923_ = t_1__923_ | t_1__925_;
  assign t_2__922_ = t_1__922_ | t_1__924_;
  assign t_2__921_ = t_1__921_ | t_1__923_;
  assign t_2__920_ = t_1__920_ | t_1__922_;
  assign t_2__919_ = t_1__919_ | t_1__921_;
  assign t_2__918_ = t_1__918_ | t_1__920_;
  assign t_2__917_ = t_1__917_ | t_1__919_;
  assign t_2__916_ = t_1__916_ | t_1__918_;
  assign t_2__915_ = t_1__915_ | t_1__917_;
  assign t_2__914_ = t_1__914_ | t_1__916_;
  assign t_2__913_ = t_1__913_ | t_1__915_;
  assign t_2__912_ = t_1__912_ | t_1__914_;
  assign t_2__911_ = t_1__911_ | t_1__913_;
  assign t_2__910_ = t_1__910_ | t_1__912_;
  assign t_2__909_ = t_1__909_ | t_1__911_;
  assign t_2__908_ = t_1__908_ | t_1__910_;
  assign t_2__907_ = t_1__907_ | t_1__909_;
  assign t_2__906_ = t_1__906_ | t_1__908_;
  assign t_2__905_ = t_1__905_ | t_1__907_;
  assign t_2__904_ = t_1__904_ | t_1__906_;
  assign t_2__903_ = t_1__903_ | t_1__905_;
  assign t_2__902_ = t_1__902_ | t_1__904_;
  assign t_2__901_ = t_1__901_ | t_1__903_;
  assign t_2__900_ = t_1__900_ | t_1__902_;
  assign t_2__899_ = t_1__899_ | t_1__901_;
  assign t_2__898_ = t_1__898_ | t_1__900_;
  assign t_2__897_ = t_1__897_ | t_1__899_;
  assign t_2__896_ = t_1__896_ | t_1__898_;
  assign t_2__895_ = t_1__895_ | t_1__897_;
  assign t_2__894_ = t_1__894_ | t_1__896_;
  assign t_2__893_ = t_1__893_ | t_1__895_;
  assign t_2__892_ = t_1__892_ | t_1__894_;
  assign t_2__891_ = t_1__891_ | t_1__893_;
  assign t_2__890_ = t_1__890_ | t_1__892_;
  assign t_2__889_ = t_1__889_ | t_1__891_;
  assign t_2__888_ = t_1__888_ | t_1__890_;
  assign t_2__887_ = t_1__887_ | t_1__889_;
  assign t_2__886_ = t_1__886_ | t_1__888_;
  assign t_2__885_ = t_1__885_ | t_1__887_;
  assign t_2__884_ = t_1__884_ | t_1__886_;
  assign t_2__883_ = t_1__883_ | t_1__885_;
  assign t_2__882_ = t_1__882_ | t_1__884_;
  assign t_2__881_ = t_1__881_ | t_1__883_;
  assign t_2__880_ = t_1__880_ | t_1__882_;
  assign t_2__879_ = t_1__879_ | t_1__881_;
  assign t_2__878_ = t_1__878_ | t_1__880_;
  assign t_2__877_ = t_1__877_ | t_1__879_;
  assign t_2__876_ = t_1__876_ | t_1__878_;
  assign t_2__875_ = t_1__875_ | t_1__877_;
  assign t_2__874_ = t_1__874_ | t_1__876_;
  assign t_2__873_ = t_1__873_ | t_1__875_;
  assign t_2__872_ = t_1__872_ | t_1__874_;
  assign t_2__871_ = t_1__871_ | t_1__873_;
  assign t_2__870_ = t_1__870_ | t_1__872_;
  assign t_2__869_ = t_1__869_ | t_1__871_;
  assign t_2__868_ = t_1__868_ | t_1__870_;
  assign t_2__867_ = t_1__867_ | t_1__869_;
  assign t_2__866_ = t_1__866_ | t_1__868_;
  assign t_2__865_ = t_1__865_ | t_1__867_;
  assign t_2__864_ = t_1__864_ | t_1__866_;
  assign t_2__863_ = t_1__863_ | t_1__865_;
  assign t_2__862_ = t_1__862_ | t_1__864_;
  assign t_2__861_ = t_1__861_ | t_1__863_;
  assign t_2__860_ = t_1__860_ | t_1__862_;
  assign t_2__859_ = t_1__859_ | t_1__861_;
  assign t_2__858_ = t_1__858_ | t_1__860_;
  assign t_2__857_ = t_1__857_ | t_1__859_;
  assign t_2__856_ = t_1__856_ | t_1__858_;
  assign t_2__855_ = t_1__855_ | t_1__857_;
  assign t_2__854_ = t_1__854_ | t_1__856_;
  assign t_2__853_ = t_1__853_ | t_1__855_;
  assign t_2__852_ = t_1__852_ | t_1__854_;
  assign t_2__851_ = t_1__851_ | t_1__853_;
  assign t_2__850_ = t_1__850_ | t_1__852_;
  assign t_2__849_ = t_1__849_ | t_1__851_;
  assign t_2__848_ = t_1__848_ | t_1__850_;
  assign t_2__847_ = t_1__847_ | t_1__849_;
  assign t_2__846_ = t_1__846_ | t_1__848_;
  assign t_2__845_ = t_1__845_ | t_1__847_;
  assign t_2__844_ = t_1__844_ | t_1__846_;
  assign t_2__843_ = t_1__843_ | t_1__845_;
  assign t_2__842_ = t_1__842_ | t_1__844_;
  assign t_2__841_ = t_1__841_ | t_1__843_;
  assign t_2__840_ = t_1__840_ | t_1__842_;
  assign t_2__839_ = t_1__839_ | t_1__841_;
  assign t_2__838_ = t_1__838_ | t_1__840_;
  assign t_2__837_ = t_1__837_ | t_1__839_;
  assign t_2__836_ = t_1__836_ | t_1__838_;
  assign t_2__835_ = t_1__835_ | t_1__837_;
  assign t_2__834_ = t_1__834_ | t_1__836_;
  assign t_2__833_ = t_1__833_ | t_1__835_;
  assign t_2__832_ = t_1__832_ | t_1__834_;
  assign t_2__831_ = t_1__831_ | t_1__833_;
  assign t_2__830_ = t_1__830_ | t_1__832_;
  assign t_2__829_ = t_1__829_ | t_1__831_;
  assign t_2__828_ = t_1__828_ | t_1__830_;
  assign t_2__827_ = t_1__827_ | t_1__829_;
  assign t_2__826_ = t_1__826_ | t_1__828_;
  assign t_2__825_ = t_1__825_ | t_1__827_;
  assign t_2__824_ = t_1__824_ | t_1__826_;
  assign t_2__823_ = t_1__823_ | t_1__825_;
  assign t_2__822_ = t_1__822_ | t_1__824_;
  assign t_2__821_ = t_1__821_ | t_1__823_;
  assign t_2__820_ = t_1__820_ | t_1__822_;
  assign t_2__819_ = t_1__819_ | t_1__821_;
  assign t_2__818_ = t_1__818_ | t_1__820_;
  assign t_2__817_ = t_1__817_ | t_1__819_;
  assign t_2__816_ = t_1__816_ | t_1__818_;
  assign t_2__815_ = t_1__815_ | t_1__817_;
  assign t_2__814_ = t_1__814_ | t_1__816_;
  assign t_2__813_ = t_1__813_ | t_1__815_;
  assign t_2__812_ = t_1__812_ | t_1__814_;
  assign t_2__811_ = t_1__811_ | t_1__813_;
  assign t_2__810_ = t_1__810_ | t_1__812_;
  assign t_2__809_ = t_1__809_ | t_1__811_;
  assign t_2__808_ = t_1__808_ | t_1__810_;
  assign t_2__807_ = t_1__807_ | t_1__809_;
  assign t_2__806_ = t_1__806_ | t_1__808_;
  assign t_2__805_ = t_1__805_ | t_1__807_;
  assign t_2__804_ = t_1__804_ | t_1__806_;
  assign t_2__803_ = t_1__803_ | t_1__805_;
  assign t_2__802_ = t_1__802_ | t_1__804_;
  assign t_2__801_ = t_1__801_ | t_1__803_;
  assign t_2__800_ = t_1__800_ | t_1__802_;
  assign t_2__799_ = t_1__799_ | t_1__801_;
  assign t_2__798_ = t_1__798_ | t_1__800_;
  assign t_2__797_ = t_1__797_ | t_1__799_;
  assign t_2__796_ = t_1__796_ | t_1__798_;
  assign t_2__795_ = t_1__795_ | t_1__797_;
  assign t_2__794_ = t_1__794_ | t_1__796_;
  assign t_2__793_ = t_1__793_ | t_1__795_;
  assign t_2__792_ = t_1__792_ | t_1__794_;
  assign t_2__791_ = t_1__791_ | t_1__793_;
  assign t_2__790_ = t_1__790_ | t_1__792_;
  assign t_2__789_ = t_1__789_ | t_1__791_;
  assign t_2__788_ = t_1__788_ | t_1__790_;
  assign t_2__787_ = t_1__787_ | t_1__789_;
  assign t_2__786_ = t_1__786_ | t_1__788_;
  assign t_2__785_ = t_1__785_ | t_1__787_;
  assign t_2__784_ = t_1__784_ | t_1__786_;
  assign t_2__783_ = t_1__783_ | t_1__785_;
  assign t_2__782_ = t_1__782_ | t_1__784_;
  assign t_2__781_ = t_1__781_ | t_1__783_;
  assign t_2__780_ = t_1__780_ | t_1__782_;
  assign t_2__779_ = t_1__779_ | t_1__781_;
  assign t_2__778_ = t_1__778_ | t_1__780_;
  assign t_2__777_ = t_1__777_ | t_1__779_;
  assign t_2__776_ = t_1__776_ | t_1__778_;
  assign t_2__775_ = t_1__775_ | t_1__777_;
  assign t_2__774_ = t_1__774_ | t_1__776_;
  assign t_2__773_ = t_1__773_ | t_1__775_;
  assign t_2__772_ = t_1__772_ | t_1__774_;
  assign t_2__771_ = t_1__771_ | t_1__773_;
  assign t_2__770_ = t_1__770_ | t_1__772_;
  assign t_2__769_ = t_1__769_ | t_1__771_;
  assign t_2__768_ = t_1__768_ | t_1__770_;
  assign t_2__767_ = t_1__767_ | t_1__769_;
  assign t_2__766_ = t_1__766_ | t_1__768_;
  assign t_2__765_ = t_1__765_ | t_1__767_;
  assign t_2__764_ = t_1__764_ | t_1__766_;
  assign t_2__763_ = t_1__763_ | t_1__765_;
  assign t_2__762_ = t_1__762_ | t_1__764_;
  assign t_2__761_ = t_1__761_ | t_1__763_;
  assign t_2__760_ = t_1__760_ | t_1__762_;
  assign t_2__759_ = t_1__759_ | t_1__761_;
  assign t_2__758_ = t_1__758_ | t_1__760_;
  assign t_2__757_ = t_1__757_ | t_1__759_;
  assign t_2__756_ = t_1__756_ | t_1__758_;
  assign t_2__755_ = t_1__755_ | t_1__757_;
  assign t_2__754_ = t_1__754_ | t_1__756_;
  assign t_2__753_ = t_1__753_ | t_1__755_;
  assign t_2__752_ = t_1__752_ | t_1__754_;
  assign t_2__751_ = t_1__751_ | t_1__753_;
  assign t_2__750_ = t_1__750_ | t_1__752_;
  assign t_2__749_ = t_1__749_ | t_1__751_;
  assign t_2__748_ = t_1__748_ | t_1__750_;
  assign t_2__747_ = t_1__747_ | t_1__749_;
  assign t_2__746_ = t_1__746_ | t_1__748_;
  assign t_2__745_ = t_1__745_ | t_1__747_;
  assign t_2__744_ = t_1__744_ | t_1__746_;
  assign t_2__743_ = t_1__743_ | t_1__745_;
  assign t_2__742_ = t_1__742_ | t_1__744_;
  assign t_2__741_ = t_1__741_ | t_1__743_;
  assign t_2__740_ = t_1__740_ | t_1__742_;
  assign t_2__739_ = t_1__739_ | t_1__741_;
  assign t_2__738_ = t_1__738_ | t_1__740_;
  assign t_2__737_ = t_1__737_ | t_1__739_;
  assign t_2__736_ = t_1__736_ | t_1__738_;
  assign t_2__735_ = t_1__735_ | t_1__737_;
  assign t_2__734_ = t_1__734_ | t_1__736_;
  assign t_2__733_ = t_1__733_ | t_1__735_;
  assign t_2__732_ = t_1__732_ | t_1__734_;
  assign t_2__731_ = t_1__731_ | t_1__733_;
  assign t_2__730_ = t_1__730_ | t_1__732_;
  assign t_2__729_ = t_1__729_ | t_1__731_;
  assign t_2__728_ = t_1__728_ | t_1__730_;
  assign t_2__727_ = t_1__727_ | t_1__729_;
  assign t_2__726_ = t_1__726_ | t_1__728_;
  assign t_2__725_ = t_1__725_ | t_1__727_;
  assign t_2__724_ = t_1__724_ | t_1__726_;
  assign t_2__723_ = t_1__723_ | t_1__725_;
  assign t_2__722_ = t_1__722_ | t_1__724_;
  assign t_2__721_ = t_1__721_ | t_1__723_;
  assign t_2__720_ = t_1__720_ | t_1__722_;
  assign t_2__719_ = t_1__719_ | t_1__721_;
  assign t_2__718_ = t_1__718_ | t_1__720_;
  assign t_2__717_ = t_1__717_ | t_1__719_;
  assign t_2__716_ = t_1__716_ | t_1__718_;
  assign t_2__715_ = t_1__715_ | t_1__717_;
  assign t_2__714_ = t_1__714_ | t_1__716_;
  assign t_2__713_ = t_1__713_ | t_1__715_;
  assign t_2__712_ = t_1__712_ | t_1__714_;
  assign t_2__711_ = t_1__711_ | t_1__713_;
  assign t_2__710_ = t_1__710_ | t_1__712_;
  assign t_2__709_ = t_1__709_ | t_1__711_;
  assign t_2__708_ = t_1__708_ | t_1__710_;
  assign t_2__707_ = t_1__707_ | t_1__709_;
  assign t_2__706_ = t_1__706_ | t_1__708_;
  assign t_2__705_ = t_1__705_ | t_1__707_;
  assign t_2__704_ = t_1__704_ | t_1__706_;
  assign t_2__703_ = t_1__703_ | t_1__705_;
  assign t_2__702_ = t_1__702_ | t_1__704_;
  assign t_2__701_ = t_1__701_ | t_1__703_;
  assign t_2__700_ = t_1__700_ | t_1__702_;
  assign t_2__699_ = t_1__699_ | t_1__701_;
  assign t_2__698_ = t_1__698_ | t_1__700_;
  assign t_2__697_ = t_1__697_ | t_1__699_;
  assign t_2__696_ = t_1__696_ | t_1__698_;
  assign t_2__695_ = t_1__695_ | t_1__697_;
  assign t_2__694_ = t_1__694_ | t_1__696_;
  assign t_2__693_ = t_1__693_ | t_1__695_;
  assign t_2__692_ = t_1__692_ | t_1__694_;
  assign t_2__691_ = t_1__691_ | t_1__693_;
  assign t_2__690_ = t_1__690_ | t_1__692_;
  assign t_2__689_ = t_1__689_ | t_1__691_;
  assign t_2__688_ = t_1__688_ | t_1__690_;
  assign t_2__687_ = t_1__687_ | t_1__689_;
  assign t_2__686_ = t_1__686_ | t_1__688_;
  assign t_2__685_ = t_1__685_ | t_1__687_;
  assign t_2__684_ = t_1__684_ | t_1__686_;
  assign t_2__683_ = t_1__683_ | t_1__685_;
  assign t_2__682_ = t_1__682_ | t_1__684_;
  assign t_2__681_ = t_1__681_ | t_1__683_;
  assign t_2__680_ = t_1__680_ | t_1__682_;
  assign t_2__679_ = t_1__679_ | t_1__681_;
  assign t_2__678_ = t_1__678_ | t_1__680_;
  assign t_2__677_ = t_1__677_ | t_1__679_;
  assign t_2__676_ = t_1__676_ | t_1__678_;
  assign t_2__675_ = t_1__675_ | t_1__677_;
  assign t_2__674_ = t_1__674_ | t_1__676_;
  assign t_2__673_ = t_1__673_ | t_1__675_;
  assign t_2__672_ = t_1__672_ | t_1__674_;
  assign t_2__671_ = t_1__671_ | t_1__673_;
  assign t_2__670_ = t_1__670_ | t_1__672_;
  assign t_2__669_ = t_1__669_ | t_1__671_;
  assign t_2__668_ = t_1__668_ | t_1__670_;
  assign t_2__667_ = t_1__667_ | t_1__669_;
  assign t_2__666_ = t_1__666_ | t_1__668_;
  assign t_2__665_ = t_1__665_ | t_1__667_;
  assign t_2__664_ = t_1__664_ | t_1__666_;
  assign t_2__663_ = t_1__663_ | t_1__665_;
  assign t_2__662_ = t_1__662_ | t_1__664_;
  assign t_2__661_ = t_1__661_ | t_1__663_;
  assign t_2__660_ = t_1__660_ | t_1__662_;
  assign t_2__659_ = t_1__659_ | t_1__661_;
  assign t_2__658_ = t_1__658_ | t_1__660_;
  assign t_2__657_ = t_1__657_ | t_1__659_;
  assign t_2__656_ = t_1__656_ | t_1__658_;
  assign t_2__655_ = t_1__655_ | t_1__657_;
  assign t_2__654_ = t_1__654_ | t_1__656_;
  assign t_2__653_ = t_1__653_ | t_1__655_;
  assign t_2__652_ = t_1__652_ | t_1__654_;
  assign t_2__651_ = t_1__651_ | t_1__653_;
  assign t_2__650_ = t_1__650_ | t_1__652_;
  assign t_2__649_ = t_1__649_ | t_1__651_;
  assign t_2__648_ = t_1__648_ | t_1__650_;
  assign t_2__647_ = t_1__647_ | t_1__649_;
  assign t_2__646_ = t_1__646_ | t_1__648_;
  assign t_2__645_ = t_1__645_ | t_1__647_;
  assign t_2__644_ = t_1__644_ | t_1__646_;
  assign t_2__643_ = t_1__643_ | t_1__645_;
  assign t_2__642_ = t_1__642_ | t_1__644_;
  assign t_2__641_ = t_1__641_ | t_1__643_;
  assign t_2__640_ = t_1__640_ | t_1__642_;
  assign t_2__639_ = t_1__639_ | t_1__641_;
  assign t_2__638_ = t_1__638_ | t_1__640_;
  assign t_2__637_ = t_1__637_ | t_1__639_;
  assign t_2__636_ = t_1__636_ | t_1__638_;
  assign t_2__635_ = t_1__635_ | t_1__637_;
  assign t_2__634_ = t_1__634_ | t_1__636_;
  assign t_2__633_ = t_1__633_ | t_1__635_;
  assign t_2__632_ = t_1__632_ | t_1__634_;
  assign t_2__631_ = t_1__631_ | t_1__633_;
  assign t_2__630_ = t_1__630_ | t_1__632_;
  assign t_2__629_ = t_1__629_ | t_1__631_;
  assign t_2__628_ = t_1__628_ | t_1__630_;
  assign t_2__627_ = t_1__627_ | t_1__629_;
  assign t_2__626_ = t_1__626_ | t_1__628_;
  assign t_2__625_ = t_1__625_ | t_1__627_;
  assign t_2__624_ = t_1__624_ | t_1__626_;
  assign t_2__623_ = t_1__623_ | t_1__625_;
  assign t_2__622_ = t_1__622_ | t_1__624_;
  assign t_2__621_ = t_1__621_ | t_1__623_;
  assign t_2__620_ = t_1__620_ | t_1__622_;
  assign t_2__619_ = t_1__619_ | t_1__621_;
  assign t_2__618_ = t_1__618_ | t_1__620_;
  assign t_2__617_ = t_1__617_ | t_1__619_;
  assign t_2__616_ = t_1__616_ | t_1__618_;
  assign t_2__615_ = t_1__615_ | t_1__617_;
  assign t_2__614_ = t_1__614_ | t_1__616_;
  assign t_2__613_ = t_1__613_ | t_1__615_;
  assign t_2__612_ = t_1__612_ | t_1__614_;
  assign t_2__611_ = t_1__611_ | t_1__613_;
  assign t_2__610_ = t_1__610_ | t_1__612_;
  assign t_2__609_ = t_1__609_ | t_1__611_;
  assign t_2__608_ = t_1__608_ | t_1__610_;
  assign t_2__607_ = t_1__607_ | t_1__609_;
  assign t_2__606_ = t_1__606_ | t_1__608_;
  assign t_2__605_ = t_1__605_ | t_1__607_;
  assign t_2__604_ = t_1__604_ | t_1__606_;
  assign t_2__603_ = t_1__603_ | t_1__605_;
  assign t_2__602_ = t_1__602_ | t_1__604_;
  assign t_2__601_ = t_1__601_ | t_1__603_;
  assign t_2__600_ = t_1__600_ | t_1__602_;
  assign t_2__599_ = t_1__599_ | t_1__601_;
  assign t_2__598_ = t_1__598_ | t_1__600_;
  assign t_2__597_ = t_1__597_ | t_1__599_;
  assign t_2__596_ = t_1__596_ | t_1__598_;
  assign t_2__595_ = t_1__595_ | t_1__597_;
  assign t_2__594_ = t_1__594_ | t_1__596_;
  assign t_2__593_ = t_1__593_ | t_1__595_;
  assign t_2__592_ = t_1__592_ | t_1__594_;
  assign t_2__591_ = t_1__591_ | t_1__593_;
  assign t_2__590_ = t_1__590_ | t_1__592_;
  assign t_2__589_ = t_1__589_ | t_1__591_;
  assign t_2__588_ = t_1__588_ | t_1__590_;
  assign t_2__587_ = t_1__587_ | t_1__589_;
  assign t_2__586_ = t_1__586_ | t_1__588_;
  assign t_2__585_ = t_1__585_ | t_1__587_;
  assign t_2__584_ = t_1__584_ | t_1__586_;
  assign t_2__583_ = t_1__583_ | t_1__585_;
  assign t_2__582_ = t_1__582_ | t_1__584_;
  assign t_2__581_ = t_1__581_ | t_1__583_;
  assign t_2__580_ = t_1__580_ | t_1__582_;
  assign t_2__579_ = t_1__579_ | t_1__581_;
  assign t_2__578_ = t_1__578_ | t_1__580_;
  assign t_2__577_ = t_1__577_ | t_1__579_;
  assign t_2__576_ = t_1__576_ | t_1__578_;
  assign t_2__575_ = t_1__575_ | t_1__577_;
  assign t_2__574_ = t_1__574_ | t_1__576_;
  assign t_2__573_ = t_1__573_ | t_1__575_;
  assign t_2__572_ = t_1__572_ | t_1__574_;
  assign t_2__571_ = t_1__571_ | t_1__573_;
  assign t_2__570_ = t_1__570_ | t_1__572_;
  assign t_2__569_ = t_1__569_ | t_1__571_;
  assign t_2__568_ = t_1__568_ | t_1__570_;
  assign t_2__567_ = t_1__567_ | t_1__569_;
  assign t_2__566_ = t_1__566_ | t_1__568_;
  assign t_2__565_ = t_1__565_ | t_1__567_;
  assign t_2__564_ = t_1__564_ | t_1__566_;
  assign t_2__563_ = t_1__563_ | t_1__565_;
  assign t_2__562_ = t_1__562_ | t_1__564_;
  assign t_2__561_ = t_1__561_ | t_1__563_;
  assign t_2__560_ = t_1__560_ | t_1__562_;
  assign t_2__559_ = t_1__559_ | t_1__561_;
  assign t_2__558_ = t_1__558_ | t_1__560_;
  assign t_2__557_ = t_1__557_ | t_1__559_;
  assign t_2__556_ = t_1__556_ | t_1__558_;
  assign t_2__555_ = t_1__555_ | t_1__557_;
  assign t_2__554_ = t_1__554_ | t_1__556_;
  assign t_2__553_ = t_1__553_ | t_1__555_;
  assign t_2__552_ = t_1__552_ | t_1__554_;
  assign t_2__551_ = t_1__551_ | t_1__553_;
  assign t_2__550_ = t_1__550_ | t_1__552_;
  assign t_2__549_ = t_1__549_ | t_1__551_;
  assign t_2__548_ = t_1__548_ | t_1__550_;
  assign t_2__547_ = t_1__547_ | t_1__549_;
  assign t_2__546_ = t_1__546_ | t_1__548_;
  assign t_2__545_ = t_1__545_ | t_1__547_;
  assign t_2__544_ = t_1__544_ | t_1__546_;
  assign t_2__543_ = t_1__543_ | t_1__545_;
  assign t_2__542_ = t_1__542_ | t_1__544_;
  assign t_2__541_ = t_1__541_ | t_1__543_;
  assign t_2__540_ = t_1__540_ | t_1__542_;
  assign t_2__539_ = t_1__539_ | t_1__541_;
  assign t_2__538_ = t_1__538_ | t_1__540_;
  assign t_2__537_ = t_1__537_ | t_1__539_;
  assign t_2__536_ = t_1__536_ | t_1__538_;
  assign t_2__535_ = t_1__535_ | t_1__537_;
  assign t_2__534_ = t_1__534_ | t_1__536_;
  assign t_2__533_ = t_1__533_ | t_1__535_;
  assign t_2__532_ = t_1__532_ | t_1__534_;
  assign t_2__531_ = t_1__531_ | t_1__533_;
  assign t_2__530_ = t_1__530_ | t_1__532_;
  assign t_2__529_ = t_1__529_ | t_1__531_;
  assign t_2__528_ = t_1__528_ | t_1__530_;
  assign t_2__527_ = t_1__527_ | t_1__529_;
  assign t_2__526_ = t_1__526_ | t_1__528_;
  assign t_2__525_ = t_1__525_ | t_1__527_;
  assign t_2__524_ = t_1__524_ | t_1__526_;
  assign t_2__523_ = t_1__523_ | t_1__525_;
  assign t_2__522_ = t_1__522_ | t_1__524_;
  assign t_2__521_ = t_1__521_ | t_1__523_;
  assign t_2__520_ = t_1__520_ | t_1__522_;
  assign t_2__519_ = t_1__519_ | t_1__521_;
  assign t_2__518_ = t_1__518_ | t_1__520_;
  assign t_2__517_ = t_1__517_ | t_1__519_;
  assign t_2__516_ = t_1__516_ | t_1__518_;
  assign t_2__515_ = t_1__515_ | t_1__517_;
  assign t_2__514_ = t_1__514_ | t_1__516_;
  assign t_2__513_ = t_1__513_ | t_1__515_;
  assign t_2__512_ = t_1__512_ | t_1__514_;
  assign t_2__511_ = t_1__511_ | t_1__513_;
  assign t_2__510_ = t_1__510_ | t_1__512_;
  assign t_2__509_ = t_1__509_ | t_1__511_;
  assign t_2__508_ = t_1__508_ | t_1__510_;
  assign t_2__507_ = t_1__507_ | t_1__509_;
  assign t_2__506_ = t_1__506_ | t_1__508_;
  assign t_2__505_ = t_1__505_ | t_1__507_;
  assign t_2__504_ = t_1__504_ | t_1__506_;
  assign t_2__503_ = t_1__503_ | t_1__505_;
  assign t_2__502_ = t_1__502_ | t_1__504_;
  assign t_2__501_ = t_1__501_ | t_1__503_;
  assign t_2__500_ = t_1__500_ | t_1__502_;
  assign t_2__499_ = t_1__499_ | t_1__501_;
  assign t_2__498_ = t_1__498_ | t_1__500_;
  assign t_2__497_ = t_1__497_ | t_1__499_;
  assign t_2__496_ = t_1__496_ | t_1__498_;
  assign t_2__495_ = t_1__495_ | t_1__497_;
  assign t_2__494_ = t_1__494_ | t_1__496_;
  assign t_2__493_ = t_1__493_ | t_1__495_;
  assign t_2__492_ = t_1__492_ | t_1__494_;
  assign t_2__491_ = t_1__491_ | t_1__493_;
  assign t_2__490_ = t_1__490_ | t_1__492_;
  assign t_2__489_ = t_1__489_ | t_1__491_;
  assign t_2__488_ = t_1__488_ | t_1__490_;
  assign t_2__487_ = t_1__487_ | t_1__489_;
  assign t_2__486_ = t_1__486_ | t_1__488_;
  assign t_2__485_ = t_1__485_ | t_1__487_;
  assign t_2__484_ = t_1__484_ | t_1__486_;
  assign t_2__483_ = t_1__483_ | t_1__485_;
  assign t_2__482_ = t_1__482_ | t_1__484_;
  assign t_2__481_ = t_1__481_ | t_1__483_;
  assign t_2__480_ = t_1__480_ | t_1__482_;
  assign t_2__479_ = t_1__479_ | t_1__481_;
  assign t_2__478_ = t_1__478_ | t_1__480_;
  assign t_2__477_ = t_1__477_ | t_1__479_;
  assign t_2__476_ = t_1__476_ | t_1__478_;
  assign t_2__475_ = t_1__475_ | t_1__477_;
  assign t_2__474_ = t_1__474_ | t_1__476_;
  assign t_2__473_ = t_1__473_ | t_1__475_;
  assign t_2__472_ = t_1__472_ | t_1__474_;
  assign t_2__471_ = t_1__471_ | t_1__473_;
  assign t_2__470_ = t_1__470_ | t_1__472_;
  assign t_2__469_ = t_1__469_ | t_1__471_;
  assign t_2__468_ = t_1__468_ | t_1__470_;
  assign t_2__467_ = t_1__467_ | t_1__469_;
  assign t_2__466_ = t_1__466_ | t_1__468_;
  assign t_2__465_ = t_1__465_ | t_1__467_;
  assign t_2__464_ = t_1__464_ | t_1__466_;
  assign t_2__463_ = t_1__463_ | t_1__465_;
  assign t_2__462_ = t_1__462_ | t_1__464_;
  assign t_2__461_ = t_1__461_ | t_1__463_;
  assign t_2__460_ = t_1__460_ | t_1__462_;
  assign t_2__459_ = t_1__459_ | t_1__461_;
  assign t_2__458_ = t_1__458_ | t_1__460_;
  assign t_2__457_ = t_1__457_ | t_1__459_;
  assign t_2__456_ = t_1__456_ | t_1__458_;
  assign t_2__455_ = t_1__455_ | t_1__457_;
  assign t_2__454_ = t_1__454_ | t_1__456_;
  assign t_2__453_ = t_1__453_ | t_1__455_;
  assign t_2__452_ = t_1__452_ | t_1__454_;
  assign t_2__451_ = t_1__451_ | t_1__453_;
  assign t_2__450_ = t_1__450_ | t_1__452_;
  assign t_2__449_ = t_1__449_ | t_1__451_;
  assign t_2__448_ = t_1__448_ | t_1__450_;
  assign t_2__447_ = t_1__447_ | t_1__449_;
  assign t_2__446_ = t_1__446_ | t_1__448_;
  assign t_2__445_ = t_1__445_ | t_1__447_;
  assign t_2__444_ = t_1__444_ | t_1__446_;
  assign t_2__443_ = t_1__443_ | t_1__445_;
  assign t_2__442_ = t_1__442_ | t_1__444_;
  assign t_2__441_ = t_1__441_ | t_1__443_;
  assign t_2__440_ = t_1__440_ | t_1__442_;
  assign t_2__439_ = t_1__439_ | t_1__441_;
  assign t_2__438_ = t_1__438_ | t_1__440_;
  assign t_2__437_ = t_1__437_ | t_1__439_;
  assign t_2__436_ = t_1__436_ | t_1__438_;
  assign t_2__435_ = t_1__435_ | t_1__437_;
  assign t_2__434_ = t_1__434_ | t_1__436_;
  assign t_2__433_ = t_1__433_ | t_1__435_;
  assign t_2__432_ = t_1__432_ | t_1__434_;
  assign t_2__431_ = t_1__431_ | t_1__433_;
  assign t_2__430_ = t_1__430_ | t_1__432_;
  assign t_2__429_ = t_1__429_ | t_1__431_;
  assign t_2__428_ = t_1__428_ | t_1__430_;
  assign t_2__427_ = t_1__427_ | t_1__429_;
  assign t_2__426_ = t_1__426_ | t_1__428_;
  assign t_2__425_ = t_1__425_ | t_1__427_;
  assign t_2__424_ = t_1__424_ | t_1__426_;
  assign t_2__423_ = t_1__423_ | t_1__425_;
  assign t_2__422_ = t_1__422_ | t_1__424_;
  assign t_2__421_ = t_1__421_ | t_1__423_;
  assign t_2__420_ = t_1__420_ | t_1__422_;
  assign t_2__419_ = t_1__419_ | t_1__421_;
  assign t_2__418_ = t_1__418_ | t_1__420_;
  assign t_2__417_ = t_1__417_ | t_1__419_;
  assign t_2__416_ = t_1__416_ | t_1__418_;
  assign t_2__415_ = t_1__415_ | t_1__417_;
  assign t_2__414_ = t_1__414_ | t_1__416_;
  assign t_2__413_ = t_1__413_ | t_1__415_;
  assign t_2__412_ = t_1__412_ | t_1__414_;
  assign t_2__411_ = t_1__411_ | t_1__413_;
  assign t_2__410_ = t_1__410_ | t_1__412_;
  assign t_2__409_ = t_1__409_ | t_1__411_;
  assign t_2__408_ = t_1__408_ | t_1__410_;
  assign t_2__407_ = t_1__407_ | t_1__409_;
  assign t_2__406_ = t_1__406_ | t_1__408_;
  assign t_2__405_ = t_1__405_ | t_1__407_;
  assign t_2__404_ = t_1__404_ | t_1__406_;
  assign t_2__403_ = t_1__403_ | t_1__405_;
  assign t_2__402_ = t_1__402_ | t_1__404_;
  assign t_2__401_ = t_1__401_ | t_1__403_;
  assign t_2__400_ = t_1__400_ | t_1__402_;
  assign t_2__399_ = t_1__399_ | t_1__401_;
  assign t_2__398_ = t_1__398_ | t_1__400_;
  assign t_2__397_ = t_1__397_ | t_1__399_;
  assign t_2__396_ = t_1__396_ | t_1__398_;
  assign t_2__395_ = t_1__395_ | t_1__397_;
  assign t_2__394_ = t_1__394_ | t_1__396_;
  assign t_2__393_ = t_1__393_ | t_1__395_;
  assign t_2__392_ = t_1__392_ | t_1__394_;
  assign t_2__391_ = t_1__391_ | t_1__393_;
  assign t_2__390_ = t_1__390_ | t_1__392_;
  assign t_2__389_ = t_1__389_ | t_1__391_;
  assign t_2__388_ = t_1__388_ | t_1__390_;
  assign t_2__387_ = t_1__387_ | t_1__389_;
  assign t_2__386_ = t_1__386_ | t_1__388_;
  assign t_2__385_ = t_1__385_ | t_1__387_;
  assign t_2__384_ = t_1__384_ | t_1__386_;
  assign t_2__383_ = t_1__383_ | t_1__385_;
  assign t_2__382_ = t_1__382_ | t_1__384_;
  assign t_2__381_ = t_1__381_ | t_1__383_;
  assign t_2__380_ = t_1__380_ | t_1__382_;
  assign t_2__379_ = t_1__379_ | t_1__381_;
  assign t_2__378_ = t_1__378_ | t_1__380_;
  assign t_2__377_ = t_1__377_ | t_1__379_;
  assign t_2__376_ = t_1__376_ | t_1__378_;
  assign t_2__375_ = t_1__375_ | t_1__377_;
  assign t_2__374_ = t_1__374_ | t_1__376_;
  assign t_2__373_ = t_1__373_ | t_1__375_;
  assign t_2__372_ = t_1__372_ | t_1__374_;
  assign t_2__371_ = t_1__371_ | t_1__373_;
  assign t_2__370_ = t_1__370_ | t_1__372_;
  assign t_2__369_ = t_1__369_ | t_1__371_;
  assign t_2__368_ = t_1__368_ | t_1__370_;
  assign t_2__367_ = t_1__367_ | t_1__369_;
  assign t_2__366_ = t_1__366_ | t_1__368_;
  assign t_2__365_ = t_1__365_ | t_1__367_;
  assign t_2__364_ = t_1__364_ | t_1__366_;
  assign t_2__363_ = t_1__363_ | t_1__365_;
  assign t_2__362_ = t_1__362_ | t_1__364_;
  assign t_2__361_ = t_1__361_ | t_1__363_;
  assign t_2__360_ = t_1__360_ | t_1__362_;
  assign t_2__359_ = t_1__359_ | t_1__361_;
  assign t_2__358_ = t_1__358_ | t_1__360_;
  assign t_2__357_ = t_1__357_ | t_1__359_;
  assign t_2__356_ = t_1__356_ | t_1__358_;
  assign t_2__355_ = t_1__355_ | t_1__357_;
  assign t_2__354_ = t_1__354_ | t_1__356_;
  assign t_2__353_ = t_1__353_ | t_1__355_;
  assign t_2__352_ = t_1__352_ | t_1__354_;
  assign t_2__351_ = t_1__351_ | t_1__353_;
  assign t_2__350_ = t_1__350_ | t_1__352_;
  assign t_2__349_ = t_1__349_ | t_1__351_;
  assign t_2__348_ = t_1__348_ | t_1__350_;
  assign t_2__347_ = t_1__347_ | t_1__349_;
  assign t_2__346_ = t_1__346_ | t_1__348_;
  assign t_2__345_ = t_1__345_ | t_1__347_;
  assign t_2__344_ = t_1__344_ | t_1__346_;
  assign t_2__343_ = t_1__343_ | t_1__345_;
  assign t_2__342_ = t_1__342_ | t_1__344_;
  assign t_2__341_ = t_1__341_ | t_1__343_;
  assign t_2__340_ = t_1__340_ | t_1__342_;
  assign t_2__339_ = t_1__339_ | t_1__341_;
  assign t_2__338_ = t_1__338_ | t_1__340_;
  assign t_2__337_ = t_1__337_ | t_1__339_;
  assign t_2__336_ = t_1__336_ | t_1__338_;
  assign t_2__335_ = t_1__335_ | t_1__337_;
  assign t_2__334_ = t_1__334_ | t_1__336_;
  assign t_2__333_ = t_1__333_ | t_1__335_;
  assign t_2__332_ = t_1__332_ | t_1__334_;
  assign t_2__331_ = t_1__331_ | t_1__333_;
  assign t_2__330_ = t_1__330_ | t_1__332_;
  assign t_2__329_ = t_1__329_ | t_1__331_;
  assign t_2__328_ = t_1__328_ | t_1__330_;
  assign t_2__327_ = t_1__327_ | t_1__329_;
  assign t_2__326_ = t_1__326_ | t_1__328_;
  assign t_2__325_ = t_1__325_ | t_1__327_;
  assign t_2__324_ = t_1__324_ | t_1__326_;
  assign t_2__323_ = t_1__323_ | t_1__325_;
  assign t_2__322_ = t_1__322_ | t_1__324_;
  assign t_2__321_ = t_1__321_ | t_1__323_;
  assign t_2__320_ = t_1__320_ | t_1__322_;
  assign t_2__319_ = t_1__319_ | t_1__321_;
  assign t_2__318_ = t_1__318_ | t_1__320_;
  assign t_2__317_ = t_1__317_ | t_1__319_;
  assign t_2__316_ = t_1__316_ | t_1__318_;
  assign t_2__315_ = t_1__315_ | t_1__317_;
  assign t_2__314_ = t_1__314_ | t_1__316_;
  assign t_2__313_ = t_1__313_ | t_1__315_;
  assign t_2__312_ = t_1__312_ | t_1__314_;
  assign t_2__311_ = t_1__311_ | t_1__313_;
  assign t_2__310_ = t_1__310_ | t_1__312_;
  assign t_2__309_ = t_1__309_ | t_1__311_;
  assign t_2__308_ = t_1__308_ | t_1__310_;
  assign t_2__307_ = t_1__307_ | t_1__309_;
  assign t_2__306_ = t_1__306_ | t_1__308_;
  assign t_2__305_ = t_1__305_ | t_1__307_;
  assign t_2__304_ = t_1__304_ | t_1__306_;
  assign t_2__303_ = t_1__303_ | t_1__305_;
  assign t_2__302_ = t_1__302_ | t_1__304_;
  assign t_2__301_ = t_1__301_ | t_1__303_;
  assign t_2__300_ = t_1__300_ | t_1__302_;
  assign t_2__299_ = t_1__299_ | t_1__301_;
  assign t_2__298_ = t_1__298_ | t_1__300_;
  assign t_2__297_ = t_1__297_ | t_1__299_;
  assign t_2__296_ = t_1__296_ | t_1__298_;
  assign t_2__295_ = t_1__295_ | t_1__297_;
  assign t_2__294_ = t_1__294_ | t_1__296_;
  assign t_2__293_ = t_1__293_ | t_1__295_;
  assign t_2__292_ = t_1__292_ | t_1__294_;
  assign t_2__291_ = t_1__291_ | t_1__293_;
  assign t_2__290_ = t_1__290_ | t_1__292_;
  assign t_2__289_ = t_1__289_ | t_1__291_;
  assign t_2__288_ = t_1__288_ | t_1__290_;
  assign t_2__287_ = t_1__287_ | t_1__289_;
  assign t_2__286_ = t_1__286_ | t_1__288_;
  assign t_2__285_ = t_1__285_ | t_1__287_;
  assign t_2__284_ = t_1__284_ | t_1__286_;
  assign t_2__283_ = t_1__283_ | t_1__285_;
  assign t_2__282_ = t_1__282_ | t_1__284_;
  assign t_2__281_ = t_1__281_ | t_1__283_;
  assign t_2__280_ = t_1__280_ | t_1__282_;
  assign t_2__279_ = t_1__279_ | t_1__281_;
  assign t_2__278_ = t_1__278_ | t_1__280_;
  assign t_2__277_ = t_1__277_ | t_1__279_;
  assign t_2__276_ = t_1__276_ | t_1__278_;
  assign t_2__275_ = t_1__275_ | t_1__277_;
  assign t_2__274_ = t_1__274_ | t_1__276_;
  assign t_2__273_ = t_1__273_ | t_1__275_;
  assign t_2__272_ = t_1__272_ | t_1__274_;
  assign t_2__271_ = t_1__271_ | t_1__273_;
  assign t_2__270_ = t_1__270_ | t_1__272_;
  assign t_2__269_ = t_1__269_ | t_1__271_;
  assign t_2__268_ = t_1__268_ | t_1__270_;
  assign t_2__267_ = t_1__267_ | t_1__269_;
  assign t_2__266_ = t_1__266_ | t_1__268_;
  assign t_2__265_ = t_1__265_ | t_1__267_;
  assign t_2__264_ = t_1__264_ | t_1__266_;
  assign t_2__263_ = t_1__263_ | t_1__265_;
  assign t_2__262_ = t_1__262_ | t_1__264_;
  assign t_2__261_ = t_1__261_ | t_1__263_;
  assign t_2__260_ = t_1__260_ | t_1__262_;
  assign t_2__259_ = t_1__259_ | t_1__261_;
  assign t_2__258_ = t_1__258_ | t_1__260_;
  assign t_2__257_ = t_1__257_ | t_1__259_;
  assign t_2__256_ = t_1__256_ | t_1__258_;
  assign t_2__255_ = t_1__255_ | t_1__257_;
  assign t_2__254_ = t_1__254_ | t_1__256_;
  assign t_2__253_ = t_1__253_ | t_1__255_;
  assign t_2__252_ = t_1__252_ | t_1__254_;
  assign t_2__251_ = t_1__251_ | t_1__253_;
  assign t_2__250_ = t_1__250_ | t_1__252_;
  assign t_2__249_ = t_1__249_ | t_1__251_;
  assign t_2__248_ = t_1__248_ | t_1__250_;
  assign t_2__247_ = t_1__247_ | t_1__249_;
  assign t_2__246_ = t_1__246_ | t_1__248_;
  assign t_2__245_ = t_1__245_ | t_1__247_;
  assign t_2__244_ = t_1__244_ | t_1__246_;
  assign t_2__243_ = t_1__243_ | t_1__245_;
  assign t_2__242_ = t_1__242_ | t_1__244_;
  assign t_2__241_ = t_1__241_ | t_1__243_;
  assign t_2__240_ = t_1__240_ | t_1__242_;
  assign t_2__239_ = t_1__239_ | t_1__241_;
  assign t_2__238_ = t_1__238_ | t_1__240_;
  assign t_2__237_ = t_1__237_ | t_1__239_;
  assign t_2__236_ = t_1__236_ | t_1__238_;
  assign t_2__235_ = t_1__235_ | t_1__237_;
  assign t_2__234_ = t_1__234_ | t_1__236_;
  assign t_2__233_ = t_1__233_ | t_1__235_;
  assign t_2__232_ = t_1__232_ | t_1__234_;
  assign t_2__231_ = t_1__231_ | t_1__233_;
  assign t_2__230_ = t_1__230_ | t_1__232_;
  assign t_2__229_ = t_1__229_ | t_1__231_;
  assign t_2__228_ = t_1__228_ | t_1__230_;
  assign t_2__227_ = t_1__227_ | t_1__229_;
  assign t_2__226_ = t_1__226_ | t_1__228_;
  assign t_2__225_ = t_1__225_ | t_1__227_;
  assign t_2__224_ = t_1__224_ | t_1__226_;
  assign t_2__223_ = t_1__223_ | t_1__225_;
  assign t_2__222_ = t_1__222_ | t_1__224_;
  assign t_2__221_ = t_1__221_ | t_1__223_;
  assign t_2__220_ = t_1__220_ | t_1__222_;
  assign t_2__219_ = t_1__219_ | t_1__221_;
  assign t_2__218_ = t_1__218_ | t_1__220_;
  assign t_2__217_ = t_1__217_ | t_1__219_;
  assign t_2__216_ = t_1__216_ | t_1__218_;
  assign t_2__215_ = t_1__215_ | t_1__217_;
  assign t_2__214_ = t_1__214_ | t_1__216_;
  assign t_2__213_ = t_1__213_ | t_1__215_;
  assign t_2__212_ = t_1__212_ | t_1__214_;
  assign t_2__211_ = t_1__211_ | t_1__213_;
  assign t_2__210_ = t_1__210_ | t_1__212_;
  assign t_2__209_ = t_1__209_ | t_1__211_;
  assign t_2__208_ = t_1__208_ | t_1__210_;
  assign t_2__207_ = t_1__207_ | t_1__209_;
  assign t_2__206_ = t_1__206_ | t_1__208_;
  assign t_2__205_ = t_1__205_ | t_1__207_;
  assign t_2__204_ = t_1__204_ | t_1__206_;
  assign t_2__203_ = t_1__203_ | t_1__205_;
  assign t_2__202_ = t_1__202_ | t_1__204_;
  assign t_2__201_ = t_1__201_ | t_1__203_;
  assign t_2__200_ = t_1__200_ | t_1__202_;
  assign t_2__199_ = t_1__199_ | t_1__201_;
  assign t_2__198_ = t_1__198_ | t_1__200_;
  assign t_2__197_ = t_1__197_ | t_1__199_;
  assign t_2__196_ = t_1__196_ | t_1__198_;
  assign t_2__195_ = t_1__195_ | t_1__197_;
  assign t_2__194_ = t_1__194_ | t_1__196_;
  assign t_2__193_ = t_1__193_ | t_1__195_;
  assign t_2__192_ = t_1__192_ | t_1__194_;
  assign t_2__191_ = t_1__191_ | t_1__193_;
  assign t_2__190_ = t_1__190_ | t_1__192_;
  assign t_2__189_ = t_1__189_ | t_1__191_;
  assign t_2__188_ = t_1__188_ | t_1__190_;
  assign t_2__187_ = t_1__187_ | t_1__189_;
  assign t_2__186_ = t_1__186_ | t_1__188_;
  assign t_2__185_ = t_1__185_ | t_1__187_;
  assign t_2__184_ = t_1__184_ | t_1__186_;
  assign t_2__183_ = t_1__183_ | t_1__185_;
  assign t_2__182_ = t_1__182_ | t_1__184_;
  assign t_2__181_ = t_1__181_ | t_1__183_;
  assign t_2__180_ = t_1__180_ | t_1__182_;
  assign t_2__179_ = t_1__179_ | t_1__181_;
  assign t_2__178_ = t_1__178_ | t_1__180_;
  assign t_2__177_ = t_1__177_ | t_1__179_;
  assign t_2__176_ = t_1__176_ | t_1__178_;
  assign t_2__175_ = t_1__175_ | t_1__177_;
  assign t_2__174_ = t_1__174_ | t_1__176_;
  assign t_2__173_ = t_1__173_ | t_1__175_;
  assign t_2__172_ = t_1__172_ | t_1__174_;
  assign t_2__171_ = t_1__171_ | t_1__173_;
  assign t_2__170_ = t_1__170_ | t_1__172_;
  assign t_2__169_ = t_1__169_ | t_1__171_;
  assign t_2__168_ = t_1__168_ | t_1__170_;
  assign t_2__167_ = t_1__167_ | t_1__169_;
  assign t_2__166_ = t_1__166_ | t_1__168_;
  assign t_2__165_ = t_1__165_ | t_1__167_;
  assign t_2__164_ = t_1__164_ | t_1__166_;
  assign t_2__163_ = t_1__163_ | t_1__165_;
  assign t_2__162_ = t_1__162_ | t_1__164_;
  assign t_2__161_ = t_1__161_ | t_1__163_;
  assign t_2__160_ = t_1__160_ | t_1__162_;
  assign t_2__159_ = t_1__159_ | t_1__161_;
  assign t_2__158_ = t_1__158_ | t_1__160_;
  assign t_2__157_ = t_1__157_ | t_1__159_;
  assign t_2__156_ = t_1__156_ | t_1__158_;
  assign t_2__155_ = t_1__155_ | t_1__157_;
  assign t_2__154_ = t_1__154_ | t_1__156_;
  assign t_2__153_ = t_1__153_ | t_1__155_;
  assign t_2__152_ = t_1__152_ | t_1__154_;
  assign t_2__151_ = t_1__151_ | t_1__153_;
  assign t_2__150_ = t_1__150_ | t_1__152_;
  assign t_2__149_ = t_1__149_ | t_1__151_;
  assign t_2__148_ = t_1__148_ | t_1__150_;
  assign t_2__147_ = t_1__147_ | t_1__149_;
  assign t_2__146_ = t_1__146_ | t_1__148_;
  assign t_2__145_ = t_1__145_ | t_1__147_;
  assign t_2__144_ = t_1__144_ | t_1__146_;
  assign t_2__143_ = t_1__143_ | t_1__145_;
  assign t_2__142_ = t_1__142_ | t_1__144_;
  assign t_2__141_ = t_1__141_ | t_1__143_;
  assign t_2__140_ = t_1__140_ | t_1__142_;
  assign t_2__139_ = t_1__139_ | t_1__141_;
  assign t_2__138_ = t_1__138_ | t_1__140_;
  assign t_2__137_ = t_1__137_ | t_1__139_;
  assign t_2__136_ = t_1__136_ | t_1__138_;
  assign t_2__135_ = t_1__135_ | t_1__137_;
  assign t_2__134_ = t_1__134_ | t_1__136_;
  assign t_2__133_ = t_1__133_ | t_1__135_;
  assign t_2__132_ = t_1__132_ | t_1__134_;
  assign t_2__131_ = t_1__131_ | t_1__133_;
  assign t_2__130_ = t_1__130_ | t_1__132_;
  assign t_2__129_ = t_1__129_ | t_1__131_;
  assign t_2__128_ = t_1__128_ | t_1__130_;
  assign t_2__127_ = t_1__127_ | t_1__129_;
  assign t_2__126_ = t_1__126_ | t_1__128_;
  assign t_2__125_ = t_1__125_ | t_1__127_;
  assign t_2__124_ = t_1__124_ | t_1__126_;
  assign t_2__123_ = t_1__123_ | t_1__125_;
  assign t_2__122_ = t_1__122_ | t_1__124_;
  assign t_2__121_ = t_1__121_ | t_1__123_;
  assign t_2__120_ = t_1__120_ | t_1__122_;
  assign t_2__119_ = t_1__119_ | t_1__121_;
  assign t_2__118_ = t_1__118_ | t_1__120_;
  assign t_2__117_ = t_1__117_ | t_1__119_;
  assign t_2__116_ = t_1__116_ | t_1__118_;
  assign t_2__115_ = t_1__115_ | t_1__117_;
  assign t_2__114_ = t_1__114_ | t_1__116_;
  assign t_2__113_ = t_1__113_ | t_1__115_;
  assign t_2__112_ = t_1__112_ | t_1__114_;
  assign t_2__111_ = t_1__111_ | t_1__113_;
  assign t_2__110_ = t_1__110_ | t_1__112_;
  assign t_2__109_ = t_1__109_ | t_1__111_;
  assign t_2__108_ = t_1__108_ | t_1__110_;
  assign t_2__107_ = t_1__107_ | t_1__109_;
  assign t_2__106_ = t_1__106_ | t_1__108_;
  assign t_2__105_ = t_1__105_ | t_1__107_;
  assign t_2__104_ = t_1__104_ | t_1__106_;
  assign t_2__103_ = t_1__103_ | t_1__105_;
  assign t_2__102_ = t_1__102_ | t_1__104_;
  assign t_2__101_ = t_1__101_ | t_1__103_;
  assign t_2__100_ = t_1__100_ | t_1__102_;
  assign t_2__99_ = t_1__99_ | t_1__101_;
  assign t_2__98_ = t_1__98_ | t_1__100_;
  assign t_2__97_ = t_1__97_ | t_1__99_;
  assign t_2__96_ = t_1__96_ | t_1__98_;
  assign t_2__95_ = t_1__95_ | t_1__97_;
  assign t_2__94_ = t_1__94_ | t_1__96_;
  assign t_2__93_ = t_1__93_ | t_1__95_;
  assign t_2__92_ = t_1__92_ | t_1__94_;
  assign t_2__91_ = t_1__91_ | t_1__93_;
  assign t_2__90_ = t_1__90_ | t_1__92_;
  assign t_2__89_ = t_1__89_ | t_1__91_;
  assign t_2__88_ = t_1__88_ | t_1__90_;
  assign t_2__87_ = t_1__87_ | t_1__89_;
  assign t_2__86_ = t_1__86_ | t_1__88_;
  assign t_2__85_ = t_1__85_ | t_1__87_;
  assign t_2__84_ = t_1__84_ | t_1__86_;
  assign t_2__83_ = t_1__83_ | t_1__85_;
  assign t_2__82_ = t_1__82_ | t_1__84_;
  assign t_2__81_ = t_1__81_ | t_1__83_;
  assign t_2__80_ = t_1__80_ | t_1__82_;
  assign t_2__79_ = t_1__79_ | t_1__81_;
  assign t_2__78_ = t_1__78_ | t_1__80_;
  assign t_2__77_ = t_1__77_ | t_1__79_;
  assign t_2__76_ = t_1__76_ | t_1__78_;
  assign t_2__75_ = t_1__75_ | t_1__77_;
  assign t_2__74_ = t_1__74_ | t_1__76_;
  assign t_2__73_ = t_1__73_ | t_1__75_;
  assign t_2__72_ = t_1__72_ | t_1__74_;
  assign t_2__71_ = t_1__71_ | t_1__73_;
  assign t_2__70_ = t_1__70_ | t_1__72_;
  assign t_2__69_ = t_1__69_ | t_1__71_;
  assign t_2__68_ = t_1__68_ | t_1__70_;
  assign t_2__67_ = t_1__67_ | t_1__69_;
  assign t_2__66_ = t_1__66_ | t_1__68_;
  assign t_2__65_ = t_1__65_ | t_1__67_;
  assign t_2__64_ = t_1__64_ | t_1__66_;
  assign t_2__63_ = t_1__63_ | t_1__65_;
  assign t_2__62_ = t_1__62_ | t_1__64_;
  assign t_2__61_ = t_1__61_ | t_1__63_;
  assign t_2__60_ = t_1__60_ | t_1__62_;
  assign t_2__59_ = t_1__59_ | t_1__61_;
  assign t_2__58_ = t_1__58_ | t_1__60_;
  assign t_2__57_ = t_1__57_ | t_1__59_;
  assign t_2__56_ = t_1__56_ | t_1__58_;
  assign t_2__55_ = t_1__55_ | t_1__57_;
  assign t_2__54_ = t_1__54_ | t_1__56_;
  assign t_2__53_ = t_1__53_ | t_1__55_;
  assign t_2__52_ = t_1__52_ | t_1__54_;
  assign t_2__51_ = t_1__51_ | t_1__53_;
  assign t_2__50_ = t_1__50_ | t_1__52_;
  assign t_2__49_ = t_1__49_ | t_1__51_;
  assign t_2__48_ = t_1__48_ | t_1__50_;
  assign t_2__47_ = t_1__47_ | t_1__49_;
  assign t_2__46_ = t_1__46_ | t_1__48_;
  assign t_2__45_ = t_1__45_ | t_1__47_;
  assign t_2__44_ = t_1__44_ | t_1__46_;
  assign t_2__43_ = t_1__43_ | t_1__45_;
  assign t_2__42_ = t_1__42_ | t_1__44_;
  assign t_2__41_ = t_1__41_ | t_1__43_;
  assign t_2__40_ = t_1__40_ | t_1__42_;
  assign t_2__39_ = t_1__39_ | t_1__41_;
  assign t_2__38_ = t_1__38_ | t_1__40_;
  assign t_2__37_ = t_1__37_ | t_1__39_;
  assign t_2__36_ = t_1__36_ | t_1__38_;
  assign t_2__35_ = t_1__35_ | t_1__37_;
  assign t_2__34_ = t_1__34_ | t_1__36_;
  assign t_2__33_ = t_1__33_ | t_1__35_;
  assign t_2__32_ = t_1__32_ | t_1__34_;
  assign t_2__31_ = t_1__31_ | t_1__33_;
  assign t_2__30_ = t_1__30_ | t_1__32_;
  assign t_2__29_ = t_1__29_ | t_1__31_;
  assign t_2__28_ = t_1__28_ | t_1__30_;
  assign t_2__27_ = t_1__27_ | t_1__29_;
  assign t_2__26_ = t_1__26_ | t_1__28_;
  assign t_2__25_ = t_1__25_ | t_1__27_;
  assign t_2__24_ = t_1__24_ | t_1__26_;
  assign t_2__23_ = t_1__23_ | t_1__25_;
  assign t_2__22_ = t_1__22_ | t_1__24_;
  assign t_2__21_ = t_1__21_ | t_1__23_;
  assign t_2__20_ = t_1__20_ | t_1__22_;
  assign t_2__19_ = t_1__19_ | t_1__21_;
  assign t_2__18_ = t_1__18_ | t_1__20_;
  assign t_2__17_ = t_1__17_ | t_1__19_;
  assign t_2__16_ = t_1__16_ | t_1__18_;
  assign t_2__15_ = t_1__15_ | t_1__17_;
  assign t_2__14_ = t_1__14_ | t_1__16_;
  assign t_2__13_ = t_1__13_ | t_1__15_;
  assign t_2__12_ = t_1__12_ | t_1__14_;
  assign t_2__11_ = t_1__11_ | t_1__13_;
  assign t_2__10_ = t_1__10_ | t_1__12_;
  assign t_2__9_ = t_1__9_ | t_1__11_;
  assign t_2__8_ = t_1__8_ | t_1__10_;
  assign t_2__7_ = t_1__7_ | t_1__9_;
  assign t_2__6_ = t_1__6_ | t_1__8_;
  assign t_2__5_ = t_1__5_ | t_1__7_;
  assign t_2__4_ = t_1__4_ | t_1__6_;
  assign t_2__3_ = t_1__3_ | t_1__5_;
  assign t_2__2_ = t_1__2_ | t_1__4_;
  assign t_2__1_ = t_1__1_ | t_1__3_;
  assign t_2__0_ = t_1__0_ | t_1__2_;
  assign t_3__1023_ = t_2__1023_ | 1'b0;
  assign t_3__1022_ = t_2__1022_ | 1'b0;
  assign t_3__1021_ = t_2__1021_ | 1'b0;
  assign t_3__1020_ = t_2__1020_ | 1'b0;
  assign t_3__1019_ = t_2__1019_ | t_2__1023_;
  assign t_3__1018_ = t_2__1018_ | t_2__1022_;
  assign t_3__1017_ = t_2__1017_ | t_2__1021_;
  assign t_3__1016_ = t_2__1016_ | t_2__1020_;
  assign t_3__1015_ = t_2__1015_ | t_2__1019_;
  assign t_3__1014_ = t_2__1014_ | t_2__1018_;
  assign t_3__1013_ = t_2__1013_ | t_2__1017_;
  assign t_3__1012_ = t_2__1012_ | t_2__1016_;
  assign t_3__1011_ = t_2__1011_ | t_2__1015_;
  assign t_3__1010_ = t_2__1010_ | t_2__1014_;
  assign t_3__1009_ = t_2__1009_ | t_2__1013_;
  assign t_3__1008_ = t_2__1008_ | t_2__1012_;
  assign t_3__1007_ = t_2__1007_ | t_2__1011_;
  assign t_3__1006_ = t_2__1006_ | t_2__1010_;
  assign t_3__1005_ = t_2__1005_ | t_2__1009_;
  assign t_3__1004_ = t_2__1004_ | t_2__1008_;
  assign t_3__1003_ = t_2__1003_ | t_2__1007_;
  assign t_3__1002_ = t_2__1002_ | t_2__1006_;
  assign t_3__1001_ = t_2__1001_ | t_2__1005_;
  assign t_3__1000_ = t_2__1000_ | t_2__1004_;
  assign t_3__999_ = t_2__999_ | t_2__1003_;
  assign t_3__998_ = t_2__998_ | t_2__1002_;
  assign t_3__997_ = t_2__997_ | t_2__1001_;
  assign t_3__996_ = t_2__996_ | t_2__1000_;
  assign t_3__995_ = t_2__995_ | t_2__999_;
  assign t_3__994_ = t_2__994_ | t_2__998_;
  assign t_3__993_ = t_2__993_ | t_2__997_;
  assign t_3__992_ = t_2__992_ | t_2__996_;
  assign t_3__991_ = t_2__991_ | t_2__995_;
  assign t_3__990_ = t_2__990_ | t_2__994_;
  assign t_3__989_ = t_2__989_ | t_2__993_;
  assign t_3__988_ = t_2__988_ | t_2__992_;
  assign t_3__987_ = t_2__987_ | t_2__991_;
  assign t_3__986_ = t_2__986_ | t_2__990_;
  assign t_3__985_ = t_2__985_ | t_2__989_;
  assign t_3__984_ = t_2__984_ | t_2__988_;
  assign t_3__983_ = t_2__983_ | t_2__987_;
  assign t_3__982_ = t_2__982_ | t_2__986_;
  assign t_3__981_ = t_2__981_ | t_2__985_;
  assign t_3__980_ = t_2__980_ | t_2__984_;
  assign t_3__979_ = t_2__979_ | t_2__983_;
  assign t_3__978_ = t_2__978_ | t_2__982_;
  assign t_3__977_ = t_2__977_ | t_2__981_;
  assign t_3__976_ = t_2__976_ | t_2__980_;
  assign t_3__975_ = t_2__975_ | t_2__979_;
  assign t_3__974_ = t_2__974_ | t_2__978_;
  assign t_3__973_ = t_2__973_ | t_2__977_;
  assign t_3__972_ = t_2__972_ | t_2__976_;
  assign t_3__971_ = t_2__971_ | t_2__975_;
  assign t_3__970_ = t_2__970_ | t_2__974_;
  assign t_3__969_ = t_2__969_ | t_2__973_;
  assign t_3__968_ = t_2__968_ | t_2__972_;
  assign t_3__967_ = t_2__967_ | t_2__971_;
  assign t_3__966_ = t_2__966_ | t_2__970_;
  assign t_3__965_ = t_2__965_ | t_2__969_;
  assign t_3__964_ = t_2__964_ | t_2__968_;
  assign t_3__963_ = t_2__963_ | t_2__967_;
  assign t_3__962_ = t_2__962_ | t_2__966_;
  assign t_3__961_ = t_2__961_ | t_2__965_;
  assign t_3__960_ = t_2__960_ | t_2__964_;
  assign t_3__959_ = t_2__959_ | t_2__963_;
  assign t_3__958_ = t_2__958_ | t_2__962_;
  assign t_3__957_ = t_2__957_ | t_2__961_;
  assign t_3__956_ = t_2__956_ | t_2__960_;
  assign t_3__955_ = t_2__955_ | t_2__959_;
  assign t_3__954_ = t_2__954_ | t_2__958_;
  assign t_3__953_ = t_2__953_ | t_2__957_;
  assign t_3__952_ = t_2__952_ | t_2__956_;
  assign t_3__951_ = t_2__951_ | t_2__955_;
  assign t_3__950_ = t_2__950_ | t_2__954_;
  assign t_3__949_ = t_2__949_ | t_2__953_;
  assign t_3__948_ = t_2__948_ | t_2__952_;
  assign t_3__947_ = t_2__947_ | t_2__951_;
  assign t_3__946_ = t_2__946_ | t_2__950_;
  assign t_3__945_ = t_2__945_ | t_2__949_;
  assign t_3__944_ = t_2__944_ | t_2__948_;
  assign t_3__943_ = t_2__943_ | t_2__947_;
  assign t_3__942_ = t_2__942_ | t_2__946_;
  assign t_3__941_ = t_2__941_ | t_2__945_;
  assign t_3__940_ = t_2__940_ | t_2__944_;
  assign t_3__939_ = t_2__939_ | t_2__943_;
  assign t_3__938_ = t_2__938_ | t_2__942_;
  assign t_3__937_ = t_2__937_ | t_2__941_;
  assign t_3__936_ = t_2__936_ | t_2__940_;
  assign t_3__935_ = t_2__935_ | t_2__939_;
  assign t_3__934_ = t_2__934_ | t_2__938_;
  assign t_3__933_ = t_2__933_ | t_2__937_;
  assign t_3__932_ = t_2__932_ | t_2__936_;
  assign t_3__931_ = t_2__931_ | t_2__935_;
  assign t_3__930_ = t_2__930_ | t_2__934_;
  assign t_3__929_ = t_2__929_ | t_2__933_;
  assign t_3__928_ = t_2__928_ | t_2__932_;
  assign t_3__927_ = t_2__927_ | t_2__931_;
  assign t_3__926_ = t_2__926_ | t_2__930_;
  assign t_3__925_ = t_2__925_ | t_2__929_;
  assign t_3__924_ = t_2__924_ | t_2__928_;
  assign t_3__923_ = t_2__923_ | t_2__927_;
  assign t_3__922_ = t_2__922_ | t_2__926_;
  assign t_3__921_ = t_2__921_ | t_2__925_;
  assign t_3__920_ = t_2__920_ | t_2__924_;
  assign t_3__919_ = t_2__919_ | t_2__923_;
  assign t_3__918_ = t_2__918_ | t_2__922_;
  assign t_3__917_ = t_2__917_ | t_2__921_;
  assign t_3__916_ = t_2__916_ | t_2__920_;
  assign t_3__915_ = t_2__915_ | t_2__919_;
  assign t_3__914_ = t_2__914_ | t_2__918_;
  assign t_3__913_ = t_2__913_ | t_2__917_;
  assign t_3__912_ = t_2__912_ | t_2__916_;
  assign t_3__911_ = t_2__911_ | t_2__915_;
  assign t_3__910_ = t_2__910_ | t_2__914_;
  assign t_3__909_ = t_2__909_ | t_2__913_;
  assign t_3__908_ = t_2__908_ | t_2__912_;
  assign t_3__907_ = t_2__907_ | t_2__911_;
  assign t_3__906_ = t_2__906_ | t_2__910_;
  assign t_3__905_ = t_2__905_ | t_2__909_;
  assign t_3__904_ = t_2__904_ | t_2__908_;
  assign t_3__903_ = t_2__903_ | t_2__907_;
  assign t_3__902_ = t_2__902_ | t_2__906_;
  assign t_3__901_ = t_2__901_ | t_2__905_;
  assign t_3__900_ = t_2__900_ | t_2__904_;
  assign t_3__899_ = t_2__899_ | t_2__903_;
  assign t_3__898_ = t_2__898_ | t_2__902_;
  assign t_3__897_ = t_2__897_ | t_2__901_;
  assign t_3__896_ = t_2__896_ | t_2__900_;
  assign t_3__895_ = t_2__895_ | t_2__899_;
  assign t_3__894_ = t_2__894_ | t_2__898_;
  assign t_3__893_ = t_2__893_ | t_2__897_;
  assign t_3__892_ = t_2__892_ | t_2__896_;
  assign t_3__891_ = t_2__891_ | t_2__895_;
  assign t_3__890_ = t_2__890_ | t_2__894_;
  assign t_3__889_ = t_2__889_ | t_2__893_;
  assign t_3__888_ = t_2__888_ | t_2__892_;
  assign t_3__887_ = t_2__887_ | t_2__891_;
  assign t_3__886_ = t_2__886_ | t_2__890_;
  assign t_3__885_ = t_2__885_ | t_2__889_;
  assign t_3__884_ = t_2__884_ | t_2__888_;
  assign t_3__883_ = t_2__883_ | t_2__887_;
  assign t_3__882_ = t_2__882_ | t_2__886_;
  assign t_3__881_ = t_2__881_ | t_2__885_;
  assign t_3__880_ = t_2__880_ | t_2__884_;
  assign t_3__879_ = t_2__879_ | t_2__883_;
  assign t_3__878_ = t_2__878_ | t_2__882_;
  assign t_3__877_ = t_2__877_ | t_2__881_;
  assign t_3__876_ = t_2__876_ | t_2__880_;
  assign t_3__875_ = t_2__875_ | t_2__879_;
  assign t_3__874_ = t_2__874_ | t_2__878_;
  assign t_3__873_ = t_2__873_ | t_2__877_;
  assign t_3__872_ = t_2__872_ | t_2__876_;
  assign t_3__871_ = t_2__871_ | t_2__875_;
  assign t_3__870_ = t_2__870_ | t_2__874_;
  assign t_3__869_ = t_2__869_ | t_2__873_;
  assign t_3__868_ = t_2__868_ | t_2__872_;
  assign t_3__867_ = t_2__867_ | t_2__871_;
  assign t_3__866_ = t_2__866_ | t_2__870_;
  assign t_3__865_ = t_2__865_ | t_2__869_;
  assign t_3__864_ = t_2__864_ | t_2__868_;
  assign t_3__863_ = t_2__863_ | t_2__867_;
  assign t_3__862_ = t_2__862_ | t_2__866_;
  assign t_3__861_ = t_2__861_ | t_2__865_;
  assign t_3__860_ = t_2__860_ | t_2__864_;
  assign t_3__859_ = t_2__859_ | t_2__863_;
  assign t_3__858_ = t_2__858_ | t_2__862_;
  assign t_3__857_ = t_2__857_ | t_2__861_;
  assign t_3__856_ = t_2__856_ | t_2__860_;
  assign t_3__855_ = t_2__855_ | t_2__859_;
  assign t_3__854_ = t_2__854_ | t_2__858_;
  assign t_3__853_ = t_2__853_ | t_2__857_;
  assign t_3__852_ = t_2__852_ | t_2__856_;
  assign t_3__851_ = t_2__851_ | t_2__855_;
  assign t_3__850_ = t_2__850_ | t_2__854_;
  assign t_3__849_ = t_2__849_ | t_2__853_;
  assign t_3__848_ = t_2__848_ | t_2__852_;
  assign t_3__847_ = t_2__847_ | t_2__851_;
  assign t_3__846_ = t_2__846_ | t_2__850_;
  assign t_3__845_ = t_2__845_ | t_2__849_;
  assign t_3__844_ = t_2__844_ | t_2__848_;
  assign t_3__843_ = t_2__843_ | t_2__847_;
  assign t_3__842_ = t_2__842_ | t_2__846_;
  assign t_3__841_ = t_2__841_ | t_2__845_;
  assign t_3__840_ = t_2__840_ | t_2__844_;
  assign t_3__839_ = t_2__839_ | t_2__843_;
  assign t_3__838_ = t_2__838_ | t_2__842_;
  assign t_3__837_ = t_2__837_ | t_2__841_;
  assign t_3__836_ = t_2__836_ | t_2__840_;
  assign t_3__835_ = t_2__835_ | t_2__839_;
  assign t_3__834_ = t_2__834_ | t_2__838_;
  assign t_3__833_ = t_2__833_ | t_2__837_;
  assign t_3__832_ = t_2__832_ | t_2__836_;
  assign t_3__831_ = t_2__831_ | t_2__835_;
  assign t_3__830_ = t_2__830_ | t_2__834_;
  assign t_3__829_ = t_2__829_ | t_2__833_;
  assign t_3__828_ = t_2__828_ | t_2__832_;
  assign t_3__827_ = t_2__827_ | t_2__831_;
  assign t_3__826_ = t_2__826_ | t_2__830_;
  assign t_3__825_ = t_2__825_ | t_2__829_;
  assign t_3__824_ = t_2__824_ | t_2__828_;
  assign t_3__823_ = t_2__823_ | t_2__827_;
  assign t_3__822_ = t_2__822_ | t_2__826_;
  assign t_3__821_ = t_2__821_ | t_2__825_;
  assign t_3__820_ = t_2__820_ | t_2__824_;
  assign t_3__819_ = t_2__819_ | t_2__823_;
  assign t_3__818_ = t_2__818_ | t_2__822_;
  assign t_3__817_ = t_2__817_ | t_2__821_;
  assign t_3__816_ = t_2__816_ | t_2__820_;
  assign t_3__815_ = t_2__815_ | t_2__819_;
  assign t_3__814_ = t_2__814_ | t_2__818_;
  assign t_3__813_ = t_2__813_ | t_2__817_;
  assign t_3__812_ = t_2__812_ | t_2__816_;
  assign t_3__811_ = t_2__811_ | t_2__815_;
  assign t_3__810_ = t_2__810_ | t_2__814_;
  assign t_3__809_ = t_2__809_ | t_2__813_;
  assign t_3__808_ = t_2__808_ | t_2__812_;
  assign t_3__807_ = t_2__807_ | t_2__811_;
  assign t_3__806_ = t_2__806_ | t_2__810_;
  assign t_3__805_ = t_2__805_ | t_2__809_;
  assign t_3__804_ = t_2__804_ | t_2__808_;
  assign t_3__803_ = t_2__803_ | t_2__807_;
  assign t_3__802_ = t_2__802_ | t_2__806_;
  assign t_3__801_ = t_2__801_ | t_2__805_;
  assign t_3__800_ = t_2__800_ | t_2__804_;
  assign t_3__799_ = t_2__799_ | t_2__803_;
  assign t_3__798_ = t_2__798_ | t_2__802_;
  assign t_3__797_ = t_2__797_ | t_2__801_;
  assign t_3__796_ = t_2__796_ | t_2__800_;
  assign t_3__795_ = t_2__795_ | t_2__799_;
  assign t_3__794_ = t_2__794_ | t_2__798_;
  assign t_3__793_ = t_2__793_ | t_2__797_;
  assign t_3__792_ = t_2__792_ | t_2__796_;
  assign t_3__791_ = t_2__791_ | t_2__795_;
  assign t_3__790_ = t_2__790_ | t_2__794_;
  assign t_3__789_ = t_2__789_ | t_2__793_;
  assign t_3__788_ = t_2__788_ | t_2__792_;
  assign t_3__787_ = t_2__787_ | t_2__791_;
  assign t_3__786_ = t_2__786_ | t_2__790_;
  assign t_3__785_ = t_2__785_ | t_2__789_;
  assign t_3__784_ = t_2__784_ | t_2__788_;
  assign t_3__783_ = t_2__783_ | t_2__787_;
  assign t_3__782_ = t_2__782_ | t_2__786_;
  assign t_3__781_ = t_2__781_ | t_2__785_;
  assign t_3__780_ = t_2__780_ | t_2__784_;
  assign t_3__779_ = t_2__779_ | t_2__783_;
  assign t_3__778_ = t_2__778_ | t_2__782_;
  assign t_3__777_ = t_2__777_ | t_2__781_;
  assign t_3__776_ = t_2__776_ | t_2__780_;
  assign t_3__775_ = t_2__775_ | t_2__779_;
  assign t_3__774_ = t_2__774_ | t_2__778_;
  assign t_3__773_ = t_2__773_ | t_2__777_;
  assign t_3__772_ = t_2__772_ | t_2__776_;
  assign t_3__771_ = t_2__771_ | t_2__775_;
  assign t_3__770_ = t_2__770_ | t_2__774_;
  assign t_3__769_ = t_2__769_ | t_2__773_;
  assign t_3__768_ = t_2__768_ | t_2__772_;
  assign t_3__767_ = t_2__767_ | t_2__771_;
  assign t_3__766_ = t_2__766_ | t_2__770_;
  assign t_3__765_ = t_2__765_ | t_2__769_;
  assign t_3__764_ = t_2__764_ | t_2__768_;
  assign t_3__763_ = t_2__763_ | t_2__767_;
  assign t_3__762_ = t_2__762_ | t_2__766_;
  assign t_3__761_ = t_2__761_ | t_2__765_;
  assign t_3__760_ = t_2__760_ | t_2__764_;
  assign t_3__759_ = t_2__759_ | t_2__763_;
  assign t_3__758_ = t_2__758_ | t_2__762_;
  assign t_3__757_ = t_2__757_ | t_2__761_;
  assign t_3__756_ = t_2__756_ | t_2__760_;
  assign t_3__755_ = t_2__755_ | t_2__759_;
  assign t_3__754_ = t_2__754_ | t_2__758_;
  assign t_3__753_ = t_2__753_ | t_2__757_;
  assign t_3__752_ = t_2__752_ | t_2__756_;
  assign t_3__751_ = t_2__751_ | t_2__755_;
  assign t_3__750_ = t_2__750_ | t_2__754_;
  assign t_3__749_ = t_2__749_ | t_2__753_;
  assign t_3__748_ = t_2__748_ | t_2__752_;
  assign t_3__747_ = t_2__747_ | t_2__751_;
  assign t_3__746_ = t_2__746_ | t_2__750_;
  assign t_3__745_ = t_2__745_ | t_2__749_;
  assign t_3__744_ = t_2__744_ | t_2__748_;
  assign t_3__743_ = t_2__743_ | t_2__747_;
  assign t_3__742_ = t_2__742_ | t_2__746_;
  assign t_3__741_ = t_2__741_ | t_2__745_;
  assign t_3__740_ = t_2__740_ | t_2__744_;
  assign t_3__739_ = t_2__739_ | t_2__743_;
  assign t_3__738_ = t_2__738_ | t_2__742_;
  assign t_3__737_ = t_2__737_ | t_2__741_;
  assign t_3__736_ = t_2__736_ | t_2__740_;
  assign t_3__735_ = t_2__735_ | t_2__739_;
  assign t_3__734_ = t_2__734_ | t_2__738_;
  assign t_3__733_ = t_2__733_ | t_2__737_;
  assign t_3__732_ = t_2__732_ | t_2__736_;
  assign t_3__731_ = t_2__731_ | t_2__735_;
  assign t_3__730_ = t_2__730_ | t_2__734_;
  assign t_3__729_ = t_2__729_ | t_2__733_;
  assign t_3__728_ = t_2__728_ | t_2__732_;
  assign t_3__727_ = t_2__727_ | t_2__731_;
  assign t_3__726_ = t_2__726_ | t_2__730_;
  assign t_3__725_ = t_2__725_ | t_2__729_;
  assign t_3__724_ = t_2__724_ | t_2__728_;
  assign t_3__723_ = t_2__723_ | t_2__727_;
  assign t_3__722_ = t_2__722_ | t_2__726_;
  assign t_3__721_ = t_2__721_ | t_2__725_;
  assign t_3__720_ = t_2__720_ | t_2__724_;
  assign t_3__719_ = t_2__719_ | t_2__723_;
  assign t_3__718_ = t_2__718_ | t_2__722_;
  assign t_3__717_ = t_2__717_ | t_2__721_;
  assign t_3__716_ = t_2__716_ | t_2__720_;
  assign t_3__715_ = t_2__715_ | t_2__719_;
  assign t_3__714_ = t_2__714_ | t_2__718_;
  assign t_3__713_ = t_2__713_ | t_2__717_;
  assign t_3__712_ = t_2__712_ | t_2__716_;
  assign t_3__711_ = t_2__711_ | t_2__715_;
  assign t_3__710_ = t_2__710_ | t_2__714_;
  assign t_3__709_ = t_2__709_ | t_2__713_;
  assign t_3__708_ = t_2__708_ | t_2__712_;
  assign t_3__707_ = t_2__707_ | t_2__711_;
  assign t_3__706_ = t_2__706_ | t_2__710_;
  assign t_3__705_ = t_2__705_ | t_2__709_;
  assign t_3__704_ = t_2__704_ | t_2__708_;
  assign t_3__703_ = t_2__703_ | t_2__707_;
  assign t_3__702_ = t_2__702_ | t_2__706_;
  assign t_3__701_ = t_2__701_ | t_2__705_;
  assign t_3__700_ = t_2__700_ | t_2__704_;
  assign t_3__699_ = t_2__699_ | t_2__703_;
  assign t_3__698_ = t_2__698_ | t_2__702_;
  assign t_3__697_ = t_2__697_ | t_2__701_;
  assign t_3__696_ = t_2__696_ | t_2__700_;
  assign t_3__695_ = t_2__695_ | t_2__699_;
  assign t_3__694_ = t_2__694_ | t_2__698_;
  assign t_3__693_ = t_2__693_ | t_2__697_;
  assign t_3__692_ = t_2__692_ | t_2__696_;
  assign t_3__691_ = t_2__691_ | t_2__695_;
  assign t_3__690_ = t_2__690_ | t_2__694_;
  assign t_3__689_ = t_2__689_ | t_2__693_;
  assign t_3__688_ = t_2__688_ | t_2__692_;
  assign t_3__687_ = t_2__687_ | t_2__691_;
  assign t_3__686_ = t_2__686_ | t_2__690_;
  assign t_3__685_ = t_2__685_ | t_2__689_;
  assign t_3__684_ = t_2__684_ | t_2__688_;
  assign t_3__683_ = t_2__683_ | t_2__687_;
  assign t_3__682_ = t_2__682_ | t_2__686_;
  assign t_3__681_ = t_2__681_ | t_2__685_;
  assign t_3__680_ = t_2__680_ | t_2__684_;
  assign t_3__679_ = t_2__679_ | t_2__683_;
  assign t_3__678_ = t_2__678_ | t_2__682_;
  assign t_3__677_ = t_2__677_ | t_2__681_;
  assign t_3__676_ = t_2__676_ | t_2__680_;
  assign t_3__675_ = t_2__675_ | t_2__679_;
  assign t_3__674_ = t_2__674_ | t_2__678_;
  assign t_3__673_ = t_2__673_ | t_2__677_;
  assign t_3__672_ = t_2__672_ | t_2__676_;
  assign t_3__671_ = t_2__671_ | t_2__675_;
  assign t_3__670_ = t_2__670_ | t_2__674_;
  assign t_3__669_ = t_2__669_ | t_2__673_;
  assign t_3__668_ = t_2__668_ | t_2__672_;
  assign t_3__667_ = t_2__667_ | t_2__671_;
  assign t_3__666_ = t_2__666_ | t_2__670_;
  assign t_3__665_ = t_2__665_ | t_2__669_;
  assign t_3__664_ = t_2__664_ | t_2__668_;
  assign t_3__663_ = t_2__663_ | t_2__667_;
  assign t_3__662_ = t_2__662_ | t_2__666_;
  assign t_3__661_ = t_2__661_ | t_2__665_;
  assign t_3__660_ = t_2__660_ | t_2__664_;
  assign t_3__659_ = t_2__659_ | t_2__663_;
  assign t_3__658_ = t_2__658_ | t_2__662_;
  assign t_3__657_ = t_2__657_ | t_2__661_;
  assign t_3__656_ = t_2__656_ | t_2__660_;
  assign t_3__655_ = t_2__655_ | t_2__659_;
  assign t_3__654_ = t_2__654_ | t_2__658_;
  assign t_3__653_ = t_2__653_ | t_2__657_;
  assign t_3__652_ = t_2__652_ | t_2__656_;
  assign t_3__651_ = t_2__651_ | t_2__655_;
  assign t_3__650_ = t_2__650_ | t_2__654_;
  assign t_3__649_ = t_2__649_ | t_2__653_;
  assign t_3__648_ = t_2__648_ | t_2__652_;
  assign t_3__647_ = t_2__647_ | t_2__651_;
  assign t_3__646_ = t_2__646_ | t_2__650_;
  assign t_3__645_ = t_2__645_ | t_2__649_;
  assign t_3__644_ = t_2__644_ | t_2__648_;
  assign t_3__643_ = t_2__643_ | t_2__647_;
  assign t_3__642_ = t_2__642_ | t_2__646_;
  assign t_3__641_ = t_2__641_ | t_2__645_;
  assign t_3__640_ = t_2__640_ | t_2__644_;
  assign t_3__639_ = t_2__639_ | t_2__643_;
  assign t_3__638_ = t_2__638_ | t_2__642_;
  assign t_3__637_ = t_2__637_ | t_2__641_;
  assign t_3__636_ = t_2__636_ | t_2__640_;
  assign t_3__635_ = t_2__635_ | t_2__639_;
  assign t_3__634_ = t_2__634_ | t_2__638_;
  assign t_3__633_ = t_2__633_ | t_2__637_;
  assign t_3__632_ = t_2__632_ | t_2__636_;
  assign t_3__631_ = t_2__631_ | t_2__635_;
  assign t_3__630_ = t_2__630_ | t_2__634_;
  assign t_3__629_ = t_2__629_ | t_2__633_;
  assign t_3__628_ = t_2__628_ | t_2__632_;
  assign t_3__627_ = t_2__627_ | t_2__631_;
  assign t_3__626_ = t_2__626_ | t_2__630_;
  assign t_3__625_ = t_2__625_ | t_2__629_;
  assign t_3__624_ = t_2__624_ | t_2__628_;
  assign t_3__623_ = t_2__623_ | t_2__627_;
  assign t_3__622_ = t_2__622_ | t_2__626_;
  assign t_3__621_ = t_2__621_ | t_2__625_;
  assign t_3__620_ = t_2__620_ | t_2__624_;
  assign t_3__619_ = t_2__619_ | t_2__623_;
  assign t_3__618_ = t_2__618_ | t_2__622_;
  assign t_3__617_ = t_2__617_ | t_2__621_;
  assign t_3__616_ = t_2__616_ | t_2__620_;
  assign t_3__615_ = t_2__615_ | t_2__619_;
  assign t_3__614_ = t_2__614_ | t_2__618_;
  assign t_3__613_ = t_2__613_ | t_2__617_;
  assign t_3__612_ = t_2__612_ | t_2__616_;
  assign t_3__611_ = t_2__611_ | t_2__615_;
  assign t_3__610_ = t_2__610_ | t_2__614_;
  assign t_3__609_ = t_2__609_ | t_2__613_;
  assign t_3__608_ = t_2__608_ | t_2__612_;
  assign t_3__607_ = t_2__607_ | t_2__611_;
  assign t_3__606_ = t_2__606_ | t_2__610_;
  assign t_3__605_ = t_2__605_ | t_2__609_;
  assign t_3__604_ = t_2__604_ | t_2__608_;
  assign t_3__603_ = t_2__603_ | t_2__607_;
  assign t_3__602_ = t_2__602_ | t_2__606_;
  assign t_3__601_ = t_2__601_ | t_2__605_;
  assign t_3__600_ = t_2__600_ | t_2__604_;
  assign t_3__599_ = t_2__599_ | t_2__603_;
  assign t_3__598_ = t_2__598_ | t_2__602_;
  assign t_3__597_ = t_2__597_ | t_2__601_;
  assign t_3__596_ = t_2__596_ | t_2__600_;
  assign t_3__595_ = t_2__595_ | t_2__599_;
  assign t_3__594_ = t_2__594_ | t_2__598_;
  assign t_3__593_ = t_2__593_ | t_2__597_;
  assign t_3__592_ = t_2__592_ | t_2__596_;
  assign t_3__591_ = t_2__591_ | t_2__595_;
  assign t_3__590_ = t_2__590_ | t_2__594_;
  assign t_3__589_ = t_2__589_ | t_2__593_;
  assign t_3__588_ = t_2__588_ | t_2__592_;
  assign t_3__587_ = t_2__587_ | t_2__591_;
  assign t_3__586_ = t_2__586_ | t_2__590_;
  assign t_3__585_ = t_2__585_ | t_2__589_;
  assign t_3__584_ = t_2__584_ | t_2__588_;
  assign t_3__583_ = t_2__583_ | t_2__587_;
  assign t_3__582_ = t_2__582_ | t_2__586_;
  assign t_3__581_ = t_2__581_ | t_2__585_;
  assign t_3__580_ = t_2__580_ | t_2__584_;
  assign t_3__579_ = t_2__579_ | t_2__583_;
  assign t_3__578_ = t_2__578_ | t_2__582_;
  assign t_3__577_ = t_2__577_ | t_2__581_;
  assign t_3__576_ = t_2__576_ | t_2__580_;
  assign t_3__575_ = t_2__575_ | t_2__579_;
  assign t_3__574_ = t_2__574_ | t_2__578_;
  assign t_3__573_ = t_2__573_ | t_2__577_;
  assign t_3__572_ = t_2__572_ | t_2__576_;
  assign t_3__571_ = t_2__571_ | t_2__575_;
  assign t_3__570_ = t_2__570_ | t_2__574_;
  assign t_3__569_ = t_2__569_ | t_2__573_;
  assign t_3__568_ = t_2__568_ | t_2__572_;
  assign t_3__567_ = t_2__567_ | t_2__571_;
  assign t_3__566_ = t_2__566_ | t_2__570_;
  assign t_3__565_ = t_2__565_ | t_2__569_;
  assign t_3__564_ = t_2__564_ | t_2__568_;
  assign t_3__563_ = t_2__563_ | t_2__567_;
  assign t_3__562_ = t_2__562_ | t_2__566_;
  assign t_3__561_ = t_2__561_ | t_2__565_;
  assign t_3__560_ = t_2__560_ | t_2__564_;
  assign t_3__559_ = t_2__559_ | t_2__563_;
  assign t_3__558_ = t_2__558_ | t_2__562_;
  assign t_3__557_ = t_2__557_ | t_2__561_;
  assign t_3__556_ = t_2__556_ | t_2__560_;
  assign t_3__555_ = t_2__555_ | t_2__559_;
  assign t_3__554_ = t_2__554_ | t_2__558_;
  assign t_3__553_ = t_2__553_ | t_2__557_;
  assign t_3__552_ = t_2__552_ | t_2__556_;
  assign t_3__551_ = t_2__551_ | t_2__555_;
  assign t_3__550_ = t_2__550_ | t_2__554_;
  assign t_3__549_ = t_2__549_ | t_2__553_;
  assign t_3__548_ = t_2__548_ | t_2__552_;
  assign t_3__547_ = t_2__547_ | t_2__551_;
  assign t_3__546_ = t_2__546_ | t_2__550_;
  assign t_3__545_ = t_2__545_ | t_2__549_;
  assign t_3__544_ = t_2__544_ | t_2__548_;
  assign t_3__543_ = t_2__543_ | t_2__547_;
  assign t_3__542_ = t_2__542_ | t_2__546_;
  assign t_3__541_ = t_2__541_ | t_2__545_;
  assign t_3__540_ = t_2__540_ | t_2__544_;
  assign t_3__539_ = t_2__539_ | t_2__543_;
  assign t_3__538_ = t_2__538_ | t_2__542_;
  assign t_3__537_ = t_2__537_ | t_2__541_;
  assign t_3__536_ = t_2__536_ | t_2__540_;
  assign t_3__535_ = t_2__535_ | t_2__539_;
  assign t_3__534_ = t_2__534_ | t_2__538_;
  assign t_3__533_ = t_2__533_ | t_2__537_;
  assign t_3__532_ = t_2__532_ | t_2__536_;
  assign t_3__531_ = t_2__531_ | t_2__535_;
  assign t_3__530_ = t_2__530_ | t_2__534_;
  assign t_3__529_ = t_2__529_ | t_2__533_;
  assign t_3__528_ = t_2__528_ | t_2__532_;
  assign t_3__527_ = t_2__527_ | t_2__531_;
  assign t_3__526_ = t_2__526_ | t_2__530_;
  assign t_3__525_ = t_2__525_ | t_2__529_;
  assign t_3__524_ = t_2__524_ | t_2__528_;
  assign t_3__523_ = t_2__523_ | t_2__527_;
  assign t_3__522_ = t_2__522_ | t_2__526_;
  assign t_3__521_ = t_2__521_ | t_2__525_;
  assign t_3__520_ = t_2__520_ | t_2__524_;
  assign t_3__519_ = t_2__519_ | t_2__523_;
  assign t_3__518_ = t_2__518_ | t_2__522_;
  assign t_3__517_ = t_2__517_ | t_2__521_;
  assign t_3__516_ = t_2__516_ | t_2__520_;
  assign t_3__515_ = t_2__515_ | t_2__519_;
  assign t_3__514_ = t_2__514_ | t_2__518_;
  assign t_3__513_ = t_2__513_ | t_2__517_;
  assign t_3__512_ = t_2__512_ | t_2__516_;
  assign t_3__511_ = t_2__511_ | t_2__515_;
  assign t_3__510_ = t_2__510_ | t_2__514_;
  assign t_3__509_ = t_2__509_ | t_2__513_;
  assign t_3__508_ = t_2__508_ | t_2__512_;
  assign t_3__507_ = t_2__507_ | t_2__511_;
  assign t_3__506_ = t_2__506_ | t_2__510_;
  assign t_3__505_ = t_2__505_ | t_2__509_;
  assign t_3__504_ = t_2__504_ | t_2__508_;
  assign t_3__503_ = t_2__503_ | t_2__507_;
  assign t_3__502_ = t_2__502_ | t_2__506_;
  assign t_3__501_ = t_2__501_ | t_2__505_;
  assign t_3__500_ = t_2__500_ | t_2__504_;
  assign t_3__499_ = t_2__499_ | t_2__503_;
  assign t_3__498_ = t_2__498_ | t_2__502_;
  assign t_3__497_ = t_2__497_ | t_2__501_;
  assign t_3__496_ = t_2__496_ | t_2__500_;
  assign t_3__495_ = t_2__495_ | t_2__499_;
  assign t_3__494_ = t_2__494_ | t_2__498_;
  assign t_3__493_ = t_2__493_ | t_2__497_;
  assign t_3__492_ = t_2__492_ | t_2__496_;
  assign t_3__491_ = t_2__491_ | t_2__495_;
  assign t_3__490_ = t_2__490_ | t_2__494_;
  assign t_3__489_ = t_2__489_ | t_2__493_;
  assign t_3__488_ = t_2__488_ | t_2__492_;
  assign t_3__487_ = t_2__487_ | t_2__491_;
  assign t_3__486_ = t_2__486_ | t_2__490_;
  assign t_3__485_ = t_2__485_ | t_2__489_;
  assign t_3__484_ = t_2__484_ | t_2__488_;
  assign t_3__483_ = t_2__483_ | t_2__487_;
  assign t_3__482_ = t_2__482_ | t_2__486_;
  assign t_3__481_ = t_2__481_ | t_2__485_;
  assign t_3__480_ = t_2__480_ | t_2__484_;
  assign t_3__479_ = t_2__479_ | t_2__483_;
  assign t_3__478_ = t_2__478_ | t_2__482_;
  assign t_3__477_ = t_2__477_ | t_2__481_;
  assign t_3__476_ = t_2__476_ | t_2__480_;
  assign t_3__475_ = t_2__475_ | t_2__479_;
  assign t_3__474_ = t_2__474_ | t_2__478_;
  assign t_3__473_ = t_2__473_ | t_2__477_;
  assign t_3__472_ = t_2__472_ | t_2__476_;
  assign t_3__471_ = t_2__471_ | t_2__475_;
  assign t_3__470_ = t_2__470_ | t_2__474_;
  assign t_3__469_ = t_2__469_ | t_2__473_;
  assign t_3__468_ = t_2__468_ | t_2__472_;
  assign t_3__467_ = t_2__467_ | t_2__471_;
  assign t_3__466_ = t_2__466_ | t_2__470_;
  assign t_3__465_ = t_2__465_ | t_2__469_;
  assign t_3__464_ = t_2__464_ | t_2__468_;
  assign t_3__463_ = t_2__463_ | t_2__467_;
  assign t_3__462_ = t_2__462_ | t_2__466_;
  assign t_3__461_ = t_2__461_ | t_2__465_;
  assign t_3__460_ = t_2__460_ | t_2__464_;
  assign t_3__459_ = t_2__459_ | t_2__463_;
  assign t_3__458_ = t_2__458_ | t_2__462_;
  assign t_3__457_ = t_2__457_ | t_2__461_;
  assign t_3__456_ = t_2__456_ | t_2__460_;
  assign t_3__455_ = t_2__455_ | t_2__459_;
  assign t_3__454_ = t_2__454_ | t_2__458_;
  assign t_3__453_ = t_2__453_ | t_2__457_;
  assign t_3__452_ = t_2__452_ | t_2__456_;
  assign t_3__451_ = t_2__451_ | t_2__455_;
  assign t_3__450_ = t_2__450_ | t_2__454_;
  assign t_3__449_ = t_2__449_ | t_2__453_;
  assign t_3__448_ = t_2__448_ | t_2__452_;
  assign t_3__447_ = t_2__447_ | t_2__451_;
  assign t_3__446_ = t_2__446_ | t_2__450_;
  assign t_3__445_ = t_2__445_ | t_2__449_;
  assign t_3__444_ = t_2__444_ | t_2__448_;
  assign t_3__443_ = t_2__443_ | t_2__447_;
  assign t_3__442_ = t_2__442_ | t_2__446_;
  assign t_3__441_ = t_2__441_ | t_2__445_;
  assign t_3__440_ = t_2__440_ | t_2__444_;
  assign t_3__439_ = t_2__439_ | t_2__443_;
  assign t_3__438_ = t_2__438_ | t_2__442_;
  assign t_3__437_ = t_2__437_ | t_2__441_;
  assign t_3__436_ = t_2__436_ | t_2__440_;
  assign t_3__435_ = t_2__435_ | t_2__439_;
  assign t_3__434_ = t_2__434_ | t_2__438_;
  assign t_3__433_ = t_2__433_ | t_2__437_;
  assign t_3__432_ = t_2__432_ | t_2__436_;
  assign t_3__431_ = t_2__431_ | t_2__435_;
  assign t_3__430_ = t_2__430_ | t_2__434_;
  assign t_3__429_ = t_2__429_ | t_2__433_;
  assign t_3__428_ = t_2__428_ | t_2__432_;
  assign t_3__427_ = t_2__427_ | t_2__431_;
  assign t_3__426_ = t_2__426_ | t_2__430_;
  assign t_3__425_ = t_2__425_ | t_2__429_;
  assign t_3__424_ = t_2__424_ | t_2__428_;
  assign t_3__423_ = t_2__423_ | t_2__427_;
  assign t_3__422_ = t_2__422_ | t_2__426_;
  assign t_3__421_ = t_2__421_ | t_2__425_;
  assign t_3__420_ = t_2__420_ | t_2__424_;
  assign t_3__419_ = t_2__419_ | t_2__423_;
  assign t_3__418_ = t_2__418_ | t_2__422_;
  assign t_3__417_ = t_2__417_ | t_2__421_;
  assign t_3__416_ = t_2__416_ | t_2__420_;
  assign t_3__415_ = t_2__415_ | t_2__419_;
  assign t_3__414_ = t_2__414_ | t_2__418_;
  assign t_3__413_ = t_2__413_ | t_2__417_;
  assign t_3__412_ = t_2__412_ | t_2__416_;
  assign t_3__411_ = t_2__411_ | t_2__415_;
  assign t_3__410_ = t_2__410_ | t_2__414_;
  assign t_3__409_ = t_2__409_ | t_2__413_;
  assign t_3__408_ = t_2__408_ | t_2__412_;
  assign t_3__407_ = t_2__407_ | t_2__411_;
  assign t_3__406_ = t_2__406_ | t_2__410_;
  assign t_3__405_ = t_2__405_ | t_2__409_;
  assign t_3__404_ = t_2__404_ | t_2__408_;
  assign t_3__403_ = t_2__403_ | t_2__407_;
  assign t_3__402_ = t_2__402_ | t_2__406_;
  assign t_3__401_ = t_2__401_ | t_2__405_;
  assign t_3__400_ = t_2__400_ | t_2__404_;
  assign t_3__399_ = t_2__399_ | t_2__403_;
  assign t_3__398_ = t_2__398_ | t_2__402_;
  assign t_3__397_ = t_2__397_ | t_2__401_;
  assign t_3__396_ = t_2__396_ | t_2__400_;
  assign t_3__395_ = t_2__395_ | t_2__399_;
  assign t_3__394_ = t_2__394_ | t_2__398_;
  assign t_3__393_ = t_2__393_ | t_2__397_;
  assign t_3__392_ = t_2__392_ | t_2__396_;
  assign t_3__391_ = t_2__391_ | t_2__395_;
  assign t_3__390_ = t_2__390_ | t_2__394_;
  assign t_3__389_ = t_2__389_ | t_2__393_;
  assign t_3__388_ = t_2__388_ | t_2__392_;
  assign t_3__387_ = t_2__387_ | t_2__391_;
  assign t_3__386_ = t_2__386_ | t_2__390_;
  assign t_3__385_ = t_2__385_ | t_2__389_;
  assign t_3__384_ = t_2__384_ | t_2__388_;
  assign t_3__383_ = t_2__383_ | t_2__387_;
  assign t_3__382_ = t_2__382_ | t_2__386_;
  assign t_3__381_ = t_2__381_ | t_2__385_;
  assign t_3__380_ = t_2__380_ | t_2__384_;
  assign t_3__379_ = t_2__379_ | t_2__383_;
  assign t_3__378_ = t_2__378_ | t_2__382_;
  assign t_3__377_ = t_2__377_ | t_2__381_;
  assign t_3__376_ = t_2__376_ | t_2__380_;
  assign t_3__375_ = t_2__375_ | t_2__379_;
  assign t_3__374_ = t_2__374_ | t_2__378_;
  assign t_3__373_ = t_2__373_ | t_2__377_;
  assign t_3__372_ = t_2__372_ | t_2__376_;
  assign t_3__371_ = t_2__371_ | t_2__375_;
  assign t_3__370_ = t_2__370_ | t_2__374_;
  assign t_3__369_ = t_2__369_ | t_2__373_;
  assign t_3__368_ = t_2__368_ | t_2__372_;
  assign t_3__367_ = t_2__367_ | t_2__371_;
  assign t_3__366_ = t_2__366_ | t_2__370_;
  assign t_3__365_ = t_2__365_ | t_2__369_;
  assign t_3__364_ = t_2__364_ | t_2__368_;
  assign t_3__363_ = t_2__363_ | t_2__367_;
  assign t_3__362_ = t_2__362_ | t_2__366_;
  assign t_3__361_ = t_2__361_ | t_2__365_;
  assign t_3__360_ = t_2__360_ | t_2__364_;
  assign t_3__359_ = t_2__359_ | t_2__363_;
  assign t_3__358_ = t_2__358_ | t_2__362_;
  assign t_3__357_ = t_2__357_ | t_2__361_;
  assign t_3__356_ = t_2__356_ | t_2__360_;
  assign t_3__355_ = t_2__355_ | t_2__359_;
  assign t_3__354_ = t_2__354_ | t_2__358_;
  assign t_3__353_ = t_2__353_ | t_2__357_;
  assign t_3__352_ = t_2__352_ | t_2__356_;
  assign t_3__351_ = t_2__351_ | t_2__355_;
  assign t_3__350_ = t_2__350_ | t_2__354_;
  assign t_3__349_ = t_2__349_ | t_2__353_;
  assign t_3__348_ = t_2__348_ | t_2__352_;
  assign t_3__347_ = t_2__347_ | t_2__351_;
  assign t_3__346_ = t_2__346_ | t_2__350_;
  assign t_3__345_ = t_2__345_ | t_2__349_;
  assign t_3__344_ = t_2__344_ | t_2__348_;
  assign t_3__343_ = t_2__343_ | t_2__347_;
  assign t_3__342_ = t_2__342_ | t_2__346_;
  assign t_3__341_ = t_2__341_ | t_2__345_;
  assign t_3__340_ = t_2__340_ | t_2__344_;
  assign t_3__339_ = t_2__339_ | t_2__343_;
  assign t_3__338_ = t_2__338_ | t_2__342_;
  assign t_3__337_ = t_2__337_ | t_2__341_;
  assign t_3__336_ = t_2__336_ | t_2__340_;
  assign t_3__335_ = t_2__335_ | t_2__339_;
  assign t_3__334_ = t_2__334_ | t_2__338_;
  assign t_3__333_ = t_2__333_ | t_2__337_;
  assign t_3__332_ = t_2__332_ | t_2__336_;
  assign t_3__331_ = t_2__331_ | t_2__335_;
  assign t_3__330_ = t_2__330_ | t_2__334_;
  assign t_3__329_ = t_2__329_ | t_2__333_;
  assign t_3__328_ = t_2__328_ | t_2__332_;
  assign t_3__327_ = t_2__327_ | t_2__331_;
  assign t_3__326_ = t_2__326_ | t_2__330_;
  assign t_3__325_ = t_2__325_ | t_2__329_;
  assign t_3__324_ = t_2__324_ | t_2__328_;
  assign t_3__323_ = t_2__323_ | t_2__327_;
  assign t_3__322_ = t_2__322_ | t_2__326_;
  assign t_3__321_ = t_2__321_ | t_2__325_;
  assign t_3__320_ = t_2__320_ | t_2__324_;
  assign t_3__319_ = t_2__319_ | t_2__323_;
  assign t_3__318_ = t_2__318_ | t_2__322_;
  assign t_3__317_ = t_2__317_ | t_2__321_;
  assign t_3__316_ = t_2__316_ | t_2__320_;
  assign t_3__315_ = t_2__315_ | t_2__319_;
  assign t_3__314_ = t_2__314_ | t_2__318_;
  assign t_3__313_ = t_2__313_ | t_2__317_;
  assign t_3__312_ = t_2__312_ | t_2__316_;
  assign t_3__311_ = t_2__311_ | t_2__315_;
  assign t_3__310_ = t_2__310_ | t_2__314_;
  assign t_3__309_ = t_2__309_ | t_2__313_;
  assign t_3__308_ = t_2__308_ | t_2__312_;
  assign t_3__307_ = t_2__307_ | t_2__311_;
  assign t_3__306_ = t_2__306_ | t_2__310_;
  assign t_3__305_ = t_2__305_ | t_2__309_;
  assign t_3__304_ = t_2__304_ | t_2__308_;
  assign t_3__303_ = t_2__303_ | t_2__307_;
  assign t_3__302_ = t_2__302_ | t_2__306_;
  assign t_3__301_ = t_2__301_ | t_2__305_;
  assign t_3__300_ = t_2__300_ | t_2__304_;
  assign t_3__299_ = t_2__299_ | t_2__303_;
  assign t_3__298_ = t_2__298_ | t_2__302_;
  assign t_3__297_ = t_2__297_ | t_2__301_;
  assign t_3__296_ = t_2__296_ | t_2__300_;
  assign t_3__295_ = t_2__295_ | t_2__299_;
  assign t_3__294_ = t_2__294_ | t_2__298_;
  assign t_3__293_ = t_2__293_ | t_2__297_;
  assign t_3__292_ = t_2__292_ | t_2__296_;
  assign t_3__291_ = t_2__291_ | t_2__295_;
  assign t_3__290_ = t_2__290_ | t_2__294_;
  assign t_3__289_ = t_2__289_ | t_2__293_;
  assign t_3__288_ = t_2__288_ | t_2__292_;
  assign t_3__287_ = t_2__287_ | t_2__291_;
  assign t_3__286_ = t_2__286_ | t_2__290_;
  assign t_3__285_ = t_2__285_ | t_2__289_;
  assign t_3__284_ = t_2__284_ | t_2__288_;
  assign t_3__283_ = t_2__283_ | t_2__287_;
  assign t_3__282_ = t_2__282_ | t_2__286_;
  assign t_3__281_ = t_2__281_ | t_2__285_;
  assign t_3__280_ = t_2__280_ | t_2__284_;
  assign t_3__279_ = t_2__279_ | t_2__283_;
  assign t_3__278_ = t_2__278_ | t_2__282_;
  assign t_3__277_ = t_2__277_ | t_2__281_;
  assign t_3__276_ = t_2__276_ | t_2__280_;
  assign t_3__275_ = t_2__275_ | t_2__279_;
  assign t_3__274_ = t_2__274_ | t_2__278_;
  assign t_3__273_ = t_2__273_ | t_2__277_;
  assign t_3__272_ = t_2__272_ | t_2__276_;
  assign t_3__271_ = t_2__271_ | t_2__275_;
  assign t_3__270_ = t_2__270_ | t_2__274_;
  assign t_3__269_ = t_2__269_ | t_2__273_;
  assign t_3__268_ = t_2__268_ | t_2__272_;
  assign t_3__267_ = t_2__267_ | t_2__271_;
  assign t_3__266_ = t_2__266_ | t_2__270_;
  assign t_3__265_ = t_2__265_ | t_2__269_;
  assign t_3__264_ = t_2__264_ | t_2__268_;
  assign t_3__263_ = t_2__263_ | t_2__267_;
  assign t_3__262_ = t_2__262_ | t_2__266_;
  assign t_3__261_ = t_2__261_ | t_2__265_;
  assign t_3__260_ = t_2__260_ | t_2__264_;
  assign t_3__259_ = t_2__259_ | t_2__263_;
  assign t_3__258_ = t_2__258_ | t_2__262_;
  assign t_3__257_ = t_2__257_ | t_2__261_;
  assign t_3__256_ = t_2__256_ | t_2__260_;
  assign t_3__255_ = t_2__255_ | t_2__259_;
  assign t_3__254_ = t_2__254_ | t_2__258_;
  assign t_3__253_ = t_2__253_ | t_2__257_;
  assign t_3__252_ = t_2__252_ | t_2__256_;
  assign t_3__251_ = t_2__251_ | t_2__255_;
  assign t_3__250_ = t_2__250_ | t_2__254_;
  assign t_3__249_ = t_2__249_ | t_2__253_;
  assign t_3__248_ = t_2__248_ | t_2__252_;
  assign t_3__247_ = t_2__247_ | t_2__251_;
  assign t_3__246_ = t_2__246_ | t_2__250_;
  assign t_3__245_ = t_2__245_ | t_2__249_;
  assign t_3__244_ = t_2__244_ | t_2__248_;
  assign t_3__243_ = t_2__243_ | t_2__247_;
  assign t_3__242_ = t_2__242_ | t_2__246_;
  assign t_3__241_ = t_2__241_ | t_2__245_;
  assign t_3__240_ = t_2__240_ | t_2__244_;
  assign t_3__239_ = t_2__239_ | t_2__243_;
  assign t_3__238_ = t_2__238_ | t_2__242_;
  assign t_3__237_ = t_2__237_ | t_2__241_;
  assign t_3__236_ = t_2__236_ | t_2__240_;
  assign t_3__235_ = t_2__235_ | t_2__239_;
  assign t_3__234_ = t_2__234_ | t_2__238_;
  assign t_3__233_ = t_2__233_ | t_2__237_;
  assign t_3__232_ = t_2__232_ | t_2__236_;
  assign t_3__231_ = t_2__231_ | t_2__235_;
  assign t_3__230_ = t_2__230_ | t_2__234_;
  assign t_3__229_ = t_2__229_ | t_2__233_;
  assign t_3__228_ = t_2__228_ | t_2__232_;
  assign t_3__227_ = t_2__227_ | t_2__231_;
  assign t_3__226_ = t_2__226_ | t_2__230_;
  assign t_3__225_ = t_2__225_ | t_2__229_;
  assign t_3__224_ = t_2__224_ | t_2__228_;
  assign t_3__223_ = t_2__223_ | t_2__227_;
  assign t_3__222_ = t_2__222_ | t_2__226_;
  assign t_3__221_ = t_2__221_ | t_2__225_;
  assign t_3__220_ = t_2__220_ | t_2__224_;
  assign t_3__219_ = t_2__219_ | t_2__223_;
  assign t_3__218_ = t_2__218_ | t_2__222_;
  assign t_3__217_ = t_2__217_ | t_2__221_;
  assign t_3__216_ = t_2__216_ | t_2__220_;
  assign t_3__215_ = t_2__215_ | t_2__219_;
  assign t_3__214_ = t_2__214_ | t_2__218_;
  assign t_3__213_ = t_2__213_ | t_2__217_;
  assign t_3__212_ = t_2__212_ | t_2__216_;
  assign t_3__211_ = t_2__211_ | t_2__215_;
  assign t_3__210_ = t_2__210_ | t_2__214_;
  assign t_3__209_ = t_2__209_ | t_2__213_;
  assign t_3__208_ = t_2__208_ | t_2__212_;
  assign t_3__207_ = t_2__207_ | t_2__211_;
  assign t_3__206_ = t_2__206_ | t_2__210_;
  assign t_3__205_ = t_2__205_ | t_2__209_;
  assign t_3__204_ = t_2__204_ | t_2__208_;
  assign t_3__203_ = t_2__203_ | t_2__207_;
  assign t_3__202_ = t_2__202_ | t_2__206_;
  assign t_3__201_ = t_2__201_ | t_2__205_;
  assign t_3__200_ = t_2__200_ | t_2__204_;
  assign t_3__199_ = t_2__199_ | t_2__203_;
  assign t_3__198_ = t_2__198_ | t_2__202_;
  assign t_3__197_ = t_2__197_ | t_2__201_;
  assign t_3__196_ = t_2__196_ | t_2__200_;
  assign t_3__195_ = t_2__195_ | t_2__199_;
  assign t_3__194_ = t_2__194_ | t_2__198_;
  assign t_3__193_ = t_2__193_ | t_2__197_;
  assign t_3__192_ = t_2__192_ | t_2__196_;
  assign t_3__191_ = t_2__191_ | t_2__195_;
  assign t_3__190_ = t_2__190_ | t_2__194_;
  assign t_3__189_ = t_2__189_ | t_2__193_;
  assign t_3__188_ = t_2__188_ | t_2__192_;
  assign t_3__187_ = t_2__187_ | t_2__191_;
  assign t_3__186_ = t_2__186_ | t_2__190_;
  assign t_3__185_ = t_2__185_ | t_2__189_;
  assign t_3__184_ = t_2__184_ | t_2__188_;
  assign t_3__183_ = t_2__183_ | t_2__187_;
  assign t_3__182_ = t_2__182_ | t_2__186_;
  assign t_3__181_ = t_2__181_ | t_2__185_;
  assign t_3__180_ = t_2__180_ | t_2__184_;
  assign t_3__179_ = t_2__179_ | t_2__183_;
  assign t_3__178_ = t_2__178_ | t_2__182_;
  assign t_3__177_ = t_2__177_ | t_2__181_;
  assign t_3__176_ = t_2__176_ | t_2__180_;
  assign t_3__175_ = t_2__175_ | t_2__179_;
  assign t_3__174_ = t_2__174_ | t_2__178_;
  assign t_3__173_ = t_2__173_ | t_2__177_;
  assign t_3__172_ = t_2__172_ | t_2__176_;
  assign t_3__171_ = t_2__171_ | t_2__175_;
  assign t_3__170_ = t_2__170_ | t_2__174_;
  assign t_3__169_ = t_2__169_ | t_2__173_;
  assign t_3__168_ = t_2__168_ | t_2__172_;
  assign t_3__167_ = t_2__167_ | t_2__171_;
  assign t_3__166_ = t_2__166_ | t_2__170_;
  assign t_3__165_ = t_2__165_ | t_2__169_;
  assign t_3__164_ = t_2__164_ | t_2__168_;
  assign t_3__163_ = t_2__163_ | t_2__167_;
  assign t_3__162_ = t_2__162_ | t_2__166_;
  assign t_3__161_ = t_2__161_ | t_2__165_;
  assign t_3__160_ = t_2__160_ | t_2__164_;
  assign t_3__159_ = t_2__159_ | t_2__163_;
  assign t_3__158_ = t_2__158_ | t_2__162_;
  assign t_3__157_ = t_2__157_ | t_2__161_;
  assign t_3__156_ = t_2__156_ | t_2__160_;
  assign t_3__155_ = t_2__155_ | t_2__159_;
  assign t_3__154_ = t_2__154_ | t_2__158_;
  assign t_3__153_ = t_2__153_ | t_2__157_;
  assign t_3__152_ = t_2__152_ | t_2__156_;
  assign t_3__151_ = t_2__151_ | t_2__155_;
  assign t_3__150_ = t_2__150_ | t_2__154_;
  assign t_3__149_ = t_2__149_ | t_2__153_;
  assign t_3__148_ = t_2__148_ | t_2__152_;
  assign t_3__147_ = t_2__147_ | t_2__151_;
  assign t_3__146_ = t_2__146_ | t_2__150_;
  assign t_3__145_ = t_2__145_ | t_2__149_;
  assign t_3__144_ = t_2__144_ | t_2__148_;
  assign t_3__143_ = t_2__143_ | t_2__147_;
  assign t_3__142_ = t_2__142_ | t_2__146_;
  assign t_3__141_ = t_2__141_ | t_2__145_;
  assign t_3__140_ = t_2__140_ | t_2__144_;
  assign t_3__139_ = t_2__139_ | t_2__143_;
  assign t_3__138_ = t_2__138_ | t_2__142_;
  assign t_3__137_ = t_2__137_ | t_2__141_;
  assign t_3__136_ = t_2__136_ | t_2__140_;
  assign t_3__135_ = t_2__135_ | t_2__139_;
  assign t_3__134_ = t_2__134_ | t_2__138_;
  assign t_3__133_ = t_2__133_ | t_2__137_;
  assign t_3__132_ = t_2__132_ | t_2__136_;
  assign t_3__131_ = t_2__131_ | t_2__135_;
  assign t_3__130_ = t_2__130_ | t_2__134_;
  assign t_3__129_ = t_2__129_ | t_2__133_;
  assign t_3__128_ = t_2__128_ | t_2__132_;
  assign t_3__127_ = t_2__127_ | t_2__131_;
  assign t_3__126_ = t_2__126_ | t_2__130_;
  assign t_3__125_ = t_2__125_ | t_2__129_;
  assign t_3__124_ = t_2__124_ | t_2__128_;
  assign t_3__123_ = t_2__123_ | t_2__127_;
  assign t_3__122_ = t_2__122_ | t_2__126_;
  assign t_3__121_ = t_2__121_ | t_2__125_;
  assign t_3__120_ = t_2__120_ | t_2__124_;
  assign t_3__119_ = t_2__119_ | t_2__123_;
  assign t_3__118_ = t_2__118_ | t_2__122_;
  assign t_3__117_ = t_2__117_ | t_2__121_;
  assign t_3__116_ = t_2__116_ | t_2__120_;
  assign t_3__115_ = t_2__115_ | t_2__119_;
  assign t_3__114_ = t_2__114_ | t_2__118_;
  assign t_3__113_ = t_2__113_ | t_2__117_;
  assign t_3__112_ = t_2__112_ | t_2__116_;
  assign t_3__111_ = t_2__111_ | t_2__115_;
  assign t_3__110_ = t_2__110_ | t_2__114_;
  assign t_3__109_ = t_2__109_ | t_2__113_;
  assign t_3__108_ = t_2__108_ | t_2__112_;
  assign t_3__107_ = t_2__107_ | t_2__111_;
  assign t_3__106_ = t_2__106_ | t_2__110_;
  assign t_3__105_ = t_2__105_ | t_2__109_;
  assign t_3__104_ = t_2__104_ | t_2__108_;
  assign t_3__103_ = t_2__103_ | t_2__107_;
  assign t_3__102_ = t_2__102_ | t_2__106_;
  assign t_3__101_ = t_2__101_ | t_2__105_;
  assign t_3__100_ = t_2__100_ | t_2__104_;
  assign t_3__99_ = t_2__99_ | t_2__103_;
  assign t_3__98_ = t_2__98_ | t_2__102_;
  assign t_3__97_ = t_2__97_ | t_2__101_;
  assign t_3__96_ = t_2__96_ | t_2__100_;
  assign t_3__95_ = t_2__95_ | t_2__99_;
  assign t_3__94_ = t_2__94_ | t_2__98_;
  assign t_3__93_ = t_2__93_ | t_2__97_;
  assign t_3__92_ = t_2__92_ | t_2__96_;
  assign t_3__91_ = t_2__91_ | t_2__95_;
  assign t_3__90_ = t_2__90_ | t_2__94_;
  assign t_3__89_ = t_2__89_ | t_2__93_;
  assign t_3__88_ = t_2__88_ | t_2__92_;
  assign t_3__87_ = t_2__87_ | t_2__91_;
  assign t_3__86_ = t_2__86_ | t_2__90_;
  assign t_3__85_ = t_2__85_ | t_2__89_;
  assign t_3__84_ = t_2__84_ | t_2__88_;
  assign t_3__83_ = t_2__83_ | t_2__87_;
  assign t_3__82_ = t_2__82_ | t_2__86_;
  assign t_3__81_ = t_2__81_ | t_2__85_;
  assign t_3__80_ = t_2__80_ | t_2__84_;
  assign t_3__79_ = t_2__79_ | t_2__83_;
  assign t_3__78_ = t_2__78_ | t_2__82_;
  assign t_3__77_ = t_2__77_ | t_2__81_;
  assign t_3__76_ = t_2__76_ | t_2__80_;
  assign t_3__75_ = t_2__75_ | t_2__79_;
  assign t_3__74_ = t_2__74_ | t_2__78_;
  assign t_3__73_ = t_2__73_ | t_2__77_;
  assign t_3__72_ = t_2__72_ | t_2__76_;
  assign t_3__71_ = t_2__71_ | t_2__75_;
  assign t_3__70_ = t_2__70_ | t_2__74_;
  assign t_3__69_ = t_2__69_ | t_2__73_;
  assign t_3__68_ = t_2__68_ | t_2__72_;
  assign t_3__67_ = t_2__67_ | t_2__71_;
  assign t_3__66_ = t_2__66_ | t_2__70_;
  assign t_3__65_ = t_2__65_ | t_2__69_;
  assign t_3__64_ = t_2__64_ | t_2__68_;
  assign t_3__63_ = t_2__63_ | t_2__67_;
  assign t_3__62_ = t_2__62_ | t_2__66_;
  assign t_3__61_ = t_2__61_ | t_2__65_;
  assign t_3__60_ = t_2__60_ | t_2__64_;
  assign t_3__59_ = t_2__59_ | t_2__63_;
  assign t_3__58_ = t_2__58_ | t_2__62_;
  assign t_3__57_ = t_2__57_ | t_2__61_;
  assign t_3__56_ = t_2__56_ | t_2__60_;
  assign t_3__55_ = t_2__55_ | t_2__59_;
  assign t_3__54_ = t_2__54_ | t_2__58_;
  assign t_3__53_ = t_2__53_ | t_2__57_;
  assign t_3__52_ = t_2__52_ | t_2__56_;
  assign t_3__51_ = t_2__51_ | t_2__55_;
  assign t_3__50_ = t_2__50_ | t_2__54_;
  assign t_3__49_ = t_2__49_ | t_2__53_;
  assign t_3__48_ = t_2__48_ | t_2__52_;
  assign t_3__47_ = t_2__47_ | t_2__51_;
  assign t_3__46_ = t_2__46_ | t_2__50_;
  assign t_3__45_ = t_2__45_ | t_2__49_;
  assign t_3__44_ = t_2__44_ | t_2__48_;
  assign t_3__43_ = t_2__43_ | t_2__47_;
  assign t_3__42_ = t_2__42_ | t_2__46_;
  assign t_3__41_ = t_2__41_ | t_2__45_;
  assign t_3__40_ = t_2__40_ | t_2__44_;
  assign t_3__39_ = t_2__39_ | t_2__43_;
  assign t_3__38_ = t_2__38_ | t_2__42_;
  assign t_3__37_ = t_2__37_ | t_2__41_;
  assign t_3__36_ = t_2__36_ | t_2__40_;
  assign t_3__35_ = t_2__35_ | t_2__39_;
  assign t_3__34_ = t_2__34_ | t_2__38_;
  assign t_3__33_ = t_2__33_ | t_2__37_;
  assign t_3__32_ = t_2__32_ | t_2__36_;
  assign t_3__31_ = t_2__31_ | t_2__35_;
  assign t_3__30_ = t_2__30_ | t_2__34_;
  assign t_3__29_ = t_2__29_ | t_2__33_;
  assign t_3__28_ = t_2__28_ | t_2__32_;
  assign t_3__27_ = t_2__27_ | t_2__31_;
  assign t_3__26_ = t_2__26_ | t_2__30_;
  assign t_3__25_ = t_2__25_ | t_2__29_;
  assign t_3__24_ = t_2__24_ | t_2__28_;
  assign t_3__23_ = t_2__23_ | t_2__27_;
  assign t_3__22_ = t_2__22_ | t_2__26_;
  assign t_3__21_ = t_2__21_ | t_2__25_;
  assign t_3__20_ = t_2__20_ | t_2__24_;
  assign t_3__19_ = t_2__19_ | t_2__23_;
  assign t_3__18_ = t_2__18_ | t_2__22_;
  assign t_3__17_ = t_2__17_ | t_2__21_;
  assign t_3__16_ = t_2__16_ | t_2__20_;
  assign t_3__15_ = t_2__15_ | t_2__19_;
  assign t_3__14_ = t_2__14_ | t_2__18_;
  assign t_3__13_ = t_2__13_ | t_2__17_;
  assign t_3__12_ = t_2__12_ | t_2__16_;
  assign t_3__11_ = t_2__11_ | t_2__15_;
  assign t_3__10_ = t_2__10_ | t_2__14_;
  assign t_3__9_ = t_2__9_ | t_2__13_;
  assign t_3__8_ = t_2__8_ | t_2__12_;
  assign t_3__7_ = t_2__7_ | t_2__11_;
  assign t_3__6_ = t_2__6_ | t_2__10_;
  assign t_3__5_ = t_2__5_ | t_2__9_;
  assign t_3__4_ = t_2__4_ | t_2__8_;
  assign t_3__3_ = t_2__3_ | t_2__7_;
  assign t_3__2_ = t_2__2_ | t_2__6_;
  assign t_3__1_ = t_2__1_ | t_2__5_;
  assign t_3__0_ = t_2__0_ | t_2__4_;
  assign t_4__1023_ = t_3__1023_ | 1'b0;
  assign t_4__1022_ = t_3__1022_ | 1'b0;
  assign t_4__1021_ = t_3__1021_ | 1'b0;
  assign t_4__1020_ = t_3__1020_ | 1'b0;
  assign t_4__1019_ = t_3__1019_ | 1'b0;
  assign t_4__1018_ = t_3__1018_ | 1'b0;
  assign t_4__1017_ = t_3__1017_ | 1'b0;
  assign t_4__1016_ = t_3__1016_ | 1'b0;
  assign t_4__1015_ = t_3__1015_ | t_3__1023_;
  assign t_4__1014_ = t_3__1014_ | t_3__1022_;
  assign t_4__1013_ = t_3__1013_ | t_3__1021_;
  assign t_4__1012_ = t_3__1012_ | t_3__1020_;
  assign t_4__1011_ = t_3__1011_ | t_3__1019_;
  assign t_4__1010_ = t_3__1010_ | t_3__1018_;
  assign t_4__1009_ = t_3__1009_ | t_3__1017_;
  assign t_4__1008_ = t_3__1008_ | t_3__1016_;
  assign t_4__1007_ = t_3__1007_ | t_3__1015_;
  assign t_4__1006_ = t_3__1006_ | t_3__1014_;
  assign t_4__1005_ = t_3__1005_ | t_3__1013_;
  assign t_4__1004_ = t_3__1004_ | t_3__1012_;
  assign t_4__1003_ = t_3__1003_ | t_3__1011_;
  assign t_4__1002_ = t_3__1002_ | t_3__1010_;
  assign t_4__1001_ = t_3__1001_ | t_3__1009_;
  assign t_4__1000_ = t_3__1000_ | t_3__1008_;
  assign t_4__999_ = t_3__999_ | t_3__1007_;
  assign t_4__998_ = t_3__998_ | t_3__1006_;
  assign t_4__997_ = t_3__997_ | t_3__1005_;
  assign t_4__996_ = t_3__996_ | t_3__1004_;
  assign t_4__995_ = t_3__995_ | t_3__1003_;
  assign t_4__994_ = t_3__994_ | t_3__1002_;
  assign t_4__993_ = t_3__993_ | t_3__1001_;
  assign t_4__992_ = t_3__992_ | t_3__1000_;
  assign t_4__991_ = t_3__991_ | t_3__999_;
  assign t_4__990_ = t_3__990_ | t_3__998_;
  assign t_4__989_ = t_3__989_ | t_3__997_;
  assign t_4__988_ = t_3__988_ | t_3__996_;
  assign t_4__987_ = t_3__987_ | t_3__995_;
  assign t_4__986_ = t_3__986_ | t_3__994_;
  assign t_4__985_ = t_3__985_ | t_3__993_;
  assign t_4__984_ = t_3__984_ | t_3__992_;
  assign t_4__983_ = t_3__983_ | t_3__991_;
  assign t_4__982_ = t_3__982_ | t_3__990_;
  assign t_4__981_ = t_3__981_ | t_3__989_;
  assign t_4__980_ = t_3__980_ | t_3__988_;
  assign t_4__979_ = t_3__979_ | t_3__987_;
  assign t_4__978_ = t_3__978_ | t_3__986_;
  assign t_4__977_ = t_3__977_ | t_3__985_;
  assign t_4__976_ = t_3__976_ | t_3__984_;
  assign t_4__975_ = t_3__975_ | t_3__983_;
  assign t_4__974_ = t_3__974_ | t_3__982_;
  assign t_4__973_ = t_3__973_ | t_3__981_;
  assign t_4__972_ = t_3__972_ | t_3__980_;
  assign t_4__971_ = t_3__971_ | t_3__979_;
  assign t_4__970_ = t_3__970_ | t_3__978_;
  assign t_4__969_ = t_3__969_ | t_3__977_;
  assign t_4__968_ = t_3__968_ | t_3__976_;
  assign t_4__967_ = t_3__967_ | t_3__975_;
  assign t_4__966_ = t_3__966_ | t_3__974_;
  assign t_4__965_ = t_3__965_ | t_3__973_;
  assign t_4__964_ = t_3__964_ | t_3__972_;
  assign t_4__963_ = t_3__963_ | t_3__971_;
  assign t_4__962_ = t_3__962_ | t_3__970_;
  assign t_4__961_ = t_3__961_ | t_3__969_;
  assign t_4__960_ = t_3__960_ | t_3__968_;
  assign t_4__959_ = t_3__959_ | t_3__967_;
  assign t_4__958_ = t_3__958_ | t_3__966_;
  assign t_4__957_ = t_3__957_ | t_3__965_;
  assign t_4__956_ = t_3__956_ | t_3__964_;
  assign t_4__955_ = t_3__955_ | t_3__963_;
  assign t_4__954_ = t_3__954_ | t_3__962_;
  assign t_4__953_ = t_3__953_ | t_3__961_;
  assign t_4__952_ = t_3__952_ | t_3__960_;
  assign t_4__951_ = t_3__951_ | t_3__959_;
  assign t_4__950_ = t_3__950_ | t_3__958_;
  assign t_4__949_ = t_3__949_ | t_3__957_;
  assign t_4__948_ = t_3__948_ | t_3__956_;
  assign t_4__947_ = t_3__947_ | t_3__955_;
  assign t_4__946_ = t_3__946_ | t_3__954_;
  assign t_4__945_ = t_3__945_ | t_3__953_;
  assign t_4__944_ = t_3__944_ | t_3__952_;
  assign t_4__943_ = t_3__943_ | t_3__951_;
  assign t_4__942_ = t_3__942_ | t_3__950_;
  assign t_4__941_ = t_3__941_ | t_3__949_;
  assign t_4__940_ = t_3__940_ | t_3__948_;
  assign t_4__939_ = t_3__939_ | t_3__947_;
  assign t_4__938_ = t_3__938_ | t_3__946_;
  assign t_4__937_ = t_3__937_ | t_3__945_;
  assign t_4__936_ = t_3__936_ | t_3__944_;
  assign t_4__935_ = t_3__935_ | t_3__943_;
  assign t_4__934_ = t_3__934_ | t_3__942_;
  assign t_4__933_ = t_3__933_ | t_3__941_;
  assign t_4__932_ = t_3__932_ | t_3__940_;
  assign t_4__931_ = t_3__931_ | t_3__939_;
  assign t_4__930_ = t_3__930_ | t_3__938_;
  assign t_4__929_ = t_3__929_ | t_3__937_;
  assign t_4__928_ = t_3__928_ | t_3__936_;
  assign t_4__927_ = t_3__927_ | t_3__935_;
  assign t_4__926_ = t_3__926_ | t_3__934_;
  assign t_4__925_ = t_3__925_ | t_3__933_;
  assign t_4__924_ = t_3__924_ | t_3__932_;
  assign t_4__923_ = t_3__923_ | t_3__931_;
  assign t_4__922_ = t_3__922_ | t_3__930_;
  assign t_4__921_ = t_3__921_ | t_3__929_;
  assign t_4__920_ = t_3__920_ | t_3__928_;
  assign t_4__919_ = t_3__919_ | t_3__927_;
  assign t_4__918_ = t_3__918_ | t_3__926_;
  assign t_4__917_ = t_3__917_ | t_3__925_;
  assign t_4__916_ = t_3__916_ | t_3__924_;
  assign t_4__915_ = t_3__915_ | t_3__923_;
  assign t_4__914_ = t_3__914_ | t_3__922_;
  assign t_4__913_ = t_3__913_ | t_3__921_;
  assign t_4__912_ = t_3__912_ | t_3__920_;
  assign t_4__911_ = t_3__911_ | t_3__919_;
  assign t_4__910_ = t_3__910_ | t_3__918_;
  assign t_4__909_ = t_3__909_ | t_3__917_;
  assign t_4__908_ = t_3__908_ | t_3__916_;
  assign t_4__907_ = t_3__907_ | t_3__915_;
  assign t_4__906_ = t_3__906_ | t_3__914_;
  assign t_4__905_ = t_3__905_ | t_3__913_;
  assign t_4__904_ = t_3__904_ | t_3__912_;
  assign t_4__903_ = t_3__903_ | t_3__911_;
  assign t_4__902_ = t_3__902_ | t_3__910_;
  assign t_4__901_ = t_3__901_ | t_3__909_;
  assign t_4__900_ = t_3__900_ | t_3__908_;
  assign t_4__899_ = t_3__899_ | t_3__907_;
  assign t_4__898_ = t_3__898_ | t_3__906_;
  assign t_4__897_ = t_3__897_ | t_3__905_;
  assign t_4__896_ = t_3__896_ | t_3__904_;
  assign t_4__895_ = t_3__895_ | t_3__903_;
  assign t_4__894_ = t_3__894_ | t_3__902_;
  assign t_4__893_ = t_3__893_ | t_3__901_;
  assign t_4__892_ = t_3__892_ | t_3__900_;
  assign t_4__891_ = t_3__891_ | t_3__899_;
  assign t_4__890_ = t_3__890_ | t_3__898_;
  assign t_4__889_ = t_3__889_ | t_3__897_;
  assign t_4__888_ = t_3__888_ | t_3__896_;
  assign t_4__887_ = t_3__887_ | t_3__895_;
  assign t_4__886_ = t_3__886_ | t_3__894_;
  assign t_4__885_ = t_3__885_ | t_3__893_;
  assign t_4__884_ = t_3__884_ | t_3__892_;
  assign t_4__883_ = t_3__883_ | t_3__891_;
  assign t_4__882_ = t_3__882_ | t_3__890_;
  assign t_4__881_ = t_3__881_ | t_3__889_;
  assign t_4__880_ = t_3__880_ | t_3__888_;
  assign t_4__879_ = t_3__879_ | t_3__887_;
  assign t_4__878_ = t_3__878_ | t_3__886_;
  assign t_4__877_ = t_3__877_ | t_3__885_;
  assign t_4__876_ = t_3__876_ | t_3__884_;
  assign t_4__875_ = t_3__875_ | t_3__883_;
  assign t_4__874_ = t_3__874_ | t_3__882_;
  assign t_4__873_ = t_3__873_ | t_3__881_;
  assign t_4__872_ = t_3__872_ | t_3__880_;
  assign t_4__871_ = t_3__871_ | t_3__879_;
  assign t_4__870_ = t_3__870_ | t_3__878_;
  assign t_4__869_ = t_3__869_ | t_3__877_;
  assign t_4__868_ = t_3__868_ | t_3__876_;
  assign t_4__867_ = t_3__867_ | t_3__875_;
  assign t_4__866_ = t_3__866_ | t_3__874_;
  assign t_4__865_ = t_3__865_ | t_3__873_;
  assign t_4__864_ = t_3__864_ | t_3__872_;
  assign t_4__863_ = t_3__863_ | t_3__871_;
  assign t_4__862_ = t_3__862_ | t_3__870_;
  assign t_4__861_ = t_3__861_ | t_3__869_;
  assign t_4__860_ = t_3__860_ | t_3__868_;
  assign t_4__859_ = t_3__859_ | t_3__867_;
  assign t_4__858_ = t_3__858_ | t_3__866_;
  assign t_4__857_ = t_3__857_ | t_3__865_;
  assign t_4__856_ = t_3__856_ | t_3__864_;
  assign t_4__855_ = t_3__855_ | t_3__863_;
  assign t_4__854_ = t_3__854_ | t_3__862_;
  assign t_4__853_ = t_3__853_ | t_3__861_;
  assign t_4__852_ = t_3__852_ | t_3__860_;
  assign t_4__851_ = t_3__851_ | t_3__859_;
  assign t_4__850_ = t_3__850_ | t_3__858_;
  assign t_4__849_ = t_3__849_ | t_3__857_;
  assign t_4__848_ = t_3__848_ | t_3__856_;
  assign t_4__847_ = t_3__847_ | t_3__855_;
  assign t_4__846_ = t_3__846_ | t_3__854_;
  assign t_4__845_ = t_3__845_ | t_3__853_;
  assign t_4__844_ = t_3__844_ | t_3__852_;
  assign t_4__843_ = t_3__843_ | t_3__851_;
  assign t_4__842_ = t_3__842_ | t_3__850_;
  assign t_4__841_ = t_3__841_ | t_3__849_;
  assign t_4__840_ = t_3__840_ | t_3__848_;
  assign t_4__839_ = t_3__839_ | t_3__847_;
  assign t_4__838_ = t_3__838_ | t_3__846_;
  assign t_4__837_ = t_3__837_ | t_3__845_;
  assign t_4__836_ = t_3__836_ | t_3__844_;
  assign t_4__835_ = t_3__835_ | t_3__843_;
  assign t_4__834_ = t_3__834_ | t_3__842_;
  assign t_4__833_ = t_3__833_ | t_3__841_;
  assign t_4__832_ = t_3__832_ | t_3__840_;
  assign t_4__831_ = t_3__831_ | t_3__839_;
  assign t_4__830_ = t_3__830_ | t_3__838_;
  assign t_4__829_ = t_3__829_ | t_3__837_;
  assign t_4__828_ = t_3__828_ | t_3__836_;
  assign t_4__827_ = t_3__827_ | t_3__835_;
  assign t_4__826_ = t_3__826_ | t_3__834_;
  assign t_4__825_ = t_3__825_ | t_3__833_;
  assign t_4__824_ = t_3__824_ | t_3__832_;
  assign t_4__823_ = t_3__823_ | t_3__831_;
  assign t_4__822_ = t_3__822_ | t_3__830_;
  assign t_4__821_ = t_3__821_ | t_3__829_;
  assign t_4__820_ = t_3__820_ | t_3__828_;
  assign t_4__819_ = t_3__819_ | t_3__827_;
  assign t_4__818_ = t_3__818_ | t_3__826_;
  assign t_4__817_ = t_3__817_ | t_3__825_;
  assign t_4__816_ = t_3__816_ | t_3__824_;
  assign t_4__815_ = t_3__815_ | t_3__823_;
  assign t_4__814_ = t_3__814_ | t_3__822_;
  assign t_4__813_ = t_3__813_ | t_3__821_;
  assign t_4__812_ = t_3__812_ | t_3__820_;
  assign t_4__811_ = t_3__811_ | t_3__819_;
  assign t_4__810_ = t_3__810_ | t_3__818_;
  assign t_4__809_ = t_3__809_ | t_3__817_;
  assign t_4__808_ = t_3__808_ | t_3__816_;
  assign t_4__807_ = t_3__807_ | t_3__815_;
  assign t_4__806_ = t_3__806_ | t_3__814_;
  assign t_4__805_ = t_3__805_ | t_3__813_;
  assign t_4__804_ = t_3__804_ | t_3__812_;
  assign t_4__803_ = t_3__803_ | t_3__811_;
  assign t_4__802_ = t_3__802_ | t_3__810_;
  assign t_4__801_ = t_3__801_ | t_3__809_;
  assign t_4__800_ = t_3__800_ | t_3__808_;
  assign t_4__799_ = t_3__799_ | t_3__807_;
  assign t_4__798_ = t_3__798_ | t_3__806_;
  assign t_4__797_ = t_3__797_ | t_3__805_;
  assign t_4__796_ = t_3__796_ | t_3__804_;
  assign t_4__795_ = t_3__795_ | t_3__803_;
  assign t_4__794_ = t_3__794_ | t_3__802_;
  assign t_4__793_ = t_3__793_ | t_3__801_;
  assign t_4__792_ = t_3__792_ | t_3__800_;
  assign t_4__791_ = t_3__791_ | t_3__799_;
  assign t_4__790_ = t_3__790_ | t_3__798_;
  assign t_4__789_ = t_3__789_ | t_3__797_;
  assign t_4__788_ = t_3__788_ | t_3__796_;
  assign t_4__787_ = t_3__787_ | t_3__795_;
  assign t_4__786_ = t_3__786_ | t_3__794_;
  assign t_4__785_ = t_3__785_ | t_3__793_;
  assign t_4__784_ = t_3__784_ | t_3__792_;
  assign t_4__783_ = t_3__783_ | t_3__791_;
  assign t_4__782_ = t_3__782_ | t_3__790_;
  assign t_4__781_ = t_3__781_ | t_3__789_;
  assign t_4__780_ = t_3__780_ | t_3__788_;
  assign t_4__779_ = t_3__779_ | t_3__787_;
  assign t_4__778_ = t_3__778_ | t_3__786_;
  assign t_4__777_ = t_3__777_ | t_3__785_;
  assign t_4__776_ = t_3__776_ | t_3__784_;
  assign t_4__775_ = t_3__775_ | t_3__783_;
  assign t_4__774_ = t_3__774_ | t_3__782_;
  assign t_4__773_ = t_3__773_ | t_3__781_;
  assign t_4__772_ = t_3__772_ | t_3__780_;
  assign t_4__771_ = t_3__771_ | t_3__779_;
  assign t_4__770_ = t_3__770_ | t_3__778_;
  assign t_4__769_ = t_3__769_ | t_3__777_;
  assign t_4__768_ = t_3__768_ | t_3__776_;
  assign t_4__767_ = t_3__767_ | t_3__775_;
  assign t_4__766_ = t_3__766_ | t_3__774_;
  assign t_4__765_ = t_3__765_ | t_3__773_;
  assign t_4__764_ = t_3__764_ | t_3__772_;
  assign t_4__763_ = t_3__763_ | t_3__771_;
  assign t_4__762_ = t_3__762_ | t_3__770_;
  assign t_4__761_ = t_3__761_ | t_3__769_;
  assign t_4__760_ = t_3__760_ | t_3__768_;
  assign t_4__759_ = t_3__759_ | t_3__767_;
  assign t_4__758_ = t_3__758_ | t_3__766_;
  assign t_4__757_ = t_3__757_ | t_3__765_;
  assign t_4__756_ = t_3__756_ | t_3__764_;
  assign t_4__755_ = t_3__755_ | t_3__763_;
  assign t_4__754_ = t_3__754_ | t_3__762_;
  assign t_4__753_ = t_3__753_ | t_3__761_;
  assign t_4__752_ = t_3__752_ | t_3__760_;
  assign t_4__751_ = t_3__751_ | t_3__759_;
  assign t_4__750_ = t_3__750_ | t_3__758_;
  assign t_4__749_ = t_3__749_ | t_3__757_;
  assign t_4__748_ = t_3__748_ | t_3__756_;
  assign t_4__747_ = t_3__747_ | t_3__755_;
  assign t_4__746_ = t_3__746_ | t_3__754_;
  assign t_4__745_ = t_3__745_ | t_3__753_;
  assign t_4__744_ = t_3__744_ | t_3__752_;
  assign t_4__743_ = t_3__743_ | t_3__751_;
  assign t_4__742_ = t_3__742_ | t_3__750_;
  assign t_4__741_ = t_3__741_ | t_3__749_;
  assign t_4__740_ = t_3__740_ | t_3__748_;
  assign t_4__739_ = t_3__739_ | t_3__747_;
  assign t_4__738_ = t_3__738_ | t_3__746_;
  assign t_4__737_ = t_3__737_ | t_3__745_;
  assign t_4__736_ = t_3__736_ | t_3__744_;
  assign t_4__735_ = t_3__735_ | t_3__743_;
  assign t_4__734_ = t_3__734_ | t_3__742_;
  assign t_4__733_ = t_3__733_ | t_3__741_;
  assign t_4__732_ = t_3__732_ | t_3__740_;
  assign t_4__731_ = t_3__731_ | t_3__739_;
  assign t_4__730_ = t_3__730_ | t_3__738_;
  assign t_4__729_ = t_3__729_ | t_3__737_;
  assign t_4__728_ = t_3__728_ | t_3__736_;
  assign t_4__727_ = t_3__727_ | t_3__735_;
  assign t_4__726_ = t_3__726_ | t_3__734_;
  assign t_4__725_ = t_3__725_ | t_3__733_;
  assign t_4__724_ = t_3__724_ | t_3__732_;
  assign t_4__723_ = t_3__723_ | t_3__731_;
  assign t_4__722_ = t_3__722_ | t_3__730_;
  assign t_4__721_ = t_3__721_ | t_3__729_;
  assign t_4__720_ = t_3__720_ | t_3__728_;
  assign t_4__719_ = t_3__719_ | t_3__727_;
  assign t_4__718_ = t_3__718_ | t_3__726_;
  assign t_4__717_ = t_3__717_ | t_3__725_;
  assign t_4__716_ = t_3__716_ | t_3__724_;
  assign t_4__715_ = t_3__715_ | t_3__723_;
  assign t_4__714_ = t_3__714_ | t_3__722_;
  assign t_4__713_ = t_3__713_ | t_3__721_;
  assign t_4__712_ = t_3__712_ | t_3__720_;
  assign t_4__711_ = t_3__711_ | t_3__719_;
  assign t_4__710_ = t_3__710_ | t_3__718_;
  assign t_4__709_ = t_3__709_ | t_3__717_;
  assign t_4__708_ = t_3__708_ | t_3__716_;
  assign t_4__707_ = t_3__707_ | t_3__715_;
  assign t_4__706_ = t_3__706_ | t_3__714_;
  assign t_4__705_ = t_3__705_ | t_3__713_;
  assign t_4__704_ = t_3__704_ | t_3__712_;
  assign t_4__703_ = t_3__703_ | t_3__711_;
  assign t_4__702_ = t_3__702_ | t_3__710_;
  assign t_4__701_ = t_3__701_ | t_3__709_;
  assign t_4__700_ = t_3__700_ | t_3__708_;
  assign t_4__699_ = t_3__699_ | t_3__707_;
  assign t_4__698_ = t_3__698_ | t_3__706_;
  assign t_4__697_ = t_3__697_ | t_3__705_;
  assign t_4__696_ = t_3__696_ | t_3__704_;
  assign t_4__695_ = t_3__695_ | t_3__703_;
  assign t_4__694_ = t_3__694_ | t_3__702_;
  assign t_4__693_ = t_3__693_ | t_3__701_;
  assign t_4__692_ = t_3__692_ | t_3__700_;
  assign t_4__691_ = t_3__691_ | t_3__699_;
  assign t_4__690_ = t_3__690_ | t_3__698_;
  assign t_4__689_ = t_3__689_ | t_3__697_;
  assign t_4__688_ = t_3__688_ | t_3__696_;
  assign t_4__687_ = t_3__687_ | t_3__695_;
  assign t_4__686_ = t_3__686_ | t_3__694_;
  assign t_4__685_ = t_3__685_ | t_3__693_;
  assign t_4__684_ = t_3__684_ | t_3__692_;
  assign t_4__683_ = t_3__683_ | t_3__691_;
  assign t_4__682_ = t_3__682_ | t_3__690_;
  assign t_4__681_ = t_3__681_ | t_3__689_;
  assign t_4__680_ = t_3__680_ | t_3__688_;
  assign t_4__679_ = t_3__679_ | t_3__687_;
  assign t_4__678_ = t_3__678_ | t_3__686_;
  assign t_4__677_ = t_3__677_ | t_3__685_;
  assign t_4__676_ = t_3__676_ | t_3__684_;
  assign t_4__675_ = t_3__675_ | t_3__683_;
  assign t_4__674_ = t_3__674_ | t_3__682_;
  assign t_4__673_ = t_3__673_ | t_3__681_;
  assign t_4__672_ = t_3__672_ | t_3__680_;
  assign t_4__671_ = t_3__671_ | t_3__679_;
  assign t_4__670_ = t_3__670_ | t_3__678_;
  assign t_4__669_ = t_3__669_ | t_3__677_;
  assign t_4__668_ = t_3__668_ | t_3__676_;
  assign t_4__667_ = t_3__667_ | t_3__675_;
  assign t_4__666_ = t_3__666_ | t_3__674_;
  assign t_4__665_ = t_3__665_ | t_3__673_;
  assign t_4__664_ = t_3__664_ | t_3__672_;
  assign t_4__663_ = t_3__663_ | t_3__671_;
  assign t_4__662_ = t_3__662_ | t_3__670_;
  assign t_4__661_ = t_3__661_ | t_3__669_;
  assign t_4__660_ = t_3__660_ | t_3__668_;
  assign t_4__659_ = t_3__659_ | t_3__667_;
  assign t_4__658_ = t_3__658_ | t_3__666_;
  assign t_4__657_ = t_3__657_ | t_3__665_;
  assign t_4__656_ = t_3__656_ | t_3__664_;
  assign t_4__655_ = t_3__655_ | t_3__663_;
  assign t_4__654_ = t_3__654_ | t_3__662_;
  assign t_4__653_ = t_3__653_ | t_3__661_;
  assign t_4__652_ = t_3__652_ | t_3__660_;
  assign t_4__651_ = t_3__651_ | t_3__659_;
  assign t_4__650_ = t_3__650_ | t_3__658_;
  assign t_4__649_ = t_3__649_ | t_3__657_;
  assign t_4__648_ = t_3__648_ | t_3__656_;
  assign t_4__647_ = t_3__647_ | t_3__655_;
  assign t_4__646_ = t_3__646_ | t_3__654_;
  assign t_4__645_ = t_3__645_ | t_3__653_;
  assign t_4__644_ = t_3__644_ | t_3__652_;
  assign t_4__643_ = t_3__643_ | t_3__651_;
  assign t_4__642_ = t_3__642_ | t_3__650_;
  assign t_4__641_ = t_3__641_ | t_3__649_;
  assign t_4__640_ = t_3__640_ | t_3__648_;
  assign t_4__639_ = t_3__639_ | t_3__647_;
  assign t_4__638_ = t_3__638_ | t_3__646_;
  assign t_4__637_ = t_3__637_ | t_3__645_;
  assign t_4__636_ = t_3__636_ | t_3__644_;
  assign t_4__635_ = t_3__635_ | t_3__643_;
  assign t_4__634_ = t_3__634_ | t_3__642_;
  assign t_4__633_ = t_3__633_ | t_3__641_;
  assign t_4__632_ = t_3__632_ | t_3__640_;
  assign t_4__631_ = t_3__631_ | t_3__639_;
  assign t_4__630_ = t_3__630_ | t_3__638_;
  assign t_4__629_ = t_3__629_ | t_3__637_;
  assign t_4__628_ = t_3__628_ | t_3__636_;
  assign t_4__627_ = t_3__627_ | t_3__635_;
  assign t_4__626_ = t_3__626_ | t_3__634_;
  assign t_4__625_ = t_3__625_ | t_3__633_;
  assign t_4__624_ = t_3__624_ | t_3__632_;
  assign t_4__623_ = t_3__623_ | t_3__631_;
  assign t_4__622_ = t_3__622_ | t_3__630_;
  assign t_4__621_ = t_3__621_ | t_3__629_;
  assign t_4__620_ = t_3__620_ | t_3__628_;
  assign t_4__619_ = t_3__619_ | t_3__627_;
  assign t_4__618_ = t_3__618_ | t_3__626_;
  assign t_4__617_ = t_3__617_ | t_3__625_;
  assign t_4__616_ = t_3__616_ | t_3__624_;
  assign t_4__615_ = t_3__615_ | t_3__623_;
  assign t_4__614_ = t_3__614_ | t_3__622_;
  assign t_4__613_ = t_3__613_ | t_3__621_;
  assign t_4__612_ = t_3__612_ | t_3__620_;
  assign t_4__611_ = t_3__611_ | t_3__619_;
  assign t_4__610_ = t_3__610_ | t_3__618_;
  assign t_4__609_ = t_3__609_ | t_3__617_;
  assign t_4__608_ = t_3__608_ | t_3__616_;
  assign t_4__607_ = t_3__607_ | t_3__615_;
  assign t_4__606_ = t_3__606_ | t_3__614_;
  assign t_4__605_ = t_3__605_ | t_3__613_;
  assign t_4__604_ = t_3__604_ | t_3__612_;
  assign t_4__603_ = t_3__603_ | t_3__611_;
  assign t_4__602_ = t_3__602_ | t_3__610_;
  assign t_4__601_ = t_3__601_ | t_3__609_;
  assign t_4__600_ = t_3__600_ | t_3__608_;
  assign t_4__599_ = t_3__599_ | t_3__607_;
  assign t_4__598_ = t_3__598_ | t_3__606_;
  assign t_4__597_ = t_3__597_ | t_3__605_;
  assign t_4__596_ = t_3__596_ | t_3__604_;
  assign t_4__595_ = t_3__595_ | t_3__603_;
  assign t_4__594_ = t_3__594_ | t_3__602_;
  assign t_4__593_ = t_3__593_ | t_3__601_;
  assign t_4__592_ = t_3__592_ | t_3__600_;
  assign t_4__591_ = t_3__591_ | t_3__599_;
  assign t_4__590_ = t_3__590_ | t_3__598_;
  assign t_4__589_ = t_3__589_ | t_3__597_;
  assign t_4__588_ = t_3__588_ | t_3__596_;
  assign t_4__587_ = t_3__587_ | t_3__595_;
  assign t_4__586_ = t_3__586_ | t_3__594_;
  assign t_4__585_ = t_3__585_ | t_3__593_;
  assign t_4__584_ = t_3__584_ | t_3__592_;
  assign t_4__583_ = t_3__583_ | t_3__591_;
  assign t_4__582_ = t_3__582_ | t_3__590_;
  assign t_4__581_ = t_3__581_ | t_3__589_;
  assign t_4__580_ = t_3__580_ | t_3__588_;
  assign t_4__579_ = t_3__579_ | t_3__587_;
  assign t_4__578_ = t_3__578_ | t_3__586_;
  assign t_4__577_ = t_3__577_ | t_3__585_;
  assign t_4__576_ = t_3__576_ | t_3__584_;
  assign t_4__575_ = t_3__575_ | t_3__583_;
  assign t_4__574_ = t_3__574_ | t_3__582_;
  assign t_4__573_ = t_3__573_ | t_3__581_;
  assign t_4__572_ = t_3__572_ | t_3__580_;
  assign t_4__571_ = t_3__571_ | t_3__579_;
  assign t_4__570_ = t_3__570_ | t_3__578_;
  assign t_4__569_ = t_3__569_ | t_3__577_;
  assign t_4__568_ = t_3__568_ | t_3__576_;
  assign t_4__567_ = t_3__567_ | t_3__575_;
  assign t_4__566_ = t_3__566_ | t_3__574_;
  assign t_4__565_ = t_3__565_ | t_3__573_;
  assign t_4__564_ = t_3__564_ | t_3__572_;
  assign t_4__563_ = t_3__563_ | t_3__571_;
  assign t_4__562_ = t_3__562_ | t_3__570_;
  assign t_4__561_ = t_3__561_ | t_3__569_;
  assign t_4__560_ = t_3__560_ | t_3__568_;
  assign t_4__559_ = t_3__559_ | t_3__567_;
  assign t_4__558_ = t_3__558_ | t_3__566_;
  assign t_4__557_ = t_3__557_ | t_3__565_;
  assign t_4__556_ = t_3__556_ | t_3__564_;
  assign t_4__555_ = t_3__555_ | t_3__563_;
  assign t_4__554_ = t_3__554_ | t_3__562_;
  assign t_4__553_ = t_3__553_ | t_3__561_;
  assign t_4__552_ = t_3__552_ | t_3__560_;
  assign t_4__551_ = t_3__551_ | t_3__559_;
  assign t_4__550_ = t_3__550_ | t_3__558_;
  assign t_4__549_ = t_3__549_ | t_3__557_;
  assign t_4__548_ = t_3__548_ | t_3__556_;
  assign t_4__547_ = t_3__547_ | t_3__555_;
  assign t_4__546_ = t_3__546_ | t_3__554_;
  assign t_4__545_ = t_3__545_ | t_3__553_;
  assign t_4__544_ = t_3__544_ | t_3__552_;
  assign t_4__543_ = t_3__543_ | t_3__551_;
  assign t_4__542_ = t_3__542_ | t_3__550_;
  assign t_4__541_ = t_3__541_ | t_3__549_;
  assign t_4__540_ = t_3__540_ | t_3__548_;
  assign t_4__539_ = t_3__539_ | t_3__547_;
  assign t_4__538_ = t_3__538_ | t_3__546_;
  assign t_4__537_ = t_3__537_ | t_3__545_;
  assign t_4__536_ = t_3__536_ | t_3__544_;
  assign t_4__535_ = t_3__535_ | t_3__543_;
  assign t_4__534_ = t_3__534_ | t_3__542_;
  assign t_4__533_ = t_3__533_ | t_3__541_;
  assign t_4__532_ = t_3__532_ | t_3__540_;
  assign t_4__531_ = t_3__531_ | t_3__539_;
  assign t_4__530_ = t_3__530_ | t_3__538_;
  assign t_4__529_ = t_3__529_ | t_3__537_;
  assign t_4__528_ = t_3__528_ | t_3__536_;
  assign t_4__527_ = t_3__527_ | t_3__535_;
  assign t_4__526_ = t_3__526_ | t_3__534_;
  assign t_4__525_ = t_3__525_ | t_3__533_;
  assign t_4__524_ = t_3__524_ | t_3__532_;
  assign t_4__523_ = t_3__523_ | t_3__531_;
  assign t_4__522_ = t_3__522_ | t_3__530_;
  assign t_4__521_ = t_3__521_ | t_3__529_;
  assign t_4__520_ = t_3__520_ | t_3__528_;
  assign t_4__519_ = t_3__519_ | t_3__527_;
  assign t_4__518_ = t_3__518_ | t_3__526_;
  assign t_4__517_ = t_3__517_ | t_3__525_;
  assign t_4__516_ = t_3__516_ | t_3__524_;
  assign t_4__515_ = t_3__515_ | t_3__523_;
  assign t_4__514_ = t_3__514_ | t_3__522_;
  assign t_4__513_ = t_3__513_ | t_3__521_;
  assign t_4__512_ = t_3__512_ | t_3__520_;
  assign t_4__511_ = t_3__511_ | t_3__519_;
  assign t_4__510_ = t_3__510_ | t_3__518_;
  assign t_4__509_ = t_3__509_ | t_3__517_;
  assign t_4__508_ = t_3__508_ | t_3__516_;
  assign t_4__507_ = t_3__507_ | t_3__515_;
  assign t_4__506_ = t_3__506_ | t_3__514_;
  assign t_4__505_ = t_3__505_ | t_3__513_;
  assign t_4__504_ = t_3__504_ | t_3__512_;
  assign t_4__503_ = t_3__503_ | t_3__511_;
  assign t_4__502_ = t_3__502_ | t_3__510_;
  assign t_4__501_ = t_3__501_ | t_3__509_;
  assign t_4__500_ = t_3__500_ | t_3__508_;
  assign t_4__499_ = t_3__499_ | t_3__507_;
  assign t_4__498_ = t_3__498_ | t_3__506_;
  assign t_4__497_ = t_3__497_ | t_3__505_;
  assign t_4__496_ = t_3__496_ | t_3__504_;
  assign t_4__495_ = t_3__495_ | t_3__503_;
  assign t_4__494_ = t_3__494_ | t_3__502_;
  assign t_4__493_ = t_3__493_ | t_3__501_;
  assign t_4__492_ = t_3__492_ | t_3__500_;
  assign t_4__491_ = t_3__491_ | t_3__499_;
  assign t_4__490_ = t_3__490_ | t_3__498_;
  assign t_4__489_ = t_3__489_ | t_3__497_;
  assign t_4__488_ = t_3__488_ | t_3__496_;
  assign t_4__487_ = t_3__487_ | t_3__495_;
  assign t_4__486_ = t_3__486_ | t_3__494_;
  assign t_4__485_ = t_3__485_ | t_3__493_;
  assign t_4__484_ = t_3__484_ | t_3__492_;
  assign t_4__483_ = t_3__483_ | t_3__491_;
  assign t_4__482_ = t_3__482_ | t_3__490_;
  assign t_4__481_ = t_3__481_ | t_3__489_;
  assign t_4__480_ = t_3__480_ | t_3__488_;
  assign t_4__479_ = t_3__479_ | t_3__487_;
  assign t_4__478_ = t_3__478_ | t_3__486_;
  assign t_4__477_ = t_3__477_ | t_3__485_;
  assign t_4__476_ = t_3__476_ | t_3__484_;
  assign t_4__475_ = t_3__475_ | t_3__483_;
  assign t_4__474_ = t_3__474_ | t_3__482_;
  assign t_4__473_ = t_3__473_ | t_3__481_;
  assign t_4__472_ = t_3__472_ | t_3__480_;
  assign t_4__471_ = t_3__471_ | t_3__479_;
  assign t_4__470_ = t_3__470_ | t_3__478_;
  assign t_4__469_ = t_3__469_ | t_3__477_;
  assign t_4__468_ = t_3__468_ | t_3__476_;
  assign t_4__467_ = t_3__467_ | t_3__475_;
  assign t_4__466_ = t_3__466_ | t_3__474_;
  assign t_4__465_ = t_3__465_ | t_3__473_;
  assign t_4__464_ = t_3__464_ | t_3__472_;
  assign t_4__463_ = t_3__463_ | t_3__471_;
  assign t_4__462_ = t_3__462_ | t_3__470_;
  assign t_4__461_ = t_3__461_ | t_3__469_;
  assign t_4__460_ = t_3__460_ | t_3__468_;
  assign t_4__459_ = t_3__459_ | t_3__467_;
  assign t_4__458_ = t_3__458_ | t_3__466_;
  assign t_4__457_ = t_3__457_ | t_3__465_;
  assign t_4__456_ = t_3__456_ | t_3__464_;
  assign t_4__455_ = t_3__455_ | t_3__463_;
  assign t_4__454_ = t_3__454_ | t_3__462_;
  assign t_4__453_ = t_3__453_ | t_3__461_;
  assign t_4__452_ = t_3__452_ | t_3__460_;
  assign t_4__451_ = t_3__451_ | t_3__459_;
  assign t_4__450_ = t_3__450_ | t_3__458_;
  assign t_4__449_ = t_3__449_ | t_3__457_;
  assign t_4__448_ = t_3__448_ | t_3__456_;
  assign t_4__447_ = t_3__447_ | t_3__455_;
  assign t_4__446_ = t_3__446_ | t_3__454_;
  assign t_4__445_ = t_3__445_ | t_3__453_;
  assign t_4__444_ = t_3__444_ | t_3__452_;
  assign t_4__443_ = t_3__443_ | t_3__451_;
  assign t_4__442_ = t_3__442_ | t_3__450_;
  assign t_4__441_ = t_3__441_ | t_3__449_;
  assign t_4__440_ = t_3__440_ | t_3__448_;
  assign t_4__439_ = t_3__439_ | t_3__447_;
  assign t_4__438_ = t_3__438_ | t_3__446_;
  assign t_4__437_ = t_3__437_ | t_3__445_;
  assign t_4__436_ = t_3__436_ | t_3__444_;
  assign t_4__435_ = t_3__435_ | t_3__443_;
  assign t_4__434_ = t_3__434_ | t_3__442_;
  assign t_4__433_ = t_3__433_ | t_3__441_;
  assign t_4__432_ = t_3__432_ | t_3__440_;
  assign t_4__431_ = t_3__431_ | t_3__439_;
  assign t_4__430_ = t_3__430_ | t_3__438_;
  assign t_4__429_ = t_3__429_ | t_3__437_;
  assign t_4__428_ = t_3__428_ | t_3__436_;
  assign t_4__427_ = t_3__427_ | t_3__435_;
  assign t_4__426_ = t_3__426_ | t_3__434_;
  assign t_4__425_ = t_3__425_ | t_3__433_;
  assign t_4__424_ = t_3__424_ | t_3__432_;
  assign t_4__423_ = t_3__423_ | t_3__431_;
  assign t_4__422_ = t_3__422_ | t_3__430_;
  assign t_4__421_ = t_3__421_ | t_3__429_;
  assign t_4__420_ = t_3__420_ | t_3__428_;
  assign t_4__419_ = t_3__419_ | t_3__427_;
  assign t_4__418_ = t_3__418_ | t_3__426_;
  assign t_4__417_ = t_3__417_ | t_3__425_;
  assign t_4__416_ = t_3__416_ | t_3__424_;
  assign t_4__415_ = t_3__415_ | t_3__423_;
  assign t_4__414_ = t_3__414_ | t_3__422_;
  assign t_4__413_ = t_3__413_ | t_3__421_;
  assign t_4__412_ = t_3__412_ | t_3__420_;
  assign t_4__411_ = t_3__411_ | t_3__419_;
  assign t_4__410_ = t_3__410_ | t_3__418_;
  assign t_4__409_ = t_3__409_ | t_3__417_;
  assign t_4__408_ = t_3__408_ | t_3__416_;
  assign t_4__407_ = t_3__407_ | t_3__415_;
  assign t_4__406_ = t_3__406_ | t_3__414_;
  assign t_4__405_ = t_3__405_ | t_3__413_;
  assign t_4__404_ = t_3__404_ | t_3__412_;
  assign t_4__403_ = t_3__403_ | t_3__411_;
  assign t_4__402_ = t_3__402_ | t_3__410_;
  assign t_4__401_ = t_3__401_ | t_3__409_;
  assign t_4__400_ = t_3__400_ | t_3__408_;
  assign t_4__399_ = t_3__399_ | t_3__407_;
  assign t_4__398_ = t_3__398_ | t_3__406_;
  assign t_4__397_ = t_3__397_ | t_3__405_;
  assign t_4__396_ = t_3__396_ | t_3__404_;
  assign t_4__395_ = t_3__395_ | t_3__403_;
  assign t_4__394_ = t_3__394_ | t_3__402_;
  assign t_4__393_ = t_3__393_ | t_3__401_;
  assign t_4__392_ = t_3__392_ | t_3__400_;
  assign t_4__391_ = t_3__391_ | t_3__399_;
  assign t_4__390_ = t_3__390_ | t_3__398_;
  assign t_4__389_ = t_3__389_ | t_3__397_;
  assign t_4__388_ = t_3__388_ | t_3__396_;
  assign t_4__387_ = t_3__387_ | t_3__395_;
  assign t_4__386_ = t_3__386_ | t_3__394_;
  assign t_4__385_ = t_3__385_ | t_3__393_;
  assign t_4__384_ = t_3__384_ | t_3__392_;
  assign t_4__383_ = t_3__383_ | t_3__391_;
  assign t_4__382_ = t_3__382_ | t_3__390_;
  assign t_4__381_ = t_3__381_ | t_3__389_;
  assign t_4__380_ = t_3__380_ | t_3__388_;
  assign t_4__379_ = t_3__379_ | t_3__387_;
  assign t_4__378_ = t_3__378_ | t_3__386_;
  assign t_4__377_ = t_3__377_ | t_3__385_;
  assign t_4__376_ = t_3__376_ | t_3__384_;
  assign t_4__375_ = t_3__375_ | t_3__383_;
  assign t_4__374_ = t_3__374_ | t_3__382_;
  assign t_4__373_ = t_3__373_ | t_3__381_;
  assign t_4__372_ = t_3__372_ | t_3__380_;
  assign t_4__371_ = t_3__371_ | t_3__379_;
  assign t_4__370_ = t_3__370_ | t_3__378_;
  assign t_4__369_ = t_3__369_ | t_3__377_;
  assign t_4__368_ = t_3__368_ | t_3__376_;
  assign t_4__367_ = t_3__367_ | t_3__375_;
  assign t_4__366_ = t_3__366_ | t_3__374_;
  assign t_4__365_ = t_3__365_ | t_3__373_;
  assign t_4__364_ = t_3__364_ | t_3__372_;
  assign t_4__363_ = t_3__363_ | t_3__371_;
  assign t_4__362_ = t_3__362_ | t_3__370_;
  assign t_4__361_ = t_3__361_ | t_3__369_;
  assign t_4__360_ = t_3__360_ | t_3__368_;
  assign t_4__359_ = t_3__359_ | t_3__367_;
  assign t_4__358_ = t_3__358_ | t_3__366_;
  assign t_4__357_ = t_3__357_ | t_3__365_;
  assign t_4__356_ = t_3__356_ | t_3__364_;
  assign t_4__355_ = t_3__355_ | t_3__363_;
  assign t_4__354_ = t_3__354_ | t_3__362_;
  assign t_4__353_ = t_3__353_ | t_3__361_;
  assign t_4__352_ = t_3__352_ | t_3__360_;
  assign t_4__351_ = t_3__351_ | t_3__359_;
  assign t_4__350_ = t_3__350_ | t_3__358_;
  assign t_4__349_ = t_3__349_ | t_3__357_;
  assign t_4__348_ = t_3__348_ | t_3__356_;
  assign t_4__347_ = t_3__347_ | t_3__355_;
  assign t_4__346_ = t_3__346_ | t_3__354_;
  assign t_4__345_ = t_3__345_ | t_3__353_;
  assign t_4__344_ = t_3__344_ | t_3__352_;
  assign t_4__343_ = t_3__343_ | t_3__351_;
  assign t_4__342_ = t_3__342_ | t_3__350_;
  assign t_4__341_ = t_3__341_ | t_3__349_;
  assign t_4__340_ = t_3__340_ | t_3__348_;
  assign t_4__339_ = t_3__339_ | t_3__347_;
  assign t_4__338_ = t_3__338_ | t_3__346_;
  assign t_4__337_ = t_3__337_ | t_3__345_;
  assign t_4__336_ = t_3__336_ | t_3__344_;
  assign t_4__335_ = t_3__335_ | t_3__343_;
  assign t_4__334_ = t_3__334_ | t_3__342_;
  assign t_4__333_ = t_3__333_ | t_3__341_;
  assign t_4__332_ = t_3__332_ | t_3__340_;
  assign t_4__331_ = t_3__331_ | t_3__339_;
  assign t_4__330_ = t_3__330_ | t_3__338_;
  assign t_4__329_ = t_3__329_ | t_3__337_;
  assign t_4__328_ = t_3__328_ | t_3__336_;
  assign t_4__327_ = t_3__327_ | t_3__335_;
  assign t_4__326_ = t_3__326_ | t_3__334_;
  assign t_4__325_ = t_3__325_ | t_3__333_;
  assign t_4__324_ = t_3__324_ | t_3__332_;
  assign t_4__323_ = t_3__323_ | t_3__331_;
  assign t_4__322_ = t_3__322_ | t_3__330_;
  assign t_4__321_ = t_3__321_ | t_3__329_;
  assign t_4__320_ = t_3__320_ | t_3__328_;
  assign t_4__319_ = t_3__319_ | t_3__327_;
  assign t_4__318_ = t_3__318_ | t_3__326_;
  assign t_4__317_ = t_3__317_ | t_3__325_;
  assign t_4__316_ = t_3__316_ | t_3__324_;
  assign t_4__315_ = t_3__315_ | t_3__323_;
  assign t_4__314_ = t_3__314_ | t_3__322_;
  assign t_4__313_ = t_3__313_ | t_3__321_;
  assign t_4__312_ = t_3__312_ | t_3__320_;
  assign t_4__311_ = t_3__311_ | t_3__319_;
  assign t_4__310_ = t_3__310_ | t_3__318_;
  assign t_4__309_ = t_3__309_ | t_3__317_;
  assign t_4__308_ = t_3__308_ | t_3__316_;
  assign t_4__307_ = t_3__307_ | t_3__315_;
  assign t_4__306_ = t_3__306_ | t_3__314_;
  assign t_4__305_ = t_3__305_ | t_3__313_;
  assign t_4__304_ = t_3__304_ | t_3__312_;
  assign t_4__303_ = t_3__303_ | t_3__311_;
  assign t_4__302_ = t_3__302_ | t_3__310_;
  assign t_4__301_ = t_3__301_ | t_3__309_;
  assign t_4__300_ = t_3__300_ | t_3__308_;
  assign t_4__299_ = t_3__299_ | t_3__307_;
  assign t_4__298_ = t_3__298_ | t_3__306_;
  assign t_4__297_ = t_3__297_ | t_3__305_;
  assign t_4__296_ = t_3__296_ | t_3__304_;
  assign t_4__295_ = t_3__295_ | t_3__303_;
  assign t_4__294_ = t_3__294_ | t_3__302_;
  assign t_4__293_ = t_3__293_ | t_3__301_;
  assign t_4__292_ = t_3__292_ | t_3__300_;
  assign t_4__291_ = t_3__291_ | t_3__299_;
  assign t_4__290_ = t_3__290_ | t_3__298_;
  assign t_4__289_ = t_3__289_ | t_3__297_;
  assign t_4__288_ = t_3__288_ | t_3__296_;
  assign t_4__287_ = t_3__287_ | t_3__295_;
  assign t_4__286_ = t_3__286_ | t_3__294_;
  assign t_4__285_ = t_3__285_ | t_3__293_;
  assign t_4__284_ = t_3__284_ | t_3__292_;
  assign t_4__283_ = t_3__283_ | t_3__291_;
  assign t_4__282_ = t_3__282_ | t_3__290_;
  assign t_4__281_ = t_3__281_ | t_3__289_;
  assign t_4__280_ = t_3__280_ | t_3__288_;
  assign t_4__279_ = t_3__279_ | t_3__287_;
  assign t_4__278_ = t_3__278_ | t_3__286_;
  assign t_4__277_ = t_3__277_ | t_3__285_;
  assign t_4__276_ = t_3__276_ | t_3__284_;
  assign t_4__275_ = t_3__275_ | t_3__283_;
  assign t_4__274_ = t_3__274_ | t_3__282_;
  assign t_4__273_ = t_3__273_ | t_3__281_;
  assign t_4__272_ = t_3__272_ | t_3__280_;
  assign t_4__271_ = t_3__271_ | t_3__279_;
  assign t_4__270_ = t_3__270_ | t_3__278_;
  assign t_4__269_ = t_3__269_ | t_3__277_;
  assign t_4__268_ = t_3__268_ | t_3__276_;
  assign t_4__267_ = t_3__267_ | t_3__275_;
  assign t_4__266_ = t_3__266_ | t_3__274_;
  assign t_4__265_ = t_3__265_ | t_3__273_;
  assign t_4__264_ = t_3__264_ | t_3__272_;
  assign t_4__263_ = t_3__263_ | t_3__271_;
  assign t_4__262_ = t_3__262_ | t_3__270_;
  assign t_4__261_ = t_3__261_ | t_3__269_;
  assign t_4__260_ = t_3__260_ | t_3__268_;
  assign t_4__259_ = t_3__259_ | t_3__267_;
  assign t_4__258_ = t_3__258_ | t_3__266_;
  assign t_4__257_ = t_3__257_ | t_3__265_;
  assign t_4__256_ = t_3__256_ | t_3__264_;
  assign t_4__255_ = t_3__255_ | t_3__263_;
  assign t_4__254_ = t_3__254_ | t_3__262_;
  assign t_4__253_ = t_3__253_ | t_3__261_;
  assign t_4__252_ = t_3__252_ | t_3__260_;
  assign t_4__251_ = t_3__251_ | t_3__259_;
  assign t_4__250_ = t_3__250_ | t_3__258_;
  assign t_4__249_ = t_3__249_ | t_3__257_;
  assign t_4__248_ = t_3__248_ | t_3__256_;
  assign t_4__247_ = t_3__247_ | t_3__255_;
  assign t_4__246_ = t_3__246_ | t_3__254_;
  assign t_4__245_ = t_3__245_ | t_3__253_;
  assign t_4__244_ = t_3__244_ | t_3__252_;
  assign t_4__243_ = t_3__243_ | t_3__251_;
  assign t_4__242_ = t_3__242_ | t_3__250_;
  assign t_4__241_ = t_3__241_ | t_3__249_;
  assign t_4__240_ = t_3__240_ | t_3__248_;
  assign t_4__239_ = t_3__239_ | t_3__247_;
  assign t_4__238_ = t_3__238_ | t_3__246_;
  assign t_4__237_ = t_3__237_ | t_3__245_;
  assign t_4__236_ = t_3__236_ | t_3__244_;
  assign t_4__235_ = t_3__235_ | t_3__243_;
  assign t_4__234_ = t_3__234_ | t_3__242_;
  assign t_4__233_ = t_3__233_ | t_3__241_;
  assign t_4__232_ = t_3__232_ | t_3__240_;
  assign t_4__231_ = t_3__231_ | t_3__239_;
  assign t_4__230_ = t_3__230_ | t_3__238_;
  assign t_4__229_ = t_3__229_ | t_3__237_;
  assign t_4__228_ = t_3__228_ | t_3__236_;
  assign t_4__227_ = t_3__227_ | t_3__235_;
  assign t_4__226_ = t_3__226_ | t_3__234_;
  assign t_4__225_ = t_3__225_ | t_3__233_;
  assign t_4__224_ = t_3__224_ | t_3__232_;
  assign t_4__223_ = t_3__223_ | t_3__231_;
  assign t_4__222_ = t_3__222_ | t_3__230_;
  assign t_4__221_ = t_3__221_ | t_3__229_;
  assign t_4__220_ = t_3__220_ | t_3__228_;
  assign t_4__219_ = t_3__219_ | t_3__227_;
  assign t_4__218_ = t_3__218_ | t_3__226_;
  assign t_4__217_ = t_3__217_ | t_3__225_;
  assign t_4__216_ = t_3__216_ | t_3__224_;
  assign t_4__215_ = t_3__215_ | t_3__223_;
  assign t_4__214_ = t_3__214_ | t_3__222_;
  assign t_4__213_ = t_3__213_ | t_3__221_;
  assign t_4__212_ = t_3__212_ | t_3__220_;
  assign t_4__211_ = t_3__211_ | t_3__219_;
  assign t_4__210_ = t_3__210_ | t_3__218_;
  assign t_4__209_ = t_3__209_ | t_3__217_;
  assign t_4__208_ = t_3__208_ | t_3__216_;
  assign t_4__207_ = t_3__207_ | t_3__215_;
  assign t_4__206_ = t_3__206_ | t_3__214_;
  assign t_4__205_ = t_3__205_ | t_3__213_;
  assign t_4__204_ = t_3__204_ | t_3__212_;
  assign t_4__203_ = t_3__203_ | t_3__211_;
  assign t_4__202_ = t_3__202_ | t_3__210_;
  assign t_4__201_ = t_3__201_ | t_3__209_;
  assign t_4__200_ = t_3__200_ | t_3__208_;
  assign t_4__199_ = t_3__199_ | t_3__207_;
  assign t_4__198_ = t_3__198_ | t_3__206_;
  assign t_4__197_ = t_3__197_ | t_3__205_;
  assign t_4__196_ = t_3__196_ | t_3__204_;
  assign t_4__195_ = t_3__195_ | t_3__203_;
  assign t_4__194_ = t_3__194_ | t_3__202_;
  assign t_4__193_ = t_3__193_ | t_3__201_;
  assign t_4__192_ = t_3__192_ | t_3__200_;
  assign t_4__191_ = t_3__191_ | t_3__199_;
  assign t_4__190_ = t_3__190_ | t_3__198_;
  assign t_4__189_ = t_3__189_ | t_3__197_;
  assign t_4__188_ = t_3__188_ | t_3__196_;
  assign t_4__187_ = t_3__187_ | t_3__195_;
  assign t_4__186_ = t_3__186_ | t_3__194_;
  assign t_4__185_ = t_3__185_ | t_3__193_;
  assign t_4__184_ = t_3__184_ | t_3__192_;
  assign t_4__183_ = t_3__183_ | t_3__191_;
  assign t_4__182_ = t_3__182_ | t_3__190_;
  assign t_4__181_ = t_3__181_ | t_3__189_;
  assign t_4__180_ = t_3__180_ | t_3__188_;
  assign t_4__179_ = t_3__179_ | t_3__187_;
  assign t_4__178_ = t_3__178_ | t_3__186_;
  assign t_4__177_ = t_3__177_ | t_3__185_;
  assign t_4__176_ = t_3__176_ | t_3__184_;
  assign t_4__175_ = t_3__175_ | t_3__183_;
  assign t_4__174_ = t_3__174_ | t_3__182_;
  assign t_4__173_ = t_3__173_ | t_3__181_;
  assign t_4__172_ = t_3__172_ | t_3__180_;
  assign t_4__171_ = t_3__171_ | t_3__179_;
  assign t_4__170_ = t_3__170_ | t_3__178_;
  assign t_4__169_ = t_3__169_ | t_3__177_;
  assign t_4__168_ = t_3__168_ | t_3__176_;
  assign t_4__167_ = t_3__167_ | t_3__175_;
  assign t_4__166_ = t_3__166_ | t_3__174_;
  assign t_4__165_ = t_3__165_ | t_3__173_;
  assign t_4__164_ = t_3__164_ | t_3__172_;
  assign t_4__163_ = t_3__163_ | t_3__171_;
  assign t_4__162_ = t_3__162_ | t_3__170_;
  assign t_4__161_ = t_3__161_ | t_3__169_;
  assign t_4__160_ = t_3__160_ | t_3__168_;
  assign t_4__159_ = t_3__159_ | t_3__167_;
  assign t_4__158_ = t_3__158_ | t_3__166_;
  assign t_4__157_ = t_3__157_ | t_3__165_;
  assign t_4__156_ = t_3__156_ | t_3__164_;
  assign t_4__155_ = t_3__155_ | t_3__163_;
  assign t_4__154_ = t_3__154_ | t_3__162_;
  assign t_4__153_ = t_3__153_ | t_3__161_;
  assign t_4__152_ = t_3__152_ | t_3__160_;
  assign t_4__151_ = t_3__151_ | t_3__159_;
  assign t_4__150_ = t_3__150_ | t_3__158_;
  assign t_4__149_ = t_3__149_ | t_3__157_;
  assign t_4__148_ = t_3__148_ | t_3__156_;
  assign t_4__147_ = t_3__147_ | t_3__155_;
  assign t_4__146_ = t_3__146_ | t_3__154_;
  assign t_4__145_ = t_3__145_ | t_3__153_;
  assign t_4__144_ = t_3__144_ | t_3__152_;
  assign t_4__143_ = t_3__143_ | t_3__151_;
  assign t_4__142_ = t_3__142_ | t_3__150_;
  assign t_4__141_ = t_3__141_ | t_3__149_;
  assign t_4__140_ = t_3__140_ | t_3__148_;
  assign t_4__139_ = t_3__139_ | t_3__147_;
  assign t_4__138_ = t_3__138_ | t_3__146_;
  assign t_4__137_ = t_3__137_ | t_3__145_;
  assign t_4__136_ = t_3__136_ | t_3__144_;
  assign t_4__135_ = t_3__135_ | t_3__143_;
  assign t_4__134_ = t_3__134_ | t_3__142_;
  assign t_4__133_ = t_3__133_ | t_3__141_;
  assign t_4__132_ = t_3__132_ | t_3__140_;
  assign t_4__131_ = t_3__131_ | t_3__139_;
  assign t_4__130_ = t_3__130_ | t_3__138_;
  assign t_4__129_ = t_3__129_ | t_3__137_;
  assign t_4__128_ = t_3__128_ | t_3__136_;
  assign t_4__127_ = t_3__127_ | t_3__135_;
  assign t_4__126_ = t_3__126_ | t_3__134_;
  assign t_4__125_ = t_3__125_ | t_3__133_;
  assign t_4__124_ = t_3__124_ | t_3__132_;
  assign t_4__123_ = t_3__123_ | t_3__131_;
  assign t_4__122_ = t_3__122_ | t_3__130_;
  assign t_4__121_ = t_3__121_ | t_3__129_;
  assign t_4__120_ = t_3__120_ | t_3__128_;
  assign t_4__119_ = t_3__119_ | t_3__127_;
  assign t_4__118_ = t_3__118_ | t_3__126_;
  assign t_4__117_ = t_3__117_ | t_3__125_;
  assign t_4__116_ = t_3__116_ | t_3__124_;
  assign t_4__115_ = t_3__115_ | t_3__123_;
  assign t_4__114_ = t_3__114_ | t_3__122_;
  assign t_4__113_ = t_3__113_ | t_3__121_;
  assign t_4__112_ = t_3__112_ | t_3__120_;
  assign t_4__111_ = t_3__111_ | t_3__119_;
  assign t_4__110_ = t_3__110_ | t_3__118_;
  assign t_4__109_ = t_3__109_ | t_3__117_;
  assign t_4__108_ = t_3__108_ | t_3__116_;
  assign t_4__107_ = t_3__107_ | t_3__115_;
  assign t_4__106_ = t_3__106_ | t_3__114_;
  assign t_4__105_ = t_3__105_ | t_3__113_;
  assign t_4__104_ = t_3__104_ | t_3__112_;
  assign t_4__103_ = t_3__103_ | t_3__111_;
  assign t_4__102_ = t_3__102_ | t_3__110_;
  assign t_4__101_ = t_3__101_ | t_3__109_;
  assign t_4__100_ = t_3__100_ | t_3__108_;
  assign t_4__99_ = t_3__99_ | t_3__107_;
  assign t_4__98_ = t_3__98_ | t_3__106_;
  assign t_4__97_ = t_3__97_ | t_3__105_;
  assign t_4__96_ = t_3__96_ | t_3__104_;
  assign t_4__95_ = t_3__95_ | t_3__103_;
  assign t_4__94_ = t_3__94_ | t_3__102_;
  assign t_4__93_ = t_3__93_ | t_3__101_;
  assign t_4__92_ = t_3__92_ | t_3__100_;
  assign t_4__91_ = t_3__91_ | t_3__99_;
  assign t_4__90_ = t_3__90_ | t_3__98_;
  assign t_4__89_ = t_3__89_ | t_3__97_;
  assign t_4__88_ = t_3__88_ | t_3__96_;
  assign t_4__87_ = t_3__87_ | t_3__95_;
  assign t_4__86_ = t_3__86_ | t_3__94_;
  assign t_4__85_ = t_3__85_ | t_3__93_;
  assign t_4__84_ = t_3__84_ | t_3__92_;
  assign t_4__83_ = t_3__83_ | t_3__91_;
  assign t_4__82_ = t_3__82_ | t_3__90_;
  assign t_4__81_ = t_3__81_ | t_3__89_;
  assign t_4__80_ = t_3__80_ | t_3__88_;
  assign t_4__79_ = t_3__79_ | t_3__87_;
  assign t_4__78_ = t_3__78_ | t_3__86_;
  assign t_4__77_ = t_3__77_ | t_3__85_;
  assign t_4__76_ = t_3__76_ | t_3__84_;
  assign t_4__75_ = t_3__75_ | t_3__83_;
  assign t_4__74_ = t_3__74_ | t_3__82_;
  assign t_4__73_ = t_3__73_ | t_3__81_;
  assign t_4__72_ = t_3__72_ | t_3__80_;
  assign t_4__71_ = t_3__71_ | t_3__79_;
  assign t_4__70_ = t_3__70_ | t_3__78_;
  assign t_4__69_ = t_3__69_ | t_3__77_;
  assign t_4__68_ = t_3__68_ | t_3__76_;
  assign t_4__67_ = t_3__67_ | t_3__75_;
  assign t_4__66_ = t_3__66_ | t_3__74_;
  assign t_4__65_ = t_3__65_ | t_3__73_;
  assign t_4__64_ = t_3__64_ | t_3__72_;
  assign t_4__63_ = t_3__63_ | t_3__71_;
  assign t_4__62_ = t_3__62_ | t_3__70_;
  assign t_4__61_ = t_3__61_ | t_3__69_;
  assign t_4__60_ = t_3__60_ | t_3__68_;
  assign t_4__59_ = t_3__59_ | t_3__67_;
  assign t_4__58_ = t_3__58_ | t_3__66_;
  assign t_4__57_ = t_3__57_ | t_3__65_;
  assign t_4__56_ = t_3__56_ | t_3__64_;
  assign t_4__55_ = t_3__55_ | t_3__63_;
  assign t_4__54_ = t_3__54_ | t_3__62_;
  assign t_4__53_ = t_3__53_ | t_3__61_;
  assign t_4__52_ = t_3__52_ | t_3__60_;
  assign t_4__51_ = t_3__51_ | t_3__59_;
  assign t_4__50_ = t_3__50_ | t_3__58_;
  assign t_4__49_ = t_3__49_ | t_3__57_;
  assign t_4__48_ = t_3__48_ | t_3__56_;
  assign t_4__47_ = t_3__47_ | t_3__55_;
  assign t_4__46_ = t_3__46_ | t_3__54_;
  assign t_4__45_ = t_3__45_ | t_3__53_;
  assign t_4__44_ = t_3__44_ | t_3__52_;
  assign t_4__43_ = t_3__43_ | t_3__51_;
  assign t_4__42_ = t_3__42_ | t_3__50_;
  assign t_4__41_ = t_3__41_ | t_3__49_;
  assign t_4__40_ = t_3__40_ | t_3__48_;
  assign t_4__39_ = t_3__39_ | t_3__47_;
  assign t_4__38_ = t_3__38_ | t_3__46_;
  assign t_4__37_ = t_3__37_ | t_3__45_;
  assign t_4__36_ = t_3__36_ | t_3__44_;
  assign t_4__35_ = t_3__35_ | t_3__43_;
  assign t_4__34_ = t_3__34_ | t_3__42_;
  assign t_4__33_ = t_3__33_ | t_3__41_;
  assign t_4__32_ = t_3__32_ | t_3__40_;
  assign t_4__31_ = t_3__31_ | t_3__39_;
  assign t_4__30_ = t_3__30_ | t_3__38_;
  assign t_4__29_ = t_3__29_ | t_3__37_;
  assign t_4__28_ = t_3__28_ | t_3__36_;
  assign t_4__27_ = t_3__27_ | t_3__35_;
  assign t_4__26_ = t_3__26_ | t_3__34_;
  assign t_4__25_ = t_3__25_ | t_3__33_;
  assign t_4__24_ = t_3__24_ | t_3__32_;
  assign t_4__23_ = t_3__23_ | t_3__31_;
  assign t_4__22_ = t_3__22_ | t_3__30_;
  assign t_4__21_ = t_3__21_ | t_3__29_;
  assign t_4__20_ = t_3__20_ | t_3__28_;
  assign t_4__19_ = t_3__19_ | t_3__27_;
  assign t_4__18_ = t_3__18_ | t_3__26_;
  assign t_4__17_ = t_3__17_ | t_3__25_;
  assign t_4__16_ = t_3__16_ | t_3__24_;
  assign t_4__15_ = t_3__15_ | t_3__23_;
  assign t_4__14_ = t_3__14_ | t_3__22_;
  assign t_4__13_ = t_3__13_ | t_3__21_;
  assign t_4__12_ = t_3__12_ | t_3__20_;
  assign t_4__11_ = t_3__11_ | t_3__19_;
  assign t_4__10_ = t_3__10_ | t_3__18_;
  assign t_4__9_ = t_3__9_ | t_3__17_;
  assign t_4__8_ = t_3__8_ | t_3__16_;
  assign t_4__7_ = t_3__7_ | t_3__15_;
  assign t_4__6_ = t_3__6_ | t_3__14_;
  assign t_4__5_ = t_3__5_ | t_3__13_;
  assign t_4__4_ = t_3__4_ | t_3__12_;
  assign t_4__3_ = t_3__3_ | t_3__11_;
  assign t_4__2_ = t_3__2_ | t_3__10_;
  assign t_4__1_ = t_3__1_ | t_3__9_;
  assign t_4__0_ = t_3__0_ | t_3__8_;
  assign t_5__1023_ = t_4__1023_ | 1'b0;
  assign t_5__1022_ = t_4__1022_ | 1'b0;
  assign t_5__1021_ = t_4__1021_ | 1'b0;
  assign t_5__1020_ = t_4__1020_ | 1'b0;
  assign t_5__1019_ = t_4__1019_ | 1'b0;
  assign t_5__1018_ = t_4__1018_ | 1'b0;
  assign t_5__1017_ = t_4__1017_ | 1'b0;
  assign t_5__1016_ = t_4__1016_ | 1'b0;
  assign t_5__1015_ = t_4__1015_ | 1'b0;
  assign t_5__1014_ = t_4__1014_ | 1'b0;
  assign t_5__1013_ = t_4__1013_ | 1'b0;
  assign t_5__1012_ = t_4__1012_ | 1'b0;
  assign t_5__1011_ = t_4__1011_ | 1'b0;
  assign t_5__1010_ = t_4__1010_ | 1'b0;
  assign t_5__1009_ = t_4__1009_ | 1'b0;
  assign t_5__1008_ = t_4__1008_ | 1'b0;
  assign t_5__1007_ = t_4__1007_ | t_4__1023_;
  assign t_5__1006_ = t_4__1006_ | t_4__1022_;
  assign t_5__1005_ = t_4__1005_ | t_4__1021_;
  assign t_5__1004_ = t_4__1004_ | t_4__1020_;
  assign t_5__1003_ = t_4__1003_ | t_4__1019_;
  assign t_5__1002_ = t_4__1002_ | t_4__1018_;
  assign t_5__1001_ = t_4__1001_ | t_4__1017_;
  assign t_5__1000_ = t_4__1000_ | t_4__1016_;
  assign t_5__999_ = t_4__999_ | t_4__1015_;
  assign t_5__998_ = t_4__998_ | t_4__1014_;
  assign t_5__997_ = t_4__997_ | t_4__1013_;
  assign t_5__996_ = t_4__996_ | t_4__1012_;
  assign t_5__995_ = t_4__995_ | t_4__1011_;
  assign t_5__994_ = t_4__994_ | t_4__1010_;
  assign t_5__993_ = t_4__993_ | t_4__1009_;
  assign t_5__992_ = t_4__992_ | t_4__1008_;
  assign t_5__991_ = t_4__991_ | t_4__1007_;
  assign t_5__990_ = t_4__990_ | t_4__1006_;
  assign t_5__989_ = t_4__989_ | t_4__1005_;
  assign t_5__988_ = t_4__988_ | t_4__1004_;
  assign t_5__987_ = t_4__987_ | t_4__1003_;
  assign t_5__986_ = t_4__986_ | t_4__1002_;
  assign t_5__985_ = t_4__985_ | t_4__1001_;
  assign t_5__984_ = t_4__984_ | t_4__1000_;
  assign t_5__983_ = t_4__983_ | t_4__999_;
  assign t_5__982_ = t_4__982_ | t_4__998_;
  assign t_5__981_ = t_4__981_ | t_4__997_;
  assign t_5__980_ = t_4__980_ | t_4__996_;
  assign t_5__979_ = t_4__979_ | t_4__995_;
  assign t_5__978_ = t_4__978_ | t_4__994_;
  assign t_5__977_ = t_4__977_ | t_4__993_;
  assign t_5__976_ = t_4__976_ | t_4__992_;
  assign t_5__975_ = t_4__975_ | t_4__991_;
  assign t_5__974_ = t_4__974_ | t_4__990_;
  assign t_5__973_ = t_4__973_ | t_4__989_;
  assign t_5__972_ = t_4__972_ | t_4__988_;
  assign t_5__971_ = t_4__971_ | t_4__987_;
  assign t_5__970_ = t_4__970_ | t_4__986_;
  assign t_5__969_ = t_4__969_ | t_4__985_;
  assign t_5__968_ = t_4__968_ | t_4__984_;
  assign t_5__967_ = t_4__967_ | t_4__983_;
  assign t_5__966_ = t_4__966_ | t_4__982_;
  assign t_5__965_ = t_4__965_ | t_4__981_;
  assign t_5__964_ = t_4__964_ | t_4__980_;
  assign t_5__963_ = t_4__963_ | t_4__979_;
  assign t_5__962_ = t_4__962_ | t_4__978_;
  assign t_5__961_ = t_4__961_ | t_4__977_;
  assign t_5__960_ = t_4__960_ | t_4__976_;
  assign t_5__959_ = t_4__959_ | t_4__975_;
  assign t_5__958_ = t_4__958_ | t_4__974_;
  assign t_5__957_ = t_4__957_ | t_4__973_;
  assign t_5__956_ = t_4__956_ | t_4__972_;
  assign t_5__955_ = t_4__955_ | t_4__971_;
  assign t_5__954_ = t_4__954_ | t_4__970_;
  assign t_5__953_ = t_4__953_ | t_4__969_;
  assign t_5__952_ = t_4__952_ | t_4__968_;
  assign t_5__951_ = t_4__951_ | t_4__967_;
  assign t_5__950_ = t_4__950_ | t_4__966_;
  assign t_5__949_ = t_4__949_ | t_4__965_;
  assign t_5__948_ = t_4__948_ | t_4__964_;
  assign t_5__947_ = t_4__947_ | t_4__963_;
  assign t_5__946_ = t_4__946_ | t_4__962_;
  assign t_5__945_ = t_4__945_ | t_4__961_;
  assign t_5__944_ = t_4__944_ | t_4__960_;
  assign t_5__943_ = t_4__943_ | t_4__959_;
  assign t_5__942_ = t_4__942_ | t_4__958_;
  assign t_5__941_ = t_4__941_ | t_4__957_;
  assign t_5__940_ = t_4__940_ | t_4__956_;
  assign t_5__939_ = t_4__939_ | t_4__955_;
  assign t_5__938_ = t_4__938_ | t_4__954_;
  assign t_5__937_ = t_4__937_ | t_4__953_;
  assign t_5__936_ = t_4__936_ | t_4__952_;
  assign t_5__935_ = t_4__935_ | t_4__951_;
  assign t_5__934_ = t_4__934_ | t_4__950_;
  assign t_5__933_ = t_4__933_ | t_4__949_;
  assign t_5__932_ = t_4__932_ | t_4__948_;
  assign t_5__931_ = t_4__931_ | t_4__947_;
  assign t_5__930_ = t_4__930_ | t_4__946_;
  assign t_5__929_ = t_4__929_ | t_4__945_;
  assign t_5__928_ = t_4__928_ | t_4__944_;
  assign t_5__927_ = t_4__927_ | t_4__943_;
  assign t_5__926_ = t_4__926_ | t_4__942_;
  assign t_5__925_ = t_4__925_ | t_4__941_;
  assign t_5__924_ = t_4__924_ | t_4__940_;
  assign t_5__923_ = t_4__923_ | t_4__939_;
  assign t_5__922_ = t_4__922_ | t_4__938_;
  assign t_5__921_ = t_4__921_ | t_4__937_;
  assign t_5__920_ = t_4__920_ | t_4__936_;
  assign t_5__919_ = t_4__919_ | t_4__935_;
  assign t_5__918_ = t_4__918_ | t_4__934_;
  assign t_5__917_ = t_4__917_ | t_4__933_;
  assign t_5__916_ = t_4__916_ | t_4__932_;
  assign t_5__915_ = t_4__915_ | t_4__931_;
  assign t_5__914_ = t_4__914_ | t_4__930_;
  assign t_5__913_ = t_4__913_ | t_4__929_;
  assign t_5__912_ = t_4__912_ | t_4__928_;
  assign t_5__911_ = t_4__911_ | t_4__927_;
  assign t_5__910_ = t_4__910_ | t_4__926_;
  assign t_5__909_ = t_4__909_ | t_4__925_;
  assign t_5__908_ = t_4__908_ | t_4__924_;
  assign t_5__907_ = t_4__907_ | t_4__923_;
  assign t_5__906_ = t_4__906_ | t_4__922_;
  assign t_5__905_ = t_4__905_ | t_4__921_;
  assign t_5__904_ = t_4__904_ | t_4__920_;
  assign t_5__903_ = t_4__903_ | t_4__919_;
  assign t_5__902_ = t_4__902_ | t_4__918_;
  assign t_5__901_ = t_4__901_ | t_4__917_;
  assign t_5__900_ = t_4__900_ | t_4__916_;
  assign t_5__899_ = t_4__899_ | t_4__915_;
  assign t_5__898_ = t_4__898_ | t_4__914_;
  assign t_5__897_ = t_4__897_ | t_4__913_;
  assign t_5__896_ = t_4__896_ | t_4__912_;
  assign t_5__895_ = t_4__895_ | t_4__911_;
  assign t_5__894_ = t_4__894_ | t_4__910_;
  assign t_5__893_ = t_4__893_ | t_4__909_;
  assign t_5__892_ = t_4__892_ | t_4__908_;
  assign t_5__891_ = t_4__891_ | t_4__907_;
  assign t_5__890_ = t_4__890_ | t_4__906_;
  assign t_5__889_ = t_4__889_ | t_4__905_;
  assign t_5__888_ = t_4__888_ | t_4__904_;
  assign t_5__887_ = t_4__887_ | t_4__903_;
  assign t_5__886_ = t_4__886_ | t_4__902_;
  assign t_5__885_ = t_4__885_ | t_4__901_;
  assign t_5__884_ = t_4__884_ | t_4__900_;
  assign t_5__883_ = t_4__883_ | t_4__899_;
  assign t_5__882_ = t_4__882_ | t_4__898_;
  assign t_5__881_ = t_4__881_ | t_4__897_;
  assign t_5__880_ = t_4__880_ | t_4__896_;
  assign t_5__879_ = t_4__879_ | t_4__895_;
  assign t_5__878_ = t_4__878_ | t_4__894_;
  assign t_5__877_ = t_4__877_ | t_4__893_;
  assign t_5__876_ = t_4__876_ | t_4__892_;
  assign t_5__875_ = t_4__875_ | t_4__891_;
  assign t_5__874_ = t_4__874_ | t_4__890_;
  assign t_5__873_ = t_4__873_ | t_4__889_;
  assign t_5__872_ = t_4__872_ | t_4__888_;
  assign t_5__871_ = t_4__871_ | t_4__887_;
  assign t_5__870_ = t_4__870_ | t_4__886_;
  assign t_5__869_ = t_4__869_ | t_4__885_;
  assign t_5__868_ = t_4__868_ | t_4__884_;
  assign t_5__867_ = t_4__867_ | t_4__883_;
  assign t_5__866_ = t_4__866_ | t_4__882_;
  assign t_5__865_ = t_4__865_ | t_4__881_;
  assign t_5__864_ = t_4__864_ | t_4__880_;
  assign t_5__863_ = t_4__863_ | t_4__879_;
  assign t_5__862_ = t_4__862_ | t_4__878_;
  assign t_5__861_ = t_4__861_ | t_4__877_;
  assign t_5__860_ = t_4__860_ | t_4__876_;
  assign t_5__859_ = t_4__859_ | t_4__875_;
  assign t_5__858_ = t_4__858_ | t_4__874_;
  assign t_5__857_ = t_4__857_ | t_4__873_;
  assign t_5__856_ = t_4__856_ | t_4__872_;
  assign t_5__855_ = t_4__855_ | t_4__871_;
  assign t_5__854_ = t_4__854_ | t_4__870_;
  assign t_5__853_ = t_4__853_ | t_4__869_;
  assign t_5__852_ = t_4__852_ | t_4__868_;
  assign t_5__851_ = t_4__851_ | t_4__867_;
  assign t_5__850_ = t_4__850_ | t_4__866_;
  assign t_5__849_ = t_4__849_ | t_4__865_;
  assign t_5__848_ = t_4__848_ | t_4__864_;
  assign t_5__847_ = t_4__847_ | t_4__863_;
  assign t_5__846_ = t_4__846_ | t_4__862_;
  assign t_5__845_ = t_4__845_ | t_4__861_;
  assign t_5__844_ = t_4__844_ | t_4__860_;
  assign t_5__843_ = t_4__843_ | t_4__859_;
  assign t_5__842_ = t_4__842_ | t_4__858_;
  assign t_5__841_ = t_4__841_ | t_4__857_;
  assign t_5__840_ = t_4__840_ | t_4__856_;
  assign t_5__839_ = t_4__839_ | t_4__855_;
  assign t_5__838_ = t_4__838_ | t_4__854_;
  assign t_5__837_ = t_4__837_ | t_4__853_;
  assign t_5__836_ = t_4__836_ | t_4__852_;
  assign t_5__835_ = t_4__835_ | t_4__851_;
  assign t_5__834_ = t_4__834_ | t_4__850_;
  assign t_5__833_ = t_4__833_ | t_4__849_;
  assign t_5__832_ = t_4__832_ | t_4__848_;
  assign t_5__831_ = t_4__831_ | t_4__847_;
  assign t_5__830_ = t_4__830_ | t_4__846_;
  assign t_5__829_ = t_4__829_ | t_4__845_;
  assign t_5__828_ = t_4__828_ | t_4__844_;
  assign t_5__827_ = t_4__827_ | t_4__843_;
  assign t_5__826_ = t_4__826_ | t_4__842_;
  assign t_5__825_ = t_4__825_ | t_4__841_;
  assign t_5__824_ = t_4__824_ | t_4__840_;
  assign t_5__823_ = t_4__823_ | t_4__839_;
  assign t_5__822_ = t_4__822_ | t_4__838_;
  assign t_5__821_ = t_4__821_ | t_4__837_;
  assign t_5__820_ = t_4__820_ | t_4__836_;
  assign t_5__819_ = t_4__819_ | t_4__835_;
  assign t_5__818_ = t_4__818_ | t_4__834_;
  assign t_5__817_ = t_4__817_ | t_4__833_;
  assign t_5__816_ = t_4__816_ | t_4__832_;
  assign t_5__815_ = t_4__815_ | t_4__831_;
  assign t_5__814_ = t_4__814_ | t_4__830_;
  assign t_5__813_ = t_4__813_ | t_4__829_;
  assign t_5__812_ = t_4__812_ | t_4__828_;
  assign t_5__811_ = t_4__811_ | t_4__827_;
  assign t_5__810_ = t_4__810_ | t_4__826_;
  assign t_5__809_ = t_4__809_ | t_4__825_;
  assign t_5__808_ = t_4__808_ | t_4__824_;
  assign t_5__807_ = t_4__807_ | t_4__823_;
  assign t_5__806_ = t_4__806_ | t_4__822_;
  assign t_5__805_ = t_4__805_ | t_4__821_;
  assign t_5__804_ = t_4__804_ | t_4__820_;
  assign t_5__803_ = t_4__803_ | t_4__819_;
  assign t_5__802_ = t_4__802_ | t_4__818_;
  assign t_5__801_ = t_4__801_ | t_4__817_;
  assign t_5__800_ = t_4__800_ | t_4__816_;
  assign t_5__799_ = t_4__799_ | t_4__815_;
  assign t_5__798_ = t_4__798_ | t_4__814_;
  assign t_5__797_ = t_4__797_ | t_4__813_;
  assign t_5__796_ = t_4__796_ | t_4__812_;
  assign t_5__795_ = t_4__795_ | t_4__811_;
  assign t_5__794_ = t_4__794_ | t_4__810_;
  assign t_5__793_ = t_4__793_ | t_4__809_;
  assign t_5__792_ = t_4__792_ | t_4__808_;
  assign t_5__791_ = t_4__791_ | t_4__807_;
  assign t_5__790_ = t_4__790_ | t_4__806_;
  assign t_5__789_ = t_4__789_ | t_4__805_;
  assign t_5__788_ = t_4__788_ | t_4__804_;
  assign t_5__787_ = t_4__787_ | t_4__803_;
  assign t_5__786_ = t_4__786_ | t_4__802_;
  assign t_5__785_ = t_4__785_ | t_4__801_;
  assign t_5__784_ = t_4__784_ | t_4__800_;
  assign t_5__783_ = t_4__783_ | t_4__799_;
  assign t_5__782_ = t_4__782_ | t_4__798_;
  assign t_5__781_ = t_4__781_ | t_4__797_;
  assign t_5__780_ = t_4__780_ | t_4__796_;
  assign t_5__779_ = t_4__779_ | t_4__795_;
  assign t_5__778_ = t_4__778_ | t_4__794_;
  assign t_5__777_ = t_4__777_ | t_4__793_;
  assign t_5__776_ = t_4__776_ | t_4__792_;
  assign t_5__775_ = t_4__775_ | t_4__791_;
  assign t_5__774_ = t_4__774_ | t_4__790_;
  assign t_5__773_ = t_4__773_ | t_4__789_;
  assign t_5__772_ = t_4__772_ | t_4__788_;
  assign t_5__771_ = t_4__771_ | t_4__787_;
  assign t_5__770_ = t_4__770_ | t_4__786_;
  assign t_5__769_ = t_4__769_ | t_4__785_;
  assign t_5__768_ = t_4__768_ | t_4__784_;
  assign t_5__767_ = t_4__767_ | t_4__783_;
  assign t_5__766_ = t_4__766_ | t_4__782_;
  assign t_5__765_ = t_4__765_ | t_4__781_;
  assign t_5__764_ = t_4__764_ | t_4__780_;
  assign t_5__763_ = t_4__763_ | t_4__779_;
  assign t_5__762_ = t_4__762_ | t_4__778_;
  assign t_5__761_ = t_4__761_ | t_4__777_;
  assign t_5__760_ = t_4__760_ | t_4__776_;
  assign t_5__759_ = t_4__759_ | t_4__775_;
  assign t_5__758_ = t_4__758_ | t_4__774_;
  assign t_5__757_ = t_4__757_ | t_4__773_;
  assign t_5__756_ = t_4__756_ | t_4__772_;
  assign t_5__755_ = t_4__755_ | t_4__771_;
  assign t_5__754_ = t_4__754_ | t_4__770_;
  assign t_5__753_ = t_4__753_ | t_4__769_;
  assign t_5__752_ = t_4__752_ | t_4__768_;
  assign t_5__751_ = t_4__751_ | t_4__767_;
  assign t_5__750_ = t_4__750_ | t_4__766_;
  assign t_5__749_ = t_4__749_ | t_4__765_;
  assign t_5__748_ = t_4__748_ | t_4__764_;
  assign t_5__747_ = t_4__747_ | t_4__763_;
  assign t_5__746_ = t_4__746_ | t_4__762_;
  assign t_5__745_ = t_4__745_ | t_4__761_;
  assign t_5__744_ = t_4__744_ | t_4__760_;
  assign t_5__743_ = t_4__743_ | t_4__759_;
  assign t_5__742_ = t_4__742_ | t_4__758_;
  assign t_5__741_ = t_4__741_ | t_4__757_;
  assign t_5__740_ = t_4__740_ | t_4__756_;
  assign t_5__739_ = t_4__739_ | t_4__755_;
  assign t_5__738_ = t_4__738_ | t_4__754_;
  assign t_5__737_ = t_4__737_ | t_4__753_;
  assign t_5__736_ = t_4__736_ | t_4__752_;
  assign t_5__735_ = t_4__735_ | t_4__751_;
  assign t_5__734_ = t_4__734_ | t_4__750_;
  assign t_5__733_ = t_4__733_ | t_4__749_;
  assign t_5__732_ = t_4__732_ | t_4__748_;
  assign t_5__731_ = t_4__731_ | t_4__747_;
  assign t_5__730_ = t_4__730_ | t_4__746_;
  assign t_5__729_ = t_4__729_ | t_4__745_;
  assign t_5__728_ = t_4__728_ | t_4__744_;
  assign t_5__727_ = t_4__727_ | t_4__743_;
  assign t_5__726_ = t_4__726_ | t_4__742_;
  assign t_5__725_ = t_4__725_ | t_4__741_;
  assign t_5__724_ = t_4__724_ | t_4__740_;
  assign t_5__723_ = t_4__723_ | t_4__739_;
  assign t_5__722_ = t_4__722_ | t_4__738_;
  assign t_5__721_ = t_4__721_ | t_4__737_;
  assign t_5__720_ = t_4__720_ | t_4__736_;
  assign t_5__719_ = t_4__719_ | t_4__735_;
  assign t_5__718_ = t_4__718_ | t_4__734_;
  assign t_5__717_ = t_4__717_ | t_4__733_;
  assign t_5__716_ = t_4__716_ | t_4__732_;
  assign t_5__715_ = t_4__715_ | t_4__731_;
  assign t_5__714_ = t_4__714_ | t_4__730_;
  assign t_5__713_ = t_4__713_ | t_4__729_;
  assign t_5__712_ = t_4__712_ | t_4__728_;
  assign t_5__711_ = t_4__711_ | t_4__727_;
  assign t_5__710_ = t_4__710_ | t_4__726_;
  assign t_5__709_ = t_4__709_ | t_4__725_;
  assign t_5__708_ = t_4__708_ | t_4__724_;
  assign t_5__707_ = t_4__707_ | t_4__723_;
  assign t_5__706_ = t_4__706_ | t_4__722_;
  assign t_5__705_ = t_4__705_ | t_4__721_;
  assign t_5__704_ = t_4__704_ | t_4__720_;
  assign t_5__703_ = t_4__703_ | t_4__719_;
  assign t_5__702_ = t_4__702_ | t_4__718_;
  assign t_5__701_ = t_4__701_ | t_4__717_;
  assign t_5__700_ = t_4__700_ | t_4__716_;
  assign t_5__699_ = t_4__699_ | t_4__715_;
  assign t_5__698_ = t_4__698_ | t_4__714_;
  assign t_5__697_ = t_4__697_ | t_4__713_;
  assign t_5__696_ = t_4__696_ | t_4__712_;
  assign t_5__695_ = t_4__695_ | t_4__711_;
  assign t_5__694_ = t_4__694_ | t_4__710_;
  assign t_5__693_ = t_4__693_ | t_4__709_;
  assign t_5__692_ = t_4__692_ | t_4__708_;
  assign t_5__691_ = t_4__691_ | t_4__707_;
  assign t_5__690_ = t_4__690_ | t_4__706_;
  assign t_5__689_ = t_4__689_ | t_4__705_;
  assign t_5__688_ = t_4__688_ | t_4__704_;
  assign t_5__687_ = t_4__687_ | t_4__703_;
  assign t_5__686_ = t_4__686_ | t_4__702_;
  assign t_5__685_ = t_4__685_ | t_4__701_;
  assign t_5__684_ = t_4__684_ | t_4__700_;
  assign t_5__683_ = t_4__683_ | t_4__699_;
  assign t_5__682_ = t_4__682_ | t_4__698_;
  assign t_5__681_ = t_4__681_ | t_4__697_;
  assign t_5__680_ = t_4__680_ | t_4__696_;
  assign t_5__679_ = t_4__679_ | t_4__695_;
  assign t_5__678_ = t_4__678_ | t_4__694_;
  assign t_5__677_ = t_4__677_ | t_4__693_;
  assign t_5__676_ = t_4__676_ | t_4__692_;
  assign t_5__675_ = t_4__675_ | t_4__691_;
  assign t_5__674_ = t_4__674_ | t_4__690_;
  assign t_5__673_ = t_4__673_ | t_4__689_;
  assign t_5__672_ = t_4__672_ | t_4__688_;
  assign t_5__671_ = t_4__671_ | t_4__687_;
  assign t_5__670_ = t_4__670_ | t_4__686_;
  assign t_5__669_ = t_4__669_ | t_4__685_;
  assign t_5__668_ = t_4__668_ | t_4__684_;
  assign t_5__667_ = t_4__667_ | t_4__683_;
  assign t_5__666_ = t_4__666_ | t_4__682_;
  assign t_5__665_ = t_4__665_ | t_4__681_;
  assign t_5__664_ = t_4__664_ | t_4__680_;
  assign t_5__663_ = t_4__663_ | t_4__679_;
  assign t_5__662_ = t_4__662_ | t_4__678_;
  assign t_5__661_ = t_4__661_ | t_4__677_;
  assign t_5__660_ = t_4__660_ | t_4__676_;
  assign t_5__659_ = t_4__659_ | t_4__675_;
  assign t_5__658_ = t_4__658_ | t_4__674_;
  assign t_5__657_ = t_4__657_ | t_4__673_;
  assign t_5__656_ = t_4__656_ | t_4__672_;
  assign t_5__655_ = t_4__655_ | t_4__671_;
  assign t_5__654_ = t_4__654_ | t_4__670_;
  assign t_5__653_ = t_4__653_ | t_4__669_;
  assign t_5__652_ = t_4__652_ | t_4__668_;
  assign t_5__651_ = t_4__651_ | t_4__667_;
  assign t_5__650_ = t_4__650_ | t_4__666_;
  assign t_5__649_ = t_4__649_ | t_4__665_;
  assign t_5__648_ = t_4__648_ | t_4__664_;
  assign t_5__647_ = t_4__647_ | t_4__663_;
  assign t_5__646_ = t_4__646_ | t_4__662_;
  assign t_5__645_ = t_4__645_ | t_4__661_;
  assign t_5__644_ = t_4__644_ | t_4__660_;
  assign t_5__643_ = t_4__643_ | t_4__659_;
  assign t_5__642_ = t_4__642_ | t_4__658_;
  assign t_5__641_ = t_4__641_ | t_4__657_;
  assign t_5__640_ = t_4__640_ | t_4__656_;
  assign t_5__639_ = t_4__639_ | t_4__655_;
  assign t_5__638_ = t_4__638_ | t_4__654_;
  assign t_5__637_ = t_4__637_ | t_4__653_;
  assign t_5__636_ = t_4__636_ | t_4__652_;
  assign t_5__635_ = t_4__635_ | t_4__651_;
  assign t_5__634_ = t_4__634_ | t_4__650_;
  assign t_5__633_ = t_4__633_ | t_4__649_;
  assign t_5__632_ = t_4__632_ | t_4__648_;
  assign t_5__631_ = t_4__631_ | t_4__647_;
  assign t_5__630_ = t_4__630_ | t_4__646_;
  assign t_5__629_ = t_4__629_ | t_4__645_;
  assign t_5__628_ = t_4__628_ | t_4__644_;
  assign t_5__627_ = t_4__627_ | t_4__643_;
  assign t_5__626_ = t_4__626_ | t_4__642_;
  assign t_5__625_ = t_4__625_ | t_4__641_;
  assign t_5__624_ = t_4__624_ | t_4__640_;
  assign t_5__623_ = t_4__623_ | t_4__639_;
  assign t_5__622_ = t_4__622_ | t_4__638_;
  assign t_5__621_ = t_4__621_ | t_4__637_;
  assign t_5__620_ = t_4__620_ | t_4__636_;
  assign t_5__619_ = t_4__619_ | t_4__635_;
  assign t_5__618_ = t_4__618_ | t_4__634_;
  assign t_5__617_ = t_4__617_ | t_4__633_;
  assign t_5__616_ = t_4__616_ | t_4__632_;
  assign t_5__615_ = t_4__615_ | t_4__631_;
  assign t_5__614_ = t_4__614_ | t_4__630_;
  assign t_5__613_ = t_4__613_ | t_4__629_;
  assign t_5__612_ = t_4__612_ | t_4__628_;
  assign t_5__611_ = t_4__611_ | t_4__627_;
  assign t_5__610_ = t_4__610_ | t_4__626_;
  assign t_5__609_ = t_4__609_ | t_4__625_;
  assign t_5__608_ = t_4__608_ | t_4__624_;
  assign t_5__607_ = t_4__607_ | t_4__623_;
  assign t_5__606_ = t_4__606_ | t_4__622_;
  assign t_5__605_ = t_4__605_ | t_4__621_;
  assign t_5__604_ = t_4__604_ | t_4__620_;
  assign t_5__603_ = t_4__603_ | t_4__619_;
  assign t_5__602_ = t_4__602_ | t_4__618_;
  assign t_5__601_ = t_4__601_ | t_4__617_;
  assign t_5__600_ = t_4__600_ | t_4__616_;
  assign t_5__599_ = t_4__599_ | t_4__615_;
  assign t_5__598_ = t_4__598_ | t_4__614_;
  assign t_5__597_ = t_4__597_ | t_4__613_;
  assign t_5__596_ = t_4__596_ | t_4__612_;
  assign t_5__595_ = t_4__595_ | t_4__611_;
  assign t_5__594_ = t_4__594_ | t_4__610_;
  assign t_5__593_ = t_4__593_ | t_4__609_;
  assign t_5__592_ = t_4__592_ | t_4__608_;
  assign t_5__591_ = t_4__591_ | t_4__607_;
  assign t_5__590_ = t_4__590_ | t_4__606_;
  assign t_5__589_ = t_4__589_ | t_4__605_;
  assign t_5__588_ = t_4__588_ | t_4__604_;
  assign t_5__587_ = t_4__587_ | t_4__603_;
  assign t_5__586_ = t_4__586_ | t_4__602_;
  assign t_5__585_ = t_4__585_ | t_4__601_;
  assign t_5__584_ = t_4__584_ | t_4__600_;
  assign t_5__583_ = t_4__583_ | t_4__599_;
  assign t_5__582_ = t_4__582_ | t_4__598_;
  assign t_5__581_ = t_4__581_ | t_4__597_;
  assign t_5__580_ = t_4__580_ | t_4__596_;
  assign t_5__579_ = t_4__579_ | t_4__595_;
  assign t_5__578_ = t_4__578_ | t_4__594_;
  assign t_5__577_ = t_4__577_ | t_4__593_;
  assign t_5__576_ = t_4__576_ | t_4__592_;
  assign t_5__575_ = t_4__575_ | t_4__591_;
  assign t_5__574_ = t_4__574_ | t_4__590_;
  assign t_5__573_ = t_4__573_ | t_4__589_;
  assign t_5__572_ = t_4__572_ | t_4__588_;
  assign t_5__571_ = t_4__571_ | t_4__587_;
  assign t_5__570_ = t_4__570_ | t_4__586_;
  assign t_5__569_ = t_4__569_ | t_4__585_;
  assign t_5__568_ = t_4__568_ | t_4__584_;
  assign t_5__567_ = t_4__567_ | t_4__583_;
  assign t_5__566_ = t_4__566_ | t_4__582_;
  assign t_5__565_ = t_4__565_ | t_4__581_;
  assign t_5__564_ = t_4__564_ | t_4__580_;
  assign t_5__563_ = t_4__563_ | t_4__579_;
  assign t_5__562_ = t_4__562_ | t_4__578_;
  assign t_5__561_ = t_4__561_ | t_4__577_;
  assign t_5__560_ = t_4__560_ | t_4__576_;
  assign t_5__559_ = t_4__559_ | t_4__575_;
  assign t_5__558_ = t_4__558_ | t_4__574_;
  assign t_5__557_ = t_4__557_ | t_4__573_;
  assign t_5__556_ = t_4__556_ | t_4__572_;
  assign t_5__555_ = t_4__555_ | t_4__571_;
  assign t_5__554_ = t_4__554_ | t_4__570_;
  assign t_5__553_ = t_4__553_ | t_4__569_;
  assign t_5__552_ = t_4__552_ | t_4__568_;
  assign t_5__551_ = t_4__551_ | t_4__567_;
  assign t_5__550_ = t_4__550_ | t_4__566_;
  assign t_5__549_ = t_4__549_ | t_4__565_;
  assign t_5__548_ = t_4__548_ | t_4__564_;
  assign t_5__547_ = t_4__547_ | t_4__563_;
  assign t_5__546_ = t_4__546_ | t_4__562_;
  assign t_5__545_ = t_4__545_ | t_4__561_;
  assign t_5__544_ = t_4__544_ | t_4__560_;
  assign t_5__543_ = t_4__543_ | t_4__559_;
  assign t_5__542_ = t_4__542_ | t_4__558_;
  assign t_5__541_ = t_4__541_ | t_4__557_;
  assign t_5__540_ = t_4__540_ | t_4__556_;
  assign t_5__539_ = t_4__539_ | t_4__555_;
  assign t_5__538_ = t_4__538_ | t_4__554_;
  assign t_5__537_ = t_4__537_ | t_4__553_;
  assign t_5__536_ = t_4__536_ | t_4__552_;
  assign t_5__535_ = t_4__535_ | t_4__551_;
  assign t_5__534_ = t_4__534_ | t_4__550_;
  assign t_5__533_ = t_4__533_ | t_4__549_;
  assign t_5__532_ = t_4__532_ | t_4__548_;
  assign t_5__531_ = t_4__531_ | t_4__547_;
  assign t_5__530_ = t_4__530_ | t_4__546_;
  assign t_5__529_ = t_4__529_ | t_4__545_;
  assign t_5__528_ = t_4__528_ | t_4__544_;
  assign t_5__527_ = t_4__527_ | t_4__543_;
  assign t_5__526_ = t_4__526_ | t_4__542_;
  assign t_5__525_ = t_4__525_ | t_4__541_;
  assign t_5__524_ = t_4__524_ | t_4__540_;
  assign t_5__523_ = t_4__523_ | t_4__539_;
  assign t_5__522_ = t_4__522_ | t_4__538_;
  assign t_5__521_ = t_4__521_ | t_4__537_;
  assign t_5__520_ = t_4__520_ | t_4__536_;
  assign t_5__519_ = t_4__519_ | t_4__535_;
  assign t_5__518_ = t_4__518_ | t_4__534_;
  assign t_5__517_ = t_4__517_ | t_4__533_;
  assign t_5__516_ = t_4__516_ | t_4__532_;
  assign t_5__515_ = t_4__515_ | t_4__531_;
  assign t_5__514_ = t_4__514_ | t_4__530_;
  assign t_5__513_ = t_4__513_ | t_4__529_;
  assign t_5__512_ = t_4__512_ | t_4__528_;
  assign t_5__511_ = t_4__511_ | t_4__527_;
  assign t_5__510_ = t_4__510_ | t_4__526_;
  assign t_5__509_ = t_4__509_ | t_4__525_;
  assign t_5__508_ = t_4__508_ | t_4__524_;
  assign t_5__507_ = t_4__507_ | t_4__523_;
  assign t_5__506_ = t_4__506_ | t_4__522_;
  assign t_5__505_ = t_4__505_ | t_4__521_;
  assign t_5__504_ = t_4__504_ | t_4__520_;
  assign t_5__503_ = t_4__503_ | t_4__519_;
  assign t_5__502_ = t_4__502_ | t_4__518_;
  assign t_5__501_ = t_4__501_ | t_4__517_;
  assign t_5__500_ = t_4__500_ | t_4__516_;
  assign t_5__499_ = t_4__499_ | t_4__515_;
  assign t_5__498_ = t_4__498_ | t_4__514_;
  assign t_5__497_ = t_4__497_ | t_4__513_;
  assign t_5__496_ = t_4__496_ | t_4__512_;
  assign t_5__495_ = t_4__495_ | t_4__511_;
  assign t_5__494_ = t_4__494_ | t_4__510_;
  assign t_5__493_ = t_4__493_ | t_4__509_;
  assign t_5__492_ = t_4__492_ | t_4__508_;
  assign t_5__491_ = t_4__491_ | t_4__507_;
  assign t_5__490_ = t_4__490_ | t_4__506_;
  assign t_5__489_ = t_4__489_ | t_4__505_;
  assign t_5__488_ = t_4__488_ | t_4__504_;
  assign t_5__487_ = t_4__487_ | t_4__503_;
  assign t_5__486_ = t_4__486_ | t_4__502_;
  assign t_5__485_ = t_4__485_ | t_4__501_;
  assign t_5__484_ = t_4__484_ | t_4__500_;
  assign t_5__483_ = t_4__483_ | t_4__499_;
  assign t_5__482_ = t_4__482_ | t_4__498_;
  assign t_5__481_ = t_4__481_ | t_4__497_;
  assign t_5__480_ = t_4__480_ | t_4__496_;
  assign t_5__479_ = t_4__479_ | t_4__495_;
  assign t_5__478_ = t_4__478_ | t_4__494_;
  assign t_5__477_ = t_4__477_ | t_4__493_;
  assign t_5__476_ = t_4__476_ | t_4__492_;
  assign t_5__475_ = t_4__475_ | t_4__491_;
  assign t_5__474_ = t_4__474_ | t_4__490_;
  assign t_5__473_ = t_4__473_ | t_4__489_;
  assign t_5__472_ = t_4__472_ | t_4__488_;
  assign t_5__471_ = t_4__471_ | t_4__487_;
  assign t_5__470_ = t_4__470_ | t_4__486_;
  assign t_5__469_ = t_4__469_ | t_4__485_;
  assign t_5__468_ = t_4__468_ | t_4__484_;
  assign t_5__467_ = t_4__467_ | t_4__483_;
  assign t_5__466_ = t_4__466_ | t_4__482_;
  assign t_5__465_ = t_4__465_ | t_4__481_;
  assign t_5__464_ = t_4__464_ | t_4__480_;
  assign t_5__463_ = t_4__463_ | t_4__479_;
  assign t_5__462_ = t_4__462_ | t_4__478_;
  assign t_5__461_ = t_4__461_ | t_4__477_;
  assign t_5__460_ = t_4__460_ | t_4__476_;
  assign t_5__459_ = t_4__459_ | t_4__475_;
  assign t_5__458_ = t_4__458_ | t_4__474_;
  assign t_5__457_ = t_4__457_ | t_4__473_;
  assign t_5__456_ = t_4__456_ | t_4__472_;
  assign t_5__455_ = t_4__455_ | t_4__471_;
  assign t_5__454_ = t_4__454_ | t_4__470_;
  assign t_5__453_ = t_4__453_ | t_4__469_;
  assign t_5__452_ = t_4__452_ | t_4__468_;
  assign t_5__451_ = t_4__451_ | t_4__467_;
  assign t_5__450_ = t_4__450_ | t_4__466_;
  assign t_5__449_ = t_4__449_ | t_4__465_;
  assign t_5__448_ = t_4__448_ | t_4__464_;
  assign t_5__447_ = t_4__447_ | t_4__463_;
  assign t_5__446_ = t_4__446_ | t_4__462_;
  assign t_5__445_ = t_4__445_ | t_4__461_;
  assign t_5__444_ = t_4__444_ | t_4__460_;
  assign t_5__443_ = t_4__443_ | t_4__459_;
  assign t_5__442_ = t_4__442_ | t_4__458_;
  assign t_5__441_ = t_4__441_ | t_4__457_;
  assign t_5__440_ = t_4__440_ | t_4__456_;
  assign t_5__439_ = t_4__439_ | t_4__455_;
  assign t_5__438_ = t_4__438_ | t_4__454_;
  assign t_5__437_ = t_4__437_ | t_4__453_;
  assign t_5__436_ = t_4__436_ | t_4__452_;
  assign t_5__435_ = t_4__435_ | t_4__451_;
  assign t_5__434_ = t_4__434_ | t_4__450_;
  assign t_5__433_ = t_4__433_ | t_4__449_;
  assign t_5__432_ = t_4__432_ | t_4__448_;
  assign t_5__431_ = t_4__431_ | t_4__447_;
  assign t_5__430_ = t_4__430_ | t_4__446_;
  assign t_5__429_ = t_4__429_ | t_4__445_;
  assign t_5__428_ = t_4__428_ | t_4__444_;
  assign t_5__427_ = t_4__427_ | t_4__443_;
  assign t_5__426_ = t_4__426_ | t_4__442_;
  assign t_5__425_ = t_4__425_ | t_4__441_;
  assign t_5__424_ = t_4__424_ | t_4__440_;
  assign t_5__423_ = t_4__423_ | t_4__439_;
  assign t_5__422_ = t_4__422_ | t_4__438_;
  assign t_5__421_ = t_4__421_ | t_4__437_;
  assign t_5__420_ = t_4__420_ | t_4__436_;
  assign t_5__419_ = t_4__419_ | t_4__435_;
  assign t_5__418_ = t_4__418_ | t_4__434_;
  assign t_5__417_ = t_4__417_ | t_4__433_;
  assign t_5__416_ = t_4__416_ | t_4__432_;
  assign t_5__415_ = t_4__415_ | t_4__431_;
  assign t_5__414_ = t_4__414_ | t_4__430_;
  assign t_5__413_ = t_4__413_ | t_4__429_;
  assign t_5__412_ = t_4__412_ | t_4__428_;
  assign t_5__411_ = t_4__411_ | t_4__427_;
  assign t_5__410_ = t_4__410_ | t_4__426_;
  assign t_5__409_ = t_4__409_ | t_4__425_;
  assign t_5__408_ = t_4__408_ | t_4__424_;
  assign t_5__407_ = t_4__407_ | t_4__423_;
  assign t_5__406_ = t_4__406_ | t_4__422_;
  assign t_5__405_ = t_4__405_ | t_4__421_;
  assign t_5__404_ = t_4__404_ | t_4__420_;
  assign t_5__403_ = t_4__403_ | t_4__419_;
  assign t_5__402_ = t_4__402_ | t_4__418_;
  assign t_5__401_ = t_4__401_ | t_4__417_;
  assign t_5__400_ = t_4__400_ | t_4__416_;
  assign t_5__399_ = t_4__399_ | t_4__415_;
  assign t_5__398_ = t_4__398_ | t_4__414_;
  assign t_5__397_ = t_4__397_ | t_4__413_;
  assign t_5__396_ = t_4__396_ | t_4__412_;
  assign t_5__395_ = t_4__395_ | t_4__411_;
  assign t_5__394_ = t_4__394_ | t_4__410_;
  assign t_5__393_ = t_4__393_ | t_4__409_;
  assign t_5__392_ = t_4__392_ | t_4__408_;
  assign t_5__391_ = t_4__391_ | t_4__407_;
  assign t_5__390_ = t_4__390_ | t_4__406_;
  assign t_5__389_ = t_4__389_ | t_4__405_;
  assign t_5__388_ = t_4__388_ | t_4__404_;
  assign t_5__387_ = t_4__387_ | t_4__403_;
  assign t_5__386_ = t_4__386_ | t_4__402_;
  assign t_5__385_ = t_4__385_ | t_4__401_;
  assign t_5__384_ = t_4__384_ | t_4__400_;
  assign t_5__383_ = t_4__383_ | t_4__399_;
  assign t_5__382_ = t_4__382_ | t_4__398_;
  assign t_5__381_ = t_4__381_ | t_4__397_;
  assign t_5__380_ = t_4__380_ | t_4__396_;
  assign t_5__379_ = t_4__379_ | t_4__395_;
  assign t_5__378_ = t_4__378_ | t_4__394_;
  assign t_5__377_ = t_4__377_ | t_4__393_;
  assign t_5__376_ = t_4__376_ | t_4__392_;
  assign t_5__375_ = t_4__375_ | t_4__391_;
  assign t_5__374_ = t_4__374_ | t_4__390_;
  assign t_5__373_ = t_4__373_ | t_4__389_;
  assign t_5__372_ = t_4__372_ | t_4__388_;
  assign t_5__371_ = t_4__371_ | t_4__387_;
  assign t_5__370_ = t_4__370_ | t_4__386_;
  assign t_5__369_ = t_4__369_ | t_4__385_;
  assign t_5__368_ = t_4__368_ | t_4__384_;
  assign t_5__367_ = t_4__367_ | t_4__383_;
  assign t_5__366_ = t_4__366_ | t_4__382_;
  assign t_5__365_ = t_4__365_ | t_4__381_;
  assign t_5__364_ = t_4__364_ | t_4__380_;
  assign t_5__363_ = t_4__363_ | t_4__379_;
  assign t_5__362_ = t_4__362_ | t_4__378_;
  assign t_5__361_ = t_4__361_ | t_4__377_;
  assign t_5__360_ = t_4__360_ | t_4__376_;
  assign t_5__359_ = t_4__359_ | t_4__375_;
  assign t_5__358_ = t_4__358_ | t_4__374_;
  assign t_5__357_ = t_4__357_ | t_4__373_;
  assign t_5__356_ = t_4__356_ | t_4__372_;
  assign t_5__355_ = t_4__355_ | t_4__371_;
  assign t_5__354_ = t_4__354_ | t_4__370_;
  assign t_5__353_ = t_4__353_ | t_4__369_;
  assign t_5__352_ = t_4__352_ | t_4__368_;
  assign t_5__351_ = t_4__351_ | t_4__367_;
  assign t_5__350_ = t_4__350_ | t_4__366_;
  assign t_5__349_ = t_4__349_ | t_4__365_;
  assign t_5__348_ = t_4__348_ | t_4__364_;
  assign t_5__347_ = t_4__347_ | t_4__363_;
  assign t_5__346_ = t_4__346_ | t_4__362_;
  assign t_5__345_ = t_4__345_ | t_4__361_;
  assign t_5__344_ = t_4__344_ | t_4__360_;
  assign t_5__343_ = t_4__343_ | t_4__359_;
  assign t_5__342_ = t_4__342_ | t_4__358_;
  assign t_5__341_ = t_4__341_ | t_4__357_;
  assign t_5__340_ = t_4__340_ | t_4__356_;
  assign t_5__339_ = t_4__339_ | t_4__355_;
  assign t_5__338_ = t_4__338_ | t_4__354_;
  assign t_5__337_ = t_4__337_ | t_4__353_;
  assign t_5__336_ = t_4__336_ | t_4__352_;
  assign t_5__335_ = t_4__335_ | t_4__351_;
  assign t_5__334_ = t_4__334_ | t_4__350_;
  assign t_5__333_ = t_4__333_ | t_4__349_;
  assign t_5__332_ = t_4__332_ | t_4__348_;
  assign t_5__331_ = t_4__331_ | t_4__347_;
  assign t_5__330_ = t_4__330_ | t_4__346_;
  assign t_5__329_ = t_4__329_ | t_4__345_;
  assign t_5__328_ = t_4__328_ | t_4__344_;
  assign t_5__327_ = t_4__327_ | t_4__343_;
  assign t_5__326_ = t_4__326_ | t_4__342_;
  assign t_5__325_ = t_4__325_ | t_4__341_;
  assign t_5__324_ = t_4__324_ | t_4__340_;
  assign t_5__323_ = t_4__323_ | t_4__339_;
  assign t_5__322_ = t_4__322_ | t_4__338_;
  assign t_5__321_ = t_4__321_ | t_4__337_;
  assign t_5__320_ = t_4__320_ | t_4__336_;
  assign t_5__319_ = t_4__319_ | t_4__335_;
  assign t_5__318_ = t_4__318_ | t_4__334_;
  assign t_5__317_ = t_4__317_ | t_4__333_;
  assign t_5__316_ = t_4__316_ | t_4__332_;
  assign t_5__315_ = t_4__315_ | t_4__331_;
  assign t_5__314_ = t_4__314_ | t_4__330_;
  assign t_5__313_ = t_4__313_ | t_4__329_;
  assign t_5__312_ = t_4__312_ | t_4__328_;
  assign t_5__311_ = t_4__311_ | t_4__327_;
  assign t_5__310_ = t_4__310_ | t_4__326_;
  assign t_5__309_ = t_4__309_ | t_4__325_;
  assign t_5__308_ = t_4__308_ | t_4__324_;
  assign t_5__307_ = t_4__307_ | t_4__323_;
  assign t_5__306_ = t_4__306_ | t_4__322_;
  assign t_5__305_ = t_4__305_ | t_4__321_;
  assign t_5__304_ = t_4__304_ | t_4__320_;
  assign t_5__303_ = t_4__303_ | t_4__319_;
  assign t_5__302_ = t_4__302_ | t_4__318_;
  assign t_5__301_ = t_4__301_ | t_4__317_;
  assign t_5__300_ = t_4__300_ | t_4__316_;
  assign t_5__299_ = t_4__299_ | t_4__315_;
  assign t_5__298_ = t_4__298_ | t_4__314_;
  assign t_5__297_ = t_4__297_ | t_4__313_;
  assign t_5__296_ = t_4__296_ | t_4__312_;
  assign t_5__295_ = t_4__295_ | t_4__311_;
  assign t_5__294_ = t_4__294_ | t_4__310_;
  assign t_5__293_ = t_4__293_ | t_4__309_;
  assign t_5__292_ = t_4__292_ | t_4__308_;
  assign t_5__291_ = t_4__291_ | t_4__307_;
  assign t_5__290_ = t_4__290_ | t_4__306_;
  assign t_5__289_ = t_4__289_ | t_4__305_;
  assign t_5__288_ = t_4__288_ | t_4__304_;
  assign t_5__287_ = t_4__287_ | t_4__303_;
  assign t_5__286_ = t_4__286_ | t_4__302_;
  assign t_5__285_ = t_4__285_ | t_4__301_;
  assign t_5__284_ = t_4__284_ | t_4__300_;
  assign t_5__283_ = t_4__283_ | t_4__299_;
  assign t_5__282_ = t_4__282_ | t_4__298_;
  assign t_5__281_ = t_4__281_ | t_4__297_;
  assign t_5__280_ = t_4__280_ | t_4__296_;
  assign t_5__279_ = t_4__279_ | t_4__295_;
  assign t_5__278_ = t_4__278_ | t_4__294_;
  assign t_5__277_ = t_4__277_ | t_4__293_;
  assign t_5__276_ = t_4__276_ | t_4__292_;
  assign t_5__275_ = t_4__275_ | t_4__291_;
  assign t_5__274_ = t_4__274_ | t_4__290_;
  assign t_5__273_ = t_4__273_ | t_4__289_;
  assign t_5__272_ = t_4__272_ | t_4__288_;
  assign t_5__271_ = t_4__271_ | t_4__287_;
  assign t_5__270_ = t_4__270_ | t_4__286_;
  assign t_5__269_ = t_4__269_ | t_4__285_;
  assign t_5__268_ = t_4__268_ | t_4__284_;
  assign t_5__267_ = t_4__267_ | t_4__283_;
  assign t_5__266_ = t_4__266_ | t_4__282_;
  assign t_5__265_ = t_4__265_ | t_4__281_;
  assign t_5__264_ = t_4__264_ | t_4__280_;
  assign t_5__263_ = t_4__263_ | t_4__279_;
  assign t_5__262_ = t_4__262_ | t_4__278_;
  assign t_5__261_ = t_4__261_ | t_4__277_;
  assign t_5__260_ = t_4__260_ | t_4__276_;
  assign t_5__259_ = t_4__259_ | t_4__275_;
  assign t_5__258_ = t_4__258_ | t_4__274_;
  assign t_5__257_ = t_4__257_ | t_4__273_;
  assign t_5__256_ = t_4__256_ | t_4__272_;
  assign t_5__255_ = t_4__255_ | t_4__271_;
  assign t_5__254_ = t_4__254_ | t_4__270_;
  assign t_5__253_ = t_4__253_ | t_4__269_;
  assign t_5__252_ = t_4__252_ | t_4__268_;
  assign t_5__251_ = t_4__251_ | t_4__267_;
  assign t_5__250_ = t_4__250_ | t_4__266_;
  assign t_5__249_ = t_4__249_ | t_4__265_;
  assign t_5__248_ = t_4__248_ | t_4__264_;
  assign t_5__247_ = t_4__247_ | t_4__263_;
  assign t_5__246_ = t_4__246_ | t_4__262_;
  assign t_5__245_ = t_4__245_ | t_4__261_;
  assign t_5__244_ = t_4__244_ | t_4__260_;
  assign t_5__243_ = t_4__243_ | t_4__259_;
  assign t_5__242_ = t_4__242_ | t_4__258_;
  assign t_5__241_ = t_4__241_ | t_4__257_;
  assign t_5__240_ = t_4__240_ | t_4__256_;
  assign t_5__239_ = t_4__239_ | t_4__255_;
  assign t_5__238_ = t_4__238_ | t_4__254_;
  assign t_5__237_ = t_4__237_ | t_4__253_;
  assign t_5__236_ = t_4__236_ | t_4__252_;
  assign t_5__235_ = t_4__235_ | t_4__251_;
  assign t_5__234_ = t_4__234_ | t_4__250_;
  assign t_5__233_ = t_4__233_ | t_4__249_;
  assign t_5__232_ = t_4__232_ | t_4__248_;
  assign t_5__231_ = t_4__231_ | t_4__247_;
  assign t_5__230_ = t_4__230_ | t_4__246_;
  assign t_5__229_ = t_4__229_ | t_4__245_;
  assign t_5__228_ = t_4__228_ | t_4__244_;
  assign t_5__227_ = t_4__227_ | t_4__243_;
  assign t_5__226_ = t_4__226_ | t_4__242_;
  assign t_5__225_ = t_4__225_ | t_4__241_;
  assign t_5__224_ = t_4__224_ | t_4__240_;
  assign t_5__223_ = t_4__223_ | t_4__239_;
  assign t_5__222_ = t_4__222_ | t_4__238_;
  assign t_5__221_ = t_4__221_ | t_4__237_;
  assign t_5__220_ = t_4__220_ | t_4__236_;
  assign t_5__219_ = t_4__219_ | t_4__235_;
  assign t_5__218_ = t_4__218_ | t_4__234_;
  assign t_5__217_ = t_4__217_ | t_4__233_;
  assign t_5__216_ = t_4__216_ | t_4__232_;
  assign t_5__215_ = t_4__215_ | t_4__231_;
  assign t_5__214_ = t_4__214_ | t_4__230_;
  assign t_5__213_ = t_4__213_ | t_4__229_;
  assign t_5__212_ = t_4__212_ | t_4__228_;
  assign t_5__211_ = t_4__211_ | t_4__227_;
  assign t_5__210_ = t_4__210_ | t_4__226_;
  assign t_5__209_ = t_4__209_ | t_4__225_;
  assign t_5__208_ = t_4__208_ | t_4__224_;
  assign t_5__207_ = t_4__207_ | t_4__223_;
  assign t_5__206_ = t_4__206_ | t_4__222_;
  assign t_5__205_ = t_4__205_ | t_4__221_;
  assign t_5__204_ = t_4__204_ | t_4__220_;
  assign t_5__203_ = t_4__203_ | t_4__219_;
  assign t_5__202_ = t_4__202_ | t_4__218_;
  assign t_5__201_ = t_4__201_ | t_4__217_;
  assign t_5__200_ = t_4__200_ | t_4__216_;
  assign t_5__199_ = t_4__199_ | t_4__215_;
  assign t_5__198_ = t_4__198_ | t_4__214_;
  assign t_5__197_ = t_4__197_ | t_4__213_;
  assign t_5__196_ = t_4__196_ | t_4__212_;
  assign t_5__195_ = t_4__195_ | t_4__211_;
  assign t_5__194_ = t_4__194_ | t_4__210_;
  assign t_5__193_ = t_4__193_ | t_4__209_;
  assign t_5__192_ = t_4__192_ | t_4__208_;
  assign t_5__191_ = t_4__191_ | t_4__207_;
  assign t_5__190_ = t_4__190_ | t_4__206_;
  assign t_5__189_ = t_4__189_ | t_4__205_;
  assign t_5__188_ = t_4__188_ | t_4__204_;
  assign t_5__187_ = t_4__187_ | t_4__203_;
  assign t_5__186_ = t_4__186_ | t_4__202_;
  assign t_5__185_ = t_4__185_ | t_4__201_;
  assign t_5__184_ = t_4__184_ | t_4__200_;
  assign t_5__183_ = t_4__183_ | t_4__199_;
  assign t_5__182_ = t_4__182_ | t_4__198_;
  assign t_5__181_ = t_4__181_ | t_4__197_;
  assign t_5__180_ = t_4__180_ | t_4__196_;
  assign t_5__179_ = t_4__179_ | t_4__195_;
  assign t_5__178_ = t_4__178_ | t_4__194_;
  assign t_5__177_ = t_4__177_ | t_4__193_;
  assign t_5__176_ = t_4__176_ | t_4__192_;
  assign t_5__175_ = t_4__175_ | t_4__191_;
  assign t_5__174_ = t_4__174_ | t_4__190_;
  assign t_5__173_ = t_4__173_ | t_4__189_;
  assign t_5__172_ = t_4__172_ | t_4__188_;
  assign t_5__171_ = t_4__171_ | t_4__187_;
  assign t_5__170_ = t_4__170_ | t_4__186_;
  assign t_5__169_ = t_4__169_ | t_4__185_;
  assign t_5__168_ = t_4__168_ | t_4__184_;
  assign t_5__167_ = t_4__167_ | t_4__183_;
  assign t_5__166_ = t_4__166_ | t_4__182_;
  assign t_5__165_ = t_4__165_ | t_4__181_;
  assign t_5__164_ = t_4__164_ | t_4__180_;
  assign t_5__163_ = t_4__163_ | t_4__179_;
  assign t_5__162_ = t_4__162_ | t_4__178_;
  assign t_5__161_ = t_4__161_ | t_4__177_;
  assign t_5__160_ = t_4__160_ | t_4__176_;
  assign t_5__159_ = t_4__159_ | t_4__175_;
  assign t_5__158_ = t_4__158_ | t_4__174_;
  assign t_5__157_ = t_4__157_ | t_4__173_;
  assign t_5__156_ = t_4__156_ | t_4__172_;
  assign t_5__155_ = t_4__155_ | t_4__171_;
  assign t_5__154_ = t_4__154_ | t_4__170_;
  assign t_5__153_ = t_4__153_ | t_4__169_;
  assign t_5__152_ = t_4__152_ | t_4__168_;
  assign t_5__151_ = t_4__151_ | t_4__167_;
  assign t_5__150_ = t_4__150_ | t_4__166_;
  assign t_5__149_ = t_4__149_ | t_4__165_;
  assign t_5__148_ = t_4__148_ | t_4__164_;
  assign t_5__147_ = t_4__147_ | t_4__163_;
  assign t_5__146_ = t_4__146_ | t_4__162_;
  assign t_5__145_ = t_4__145_ | t_4__161_;
  assign t_5__144_ = t_4__144_ | t_4__160_;
  assign t_5__143_ = t_4__143_ | t_4__159_;
  assign t_5__142_ = t_4__142_ | t_4__158_;
  assign t_5__141_ = t_4__141_ | t_4__157_;
  assign t_5__140_ = t_4__140_ | t_4__156_;
  assign t_5__139_ = t_4__139_ | t_4__155_;
  assign t_5__138_ = t_4__138_ | t_4__154_;
  assign t_5__137_ = t_4__137_ | t_4__153_;
  assign t_5__136_ = t_4__136_ | t_4__152_;
  assign t_5__135_ = t_4__135_ | t_4__151_;
  assign t_5__134_ = t_4__134_ | t_4__150_;
  assign t_5__133_ = t_4__133_ | t_4__149_;
  assign t_5__132_ = t_4__132_ | t_4__148_;
  assign t_5__131_ = t_4__131_ | t_4__147_;
  assign t_5__130_ = t_4__130_ | t_4__146_;
  assign t_5__129_ = t_4__129_ | t_4__145_;
  assign t_5__128_ = t_4__128_ | t_4__144_;
  assign t_5__127_ = t_4__127_ | t_4__143_;
  assign t_5__126_ = t_4__126_ | t_4__142_;
  assign t_5__125_ = t_4__125_ | t_4__141_;
  assign t_5__124_ = t_4__124_ | t_4__140_;
  assign t_5__123_ = t_4__123_ | t_4__139_;
  assign t_5__122_ = t_4__122_ | t_4__138_;
  assign t_5__121_ = t_4__121_ | t_4__137_;
  assign t_5__120_ = t_4__120_ | t_4__136_;
  assign t_5__119_ = t_4__119_ | t_4__135_;
  assign t_5__118_ = t_4__118_ | t_4__134_;
  assign t_5__117_ = t_4__117_ | t_4__133_;
  assign t_5__116_ = t_4__116_ | t_4__132_;
  assign t_5__115_ = t_4__115_ | t_4__131_;
  assign t_5__114_ = t_4__114_ | t_4__130_;
  assign t_5__113_ = t_4__113_ | t_4__129_;
  assign t_5__112_ = t_4__112_ | t_4__128_;
  assign t_5__111_ = t_4__111_ | t_4__127_;
  assign t_5__110_ = t_4__110_ | t_4__126_;
  assign t_5__109_ = t_4__109_ | t_4__125_;
  assign t_5__108_ = t_4__108_ | t_4__124_;
  assign t_5__107_ = t_4__107_ | t_4__123_;
  assign t_5__106_ = t_4__106_ | t_4__122_;
  assign t_5__105_ = t_4__105_ | t_4__121_;
  assign t_5__104_ = t_4__104_ | t_4__120_;
  assign t_5__103_ = t_4__103_ | t_4__119_;
  assign t_5__102_ = t_4__102_ | t_4__118_;
  assign t_5__101_ = t_4__101_ | t_4__117_;
  assign t_5__100_ = t_4__100_ | t_4__116_;
  assign t_5__99_ = t_4__99_ | t_4__115_;
  assign t_5__98_ = t_4__98_ | t_4__114_;
  assign t_5__97_ = t_4__97_ | t_4__113_;
  assign t_5__96_ = t_4__96_ | t_4__112_;
  assign t_5__95_ = t_4__95_ | t_4__111_;
  assign t_5__94_ = t_4__94_ | t_4__110_;
  assign t_5__93_ = t_4__93_ | t_4__109_;
  assign t_5__92_ = t_4__92_ | t_4__108_;
  assign t_5__91_ = t_4__91_ | t_4__107_;
  assign t_5__90_ = t_4__90_ | t_4__106_;
  assign t_5__89_ = t_4__89_ | t_4__105_;
  assign t_5__88_ = t_4__88_ | t_4__104_;
  assign t_5__87_ = t_4__87_ | t_4__103_;
  assign t_5__86_ = t_4__86_ | t_4__102_;
  assign t_5__85_ = t_4__85_ | t_4__101_;
  assign t_5__84_ = t_4__84_ | t_4__100_;
  assign t_5__83_ = t_4__83_ | t_4__99_;
  assign t_5__82_ = t_4__82_ | t_4__98_;
  assign t_5__81_ = t_4__81_ | t_4__97_;
  assign t_5__80_ = t_4__80_ | t_4__96_;
  assign t_5__79_ = t_4__79_ | t_4__95_;
  assign t_5__78_ = t_4__78_ | t_4__94_;
  assign t_5__77_ = t_4__77_ | t_4__93_;
  assign t_5__76_ = t_4__76_ | t_4__92_;
  assign t_5__75_ = t_4__75_ | t_4__91_;
  assign t_5__74_ = t_4__74_ | t_4__90_;
  assign t_5__73_ = t_4__73_ | t_4__89_;
  assign t_5__72_ = t_4__72_ | t_4__88_;
  assign t_5__71_ = t_4__71_ | t_4__87_;
  assign t_5__70_ = t_4__70_ | t_4__86_;
  assign t_5__69_ = t_4__69_ | t_4__85_;
  assign t_5__68_ = t_4__68_ | t_4__84_;
  assign t_5__67_ = t_4__67_ | t_4__83_;
  assign t_5__66_ = t_4__66_ | t_4__82_;
  assign t_5__65_ = t_4__65_ | t_4__81_;
  assign t_5__64_ = t_4__64_ | t_4__80_;
  assign t_5__63_ = t_4__63_ | t_4__79_;
  assign t_5__62_ = t_4__62_ | t_4__78_;
  assign t_5__61_ = t_4__61_ | t_4__77_;
  assign t_5__60_ = t_4__60_ | t_4__76_;
  assign t_5__59_ = t_4__59_ | t_4__75_;
  assign t_5__58_ = t_4__58_ | t_4__74_;
  assign t_5__57_ = t_4__57_ | t_4__73_;
  assign t_5__56_ = t_4__56_ | t_4__72_;
  assign t_5__55_ = t_4__55_ | t_4__71_;
  assign t_5__54_ = t_4__54_ | t_4__70_;
  assign t_5__53_ = t_4__53_ | t_4__69_;
  assign t_5__52_ = t_4__52_ | t_4__68_;
  assign t_5__51_ = t_4__51_ | t_4__67_;
  assign t_5__50_ = t_4__50_ | t_4__66_;
  assign t_5__49_ = t_4__49_ | t_4__65_;
  assign t_5__48_ = t_4__48_ | t_4__64_;
  assign t_5__47_ = t_4__47_ | t_4__63_;
  assign t_5__46_ = t_4__46_ | t_4__62_;
  assign t_5__45_ = t_4__45_ | t_4__61_;
  assign t_5__44_ = t_4__44_ | t_4__60_;
  assign t_5__43_ = t_4__43_ | t_4__59_;
  assign t_5__42_ = t_4__42_ | t_4__58_;
  assign t_5__41_ = t_4__41_ | t_4__57_;
  assign t_5__40_ = t_4__40_ | t_4__56_;
  assign t_5__39_ = t_4__39_ | t_4__55_;
  assign t_5__38_ = t_4__38_ | t_4__54_;
  assign t_5__37_ = t_4__37_ | t_4__53_;
  assign t_5__36_ = t_4__36_ | t_4__52_;
  assign t_5__35_ = t_4__35_ | t_4__51_;
  assign t_5__34_ = t_4__34_ | t_4__50_;
  assign t_5__33_ = t_4__33_ | t_4__49_;
  assign t_5__32_ = t_4__32_ | t_4__48_;
  assign t_5__31_ = t_4__31_ | t_4__47_;
  assign t_5__30_ = t_4__30_ | t_4__46_;
  assign t_5__29_ = t_4__29_ | t_4__45_;
  assign t_5__28_ = t_4__28_ | t_4__44_;
  assign t_5__27_ = t_4__27_ | t_4__43_;
  assign t_5__26_ = t_4__26_ | t_4__42_;
  assign t_5__25_ = t_4__25_ | t_4__41_;
  assign t_5__24_ = t_4__24_ | t_4__40_;
  assign t_5__23_ = t_4__23_ | t_4__39_;
  assign t_5__22_ = t_4__22_ | t_4__38_;
  assign t_5__21_ = t_4__21_ | t_4__37_;
  assign t_5__20_ = t_4__20_ | t_4__36_;
  assign t_5__19_ = t_4__19_ | t_4__35_;
  assign t_5__18_ = t_4__18_ | t_4__34_;
  assign t_5__17_ = t_4__17_ | t_4__33_;
  assign t_5__16_ = t_4__16_ | t_4__32_;
  assign t_5__15_ = t_4__15_ | t_4__31_;
  assign t_5__14_ = t_4__14_ | t_4__30_;
  assign t_5__13_ = t_4__13_ | t_4__29_;
  assign t_5__12_ = t_4__12_ | t_4__28_;
  assign t_5__11_ = t_4__11_ | t_4__27_;
  assign t_5__10_ = t_4__10_ | t_4__26_;
  assign t_5__9_ = t_4__9_ | t_4__25_;
  assign t_5__8_ = t_4__8_ | t_4__24_;
  assign t_5__7_ = t_4__7_ | t_4__23_;
  assign t_5__6_ = t_4__6_ | t_4__22_;
  assign t_5__5_ = t_4__5_ | t_4__21_;
  assign t_5__4_ = t_4__4_ | t_4__20_;
  assign t_5__3_ = t_4__3_ | t_4__19_;
  assign t_5__2_ = t_4__2_ | t_4__18_;
  assign t_5__1_ = t_4__1_ | t_4__17_;
  assign t_5__0_ = t_4__0_ | t_4__16_;
  assign t_6__1023_ = t_5__1023_ | 1'b0;
  assign t_6__1022_ = t_5__1022_ | 1'b0;
  assign t_6__1021_ = t_5__1021_ | 1'b0;
  assign t_6__1020_ = t_5__1020_ | 1'b0;
  assign t_6__1019_ = t_5__1019_ | 1'b0;
  assign t_6__1018_ = t_5__1018_ | 1'b0;
  assign t_6__1017_ = t_5__1017_ | 1'b0;
  assign t_6__1016_ = t_5__1016_ | 1'b0;
  assign t_6__1015_ = t_5__1015_ | 1'b0;
  assign t_6__1014_ = t_5__1014_ | 1'b0;
  assign t_6__1013_ = t_5__1013_ | 1'b0;
  assign t_6__1012_ = t_5__1012_ | 1'b0;
  assign t_6__1011_ = t_5__1011_ | 1'b0;
  assign t_6__1010_ = t_5__1010_ | 1'b0;
  assign t_6__1009_ = t_5__1009_ | 1'b0;
  assign t_6__1008_ = t_5__1008_ | 1'b0;
  assign t_6__1007_ = t_5__1007_ | 1'b0;
  assign t_6__1006_ = t_5__1006_ | 1'b0;
  assign t_6__1005_ = t_5__1005_ | 1'b0;
  assign t_6__1004_ = t_5__1004_ | 1'b0;
  assign t_6__1003_ = t_5__1003_ | 1'b0;
  assign t_6__1002_ = t_5__1002_ | 1'b0;
  assign t_6__1001_ = t_5__1001_ | 1'b0;
  assign t_6__1000_ = t_5__1000_ | 1'b0;
  assign t_6__999_ = t_5__999_ | 1'b0;
  assign t_6__998_ = t_5__998_ | 1'b0;
  assign t_6__997_ = t_5__997_ | 1'b0;
  assign t_6__996_ = t_5__996_ | 1'b0;
  assign t_6__995_ = t_5__995_ | 1'b0;
  assign t_6__994_ = t_5__994_ | 1'b0;
  assign t_6__993_ = t_5__993_ | 1'b0;
  assign t_6__992_ = t_5__992_ | 1'b0;
  assign t_6__991_ = t_5__991_ | t_5__1023_;
  assign t_6__990_ = t_5__990_ | t_5__1022_;
  assign t_6__989_ = t_5__989_ | t_5__1021_;
  assign t_6__988_ = t_5__988_ | t_5__1020_;
  assign t_6__987_ = t_5__987_ | t_5__1019_;
  assign t_6__986_ = t_5__986_ | t_5__1018_;
  assign t_6__985_ = t_5__985_ | t_5__1017_;
  assign t_6__984_ = t_5__984_ | t_5__1016_;
  assign t_6__983_ = t_5__983_ | t_5__1015_;
  assign t_6__982_ = t_5__982_ | t_5__1014_;
  assign t_6__981_ = t_5__981_ | t_5__1013_;
  assign t_6__980_ = t_5__980_ | t_5__1012_;
  assign t_6__979_ = t_5__979_ | t_5__1011_;
  assign t_6__978_ = t_5__978_ | t_5__1010_;
  assign t_6__977_ = t_5__977_ | t_5__1009_;
  assign t_6__976_ = t_5__976_ | t_5__1008_;
  assign t_6__975_ = t_5__975_ | t_5__1007_;
  assign t_6__974_ = t_5__974_ | t_5__1006_;
  assign t_6__973_ = t_5__973_ | t_5__1005_;
  assign t_6__972_ = t_5__972_ | t_5__1004_;
  assign t_6__971_ = t_5__971_ | t_5__1003_;
  assign t_6__970_ = t_5__970_ | t_5__1002_;
  assign t_6__969_ = t_5__969_ | t_5__1001_;
  assign t_6__968_ = t_5__968_ | t_5__1000_;
  assign t_6__967_ = t_5__967_ | t_5__999_;
  assign t_6__966_ = t_5__966_ | t_5__998_;
  assign t_6__965_ = t_5__965_ | t_5__997_;
  assign t_6__964_ = t_5__964_ | t_5__996_;
  assign t_6__963_ = t_5__963_ | t_5__995_;
  assign t_6__962_ = t_5__962_ | t_5__994_;
  assign t_6__961_ = t_5__961_ | t_5__993_;
  assign t_6__960_ = t_5__960_ | t_5__992_;
  assign t_6__959_ = t_5__959_ | t_5__991_;
  assign t_6__958_ = t_5__958_ | t_5__990_;
  assign t_6__957_ = t_5__957_ | t_5__989_;
  assign t_6__956_ = t_5__956_ | t_5__988_;
  assign t_6__955_ = t_5__955_ | t_5__987_;
  assign t_6__954_ = t_5__954_ | t_5__986_;
  assign t_6__953_ = t_5__953_ | t_5__985_;
  assign t_6__952_ = t_5__952_ | t_5__984_;
  assign t_6__951_ = t_5__951_ | t_5__983_;
  assign t_6__950_ = t_5__950_ | t_5__982_;
  assign t_6__949_ = t_5__949_ | t_5__981_;
  assign t_6__948_ = t_5__948_ | t_5__980_;
  assign t_6__947_ = t_5__947_ | t_5__979_;
  assign t_6__946_ = t_5__946_ | t_5__978_;
  assign t_6__945_ = t_5__945_ | t_5__977_;
  assign t_6__944_ = t_5__944_ | t_5__976_;
  assign t_6__943_ = t_5__943_ | t_5__975_;
  assign t_6__942_ = t_5__942_ | t_5__974_;
  assign t_6__941_ = t_5__941_ | t_5__973_;
  assign t_6__940_ = t_5__940_ | t_5__972_;
  assign t_6__939_ = t_5__939_ | t_5__971_;
  assign t_6__938_ = t_5__938_ | t_5__970_;
  assign t_6__937_ = t_5__937_ | t_5__969_;
  assign t_6__936_ = t_5__936_ | t_5__968_;
  assign t_6__935_ = t_5__935_ | t_5__967_;
  assign t_6__934_ = t_5__934_ | t_5__966_;
  assign t_6__933_ = t_5__933_ | t_5__965_;
  assign t_6__932_ = t_5__932_ | t_5__964_;
  assign t_6__931_ = t_5__931_ | t_5__963_;
  assign t_6__930_ = t_5__930_ | t_5__962_;
  assign t_6__929_ = t_5__929_ | t_5__961_;
  assign t_6__928_ = t_5__928_ | t_5__960_;
  assign t_6__927_ = t_5__927_ | t_5__959_;
  assign t_6__926_ = t_5__926_ | t_5__958_;
  assign t_6__925_ = t_5__925_ | t_5__957_;
  assign t_6__924_ = t_5__924_ | t_5__956_;
  assign t_6__923_ = t_5__923_ | t_5__955_;
  assign t_6__922_ = t_5__922_ | t_5__954_;
  assign t_6__921_ = t_5__921_ | t_5__953_;
  assign t_6__920_ = t_5__920_ | t_5__952_;
  assign t_6__919_ = t_5__919_ | t_5__951_;
  assign t_6__918_ = t_5__918_ | t_5__950_;
  assign t_6__917_ = t_5__917_ | t_5__949_;
  assign t_6__916_ = t_5__916_ | t_5__948_;
  assign t_6__915_ = t_5__915_ | t_5__947_;
  assign t_6__914_ = t_5__914_ | t_5__946_;
  assign t_6__913_ = t_5__913_ | t_5__945_;
  assign t_6__912_ = t_5__912_ | t_5__944_;
  assign t_6__911_ = t_5__911_ | t_5__943_;
  assign t_6__910_ = t_5__910_ | t_5__942_;
  assign t_6__909_ = t_5__909_ | t_5__941_;
  assign t_6__908_ = t_5__908_ | t_5__940_;
  assign t_6__907_ = t_5__907_ | t_5__939_;
  assign t_6__906_ = t_5__906_ | t_5__938_;
  assign t_6__905_ = t_5__905_ | t_5__937_;
  assign t_6__904_ = t_5__904_ | t_5__936_;
  assign t_6__903_ = t_5__903_ | t_5__935_;
  assign t_6__902_ = t_5__902_ | t_5__934_;
  assign t_6__901_ = t_5__901_ | t_5__933_;
  assign t_6__900_ = t_5__900_ | t_5__932_;
  assign t_6__899_ = t_5__899_ | t_5__931_;
  assign t_6__898_ = t_5__898_ | t_5__930_;
  assign t_6__897_ = t_5__897_ | t_5__929_;
  assign t_6__896_ = t_5__896_ | t_5__928_;
  assign t_6__895_ = t_5__895_ | t_5__927_;
  assign t_6__894_ = t_5__894_ | t_5__926_;
  assign t_6__893_ = t_5__893_ | t_5__925_;
  assign t_6__892_ = t_5__892_ | t_5__924_;
  assign t_6__891_ = t_5__891_ | t_5__923_;
  assign t_6__890_ = t_5__890_ | t_5__922_;
  assign t_6__889_ = t_5__889_ | t_5__921_;
  assign t_6__888_ = t_5__888_ | t_5__920_;
  assign t_6__887_ = t_5__887_ | t_5__919_;
  assign t_6__886_ = t_5__886_ | t_5__918_;
  assign t_6__885_ = t_5__885_ | t_5__917_;
  assign t_6__884_ = t_5__884_ | t_5__916_;
  assign t_6__883_ = t_5__883_ | t_5__915_;
  assign t_6__882_ = t_5__882_ | t_5__914_;
  assign t_6__881_ = t_5__881_ | t_5__913_;
  assign t_6__880_ = t_5__880_ | t_5__912_;
  assign t_6__879_ = t_5__879_ | t_5__911_;
  assign t_6__878_ = t_5__878_ | t_5__910_;
  assign t_6__877_ = t_5__877_ | t_5__909_;
  assign t_6__876_ = t_5__876_ | t_5__908_;
  assign t_6__875_ = t_5__875_ | t_5__907_;
  assign t_6__874_ = t_5__874_ | t_5__906_;
  assign t_6__873_ = t_5__873_ | t_5__905_;
  assign t_6__872_ = t_5__872_ | t_5__904_;
  assign t_6__871_ = t_5__871_ | t_5__903_;
  assign t_6__870_ = t_5__870_ | t_5__902_;
  assign t_6__869_ = t_5__869_ | t_5__901_;
  assign t_6__868_ = t_5__868_ | t_5__900_;
  assign t_6__867_ = t_5__867_ | t_5__899_;
  assign t_6__866_ = t_5__866_ | t_5__898_;
  assign t_6__865_ = t_5__865_ | t_5__897_;
  assign t_6__864_ = t_5__864_ | t_5__896_;
  assign t_6__863_ = t_5__863_ | t_5__895_;
  assign t_6__862_ = t_5__862_ | t_5__894_;
  assign t_6__861_ = t_5__861_ | t_5__893_;
  assign t_6__860_ = t_5__860_ | t_5__892_;
  assign t_6__859_ = t_5__859_ | t_5__891_;
  assign t_6__858_ = t_5__858_ | t_5__890_;
  assign t_6__857_ = t_5__857_ | t_5__889_;
  assign t_6__856_ = t_5__856_ | t_5__888_;
  assign t_6__855_ = t_5__855_ | t_5__887_;
  assign t_6__854_ = t_5__854_ | t_5__886_;
  assign t_6__853_ = t_5__853_ | t_5__885_;
  assign t_6__852_ = t_5__852_ | t_5__884_;
  assign t_6__851_ = t_5__851_ | t_5__883_;
  assign t_6__850_ = t_5__850_ | t_5__882_;
  assign t_6__849_ = t_5__849_ | t_5__881_;
  assign t_6__848_ = t_5__848_ | t_5__880_;
  assign t_6__847_ = t_5__847_ | t_5__879_;
  assign t_6__846_ = t_5__846_ | t_5__878_;
  assign t_6__845_ = t_5__845_ | t_5__877_;
  assign t_6__844_ = t_5__844_ | t_5__876_;
  assign t_6__843_ = t_5__843_ | t_5__875_;
  assign t_6__842_ = t_5__842_ | t_5__874_;
  assign t_6__841_ = t_5__841_ | t_5__873_;
  assign t_6__840_ = t_5__840_ | t_5__872_;
  assign t_6__839_ = t_5__839_ | t_5__871_;
  assign t_6__838_ = t_5__838_ | t_5__870_;
  assign t_6__837_ = t_5__837_ | t_5__869_;
  assign t_6__836_ = t_5__836_ | t_5__868_;
  assign t_6__835_ = t_5__835_ | t_5__867_;
  assign t_6__834_ = t_5__834_ | t_5__866_;
  assign t_6__833_ = t_5__833_ | t_5__865_;
  assign t_6__832_ = t_5__832_ | t_5__864_;
  assign t_6__831_ = t_5__831_ | t_5__863_;
  assign t_6__830_ = t_5__830_ | t_5__862_;
  assign t_6__829_ = t_5__829_ | t_5__861_;
  assign t_6__828_ = t_5__828_ | t_5__860_;
  assign t_6__827_ = t_5__827_ | t_5__859_;
  assign t_6__826_ = t_5__826_ | t_5__858_;
  assign t_6__825_ = t_5__825_ | t_5__857_;
  assign t_6__824_ = t_5__824_ | t_5__856_;
  assign t_6__823_ = t_5__823_ | t_5__855_;
  assign t_6__822_ = t_5__822_ | t_5__854_;
  assign t_6__821_ = t_5__821_ | t_5__853_;
  assign t_6__820_ = t_5__820_ | t_5__852_;
  assign t_6__819_ = t_5__819_ | t_5__851_;
  assign t_6__818_ = t_5__818_ | t_5__850_;
  assign t_6__817_ = t_5__817_ | t_5__849_;
  assign t_6__816_ = t_5__816_ | t_5__848_;
  assign t_6__815_ = t_5__815_ | t_5__847_;
  assign t_6__814_ = t_5__814_ | t_5__846_;
  assign t_6__813_ = t_5__813_ | t_5__845_;
  assign t_6__812_ = t_5__812_ | t_5__844_;
  assign t_6__811_ = t_5__811_ | t_5__843_;
  assign t_6__810_ = t_5__810_ | t_5__842_;
  assign t_6__809_ = t_5__809_ | t_5__841_;
  assign t_6__808_ = t_5__808_ | t_5__840_;
  assign t_6__807_ = t_5__807_ | t_5__839_;
  assign t_6__806_ = t_5__806_ | t_5__838_;
  assign t_6__805_ = t_5__805_ | t_5__837_;
  assign t_6__804_ = t_5__804_ | t_5__836_;
  assign t_6__803_ = t_5__803_ | t_5__835_;
  assign t_6__802_ = t_5__802_ | t_5__834_;
  assign t_6__801_ = t_5__801_ | t_5__833_;
  assign t_6__800_ = t_5__800_ | t_5__832_;
  assign t_6__799_ = t_5__799_ | t_5__831_;
  assign t_6__798_ = t_5__798_ | t_5__830_;
  assign t_6__797_ = t_5__797_ | t_5__829_;
  assign t_6__796_ = t_5__796_ | t_5__828_;
  assign t_6__795_ = t_5__795_ | t_5__827_;
  assign t_6__794_ = t_5__794_ | t_5__826_;
  assign t_6__793_ = t_5__793_ | t_5__825_;
  assign t_6__792_ = t_5__792_ | t_5__824_;
  assign t_6__791_ = t_5__791_ | t_5__823_;
  assign t_6__790_ = t_5__790_ | t_5__822_;
  assign t_6__789_ = t_5__789_ | t_5__821_;
  assign t_6__788_ = t_5__788_ | t_5__820_;
  assign t_6__787_ = t_5__787_ | t_5__819_;
  assign t_6__786_ = t_5__786_ | t_5__818_;
  assign t_6__785_ = t_5__785_ | t_5__817_;
  assign t_6__784_ = t_5__784_ | t_5__816_;
  assign t_6__783_ = t_5__783_ | t_5__815_;
  assign t_6__782_ = t_5__782_ | t_5__814_;
  assign t_6__781_ = t_5__781_ | t_5__813_;
  assign t_6__780_ = t_5__780_ | t_5__812_;
  assign t_6__779_ = t_5__779_ | t_5__811_;
  assign t_6__778_ = t_5__778_ | t_5__810_;
  assign t_6__777_ = t_5__777_ | t_5__809_;
  assign t_6__776_ = t_5__776_ | t_5__808_;
  assign t_6__775_ = t_5__775_ | t_5__807_;
  assign t_6__774_ = t_5__774_ | t_5__806_;
  assign t_6__773_ = t_5__773_ | t_5__805_;
  assign t_6__772_ = t_5__772_ | t_5__804_;
  assign t_6__771_ = t_5__771_ | t_5__803_;
  assign t_6__770_ = t_5__770_ | t_5__802_;
  assign t_6__769_ = t_5__769_ | t_5__801_;
  assign t_6__768_ = t_5__768_ | t_5__800_;
  assign t_6__767_ = t_5__767_ | t_5__799_;
  assign t_6__766_ = t_5__766_ | t_5__798_;
  assign t_6__765_ = t_5__765_ | t_5__797_;
  assign t_6__764_ = t_5__764_ | t_5__796_;
  assign t_6__763_ = t_5__763_ | t_5__795_;
  assign t_6__762_ = t_5__762_ | t_5__794_;
  assign t_6__761_ = t_5__761_ | t_5__793_;
  assign t_6__760_ = t_5__760_ | t_5__792_;
  assign t_6__759_ = t_5__759_ | t_5__791_;
  assign t_6__758_ = t_5__758_ | t_5__790_;
  assign t_6__757_ = t_5__757_ | t_5__789_;
  assign t_6__756_ = t_5__756_ | t_5__788_;
  assign t_6__755_ = t_5__755_ | t_5__787_;
  assign t_6__754_ = t_5__754_ | t_5__786_;
  assign t_6__753_ = t_5__753_ | t_5__785_;
  assign t_6__752_ = t_5__752_ | t_5__784_;
  assign t_6__751_ = t_5__751_ | t_5__783_;
  assign t_6__750_ = t_5__750_ | t_5__782_;
  assign t_6__749_ = t_5__749_ | t_5__781_;
  assign t_6__748_ = t_5__748_ | t_5__780_;
  assign t_6__747_ = t_5__747_ | t_5__779_;
  assign t_6__746_ = t_5__746_ | t_5__778_;
  assign t_6__745_ = t_5__745_ | t_5__777_;
  assign t_6__744_ = t_5__744_ | t_5__776_;
  assign t_6__743_ = t_5__743_ | t_5__775_;
  assign t_6__742_ = t_5__742_ | t_5__774_;
  assign t_6__741_ = t_5__741_ | t_5__773_;
  assign t_6__740_ = t_5__740_ | t_5__772_;
  assign t_6__739_ = t_5__739_ | t_5__771_;
  assign t_6__738_ = t_5__738_ | t_5__770_;
  assign t_6__737_ = t_5__737_ | t_5__769_;
  assign t_6__736_ = t_5__736_ | t_5__768_;
  assign t_6__735_ = t_5__735_ | t_5__767_;
  assign t_6__734_ = t_5__734_ | t_5__766_;
  assign t_6__733_ = t_5__733_ | t_5__765_;
  assign t_6__732_ = t_5__732_ | t_5__764_;
  assign t_6__731_ = t_5__731_ | t_5__763_;
  assign t_6__730_ = t_5__730_ | t_5__762_;
  assign t_6__729_ = t_5__729_ | t_5__761_;
  assign t_6__728_ = t_5__728_ | t_5__760_;
  assign t_6__727_ = t_5__727_ | t_5__759_;
  assign t_6__726_ = t_5__726_ | t_5__758_;
  assign t_6__725_ = t_5__725_ | t_5__757_;
  assign t_6__724_ = t_5__724_ | t_5__756_;
  assign t_6__723_ = t_5__723_ | t_5__755_;
  assign t_6__722_ = t_5__722_ | t_5__754_;
  assign t_6__721_ = t_5__721_ | t_5__753_;
  assign t_6__720_ = t_5__720_ | t_5__752_;
  assign t_6__719_ = t_5__719_ | t_5__751_;
  assign t_6__718_ = t_5__718_ | t_5__750_;
  assign t_6__717_ = t_5__717_ | t_5__749_;
  assign t_6__716_ = t_5__716_ | t_5__748_;
  assign t_6__715_ = t_5__715_ | t_5__747_;
  assign t_6__714_ = t_5__714_ | t_5__746_;
  assign t_6__713_ = t_5__713_ | t_5__745_;
  assign t_6__712_ = t_5__712_ | t_5__744_;
  assign t_6__711_ = t_5__711_ | t_5__743_;
  assign t_6__710_ = t_5__710_ | t_5__742_;
  assign t_6__709_ = t_5__709_ | t_5__741_;
  assign t_6__708_ = t_5__708_ | t_5__740_;
  assign t_6__707_ = t_5__707_ | t_5__739_;
  assign t_6__706_ = t_5__706_ | t_5__738_;
  assign t_6__705_ = t_5__705_ | t_5__737_;
  assign t_6__704_ = t_5__704_ | t_5__736_;
  assign t_6__703_ = t_5__703_ | t_5__735_;
  assign t_6__702_ = t_5__702_ | t_5__734_;
  assign t_6__701_ = t_5__701_ | t_5__733_;
  assign t_6__700_ = t_5__700_ | t_5__732_;
  assign t_6__699_ = t_5__699_ | t_5__731_;
  assign t_6__698_ = t_5__698_ | t_5__730_;
  assign t_6__697_ = t_5__697_ | t_5__729_;
  assign t_6__696_ = t_5__696_ | t_5__728_;
  assign t_6__695_ = t_5__695_ | t_5__727_;
  assign t_6__694_ = t_5__694_ | t_5__726_;
  assign t_6__693_ = t_5__693_ | t_5__725_;
  assign t_6__692_ = t_5__692_ | t_5__724_;
  assign t_6__691_ = t_5__691_ | t_5__723_;
  assign t_6__690_ = t_5__690_ | t_5__722_;
  assign t_6__689_ = t_5__689_ | t_5__721_;
  assign t_6__688_ = t_5__688_ | t_5__720_;
  assign t_6__687_ = t_5__687_ | t_5__719_;
  assign t_6__686_ = t_5__686_ | t_5__718_;
  assign t_6__685_ = t_5__685_ | t_5__717_;
  assign t_6__684_ = t_5__684_ | t_5__716_;
  assign t_6__683_ = t_5__683_ | t_5__715_;
  assign t_6__682_ = t_5__682_ | t_5__714_;
  assign t_6__681_ = t_5__681_ | t_5__713_;
  assign t_6__680_ = t_5__680_ | t_5__712_;
  assign t_6__679_ = t_5__679_ | t_5__711_;
  assign t_6__678_ = t_5__678_ | t_5__710_;
  assign t_6__677_ = t_5__677_ | t_5__709_;
  assign t_6__676_ = t_5__676_ | t_5__708_;
  assign t_6__675_ = t_5__675_ | t_5__707_;
  assign t_6__674_ = t_5__674_ | t_5__706_;
  assign t_6__673_ = t_5__673_ | t_5__705_;
  assign t_6__672_ = t_5__672_ | t_5__704_;
  assign t_6__671_ = t_5__671_ | t_5__703_;
  assign t_6__670_ = t_5__670_ | t_5__702_;
  assign t_6__669_ = t_5__669_ | t_5__701_;
  assign t_6__668_ = t_5__668_ | t_5__700_;
  assign t_6__667_ = t_5__667_ | t_5__699_;
  assign t_6__666_ = t_5__666_ | t_5__698_;
  assign t_6__665_ = t_5__665_ | t_5__697_;
  assign t_6__664_ = t_5__664_ | t_5__696_;
  assign t_6__663_ = t_5__663_ | t_5__695_;
  assign t_6__662_ = t_5__662_ | t_5__694_;
  assign t_6__661_ = t_5__661_ | t_5__693_;
  assign t_6__660_ = t_5__660_ | t_5__692_;
  assign t_6__659_ = t_5__659_ | t_5__691_;
  assign t_6__658_ = t_5__658_ | t_5__690_;
  assign t_6__657_ = t_5__657_ | t_5__689_;
  assign t_6__656_ = t_5__656_ | t_5__688_;
  assign t_6__655_ = t_5__655_ | t_5__687_;
  assign t_6__654_ = t_5__654_ | t_5__686_;
  assign t_6__653_ = t_5__653_ | t_5__685_;
  assign t_6__652_ = t_5__652_ | t_5__684_;
  assign t_6__651_ = t_5__651_ | t_5__683_;
  assign t_6__650_ = t_5__650_ | t_5__682_;
  assign t_6__649_ = t_5__649_ | t_5__681_;
  assign t_6__648_ = t_5__648_ | t_5__680_;
  assign t_6__647_ = t_5__647_ | t_5__679_;
  assign t_6__646_ = t_5__646_ | t_5__678_;
  assign t_6__645_ = t_5__645_ | t_5__677_;
  assign t_6__644_ = t_5__644_ | t_5__676_;
  assign t_6__643_ = t_5__643_ | t_5__675_;
  assign t_6__642_ = t_5__642_ | t_5__674_;
  assign t_6__641_ = t_5__641_ | t_5__673_;
  assign t_6__640_ = t_5__640_ | t_5__672_;
  assign t_6__639_ = t_5__639_ | t_5__671_;
  assign t_6__638_ = t_5__638_ | t_5__670_;
  assign t_6__637_ = t_5__637_ | t_5__669_;
  assign t_6__636_ = t_5__636_ | t_5__668_;
  assign t_6__635_ = t_5__635_ | t_5__667_;
  assign t_6__634_ = t_5__634_ | t_5__666_;
  assign t_6__633_ = t_5__633_ | t_5__665_;
  assign t_6__632_ = t_5__632_ | t_5__664_;
  assign t_6__631_ = t_5__631_ | t_5__663_;
  assign t_6__630_ = t_5__630_ | t_5__662_;
  assign t_6__629_ = t_5__629_ | t_5__661_;
  assign t_6__628_ = t_5__628_ | t_5__660_;
  assign t_6__627_ = t_5__627_ | t_5__659_;
  assign t_6__626_ = t_5__626_ | t_5__658_;
  assign t_6__625_ = t_5__625_ | t_5__657_;
  assign t_6__624_ = t_5__624_ | t_5__656_;
  assign t_6__623_ = t_5__623_ | t_5__655_;
  assign t_6__622_ = t_5__622_ | t_5__654_;
  assign t_6__621_ = t_5__621_ | t_5__653_;
  assign t_6__620_ = t_5__620_ | t_5__652_;
  assign t_6__619_ = t_5__619_ | t_5__651_;
  assign t_6__618_ = t_5__618_ | t_5__650_;
  assign t_6__617_ = t_5__617_ | t_5__649_;
  assign t_6__616_ = t_5__616_ | t_5__648_;
  assign t_6__615_ = t_5__615_ | t_5__647_;
  assign t_6__614_ = t_5__614_ | t_5__646_;
  assign t_6__613_ = t_5__613_ | t_5__645_;
  assign t_6__612_ = t_5__612_ | t_5__644_;
  assign t_6__611_ = t_5__611_ | t_5__643_;
  assign t_6__610_ = t_5__610_ | t_5__642_;
  assign t_6__609_ = t_5__609_ | t_5__641_;
  assign t_6__608_ = t_5__608_ | t_5__640_;
  assign t_6__607_ = t_5__607_ | t_5__639_;
  assign t_6__606_ = t_5__606_ | t_5__638_;
  assign t_6__605_ = t_5__605_ | t_5__637_;
  assign t_6__604_ = t_5__604_ | t_5__636_;
  assign t_6__603_ = t_5__603_ | t_5__635_;
  assign t_6__602_ = t_5__602_ | t_5__634_;
  assign t_6__601_ = t_5__601_ | t_5__633_;
  assign t_6__600_ = t_5__600_ | t_5__632_;
  assign t_6__599_ = t_5__599_ | t_5__631_;
  assign t_6__598_ = t_5__598_ | t_5__630_;
  assign t_6__597_ = t_5__597_ | t_5__629_;
  assign t_6__596_ = t_5__596_ | t_5__628_;
  assign t_6__595_ = t_5__595_ | t_5__627_;
  assign t_6__594_ = t_5__594_ | t_5__626_;
  assign t_6__593_ = t_5__593_ | t_5__625_;
  assign t_6__592_ = t_5__592_ | t_5__624_;
  assign t_6__591_ = t_5__591_ | t_5__623_;
  assign t_6__590_ = t_5__590_ | t_5__622_;
  assign t_6__589_ = t_5__589_ | t_5__621_;
  assign t_6__588_ = t_5__588_ | t_5__620_;
  assign t_6__587_ = t_5__587_ | t_5__619_;
  assign t_6__586_ = t_5__586_ | t_5__618_;
  assign t_6__585_ = t_5__585_ | t_5__617_;
  assign t_6__584_ = t_5__584_ | t_5__616_;
  assign t_6__583_ = t_5__583_ | t_5__615_;
  assign t_6__582_ = t_5__582_ | t_5__614_;
  assign t_6__581_ = t_5__581_ | t_5__613_;
  assign t_6__580_ = t_5__580_ | t_5__612_;
  assign t_6__579_ = t_5__579_ | t_5__611_;
  assign t_6__578_ = t_5__578_ | t_5__610_;
  assign t_6__577_ = t_5__577_ | t_5__609_;
  assign t_6__576_ = t_5__576_ | t_5__608_;
  assign t_6__575_ = t_5__575_ | t_5__607_;
  assign t_6__574_ = t_5__574_ | t_5__606_;
  assign t_6__573_ = t_5__573_ | t_5__605_;
  assign t_6__572_ = t_5__572_ | t_5__604_;
  assign t_6__571_ = t_5__571_ | t_5__603_;
  assign t_6__570_ = t_5__570_ | t_5__602_;
  assign t_6__569_ = t_5__569_ | t_5__601_;
  assign t_6__568_ = t_5__568_ | t_5__600_;
  assign t_6__567_ = t_5__567_ | t_5__599_;
  assign t_6__566_ = t_5__566_ | t_5__598_;
  assign t_6__565_ = t_5__565_ | t_5__597_;
  assign t_6__564_ = t_5__564_ | t_5__596_;
  assign t_6__563_ = t_5__563_ | t_5__595_;
  assign t_6__562_ = t_5__562_ | t_5__594_;
  assign t_6__561_ = t_5__561_ | t_5__593_;
  assign t_6__560_ = t_5__560_ | t_5__592_;
  assign t_6__559_ = t_5__559_ | t_5__591_;
  assign t_6__558_ = t_5__558_ | t_5__590_;
  assign t_6__557_ = t_5__557_ | t_5__589_;
  assign t_6__556_ = t_5__556_ | t_5__588_;
  assign t_6__555_ = t_5__555_ | t_5__587_;
  assign t_6__554_ = t_5__554_ | t_5__586_;
  assign t_6__553_ = t_5__553_ | t_5__585_;
  assign t_6__552_ = t_5__552_ | t_5__584_;
  assign t_6__551_ = t_5__551_ | t_5__583_;
  assign t_6__550_ = t_5__550_ | t_5__582_;
  assign t_6__549_ = t_5__549_ | t_5__581_;
  assign t_6__548_ = t_5__548_ | t_5__580_;
  assign t_6__547_ = t_5__547_ | t_5__579_;
  assign t_6__546_ = t_5__546_ | t_5__578_;
  assign t_6__545_ = t_5__545_ | t_5__577_;
  assign t_6__544_ = t_5__544_ | t_5__576_;
  assign t_6__543_ = t_5__543_ | t_5__575_;
  assign t_6__542_ = t_5__542_ | t_5__574_;
  assign t_6__541_ = t_5__541_ | t_5__573_;
  assign t_6__540_ = t_5__540_ | t_5__572_;
  assign t_6__539_ = t_5__539_ | t_5__571_;
  assign t_6__538_ = t_5__538_ | t_5__570_;
  assign t_6__537_ = t_5__537_ | t_5__569_;
  assign t_6__536_ = t_5__536_ | t_5__568_;
  assign t_6__535_ = t_5__535_ | t_5__567_;
  assign t_6__534_ = t_5__534_ | t_5__566_;
  assign t_6__533_ = t_5__533_ | t_5__565_;
  assign t_6__532_ = t_5__532_ | t_5__564_;
  assign t_6__531_ = t_5__531_ | t_5__563_;
  assign t_6__530_ = t_5__530_ | t_5__562_;
  assign t_6__529_ = t_5__529_ | t_5__561_;
  assign t_6__528_ = t_5__528_ | t_5__560_;
  assign t_6__527_ = t_5__527_ | t_5__559_;
  assign t_6__526_ = t_5__526_ | t_5__558_;
  assign t_6__525_ = t_5__525_ | t_5__557_;
  assign t_6__524_ = t_5__524_ | t_5__556_;
  assign t_6__523_ = t_5__523_ | t_5__555_;
  assign t_6__522_ = t_5__522_ | t_5__554_;
  assign t_6__521_ = t_5__521_ | t_5__553_;
  assign t_6__520_ = t_5__520_ | t_5__552_;
  assign t_6__519_ = t_5__519_ | t_5__551_;
  assign t_6__518_ = t_5__518_ | t_5__550_;
  assign t_6__517_ = t_5__517_ | t_5__549_;
  assign t_6__516_ = t_5__516_ | t_5__548_;
  assign t_6__515_ = t_5__515_ | t_5__547_;
  assign t_6__514_ = t_5__514_ | t_5__546_;
  assign t_6__513_ = t_5__513_ | t_5__545_;
  assign t_6__512_ = t_5__512_ | t_5__544_;
  assign t_6__511_ = t_5__511_ | t_5__543_;
  assign t_6__510_ = t_5__510_ | t_5__542_;
  assign t_6__509_ = t_5__509_ | t_5__541_;
  assign t_6__508_ = t_5__508_ | t_5__540_;
  assign t_6__507_ = t_5__507_ | t_5__539_;
  assign t_6__506_ = t_5__506_ | t_5__538_;
  assign t_6__505_ = t_5__505_ | t_5__537_;
  assign t_6__504_ = t_5__504_ | t_5__536_;
  assign t_6__503_ = t_5__503_ | t_5__535_;
  assign t_6__502_ = t_5__502_ | t_5__534_;
  assign t_6__501_ = t_5__501_ | t_5__533_;
  assign t_6__500_ = t_5__500_ | t_5__532_;
  assign t_6__499_ = t_5__499_ | t_5__531_;
  assign t_6__498_ = t_5__498_ | t_5__530_;
  assign t_6__497_ = t_5__497_ | t_5__529_;
  assign t_6__496_ = t_5__496_ | t_5__528_;
  assign t_6__495_ = t_5__495_ | t_5__527_;
  assign t_6__494_ = t_5__494_ | t_5__526_;
  assign t_6__493_ = t_5__493_ | t_5__525_;
  assign t_6__492_ = t_5__492_ | t_5__524_;
  assign t_6__491_ = t_5__491_ | t_5__523_;
  assign t_6__490_ = t_5__490_ | t_5__522_;
  assign t_6__489_ = t_5__489_ | t_5__521_;
  assign t_6__488_ = t_5__488_ | t_5__520_;
  assign t_6__487_ = t_5__487_ | t_5__519_;
  assign t_6__486_ = t_5__486_ | t_5__518_;
  assign t_6__485_ = t_5__485_ | t_5__517_;
  assign t_6__484_ = t_5__484_ | t_5__516_;
  assign t_6__483_ = t_5__483_ | t_5__515_;
  assign t_6__482_ = t_5__482_ | t_5__514_;
  assign t_6__481_ = t_5__481_ | t_5__513_;
  assign t_6__480_ = t_5__480_ | t_5__512_;
  assign t_6__479_ = t_5__479_ | t_5__511_;
  assign t_6__478_ = t_5__478_ | t_5__510_;
  assign t_6__477_ = t_5__477_ | t_5__509_;
  assign t_6__476_ = t_5__476_ | t_5__508_;
  assign t_6__475_ = t_5__475_ | t_5__507_;
  assign t_6__474_ = t_5__474_ | t_5__506_;
  assign t_6__473_ = t_5__473_ | t_5__505_;
  assign t_6__472_ = t_5__472_ | t_5__504_;
  assign t_6__471_ = t_5__471_ | t_5__503_;
  assign t_6__470_ = t_5__470_ | t_5__502_;
  assign t_6__469_ = t_5__469_ | t_5__501_;
  assign t_6__468_ = t_5__468_ | t_5__500_;
  assign t_6__467_ = t_5__467_ | t_5__499_;
  assign t_6__466_ = t_5__466_ | t_5__498_;
  assign t_6__465_ = t_5__465_ | t_5__497_;
  assign t_6__464_ = t_5__464_ | t_5__496_;
  assign t_6__463_ = t_5__463_ | t_5__495_;
  assign t_6__462_ = t_5__462_ | t_5__494_;
  assign t_6__461_ = t_5__461_ | t_5__493_;
  assign t_6__460_ = t_5__460_ | t_5__492_;
  assign t_6__459_ = t_5__459_ | t_5__491_;
  assign t_6__458_ = t_5__458_ | t_5__490_;
  assign t_6__457_ = t_5__457_ | t_5__489_;
  assign t_6__456_ = t_5__456_ | t_5__488_;
  assign t_6__455_ = t_5__455_ | t_5__487_;
  assign t_6__454_ = t_5__454_ | t_5__486_;
  assign t_6__453_ = t_5__453_ | t_5__485_;
  assign t_6__452_ = t_5__452_ | t_5__484_;
  assign t_6__451_ = t_5__451_ | t_5__483_;
  assign t_6__450_ = t_5__450_ | t_5__482_;
  assign t_6__449_ = t_5__449_ | t_5__481_;
  assign t_6__448_ = t_5__448_ | t_5__480_;
  assign t_6__447_ = t_5__447_ | t_5__479_;
  assign t_6__446_ = t_5__446_ | t_5__478_;
  assign t_6__445_ = t_5__445_ | t_5__477_;
  assign t_6__444_ = t_5__444_ | t_5__476_;
  assign t_6__443_ = t_5__443_ | t_5__475_;
  assign t_6__442_ = t_5__442_ | t_5__474_;
  assign t_6__441_ = t_5__441_ | t_5__473_;
  assign t_6__440_ = t_5__440_ | t_5__472_;
  assign t_6__439_ = t_5__439_ | t_5__471_;
  assign t_6__438_ = t_5__438_ | t_5__470_;
  assign t_6__437_ = t_5__437_ | t_5__469_;
  assign t_6__436_ = t_5__436_ | t_5__468_;
  assign t_6__435_ = t_5__435_ | t_5__467_;
  assign t_6__434_ = t_5__434_ | t_5__466_;
  assign t_6__433_ = t_5__433_ | t_5__465_;
  assign t_6__432_ = t_5__432_ | t_5__464_;
  assign t_6__431_ = t_5__431_ | t_5__463_;
  assign t_6__430_ = t_5__430_ | t_5__462_;
  assign t_6__429_ = t_5__429_ | t_5__461_;
  assign t_6__428_ = t_5__428_ | t_5__460_;
  assign t_6__427_ = t_5__427_ | t_5__459_;
  assign t_6__426_ = t_5__426_ | t_5__458_;
  assign t_6__425_ = t_5__425_ | t_5__457_;
  assign t_6__424_ = t_5__424_ | t_5__456_;
  assign t_6__423_ = t_5__423_ | t_5__455_;
  assign t_6__422_ = t_5__422_ | t_5__454_;
  assign t_6__421_ = t_5__421_ | t_5__453_;
  assign t_6__420_ = t_5__420_ | t_5__452_;
  assign t_6__419_ = t_5__419_ | t_5__451_;
  assign t_6__418_ = t_5__418_ | t_5__450_;
  assign t_6__417_ = t_5__417_ | t_5__449_;
  assign t_6__416_ = t_5__416_ | t_5__448_;
  assign t_6__415_ = t_5__415_ | t_5__447_;
  assign t_6__414_ = t_5__414_ | t_5__446_;
  assign t_6__413_ = t_5__413_ | t_5__445_;
  assign t_6__412_ = t_5__412_ | t_5__444_;
  assign t_6__411_ = t_5__411_ | t_5__443_;
  assign t_6__410_ = t_5__410_ | t_5__442_;
  assign t_6__409_ = t_5__409_ | t_5__441_;
  assign t_6__408_ = t_5__408_ | t_5__440_;
  assign t_6__407_ = t_5__407_ | t_5__439_;
  assign t_6__406_ = t_5__406_ | t_5__438_;
  assign t_6__405_ = t_5__405_ | t_5__437_;
  assign t_6__404_ = t_5__404_ | t_5__436_;
  assign t_6__403_ = t_5__403_ | t_5__435_;
  assign t_6__402_ = t_5__402_ | t_5__434_;
  assign t_6__401_ = t_5__401_ | t_5__433_;
  assign t_6__400_ = t_5__400_ | t_5__432_;
  assign t_6__399_ = t_5__399_ | t_5__431_;
  assign t_6__398_ = t_5__398_ | t_5__430_;
  assign t_6__397_ = t_5__397_ | t_5__429_;
  assign t_6__396_ = t_5__396_ | t_5__428_;
  assign t_6__395_ = t_5__395_ | t_5__427_;
  assign t_6__394_ = t_5__394_ | t_5__426_;
  assign t_6__393_ = t_5__393_ | t_5__425_;
  assign t_6__392_ = t_5__392_ | t_5__424_;
  assign t_6__391_ = t_5__391_ | t_5__423_;
  assign t_6__390_ = t_5__390_ | t_5__422_;
  assign t_6__389_ = t_5__389_ | t_5__421_;
  assign t_6__388_ = t_5__388_ | t_5__420_;
  assign t_6__387_ = t_5__387_ | t_5__419_;
  assign t_6__386_ = t_5__386_ | t_5__418_;
  assign t_6__385_ = t_5__385_ | t_5__417_;
  assign t_6__384_ = t_5__384_ | t_5__416_;
  assign t_6__383_ = t_5__383_ | t_5__415_;
  assign t_6__382_ = t_5__382_ | t_5__414_;
  assign t_6__381_ = t_5__381_ | t_5__413_;
  assign t_6__380_ = t_5__380_ | t_5__412_;
  assign t_6__379_ = t_5__379_ | t_5__411_;
  assign t_6__378_ = t_5__378_ | t_5__410_;
  assign t_6__377_ = t_5__377_ | t_5__409_;
  assign t_6__376_ = t_5__376_ | t_5__408_;
  assign t_6__375_ = t_5__375_ | t_5__407_;
  assign t_6__374_ = t_5__374_ | t_5__406_;
  assign t_6__373_ = t_5__373_ | t_5__405_;
  assign t_6__372_ = t_5__372_ | t_5__404_;
  assign t_6__371_ = t_5__371_ | t_5__403_;
  assign t_6__370_ = t_5__370_ | t_5__402_;
  assign t_6__369_ = t_5__369_ | t_5__401_;
  assign t_6__368_ = t_5__368_ | t_5__400_;
  assign t_6__367_ = t_5__367_ | t_5__399_;
  assign t_6__366_ = t_5__366_ | t_5__398_;
  assign t_6__365_ = t_5__365_ | t_5__397_;
  assign t_6__364_ = t_5__364_ | t_5__396_;
  assign t_6__363_ = t_5__363_ | t_5__395_;
  assign t_6__362_ = t_5__362_ | t_5__394_;
  assign t_6__361_ = t_5__361_ | t_5__393_;
  assign t_6__360_ = t_5__360_ | t_5__392_;
  assign t_6__359_ = t_5__359_ | t_5__391_;
  assign t_6__358_ = t_5__358_ | t_5__390_;
  assign t_6__357_ = t_5__357_ | t_5__389_;
  assign t_6__356_ = t_5__356_ | t_5__388_;
  assign t_6__355_ = t_5__355_ | t_5__387_;
  assign t_6__354_ = t_5__354_ | t_5__386_;
  assign t_6__353_ = t_5__353_ | t_5__385_;
  assign t_6__352_ = t_5__352_ | t_5__384_;
  assign t_6__351_ = t_5__351_ | t_5__383_;
  assign t_6__350_ = t_5__350_ | t_5__382_;
  assign t_6__349_ = t_5__349_ | t_5__381_;
  assign t_6__348_ = t_5__348_ | t_5__380_;
  assign t_6__347_ = t_5__347_ | t_5__379_;
  assign t_6__346_ = t_5__346_ | t_5__378_;
  assign t_6__345_ = t_5__345_ | t_5__377_;
  assign t_6__344_ = t_5__344_ | t_5__376_;
  assign t_6__343_ = t_5__343_ | t_5__375_;
  assign t_6__342_ = t_5__342_ | t_5__374_;
  assign t_6__341_ = t_5__341_ | t_5__373_;
  assign t_6__340_ = t_5__340_ | t_5__372_;
  assign t_6__339_ = t_5__339_ | t_5__371_;
  assign t_6__338_ = t_5__338_ | t_5__370_;
  assign t_6__337_ = t_5__337_ | t_5__369_;
  assign t_6__336_ = t_5__336_ | t_5__368_;
  assign t_6__335_ = t_5__335_ | t_5__367_;
  assign t_6__334_ = t_5__334_ | t_5__366_;
  assign t_6__333_ = t_5__333_ | t_5__365_;
  assign t_6__332_ = t_5__332_ | t_5__364_;
  assign t_6__331_ = t_5__331_ | t_5__363_;
  assign t_6__330_ = t_5__330_ | t_5__362_;
  assign t_6__329_ = t_5__329_ | t_5__361_;
  assign t_6__328_ = t_5__328_ | t_5__360_;
  assign t_6__327_ = t_5__327_ | t_5__359_;
  assign t_6__326_ = t_5__326_ | t_5__358_;
  assign t_6__325_ = t_5__325_ | t_5__357_;
  assign t_6__324_ = t_5__324_ | t_5__356_;
  assign t_6__323_ = t_5__323_ | t_5__355_;
  assign t_6__322_ = t_5__322_ | t_5__354_;
  assign t_6__321_ = t_5__321_ | t_5__353_;
  assign t_6__320_ = t_5__320_ | t_5__352_;
  assign t_6__319_ = t_5__319_ | t_5__351_;
  assign t_6__318_ = t_5__318_ | t_5__350_;
  assign t_6__317_ = t_5__317_ | t_5__349_;
  assign t_6__316_ = t_5__316_ | t_5__348_;
  assign t_6__315_ = t_5__315_ | t_5__347_;
  assign t_6__314_ = t_5__314_ | t_5__346_;
  assign t_6__313_ = t_5__313_ | t_5__345_;
  assign t_6__312_ = t_5__312_ | t_5__344_;
  assign t_6__311_ = t_5__311_ | t_5__343_;
  assign t_6__310_ = t_5__310_ | t_5__342_;
  assign t_6__309_ = t_5__309_ | t_5__341_;
  assign t_6__308_ = t_5__308_ | t_5__340_;
  assign t_6__307_ = t_5__307_ | t_5__339_;
  assign t_6__306_ = t_5__306_ | t_5__338_;
  assign t_6__305_ = t_5__305_ | t_5__337_;
  assign t_6__304_ = t_5__304_ | t_5__336_;
  assign t_6__303_ = t_5__303_ | t_5__335_;
  assign t_6__302_ = t_5__302_ | t_5__334_;
  assign t_6__301_ = t_5__301_ | t_5__333_;
  assign t_6__300_ = t_5__300_ | t_5__332_;
  assign t_6__299_ = t_5__299_ | t_5__331_;
  assign t_6__298_ = t_5__298_ | t_5__330_;
  assign t_6__297_ = t_5__297_ | t_5__329_;
  assign t_6__296_ = t_5__296_ | t_5__328_;
  assign t_6__295_ = t_5__295_ | t_5__327_;
  assign t_6__294_ = t_5__294_ | t_5__326_;
  assign t_6__293_ = t_5__293_ | t_5__325_;
  assign t_6__292_ = t_5__292_ | t_5__324_;
  assign t_6__291_ = t_5__291_ | t_5__323_;
  assign t_6__290_ = t_5__290_ | t_5__322_;
  assign t_6__289_ = t_5__289_ | t_5__321_;
  assign t_6__288_ = t_5__288_ | t_5__320_;
  assign t_6__287_ = t_5__287_ | t_5__319_;
  assign t_6__286_ = t_5__286_ | t_5__318_;
  assign t_6__285_ = t_5__285_ | t_5__317_;
  assign t_6__284_ = t_5__284_ | t_5__316_;
  assign t_6__283_ = t_5__283_ | t_5__315_;
  assign t_6__282_ = t_5__282_ | t_5__314_;
  assign t_6__281_ = t_5__281_ | t_5__313_;
  assign t_6__280_ = t_5__280_ | t_5__312_;
  assign t_6__279_ = t_5__279_ | t_5__311_;
  assign t_6__278_ = t_5__278_ | t_5__310_;
  assign t_6__277_ = t_5__277_ | t_5__309_;
  assign t_6__276_ = t_5__276_ | t_5__308_;
  assign t_6__275_ = t_5__275_ | t_5__307_;
  assign t_6__274_ = t_5__274_ | t_5__306_;
  assign t_6__273_ = t_5__273_ | t_5__305_;
  assign t_6__272_ = t_5__272_ | t_5__304_;
  assign t_6__271_ = t_5__271_ | t_5__303_;
  assign t_6__270_ = t_5__270_ | t_5__302_;
  assign t_6__269_ = t_5__269_ | t_5__301_;
  assign t_6__268_ = t_5__268_ | t_5__300_;
  assign t_6__267_ = t_5__267_ | t_5__299_;
  assign t_6__266_ = t_5__266_ | t_5__298_;
  assign t_6__265_ = t_5__265_ | t_5__297_;
  assign t_6__264_ = t_5__264_ | t_5__296_;
  assign t_6__263_ = t_5__263_ | t_5__295_;
  assign t_6__262_ = t_5__262_ | t_5__294_;
  assign t_6__261_ = t_5__261_ | t_5__293_;
  assign t_6__260_ = t_5__260_ | t_5__292_;
  assign t_6__259_ = t_5__259_ | t_5__291_;
  assign t_6__258_ = t_5__258_ | t_5__290_;
  assign t_6__257_ = t_5__257_ | t_5__289_;
  assign t_6__256_ = t_5__256_ | t_5__288_;
  assign t_6__255_ = t_5__255_ | t_5__287_;
  assign t_6__254_ = t_5__254_ | t_5__286_;
  assign t_6__253_ = t_5__253_ | t_5__285_;
  assign t_6__252_ = t_5__252_ | t_5__284_;
  assign t_6__251_ = t_5__251_ | t_5__283_;
  assign t_6__250_ = t_5__250_ | t_5__282_;
  assign t_6__249_ = t_5__249_ | t_5__281_;
  assign t_6__248_ = t_5__248_ | t_5__280_;
  assign t_6__247_ = t_5__247_ | t_5__279_;
  assign t_6__246_ = t_5__246_ | t_5__278_;
  assign t_6__245_ = t_5__245_ | t_5__277_;
  assign t_6__244_ = t_5__244_ | t_5__276_;
  assign t_6__243_ = t_5__243_ | t_5__275_;
  assign t_6__242_ = t_5__242_ | t_5__274_;
  assign t_6__241_ = t_5__241_ | t_5__273_;
  assign t_6__240_ = t_5__240_ | t_5__272_;
  assign t_6__239_ = t_5__239_ | t_5__271_;
  assign t_6__238_ = t_5__238_ | t_5__270_;
  assign t_6__237_ = t_5__237_ | t_5__269_;
  assign t_6__236_ = t_5__236_ | t_5__268_;
  assign t_6__235_ = t_5__235_ | t_5__267_;
  assign t_6__234_ = t_5__234_ | t_5__266_;
  assign t_6__233_ = t_5__233_ | t_5__265_;
  assign t_6__232_ = t_5__232_ | t_5__264_;
  assign t_6__231_ = t_5__231_ | t_5__263_;
  assign t_6__230_ = t_5__230_ | t_5__262_;
  assign t_6__229_ = t_5__229_ | t_5__261_;
  assign t_6__228_ = t_5__228_ | t_5__260_;
  assign t_6__227_ = t_5__227_ | t_5__259_;
  assign t_6__226_ = t_5__226_ | t_5__258_;
  assign t_6__225_ = t_5__225_ | t_5__257_;
  assign t_6__224_ = t_5__224_ | t_5__256_;
  assign t_6__223_ = t_5__223_ | t_5__255_;
  assign t_6__222_ = t_5__222_ | t_5__254_;
  assign t_6__221_ = t_5__221_ | t_5__253_;
  assign t_6__220_ = t_5__220_ | t_5__252_;
  assign t_6__219_ = t_5__219_ | t_5__251_;
  assign t_6__218_ = t_5__218_ | t_5__250_;
  assign t_6__217_ = t_5__217_ | t_5__249_;
  assign t_6__216_ = t_5__216_ | t_5__248_;
  assign t_6__215_ = t_5__215_ | t_5__247_;
  assign t_6__214_ = t_5__214_ | t_5__246_;
  assign t_6__213_ = t_5__213_ | t_5__245_;
  assign t_6__212_ = t_5__212_ | t_5__244_;
  assign t_6__211_ = t_5__211_ | t_5__243_;
  assign t_6__210_ = t_5__210_ | t_5__242_;
  assign t_6__209_ = t_5__209_ | t_5__241_;
  assign t_6__208_ = t_5__208_ | t_5__240_;
  assign t_6__207_ = t_5__207_ | t_5__239_;
  assign t_6__206_ = t_5__206_ | t_5__238_;
  assign t_6__205_ = t_5__205_ | t_5__237_;
  assign t_6__204_ = t_5__204_ | t_5__236_;
  assign t_6__203_ = t_5__203_ | t_5__235_;
  assign t_6__202_ = t_5__202_ | t_5__234_;
  assign t_6__201_ = t_5__201_ | t_5__233_;
  assign t_6__200_ = t_5__200_ | t_5__232_;
  assign t_6__199_ = t_5__199_ | t_5__231_;
  assign t_6__198_ = t_5__198_ | t_5__230_;
  assign t_6__197_ = t_5__197_ | t_5__229_;
  assign t_6__196_ = t_5__196_ | t_5__228_;
  assign t_6__195_ = t_5__195_ | t_5__227_;
  assign t_6__194_ = t_5__194_ | t_5__226_;
  assign t_6__193_ = t_5__193_ | t_5__225_;
  assign t_6__192_ = t_5__192_ | t_5__224_;
  assign t_6__191_ = t_5__191_ | t_5__223_;
  assign t_6__190_ = t_5__190_ | t_5__222_;
  assign t_6__189_ = t_5__189_ | t_5__221_;
  assign t_6__188_ = t_5__188_ | t_5__220_;
  assign t_6__187_ = t_5__187_ | t_5__219_;
  assign t_6__186_ = t_5__186_ | t_5__218_;
  assign t_6__185_ = t_5__185_ | t_5__217_;
  assign t_6__184_ = t_5__184_ | t_5__216_;
  assign t_6__183_ = t_5__183_ | t_5__215_;
  assign t_6__182_ = t_5__182_ | t_5__214_;
  assign t_6__181_ = t_5__181_ | t_5__213_;
  assign t_6__180_ = t_5__180_ | t_5__212_;
  assign t_6__179_ = t_5__179_ | t_5__211_;
  assign t_6__178_ = t_5__178_ | t_5__210_;
  assign t_6__177_ = t_5__177_ | t_5__209_;
  assign t_6__176_ = t_5__176_ | t_5__208_;
  assign t_6__175_ = t_5__175_ | t_5__207_;
  assign t_6__174_ = t_5__174_ | t_5__206_;
  assign t_6__173_ = t_5__173_ | t_5__205_;
  assign t_6__172_ = t_5__172_ | t_5__204_;
  assign t_6__171_ = t_5__171_ | t_5__203_;
  assign t_6__170_ = t_5__170_ | t_5__202_;
  assign t_6__169_ = t_5__169_ | t_5__201_;
  assign t_6__168_ = t_5__168_ | t_5__200_;
  assign t_6__167_ = t_5__167_ | t_5__199_;
  assign t_6__166_ = t_5__166_ | t_5__198_;
  assign t_6__165_ = t_5__165_ | t_5__197_;
  assign t_6__164_ = t_5__164_ | t_5__196_;
  assign t_6__163_ = t_5__163_ | t_5__195_;
  assign t_6__162_ = t_5__162_ | t_5__194_;
  assign t_6__161_ = t_5__161_ | t_5__193_;
  assign t_6__160_ = t_5__160_ | t_5__192_;
  assign t_6__159_ = t_5__159_ | t_5__191_;
  assign t_6__158_ = t_5__158_ | t_5__190_;
  assign t_6__157_ = t_5__157_ | t_5__189_;
  assign t_6__156_ = t_5__156_ | t_5__188_;
  assign t_6__155_ = t_5__155_ | t_5__187_;
  assign t_6__154_ = t_5__154_ | t_5__186_;
  assign t_6__153_ = t_5__153_ | t_5__185_;
  assign t_6__152_ = t_5__152_ | t_5__184_;
  assign t_6__151_ = t_5__151_ | t_5__183_;
  assign t_6__150_ = t_5__150_ | t_5__182_;
  assign t_6__149_ = t_5__149_ | t_5__181_;
  assign t_6__148_ = t_5__148_ | t_5__180_;
  assign t_6__147_ = t_5__147_ | t_5__179_;
  assign t_6__146_ = t_5__146_ | t_5__178_;
  assign t_6__145_ = t_5__145_ | t_5__177_;
  assign t_6__144_ = t_5__144_ | t_5__176_;
  assign t_6__143_ = t_5__143_ | t_5__175_;
  assign t_6__142_ = t_5__142_ | t_5__174_;
  assign t_6__141_ = t_5__141_ | t_5__173_;
  assign t_6__140_ = t_5__140_ | t_5__172_;
  assign t_6__139_ = t_5__139_ | t_5__171_;
  assign t_6__138_ = t_5__138_ | t_5__170_;
  assign t_6__137_ = t_5__137_ | t_5__169_;
  assign t_6__136_ = t_5__136_ | t_5__168_;
  assign t_6__135_ = t_5__135_ | t_5__167_;
  assign t_6__134_ = t_5__134_ | t_5__166_;
  assign t_6__133_ = t_5__133_ | t_5__165_;
  assign t_6__132_ = t_5__132_ | t_5__164_;
  assign t_6__131_ = t_5__131_ | t_5__163_;
  assign t_6__130_ = t_5__130_ | t_5__162_;
  assign t_6__129_ = t_5__129_ | t_5__161_;
  assign t_6__128_ = t_5__128_ | t_5__160_;
  assign t_6__127_ = t_5__127_ | t_5__159_;
  assign t_6__126_ = t_5__126_ | t_5__158_;
  assign t_6__125_ = t_5__125_ | t_5__157_;
  assign t_6__124_ = t_5__124_ | t_5__156_;
  assign t_6__123_ = t_5__123_ | t_5__155_;
  assign t_6__122_ = t_5__122_ | t_5__154_;
  assign t_6__121_ = t_5__121_ | t_5__153_;
  assign t_6__120_ = t_5__120_ | t_5__152_;
  assign t_6__119_ = t_5__119_ | t_5__151_;
  assign t_6__118_ = t_5__118_ | t_5__150_;
  assign t_6__117_ = t_5__117_ | t_5__149_;
  assign t_6__116_ = t_5__116_ | t_5__148_;
  assign t_6__115_ = t_5__115_ | t_5__147_;
  assign t_6__114_ = t_5__114_ | t_5__146_;
  assign t_6__113_ = t_5__113_ | t_5__145_;
  assign t_6__112_ = t_5__112_ | t_5__144_;
  assign t_6__111_ = t_5__111_ | t_5__143_;
  assign t_6__110_ = t_5__110_ | t_5__142_;
  assign t_6__109_ = t_5__109_ | t_5__141_;
  assign t_6__108_ = t_5__108_ | t_5__140_;
  assign t_6__107_ = t_5__107_ | t_5__139_;
  assign t_6__106_ = t_5__106_ | t_5__138_;
  assign t_6__105_ = t_5__105_ | t_5__137_;
  assign t_6__104_ = t_5__104_ | t_5__136_;
  assign t_6__103_ = t_5__103_ | t_5__135_;
  assign t_6__102_ = t_5__102_ | t_5__134_;
  assign t_6__101_ = t_5__101_ | t_5__133_;
  assign t_6__100_ = t_5__100_ | t_5__132_;
  assign t_6__99_ = t_5__99_ | t_5__131_;
  assign t_6__98_ = t_5__98_ | t_5__130_;
  assign t_6__97_ = t_5__97_ | t_5__129_;
  assign t_6__96_ = t_5__96_ | t_5__128_;
  assign t_6__95_ = t_5__95_ | t_5__127_;
  assign t_6__94_ = t_5__94_ | t_5__126_;
  assign t_6__93_ = t_5__93_ | t_5__125_;
  assign t_6__92_ = t_5__92_ | t_5__124_;
  assign t_6__91_ = t_5__91_ | t_5__123_;
  assign t_6__90_ = t_5__90_ | t_5__122_;
  assign t_6__89_ = t_5__89_ | t_5__121_;
  assign t_6__88_ = t_5__88_ | t_5__120_;
  assign t_6__87_ = t_5__87_ | t_5__119_;
  assign t_6__86_ = t_5__86_ | t_5__118_;
  assign t_6__85_ = t_5__85_ | t_5__117_;
  assign t_6__84_ = t_5__84_ | t_5__116_;
  assign t_6__83_ = t_5__83_ | t_5__115_;
  assign t_6__82_ = t_5__82_ | t_5__114_;
  assign t_6__81_ = t_5__81_ | t_5__113_;
  assign t_6__80_ = t_5__80_ | t_5__112_;
  assign t_6__79_ = t_5__79_ | t_5__111_;
  assign t_6__78_ = t_5__78_ | t_5__110_;
  assign t_6__77_ = t_5__77_ | t_5__109_;
  assign t_6__76_ = t_5__76_ | t_5__108_;
  assign t_6__75_ = t_5__75_ | t_5__107_;
  assign t_6__74_ = t_5__74_ | t_5__106_;
  assign t_6__73_ = t_5__73_ | t_5__105_;
  assign t_6__72_ = t_5__72_ | t_5__104_;
  assign t_6__71_ = t_5__71_ | t_5__103_;
  assign t_6__70_ = t_5__70_ | t_5__102_;
  assign t_6__69_ = t_5__69_ | t_5__101_;
  assign t_6__68_ = t_5__68_ | t_5__100_;
  assign t_6__67_ = t_5__67_ | t_5__99_;
  assign t_6__66_ = t_5__66_ | t_5__98_;
  assign t_6__65_ = t_5__65_ | t_5__97_;
  assign t_6__64_ = t_5__64_ | t_5__96_;
  assign t_6__63_ = t_5__63_ | t_5__95_;
  assign t_6__62_ = t_5__62_ | t_5__94_;
  assign t_6__61_ = t_5__61_ | t_5__93_;
  assign t_6__60_ = t_5__60_ | t_5__92_;
  assign t_6__59_ = t_5__59_ | t_5__91_;
  assign t_6__58_ = t_5__58_ | t_5__90_;
  assign t_6__57_ = t_5__57_ | t_5__89_;
  assign t_6__56_ = t_5__56_ | t_5__88_;
  assign t_6__55_ = t_5__55_ | t_5__87_;
  assign t_6__54_ = t_5__54_ | t_5__86_;
  assign t_6__53_ = t_5__53_ | t_5__85_;
  assign t_6__52_ = t_5__52_ | t_5__84_;
  assign t_6__51_ = t_5__51_ | t_5__83_;
  assign t_6__50_ = t_5__50_ | t_5__82_;
  assign t_6__49_ = t_5__49_ | t_5__81_;
  assign t_6__48_ = t_5__48_ | t_5__80_;
  assign t_6__47_ = t_5__47_ | t_5__79_;
  assign t_6__46_ = t_5__46_ | t_5__78_;
  assign t_6__45_ = t_5__45_ | t_5__77_;
  assign t_6__44_ = t_5__44_ | t_5__76_;
  assign t_6__43_ = t_5__43_ | t_5__75_;
  assign t_6__42_ = t_5__42_ | t_5__74_;
  assign t_6__41_ = t_5__41_ | t_5__73_;
  assign t_6__40_ = t_5__40_ | t_5__72_;
  assign t_6__39_ = t_5__39_ | t_5__71_;
  assign t_6__38_ = t_5__38_ | t_5__70_;
  assign t_6__37_ = t_5__37_ | t_5__69_;
  assign t_6__36_ = t_5__36_ | t_5__68_;
  assign t_6__35_ = t_5__35_ | t_5__67_;
  assign t_6__34_ = t_5__34_ | t_5__66_;
  assign t_6__33_ = t_5__33_ | t_5__65_;
  assign t_6__32_ = t_5__32_ | t_5__64_;
  assign t_6__31_ = t_5__31_ | t_5__63_;
  assign t_6__30_ = t_5__30_ | t_5__62_;
  assign t_6__29_ = t_5__29_ | t_5__61_;
  assign t_6__28_ = t_5__28_ | t_5__60_;
  assign t_6__27_ = t_5__27_ | t_5__59_;
  assign t_6__26_ = t_5__26_ | t_5__58_;
  assign t_6__25_ = t_5__25_ | t_5__57_;
  assign t_6__24_ = t_5__24_ | t_5__56_;
  assign t_6__23_ = t_5__23_ | t_5__55_;
  assign t_6__22_ = t_5__22_ | t_5__54_;
  assign t_6__21_ = t_5__21_ | t_5__53_;
  assign t_6__20_ = t_5__20_ | t_5__52_;
  assign t_6__19_ = t_5__19_ | t_5__51_;
  assign t_6__18_ = t_5__18_ | t_5__50_;
  assign t_6__17_ = t_5__17_ | t_5__49_;
  assign t_6__16_ = t_5__16_ | t_5__48_;
  assign t_6__15_ = t_5__15_ | t_5__47_;
  assign t_6__14_ = t_5__14_ | t_5__46_;
  assign t_6__13_ = t_5__13_ | t_5__45_;
  assign t_6__12_ = t_5__12_ | t_5__44_;
  assign t_6__11_ = t_5__11_ | t_5__43_;
  assign t_6__10_ = t_5__10_ | t_5__42_;
  assign t_6__9_ = t_5__9_ | t_5__41_;
  assign t_6__8_ = t_5__8_ | t_5__40_;
  assign t_6__7_ = t_5__7_ | t_5__39_;
  assign t_6__6_ = t_5__6_ | t_5__38_;
  assign t_6__5_ = t_5__5_ | t_5__37_;
  assign t_6__4_ = t_5__4_ | t_5__36_;
  assign t_6__3_ = t_5__3_ | t_5__35_;
  assign t_6__2_ = t_5__2_ | t_5__34_;
  assign t_6__1_ = t_5__1_ | t_5__33_;
  assign t_6__0_ = t_5__0_ | t_5__32_;
  assign t_7__1023_ = t_6__1023_ | 1'b0;
  assign t_7__1022_ = t_6__1022_ | 1'b0;
  assign t_7__1021_ = t_6__1021_ | 1'b0;
  assign t_7__1020_ = t_6__1020_ | 1'b0;
  assign t_7__1019_ = t_6__1019_ | 1'b0;
  assign t_7__1018_ = t_6__1018_ | 1'b0;
  assign t_7__1017_ = t_6__1017_ | 1'b0;
  assign t_7__1016_ = t_6__1016_ | 1'b0;
  assign t_7__1015_ = t_6__1015_ | 1'b0;
  assign t_7__1014_ = t_6__1014_ | 1'b0;
  assign t_7__1013_ = t_6__1013_ | 1'b0;
  assign t_7__1012_ = t_6__1012_ | 1'b0;
  assign t_7__1011_ = t_6__1011_ | 1'b0;
  assign t_7__1010_ = t_6__1010_ | 1'b0;
  assign t_7__1009_ = t_6__1009_ | 1'b0;
  assign t_7__1008_ = t_6__1008_ | 1'b0;
  assign t_7__1007_ = t_6__1007_ | 1'b0;
  assign t_7__1006_ = t_6__1006_ | 1'b0;
  assign t_7__1005_ = t_6__1005_ | 1'b0;
  assign t_7__1004_ = t_6__1004_ | 1'b0;
  assign t_7__1003_ = t_6__1003_ | 1'b0;
  assign t_7__1002_ = t_6__1002_ | 1'b0;
  assign t_7__1001_ = t_6__1001_ | 1'b0;
  assign t_7__1000_ = t_6__1000_ | 1'b0;
  assign t_7__999_ = t_6__999_ | 1'b0;
  assign t_7__998_ = t_6__998_ | 1'b0;
  assign t_7__997_ = t_6__997_ | 1'b0;
  assign t_7__996_ = t_6__996_ | 1'b0;
  assign t_7__995_ = t_6__995_ | 1'b0;
  assign t_7__994_ = t_6__994_ | 1'b0;
  assign t_7__993_ = t_6__993_ | 1'b0;
  assign t_7__992_ = t_6__992_ | 1'b0;
  assign t_7__991_ = t_6__991_ | 1'b0;
  assign t_7__990_ = t_6__990_ | 1'b0;
  assign t_7__989_ = t_6__989_ | 1'b0;
  assign t_7__988_ = t_6__988_ | 1'b0;
  assign t_7__987_ = t_6__987_ | 1'b0;
  assign t_7__986_ = t_6__986_ | 1'b0;
  assign t_7__985_ = t_6__985_ | 1'b0;
  assign t_7__984_ = t_6__984_ | 1'b0;
  assign t_7__983_ = t_6__983_ | 1'b0;
  assign t_7__982_ = t_6__982_ | 1'b0;
  assign t_7__981_ = t_6__981_ | 1'b0;
  assign t_7__980_ = t_6__980_ | 1'b0;
  assign t_7__979_ = t_6__979_ | 1'b0;
  assign t_7__978_ = t_6__978_ | 1'b0;
  assign t_7__977_ = t_6__977_ | 1'b0;
  assign t_7__976_ = t_6__976_ | 1'b0;
  assign t_7__975_ = t_6__975_ | 1'b0;
  assign t_7__974_ = t_6__974_ | 1'b0;
  assign t_7__973_ = t_6__973_ | 1'b0;
  assign t_7__972_ = t_6__972_ | 1'b0;
  assign t_7__971_ = t_6__971_ | 1'b0;
  assign t_7__970_ = t_6__970_ | 1'b0;
  assign t_7__969_ = t_6__969_ | 1'b0;
  assign t_7__968_ = t_6__968_ | 1'b0;
  assign t_7__967_ = t_6__967_ | 1'b0;
  assign t_7__966_ = t_6__966_ | 1'b0;
  assign t_7__965_ = t_6__965_ | 1'b0;
  assign t_7__964_ = t_6__964_ | 1'b0;
  assign t_7__963_ = t_6__963_ | 1'b0;
  assign t_7__962_ = t_6__962_ | 1'b0;
  assign t_7__961_ = t_6__961_ | 1'b0;
  assign t_7__960_ = t_6__960_ | 1'b0;
  assign t_7__959_ = t_6__959_ | t_6__1023_;
  assign t_7__958_ = t_6__958_ | t_6__1022_;
  assign t_7__957_ = t_6__957_ | t_6__1021_;
  assign t_7__956_ = t_6__956_ | t_6__1020_;
  assign t_7__955_ = t_6__955_ | t_6__1019_;
  assign t_7__954_ = t_6__954_ | t_6__1018_;
  assign t_7__953_ = t_6__953_ | t_6__1017_;
  assign t_7__952_ = t_6__952_ | t_6__1016_;
  assign t_7__951_ = t_6__951_ | t_6__1015_;
  assign t_7__950_ = t_6__950_ | t_6__1014_;
  assign t_7__949_ = t_6__949_ | t_6__1013_;
  assign t_7__948_ = t_6__948_ | t_6__1012_;
  assign t_7__947_ = t_6__947_ | t_6__1011_;
  assign t_7__946_ = t_6__946_ | t_6__1010_;
  assign t_7__945_ = t_6__945_ | t_6__1009_;
  assign t_7__944_ = t_6__944_ | t_6__1008_;
  assign t_7__943_ = t_6__943_ | t_6__1007_;
  assign t_7__942_ = t_6__942_ | t_6__1006_;
  assign t_7__941_ = t_6__941_ | t_6__1005_;
  assign t_7__940_ = t_6__940_ | t_6__1004_;
  assign t_7__939_ = t_6__939_ | t_6__1003_;
  assign t_7__938_ = t_6__938_ | t_6__1002_;
  assign t_7__937_ = t_6__937_ | t_6__1001_;
  assign t_7__936_ = t_6__936_ | t_6__1000_;
  assign t_7__935_ = t_6__935_ | t_6__999_;
  assign t_7__934_ = t_6__934_ | t_6__998_;
  assign t_7__933_ = t_6__933_ | t_6__997_;
  assign t_7__932_ = t_6__932_ | t_6__996_;
  assign t_7__931_ = t_6__931_ | t_6__995_;
  assign t_7__930_ = t_6__930_ | t_6__994_;
  assign t_7__929_ = t_6__929_ | t_6__993_;
  assign t_7__928_ = t_6__928_ | t_6__992_;
  assign t_7__927_ = t_6__927_ | t_6__991_;
  assign t_7__926_ = t_6__926_ | t_6__990_;
  assign t_7__925_ = t_6__925_ | t_6__989_;
  assign t_7__924_ = t_6__924_ | t_6__988_;
  assign t_7__923_ = t_6__923_ | t_6__987_;
  assign t_7__922_ = t_6__922_ | t_6__986_;
  assign t_7__921_ = t_6__921_ | t_6__985_;
  assign t_7__920_ = t_6__920_ | t_6__984_;
  assign t_7__919_ = t_6__919_ | t_6__983_;
  assign t_7__918_ = t_6__918_ | t_6__982_;
  assign t_7__917_ = t_6__917_ | t_6__981_;
  assign t_7__916_ = t_6__916_ | t_6__980_;
  assign t_7__915_ = t_6__915_ | t_6__979_;
  assign t_7__914_ = t_6__914_ | t_6__978_;
  assign t_7__913_ = t_6__913_ | t_6__977_;
  assign t_7__912_ = t_6__912_ | t_6__976_;
  assign t_7__911_ = t_6__911_ | t_6__975_;
  assign t_7__910_ = t_6__910_ | t_6__974_;
  assign t_7__909_ = t_6__909_ | t_6__973_;
  assign t_7__908_ = t_6__908_ | t_6__972_;
  assign t_7__907_ = t_6__907_ | t_6__971_;
  assign t_7__906_ = t_6__906_ | t_6__970_;
  assign t_7__905_ = t_6__905_ | t_6__969_;
  assign t_7__904_ = t_6__904_ | t_6__968_;
  assign t_7__903_ = t_6__903_ | t_6__967_;
  assign t_7__902_ = t_6__902_ | t_6__966_;
  assign t_7__901_ = t_6__901_ | t_6__965_;
  assign t_7__900_ = t_6__900_ | t_6__964_;
  assign t_7__899_ = t_6__899_ | t_6__963_;
  assign t_7__898_ = t_6__898_ | t_6__962_;
  assign t_7__897_ = t_6__897_ | t_6__961_;
  assign t_7__896_ = t_6__896_ | t_6__960_;
  assign t_7__895_ = t_6__895_ | t_6__959_;
  assign t_7__894_ = t_6__894_ | t_6__958_;
  assign t_7__893_ = t_6__893_ | t_6__957_;
  assign t_7__892_ = t_6__892_ | t_6__956_;
  assign t_7__891_ = t_6__891_ | t_6__955_;
  assign t_7__890_ = t_6__890_ | t_6__954_;
  assign t_7__889_ = t_6__889_ | t_6__953_;
  assign t_7__888_ = t_6__888_ | t_6__952_;
  assign t_7__887_ = t_6__887_ | t_6__951_;
  assign t_7__886_ = t_6__886_ | t_6__950_;
  assign t_7__885_ = t_6__885_ | t_6__949_;
  assign t_7__884_ = t_6__884_ | t_6__948_;
  assign t_7__883_ = t_6__883_ | t_6__947_;
  assign t_7__882_ = t_6__882_ | t_6__946_;
  assign t_7__881_ = t_6__881_ | t_6__945_;
  assign t_7__880_ = t_6__880_ | t_6__944_;
  assign t_7__879_ = t_6__879_ | t_6__943_;
  assign t_7__878_ = t_6__878_ | t_6__942_;
  assign t_7__877_ = t_6__877_ | t_6__941_;
  assign t_7__876_ = t_6__876_ | t_6__940_;
  assign t_7__875_ = t_6__875_ | t_6__939_;
  assign t_7__874_ = t_6__874_ | t_6__938_;
  assign t_7__873_ = t_6__873_ | t_6__937_;
  assign t_7__872_ = t_6__872_ | t_6__936_;
  assign t_7__871_ = t_6__871_ | t_6__935_;
  assign t_7__870_ = t_6__870_ | t_6__934_;
  assign t_7__869_ = t_6__869_ | t_6__933_;
  assign t_7__868_ = t_6__868_ | t_6__932_;
  assign t_7__867_ = t_6__867_ | t_6__931_;
  assign t_7__866_ = t_6__866_ | t_6__930_;
  assign t_7__865_ = t_6__865_ | t_6__929_;
  assign t_7__864_ = t_6__864_ | t_6__928_;
  assign t_7__863_ = t_6__863_ | t_6__927_;
  assign t_7__862_ = t_6__862_ | t_6__926_;
  assign t_7__861_ = t_6__861_ | t_6__925_;
  assign t_7__860_ = t_6__860_ | t_6__924_;
  assign t_7__859_ = t_6__859_ | t_6__923_;
  assign t_7__858_ = t_6__858_ | t_6__922_;
  assign t_7__857_ = t_6__857_ | t_6__921_;
  assign t_7__856_ = t_6__856_ | t_6__920_;
  assign t_7__855_ = t_6__855_ | t_6__919_;
  assign t_7__854_ = t_6__854_ | t_6__918_;
  assign t_7__853_ = t_6__853_ | t_6__917_;
  assign t_7__852_ = t_6__852_ | t_6__916_;
  assign t_7__851_ = t_6__851_ | t_6__915_;
  assign t_7__850_ = t_6__850_ | t_6__914_;
  assign t_7__849_ = t_6__849_ | t_6__913_;
  assign t_7__848_ = t_6__848_ | t_6__912_;
  assign t_7__847_ = t_6__847_ | t_6__911_;
  assign t_7__846_ = t_6__846_ | t_6__910_;
  assign t_7__845_ = t_6__845_ | t_6__909_;
  assign t_7__844_ = t_6__844_ | t_6__908_;
  assign t_7__843_ = t_6__843_ | t_6__907_;
  assign t_7__842_ = t_6__842_ | t_6__906_;
  assign t_7__841_ = t_6__841_ | t_6__905_;
  assign t_7__840_ = t_6__840_ | t_6__904_;
  assign t_7__839_ = t_6__839_ | t_6__903_;
  assign t_7__838_ = t_6__838_ | t_6__902_;
  assign t_7__837_ = t_6__837_ | t_6__901_;
  assign t_7__836_ = t_6__836_ | t_6__900_;
  assign t_7__835_ = t_6__835_ | t_6__899_;
  assign t_7__834_ = t_6__834_ | t_6__898_;
  assign t_7__833_ = t_6__833_ | t_6__897_;
  assign t_7__832_ = t_6__832_ | t_6__896_;
  assign t_7__831_ = t_6__831_ | t_6__895_;
  assign t_7__830_ = t_6__830_ | t_6__894_;
  assign t_7__829_ = t_6__829_ | t_6__893_;
  assign t_7__828_ = t_6__828_ | t_6__892_;
  assign t_7__827_ = t_6__827_ | t_6__891_;
  assign t_7__826_ = t_6__826_ | t_6__890_;
  assign t_7__825_ = t_6__825_ | t_6__889_;
  assign t_7__824_ = t_6__824_ | t_6__888_;
  assign t_7__823_ = t_6__823_ | t_6__887_;
  assign t_7__822_ = t_6__822_ | t_6__886_;
  assign t_7__821_ = t_6__821_ | t_6__885_;
  assign t_7__820_ = t_6__820_ | t_6__884_;
  assign t_7__819_ = t_6__819_ | t_6__883_;
  assign t_7__818_ = t_6__818_ | t_6__882_;
  assign t_7__817_ = t_6__817_ | t_6__881_;
  assign t_7__816_ = t_6__816_ | t_6__880_;
  assign t_7__815_ = t_6__815_ | t_6__879_;
  assign t_7__814_ = t_6__814_ | t_6__878_;
  assign t_7__813_ = t_6__813_ | t_6__877_;
  assign t_7__812_ = t_6__812_ | t_6__876_;
  assign t_7__811_ = t_6__811_ | t_6__875_;
  assign t_7__810_ = t_6__810_ | t_6__874_;
  assign t_7__809_ = t_6__809_ | t_6__873_;
  assign t_7__808_ = t_6__808_ | t_6__872_;
  assign t_7__807_ = t_6__807_ | t_6__871_;
  assign t_7__806_ = t_6__806_ | t_6__870_;
  assign t_7__805_ = t_6__805_ | t_6__869_;
  assign t_7__804_ = t_6__804_ | t_6__868_;
  assign t_7__803_ = t_6__803_ | t_6__867_;
  assign t_7__802_ = t_6__802_ | t_6__866_;
  assign t_7__801_ = t_6__801_ | t_6__865_;
  assign t_7__800_ = t_6__800_ | t_6__864_;
  assign t_7__799_ = t_6__799_ | t_6__863_;
  assign t_7__798_ = t_6__798_ | t_6__862_;
  assign t_7__797_ = t_6__797_ | t_6__861_;
  assign t_7__796_ = t_6__796_ | t_6__860_;
  assign t_7__795_ = t_6__795_ | t_6__859_;
  assign t_7__794_ = t_6__794_ | t_6__858_;
  assign t_7__793_ = t_6__793_ | t_6__857_;
  assign t_7__792_ = t_6__792_ | t_6__856_;
  assign t_7__791_ = t_6__791_ | t_6__855_;
  assign t_7__790_ = t_6__790_ | t_6__854_;
  assign t_7__789_ = t_6__789_ | t_6__853_;
  assign t_7__788_ = t_6__788_ | t_6__852_;
  assign t_7__787_ = t_6__787_ | t_6__851_;
  assign t_7__786_ = t_6__786_ | t_6__850_;
  assign t_7__785_ = t_6__785_ | t_6__849_;
  assign t_7__784_ = t_6__784_ | t_6__848_;
  assign t_7__783_ = t_6__783_ | t_6__847_;
  assign t_7__782_ = t_6__782_ | t_6__846_;
  assign t_7__781_ = t_6__781_ | t_6__845_;
  assign t_7__780_ = t_6__780_ | t_6__844_;
  assign t_7__779_ = t_6__779_ | t_6__843_;
  assign t_7__778_ = t_6__778_ | t_6__842_;
  assign t_7__777_ = t_6__777_ | t_6__841_;
  assign t_7__776_ = t_6__776_ | t_6__840_;
  assign t_7__775_ = t_6__775_ | t_6__839_;
  assign t_7__774_ = t_6__774_ | t_6__838_;
  assign t_7__773_ = t_6__773_ | t_6__837_;
  assign t_7__772_ = t_6__772_ | t_6__836_;
  assign t_7__771_ = t_6__771_ | t_6__835_;
  assign t_7__770_ = t_6__770_ | t_6__834_;
  assign t_7__769_ = t_6__769_ | t_6__833_;
  assign t_7__768_ = t_6__768_ | t_6__832_;
  assign t_7__767_ = t_6__767_ | t_6__831_;
  assign t_7__766_ = t_6__766_ | t_6__830_;
  assign t_7__765_ = t_6__765_ | t_6__829_;
  assign t_7__764_ = t_6__764_ | t_6__828_;
  assign t_7__763_ = t_6__763_ | t_6__827_;
  assign t_7__762_ = t_6__762_ | t_6__826_;
  assign t_7__761_ = t_6__761_ | t_6__825_;
  assign t_7__760_ = t_6__760_ | t_6__824_;
  assign t_7__759_ = t_6__759_ | t_6__823_;
  assign t_7__758_ = t_6__758_ | t_6__822_;
  assign t_7__757_ = t_6__757_ | t_6__821_;
  assign t_7__756_ = t_6__756_ | t_6__820_;
  assign t_7__755_ = t_6__755_ | t_6__819_;
  assign t_7__754_ = t_6__754_ | t_6__818_;
  assign t_7__753_ = t_6__753_ | t_6__817_;
  assign t_7__752_ = t_6__752_ | t_6__816_;
  assign t_7__751_ = t_6__751_ | t_6__815_;
  assign t_7__750_ = t_6__750_ | t_6__814_;
  assign t_7__749_ = t_6__749_ | t_6__813_;
  assign t_7__748_ = t_6__748_ | t_6__812_;
  assign t_7__747_ = t_6__747_ | t_6__811_;
  assign t_7__746_ = t_6__746_ | t_6__810_;
  assign t_7__745_ = t_6__745_ | t_6__809_;
  assign t_7__744_ = t_6__744_ | t_6__808_;
  assign t_7__743_ = t_6__743_ | t_6__807_;
  assign t_7__742_ = t_6__742_ | t_6__806_;
  assign t_7__741_ = t_6__741_ | t_6__805_;
  assign t_7__740_ = t_6__740_ | t_6__804_;
  assign t_7__739_ = t_6__739_ | t_6__803_;
  assign t_7__738_ = t_6__738_ | t_6__802_;
  assign t_7__737_ = t_6__737_ | t_6__801_;
  assign t_7__736_ = t_6__736_ | t_6__800_;
  assign t_7__735_ = t_6__735_ | t_6__799_;
  assign t_7__734_ = t_6__734_ | t_6__798_;
  assign t_7__733_ = t_6__733_ | t_6__797_;
  assign t_7__732_ = t_6__732_ | t_6__796_;
  assign t_7__731_ = t_6__731_ | t_6__795_;
  assign t_7__730_ = t_6__730_ | t_6__794_;
  assign t_7__729_ = t_6__729_ | t_6__793_;
  assign t_7__728_ = t_6__728_ | t_6__792_;
  assign t_7__727_ = t_6__727_ | t_6__791_;
  assign t_7__726_ = t_6__726_ | t_6__790_;
  assign t_7__725_ = t_6__725_ | t_6__789_;
  assign t_7__724_ = t_6__724_ | t_6__788_;
  assign t_7__723_ = t_6__723_ | t_6__787_;
  assign t_7__722_ = t_6__722_ | t_6__786_;
  assign t_7__721_ = t_6__721_ | t_6__785_;
  assign t_7__720_ = t_6__720_ | t_6__784_;
  assign t_7__719_ = t_6__719_ | t_6__783_;
  assign t_7__718_ = t_6__718_ | t_6__782_;
  assign t_7__717_ = t_6__717_ | t_6__781_;
  assign t_7__716_ = t_6__716_ | t_6__780_;
  assign t_7__715_ = t_6__715_ | t_6__779_;
  assign t_7__714_ = t_6__714_ | t_6__778_;
  assign t_7__713_ = t_6__713_ | t_6__777_;
  assign t_7__712_ = t_6__712_ | t_6__776_;
  assign t_7__711_ = t_6__711_ | t_6__775_;
  assign t_7__710_ = t_6__710_ | t_6__774_;
  assign t_7__709_ = t_6__709_ | t_6__773_;
  assign t_7__708_ = t_6__708_ | t_6__772_;
  assign t_7__707_ = t_6__707_ | t_6__771_;
  assign t_7__706_ = t_6__706_ | t_6__770_;
  assign t_7__705_ = t_6__705_ | t_6__769_;
  assign t_7__704_ = t_6__704_ | t_6__768_;
  assign t_7__703_ = t_6__703_ | t_6__767_;
  assign t_7__702_ = t_6__702_ | t_6__766_;
  assign t_7__701_ = t_6__701_ | t_6__765_;
  assign t_7__700_ = t_6__700_ | t_6__764_;
  assign t_7__699_ = t_6__699_ | t_6__763_;
  assign t_7__698_ = t_6__698_ | t_6__762_;
  assign t_7__697_ = t_6__697_ | t_6__761_;
  assign t_7__696_ = t_6__696_ | t_6__760_;
  assign t_7__695_ = t_6__695_ | t_6__759_;
  assign t_7__694_ = t_6__694_ | t_6__758_;
  assign t_7__693_ = t_6__693_ | t_6__757_;
  assign t_7__692_ = t_6__692_ | t_6__756_;
  assign t_7__691_ = t_6__691_ | t_6__755_;
  assign t_7__690_ = t_6__690_ | t_6__754_;
  assign t_7__689_ = t_6__689_ | t_6__753_;
  assign t_7__688_ = t_6__688_ | t_6__752_;
  assign t_7__687_ = t_6__687_ | t_6__751_;
  assign t_7__686_ = t_6__686_ | t_6__750_;
  assign t_7__685_ = t_6__685_ | t_6__749_;
  assign t_7__684_ = t_6__684_ | t_6__748_;
  assign t_7__683_ = t_6__683_ | t_6__747_;
  assign t_7__682_ = t_6__682_ | t_6__746_;
  assign t_7__681_ = t_6__681_ | t_6__745_;
  assign t_7__680_ = t_6__680_ | t_6__744_;
  assign t_7__679_ = t_6__679_ | t_6__743_;
  assign t_7__678_ = t_6__678_ | t_6__742_;
  assign t_7__677_ = t_6__677_ | t_6__741_;
  assign t_7__676_ = t_6__676_ | t_6__740_;
  assign t_7__675_ = t_6__675_ | t_6__739_;
  assign t_7__674_ = t_6__674_ | t_6__738_;
  assign t_7__673_ = t_6__673_ | t_6__737_;
  assign t_7__672_ = t_6__672_ | t_6__736_;
  assign t_7__671_ = t_6__671_ | t_6__735_;
  assign t_7__670_ = t_6__670_ | t_6__734_;
  assign t_7__669_ = t_6__669_ | t_6__733_;
  assign t_7__668_ = t_6__668_ | t_6__732_;
  assign t_7__667_ = t_6__667_ | t_6__731_;
  assign t_7__666_ = t_6__666_ | t_6__730_;
  assign t_7__665_ = t_6__665_ | t_6__729_;
  assign t_7__664_ = t_6__664_ | t_6__728_;
  assign t_7__663_ = t_6__663_ | t_6__727_;
  assign t_7__662_ = t_6__662_ | t_6__726_;
  assign t_7__661_ = t_6__661_ | t_6__725_;
  assign t_7__660_ = t_6__660_ | t_6__724_;
  assign t_7__659_ = t_6__659_ | t_6__723_;
  assign t_7__658_ = t_6__658_ | t_6__722_;
  assign t_7__657_ = t_6__657_ | t_6__721_;
  assign t_7__656_ = t_6__656_ | t_6__720_;
  assign t_7__655_ = t_6__655_ | t_6__719_;
  assign t_7__654_ = t_6__654_ | t_6__718_;
  assign t_7__653_ = t_6__653_ | t_6__717_;
  assign t_7__652_ = t_6__652_ | t_6__716_;
  assign t_7__651_ = t_6__651_ | t_6__715_;
  assign t_7__650_ = t_6__650_ | t_6__714_;
  assign t_7__649_ = t_6__649_ | t_6__713_;
  assign t_7__648_ = t_6__648_ | t_6__712_;
  assign t_7__647_ = t_6__647_ | t_6__711_;
  assign t_7__646_ = t_6__646_ | t_6__710_;
  assign t_7__645_ = t_6__645_ | t_6__709_;
  assign t_7__644_ = t_6__644_ | t_6__708_;
  assign t_7__643_ = t_6__643_ | t_6__707_;
  assign t_7__642_ = t_6__642_ | t_6__706_;
  assign t_7__641_ = t_6__641_ | t_6__705_;
  assign t_7__640_ = t_6__640_ | t_6__704_;
  assign t_7__639_ = t_6__639_ | t_6__703_;
  assign t_7__638_ = t_6__638_ | t_6__702_;
  assign t_7__637_ = t_6__637_ | t_6__701_;
  assign t_7__636_ = t_6__636_ | t_6__700_;
  assign t_7__635_ = t_6__635_ | t_6__699_;
  assign t_7__634_ = t_6__634_ | t_6__698_;
  assign t_7__633_ = t_6__633_ | t_6__697_;
  assign t_7__632_ = t_6__632_ | t_6__696_;
  assign t_7__631_ = t_6__631_ | t_6__695_;
  assign t_7__630_ = t_6__630_ | t_6__694_;
  assign t_7__629_ = t_6__629_ | t_6__693_;
  assign t_7__628_ = t_6__628_ | t_6__692_;
  assign t_7__627_ = t_6__627_ | t_6__691_;
  assign t_7__626_ = t_6__626_ | t_6__690_;
  assign t_7__625_ = t_6__625_ | t_6__689_;
  assign t_7__624_ = t_6__624_ | t_6__688_;
  assign t_7__623_ = t_6__623_ | t_6__687_;
  assign t_7__622_ = t_6__622_ | t_6__686_;
  assign t_7__621_ = t_6__621_ | t_6__685_;
  assign t_7__620_ = t_6__620_ | t_6__684_;
  assign t_7__619_ = t_6__619_ | t_6__683_;
  assign t_7__618_ = t_6__618_ | t_6__682_;
  assign t_7__617_ = t_6__617_ | t_6__681_;
  assign t_7__616_ = t_6__616_ | t_6__680_;
  assign t_7__615_ = t_6__615_ | t_6__679_;
  assign t_7__614_ = t_6__614_ | t_6__678_;
  assign t_7__613_ = t_6__613_ | t_6__677_;
  assign t_7__612_ = t_6__612_ | t_6__676_;
  assign t_7__611_ = t_6__611_ | t_6__675_;
  assign t_7__610_ = t_6__610_ | t_6__674_;
  assign t_7__609_ = t_6__609_ | t_6__673_;
  assign t_7__608_ = t_6__608_ | t_6__672_;
  assign t_7__607_ = t_6__607_ | t_6__671_;
  assign t_7__606_ = t_6__606_ | t_6__670_;
  assign t_7__605_ = t_6__605_ | t_6__669_;
  assign t_7__604_ = t_6__604_ | t_6__668_;
  assign t_7__603_ = t_6__603_ | t_6__667_;
  assign t_7__602_ = t_6__602_ | t_6__666_;
  assign t_7__601_ = t_6__601_ | t_6__665_;
  assign t_7__600_ = t_6__600_ | t_6__664_;
  assign t_7__599_ = t_6__599_ | t_6__663_;
  assign t_7__598_ = t_6__598_ | t_6__662_;
  assign t_7__597_ = t_6__597_ | t_6__661_;
  assign t_7__596_ = t_6__596_ | t_6__660_;
  assign t_7__595_ = t_6__595_ | t_6__659_;
  assign t_7__594_ = t_6__594_ | t_6__658_;
  assign t_7__593_ = t_6__593_ | t_6__657_;
  assign t_7__592_ = t_6__592_ | t_6__656_;
  assign t_7__591_ = t_6__591_ | t_6__655_;
  assign t_7__590_ = t_6__590_ | t_6__654_;
  assign t_7__589_ = t_6__589_ | t_6__653_;
  assign t_7__588_ = t_6__588_ | t_6__652_;
  assign t_7__587_ = t_6__587_ | t_6__651_;
  assign t_7__586_ = t_6__586_ | t_6__650_;
  assign t_7__585_ = t_6__585_ | t_6__649_;
  assign t_7__584_ = t_6__584_ | t_6__648_;
  assign t_7__583_ = t_6__583_ | t_6__647_;
  assign t_7__582_ = t_6__582_ | t_6__646_;
  assign t_7__581_ = t_6__581_ | t_6__645_;
  assign t_7__580_ = t_6__580_ | t_6__644_;
  assign t_7__579_ = t_6__579_ | t_6__643_;
  assign t_7__578_ = t_6__578_ | t_6__642_;
  assign t_7__577_ = t_6__577_ | t_6__641_;
  assign t_7__576_ = t_6__576_ | t_6__640_;
  assign t_7__575_ = t_6__575_ | t_6__639_;
  assign t_7__574_ = t_6__574_ | t_6__638_;
  assign t_7__573_ = t_6__573_ | t_6__637_;
  assign t_7__572_ = t_6__572_ | t_6__636_;
  assign t_7__571_ = t_6__571_ | t_6__635_;
  assign t_7__570_ = t_6__570_ | t_6__634_;
  assign t_7__569_ = t_6__569_ | t_6__633_;
  assign t_7__568_ = t_6__568_ | t_6__632_;
  assign t_7__567_ = t_6__567_ | t_6__631_;
  assign t_7__566_ = t_6__566_ | t_6__630_;
  assign t_7__565_ = t_6__565_ | t_6__629_;
  assign t_7__564_ = t_6__564_ | t_6__628_;
  assign t_7__563_ = t_6__563_ | t_6__627_;
  assign t_7__562_ = t_6__562_ | t_6__626_;
  assign t_7__561_ = t_6__561_ | t_6__625_;
  assign t_7__560_ = t_6__560_ | t_6__624_;
  assign t_7__559_ = t_6__559_ | t_6__623_;
  assign t_7__558_ = t_6__558_ | t_6__622_;
  assign t_7__557_ = t_6__557_ | t_6__621_;
  assign t_7__556_ = t_6__556_ | t_6__620_;
  assign t_7__555_ = t_6__555_ | t_6__619_;
  assign t_7__554_ = t_6__554_ | t_6__618_;
  assign t_7__553_ = t_6__553_ | t_6__617_;
  assign t_7__552_ = t_6__552_ | t_6__616_;
  assign t_7__551_ = t_6__551_ | t_6__615_;
  assign t_7__550_ = t_6__550_ | t_6__614_;
  assign t_7__549_ = t_6__549_ | t_6__613_;
  assign t_7__548_ = t_6__548_ | t_6__612_;
  assign t_7__547_ = t_6__547_ | t_6__611_;
  assign t_7__546_ = t_6__546_ | t_6__610_;
  assign t_7__545_ = t_6__545_ | t_6__609_;
  assign t_7__544_ = t_6__544_ | t_6__608_;
  assign t_7__543_ = t_6__543_ | t_6__607_;
  assign t_7__542_ = t_6__542_ | t_6__606_;
  assign t_7__541_ = t_6__541_ | t_6__605_;
  assign t_7__540_ = t_6__540_ | t_6__604_;
  assign t_7__539_ = t_6__539_ | t_6__603_;
  assign t_7__538_ = t_6__538_ | t_6__602_;
  assign t_7__537_ = t_6__537_ | t_6__601_;
  assign t_7__536_ = t_6__536_ | t_6__600_;
  assign t_7__535_ = t_6__535_ | t_6__599_;
  assign t_7__534_ = t_6__534_ | t_6__598_;
  assign t_7__533_ = t_6__533_ | t_6__597_;
  assign t_7__532_ = t_6__532_ | t_6__596_;
  assign t_7__531_ = t_6__531_ | t_6__595_;
  assign t_7__530_ = t_6__530_ | t_6__594_;
  assign t_7__529_ = t_6__529_ | t_6__593_;
  assign t_7__528_ = t_6__528_ | t_6__592_;
  assign t_7__527_ = t_6__527_ | t_6__591_;
  assign t_7__526_ = t_6__526_ | t_6__590_;
  assign t_7__525_ = t_6__525_ | t_6__589_;
  assign t_7__524_ = t_6__524_ | t_6__588_;
  assign t_7__523_ = t_6__523_ | t_6__587_;
  assign t_7__522_ = t_6__522_ | t_6__586_;
  assign t_7__521_ = t_6__521_ | t_6__585_;
  assign t_7__520_ = t_6__520_ | t_6__584_;
  assign t_7__519_ = t_6__519_ | t_6__583_;
  assign t_7__518_ = t_6__518_ | t_6__582_;
  assign t_7__517_ = t_6__517_ | t_6__581_;
  assign t_7__516_ = t_6__516_ | t_6__580_;
  assign t_7__515_ = t_6__515_ | t_6__579_;
  assign t_7__514_ = t_6__514_ | t_6__578_;
  assign t_7__513_ = t_6__513_ | t_6__577_;
  assign t_7__512_ = t_6__512_ | t_6__576_;
  assign t_7__511_ = t_6__511_ | t_6__575_;
  assign t_7__510_ = t_6__510_ | t_6__574_;
  assign t_7__509_ = t_6__509_ | t_6__573_;
  assign t_7__508_ = t_6__508_ | t_6__572_;
  assign t_7__507_ = t_6__507_ | t_6__571_;
  assign t_7__506_ = t_6__506_ | t_6__570_;
  assign t_7__505_ = t_6__505_ | t_6__569_;
  assign t_7__504_ = t_6__504_ | t_6__568_;
  assign t_7__503_ = t_6__503_ | t_6__567_;
  assign t_7__502_ = t_6__502_ | t_6__566_;
  assign t_7__501_ = t_6__501_ | t_6__565_;
  assign t_7__500_ = t_6__500_ | t_6__564_;
  assign t_7__499_ = t_6__499_ | t_6__563_;
  assign t_7__498_ = t_6__498_ | t_6__562_;
  assign t_7__497_ = t_6__497_ | t_6__561_;
  assign t_7__496_ = t_6__496_ | t_6__560_;
  assign t_7__495_ = t_6__495_ | t_6__559_;
  assign t_7__494_ = t_6__494_ | t_6__558_;
  assign t_7__493_ = t_6__493_ | t_6__557_;
  assign t_7__492_ = t_6__492_ | t_6__556_;
  assign t_7__491_ = t_6__491_ | t_6__555_;
  assign t_7__490_ = t_6__490_ | t_6__554_;
  assign t_7__489_ = t_6__489_ | t_6__553_;
  assign t_7__488_ = t_6__488_ | t_6__552_;
  assign t_7__487_ = t_6__487_ | t_6__551_;
  assign t_7__486_ = t_6__486_ | t_6__550_;
  assign t_7__485_ = t_6__485_ | t_6__549_;
  assign t_7__484_ = t_6__484_ | t_6__548_;
  assign t_7__483_ = t_6__483_ | t_6__547_;
  assign t_7__482_ = t_6__482_ | t_6__546_;
  assign t_7__481_ = t_6__481_ | t_6__545_;
  assign t_7__480_ = t_6__480_ | t_6__544_;
  assign t_7__479_ = t_6__479_ | t_6__543_;
  assign t_7__478_ = t_6__478_ | t_6__542_;
  assign t_7__477_ = t_6__477_ | t_6__541_;
  assign t_7__476_ = t_6__476_ | t_6__540_;
  assign t_7__475_ = t_6__475_ | t_6__539_;
  assign t_7__474_ = t_6__474_ | t_6__538_;
  assign t_7__473_ = t_6__473_ | t_6__537_;
  assign t_7__472_ = t_6__472_ | t_6__536_;
  assign t_7__471_ = t_6__471_ | t_6__535_;
  assign t_7__470_ = t_6__470_ | t_6__534_;
  assign t_7__469_ = t_6__469_ | t_6__533_;
  assign t_7__468_ = t_6__468_ | t_6__532_;
  assign t_7__467_ = t_6__467_ | t_6__531_;
  assign t_7__466_ = t_6__466_ | t_6__530_;
  assign t_7__465_ = t_6__465_ | t_6__529_;
  assign t_7__464_ = t_6__464_ | t_6__528_;
  assign t_7__463_ = t_6__463_ | t_6__527_;
  assign t_7__462_ = t_6__462_ | t_6__526_;
  assign t_7__461_ = t_6__461_ | t_6__525_;
  assign t_7__460_ = t_6__460_ | t_6__524_;
  assign t_7__459_ = t_6__459_ | t_6__523_;
  assign t_7__458_ = t_6__458_ | t_6__522_;
  assign t_7__457_ = t_6__457_ | t_6__521_;
  assign t_7__456_ = t_6__456_ | t_6__520_;
  assign t_7__455_ = t_6__455_ | t_6__519_;
  assign t_7__454_ = t_6__454_ | t_6__518_;
  assign t_7__453_ = t_6__453_ | t_6__517_;
  assign t_7__452_ = t_6__452_ | t_6__516_;
  assign t_7__451_ = t_6__451_ | t_6__515_;
  assign t_7__450_ = t_6__450_ | t_6__514_;
  assign t_7__449_ = t_6__449_ | t_6__513_;
  assign t_7__448_ = t_6__448_ | t_6__512_;
  assign t_7__447_ = t_6__447_ | t_6__511_;
  assign t_7__446_ = t_6__446_ | t_6__510_;
  assign t_7__445_ = t_6__445_ | t_6__509_;
  assign t_7__444_ = t_6__444_ | t_6__508_;
  assign t_7__443_ = t_6__443_ | t_6__507_;
  assign t_7__442_ = t_6__442_ | t_6__506_;
  assign t_7__441_ = t_6__441_ | t_6__505_;
  assign t_7__440_ = t_6__440_ | t_6__504_;
  assign t_7__439_ = t_6__439_ | t_6__503_;
  assign t_7__438_ = t_6__438_ | t_6__502_;
  assign t_7__437_ = t_6__437_ | t_6__501_;
  assign t_7__436_ = t_6__436_ | t_6__500_;
  assign t_7__435_ = t_6__435_ | t_6__499_;
  assign t_7__434_ = t_6__434_ | t_6__498_;
  assign t_7__433_ = t_6__433_ | t_6__497_;
  assign t_7__432_ = t_6__432_ | t_6__496_;
  assign t_7__431_ = t_6__431_ | t_6__495_;
  assign t_7__430_ = t_6__430_ | t_6__494_;
  assign t_7__429_ = t_6__429_ | t_6__493_;
  assign t_7__428_ = t_6__428_ | t_6__492_;
  assign t_7__427_ = t_6__427_ | t_6__491_;
  assign t_7__426_ = t_6__426_ | t_6__490_;
  assign t_7__425_ = t_6__425_ | t_6__489_;
  assign t_7__424_ = t_6__424_ | t_6__488_;
  assign t_7__423_ = t_6__423_ | t_6__487_;
  assign t_7__422_ = t_6__422_ | t_6__486_;
  assign t_7__421_ = t_6__421_ | t_6__485_;
  assign t_7__420_ = t_6__420_ | t_6__484_;
  assign t_7__419_ = t_6__419_ | t_6__483_;
  assign t_7__418_ = t_6__418_ | t_6__482_;
  assign t_7__417_ = t_6__417_ | t_6__481_;
  assign t_7__416_ = t_6__416_ | t_6__480_;
  assign t_7__415_ = t_6__415_ | t_6__479_;
  assign t_7__414_ = t_6__414_ | t_6__478_;
  assign t_7__413_ = t_6__413_ | t_6__477_;
  assign t_7__412_ = t_6__412_ | t_6__476_;
  assign t_7__411_ = t_6__411_ | t_6__475_;
  assign t_7__410_ = t_6__410_ | t_6__474_;
  assign t_7__409_ = t_6__409_ | t_6__473_;
  assign t_7__408_ = t_6__408_ | t_6__472_;
  assign t_7__407_ = t_6__407_ | t_6__471_;
  assign t_7__406_ = t_6__406_ | t_6__470_;
  assign t_7__405_ = t_6__405_ | t_6__469_;
  assign t_7__404_ = t_6__404_ | t_6__468_;
  assign t_7__403_ = t_6__403_ | t_6__467_;
  assign t_7__402_ = t_6__402_ | t_6__466_;
  assign t_7__401_ = t_6__401_ | t_6__465_;
  assign t_7__400_ = t_6__400_ | t_6__464_;
  assign t_7__399_ = t_6__399_ | t_6__463_;
  assign t_7__398_ = t_6__398_ | t_6__462_;
  assign t_7__397_ = t_6__397_ | t_6__461_;
  assign t_7__396_ = t_6__396_ | t_6__460_;
  assign t_7__395_ = t_6__395_ | t_6__459_;
  assign t_7__394_ = t_6__394_ | t_6__458_;
  assign t_7__393_ = t_6__393_ | t_6__457_;
  assign t_7__392_ = t_6__392_ | t_6__456_;
  assign t_7__391_ = t_6__391_ | t_6__455_;
  assign t_7__390_ = t_6__390_ | t_6__454_;
  assign t_7__389_ = t_6__389_ | t_6__453_;
  assign t_7__388_ = t_6__388_ | t_6__452_;
  assign t_7__387_ = t_6__387_ | t_6__451_;
  assign t_7__386_ = t_6__386_ | t_6__450_;
  assign t_7__385_ = t_6__385_ | t_6__449_;
  assign t_7__384_ = t_6__384_ | t_6__448_;
  assign t_7__383_ = t_6__383_ | t_6__447_;
  assign t_7__382_ = t_6__382_ | t_6__446_;
  assign t_7__381_ = t_6__381_ | t_6__445_;
  assign t_7__380_ = t_6__380_ | t_6__444_;
  assign t_7__379_ = t_6__379_ | t_6__443_;
  assign t_7__378_ = t_6__378_ | t_6__442_;
  assign t_7__377_ = t_6__377_ | t_6__441_;
  assign t_7__376_ = t_6__376_ | t_6__440_;
  assign t_7__375_ = t_6__375_ | t_6__439_;
  assign t_7__374_ = t_6__374_ | t_6__438_;
  assign t_7__373_ = t_6__373_ | t_6__437_;
  assign t_7__372_ = t_6__372_ | t_6__436_;
  assign t_7__371_ = t_6__371_ | t_6__435_;
  assign t_7__370_ = t_6__370_ | t_6__434_;
  assign t_7__369_ = t_6__369_ | t_6__433_;
  assign t_7__368_ = t_6__368_ | t_6__432_;
  assign t_7__367_ = t_6__367_ | t_6__431_;
  assign t_7__366_ = t_6__366_ | t_6__430_;
  assign t_7__365_ = t_6__365_ | t_6__429_;
  assign t_7__364_ = t_6__364_ | t_6__428_;
  assign t_7__363_ = t_6__363_ | t_6__427_;
  assign t_7__362_ = t_6__362_ | t_6__426_;
  assign t_7__361_ = t_6__361_ | t_6__425_;
  assign t_7__360_ = t_6__360_ | t_6__424_;
  assign t_7__359_ = t_6__359_ | t_6__423_;
  assign t_7__358_ = t_6__358_ | t_6__422_;
  assign t_7__357_ = t_6__357_ | t_6__421_;
  assign t_7__356_ = t_6__356_ | t_6__420_;
  assign t_7__355_ = t_6__355_ | t_6__419_;
  assign t_7__354_ = t_6__354_ | t_6__418_;
  assign t_7__353_ = t_6__353_ | t_6__417_;
  assign t_7__352_ = t_6__352_ | t_6__416_;
  assign t_7__351_ = t_6__351_ | t_6__415_;
  assign t_7__350_ = t_6__350_ | t_6__414_;
  assign t_7__349_ = t_6__349_ | t_6__413_;
  assign t_7__348_ = t_6__348_ | t_6__412_;
  assign t_7__347_ = t_6__347_ | t_6__411_;
  assign t_7__346_ = t_6__346_ | t_6__410_;
  assign t_7__345_ = t_6__345_ | t_6__409_;
  assign t_7__344_ = t_6__344_ | t_6__408_;
  assign t_7__343_ = t_6__343_ | t_6__407_;
  assign t_7__342_ = t_6__342_ | t_6__406_;
  assign t_7__341_ = t_6__341_ | t_6__405_;
  assign t_7__340_ = t_6__340_ | t_6__404_;
  assign t_7__339_ = t_6__339_ | t_6__403_;
  assign t_7__338_ = t_6__338_ | t_6__402_;
  assign t_7__337_ = t_6__337_ | t_6__401_;
  assign t_7__336_ = t_6__336_ | t_6__400_;
  assign t_7__335_ = t_6__335_ | t_6__399_;
  assign t_7__334_ = t_6__334_ | t_6__398_;
  assign t_7__333_ = t_6__333_ | t_6__397_;
  assign t_7__332_ = t_6__332_ | t_6__396_;
  assign t_7__331_ = t_6__331_ | t_6__395_;
  assign t_7__330_ = t_6__330_ | t_6__394_;
  assign t_7__329_ = t_6__329_ | t_6__393_;
  assign t_7__328_ = t_6__328_ | t_6__392_;
  assign t_7__327_ = t_6__327_ | t_6__391_;
  assign t_7__326_ = t_6__326_ | t_6__390_;
  assign t_7__325_ = t_6__325_ | t_6__389_;
  assign t_7__324_ = t_6__324_ | t_6__388_;
  assign t_7__323_ = t_6__323_ | t_6__387_;
  assign t_7__322_ = t_6__322_ | t_6__386_;
  assign t_7__321_ = t_6__321_ | t_6__385_;
  assign t_7__320_ = t_6__320_ | t_6__384_;
  assign t_7__319_ = t_6__319_ | t_6__383_;
  assign t_7__318_ = t_6__318_ | t_6__382_;
  assign t_7__317_ = t_6__317_ | t_6__381_;
  assign t_7__316_ = t_6__316_ | t_6__380_;
  assign t_7__315_ = t_6__315_ | t_6__379_;
  assign t_7__314_ = t_6__314_ | t_6__378_;
  assign t_7__313_ = t_6__313_ | t_6__377_;
  assign t_7__312_ = t_6__312_ | t_6__376_;
  assign t_7__311_ = t_6__311_ | t_6__375_;
  assign t_7__310_ = t_6__310_ | t_6__374_;
  assign t_7__309_ = t_6__309_ | t_6__373_;
  assign t_7__308_ = t_6__308_ | t_6__372_;
  assign t_7__307_ = t_6__307_ | t_6__371_;
  assign t_7__306_ = t_6__306_ | t_6__370_;
  assign t_7__305_ = t_6__305_ | t_6__369_;
  assign t_7__304_ = t_6__304_ | t_6__368_;
  assign t_7__303_ = t_6__303_ | t_6__367_;
  assign t_7__302_ = t_6__302_ | t_6__366_;
  assign t_7__301_ = t_6__301_ | t_6__365_;
  assign t_7__300_ = t_6__300_ | t_6__364_;
  assign t_7__299_ = t_6__299_ | t_6__363_;
  assign t_7__298_ = t_6__298_ | t_6__362_;
  assign t_7__297_ = t_6__297_ | t_6__361_;
  assign t_7__296_ = t_6__296_ | t_6__360_;
  assign t_7__295_ = t_6__295_ | t_6__359_;
  assign t_7__294_ = t_6__294_ | t_6__358_;
  assign t_7__293_ = t_6__293_ | t_6__357_;
  assign t_7__292_ = t_6__292_ | t_6__356_;
  assign t_7__291_ = t_6__291_ | t_6__355_;
  assign t_7__290_ = t_6__290_ | t_6__354_;
  assign t_7__289_ = t_6__289_ | t_6__353_;
  assign t_7__288_ = t_6__288_ | t_6__352_;
  assign t_7__287_ = t_6__287_ | t_6__351_;
  assign t_7__286_ = t_6__286_ | t_6__350_;
  assign t_7__285_ = t_6__285_ | t_6__349_;
  assign t_7__284_ = t_6__284_ | t_6__348_;
  assign t_7__283_ = t_6__283_ | t_6__347_;
  assign t_7__282_ = t_6__282_ | t_6__346_;
  assign t_7__281_ = t_6__281_ | t_6__345_;
  assign t_7__280_ = t_6__280_ | t_6__344_;
  assign t_7__279_ = t_6__279_ | t_6__343_;
  assign t_7__278_ = t_6__278_ | t_6__342_;
  assign t_7__277_ = t_6__277_ | t_6__341_;
  assign t_7__276_ = t_6__276_ | t_6__340_;
  assign t_7__275_ = t_6__275_ | t_6__339_;
  assign t_7__274_ = t_6__274_ | t_6__338_;
  assign t_7__273_ = t_6__273_ | t_6__337_;
  assign t_7__272_ = t_6__272_ | t_6__336_;
  assign t_7__271_ = t_6__271_ | t_6__335_;
  assign t_7__270_ = t_6__270_ | t_6__334_;
  assign t_7__269_ = t_6__269_ | t_6__333_;
  assign t_7__268_ = t_6__268_ | t_6__332_;
  assign t_7__267_ = t_6__267_ | t_6__331_;
  assign t_7__266_ = t_6__266_ | t_6__330_;
  assign t_7__265_ = t_6__265_ | t_6__329_;
  assign t_7__264_ = t_6__264_ | t_6__328_;
  assign t_7__263_ = t_6__263_ | t_6__327_;
  assign t_7__262_ = t_6__262_ | t_6__326_;
  assign t_7__261_ = t_6__261_ | t_6__325_;
  assign t_7__260_ = t_6__260_ | t_6__324_;
  assign t_7__259_ = t_6__259_ | t_6__323_;
  assign t_7__258_ = t_6__258_ | t_6__322_;
  assign t_7__257_ = t_6__257_ | t_6__321_;
  assign t_7__256_ = t_6__256_ | t_6__320_;
  assign t_7__255_ = t_6__255_ | t_6__319_;
  assign t_7__254_ = t_6__254_ | t_6__318_;
  assign t_7__253_ = t_6__253_ | t_6__317_;
  assign t_7__252_ = t_6__252_ | t_6__316_;
  assign t_7__251_ = t_6__251_ | t_6__315_;
  assign t_7__250_ = t_6__250_ | t_6__314_;
  assign t_7__249_ = t_6__249_ | t_6__313_;
  assign t_7__248_ = t_6__248_ | t_6__312_;
  assign t_7__247_ = t_6__247_ | t_6__311_;
  assign t_7__246_ = t_6__246_ | t_6__310_;
  assign t_7__245_ = t_6__245_ | t_6__309_;
  assign t_7__244_ = t_6__244_ | t_6__308_;
  assign t_7__243_ = t_6__243_ | t_6__307_;
  assign t_7__242_ = t_6__242_ | t_6__306_;
  assign t_7__241_ = t_6__241_ | t_6__305_;
  assign t_7__240_ = t_6__240_ | t_6__304_;
  assign t_7__239_ = t_6__239_ | t_6__303_;
  assign t_7__238_ = t_6__238_ | t_6__302_;
  assign t_7__237_ = t_6__237_ | t_6__301_;
  assign t_7__236_ = t_6__236_ | t_6__300_;
  assign t_7__235_ = t_6__235_ | t_6__299_;
  assign t_7__234_ = t_6__234_ | t_6__298_;
  assign t_7__233_ = t_6__233_ | t_6__297_;
  assign t_7__232_ = t_6__232_ | t_6__296_;
  assign t_7__231_ = t_6__231_ | t_6__295_;
  assign t_7__230_ = t_6__230_ | t_6__294_;
  assign t_7__229_ = t_6__229_ | t_6__293_;
  assign t_7__228_ = t_6__228_ | t_6__292_;
  assign t_7__227_ = t_6__227_ | t_6__291_;
  assign t_7__226_ = t_6__226_ | t_6__290_;
  assign t_7__225_ = t_6__225_ | t_6__289_;
  assign t_7__224_ = t_6__224_ | t_6__288_;
  assign t_7__223_ = t_6__223_ | t_6__287_;
  assign t_7__222_ = t_6__222_ | t_6__286_;
  assign t_7__221_ = t_6__221_ | t_6__285_;
  assign t_7__220_ = t_6__220_ | t_6__284_;
  assign t_7__219_ = t_6__219_ | t_6__283_;
  assign t_7__218_ = t_6__218_ | t_6__282_;
  assign t_7__217_ = t_6__217_ | t_6__281_;
  assign t_7__216_ = t_6__216_ | t_6__280_;
  assign t_7__215_ = t_6__215_ | t_6__279_;
  assign t_7__214_ = t_6__214_ | t_6__278_;
  assign t_7__213_ = t_6__213_ | t_6__277_;
  assign t_7__212_ = t_6__212_ | t_6__276_;
  assign t_7__211_ = t_6__211_ | t_6__275_;
  assign t_7__210_ = t_6__210_ | t_6__274_;
  assign t_7__209_ = t_6__209_ | t_6__273_;
  assign t_7__208_ = t_6__208_ | t_6__272_;
  assign t_7__207_ = t_6__207_ | t_6__271_;
  assign t_7__206_ = t_6__206_ | t_6__270_;
  assign t_7__205_ = t_6__205_ | t_6__269_;
  assign t_7__204_ = t_6__204_ | t_6__268_;
  assign t_7__203_ = t_6__203_ | t_6__267_;
  assign t_7__202_ = t_6__202_ | t_6__266_;
  assign t_7__201_ = t_6__201_ | t_6__265_;
  assign t_7__200_ = t_6__200_ | t_6__264_;
  assign t_7__199_ = t_6__199_ | t_6__263_;
  assign t_7__198_ = t_6__198_ | t_6__262_;
  assign t_7__197_ = t_6__197_ | t_6__261_;
  assign t_7__196_ = t_6__196_ | t_6__260_;
  assign t_7__195_ = t_6__195_ | t_6__259_;
  assign t_7__194_ = t_6__194_ | t_6__258_;
  assign t_7__193_ = t_6__193_ | t_6__257_;
  assign t_7__192_ = t_6__192_ | t_6__256_;
  assign t_7__191_ = t_6__191_ | t_6__255_;
  assign t_7__190_ = t_6__190_ | t_6__254_;
  assign t_7__189_ = t_6__189_ | t_6__253_;
  assign t_7__188_ = t_6__188_ | t_6__252_;
  assign t_7__187_ = t_6__187_ | t_6__251_;
  assign t_7__186_ = t_6__186_ | t_6__250_;
  assign t_7__185_ = t_6__185_ | t_6__249_;
  assign t_7__184_ = t_6__184_ | t_6__248_;
  assign t_7__183_ = t_6__183_ | t_6__247_;
  assign t_7__182_ = t_6__182_ | t_6__246_;
  assign t_7__181_ = t_6__181_ | t_6__245_;
  assign t_7__180_ = t_6__180_ | t_6__244_;
  assign t_7__179_ = t_6__179_ | t_6__243_;
  assign t_7__178_ = t_6__178_ | t_6__242_;
  assign t_7__177_ = t_6__177_ | t_6__241_;
  assign t_7__176_ = t_6__176_ | t_6__240_;
  assign t_7__175_ = t_6__175_ | t_6__239_;
  assign t_7__174_ = t_6__174_ | t_6__238_;
  assign t_7__173_ = t_6__173_ | t_6__237_;
  assign t_7__172_ = t_6__172_ | t_6__236_;
  assign t_7__171_ = t_6__171_ | t_6__235_;
  assign t_7__170_ = t_6__170_ | t_6__234_;
  assign t_7__169_ = t_6__169_ | t_6__233_;
  assign t_7__168_ = t_6__168_ | t_6__232_;
  assign t_7__167_ = t_6__167_ | t_6__231_;
  assign t_7__166_ = t_6__166_ | t_6__230_;
  assign t_7__165_ = t_6__165_ | t_6__229_;
  assign t_7__164_ = t_6__164_ | t_6__228_;
  assign t_7__163_ = t_6__163_ | t_6__227_;
  assign t_7__162_ = t_6__162_ | t_6__226_;
  assign t_7__161_ = t_6__161_ | t_6__225_;
  assign t_7__160_ = t_6__160_ | t_6__224_;
  assign t_7__159_ = t_6__159_ | t_6__223_;
  assign t_7__158_ = t_6__158_ | t_6__222_;
  assign t_7__157_ = t_6__157_ | t_6__221_;
  assign t_7__156_ = t_6__156_ | t_6__220_;
  assign t_7__155_ = t_6__155_ | t_6__219_;
  assign t_7__154_ = t_6__154_ | t_6__218_;
  assign t_7__153_ = t_6__153_ | t_6__217_;
  assign t_7__152_ = t_6__152_ | t_6__216_;
  assign t_7__151_ = t_6__151_ | t_6__215_;
  assign t_7__150_ = t_6__150_ | t_6__214_;
  assign t_7__149_ = t_6__149_ | t_6__213_;
  assign t_7__148_ = t_6__148_ | t_6__212_;
  assign t_7__147_ = t_6__147_ | t_6__211_;
  assign t_7__146_ = t_6__146_ | t_6__210_;
  assign t_7__145_ = t_6__145_ | t_6__209_;
  assign t_7__144_ = t_6__144_ | t_6__208_;
  assign t_7__143_ = t_6__143_ | t_6__207_;
  assign t_7__142_ = t_6__142_ | t_6__206_;
  assign t_7__141_ = t_6__141_ | t_6__205_;
  assign t_7__140_ = t_6__140_ | t_6__204_;
  assign t_7__139_ = t_6__139_ | t_6__203_;
  assign t_7__138_ = t_6__138_ | t_6__202_;
  assign t_7__137_ = t_6__137_ | t_6__201_;
  assign t_7__136_ = t_6__136_ | t_6__200_;
  assign t_7__135_ = t_6__135_ | t_6__199_;
  assign t_7__134_ = t_6__134_ | t_6__198_;
  assign t_7__133_ = t_6__133_ | t_6__197_;
  assign t_7__132_ = t_6__132_ | t_6__196_;
  assign t_7__131_ = t_6__131_ | t_6__195_;
  assign t_7__130_ = t_6__130_ | t_6__194_;
  assign t_7__129_ = t_6__129_ | t_6__193_;
  assign t_7__128_ = t_6__128_ | t_6__192_;
  assign t_7__127_ = t_6__127_ | t_6__191_;
  assign t_7__126_ = t_6__126_ | t_6__190_;
  assign t_7__125_ = t_6__125_ | t_6__189_;
  assign t_7__124_ = t_6__124_ | t_6__188_;
  assign t_7__123_ = t_6__123_ | t_6__187_;
  assign t_7__122_ = t_6__122_ | t_6__186_;
  assign t_7__121_ = t_6__121_ | t_6__185_;
  assign t_7__120_ = t_6__120_ | t_6__184_;
  assign t_7__119_ = t_6__119_ | t_6__183_;
  assign t_7__118_ = t_6__118_ | t_6__182_;
  assign t_7__117_ = t_6__117_ | t_6__181_;
  assign t_7__116_ = t_6__116_ | t_6__180_;
  assign t_7__115_ = t_6__115_ | t_6__179_;
  assign t_7__114_ = t_6__114_ | t_6__178_;
  assign t_7__113_ = t_6__113_ | t_6__177_;
  assign t_7__112_ = t_6__112_ | t_6__176_;
  assign t_7__111_ = t_6__111_ | t_6__175_;
  assign t_7__110_ = t_6__110_ | t_6__174_;
  assign t_7__109_ = t_6__109_ | t_6__173_;
  assign t_7__108_ = t_6__108_ | t_6__172_;
  assign t_7__107_ = t_6__107_ | t_6__171_;
  assign t_7__106_ = t_6__106_ | t_6__170_;
  assign t_7__105_ = t_6__105_ | t_6__169_;
  assign t_7__104_ = t_6__104_ | t_6__168_;
  assign t_7__103_ = t_6__103_ | t_6__167_;
  assign t_7__102_ = t_6__102_ | t_6__166_;
  assign t_7__101_ = t_6__101_ | t_6__165_;
  assign t_7__100_ = t_6__100_ | t_6__164_;
  assign t_7__99_ = t_6__99_ | t_6__163_;
  assign t_7__98_ = t_6__98_ | t_6__162_;
  assign t_7__97_ = t_6__97_ | t_6__161_;
  assign t_7__96_ = t_6__96_ | t_6__160_;
  assign t_7__95_ = t_6__95_ | t_6__159_;
  assign t_7__94_ = t_6__94_ | t_6__158_;
  assign t_7__93_ = t_6__93_ | t_6__157_;
  assign t_7__92_ = t_6__92_ | t_6__156_;
  assign t_7__91_ = t_6__91_ | t_6__155_;
  assign t_7__90_ = t_6__90_ | t_6__154_;
  assign t_7__89_ = t_6__89_ | t_6__153_;
  assign t_7__88_ = t_6__88_ | t_6__152_;
  assign t_7__87_ = t_6__87_ | t_6__151_;
  assign t_7__86_ = t_6__86_ | t_6__150_;
  assign t_7__85_ = t_6__85_ | t_6__149_;
  assign t_7__84_ = t_6__84_ | t_6__148_;
  assign t_7__83_ = t_6__83_ | t_6__147_;
  assign t_7__82_ = t_6__82_ | t_6__146_;
  assign t_7__81_ = t_6__81_ | t_6__145_;
  assign t_7__80_ = t_6__80_ | t_6__144_;
  assign t_7__79_ = t_6__79_ | t_6__143_;
  assign t_7__78_ = t_6__78_ | t_6__142_;
  assign t_7__77_ = t_6__77_ | t_6__141_;
  assign t_7__76_ = t_6__76_ | t_6__140_;
  assign t_7__75_ = t_6__75_ | t_6__139_;
  assign t_7__74_ = t_6__74_ | t_6__138_;
  assign t_7__73_ = t_6__73_ | t_6__137_;
  assign t_7__72_ = t_6__72_ | t_6__136_;
  assign t_7__71_ = t_6__71_ | t_6__135_;
  assign t_7__70_ = t_6__70_ | t_6__134_;
  assign t_7__69_ = t_6__69_ | t_6__133_;
  assign t_7__68_ = t_6__68_ | t_6__132_;
  assign t_7__67_ = t_6__67_ | t_6__131_;
  assign t_7__66_ = t_6__66_ | t_6__130_;
  assign t_7__65_ = t_6__65_ | t_6__129_;
  assign t_7__64_ = t_6__64_ | t_6__128_;
  assign t_7__63_ = t_6__63_ | t_6__127_;
  assign t_7__62_ = t_6__62_ | t_6__126_;
  assign t_7__61_ = t_6__61_ | t_6__125_;
  assign t_7__60_ = t_6__60_ | t_6__124_;
  assign t_7__59_ = t_6__59_ | t_6__123_;
  assign t_7__58_ = t_6__58_ | t_6__122_;
  assign t_7__57_ = t_6__57_ | t_6__121_;
  assign t_7__56_ = t_6__56_ | t_6__120_;
  assign t_7__55_ = t_6__55_ | t_6__119_;
  assign t_7__54_ = t_6__54_ | t_6__118_;
  assign t_7__53_ = t_6__53_ | t_6__117_;
  assign t_7__52_ = t_6__52_ | t_6__116_;
  assign t_7__51_ = t_6__51_ | t_6__115_;
  assign t_7__50_ = t_6__50_ | t_6__114_;
  assign t_7__49_ = t_6__49_ | t_6__113_;
  assign t_7__48_ = t_6__48_ | t_6__112_;
  assign t_7__47_ = t_6__47_ | t_6__111_;
  assign t_7__46_ = t_6__46_ | t_6__110_;
  assign t_7__45_ = t_6__45_ | t_6__109_;
  assign t_7__44_ = t_6__44_ | t_6__108_;
  assign t_7__43_ = t_6__43_ | t_6__107_;
  assign t_7__42_ = t_6__42_ | t_6__106_;
  assign t_7__41_ = t_6__41_ | t_6__105_;
  assign t_7__40_ = t_6__40_ | t_6__104_;
  assign t_7__39_ = t_6__39_ | t_6__103_;
  assign t_7__38_ = t_6__38_ | t_6__102_;
  assign t_7__37_ = t_6__37_ | t_6__101_;
  assign t_7__36_ = t_6__36_ | t_6__100_;
  assign t_7__35_ = t_6__35_ | t_6__99_;
  assign t_7__34_ = t_6__34_ | t_6__98_;
  assign t_7__33_ = t_6__33_ | t_6__97_;
  assign t_7__32_ = t_6__32_ | t_6__96_;
  assign t_7__31_ = t_6__31_ | t_6__95_;
  assign t_7__30_ = t_6__30_ | t_6__94_;
  assign t_7__29_ = t_6__29_ | t_6__93_;
  assign t_7__28_ = t_6__28_ | t_6__92_;
  assign t_7__27_ = t_6__27_ | t_6__91_;
  assign t_7__26_ = t_6__26_ | t_6__90_;
  assign t_7__25_ = t_6__25_ | t_6__89_;
  assign t_7__24_ = t_6__24_ | t_6__88_;
  assign t_7__23_ = t_6__23_ | t_6__87_;
  assign t_7__22_ = t_6__22_ | t_6__86_;
  assign t_7__21_ = t_6__21_ | t_6__85_;
  assign t_7__20_ = t_6__20_ | t_6__84_;
  assign t_7__19_ = t_6__19_ | t_6__83_;
  assign t_7__18_ = t_6__18_ | t_6__82_;
  assign t_7__17_ = t_6__17_ | t_6__81_;
  assign t_7__16_ = t_6__16_ | t_6__80_;
  assign t_7__15_ = t_6__15_ | t_6__79_;
  assign t_7__14_ = t_6__14_ | t_6__78_;
  assign t_7__13_ = t_6__13_ | t_6__77_;
  assign t_7__12_ = t_6__12_ | t_6__76_;
  assign t_7__11_ = t_6__11_ | t_6__75_;
  assign t_7__10_ = t_6__10_ | t_6__74_;
  assign t_7__9_ = t_6__9_ | t_6__73_;
  assign t_7__8_ = t_6__8_ | t_6__72_;
  assign t_7__7_ = t_6__7_ | t_6__71_;
  assign t_7__6_ = t_6__6_ | t_6__70_;
  assign t_7__5_ = t_6__5_ | t_6__69_;
  assign t_7__4_ = t_6__4_ | t_6__68_;
  assign t_7__3_ = t_6__3_ | t_6__67_;
  assign t_7__2_ = t_6__2_ | t_6__66_;
  assign t_7__1_ = t_6__1_ | t_6__65_;
  assign t_7__0_ = t_6__0_ | t_6__64_;
  assign t_8__1023_ = t_7__1023_ | 1'b0;
  assign t_8__1022_ = t_7__1022_ | 1'b0;
  assign t_8__1021_ = t_7__1021_ | 1'b0;
  assign t_8__1020_ = t_7__1020_ | 1'b0;
  assign t_8__1019_ = t_7__1019_ | 1'b0;
  assign t_8__1018_ = t_7__1018_ | 1'b0;
  assign t_8__1017_ = t_7__1017_ | 1'b0;
  assign t_8__1016_ = t_7__1016_ | 1'b0;
  assign t_8__1015_ = t_7__1015_ | 1'b0;
  assign t_8__1014_ = t_7__1014_ | 1'b0;
  assign t_8__1013_ = t_7__1013_ | 1'b0;
  assign t_8__1012_ = t_7__1012_ | 1'b0;
  assign t_8__1011_ = t_7__1011_ | 1'b0;
  assign t_8__1010_ = t_7__1010_ | 1'b0;
  assign t_8__1009_ = t_7__1009_ | 1'b0;
  assign t_8__1008_ = t_7__1008_ | 1'b0;
  assign t_8__1007_ = t_7__1007_ | 1'b0;
  assign t_8__1006_ = t_7__1006_ | 1'b0;
  assign t_8__1005_ = t_7__1005_ | 1'b0;
  assign t_8__1004_ = t_7__1004_ | 1'b0;
  assign t_8__1003_ = t_7__1003_ | 1'b0;
  assign t_8__1002_ = t_7__1002_ | 1'b0;
  assign t_8__1001_ = t_7__1001_ | 1'b0;
  assign t_8__1000_ = t_7__1000_ | 1'b0;
  assign t_8__999_ = t_7__999_ | 1'b0;
  assign t_8__998_ = t_7__998_ | 1'b0;
  assign t_8__997_ = t_7__997_ | 1'b0;
  assign t_8__996_ = t_7__996_ | 1'b0;
  assign t_8__995_ = t_7__995_ | 1'b0;
  assign t_8__994_ = t_7__994_ | 1'b0;
  assign t_8__993_ = t_7__993_ | 1'b0;
  assign t_8__992_ = t_7__992_ | 1'b0;
  assign t_8__991_ = t_7__991_ | 1'b0;
  assign t_8__990_ = t_7__990_ | 1'b0;
  assign t_8__989_ = t_7__989_ | 1'b0;
  assign t_8__988_ = t_7__988_ | 1'b0;
  assign t_8__987_ = t_7__987_ | 1'b0;
  assign t_8__986_ = t_7__986_ | 1'b0;
  assign t_8__985_ = t_7__985_ | 1'b0;
  assign t_8__984_ = t_7__984_ | 1'b0;
  assign t_8__983_ = t_7__983_ | 1'b0;
  assign t_8__982_ = t_7__982_ | 1'b0;
  assign t_8__981_ = t_7__981_ | 1'b0;
  assign t_8__980_ = t_7__980_ | 1'b0;
  assign t_8__979_ = t_7__979_ | 1'b0;
  assign t_8__978_ = t_7__978_ | 1'b0;
  assign t_8__977_ = t_7__977_ | 1'b0;
  assign t_8__976_ = t_7__976_ | 1'b0;
  assign t_8__975_ = t_7__975_ | 1'b0;
  assign t_8__974_ = t_7__974_ | 1'b0;
  assign t_8__973_ = t_7__973_ | 1'b0;
  assign t_8__972_ = t_7__972_ | 1'b0;
  assign t_8__971_ = t_7__971_ | 1'b0;
  assign t_8__970_ = t_7__970_ | 1'b0;
  assign t_8__969_ = t_7__969_ | 1'b0;
  assign t_8__968_ = t_7__968_ | 1'b0;
  assign t_8__967_ = t_7__967_ | 1'b0;
  assign t_8__966_ = t_7__966_ | 1'b0;
  assign t_8__965_ = t_7__965_ | 1'b0;
  assign t_8__964_ = t_7__964_ | 1'b0;
  assign t_8__963_ = t_7__963_ | 1'b0;
  assign t_8__962_ = t_7__962_ | 1'b0;
  assign t_8__961_ = t_7__961_ | 1'b0;
  assign t_8__960_ = t_7__960_ | 1'b0;
  assign t_8__959_ = t_7__959_ | 1'b0;
  assign t_8__958_ = t_7__958_ | 1'b0;
  assign t_8__957_ = t_7__957_ | 1'b0;
  assign t_8__956_ = t_7__956_ | 1'b0;
  assign t_8__955_ = t_7__955_ | 1'b0;
  assign t_8__954_ = t_7__954_ | 1'b0;
  assign t_8__953_ = t_7__953_ | 1'b0;
  assign t_8__952_ = t_7__952_ | 1'b0;
  assign t_8__951_ = t_7__951_ | 1'b0;
  assign t_8__950_ = t_7__950_ | 1'b0;
  assign t_8__949_ = t_7__949_ | 1'b0;
  assign t_8__948_ = t_7__948_ | 1'b0;
  assign t_8__947_ = t_7__947_ | 1'b0;
  assign t_8__946_ = t_7__946_ | 1'b0;
  assign t_8__945_ = t_7__945_ | 1'b0;
  assign t_8__944_ = t_7__944_ | 1'b0;
  assign t_8__943_ = t_7__943_ | 1'b0;
  assign t_8__942_ = t_7__942_ | 1'b0;
  assign t_8__941_ = t_7__941_ | 1'b0;
  assign t_8__940_ = t_7__940_ | 1'b0;
  assign t_8__939_ = t_7__939_ | 1'b0;
  assign t_8__938_ = t_7__938_ | 1'b0;
  assign t_8__937_ = t_7__937_ | 1'b0;
  assign t_8__936_ = t_7__936_ | 1'b0;
  assign t_8__935_ = t_7__935_ | 1'b0;
  assign t_8__934_ = t_7__934_ | 1'b0;
  assign t_8__933_ = t_7__933_ | 1'b0;
  assign t_8__932_ = t_7__932_ | 1'b0;
  assign t_8__931_ = t_7__931_ | 1'b0;
  assign t_8__930_ = t_7__930_ | 1'b0;
  assign t_8__929_ = t_7__929_ | 1'b0;
  assign t_8__928_ = t_7__928_ | 1'b0;
  assign t_8__927_ = t_7__927_ | 1'b0;
  assign t_8__926_ = t_7__926_ | 1'b0;
  assign t_8__925_ = t_7__925_ | 1'b0;
  assign t_8__924_ = t_7__924_ | 1'b0;
  assign t_8__923_ = t_7__923_ | 1'b0;
  assign t_8__922_ = t_7__922_ | 1'b0;
  assign t_8__921_ = t_7__921_ | 1'b0;
  assign t_8__920_ = t_7__920_ | 1'b0;
  assign t_8__919_ = t_7__919_ | 1'b0;
  assign t_8__918_ = t_7__918_ | 1'b0;
  assign t_8__917_ = t_7__917_ | 1'b0;
  assign t_8__916_ = t_7__916_ | 1'b0;
  assign t_8__915_ = t_7__915_ | 1'b0;
  assign t_8__914_ = t_7__914_ | 1'b0;
  assign t_8__913_ = t_7__913_ | 1'b0;
  assign t_8__912_ = t_7__912_ | 1'b0;
  assign t_8__911_ = t_7__911_ | 1'b0;
  assign t_8__910_ = t_7__910_ | 1'b0;
  assign t_8__909_ = t_7__909_ | 1'b0;
  assign t_8__908_ = t_7__908_ | 1'b0;
  assign t_8__907_ = t_7__907_ | 1'b0;
  assign t_8__906_ = t_7__906_ | 1'b0;
  assign t_8__905_ = t_7__905_ | 1'b0;
  assign t_8__904_ = t_7__904_ | 1'b0;
  assign t_8__903_ = t_7__903_ | 1'b0;
  assign t_8__902_ = t_7__902_ | 1'b0;
  assign t_8__901_ = t_7__901_ | 1'b0;
  assign t_8__900_ = t_7__900_ | 1'b0;
  assign t_8__899_ = t_7__899_ | 1'b0;
  assign t_8__898_ = t_7__898_ | 1'b0;
  assign t_8__897_ = t_7__897_ | 1'b0;
  assign t_8__896_ = t_7__896_ | 1'b0;
  assign t_8__895_ = t_7__895_ | t_7__1023_;
  assign t_8__894_ = t_7__894_ | t_7__1022_;
  assign t_8__893_ = t_7__893_ | t_7__1021_;
  assign t_8__892_ = t_7__892_ | t_7__1020_;
  assign t_8__891_ = t_7__891_ | t_7__1019_;
  assign t_8__890_ = t_7__890_ | t_7__1018_;
  assign t_8__889_ = t_7__889_ | t_7__1017_;
  assign t_8__888_ = t_7__888_ | t_7__1016_;
  assign t_8__887_ = t_7__887_ | t_7__1015_;
  assign t_8__886_ = t_7__886_ | t_7__1014_;
  assign t_8__885_ = t_7__885_ | t_7__1013_;
  assign t_8__884_ = t_7__884_ | t_7__1012_;
  assign t_8__883_ = t_7__883_ | t_7__1011_;
  assign t_8__882_ = t_7__882_ | t_7__1010_;
  assign t_8__881_ = t_7__881_ | t_7__1009_;
  assign t_8__880_ = t_7__880_ | t_7__1008_;
  assign t_8__879_ = t_7__879_ | t_7__1007_;
  assign t_8__878_ = t_7__878_ | t_7__1006_;
  assign t_8__877_ = t_7__877_ | t_7__1005_;
  assign t_8__876_ = t_7__876_ | t_7__1004_;
  assign t_8__875_ = t_7__875_ | t_7__1003_;
  assign t_8__874_ = t_7__874_ | t_7__1002_;
  assign t_8__873_ = t_7__873_ | t_7__1001_;
  assign t_8__872_ = t_7__872_ | t_7__1000_;
  assign t_8__871_ = t_7__871_ | t_7__999_;
  assign t_8__870_ = t_7__870_ | t_7__998_;
  assign t_8__869_ = t_7__869_ | t_7__997_;
  assign t_8__868_ = t_7__868_ | t_7__996_;
  assign t_8__867_ = t_7__867_ | t_7__995_;
  assign t_8__866_ = t_7__866_ | t_7__994_;
  assign t_8__865_ = t_7__865_ | t_7__993_;
  assign t_8__864_ = t_7__864_ | t_7__992_;
  assign t_8__863_ = t_7__863_ | t_7__991_;
  assign t_8__862_ = t_7__862_ | t_7__990_;
  assign t_8__861_ = t_7__861_ | t_7__989_;
  assign t_8__860_ = t_7__860_ | t_7__988_;
  assign t_8__859_ = t_7__859_ | t_7__987_;
  assign t_8__858_ = t_7__858_ | t_7__986_;
  assign t_8__857_ = t_7__857_ | t_7__985_;
  assign t_8__856_ = t_7__856_ | t_7__984_;
  assign t_8__855_ = t_7__855_ | t_7__983_;
  assign t_8__854_ = t_7__854_ | t_7__982_;
  assign t_8__853_ = t_7__853_ | t_7__981_;
  assign t_8__852_ = t_7__852_ | t_7__980_;
  assign t_8__851_ = t_7__851_ | t_7__979_;
  assign t_8__850_ = t_7__850_ | t_7__978_;
  assign t_8__849_ = t_7__849_ | t_7__977_;
  assign t_8__848_ = t_7__848_ | t_7__976_;
  assign t_8__847_ = t_7__847_ | t_7__975_;
  assign t_8__846_ = t_7__846_ | t_7__974_;
  assign t_8__845_ = t_7__845_ | t_7__973_;
  assign t_8__844_ = t_7__844_ | t_7__972_;
  assign t_8__843_ = t_7__843_ | t_7__971_;
  assign t_8__842_ = t_7__842_ | t_7__970_;
  assign t_8__841_ = t_7__841_ | t_7__969_;
  assign t_8__840_ = t_7__840_ | t_7__968_;
  assign t_8__839_ = t_7__839_ | t_7__967_;
  assign t_8__838_ = t_7__838_ | t_7__966_;
  assign t_8__837_ = t_7__837_ | t_7__965_;
  assign t_8__836_ = t_7__836_ | t_7__964_;
  assign t_8__835_ = t_7__835_ | t_7__963_;
  assign t_8__834_ = t_7__834_ | t_7__962_;
  assign t_8__833_ = t_7__833_ | t_7__961_;
  assign t_8__832_ = t_7__832_ | t_7__960_;
  assign t_8__831_ = t_7__831_ | t_7__959_;
  assign t_8__830_ = t_7__830_ | t_7__958_;
  assign t_8__829_ = t_7__829_ | t_7__957_;
  assign t_8__828_ = t_7__828_ | t_7__956_;
  assign t_8__827_ = t_7__827_ | t_7__955_;
  assign t_8__826_ = t_7__826_ | t_7__954_;
  assign t_8__825_ = t_7__825_ | t_7__953_;
  assign t_8__824_ = t_7__824_ | t_7__952_;
  assign t_8__823_ = t_7__823_ | t_7__951_;
  assign t_8__822_ = t_7__822_ | t_7__950_;
  assign t_8__821_ = t_7__821_ | t_7__949_;
  assign t_8__820_ = t_7__820_ | t_7__948_;
  assign t_8__819_ = t_7__819_ | t_7__947_;
  assign t_8__818_ = t_7__818_ | t_7__946_;
  assign t_8__817_ = t_7__817_ | t_7__945_;
  assign t_8__816_ = t_7__816_ | t_7__944_;
  assign t_8__815_ = t_7__815_ | t_7__943_;
  assign t_8__814_ = t_7__814_ | t_7__942_;
  assign t_8__813_ = t_7__813_ | t_7__941_;
  assign t_8__812_ = t_7__812_ | t_7__940_;
  assign t_8__811_ = t_7__811_ | t_7__939_;
  assign t_8__810_ = t_7__810_ | t_7__938_;
  assign t_8__809_ = t_7__809_ | t_7__937_;
  assign t_8__808_ = t_7__808_ | t_7__936_;
  assign t_8__807_ = t_7__807_ | t_7__935_;
  assign t_8__806_ = t_7__806_ | t_7__934_;
  assign t_8__805_ = t_7__805_ | t_7__933_;
  assign t_8__804_ = t_7__804_ | t_7__932_;
  assign t_8__803_ = t_7__803_ | t_7__931_;
  assign t_8__802_ = t_7__802_ | t_7__930_;
  assign t_8__801_ = t_7__801_ | t_7__929_;
  assign t_8__800_ = t_7__800_ | t_7__928_;
  assign t_8__799_ = t_7__799_ | t_7__927_;
  assign t_8__798_ = t_7__798_ | t_7__926_;
  assign t_8__797_ = t_7__797_ | t_7__925_;
  assign t_8__796_ = t_7__796_ | t_7__924_;
  assign t_8__795_ = t_7__795_ | t_7__923_;
  assign t_8__794_ = t_7__794_ | t_7__922_;
  assign t_8__793_ = t_7__793_ | t_7__921_;
  assign t_8__792_ = t_7__792_ | t_7__920_;
  assign t_8__791_ = t_7__791_ | t_7__919_;
  assign t_8__790_ = t_7__790_ | t_7__918_;
  assign t_8__789_ = t_7__789_ | t_7__917_;
  assign t_8__788_ = t_7__788_ | t_7__916_;
  assign t_8__787_ = t_7__787_ | t_7__915_;
  assign t_8__786_ = t_7__786_ | t_7__914_;
  assign t_8__785_ = t_7__785_ | t_7__913_;
  assign t_8__784_ = t_7__784_ | t_7__912_;
  assign t_8__783_ = t_7__783_ | t_7__911_;
  assign t_8__782_ = t_7__782_ | t_7__910_;
  assign t_8__781_ = t_7__781_ | t_7__909_;
  assign t_8__780_ = t_7__780_ | t_7__908_;
  assign t_8__779_ = t_7__779_ | t_7__907_;
  assign t_8__778_ = t_7__778_ | t_7__906_;
  assign t_8__777_ = t_7__777_ | t_7__905_;
  assign t_8__776_ = t_7__776_ | t_7__904_;
  assign t_8__775_ = t_7__775_ | t_7__903_;
  assign t_8__774_ = t_7__774_ | t_7__902_;
  assign t_8__773_ = t_7__773_ | t_7__901_;
  assign t_8__772_ = t_7__772_ | t_7__900_;
  assign t_8__771_ = t_7__771_ | t_7__899_;
  assign t_8__770_ = t_7__770_ | t_7__898_;
  assign t_8__769_ = t_7__769_ | t_7__897_;
  assign t_8__768_ = t_7__768_ | t_7__896_;
  assign t_8__767_ = t_7__767_ | t_7__895_;
  assign t_8__766_ = t_7__766_ | t_7__894_;
  assign t_8__765_ = t_7__765_ | t_7__893_;
  assign t_8__764_ = t_7__764_ | t_7__892_;
  assign t_8__763_ = t_7__763_ | t_7__891_;
  assign t_8__762_ = t_7__762_ | t_7__890_;
  assign t_8__761_ = t_7__761_ | t_7__889_;
  assign t_8__760_ = t_7__760_ | t_7__888_;
  assign t_8__759_ = t_7__759_ | t_7__887_;
  assign t_8__758_ = t_7__758_ | t_7__886_;
  assign t_8__757_ = t_7__757_ | t_7__885_;
  assign t_8__756_ = t_7__756_ | t_7__884_;
  assign t_8__755_ = t_7__755_ | t_7__883_;
  assign t_8__754_ = t_7__754_ | t_7__882_;
  assign t_8__753_ = t_7__753_ | t_7__881_;
  assign t_8__752_ = t_7__752_ | t_7__880_;
  assign t_8__751_ = t_7__751_ | t_7__879_;
  assign t_8__750_ = t_7__750_ | t_7__878_;
  assign t_8__749_ = t_7__749_ | t_7__877_;
  assign t_8__748_ = t_7__748_ | t_7__876_;
  assign t_8__747_ = t_7__747_ | t_7__875_;
  assign t_8__746_ = t_7__746_ | t_7__874_;
  assign t_8__745_ = t_7__745_ | t_7__873_;
  assign t_8__744_ = t_7__744_ | t_7__872_;
  assign t_8__743_ = t_7__743_ | t_7__871_;
  assign t_8__742_ = t_7__742_ | t_7__870_;
  assign t_8__741_ = t_7__741_ | t_7__869_;
  assign t_8__740_ = t_7__740_ | t_7__868_;
  assign t_8__739_ = t_7__739_ | t_7__867_;
  assign t_8__738_ = t_7__738_ | t_7__866_;
  assign t_8__737_ = t_7__737_ | t_7__865_;
  assign t_8__736_ = t_7__736_ | t_7__864_;
  assign t_8__735_ = t_7__735_ | t_7__863_;
  assign t_8__734_ = t_7__734_ | t_7__862_;
  assign t_8__733_ = t_7__733_ | t_7__861_;
  assign t_8__732_ = t_7__732_ | t_7__860_;
  assign t_8__731_ = t_7__731_ | t_7__859_;
  assign t_8__730_ = t_7__730_ | t_7__858_;
  assign t_8__729_ = t_7__729_ | t_7__857_;
  assign t_8__728_ = t_7__728_ | t_7__856_;
  assign t_8__727_ = t_7__727_ | t_7__855_;
  assign t_8__726_ = t_7__726_ | t_7__854_;
  assign t_8__725_ = t_7__725_ | t_7__853_;
  assign t_8__724_ = t_7__724_ | t_7__852_;
  assign t_8__723_ = t_7__723_ | t_7__851_;
  assign t_8__722_ = t_7__722_ | t_7__850_;
  assign t_8__721_ = t_7__721_ | t_7__849_;
  assign t_8__720_ = t_7__720_ | t_7__848_;
  assign t_8__719_ = t_7__719_ | t_7__847_;
  assign t_8__718_ = t_7__718_ | t_7__846_;
  assign t_8__717_ = t_7__717_ | t_7__845_;
  assign t_8__716_ = t_7__716_ | t_7__844_;
  assign t_8__715_ = t_7__715_ | t_7__843_;
  assign t_8__714_ = t_7__714_ | t_7__842_;
  assign t_8__713_ = t_7__713_ | t_7__841_;
  assign t_8__712_ = t_7__712_ | t_7__840_;
  assign t_8__711_ = t_7__711_ | t_7__839_;
  assign t_8__710_ = t_7__710_ | t_7__838_;
  assign t_8__709_ = t_7__709_ | t_7__837_;
  assign t_8__708_ = t_7__708_ | t_7__836_;
  assign t_8__707_ = t_7__707_ | t_7__835_;
  assign t_8__706_ = t_7__706_ | t_7__834_;
  assign t_8__705_ = t_7__705_ | t_7__833_;
  assign t_8__704_ = t_7__704_ | t_7__832_;
  assign t_8__703_ = t_7__703_ | t_7__831_;
  assign t_8__702_ = t_7__702_ | t_7__830_;
  assign t_8__701_ = t_7__701_ | t_7__829_;
  assign t_8__700_ = t_7__700_ | t_7__828_;
  assign t_8__699_ = t_7__699_ | t_7__827_;
  assign t_8__698_ = t_7__698_ | t_7__826_;
  assign t_8__697_ = t_7__697_ | t_7__825_;
  assign t_8__696_ = t_7__696_ | t_7__824_;
  assign t_8__695_ = t_7__695_ | t_7__823_;
  assign t_8__694_ = t_7__694_ | t_7__822_;
  assign t_8__693_ = t_7__693_ | t_7__821_;
  assign t_8__692_ = t_7__692_ | t_7__820_;
  assign t_8__691_ = t_7__691_ | t_7__819_;
  assign t_8__690_ = t_7__690_ | t_7__818_;
  assign t_8__689_ = t_7__689_ | t_7__817_;
  assign t_8__688_ = t_7__688_ | t_7__816_;
  assign t_8__687_ = t_7__687_ | t_7__815_;
  assign t_8__686_ = t_7__686_ | t_7__814_;
  assign t_8__685_ = t_7__685_ | t_7__813_;
  assign t_8__684_ = t_7__684_ | t_7__812_;
  assign t_8__683_ = t_7__683_ | t_7__811_;
  assign t_8__682_ = t_7__682_ | t_7__810_;
  assign t_8__681_ = t_7__681_ | t_7__809_;
  assign t_8__680_ = t_7__680_ | t_7__808_;
  assign t_8__679_ = t_7__679_ | t_7__807_;
  assign t_8__678_ = t_7__678_ | t_7__806_;
  assign t_8__677_ = t_7__677_ | t_7__805_;
  assign t_8__676_ = t_7__676_ | t_7__804_;
  assign t_8__675_ = t_7__675_ | t_7__803_;
  assign t_8__674_ = t_7__674_ | t_7__802_;
  assign t_8__673_ = t_7__673_ | t_7__801_;
  assign t_8__672_ = t_7__672_ | t_7__800_;
  assign t_8__671_ = t_7__671_ | t_7__799_;
  assign t_8__670_ = t_7__670_ | t_7__798_;
  assign t_8__669_ = t_7__669_ | t_7__797_;
  assign t_8__668_ = t_7__668_ | t_7__796_;
  assign t_8__667_ = t_7__667_ | t_7__795_;
  assign t_8__666_ = t_7__666_ | t_7__794_;
  assign t_8__665_ = t_7__665_ | t_7__793_;
  assign t_8__664_ = t_7__664_ | t_7__792_;
  assign t_8__663_ = t_7__663_ | t_7__791_;
  assign t_8__662_ = t_7__662_ | t_7__790_;
  assign t_8__661_ = t_7__661_ | t_7__789_;
  assign t_8__660_ = t_7__660_ | t_7__788_;
  assign t_8__659_ = t_7__659_ | t_7__787_;
  assign t_8__658_ = t_7__658_ | t_7__786_;
  assign t_8__657_ = t_7__657_ | t_7__785_;
  assign t_8__656_ = t_7__656_ | t_7__784_;
  assign t_8__655_ = t_7__655_ | t_7__783_;
  assign t_8__654_ = t_7__654_ | t_7__782_;
  assign t_8__653_ = t_7__653_ | t_7__781_;
  assign t_8__652_ = t_7__652_ | t_7__780_;
  assign t_8__651_ = t_7__651_ | t_7__779_;
  assign t_8__650_ = t_7__650_ | t_7__778_;
  assign t_8__649_ = t_7__649_ | t_7__777_;
  assign t_8__648_ = t_7__648_ | t_7__776_;
  assign t_8__647_ = t_7__647_ | t_7__775_;
  assign t_8__646_ = t_7__646_ | t_7__774_;
  assign t_8__645_ = t_7__645_ | t_7__773_;
  assign t_8__644_ = t_7__644_ | t_7__772_;
  assign t_8__643_ = t_7__643_ | t_7__771_;
  assign t_8__642_ = t_7__642_ | t_7__770_;
  assign t_8__641_ = t_7__641_ | t_7__769_;
  assign t_8__640_ = t_7__640_ | t_7__768_;
  assign t_8__639_ = t_7__639_ | t_7__767_;
  assign t_8__638_ = t_7__638_ | t_7__766_;
  assign t_8__637_ = t_7__637_ | t_7__765_;
  assign t_8__636_ = t_7__636_ | t_7__764_;
  assign t_8__635_ = t_7__635_ | t_7__763_;
  assign t_8__634_ = t_7__634_ | t_7__762_;
  assign t_8__633_ = t_7__633_ | t_7__761_;
  assign t_8__632_ = t_7__632_ | t_7__760_;
  assign t_8__631_ = t_7__631_ | t_7__759_;
  assign t_8__630_ = t_7__630_ | t_7__758_;
  assign t_8__629_ = t_7__629_ | t_7__757_;
  assign t_8__628_ = t_7__628_ | t_7__756_;
  assign t_8__627_ = t_7__627_ | t_7__755_;
  assign t_8__626_ = t_7__626_ | t_7__754_;
  assign t_8__625_ = t_7__625_ | t_7__753_;
  assign t_8__624_ = t_7__624_ | t_7__752_;
  assign t_8__623_ = t_7__623_ | t_7__751_;
  assign t_8__622_ = t_7__622_ | t_7__750_;
  assign t_8__621_ = t_7__621_ | t_7__749_;
  assign t_8__620_ = t_7__620_ | t_7__748_;
  assign t_8__619_ = t_7__619_ | t_7__747_;
  assign t_8__618_ = t_7__618_ | t_7__746_;
  assign t_8__617_ = t_7__617_ | t_7__745_;
  assign t_8__616_ = t_7__616_ | t_7__744_;
  assign t_8__615_ = t_7__615_ | t_7__743_;
  assign t_8__614_ = t_7__614_ | t_7__742_;
  assign t_8__613_ = t_7__613_ | t_7__741_;
  assign t_8__612_ = t_7__612_ | t_7__740_;
  assign t_8__611_ = t_7__611_ | t_7__739_;
  assign t_8__610_ = t_7__610_ | t_7__738_;
  assign t_8__609_ = t_7__609_ | t_7__737_;
  assign t_8__608_ = t_7__608_ | t_7__736_;
  assign t_8__607_ = t_7__607_ | t_7__735_;
  assign t_8__606_ = t_7__606_ | t_7__734_;
  assign t_8__605_ = t_7__605_ | t_7__733_;
  assign t_8__604_ = t_7__604_ | t_7__732_;
  assign t_8__603_ = t_7__603_ | t_7__731_;
  assign t_8__602_ = t_7__602_ | t_7__730_;
  assign t_8__601_ = t_7__601_ | t_7__729_;
  assign t_8__600_ = t_7__600_ | t_7__728_;
  assign t_8__599_ = t_7__599_ | t_7__727_;
  assign t_8__598_ = t_7__598_ | t_7__726_;
  assign t_8__597_ = t_7__597_ | t_7__725_;
  assign t_8__596_ = t_7__596_ | t_7__724_;
  assign t_8__595_ = t_7__595_ | t_7__723_;
  assign t_8__594_ = t_7__594_ | t_7__722_;
  assign t_8__593_ = t_7__593_ | t_7__721_;
  assign t_8__592_ = t_7__592_ | t_7__720_;
  assign t_8__591_ = t_7__591_ | t_7__719_;
  assign t_8__590_ = t_7__590_ | t_7__718_;
  assign t_8__589_ = t_7__589_ | t_7__717_;
  assign t_8__588_ = t_7__588_ | t_7__716_;
  assign t_8__587_ = t_7__587_ | t_7__715_;
  assign t_8__586_ = t_7__586_ | t_7__714_;
  assign t_8__585_ = t_7__585_ | t_7__713_;
  assign t_8__584_ = t_7__584_ | t_7__712_;
  assign t_8__583_ = t_7__583_ | t_7__711_;
  assign t_8__582_ = t_7__582_ | t_7__710_;
  assign t_8__581_ = t_7__581_ | t_7__709_;
  assign t_8__580_ = t_7__580_ | t_7__708_;
  assign t_8__579_ = t_7__579_ | t_7__707_;
  assign t_8__578_ = t_7__578_ | t_7__706_;
  assign t_8__577_ = t_7__577_ | t_7__705_;
  assign t_8__576_ = t_7__576_ | t_7__704_;
  assign t_8__575_ = t_7__575_ | t_7__703_;
  assign t_8__574_ = t_7__574_ | t_7__702_;
  assign t_8__573_ = t_7__573_ | t_7__701_;
  assign t_8__572_ = t_7__572_ | t_7__700_;
  assign t_8__571_ = t_7__571_ | t_7__699_;
  assign t_8__570_ = t_7__570_ | t_7__698_;
  assign t_8__569_ = t_7__569_ | t_7__697_;
  assign t_8__568_ = t_7__568_ | t_7__696_;
  assign t_8__567_ = t_7__567_ | t_7__695_;
  assign t_8__566_ = t_7__566_ | t_7__694_;
  assign t_8__565_ = t_7__565_ | t_7__693_;
  assign t_8__564_ = t_7__564_ | t_7__692_;
  assign t_8__563_ = t_7__563_ | t_7__691_;
  assign t_8__562_ = t_7__562_ | t_7__690_;
  assign t_8__561_ = t_7__561_ | t_7__689_;
  assign t_8__560_ = t_7__560_ | t_7__688_;
  assign t_8__559_ = t_7__559_ | t_7__687_;
  assign t_8__558_ = t_7__558_ | t_7__686_;
  assign t_8__557_ = t_7__557_ | t_7__685_;
  assign t_8__556_ = t_7__556_ | t_7__684_;
  assign t_8__555_ = t_7__555_ | t_7__683_;
  assign t_8__554_ = t_7__554_ | t_7__682_;
  assign t_8__553_ = t_7__553_ | t_7__681_;
  assign t_8__552_ = t_7__552_ | t_7__680_;
  assign t_8__551_ = t_7__551_ | t_7__679_;
  assign t_8__550_ = t_7__550_ | t_7__678_;
  assign t_8__549_ = t_7__549_ | t_7__677_;
  assign t_8__548_ = t_7__548_ | t_7__676_;
  assign t_8__547_ = t_7__547_ | t_7__675_;
  assign t_8__546_ = t_7__546_ | t_7__674_;
  assign t_8__545_ = t_7__545_ | t_7__673_;
  assign t_8__544_ = t_7__544_ | t_7__672_;
  assign t_8__543_ = t_7__543_ | t_7__671_;
  assign t_8__542_ = t_7__542_ | t_7__670_;
  assign t_8__541_ = t_7__541_ | t_7__669_;
  assign t_8__540_ = t_7__540_ | t_7__668_;
  assign t_8__539_ = t_7__539_ | t_7__667_;
  assign t_8__538_ = t_7__538_ | t_7__666_;
  assign t_8__537_ = t_7__537_ | t_7__665_;
  assign t_8__536_ = t_7__536_ | t_7__664_;
  assign t_8__535_ = t_7__535_ | t_7__663_;
  assign t_8__534_ = t_7__534_ | t_7__662_;
  assign t_8__533_ = t_7__533_ | t_7__661_;
  assign t_8__532_ = t_7__532_ | t_7__660_;
  assign t_8__531_ = t_7__531_ | t_7__659_;
  assign t_8__530_ = t_7__530_ | t_7__658_;
  assign t_8__529_ = t_7__529_ | t_7__657_;
  assign t_8__528_ = t_7__528_ | t_7__656_;
  assign t_8__527_ = t_7__527_ | t_7__655_;
  assign t_8__526_ = t_7__526_ | t_7__654_;
  assign t_8__525_ = t_7__525_ | t_7__653_;
  assign t_8__524_ = t_7__524_ | t_7__652_;
  assign t_8__523_ = t_7__523_ | t_7__651_;
  assign t_8__522_ = t_7__522_ | t_7__650_;
  assign t_8__521_ = t_7__521_ | t_7__649_;
  assign t_8__520_ = t_7__520_ | t_7__648_;
  assign t_8__519_ = t_7__519_ | t_7__647_;
  assign t_8__518_ = t_7__518_ | t_7__646_;
  assign t_8__517_ = t_7__517_ | t_7__645_;
  assign t_8__516_ = t_7__516_ | t_7__644_;
  assign t_8__515_ = t_7__515_ | t_7__643_;
  assign t_8__514_ = t_7__514_ | t_7__642_;
  assign t_8__513_ = t_7__513_ | t_7__641_;
  assign t_8__512_ = t_7__512_ | t_7__640_;
  assign t_8__511_ = t_7__511_ | t_7__639_;
  assign t_8__510_ = t_7__510_ | t_7__638_;
  assign t_8__509_ = t_7__509_ | t_7__637_;
  assign t_8__508_ = t_7__508_ | t_7__636_;
  assign t_8__507_ = t_7__507_ | t_7__635_;
  assign t_8__506_ = t_7__506_ | t_7__634_;
  assign t_8__505_ = t_7__505_ | t_7__633_;
  assign t_8__504_ = t_7__504_ | t_7__632_;
  assign t_8__503_ = t_7__503_ | t_7__631_;
  assign t_8__502_ = t_7__502_ | t_7__630_;
  assign t_8__501_ = t_7__501_ | t_7__629_;
  assign t_8__500_ = t_7__500_ | t_7__628_;
  assign t_8__499_ = t_7__499_ | t_7__627_;
  assign t_8__498_ = t_7__498_ | t_7__626_;
  assign t_8__497_ = t_7__497_ | t_7__625_;
  assign t_8__496_ = t_7__496_ | t_7__624_;
  assign t_8__495_ = t_7__495_ | t_7__623_;
  assign t_8__494_ = t_7__494_ | t_7__622_;
  assign t_8__493_ = t_7__493_ | t_7__621_;
  assign t_8__492_ = t_7__492_ | t_7__620_;
  assign t_8__491_ = t_7__491_ | t_7__619_;
  assign t_8__490_ = t_7__490_ | t_7__618_;
  assign t_8__489_ = t_7__489_ | t_7__617_;
  assign t_8__488_ = t_7__488_ | t_7__616_;
  assign t_8__487_ = t_7__487_ | t_7__615_;
  assign t_8__486_ = t_7__486_ | t_7__614_;
  assign t_8__485_ = t_7__485_ | t_7__613_;
  assign t_8__484_ = t_7__484_ | t_7__612_;
  assign t_8__483_ = t_7__483_ | t_7__611_;
  assign t_8__482_ = t_7__482_ | t_7__610_;
  assign t_8__481_ = t_7__481_ | t_7__609_;
  assign t_8__480_ = t_7__480_ | t_7__608_;
  assign t_8__479_ = t_7__479_ | t_7__607_;
  assign t_8__478_ = t_7__478_ | t_7__606_;
  assign t_8__477_ = t_7__477_ | t_7__605_;
  assign t_8__476_ = t_7__476_ | t_7__604_;
  assign t_8__475_ = t_7__475_ | t_7__603_;
  assign t_8__474_ = t_7__474_ | t_7__602_;
  assign t_8__473_ = t_7__473_ | t_7__601_;
  assign t_8__472_ = t_7__472_ | t_7__600_;
  assign t_8__471_ = t_7__471_ | t_7__599_;
  assign t_8__470_ = t_7__470_ | t_7__598_;
  assign t_8__469_ = t_7__469_ | t_7__597_;
  assign t_8__468_ = t_7__468_ | t_7__596_;
  assign t_8__467_ = t_7__467_ | t_7__595_;
  assign t_8__466_ = t_7__466_ | t_7__594_;
  assign t_8__465_ = t_7__465_ | t_7__593_;
  assign t_8__464_ = t_7__464_ | t_7__592_;
  assign t_8__463_ = t_7__463_ | t_7__591_;
  assign t_8__462_ = t_7__462_ | t_7__590_;
  assign t_8__461_ = t_7__461_ | t_7__589_;
  assign t_8__460_ = t_7__460_ | t_7__588_;
  assign t_8__459_ = t_7__459_ | t_7__587_;
  assign t_8__458_ = t_7__458_ | t_7__586_;
  assign t_8__457_ = t_7__457_ | t_7__585_;
  assign t_8__456_ = t_7__456_ | t_7__584_;
  assign t_8__455_ = t_7__455_ | t_7__583_;
  assign t_8__454_ = t_7__454_ | t_7__582_;
  assign t_8__453_ = t_7__453_ | t_7__581_;
  assign t_8__452_ = t_7__452_ | t_7__580_;
  assign t_8__451_ = t_7__451_ | t_7__579_;
  assign t_8__450_ = t_7__450_ | t_7__578_;
  assign t_8__449_ = t_7__449_ | t_7__577_;
  assign t_8__448_ = t_7__448_ | t_7__576_;
  assign t_8__447_ = t_7__447_ | t_7__575_;
  assign t_8__446_ = t_7__446_ | t_7__574_;
  assign t_8__445_ = t_7__445_ | t_7__573_;
  assign t_8__444_ = t_7__444_ | t_7__572_;
  assign t_8__443_ = t_7__443_ | t_7__571_;
  assign t_8__442_ = t_7__442_ | t_7__570_;
  assign t_8__441_ = t_7__441_ | t_7__569_;
  assign t_8__440_ = t_7__440_ | t_7__568_;
  assign t_8__439_ = t_7__439_ | t_7__567_;
  assign t_8__438_ = t_7__438_ | t_7__566_;
  assign t_8__437_ = t_7__437_ | t_7__565_;
  assign t_8__436_ = t_7__436_ | t_7__564_;
  assign t_8__435_ = t_7__435_ | t_7__563_;
  assign t_8__434_ = t_7__434_ | t_7__562_;
  assign t_8__433_ = t_7__433_ | t_7__561_;
  assign t_8__432_ = t_7__432_ | t_7__560_;
  assign t_8__431_ = t_7__431_ | t_7__559_;
  assign t_8__430_ = t_7__430_ | t_7__558_;
  assign t_8__429_ = t_7__429_ | t_7__557_;
  assign t_8__428_ = t_7__428_ | t_7__556_;
  assign t_8__427_ = t_7__427_ | t_7__555_;
  assign t_8__426_ = t_7__426_ | t_7__554_;
  assign t_8__425_ = t_7__425_ | t_7__553_;
  assign t_8__424_ = t_7__424_ | t_7__552_;
  assign t_8__423_ = t_7__423_ | t_7__551_;
  assign t_8__422_ = t_7__422_ | t_7__550_;
  assign t_8__421_ = t_7__421_ | t_7__549_;
  assign t_8__420_ = t_7__420_ | t_7__548_;
  assign t_8__419_ = t_7__419_ | t_7__547_;
  assign t_8__418_ = t_7__418_ | t_7__546_;
  assign t_8__417_ = t_7__417_ | t_7__545_;
  assign t_8__416_ = t_7__416_ | t_7__544_;
  assign t_8__415_ = t_7__415_ | t_7__543_;
  assign t_8__414_ = t_7__414_ | t_7__542_;
  assign t_8__413_ = t_7__413_ | t_7__541_;
  assign t_8__412_ = t_7__412_ | t_7__540_;
  assign t_8__411_ = t_7__411_ | t_7__539_;
  assign t_8__410_ = t_7__410_ | t_7__538_;
  assign t_8__409_ = t_7__409_ | t_7__537_;
  assign t_8__408_ = t_7__408_ | t_7__536_;
  assign t_8__407_ = t_7__407_ | t_7__535_;
  assign t_8__406_ = t_7__406_ | t_7__534_;
  assign t_8__405_ = t_7__405_ | t_7__533_;
  assign t_8__404_ = t_7__404_ | t_7__532_;
  assign t_8__403_ = t_7__403_ | t_7__531_;
  assign t_8__402_ = t_7__402_ | t_7__530_;
  assign t_8__401_ = t_7__401_ | t_7__529_;
  assign t_8__400_ = t_7__400_ | t_7__528_;
  assign t_8__399_ = t_7__399_ | t_7__527_;
  assign t_8__398_ = t_7__398_ | t_7__526_;
  assign t_8__397_ = t_7__397_ | t_7__525_;
  assign t_8__396_ = t_7__396_ | t_7__524_;
  assign t_8__395_ = t_7__395_ | t_7__523_;
  assign t_8__394_ = t_7__394_ | t_7__522_;
  assign t_8__393_ = t_7__393_ | t_7__521_;
  assign t_8__392_ = t_7__392_ | t_7__520_;
  assign t_8__391_ = t_7__391_ | t_7__519_;
  assign t_8__390_ = t_7__390_ | t_7__518_;
  assign t_8__389_ = t_7__389_ | t_7__517_;
  assign t_8__388_ = t_7__388_ | t_7__516_;
  assign t_8__387_ = t_7__387_ | t_7__515_;
  assign t_8__386_ = t_7__386_ | t_7__514_;
  assign t_8__385_ = t_7__385_ | t_7__513_;
  assign t_8__384_ = t_7__384_ | t_7__512_;
  assign t_8__383_ = t_7__383_ | t_7__511_;
  assign t_8__382_ = t_7__382_ | t_7__510_;
  assign t_8__381_ = t_7__381_ | t_7__509_;
  assign t_8__380_ = t_7__380_ | t_7__508_;
  assign t_8__379_ = t_7__379_ | t_7__507_;
  assign t_8__378_ = t_7__378_ | t_7__506_;
  assign t_8__377_ = t_7__377_ | t_7__505_;
  assign t_8__376_ = t_7__376_ | t_7__504_;
  assign t_8__375_ = t_7__375_ | t_7__503_;
  assign t_8__374_ = t_7__374_ | t_7__502_;
  assign t_8__373_ = t_7__373_ | t_7__501_;
  assign t_8__372_ = t_7__372_ | t_7__500_;
  assign t_8__371_ = t_7__371_ | t_7__499_;
  assign t_8__370_ = t_7__370_ | t_7__498_;
  assign t_8__369_ = t_7__369_ | t_7__497_;
  assign t_8__368_ = t_7__368_ | t_7__496_;
  assign t_8__367_ = t_7__367_ | t_7__495_;
  assign t_8__366_ = t_7__366_ | t_7__494_;
  assign t_8__365_ = t_7__365_ | t_7__493_;
  assign t_8__364_ = t_7__364_ | t_7__492_;
  assign t_8__363_ = t_7__363_ | t_7__491_;
  assign t_8__362_ = t_7__362_ | t_7__490_;
  assign t_8__361_ = t_7__361_ | t_7__489_;
  assign t_8__360_ = t_7__360_ | t_7__488_;
  assign t_8__359_ = t_7__359_ | t_7__487_;
  assign t_8__358_ = t_7__358_ | t_7__486_;
  assign t_8__357_ = t_7__357_ | t_7__485_;
  assign t_8__356_ = t_7__356_ | t_7__484_;
  assign t_8__355_ = t_7__355_ | t_7__483_;
  assign t_8__354_ = t_7__354_ | t_7__482_;
  assign t_8__353_ = t_7__353_ | t_7__481_;
  assign t_8__352_ = t_7__352_ | t_7__480_;
  assign t_8__351_ = t_7__351_ | t_7__479_;
  assign t_8__350_ = t_7__350_ | t_7__478_;
  assign t_8__349_ = t_7__349_ | t_7__477_;
  assign t_8__348_ = t_7__348_ | t_7__476_;
  assign t_8__347_ = t_7__347_ | t_7__475_;
  assign t_8__346_ = t_7__346_ | t_7__474_;
  assign t_8__345_ = t_7__345_ | t_7__473_;
  assign t_8__344_ = t_7__344_ | t_7__472_;
  assign t_8__343_ = t_7__343_ | t_7__471_;
  assign t_8__342_ = t_7__342_ | t_7__470_;
  assign t_8__341_ = t_7__341_ | t_7__469_;
  assign t_8__340_ = t_7__340_ | t_7__468_;
  assign t_8__339_ = t_7__339_ | t_7__467_;
  assign t_8__338_ = t_7__338_ | t_7__466_;
  assign t_8__337_ = t_7__337_ | t_7__465_;
  assign t_8__336_ = t_7__336_ | t_7__464_;
  assign t_8__335_ = t_7__335_ | t_7__463_;
  assign t_8__334_ = t_7__334_ | t_7__462_;
  assign t_8__333_ = t_7__333_ | t_7__461_;
  assign t_8__332_ = t_7__332_ | t_7__460_;
  assign t_8__331_ = t_7__331_ | t_7__459_;
  assign t_8__330_ = t_7__330_ | t_7__458_;
  assign t_8__329_ = t_7__329_ | t_7__457_;
  assign t_8__328_ = t_7__328_ | t_7__456_;
  assign t_8__327_ = t_7__327_ | t_7__455_;
  assign t_8__326_ = t_7__326_ | t_7__454_;
  assign t_8__325_ = t_7__325_ | t_7__453_;
  assign t_8__324_ = t_7__324_ | t_7__452_;
  assign t_8__323_ = t_7__323_ | t_7__451_;
  assign t_8__322_ = t_7__322_ | t_7__450_;
  assign t_8__321_ = t_7__321_ | t_7__449_;
  assign t_8__320_ = t_7__320_ | t_7__448_;
  assign t_8__319_ = t_7__319_ | t_7__447_;
  assign t_8__318_ = t_7__318_ | t_7__446_;
  assign t_8__317_ = t_7__317_ | t_7__445_;
  assign t_8__316_ = t_7__316_ | t_7__444_;
  assign t_8__315_ = t_7__315_ | t_7__443_;
  assign t_8__314_ = t_7__314_ | t_7__442_;
  assign t_8__313_ = t_7__313_ | t_7__441_;
  assign t_8__312_ = t_7__312_ | t_7__440_;
  assign t_8__311_ = t_7__311_ | t_7__439_;
  assign t_8__310_ = t_7__310_ | t_7__438_;
  assign t_8__309_ = t_7__309_ | t_7__437_;
  assign t_8__308_ = t_7__308_ | t_7__436_;
  assign t_8__307_ = t_7__307_ | t_7__435_;
  assign t_8__306_ = t_7__306_ | t_7__434_;
  assign t_8__305_ = t_7__305_ | t_7__433_;
  assign t_8__304_ = t_7__304_ | t_7__432_;
  assign t_8__303_ = t_7__303_ | t_7__431_;
  assign t_8__302_ = t_7__302_ | t_7__430_;
  assign t_8__301_ = t_7__301_ | t_7__429_;
  assign t_8__300_ = t_7__300_ | t_7__428_;
  assign t_8__299_ = t_7__299_ | t_7__427_;
  assign t_8__298_ = t_7__298_ | t_7__426_;
  assign t_8__297_ = t_7__297_ | t_7__425_;
  assign t_8__296_ = t_7__296_ | t_7__424_;
  assign t_8__295_ = t_7__295_ | t_7__423_;
  assign t_8__294_ = t_7__294_ | t_7__422_;
  assign t_8__293_ = t_7__293_ | t_7__421_;
  assign t_8__292_ = t_7__292_ | t_7__420_;
  assign t_8__291_ = t_7__291_ | t_7__419_;
  assign t_8__290_ = t_7__290_ | t_7__418_;
  assign t_8__289_ = t_7__289_ | t_7__417_;
  assign t_8__288_ = t_7__288_ | t_7__416_;
  assign t_8__287_ = t_7__287_ | t_7__415_;
  assign t_8__286_ = t_7__286_ | t_7__414_;
  assign t_8__285_ = t_7__285_ | t_7__413_;
  assign t_8__284_ = t_7__284_ | t_7__412_;
  assign t_8__283_ = t_7__283_ | t_7__411_;
  assign t_8__282_ = t_7__282_ | t_7__410_;
  assign t_8__281_ = t_7__281_ | t_7__409_;
  assign t_8__280_ = t_7__280_ | t_7__408_;
  assign t_8__279_ = t_7__279_ | t_7__407_;
  assign t_8__278_ = t_7__278_ | t_7__406_;
  assign t_8__277_ = t_7__277_ | t_7__405_;
  assign t_8__276_ = t_7__276_ | t_7__404_;
  assign t_8__275_ = t_7__275_ | t_7__403_;
  assign t_8__274_ = t_7__274_ | t_7__402_;
  assign t_8__273_ = t_7__273_ | t_7__401_;
  assign t_8__272_ = t_7__272_ | t_7__400_;
  assign t_8__271_ = t_7__271_ | t_7__399_;
  assign t_8__270_ = t_7__270_ | t_7__398_;
  assign t_8__269_ = t_7__269_ | t_7__397_;
  assign t_8__268_ = t_7__268_ | t_7__396_;
  assign t_8__267_ = t_7__267_ | t_7__395_;
  assign t_8__266_ = t_7__266_ | t_7__394_;
  assign t_8__265_ = t_7__265_ | t_7__393_;
  assign t_8__264_ = t_7__264_ | t_7__392_;
  assign t_8__263_ = t_7__263_ | t_7__391_;
  assign t_8__262_ = t_7__262_ | t_7__390_;
  assign t_8__261_ = t_7__261_ | t_7__389_;
  assign t_8__260_ = t_7__260_ | t_7__388_;
  assign t_8__259_ = t_7__259_ | t_7__387_;
  assign t_8__258_ = t_7__258_ | t_7__386_;
  assign t_8__257_ = t_7__257_ | t_7__385_;
  assign t_8__256_ = t_7__256_ | t_7__384_;
  assign t_8__255_ = t_7__255_ | t_7__383_;
  assign t_8__254_ = t_7__254_ | t_7__382_;
  assign t_8__253_ = t_7__253_ | t_7__381_;
  assign t_8__252_ = t_7__252_ | t_7__380_;
  assign t_8__251_ = t_7__251_ | t_7__379_;
  assign t_8__250_ = t_7__250_ | t_7__378_;
  assign t_8__249_ = t_7__249_ | t_7__377_;
  assign t_8__248_ = t_7__248_ | t_7__376_;
  assign t_8__247_ = t_7__247_ | t_7__375_;
  assign t_8__246_ = t_7__246_ | t_7__374_;
  assign t_8__245_ = t_7__245_ | t_7__373_;
  assign t_8__244_ = t_7__244_ | t_7__372_;
  assign t_8__243_ = t_7__243_ | t_7__371_;
  assign t_8__242_ = t_7__242_ | t_7__370_;
  assign t_8__241_ = t_7__241_ | t_7__369_;
  assign t_8__240_ = t_7__240_ | t_7__368_;
  assign t_8__239_ = t_7__239_ | t_7__367_;
  assign t_8__238_ = t_7__238_ | t_7__366_;
  assign t_8__237_ = t_7__237_ | t_7__365_;
  assign t_8__236_ = t_7__236_ | t_7__364_;
  assign t_8__235_ = t_7__235_ | t_7__363_;
  assign t_8__234_ = t_7__234_ | t_7__362_;
  assign t_8__233_ = t_7__233_ | t_7__361_;
  assign t_8__232_ = t_7__232_ | t_7__360_;
  assign t_8__231_ = t_7__231_ | t_7__359_;
  assign t_8__230_ = t_7__230_ | t_7__358_;
  assign t_8__229_ = t_7__229_ | t_7__357_;
  assign t_8__228_ = t_7__228_ | t_7__356_;
  assign t_8__227_ = t_7__227_ | t_7__355_;
  assign t_8__226_ = t_7__226_ | t_7__354_;
  assign t_8__225_ = t_7__225_ | t_7__353_;
  assign t_8__224_ = t_7__224_ | t_7__352_;
  assign t_8__223_ = t_7__223_ | t_7__351_;
  assign t_8__222_ = t_7__222_ | t_7__350_;
  assign t_8__221_ = t_7__221_ | t_7__349_;
  assign t_8__220_ = t_7__220_ | t_7__348_;
  assign t_8__219_ = t_7__219_ | t_7__347_;
  assign t_8__218_ = t_7__218_ | t_7__346_;
  assign t_8__217_ = t_7__217_ | t_7__345_;
  assign t_8__216_ = t_7__216_ | t_7__344_;
  assign t_8__215_ = t_7__215_ | t_7__343_;
  assign t_8__214_ = t_7__214_ | t_7__342_;
  assign t_8__213_ = t_7__213_ | t_7__341_;
  assign t_8__212_ = t_7__212_ | t_7__340_;
  assign t_8__211_ = t_7__211_ | t_7__339_;
  assign t_8__210_ = t_7__210_ | t_7__338_;
  assign t_8__209_ = t_7__209_ | t_7__337_;
  assign t_8__208_ = t_7__208_ | t_7__336_;
  assign t_8__207_ = t_7__207_ | t_7__335_;
  assign t_8__206_ = t_7__206_ | t_7__334_;
  assign t_8__205_ = t_7__205_ | t_7__333_;
  assign t_8__204_ = t_7__204_ | t_7__332_;
  assign t_8__203_ = t_7__203_ | t_7__331_;
  assign t_8__202_ = t_7__202_ | t_7__330_;
  assign t_8__201_ = t_7__201_ | t_7__329_;
  assign t_8__200_ = t_7__200_ | t_7__328_;
  assign t_8__199_ = t_7__199_ | t_7__327_;
  assign t_8__198_ = t_7__198_ | t_7__326_;
  assign t_8__197_ = t_7__197_ | t_7__325_;
  assign t_8__196_ = t_7__196_ | t_7__324_;
  assign t_8__195_ = t_7__195_ | t_7__323_;
  assign t_8__194_ = t_7__194_ | t_7__322_;
  assign t_8__193_ = t_7__193_ | t_7__321_;
  assign t_8__192_ = t_7__192_ | t_7__320_;
  assign t_8__191_ = t_7__191_ | t_7__319_;
  assign t_8__190_ = t_7__190_ | t_7__318_;
  assign t_8__189_ = t_7__189_ | t_7__317_;
  assign t_8__188_ = t_7__188_ | t_7__316_;
  assign t_8__187_ = t_7__187_ | t_7__315_;
  assign t_8__186_ = t_7__186_ | t_7__314_;
  assign t_8__185_ = t_7__185_ | t_7__313_;
  assign t_8__184_ = t_7__184_ | t_7__312_;
  assign t_8__183_ = t_7__183_ | t_7__311_;
  assign t_8__182_ = t_7__182_ | t_7__310_;
  assign t_8__181_ = t_7__181_ | t_7__309_;
  assign t_8__180_ = t_7__180_ | t_7__308_;
  assign t_8__179_ = t_7__179_ | t_7__307_;
  assign t_8__178_ = t_7__178_ | t_7__306_;
  assign t_8__177_ = t_7__177_ | t_7__305_;
  assign t_8__176_ = t_7__176_ | t_7__304_;
  assign t_8__175_ = t_7__175_ | t_7__303_;
  assign t_8__174_ = t_7__174_ | t_7__302_;
  assign t_8__173_ = t_7__173_ | t_7__301_;
  assign t_8__172_ = t_7__172_ | t_7__300_;
  assign t_8__171_ = t_7__171_ | t_7__299_;
  assign t_8__170_ = t_7__170_ | t_7__298_;
  assign t_8__169_ = t_7__169_ | t_7__297_;
  assign t_8__168_ = t_7__168_ | t_7__296_;
  assign t_8__167_ = t_7__167_ | t_7__295_;
  assign t_8__166_ = t_7__166_ | t_7__294_;
  assign t_8__165_ = t_7__165_ | t_7__293_;
  assign t_8__164_ = t_7__164_ | t_7__292_;
  assign t_8__163_ = t_7__163_ | t_7__291_;
  assign t_8__162_ = t_7__162_ | t_7__290_;
  assign t_8__161_ = t_7__161_ | t_7__289_;
  assign t_8__160_ = t_7__160_ | t_7__288_;
  assign t_8__159_ = t_7__159_ | t_7__287_;
  assign t_8__158_ = t_7__158_ | t_7__286_;
  assign t_8__157_ = t_7__157_ | t_7__285_;
  assign t_8__156_ = t_7__156_ | t_7__284_;
  assign t_8__155_ = t_7__155_ | t_7__283_;
  assign t_8__154_ = t_7__154_ | t_7__282_;
  assign t_8__153_ = t_7__153_ | t_7__281_;
  assign t_8__152_ = t_7__152_ | t_7__280_;
  assign t_8__151_ = t_7__151_ | t_7__279_;
  assign t_8__150_ = t_7__150_ | t_7__278_;
  assign t_8__149_ = t_7__149_ | t_7__277_;
  assign t_8__148_ = t_7__148_ | t_7__276_;
  assign t_8__147_ = t_7__147_ | t_7__275_;
  assign t_8__146_ = t_7__146_ | t_7__274_;
  assign t_8__145_ = t_7__145_ | t_7__273_;
  assign t_8__144_ = t_7__144_ | t_7__272_;
  assign t_8__143_ = t_7__143_ | t_7__271_;
  assign t_8__142_ = t_7__142_ | t_7__270_;
  assign t_8__141_ = t_7__141_ | t_7__269_;
  assign t_8__140_ = t_7__140_ | t_7__268_;
  assign t_8__139_ = t_7__139_ | t_7__267_;
  assign t_8__138_ = t_7__138_ | t_7__266_;
  assign t_8__137_ = t_7__137_ | t_7__265_;
  assign t_8__136_ = t_7__136_ | t_7__264_;
  assign t_8__135_ = t_7__135_ | t_7__263_;
  assign t_8__134_ = t_7__134_ | t_7__262_;
  assign t_8__133_ = t_7__133_ | t_7__261_;
  assign t_8__132_ = t_7__132_ | t_7__260_;
  assign t_8__131_ = t_7__131_ | t_7__259_;
  assign t_8__130_ = t_7__130_ | t_7__258_;
  assign t_8__129_ = t_7__129_ | t_7__257_;
  assign t_8__128_ = t_7__128_ | t_7__256_;
  assign t_8__127_ = t_7__127_ | t_7__255_;
  assign t_8__126_ = t_7__126_ | t_7__254_;
  assign t_8__125_ = t_7__125_ | t_7__253_;
  assign t_8__124_ = t_7__124_ | t_7__252_;
  assign t_8__123_ = t_7__123_ | t_7__251_;
  assign t_8__122_ = t_7__122_ | t_7__250_;
  assign t_8__121_ = t_7__121_ | t_7__249_;
  assign t_8__120_ = t_7__120_ | t_7__248_;
  assign t_8__119_ = t_7__119_ | t_7__247_;
  assign t_8__118_ = t_7__118_ | t_7__246_;
  assign t_8__117_ = t_7__117_ | t_7__245_;
  assign t_8__116_ = t_7__116_ | t_7__244_;
  assign t_8__115_ = t_7__115_ | t_7__243_;
  assign t_8__114_ = t_7__114_ | t_7__242_;
  assign t_8__113_ = t_7__113_ | t_7__241_;
  assign t_8__112_ = t_7__112_ | t_7__240_;
  assign t_8__111_ = t_7__111_ | t_7__239_;
  assign t_8__110_ = t_7__110_ | t_7__238_;
  assign t_8__109_ = t_7__109_ | t_7__237_;
  assign t_8__108_ = t_7__108_ | t_7__236_;
  assign t_8__107_ = t_7__107_ | t_7__235_;
  assign t_8__106_ = t_7__106_ | t_7__234_;
  assign t_8__105_ = t_7__105_ | t_7__233_;
  assign t_8__104_ = t_7__104_ | t_7__232_;
  assign t_8__103_ = t_7__103_ | t_7__231_;
  assign t_8__102_ = t_7__102_ | t_7__230_;
  assign t_8__101_ = t_7__101_ | t_7__229_;
  assign t_8__100_ = t_7__100_ | t_7__228_;
  assign t_8__99_ = t_7__99_ | t_7__227_;
  assign t_8__98_ = t_7__98_ | t_7__226_;
  assign t_8__97_ = t_7__97_ | t_7__225_;
  assign t_8__96_ = t_7__96_ | t_7__224_;
  assign t_8__95_ = t_7__95_ | t_7__223_;
  assign t_8__94_ = t_7__94_ | t_7__222_;
  assign t_8__93_ = t_7__93_ | t_7__221_;
  assign t_8__92_ = t_7__92_ | t_7__220_;
  assign t_8__91_ = t_7__91_ | t_7__219_;
  assign t_8__90_ = t_7__90_ | t_7__218_;
  assign t_8__89_ = t_7__89_ | t_7__217_;
  assign t_8__88_ = t_7__88_ | t_7__216_;
  assign t_8__87_ = t_7__87_ | t_7__215_;
  assign t_8__86_ = t_7__86_ | t_7__214_;
  assign t_8__85_ = t_7__85_ | t_7__213_;
  assign t_8__84_ = t_7__84_ | t_7__212_;
  assign t_8__83_ = t_7__83_ | t_7__211_;
  assign t_8__82_ = t_7__82_ | t_7__210_;
  assign t_8__81_ = t_7__81_ | t_7__209_;
  assign t_8__80_ = t_7__80_ | t_7__208_;
  assign t_8__79_ = t_7__79_ | t_7__207_;
  assign t_8__78_ = t_7__78_ | t_7__206_;
  assign t_8__77_ = t_7__77_ | t_7__205_;
  assign t_8__76_ = t_7__76_ | t_7__204_;
  assign t_8__75_ = t_7__75_ | t_7__203_;
  assign t_8__74_ = t_7__74_ | t_7__202_;
  assign t_8__73_ = t_7__73_ | t_7__201_;
  assign t_8__72_ = t_7__72_ | t_7__200_;
  assign t_8__71_ = t_7__71_ | t_7__199_;
  assign t_8__70_ = t_7__70_ | t_7__198_;
  assign t_8__69_ = t_7__69_ | t_7__197_;
  assign t_8__68_ = t_7__68_ | t_7__196_;
  assign t_8__67_ = t_7__67_ | t_7__195_;
  assign t_8__66_ = t_7__66_ | t_7__194_;
  assign t_8__65_ = t_7__65_ | t_7__193_;
  assign t_8__64_ = t_7__64_ | t_7__192_;
  assign t_8__63_ = t_7__63_ | t_7__191_;
  assign t_8__62_ = t_7__62_ | t_7__190_;
  assign t_8__61_ = t_7__61_ | t_7__189_;
  assign t_8__60_ = t_7__60_ | t_7__188_;
  assign t_8__59_ = t_7__59_ | t_7__187_;
  assign t_8__58_ = t_7__58_ | t_7__186_;
  assign t_8__57_ = t_7__57_ | t_7__185_;
  assign t_8__56_ = t_7__56_ | t_7__184_;
  assign t_8__55_ = t_7__55_ | t_7__183_;
  assign t_8__54_ = t_7__54_ | t_7__182_;
  assign t_8__53_ = t_7__53_ | t_7__181_;
  assign t_8__52_ = t_7__52_ | t_7__180_;
  assign t_8__51_ = t_7__51_ | t_7__179_;
  assign t_8__50_ = t_7__50_ | t_7__178_;
  assign t_8__49_ = t_7__49_ | t_7__177_;
  assign t_8__48_ = t_7__48_ | t_7__176_;
  assign t_8__47_ = t_7__47_ | t_7__175_;
  assign t_8__46_ = t_7__46_ | t_7__174_;
  assign t_8__45_ = t_7__45_ | t_7__173_;
  assign t_8__44_ = t_7__44_ | t_7__172_;
  assign t_8__43_ = t_7__43_ | t_7__171_;
  assign t_8__42_ = t_7__42_ | t_7__170_;
  assign t_8__41_ = t_7__41_ | t_7__169_;
  assign t_8__40_ = t_7__40_ | t_7__168_;
  assign t_8__39_ = t_7__39_ | t_7__167_;
  assign t_8__38_ = t_7__38_ | t_7__166_;
  assign t_8__37_ = t_7__37_ | t_7__165_;
  assign t_8__36_ = t_7__36_ | t_7__164_;
  assign t_8__35_ = t_7__35_ | t_7__163_;
  assign t_8__34_ = t_7__34_ | t_7__162_;
  assign t_8__33_ = t_7__33_ | t_7__161_;
  assign t_8__32_ = t_7__32_ | t_7__160_;
  assign t_8__31_ = t_7__31_ | t_7__159_;
  assign t_8__30_ = t_7__30_ | t_7__158_;
  assign t_8__29_ = t_7__29_ | t_7__157_;
  assign t_8__28_ = t_7__28_ | t_7__156_;
  assign t_8__27_ = t_7__27_ | t_7__155_;
  assign t_8__26_ = t_7__26_ | t_7__154_;
  assign t_8__25_ = t_7__25_ | t_7__153_;
  assign t_8__24_ = t_7__24_ | t_7__152_;
  assign t_8__23_ = t_7__23_ | t_7__151_;
  assign t_8__22_ = t_7__22_ | t_7__150_;
  assign t_8__21_ = t_7__21_ | t_7__149_;
  assign t_8__20_ = t_7__20_ | t_7__148_;
  assign t_8__19_ = t_7__19_ | t_7__147_;
  assign t_8__18_ = t_7__18_ | t_7__146_;
  assign t_8__17_ = t_7__17_ | t_7__145_;
  assign t_8__16_ = t_7__16_ | t_7__144_;
  assign t_8__15_ = t_7__15_ | t_7__143_;
  assign t_8__14_ = t_7__14_ | t_7__142_;
  assign t_8__13_ = t_7__13_ | t_7__141_;
  assign t_8__12_ = t_7__12_ | t_7__140_;
  assign t_8__11_ = t_7__11_ | t_7__139_;
  assign t_8__10_ = t_7__10_ | t_7__138_;
  assign t_8__9_ = t_7__9_ | t_7__137_;
  assign t_8__8_ = t_7__8_ | t_7__136_;
  assign t_8__7_ = t_7__7_ | t_7__135_;
  assign t_8__6_ = t_7__6_ | t_7__134_;
  assign t_8__5_ = t_7__5_ | t_7__133_;
  assign t_8__4_ = t_7__4_ | t_7__132_;
  assign t_8__3_ = t_7__3_ | t_7__131_;
  assign t_8__2_ = t_7__2_ | t_7__130_;
  assign t_8__1_ = t_7__1_ | t_7__129_;
  assign t_8__0_ = t_7__0_ | t_7__128_;
  assign t_9__1023_ = t_8__1023_ | 1'b0;
  assign t_9__1022_ = t_8__1022_ | 1'b0;
  assign t_9__1021_ = t_8__1021_ | 1'b0;
  assign t_9__1020_ = t_8__1020_ | 1'b0;
  assign t_9__1019_ = t_8__1019_ | 1'b0;
  assign t_9__1018_ = t_8__1018_ | 1'b0;
  assign t_9__1017_ = t_8__1017_ | 1'b0;
  assign t_9__1016_ = t_8__1016_ | 1'b0;
  assign t_9__1015_ = t_8__1015_ | 1'b0;
  assign t_9__1014_ = t_8__1014_ | 1'b0;
  assign t_9__1013_ = t_8__1013_ | 1'b0;
  assign t_9__1012_ = t_8__1012_ | 1'b0;
  assign t_9__1011_ = t_8__1011_ | 1'b0;
  assign t_9__1010_ = t_8__1010_ | 1'b0;
  assign t_9__1009_ = t_8__1009_ | 1'b0;
  assign t_9__1008_ = t_8__1008_ | 1'b0;
  assign t_9__1007_ = t_8__1007_ | 1'b0;
  assign t_9__1006_ = t_8__1006_ | 1'b0;
  assign t_9__1005_ = t_8__1005_ | 1'b0;
  assign t_9__1004_ = t_8__1004_ | 1'b0;
  assign t_9__1003_ = t_8__1003_ | 1'b0;
  assign t_9__1002_ = t_8__1002_ | 1'b0;
  assign t_9__1001_ = t_8__1001_ | 1'b0;
  assign t_9__1000_ = t_8__1000_ | 1'b0;
  assign t_9__999_ = t_8__999_ | 1'b0;
  assign t_9__998_ = t_8__998_ | 1'b0;
  assign t_9__997_ = t_8__997_ | 1'b0;
  assign t_9__996_ = t_8__996_ | 1'b0;
  assign t_9__995_ = t_8__995_ | 1'b0;
  assign t_9__994_ = t_8__994_ | 1'b0;
  assign t_9__993_ = t_8__993_ | 1'b0;
  assign t_9__992_ = t_8__992_ | 1'b0;
  assign t_9__991_ = t_8__991_ | 1'b0;
  assign t_9__990_ = t_8__990_ | 1'b0;
  assign t_9__989_ = t_8__989_ | 1'b0;
  assign t_9__988_ = t_8__988_ | 1'b0;
  assign t_9__987_ = t_8__987_ | 1'b0;
  assign t_9__986_ = t_8__986_ | 1'b0;
  assign t_9__985_ = t_8__985_ | 1'b0;
  assign t_9__984_ = t_8__984_ | 1'b0;
  assign t_9__983_ = t_8__983_ | 1'b0;
  assign t_9__982_ = t_8__982_ | 1'b0;
  assign t_9__981_ = t_8__981_ | 1'b0;
  assign t_9__980_ = t_8__980_ | 1'b0;
  assign t_9__979_ = t_8__979_ | 1'b0;
  assign t_9__978_ = t_8__978_ | 1'b0;
  assign t_9__977_ = t_8__977_ | 1'b0;
  assign t_9__976_ = t_8__976_ | 1'b0;
  assign t_9__975_ = t_8__975_ | 1'b0;
  assign t_9__974_ = t_8__974_ | 1'b0;
  assign t_9__973_ = t_8__973_ | 1'b0;
  assign t_9__972_ = t_8__972_ | 1'b0;
  assign t_9__971_ = t_8__971_ | 1'b0;
  assign t_9__970_ = t_8__970_ | 1'b0;
  assign t_9__969_ = t_8__969_ | 1'b0;
  assign t_9__968_ = t_8__968_ | 1'b0;
  assign t_9__967_ = t_8__967_ | 1'b0;
  assign t_9__966_ = t_8__966_ | 1'b0;
  assign t_9__965_ = t_8__965_ | 1'b0;
  assign t_9__964_ = t_8__964_ | 1'b0;
  assign t_9__963_ = t_8__963_ | 1'b0;
  assign t_9__962_ = t_8__962_ | 1'b0;
  assign t_9__961_ = t_8__961_ | 1'b0;
  assign t_9__960_ = t_8__960_ | 1'b0;
  assign t_9__959_ = t_8__959_ | 1'b0;
  assign t_9__958_ = t_8__958_ | 1'b0;
  assign t_9__957_ = t_8__957_ | 1'b0;
  assign t_9__956_ = t_8__956_ | 1'b0;
  assign t_9__955_ = t_8__955_ | 1'b0;
  assign t_9__954_ = t_8__954_ | 1'b0;
  assign t_9__953_ = t_8__953_ | 1'b0;
  assign t_9__952_ = t_8__952_ | 1'b0;
  assign t_9__951_ = t_8__951_ | 1'b0;
  assign t_9__950_ = t_8__950_ | 1'b0;
  assign t_9__949_ = t_8__949_ | 1'b0;
  assign t_9__948_ = t_8__948_ | 1'b0;
  assign t_9__947_ = t_8__947_ | 1'b0;
  assign t_9__946_ = t_8__946_ | 1'b0;
  assign t_9__945_ = t_8__945_ | 1'b0;
  assign t_9__944_ = t_8__944_ | 1'b0;
  assign t_9__943_ = t_8__943_ | 1'b0;
  assign t_9__942_ = t_8__942_ | 1'b0;
  assign t_9__941_ = t_8__941_ | 1'b0;
  assign t_9__940_ = t_8__940_ | 1'b0;
  assign t_9__939_ = t_8__939_ | 1'b0;
  assign t_9__938_ = t_8__938_ | 1'b0;
  assign t_9__937_ = t_8__937_ | 1'b0;
  assign t_9__936_ = t_8__936_ | 1'b0;
  assign t_9__935_ = t_8__935_ | 1'b0;
  assign t_9__934_ = t_8__934_ | 1'b0;
  assign t_9__933_ = t_8__933_ | 1'b0;
  assign t_9__932_ = t_8__932_ | 1'b0;
  assign t_9__931_ = t_8__931_ | 1'b0;
  assign t_9__930_ = t_8__930_ | 1'b0;
  assign t_9__929_ = t_8__929_ | 1'b0;
  assign t_9__928_ = t_8__928_ | 1'b0;
  assign t_9__927_ = t_8__927_ | 1'b0;
  assign t_9__926_ = t_8__926_ | 1'b0;
  assign t_9__925_ = t_8__925_ | 1'b0;
  assign t_9__924_ = t_8__924_ | 1'b0;
  assign t_9__923_ = t_8__923_ | 1'b0;
  assign t_9__922_ = t_8__922_ | 1'b0;
  assign t_9__921_ = t_8__921_ | 1'b0;
  assign t_9__920_ = t_8__920_ | 1'b0;
  assign t_9__919_ = t_8__919_ | 1'b0;
  assign t_9__918_ = t_8__918_ | 1'b0;
  assign t_9__917_ = t_8__917_ | 1'b0;
  assign t_9__916_ = t_8__916_ | 1'b0;
  assign t_9__915_ = t_8__915_ | 1'b0;
  assign t_9__914_ = t_8__914_ | 1'b0;
  assign t_9__913_ = t_8__913_ | 1'b0;
  assign t_9__912_ = t_8__912_ | 1'b0;
  assign t_9__911_ = t_8__911_ | 1'b0;
  assign t_9__910_ = t_8__910_ | 1'b0;
  assign t_9__909_ = t_8__909_ | 1'b0;
  assign t_9__908_ = t_8__908_ | 1'b0;
  assign t_9__907_ = t_8__907_ | 1'b0;
  assign t_9__906_ = t_8__906_ | 1'b0;
  assign t_9__905_ = t_8__905_ | 1'b0;
  assign t_9__904_ = t_8__904_ | 1'b0;
  assign t_9__903_ = t_8__903_ | 1'b0;
  assign t_9__902_ = t_8__902_ | 1'b0;
  assign t_9__901_ = t_8__901_ | 1'b0;
  assign t_9__900_ = t_8__900_ | 1'b0;
  assign t_9__899_ = t_8__899_ | 1'b0;
  assign t_9__898_ = t_8__898_ | 1'b0;
  assign t_9__897_ = t_8__897_ | 1'b0;
  assign t_9__896_ = t_8__896_ | 1'b0;
  assign t_9__895_ = t_8__895_ | 1'b0;
  assign t_9__894_ = t_8__894_ | 1'b0;
  assign t_9__893_ = t_8__893_ | 1'b0;
  assign t_9__892_ = t_8__892_ | 1'b0;
  assign t_9__891_ = t_8__891_ | 1'b0;
  assign t_9__890_ = t_8__890_ | 1'b0;
  assign t_9__889_ = t_8__889_ | 1'b0;
  assign t_9__888_ = t_8__888_ | 1'b0;
  assign t_9__887_ = t_8__887_ | 1'b0;
  assign t_9__886_ = t_8__886_ | 1'b0;
  assign t_9__885_ = t_8__885_ | 1'b0;
  assign t_9__884_ = t_8__884_ | 1'b0;
  assign t_9__883_ = t_8__883_ | 1'b0;
  assign t_9__882_ = t_8__882_ | 1'b0;
  assign t_9__881_ = t_8__881_ | 1'b0;
  assign t_9__880_ = t_8__880_ | 1'b0;
  assign t_9__879_ = t_8__879_ | 1'b0;
  assign t_9__878_ = t_8__878_ | 1'b0;
  assign t_9__877_ = t_8__877_ | 1'b0;
  assign t_9__876_ = t_8__876_ | 1'b0;
  assign t_9__875_ = t_8__875_ | 1'b0;
  assign t_9__874_ = t_8__874_ | 1'b0;
  assign t_9__873_ = t_8__873_ | 1'b0;
  assign t_9__872_ = t_8__872_ | 1'b0;
  assign t_9__871_ = t_8__871_ | 1'b0;
  assign t_9__870_ = t_8__870_ | 1'b0;
  assign t_9__869_ = t_8__869_ | 1'b0;
  assign t_9__868_ = t_8__868_ | 1'b0;
  assign t_9__867_ = t_8__867_ | 1'b0;
  assign t_9__866_ = t_8__866_ | 1'b0;
  assign t_9__865_ = t_8__865_ | 1'b0;
  assign t_9__864_ = t_8__864_ | 1'b0;
  assign t_9__863_ = t_8__863_ | 1'b0;
  assign t_9__862_ = t_8__862_ | 1'b0;
  assign t_9__861_ = t_8__861_ | 1'b0;
  assign t_9__860_ = t_8__860_ | 1'b0;
  assign t_9__859_ = t_8__859_ | 1'b0;
  assign t_9__858_ = t_8__858_ | 1'b0;
  assign t_9__857_ = t_8__857_ | 1'b0;
  assign t_9__856_ = t_8__856_ | 1'b0;
  assign t_9__855_ = t_8__855_ | 1'b0;
  assign t_9__854_ = t_8__854_ | 1'b0;
  assign t_9__853_ = t_8__853_ | 1'b0;
  assign t_9__852_ = t_8__852_ | 1'b0;
  assign t_9__851_ = t_8__851_ | 1'b0;
  assign t_9__850_ = t_8__850_ | 1'b0;
  assign t_9__849_ = t_8__849_ | 1'b0;
  assign t_9__848_ = t_8__848_ | 1'b0;
  assign t_9__847_ = t_8__847_ | 1'b0;
  assign t_9__846_ = t_8__846_ | 1'b0;
  assign t_9__845_ = t_8__845_ | 1'b0;
  assign t_9__844_ = t_8__844_ | 1'b0;
  assign t_9__843_ = t_8__843_ | 1'b0;
  assign t_9__842_ = t_8__842_ | 1'b0;
  assign t_9__841_ = t_8__841_ | 1'b0;
  assign t_9__840_ = t_8__840_ | 1'b0;
  assign t_9__839_ = t_8__839_ | 1'b0;
  assign t_9__838_ = t_8__838_ | 1'b0;
  assign t_9__837_ = t_8__837_ | 1'b0;
  assign t_9__836_ = t_8__836_ | 1'b0;
  assign t_9__835_ = t_8__835_ | 1'b0;
  assign t_9__834_ = t_8__834_ | 1'b0;
  assign t_9__833_ = t_8__833_ | 1'b0;
  assign t_9__832_ = t_8__832_ | 1'b0;
  assign t_9__831_ = t_8__831_ | 1'b0;
  assign t_9__830_ = t_8__830_ | 1'b0;
  assign t_9__829_ = t_8__829_ | 1'b0;
  assign t_9__828_ = t_8__828_ | 1'b0;
  assign t_9__827_ = t_8__827_ | 1'b0;
  assign t_9__826_ = t_8__826_ | 1'b0;
  assign t_9__825_ = t_8__825_ | 1'b0;
  assign t_9__824_ = t_8__824_ | 1'b0;
  assign t_9__823_ = t_8__823_ | 1'b0;
  assign t_9__822_ = t_8__822_ | 1'b0;
  assign t_9__821_ = t_8__821_ | 1'b0;
  assign t_9__820_ = t_8__820_ | 1'b0;
  assign t_9__819_ = t_8__819_ | 1'b0;
  assign t_9__818_ = t_8__818_ | 1'b0;
  assign t_9__817_ = t_8__817_ | 1'b0;
  assign t_9__816_ = t_8__816_ | 1'b0;
  assign t_9__815_ = t_8__815_ | 1'b0;
  assign t_9__814_ = t_8__814_ | 1'b0;
  assign t_9__813_ = t_8__813_ | 1'b0;
  assign t_9__812_ = t_8__812_ | 1'b0;
  assign t_9__811_ = t_8__811_ | 1'b0;
  assign t_9__810_ = t_8__810_ | 1'b0;
  assign t_9__809_ = t_8__809_ | 1'b0;
  assign t_9__808_ = t_8__808_ | 1'b0;
  assign t_9__807_ = t_8__807_ | 1'b0;
  assign t_9__806_ = t_8__806_ | 1'b0;
  assign t_9__805_ = t_8__805_ | 1'b0;
  assign t_9__804_ = t_8__804_ | 1'b0;
  assign t_9__803_ = t_8__803_ | 1'b0;
  assign t_9__802_ = t_8__802_ | 1'b0;
  assign t_9__801_ = t_8__801_ | 1'b0;
  assign t_9__800_ = t_8__800_ | 1'b0;
  assign t_9__799_ = t_8__799_ | 1'b0;
  assign t_9__798_ = t_8__798_ | 1'b0;
  assign t_9__797_ = t_8__797_ | 1'b0;
  assign t_9__796_ = t_8__796_ | 1'b0;
  assign t_9__795_ = t_8__795_ | 1'b0;
  assign t_9__794_ = t_8__794_ | 1'b0;
  assign t_9__793_ = t_8__793_ | 1'b0;
  assign t_9__792_ = t_8__792_ | 1'b0;
  assign t_9__791_ = t_8__791_ | 1'b0;
  assign t_9__790_ = t_8__790_ | 1'b0;
  assign t_9__789_ = t_8__789_ | 1'b0;
  assign t_9__788_ = t_8__788_ | 1'b0;
  assign t_9__787_ = t_8__787_ | 1'b0;
  assign t_9__786_ = t_8__786_ | 1'b0;
  assign t_9__785_ = t_8__785_ | 1'b0;
  assign t_9__784_ = t_8__784_ | 1'b0;
  assign t_9__783_ = t_8__783_ | 1'b0;
  assign t_9__782_ = t_8__782_ | 1'b0;
  assign t_9__781_ = t_8__781_ | 1'b0;
  assign t_9__780_ = t_8__780_ | 1'b0;
  assign t_9__779_ = t_8__779_ | 1'b0;
  assign t_9__778_ = t_8__778_ | 1'b0;
  assign t_9__777_ = t_8__777_ | 1'b0;
  assign t_9__776_ = t_8__776_ | 1'b0;
  assign t_9__775_ = t_8__775_ | 1'b0;
  assign t_9__774_ = t_8__774_ | 1'b0;
  assign t_9__773_ = t_8__773_ | 1'b0;
  assign t_9__772_ = t_8__772_ | 1'b0;
  assign t_9__771_ = t_8__771_ | 1'b0;
  assign t_9__770_ = t_8__770_ | 1'b0;
  assign t_9__769_ = t_8__769_ | 1'b0;
  assign t_9__768_ = t_8__768_ | 1'b0;
  assign t_9__767_ = t_8__767_ | t_8__1023_;
  assign t_9__766_ = t_8__766_ | t_8__1022_;
  assign t_9__765_ = t_8__765_ | t_8__1021_;
  assign t_9__764_ = t_8__764_ | t_8__1020_;
  assign t_9__763_ = t_8__763_ | t_8__1019_;
  assign t_9__762_ = t_8__762_ | t_8__1018_;
  assign t_9__761_ = t_8__761_ | t_8__1017_;
  assign t_9__760_ = t_8__760_ | t_8__1016_;
  assign t_9__759_ = t_8__759_ | t_8__1015_;
  assign t_9__758_ = t_8__758_ | t_8__1014_;
  assign t_9__757_ = t_8__757_ | t_8__1013_;
  assign t_9__756_ = t_8__756_ | t_8__1012_;
  assign t_9__755_ = t_8__755_ | t_8__1011_;
  assign t_9__754_ = t_8__754_ | t_8__1010_;
  assign t_9__753_ = t_8__753_ | t_8__1009_;
  assign t_9__752_ = t_8__752_ | t_8__1008_;
  assign t_9__751_ = t_8__751_ | t_8__1007_;
  assign t_9__750_ = t_8__750_ | t_8__1006_;
  assign t_9__749_ = t_8__749_ | t_8__1005_;
  assign t_9__748_ = t_8__748_ | t_8__1004_;
  assign t_9__747_ = t_8__747_ | t_8__1003_;
  assign t_9__746_ = t_8__746_ | t_8__1002_;
  assign t_9__745_ = t_8__745_ | t_8__1001_;
  assign t_9__744_ = t_8__744_ | t_8__1000_;
  assign t_9__743_ = t_8__743_ | t_8__999_;
  assign t_9__742_ = t_8__742_ | t_8__998_;
  assign t_9__741_ = t_8__741_ | t_8__997_;
  assign t_9__740_ = t_8__740_ | t_8__996_;
  assign t_9__739_ = t_8__739_ | t_8__995_;
  assign t_9__738_ = t_8__738_ | t_8__994_;
  assign t_9__737_ = t_8__737_ | t_8__993_;
  assign t_9__736_ = t_8__736_ | t_8__992_;
  assign t_9__735_ = t_8__735_ | t_8__991_;
  assign t_9__734_ = t_8__734_ | t_8__990_;
  assign t_9__733_ = t_8__733_ | t_8__989_;
  assign t_9__732_ = t_8__732_ | t_8__988_;
  assign t_9__731_ = t_8__731_ | t_8__987_;
  assign t_9__730_ = t_8__730_ | t_8__986_;
  assign t_9__729_ = t_8__729_ | t_8__985_;
  assign t_9__728_ = t_8__728_ | t_8__984_;
  assign t_9__727_ = t_8__727_ | t_8__983_;
  assign t_9__726_ = t_8__726_ | t_8__982_;
  assign t_9__725_ = t_8__725_ | t_8__981_;
  assign t_9__724_ = t_8__724_ | t_8__980_;
  assign t_9__723_ = t_8__723_ | t_8__979_;
  assign t_9__722_ = t_8__722_ | t_8__978_;
  assign t_9__721_ = t_8__721_ | t_8__977_;
  assign t_9__720_ = t_8__720_ | t_8__976_;
  assign t_9__719_ = t_8__719_ | t_8__975_;
  assign t_9__718_ = t_8__718_ | t_8__974_;
  assign t_9__717_ = t_8__717_ | t_8__973_;
  assign t_9__716_ = t_8__716_ | t_8__972_;
  assign t_9__715_ = t_8__715_ | t_8__971_;
  assign t_9__714_ = t_8__714_ | t_8__970_;
  assign t_9__713_ = t_8__713_ | t_8__969_;
  assign t_9__712_ = t_8__712_ | t_8__968_;
  assign t_9__711_ = t_8__711_ | t_8__967_;
  assign t_9__710_ = t_8__710_ | t_8__966_;
  assign t_9__709_ = t_8__709_ | t_8__965_;
  assign t_9__708_ = t_8__708_ | t_8__964_;
  assign t_9__707_ = t_8__707_ | t_8__963_;
  assign t_9__706_ = t_8__706_ | t_8__962_;
  assign t_9__705_ = t_8__705_ | t_8__961_;
  assign t_9__704_ = t_8__704_ | t_8__960_;
  assign t_9__703_ = t_8__703_ | t_8__959_;
  assign t_9__702_ = t_8__702_ | t_8__958_;
  assign t_9__701_ = t_8__701_ | t_8__957_;
  assign t_9__700_ = t_8__700_ | t_8__956_;
  assign t_9__699_ = t_8__699_ | t_8__955_;
  assign t_9__698_ = t_8__698_ | t_8__954_;
  assign t_9__697_ = t_8__697_ | t_8__953_;
  assign t_9__696_ = t_8__696_ | t_8__952_;
  assign t_9__695_ = t_8__695_ | t_8__951_;
  assign t_9__694_ = t_8__694_ | t_8__950_;
  assign t_9__693_ = t_8__693_ | t_8__949_;
  assign t_9__692_ = t_8__692_ | t_8__948_;
  assign t_9__691_ = t_8__691_ | t_8__947_;
  assign t_9__690_ = t_8__690_ | t_8__946_;
  assign t_9__689_ = t_8__689_ | t_8__945_;
  assign t_9__688_ = t_8__688_ | t_8__944_;
  assign t_9__687_ = t_8__687_ | t_8__943_;
  assign t_9__686_ = t_8__686_ | t_8__942_;
  assign t_9__685_ = t_8__685_ | t_8__941_;
  assign t_9__684_ = t_8__684_ | t_8__940_;
  assign t_9__683_ = t_8__683_ | t_8__939_;
  assign t_9__682_ = t_8__682_ | t_8__938_;
  assign t_9__681_ = t_8__681_ | t_8__937_;
  assign t_9__680_ = t_8__680_ | t_8__936_;
  assign t_9__679_ = t_8__679_ | t_8__935_;
  assign t_9__678_ = t_8__678_ | t_8__934_;
  assign t_9__677_ = t_8__677_ | t_8__933_;
  assign t_9__676_ = t_8__676_ | t_8__932_;
  assign t_9__675_ = t_8__675_ | t_8__931_;
  assign t_9__674_ = t_8__674_ | t_8__930_;
  assign t_9__673_ = t_8__673_ | t_8__929_;
  assign t_9__672_ = t_8__672_ | t_8__928_;
  assign t_9__671_ = t_8__671_ | t_8__927_;
  assign t_9__670_ = t_8__670_ | t_8__926_;
  assign t_9__669_ = t_8__669_ | t_8__925_;
  assign t_9__668_ = t_8__668_ | t_8__924_;
  assign t_9__667_ = t_8__667_ | t_8__923_;
  assign t_9__666_ = t_8__666_ | t_8__922_;
  assign t_9__665_ = t_8__665_ | t_8__921_;
  assign t_9__664_ = t_8__664_ | t_8__920_;
  assign t_9__663_ = t_8__663_ | t_8__919_;
  assign t_9__662_ = t_8__662_ | t_8__918_;
  assign t_9__661_ = t_8__661_ | t_8__917_;
  assign t_9__660_ = t_8__660_ | t_8__916_;
  assign t_9__659_ = t_8__659_ | t_8__915_;
  assign t_9__658_ = t_8__658_ | t_8__914_;
  assign t_9__657_ = t_8__657_ | t_8__913_;
  assign t_9__656_ = t_8__656_ | t_8__912_;
  assign t_9__655_ = t_8__655_ | t_8__911_;
  assign t_9__654_ = t_8__654_ | t_8__910_;
  assign t_9__653_ = t_8__653_ | t_8__909_;
  assign t_9__652_ = t_8__652_ | t_8__908_;
  assign t_9__651_ = t_8__651_ | t_8__907_;
  assign t_9__650_ = t_8__650_ | t_8__906_;
  assign t_9__649_ = t_8__649_ | t_8__905_;
  assign t_9__648_ = t_8__648_ | t_8__904_;
  assign t_9__647_ = t_8__647_ | t_8__903_;
  assign t_9__646_ = t_8__646_ | t_8__902_;
  assign t_9__645_ = t_8__645_ | t_8__901_;
  assign t_9__644_ = t_8__644_ | t_8__900_;
  assign t_9__643_ = t_8__643_ | t_8__899_;
  assign t_9__642_ = t_8__642_ | t_8__898_;
  assign t_9__641_ = t_8__641_ | t_8__897_;
  assign t_9__640_ = t_8__640_ | t_8__896_;
  assign t_9__639_ = t_8__639_ | t_8__895_;
  assign t_9__638_ = t_8__638_ | t_8__894_;
  assign t_9__637_ = t_8__637_ | t_8__893_;
  assign t_9__636_ = t_8__636_ | t_8__892_;
  assign t_9__635_ = t_8__635_ | t_8__891_;
  assign t_9__634_ = t_8__634_ | t_8__890_;
  assign t_9__633_ = t_8__633_ | t_8__889_;
  assign t_9__632_ = t_8__632_ | t_8__888_;
  assign t_9__631_ = t_8__631_ | t_8__887_;
  assign t_9__630_ = t_8__630_ | t_8__886_;
  assign t_9__629_ = t_8__629_ | t_8__885_;
  assign t_9__628_ = t_8__628_ | t_8__884_;
  assign t_9__627_ = t_8__627_ | t_8__883_;
  assign t_9__626_ = t_8__626_ | t_8__882_;
  assign t_9__625_ = t_8__625_ | t_8__881_;
  assign t_9__624_ = t_8__624_ | t_8__880_;
  assign t_9__623_ = t_8__623_ | t_8__879_;
  assign t_9__622_ = t_8__622_ | t_8__878_;
  assign t_9__621_ = t_8__621_ | t_8__877_;
  assign t_9__620_ = t_8__620_ | t_8__876_;
  assign t_9__619_ = t_8__619_ | t_8__875_;
  assign t_9__618_ = t_8__618_ | t_8__874_;
  assign t_9__617_ = t_8__617_ | t_8__873_;
  assign t_9__616_ = t_8__616_ | t_8__872_;
  assign t_9__615_ = t_8__615_ | t_8__871_;
  assign t_9__614_ = t_8__614_ | t_8__870_;
  assign t_9__613_ = t_8__613_ | t_8__869_;
  assign t_9__612_ = t_8__612_ | t_8__868_;
  assign t_9__611_ = t_8__611_ | t_8__867_;
  assign t_9__610_ = t_8__610_ | t_8__866_;
  assign t_9__609_ = t_8__609_ | t_8__865_;
  assign t_9__608_ = t_8__608_ | t_8__864_;
  assign t_9__607_ = t_8__607_ | t_8__863_;
  assign t_9__606_ = t_8__606_ | t_8__862_;
  assign t_9__605_ = t_8__605_ | t_8__861_;
  assign t_9__604_ = t_8__604_ | t_8__860_;
  assign t_9__603_ = t_8__603_ | t_8__859_;
  assign t_9__602_ = t_8__602_ | t_8__858_;
  assign t_9__601_ = t_8__601_ | t_8__857_;
  assign t_9__600_ = t_8__600_ | t_8__856_;
  assign t_9__599_ = t_8__599_ | t_8__855_;
  assign t_9__598_ = t_8__598_ | t_8__854_;
  assign t_9__597_ = t_8__597_ | t_8__853_;
  assign t_9__596_ = t_8__596_ | t_8__852_;
  assign t_9__595_ = t_8__595_ | t_8__851_;
  assign t_9__594_ = t_8__594_ | t_8__850_;
  assign t_9__593_ = t_8__593_ | t_8__849_;
  assign t_9__592_ = t_8__592_ | t_8__848_;
  assign t_9__591_ = t_8__591_ | t_8__847_;
  assign t_9__590_ = t_8__590_ | t_8__846_;
  assign t_9__589_ = t_8__589_ | t_8__845_;
  assign t_9__588_ = t_8__588_ | t_8__844_;
  assign t_9__587_ = t_8__587_ | t_8__843_;
  assign t_9__586_ = t_8__586_ | t_8__842_;
  assign t_9__585_ = t_8__585_ | t_8__841_;
  assign t_9__584_ = t_8__584_ | t_8__840_;
  assign t_9__583_ = t_8__583_ | t_8__839_;
  assign t_9__582_ = t_8__582_ | t_8__838_;
  assign t_9__581_ = t_8__581_ | t_8__837_;
  assign t_9__580_ = t_8__580_ | t_8__836_;
  assign t_9__579_ = t_8__579_ | t_8__835_;
  assign t_9__578_ = t_8__578_ | t_8__834_;
  assign t_9__577_ = t_8__577_ | t_8__833_;
  assign t_9__576_ = t_8__576_ | t_8__832_;
  assign t_9__575_ = t_8__575_ | t_8__831_;
  assign t_9__574_ = t_8__574_ | t_8__830_;
  assign t_9__573_ = t_8__573_ | t_8__829_;
  assign t_9__572_ = t_8__572_ | t_8__828_;
  assign t_9__571_ = t_8__571_ | t_8__827_;
  assign t_9__570_ = t_8__570_ | t_8__826_;
  assign t_9__569_ = t_8__569_ | t_8__825_;
  assign t_9__568_ = t_8__568_ | t_8__824_;
  assign t_9__567_ = t_8__567_ | t_8__823_;
  assign t_9__566_ = t_8__566_ | t_8__822_;
  assign t_9__565_ = t_8__565_ | t_8__821_;
  assign t_9__564_ = t_8__564_ | t_8__820_;
  assign t_9__563_ = t_8__563_ | t_8__819_;
  assign t_9__562_ = t_8__562_ | t_8__818_;
  assign t_9__561_ = t_8__561_ | t_8__817_;
  assign t_9__560_ = t_8__560_ | t_8__816_;
  assign t_9__559_ = t_8__559_ | t_8__815_;
  assign t_9__558_ = t_8__558_ | t_8__814_;
  assign t_9__557_ = t_8__557_ | t_8__813_;
  assign t_9__556_ = t_8__556_ | t_8__812_;
  assign t_9__555_ = t_8__555_ | t_8__811_;
  assign t_9__554_ = t_8__554_ | t_8__810_;
  assign t_9__553_ = t_8__553_ | t_8__809_;
  assign t_9__552_ = t_8__552_ | t_8__808_;
  assign t_9__551_ = t_8__551_ | t_8__807_;
  assign t_9__550_ = t_8__550_ | t_8__806_;
  assign t_9__549_ = t_8__549_ | t_8__805_;
  assign t_9__548_ = t_8__548_ | t_8__804_;
  assign t_9__547_ = t_8__547_ | t_8__803_;
  assign t_9__546_ = t_8__546_ | t_8__802_;
  assign t_9__545_ = t_8__545_ | t_8__801_;
  assign t_9__544_ = t_8__544_ | t_8__800_;
  assign t_9__543_ = t_8__543_ | t_8__799_;
  assign t_9__542_ = t_8__542_ | t_8__798_;
  assign t_9__541_ = t_8__541_ | t_8__797_;
  assign t_9__540_ = t_8__540_ | t_8__796_;
  assign t_9__539_ = t_8__539_ | t_8__795_;
  assign t_9__538_ = t_8__538_ | t_8__794_;
  assign t_9__537_ = t_8__537_ | t_8__793_;
  assign t_9__536_ = t_8__536_ | t_8__792_;
  assign t_9__535_ = t_8__535_ | t_8__791_;
  assign t_9__534_ = t_8__534_ | t_8__790_;
  assign t_9__533_ = t_8__533_ | t_8__789_;
  assign t_9__532_ = t_8__532_ | t_8__788_;
  assign t_9__531_ = t_8__531_ | t_8__787_;
  assign t_9__530_ = t_8__530_ | t_8__786_;
  assign t_9__529_ = t_8__529_ | t_8__785_;
  assign t_9__528_ = t_8__528_ | t_8__784_;
  assign t_9__527_ = t_8__527_ | t_8__783_;
  assign t_9__526_ = t_8__526_ | t_8__782_;
  assign t_9__525_ = t_8__525_ | t_8__781_;
  assign t_9__524_ = t_8__524_ | t_8__780_;
  assign t_9__523_ = t_8__523_ | t_8__779_;
  assign t_9__522_ = t_8__522_ | t_8__778_;
  assign t_9__521_ = t_8__521_ | t_8__777_;
  assign t_9__520_ = t_8__520_ | t_8__776_;
  assign t_9__519_ = t_8__519_ | t_8__775_;
  assign t_9__518_ = t_8__518_ | t_8__774_;
  assign t_9__517_ = t_8__517_ | t_8__773_;
  assign t_9__516_ = t_8__516_ | t_8__772_;
  assign t_9__515_ = t_8__515_ | t_8__771_;
  assign t_9__514_ = t_8__514_ | t_8__770_;
  assign t_9__513_ = t_8__513_ | t_8__769_;
  assign t_9__512_ = t_8__512_ | t_8__768_;
  assign t_9__511_ = t_8__511_ | t_8__767_;
  assign t_9__510_ = t_8__510_ | t_8__766_;
  assign t_9__509_ = t_8__509_ | t_8__765_;
  assign t_9__508_ = t_8__508_ | t_8__764_;
  assign t_9__507_ = t_8__507_ | t_8__763_;
  assign t_9__506_ = t_8__506_ | t_8__762_;
  assign t_9__505_ = t_8__505_ | t_8__761_;
  assign t_9__504_ = t_8__504_ | t_8__760_;
  assign t_9__503_ = t_8__503_ | t_8__759_;
  assign t_9__502_ = t_8__502_ | t_8__758_;
  assign t_9__501_ = t_8__501_ | t_8__757_;
  assign t_9__500_ = t_8__500_ | t_8__756_;
  assign t_9__499_ = t_8__499_ | t_8__755_;
  assign t_9__498_ = t_8__498_ | t_8__754_;
  assign t_9__497_ = t_8__497_ | t_8__753_;
  assign t_9__496_ = t_8__496_ | t_8__752_;
  assign t_9__495_ = t_8__495_ | t_8__751_;
  assign t_9__494_ = t_8__494_ | t_8__750_;
  assign t_9__493_ = t_8__493_ | t_8__749_;
  assign t_9__492_ = t_8__492_ | t_8__748_;
  assign t_9__491_ = t_8__491_ | t_8__747_;
  assign t_9__490_ = t_8__490_ | t_8__746_;
  assign t_9__489_ = t_8__489_ | t_8__745_;
  assign t_9__488_ = t_8__488_ | t_8__744_;
  assign t_9__487_ = t_8__487_ | t_8__743_;
  assign t_9__486_ = t_8__486_ | t_8__742_;
  assign t_9__485_ = t_8__485_ | t_8__741_;
  assign t_9__484_ = t_8__484_ | t_8__740_;
  assign t_9__483_ = t_8__483_ | t_8__739_;
  assign t_9__482_ = t_8__482_ | t_8__738_;
  assign t_9__481_ = t_8__481_ | t_8__737_;
  assign t_9__480_ = t_8__480_ | t_8__736_;
  assign t_9__479_ = t_8__479_ | t_8__735_;
  assign t_9__478_ = t_8__478_ | t_8__734_;
  assign t_9__477_ = t_8__477_ | t_8__733_;
  assign t_9__476_ = t_8__476_ | t_8__732_;
  assign t_9__475_ = t_8__475_ | t_8__731_;
  assign t_9__474_ = t_8__474_ | t_8__730_;
  assign t_9__473_ = t_8__473_ | t_8__729_;
  assign t_9__472_ = t_8__472_ | t_8__728_;
  assign t_9__471_ = t_8__471_ | t_8__727_;
  assign t_9__470_ = t_8__470_ | t_8__726_;
  assign t_9__469_ = t_8__469_ | t_8__725_;
  assign t_9__468_ = t_8__468_ | t_8__724_;
  assign t_9__467_ = t_8__467_ | t_8__723_;
  assign t_9__466_ = t_8__466_ | t_8__722_;
  assign t_9__465_ = t_8__465_ | t_8__721_;
  assign t_9__464_ = t_8__464_ | t_8__720_;
  assign t_9__463_ = t_8__463_ | t_8__719_;
  assign t_9__462_ = t_8__462_ | t_8__718_;
  assign t_9__461_ = t_8__461_ | t_8__717_;
  assign t_9__460_ = t_8__460_ | t_8__716_;
  assign t_9__459_ = t_8__459_ | t_8__715_;
  assign t_9__458_ = t_8__458_ | t_8__714_;
  assign t_9__457_ = t_8__457_ | t_8__713_;
  assign t_9__456_ = t_8__456_ | t_8__712_;
  assign t_9__455_ = t_8__455_ | t_8__711_;
  assign t_9__454_ = t_8__454_ | t_8__710_;
  assign t_9__453_ = t_8__453_ | t_8__709_;
  assign t_9__452_ = t_8__452_ | t_8__708_;
  assign t_9__451_ = t_8__451_ | t_8__707_;
  assign t_9__450_ = t_8__450_ | t_8__706_;
  assign t_9__449_ = t_8__449_ | t_8__705_;
  assign t_9__448_ = t_8__448_ | t_8__704_;
  assign t_9__447_ = t_8__447_ | t_8__703_;
  assign t_9__446_ = t_8__446_ | t_8__702_;
  assign t_9__445_ = t_8__445_ | t_8__701_;
  assign t_9__444_ = t_8__444_ | t_8__700_;
  assign t_9__443_ = t_8__443_ | t_8__699_;
  assign t_9__442_ = t_8__442_ | t_8__698_;
  assign t_9__441_ = t_8__441_ | t_8__697_;
  assign t_9__440_ = t_8__440_ | t_8__696_;
  assign t_9__439_ = t_8__439_ | t_8__695_;
  assign t_9__438_ = t_8__438_ | t_8__694_;
  assign t_9__437_ = t_8__437_ | t_8__693_;
  assign t_9__436_ = t_8__436_ | t_8__692_;
  assign t_9__435_ = t_8__435_ | t_8__691_;
  assign t_9__434_ = t_8__434_ | t_8__690_;
  assign t_9__433_ = t_8__433_ | t_8__689_;
  assign t_9__432_ = t_8__432_ | t_8__688_;
  assign t_9__431_ = t_8__431_ | t_8__687_;
  assign t_9__430_ = t_8__430_ | t_8__686_;
  assign t_9__429_ = t_8__429_ | t_8__685_;
  assign t_9__428_ = t_8__428_ | t_8__684_;
  assign t_9__427_ = t_8__427_ | t_8__683_;
  assign t_9__426_ = t_8__426_ | t_8__682_;
  assign t_9__425_ = t_8__425_ | t_8__681_;
  assign t_9__424_ = t_8__424_ | t_8__680_;
  assign t_9__423_ = t_8__423_ | t_8__679_;
  assign t_9__422_ = t_8__422_ | t_8__678_;
  assign t_9__421_ = t_8__421_ | t_8__677_;
  assign t_9__420_ = t_8__420_ | t_8__676_;
  assign t_9__419_ = t_8__419_ | t_8__675_;
  assign t_9__418_ = t_8__418_ | t_8__674_;
  assign t_9__417_ = t_8__417_ | t_8__673_;
  assign t_9__416_ = t_8__416_ | t_8__672_;
  assign t_9__415_ = t_8__415_ | t_8__671_;
  assign t_9__414_ = t_8__414_ | t_8__670_;
  assign t_9__413_ = t_8__413_ | t_8__669_;
  assign t_9__412_ = t_8__412_ | t_8__668_;
  assign t_9__411_ = t_8__411_ | t_8__667_;
  assign t_9__410_ = t_8__410_ | t_8__666_;
  assign t_9__409_ = t_8__409_ | t_8__665_;
  assign t_9__408_ = t_8__408_ | t_8__664_;
  assign t_9__407_ = t_8__407_ | t_8__663_;
  assign t_9__406_ = t_8__406_ | t_8__662_;
  assign t_9__405_ = t_8__405_ | t_8__661_;
  assign t_9__404_ = t_8__404_ | t_8__660_;
  assign t_9__403_ = t_8__403_ | t_8__659_;
  assign t_9__402_ = t_8__402_ | t_8__658_;
  assign t_9__401_ = t_8__401_ | t_8__657_;
  assign t_9__400_ = t_8__400_ | t_8__656_;
  assign t_9__399_ = t_8__399_ | t_8__655_;
  assign t_9__398_ = t_8__398_ | t_8__654_;
  assign t_9__397_ = t_8__397_ | t_8__653_;
  assign t_9__396_ = t_8__396_ | t_8__652_;
  assign t_9__395_ = t_8__395_ | t_8__651_;
  assign t_9__394_ = t_8__394_ | t_8__650_;
  assign t_9__393_ = t_8__393_ | t_8__649_;
  assign t_9__392_ = t_8__392_ | t_8__648_;
  assign t_9__391_ = t_8__391_ | t_8__647_;
  assign t_9__390_ = t_8__390_ | t_8__646_;
  assign t_9__389_ = t_8__389_ | t_8__645_;
  assign t_9__388_ = t_8__388_ | t_8__644_;
  assign t_9__387_ = t_8__387_ | t_8__643_;
  assign t_9__386_ = t_8__386_ | t_8__642_;
  assign t_9__385_ = t_8__385_ | t_8__641_;
  assign t_9__384_ = t_8__384_ | t_8__640_;
  assign t_9__383_ = t_8__383_ | t_8__639_;
  assign t_9__382_ = t_8__382_ | t_8__638_;
  assign t_9__381_ = t_8__381_ | t_8__637_;
  assign t_9__380_ = t_8__380_ | t_8__636_;
  assign t_9__379_ = t_8__379_ | t_8__635_;
  assign t_9__378_ = t_8__378_ | t_8__634_;
  assign t_9__377_ = t_8__377_ | t_8__633_;
  assign t_9__376_ = t_8__376_ | t_8__632_;
  assign t_9__375_ = t_8__375_ | t_8__631_;
  assign t_9__374_ = t_8__374_ | t_8__630_;
  assign t_9__373_ = t_8__373_ | t_8__629_;
  assign t_9__372_ = t_8__372_ | t_8__628_;
  assign t_9__371_ = t_8__371_ | t_8__627_;
  assign t_9__370_ = t_8__370_ | t_8__626_;
  assign t_9__369_ = t_8__369_ | t_8__625_;
  assign t_9__368_ = t_8__368_ | t_8__624_;
  assign t_9__367_ = t_8__367_ | t_8__623_;
  assign t_9__366_ = t_8__366_ | t_8__622_;
  assign t_9__365_ = t_8__365_ | t_8__621_;
  assign t_9__364_ = t_8__364_ | t_8__620_;
  assign t_9__363_ = t_8__363_ | t_8__619_;
  assign t_9__362_ = t_8__362_ | t_8__618_;
  assign t_9__361_ = t_8__361_ | t_8__617_;
  assign t_9__360_ = t_8__360_ | t_8__616_;
  assign t_9__359_ = t_8__359_ | t_8__615_;
  assign t_9__358_ = t_8__358_ | t_8__614_;
  assign t_9__357_ = t_8__357_ | t_8__613_;
  assign t_9__356_ = t_8__356_ | t_8__612_;
  assign t_9__355_ = t_8__355_ | t_8__611_;
  assign t_9__354_ = t_8__354_ | t_8__610_;
  assign t_9__353_ = t_8__353_ | t_8__609_;
  assign t_9__352_ = t_8__352_ | t_8__608_;
  assign t_9__351_ = t_8__351_ | t_8__607_;
  assign t_9__350_ = t_8__350_ | t_8__606_;
  assign t_9__349_ = t_8__349_ | t_8__605_;
  assign t_9__348_ = t_8__348_ | t_8__604_;
  assign t_9__347_ = t_8__347_ | t_8__603_;
  assign t_9__346_ = t_8__346_ | t_8__602_;
  assign t_9__345_ = t_8__345_ | t_8__601_;
  assign t_9__344_ = t_8__344_ | t_8__600_;
  assign t_9__343_ = t_8__343_ | t_8__599_;
  assign t_9__342_ = t_8__342_ | t_8__598_;
  assign t_9__341_ = t_8__341_ | t_8__597_;
  assign t_9__340_ = t_8__340_ | t_8__596_;
  assign t_9__339_ = t_8__339_ | t_8__595_;
  assign t_9__338_ = t_8__338_ | t_8__594_;
  assign t_9__337_ = t_8__337_ | t_8__593_;
  assign t_9__336_ = t_8__336_ | t_8__592_;
  assign t_9__335_ = t_8__335_ | t_8__591_;
  assign t_9__334_ = t_8__334_ | t_8__590_;
  assign t_9__333_ = t_8__333_ | t_8__589_;
  assign t_9__332_ = t_8__332_ | t_8__588_;
  assign t_9__331_ = t_8__331_ | t_8__587_;
  assign t_9__330_ = t_8__330_ | t_8__586_;
  assign t_9__329_ = t_8__329_ | t_8__585_;
  assign t_9__328_ = t_8__328_ | t_8__584_;
  assign t_9__327_ = t_8__327_ | t_8__583_;
  assign t_9__326_ = t_8__326_ | t_8__582_;
  assign t_9__325_ = t_8__325_ | t_8__581_;
  assign t_9__324_ = t_8__324_ | t_8__580_;
  assign t_9__323_ = t_8__323_ | t_8__579_;
  assign t_9__322_ = t_8__322_ | t_8__578_;
  assign t_9__321_ = t_8__321_ | t_8__577_;
  assign t_9__320_ = t_8__320_ | t_8__576_;
  assign t_9__319_ = t_8__319_ | t_8__575_;
  assign t_9__318_ = t_8__318_ | t_8__574_;
  assign t_9__317_ = t_8__317_ | t_8__573_;
  assign t_9__316_ = t_8__316_ | t_8__572_;
  assign t_9__315_ = t_8__315_ | t_8__571_;
  assign t_9__314_ = t_8__314_ | t_8__570_;
  assign t_9__313_ = t_8__313_ | t_8__569_;
  assign t_9__312_ = t_8__312_ | t_8__568_;
  assign t_9__311_ = t_8__311_ | t_8__567_;
  assign t_9__310_ = t_8__310_ | t_8__566_;
  assign t_9__309_ = t_8__309_ | t_8__565_;
  assign t_9__308_ = t_8__308_ | t_8__564_;
  assign t_9__307_ = t_8__307_ | t_8__563_;
  assign t_9__306_ = t_8__306_ | t_8__562_;
  assign t_9__305_ = t_8__305_ | t_8__561_;
  assign t_9__304_ = t_8__304_ | t_8__560_;
  assign t_9__303_ = t_8__303_ | t_8__559_;
  assign t_9__302_ = t_8__302_ | t_8__558_;
  assign t_9__301_ = t_8__301_ | t_8__557_;
  assign t_9__300_ = t_8__300_ | t_8__556_;
  assign t_9__299_ = t_8__299_ | t_8__555_;
  assign t_9__298_ = t_8__298_ | t_8__554_;
  assign t_9__297_ = t_8__297_ | t_8__553_;
  assign t_9__296_ = t_8__296_ | t_8__552_;
  assign t_9__295_ = t_8__295_ | t_8__551_;
  assign t_9__294_ = t_8__294_ | t_8__550_;
  assign t_9__293_ = t_8__293_ | t_8__549_;
  assign t_9__292_ = t_8__292_ | t_8__548_;
  assign t_9__291_ = t_8__291_ | t_8__547_;
  assign t_9__290_ = t_8__290_ | t_8__546_;
  assign t_9__289_ = t_8__289_ | t_8__545_;
  assign t_9__288_ = t_8__288_ | t_8__544_;
  assign t_9__287_ = t_8__287_ | t_8__543_;
  assign t_9__286_ = t_8__286_ | t_8__542_;
  assign t_9__285_ = t_8__285_ | t_8__541_;
  assign t_9__284_ = t_8__284_ | t_8__540_;
  assign t_9__283_ = t_8__283_ | t_8__539_;
  assign t_9__282_ = t_8__282_ | t_8__538_;
  assign t_9__281_ = t_8__281_ | t_8__537_;
  assign t_9__280_ = t_8__280_ | t_8__536_;
  assign t_9__279_ = t_8__279_ | t_8__535_;
  assign t_9__278_ = t_8__278_ | t_8__534_;
  assign t_9__277_ = t_8__277_ | t_8__533_;
  assign t_9__276_ = t_8__276_ | t_8__532_;
  assign t_9__275_ = t_8__275_ | t_8__531_;
  assign t_9__274_ = t_8__274_ | t_8__530_;
  assign t_9__273_ = t_8__273_ | t_8__529_;
  assign t_9__272_ = t_8__272_ | t_8__528_;
  assign t_9__271_ = t_8__271_ | t_8__527_;
  assign t_9__270_ = t_8__270_ | t_8__526_;
  assign t_9__269_ = t_8__269_ | t_8__525_;
  assign t_9__268_ = t_8__268_ | t_8__524_;
  assign t_9__267_ = t_8__267_ | t_8__523_;
  assign t_9__266_ = t_8__266_ | t_8__522_;
  assign t_9__265_ = t_8__265_ | t_8__521_;
  assign t_9__264_ = t_8__264_ | t_8__520_;
  assign t_9__263_ = t_8__263_ | t_8__519_;
  assign t_9__262_ = t_8__262_ | t_8__518_;
  assign t_9__261_ = t_8__261_ | t_8__517_;
  assign t_9__260_ = t_8__260_ | t_8__516_;
  assign t_9__259_ = t_8__259_ | t_8__515_;
  assign t_9__258_ = t_8__258_ | t_8__514_;
  assign t_9__257_ = t_8__257_ | t_8__513_;
  assign t_9__256_ = t_8__256_ | t_8__512_;
  assign t_9__255_ = t_8__255_ | t_8__511_;
  assign t_9__254_ = t_8__254_ | t_8__510_;
  assign t_9__253_ = t_8__253_ | t_8__509_;
  assign t_9__252_ = t_8__252_ | t_8__508_;
  assign t_9__251_ = t_8__251_ | t_8__507_;
  assign t_9__250_ = t_8__250_ | t_8__506_;
  assign t_9__249_ = t_8__249_ | t_8__505_;
  assign t_9__248_ = t_8__248_ | t_8__504_;
  assign t_9__247_ = t_8__247_ | t_8__503_;
  assign t_9__246_ = t_8__246_ | t_8__502_;
  assign t_9__245_ = t_8__245_ | t_8__501_;
  assign t_9__244_ = t_8__244_ | t_8__500_;
  assign t_9__243_ = t_8__243_ | t_8__499_;
  assign t_9__242_ = t_8__242_ | t_8__498_;
  assign t_9__241_ = t_8__241_ | t_8__497_;
  assign t_9__240_ = t_8__240_ | t_8__496_;
  assign t_9__239_ = t_8__239_ | t_8__495_;
  assign t_9__238_ = t_8__238_ | t_8__494_;
  assign t_9__237_ = t_8__237_ | t_8__493_;
  assign t_9__236_ = t_8__236_ | t_8__492_;
  assign t_9__235_ = t_8__235_ | t_8__491_;
  assign t_9__234_ = t_8__234_ | t_8__490_;
  assign t_9__233_ = t_8__233_ | t_8__489_;
  assign t_9__232_ = t_8__232_ | t_8__488_;
  assign t_9__231_ = t_8__231_ | t_8__487_;
  assign t_9__230_ = t_8__230_ | t_8__486_;
  assign t_9__229_ = t_8__229_ | t_8__485_;
  assign t_9__228_ = t_8__228_ | t_8__484_;
  assign t_9__227_ = t_8__227_ | t_8__483_;
  assign t_9__226_ = t_8__226_ | t_8__482_;
  assign t_9__225_ = t_8__225_ | t_8__481_;
  assign t_9__224_ = t_8__224_ | t_8__480_;
  assign t_9__223_ = t_8__223_ | t_8__479_;
  assign t_9__222_ = t_8__222_ | t_8__478_;
  assign t_9__221_ = t_8__221_ | t_8__477_;
  assign t_9__220_ = t_8__220_ | t_8__476_;
  assign t_9__219_ = t_8__219_ | t_8__475_;
  assign t_9__218_ = t_8__218_ | t_8__474_;
  assign t_9__217_ = t_8__217_ | t_8__473_;
  assign t_9__216_ = t_8__216_ | t_8__472_;
  assign t_9__215_ = t_8__215_ | t_8__471_;
  assign t_9__214_ = t_8__214_ | t_8__470_;
  assign t_9__213_ = t_8__213_ | t_8__469_;
  assign t_9__212_ = t_8__212_ | t_8__468_;
  assign t_9__211_ = t_8__211_ | t_8__467_;
  assign t_9__210_ = t_8__210_ | t_8__466_;
  assign t_9__209_ = t_8__209_ | t_8__465_;
  assign t_9__208_ = t_8__208_ | t_8__464_;
  assign t_9__207_ = t_8__207_ | t_8__463_;
  assign t_9__206_ = t_8__206_ | t_8__462_;
  assign t_9__205_ = t_8__205_ | t_8__461_;
  assign t_9__204_ = t_8__204_ | t_8__460_;
  assign t_9__203_ = t_8__203_ | t_8__459_;
  assign t_9__202_ = t_8__202_ | t_8__458_;
  assign t_9__201_ = t_8__201_ | t_8__457_;
  assign t_9__200_ = t_8__200_ | t_8__456_;
  assign t_9__199_ = t_8__199_ | t_8__455_;
  assign t_9__198_ = t_8__198_ | t_8__454_;
  assign t_9__197_ = t_8__197_ | t_8__453_;
  assign t_9__196_ = t_8__196_ | t_8__452_;
  assign t_9__195_ = t_8__195_ | t_8__451_;
  assign t_9__194_ = t_8__194_ | t_8__450_;
  assign t_9__193_ = t_8__193_ | t_8__449_;
  assign t_9__192_ = t_8__192_ | t_8__448_;
  assign t_9__191_ = t_8__191_ | t_8__447_;
  assign t_9__190_ = t_8__190_ | t_8__446_;
  assign t_9__189_ = t_8__189_ | t_8__445_;
  assign t_9__188_ = t_8__188_ | t_8__444_;
  assign t_9__187_ = t_8__187_ | t_8__443_;
  assign t_9__186_ = t_8__186_ | t_8__442_;
  assign t_9__185_ = t_8__185_ | t_8__441_;
  assign t_9__184_ = t_8__184_ | t_8__440_;
  assign t_9__183_ = t_8__183_ | t_8__439_;
  assign t_9__182_ = t_8__182_ | t_8__438_;
  assign t_9__181_ = t_8__181_ | t_8__437_;
  assign t_9__180_ = t_8__180_ | t_8__436_;
  assign t_9__179_ = t_8__179_ | t_8__435_;
  assign t_9__178_ = t_8__178_ | t_8__434_;
  assign t_9__177_ = t_8__177_ | t_8__433_;
  assign t_9__176_ = t_8__176_ | t_8__432_;
  assign t_9__175_ = t_8__175_ | t_8__431_;
  assign t_9__174_ = t_8__174_ | t_8__430_;
  assign t_9__173_ = t_8__173_ | t_8__429_;
  assign t_9__172_ = t_8__172_ | t_8__428_;
  assign t_9__171_ = t_8__171_ | t_8__427_;
  assign t_9__170_ = t_8__170_ | t_8__426_;
  assign t_9__169_ = t_8__169_ | t_8__425_;
  assign t_9__168_ = t_8__168_ | t_8__424_;
  assign t_9__167_ = t_8__167_ | t_8__423_;
  assign t_9__166_ = t_8__166_ | t_8__422_;
  assign t_9__165_ = t_8__165_ | t_8__421_;
  assign t_9__164_ = t_8__164_ | t_8__420_;
  assign t_9__163_ = t_8__163_ | t_8__419_;
  assign t_9__162_ = t_8__162_ | t_8__418_;
  assign t_9__161_ = t_8__161_ | t_8__417_;
  assign t_9__160_ = t_8__160_ | t_8__416_;
  assign t_9__159_ = t_8__159_ | t_8__415_;
  assign t_9__158_ = t_8__158_ | t_8__414_;
  assign t_9__157_ = t_8__157_ | t_8__413_;
  assign t_9__156_ = t_8__156_ | t_8__412_;
  assign t_9__155_ = t_8__155_ | t_8__411_;
  assign t_9__154_ = t_8__154_ | t_8__410_;
  assign t_9__153_ = t_8__153_ | t_8__409_;
  assign t_9__152_ = t_8__152_ | t_8__408_;
  assign t_9__151_ = t_8__151_ | t_8__407_;
  assign t_9__150_ = t_8__150_ | t_8__406_;
  assign t_9__149_ = t_8__149_ | t_8__405_;
  assign t_9__148_ = t_8__148_ | t_8__404_;
  assign t_9__147_ = t_8__147_ | t_8__403_;
  assign t_9__146_ = t_8__146_ | t_8__402_;
  assign t_9__145_ = t_8__145_ | t_8__401_;
  assign t_9__144_ = t_8__144_ | t_8__400_;
  assign t_9__143_ = t_8__143_ | t_8__399_;
  assign t_9__142_ = t_8__142_ | t_8__398_;
  assign t_9__141_ = t_8__141_ | t_8__397_;
  assign t_9__140_ = t_8__140_ | t_8__396_;
  assign t_9__139_ = t_8__139_ | t_8__395_;
  assign t_9__138_ = t_8__138_ | t_8__394_;
  assign t_9__137_ = t_8__137_ | t_8__393_;
  assign t_9__136_ = t_8__136_ | t_8__392_;
  assign t_9__135_ = t_8__135_ | t_8__391_;
  assign t_9__134_ = t_8__134_ | t_8__390_;
  assign t_9__133_ = t_8__133_ | t_8__389_;
  assign t_9__132_ = t_8__132_ | t_8__388_;
  assign t_9__131_ = t_8__131_ | t_8__387_;
  assign t_9__130_ = t_8__130_ | t_8__386_;
  assign t_9__129_ = t_8__129_ | t_8__385_;
  assign t_9__128_ = t_8__128_ | t_8__384_;
  assign t_9__127_ = t_8__127_ | t_8__383_;
  assign t_9__126_ = t_8__126_ | t_8__382_;
  assign t_9__125_ = t_8__125_ | t_8__381_;
  assign t_9__124_ = t_8__124_ | t_8__380_;
  assign t_9__123_ = t_8__123_ | t_8__379_;
  assign t_9__122_ = t_8__122_ | t_8__378_;
  assign t_9__121_ = t_8__121_ | t_8__377_;
  assign t_9__120_ = t_8__120_ | t_8__376_;
  assign t_9__119_ = t_8__119_ | t_8__375_;
  assign t_9__118_ = t_8__118_ | t_8__374_;
  assign t_9__117_ = t_8__117_ | t_8__373_;
  assign t_9__116_ = t_8__116_ | t_8__372_;
  assign t_9__115_ = t_8__115_ | t_8__371_;
  assign t_9__114_ = t_8__114_ | t_8__370_;
  assign t_9__113_ = t_8__113_ | t_8__369_;
  assign t_9__112_ = t_8__112_ | t_8__368_;
  assign t_9__111_ = t_8__111_ | t_8__367_;
  assign t_9__110_ = t_8__110_ | t_8__366_;
  assign t_9__109_ = t_8__109_ | t_8__365_;
  assign t_9__108_ = t_8__108_ | t_8__364_;
  assign t_9__107_ = t_8__107_ | t_8__363_;
  assign t_9__106_ = t_8__106_ | t_8__362_;
  assign t_9__105_ = t_8__105_ | t_8__361_;
  assign t_9__104_ = t_8__104_ | t_8__360_;
  assign t_9__103_ = t_8__103_ | t_8__359_;
  assign t_9__102_ = t_8__102_ | t_8__358_;
  assign t_9__101_ = t_8__101_ | t_8__357_;
  assign t_9__100_ = t_8__100_ | t_8__356_;
  assign t_9__99_ = t_8__99_ | t_8__355_;
  assign t_9__98_ = t_8__98_ | t_8__354_;
  assign t_9__97_ = t_8__97_ | t_8__353_;
  assign t_9__96_ = t_8__96_ | t_8__352_;
  assign t_9__95_ = t_8__95_ | t_8__351_;
  assign t_9__94_ = t_8__94_ | t_8__350_;
  assign t_9__93_ = t_8__93_ | t_8__349_;
  assign t_9__92_ = t_8__92_ | t_8__348_;
  assign t_9__91_ = t_8__91_ | t_8__347_;
  assign t_9__90_ = t_8__90_ | t_8__346_;
  assign t_9__89_ = t_8__89_ | t_8__345_;
  assign t_9__88_ = t_8__88_ | t_8__344_;
  assign t_9__87_ = t_8__87_ | t_8__343_;
  assign t_9__86_ = t_8__86_ | t_8__342_;
  assign t_9__85_ = t_8__85_ | t_8__341_;
  assign t_9__84_ = t_8__84_ | t_8__340_;
  assign t_9__83_ = t_8__83_ | t_8__339_;
  assign t_9__82_ = t_8__82_ | t_8__338_;
  assign t_9__81_ = t_8__81_ | t_8__337_;
  assign t_9__80_ = t_8__80_ | t_8__336_;
  assign t_9__79_ = t_8__79_ | t_8__335_;
  assign t_9__78_ = t_8__78_ | t_8__334_;
  assign t_9__77_ = t_8__77_ | t_8__333_;
  assign t_9__76_ = t_8__76_ | t_8__332_;
  assign t_9__75_ = t_8__75_ | t_8__331_;
  assign t_9__74_ = t_8__74_ | t_8__330_;
  assign t_9__73_ = t_8__73_ | t_8__329_;
  assign t_9__72_ = t_8__72_ | t_8__328_;
  assign t_9__71_ = t_8__71_ | t_8__327_;
  assign t_9__70_ = t_8__70_ | t_8__326_;
  assign t_9__69_ = t_8__69_ | t_8__325_;
  assign t_9__68_ = t_8__68_ | t_8__324_;
  assign t_9__67_ = t_8__67_ | t_8__323_;
  assign t_9__66_ = t_8__66_ | t_8__322_;
  assign t_9__65_ = t_8__65_ | t_8__321_;
  assign t_9__64_ = t_8__64_ | t_8__320_;
  assign t_9__63_ = t_8__63_ | t_8__319_;
  assign t_9__62_ = t_8__62_ | t_8__318_;
  assign t_9__61_ = t_8__61_ | t_8__317_;
  assign t_9__60_ = t_8__60_ | t_8__316_;
  assign t_9__59_ = t_8__59_ | t_8__315_;
  assign t_9__58_ = t_8__58_ | t_8__314_;
  assign t_9__57_ = t_8__57_ | t_8__313_;
  assign t_9__56_ = t_8__56_ | t_8__312_;
  assign t_9__55_ = t_8__55_ | t_8__311_;
  assign t_9__54_ = t_8__54_ | t_8__310_;
  assign t_9__53_ = t_8__53_ | t_8__309_;
  assign t_9__52_ = t_8__52_ | t_8__308_;
  assign t_9__51_ = t_8__51_ | t_8__307_;
  assign t_9__50_ = t_8__50_ | t_8__306_;
  assign t_9__49_ = t_8__49_ | t_8__305_;
  assign t_9__48_ = t_8__48_ | t_8__304_;
  assign t_9__47_ = t_8__47_ | t_8__303_;
  assign t_9__46_ = t_8__46_ | t_8__302_;
  assign t_9__45_ = t_8__45_ | t_8__301_;
  assign t_9__44_ = t_8__44_ | t_8__300_;
  assign t_9__43_ = t_8__43_ | t_8__299_;
  assign t_9__42_ = t_8__42_ | t_8__298_;
  assign t_9__41_ = t_8__41_ | t_8__297_;
  assign t_9__40_ = t_8__40_ | t_8__296_;
  assign t_9__39_ = t_8__39_ | t_8__295_;
  assign t_9__38_ = t_8__38_ | t_8__294_;
  assign t_9__37_ = t_8__37_ | t_8__293_;
  assign t_9__36_ = t_8__36_ | t_8__292_;
  assign t_9__35_ = t_8__35_ | t_8__291_;
  assign t_9__34_ = t_8__34_ | t_8__290_;
  assign t_9__33_ = t_8__33_ | t_8__289_;
  assign t_9__32_ = t_8__32_ | t_8__288_;
  assign t_9__31_ = t_8__31_ | t_8__287_;
  assign t_9__30_ = t_8__30_ | t_8__286_;
  assign t_9__29_ = t_8__29_ | t_8__285_;
  assign t_9__28_ = t_8__28_ | t_8__284_;
  assign t_9__27_ = t_8__27_ | t_8__283_;
  assign t_9__26_ = t_8__26_ | t_8__282_;
  assign t_9__25_ = t_8__25_ | t_8__281_;
  assign t_9__24_ = t_8__24_ | t_8__280_;
  assign t_9__23_ = t_8__23_ | t_8__279_;
  assign t_9__22_ = t_8__22_ | t_8__278_;
  assign t_9__21_ = t_8__21_ | t_8__277_;
  assign t_9__20_ = t_8__20_ | t_8__276_;
  assign t_9__19_ = t_8__19_ | t_8__275_;
  assign t_9__18_ = t_8__18_ | t_8__274_;
  assign t_9__17_ = t_8__17_ | t_8__273_;
  assign t_9__16_ = t_8__16_ | t_8__272_;
  assign t_9__15_ = t_8__15_ | t_8__271_;
  assign t_9__14_ = t_8__14_ | t_8__270_;
  assign t_9__13_ = t_8__13_ | t_8__269_;
  assign t_9__12_ = t_8__12_ | t_8__268_;
  assign t_9__11_ = t_8__11_ | t_8__267_;
  assign t_9__10_ = t_8__10_ | t_8__266_;
  assign t_9__9_ = t_8__9_ | t_8__265_;
  assign t_9__8_ = t_8__8_ | t_8__264_;
  assign t_9__7_ = t_8__7_ | t_8__263_;
  assign t_9__6_ = t_8__6_ | t_8__262_;
  assign t_9__5_ = t_8__5_ | t_8__261_;
  assign t_9__4_ = t_8__4_ | t_8__260_;
  assign t_9__3_ = t_8__3_ | t_8__259_;
  assign t_9__2_ = t_8__2_ | t_8__258_;
  assign t_9__1_ = t_8__1_ | t_8__257_;
  assign t_9__0_ = t_8__0_ | t_8__256_;
  assign o[0] = t_9__1023_ | 1'b0;
  assign o[1] = t_9__1022_ | 1'b0;
  assign o[2] = t_9__1021_ | 1'b0;
  assign o[3] = t_9__1020_ | 1'b0;
  assign o[4] = t_9__1019_ | 1'b0;
  assign o[5] = t_9__1018_ | 1'b0;
  assign o[6] = t_9__1017_ | 1'b0;
  assign o[7] = t_9__1016_ | 1'b0;
  assign o[8] = t_9__1015_ | 1'b0;
  assign o[9] = t_9__1014_ | 1'b0;
  assign o[10] = t_9__1013_ | 1'b0;
  assign o[11] = t_9__1012_ | 1'b0;
  assign o[12] = t_9__1011_ | 1'b0;
  assign o[13] = t_9__1010_ | 1'b0;
  assign o[14] = t_9__1009_ | 1'b0;
  assign o[15] = t_9__1008_ | 1'b0;
  assign o[16] = t_9__1007_ | 1'b0;
  assign o[17] = t_9__1006_ | 1'b0;
  assign o[18] = t_9__1005_ | 1'b0;
  assign o[19] = t_9__1004_ | 1'b0;
  assign o[20] = t_9__1003_ | 1'b0;
  assign o[21] = t_9__1002_ | 1'b0;
  assign o[22] = t_9__1001_ | 1'b0;
  assign o[23] = t_9__1000_ | 1'b0;
  assign o[24] = t_9__999_ | 1'b0;
  assign o[25] = t_9__998_ | 1'b0;
  assign o[26] = t_9__997_ | 1'b0;
  assign o[27] = t_9__996_ | 1'b0;
  assign o[28] = t_9__995_ | 1'b0;
  assign o[29] = t_9__994_ | 1'b0;
  assign o[30] = t_9__993_ | 1'b0;
  assign o[31] = t_9__992_ | 1'b0;
  assign o[32] = t_9__991_ | 1'b0;
  assign o[33] = t_9__990_ | 1'b0;
  assign o[34] = t_9__989_ | 1'b0;
  assign o[35] = t_9__988_ | 1'b0;
  assign o[36] = t_9__987_ | 1'b0;
  assign o[37] = t_9__986_ | 1'b0;
  assign o[38] = t_9__985_ | 1'b0;
  assign o[39] = t_9__984_ | 1'b0;
  assign o[40] = t_9__983_ | 1'b0;
  assign o[41] = t_9__982_ | 1'b0;
  assign o[42] = t_9__981_ | 1'b0;
  assign o[43] = t_9__980_ | 1'b0;
  assign o[44] = t_9__979_ | 1'b0;
  assign o[45] = t_9__978_ | 1'b0;
  assign o[46] = t_9__977_ | 1'b0;
  assign o[47] = t_9__976_ | 1'b0;
  assign o[48] = t_9__975_ | 1'b0;
  assign o[49] = t_9__974_ | 1'b0;
  assign o[50] = t_9__973_ | 1'b0;
  assign o[51] = t_9__972_ | 1'b0;
  assign o[52] = t_9__971_ | 1'b0;
  assign o[53] = t_9__970_ | 1'b0;
  assign o[54] = t_9__969_ | 1'b0;
  assign o[55] = t_9__968_ | 1'b0;
  assign o[56] = t_9__967_ | 1'b0;
  assign o[57] = t_9__966_ | 1'b0;
  assign o[58] = t_9__965_ | 1'b0;
  assign o[59] = t_9__964_ | 1'b0;
  assign o[60] = t_9__963_ | 1'b0;
  assign o[61] = t_9__962_ | 1'b0;
  assign o[62] = t_9__961_ | 1'b0;
  assign o[63] = t_9__960_ | 1'b0;
  assign o[64] = t_9__959_ | 1'b0;
  assign o[65] = t_9__958_ | 1'b0;
  assign o[66] = t_9__957_ | 1'b0;
  assign o[67] = t_9__956_ | 1'b0;
  assign o[68] = t_9__955_ | 1'b0;
  assign o[69] = t_9__954_ | 1'b0;
  assign o[70] = t_9__953_ | 1'b0;
  assign o[71] = t_9__952_ | 1'b0;
  assign o[72] = t_9__951_ | 1'b0;
  assign o[73] = t_9__950_ | 1'b0;
  assign o[74] = t_9__949_ | 1'b0;
  assign o[75] = t_9__948_ | 1'b0;
  assign o[76] = t_9__947_ | 1'b0;
  assign o[77] = t_9__946_ | 1'b0;
  assign o[78] = t_9__945_ | 1'b0;
  assign o[79] = t_9__944_ | 1'b0;
  assign o[80] = t_9__943_ | 1'b0;
  assign o[81] = t_9__942_ | 1'b0;
  assign o[82] = t_9__941_ | 1'b0;
  assign o[83] = t_9__940_ | 1'b0;
  assign o[84] = t_9__939_ | 1'b0;
  assign o[85] = t_9__938_ | 1'b0;
  assign o[86] = t_9__937_ | 1'b0;
  assign o[87] = t_9__936_ | 1'b0;
  assign o[88] = t_9__935_ | 1'b0;
  assign o[89] = t_9__934_ | 1'b0;
  assign o[90] = t_9__933_ | 1'b0;
  assign o[91] = t_9__932_ | 1'b0;
  assign o[92] = t_9__931_ | 1'b0;
  assign o[93] = t_9__930_ | 1'b0;
  assign o[94] = t_9__929_ | 1'b0;
  assign o[95] = t_9__928_ | 1'b0;
  assign o[96] = t_9__927_ | 1'b0;
  assign o[97] = t_9__926_ | 1'b0;
  assign o[98] = t_9__925_ | 1'b0;
  assign o[99] = t_9__924_ | 1'b0;
  assign o[100] = t_9__923_ | 1'b0;
  assign o[101] = t_9__922_ | 1'b0;
  assign o[102] = t_9__921_ | 1'b0;
  assign o[103] = t_9__920_ | 1'b0;
  assign o[104] = t_9__919_ | 1'b0;
  assign o[105] = t_9__918_ | 1'b0;
  assign o[106] = t_9__917_ | 1'b0;
  assign o[107] = t_9__916_ | 1'b0;
  assign o[108] = t_9__915_ | 1'b0;
  assign o[109] = t_9__914_ | 1'b0;
  assign o[110] = t_9__913_ | 1'b0;
  assign o[111] = t_9__912_ | 1'b0;
  assign o[112] = t_9__911_ | 1'b0;
  assign o[113] = t_9__910_ | 1'b0;
  assign o[114] = t_9__909_ | 1'b0;
  assign o[115] = t_9__908_ | 1'b0;
  assign o[116] = t_9__907_ | 1'b0;
  assign o[117] = t_9__906_ | 1'b0;
  assign o[118] = t_9__905_ | 1'b0;
  assign o[119] = t_9__904_ | 1'b0;
  assign o[120] = t_9__903_ | 1'b0;
  assign o[121] = t_9__902_ | 1'b0;
  assign o[122] = t_9__901_ | 1'b0;
  assign o[123] = t_9__900_ | 1'b0;
  assign o[124] = t_9__899_ | 1'b0;
  assign o[125] = t_9__898_ | 1'b0;
  assign o[126] = t_9__897_ | 1'b0;
  assign o[127] = t_9__896_ | 1'b0;
  assign o[128] = t_9__895_ | 1'b0;
  assign o[129] = t_9__894_ | 1'b0;
  assign o[130] = t_9__893_ | 1'b0;
  assign o[131] = t_9__892_ | 1'b0;
  assign o[132] = t_9__891_ | 1'b0;
  assign o[133] = t_9__890_ | 1'b0;
  assign o[134] = t_9__889_ | 1'b0;
  assign o[135] = t_9__888_ | 1'b0;
  assign o[136] = t_9__887_ | 1'b0;
  assign o[137] = t_9__886_ | 1'b0;
  assign o[138] = t_9__885_ | 1'b0;
  assign o[139] = t_9__884_ | 1'b0;
  assign o[140] = t_9__883_ | 1'b0;
  assign o[141] = t_9__882_ | 1'b0;
  assign o[142] = t_9__881_ | 1'b0;
  assign o[143] = t_9__880_ | 1'b0;
  assign o[144] = t_9__879_ | 1'b0;
  assign o[145] = t_9__878_ | 1'b0;
  assign o[146] = t_9__877_ | 1'b0;
  assign o[147] = t_9__876_ | 1'b0;
  assign o[148] = t_9__875_ | 1'b0;
  assign o[149] = t_9__874_ | 1'b0;
  assign o[150] = t_9__873_ | 1'b0;
  assign o[151] = t_9__872_ | 1'b0;
  assign o[152] = t_9__871_ | 1'b0;
  assign o[153] = t_9__870_ | 1'b0;
  assign o[154] = t_9__869_ | 1'b0;
  assign o[155] = t_9__868_ | 1'b0;
  assign o[156] = t_9__867_ | 1'b0;
  assign o[157] = t_9__866_ | 1'b0;
  assign o[158] = t_9__865_ | 1'b0;
  assign o[159] = t_9__864_ | 1'b0;
  assign o[160] = t_9__863_ | 1'b0;
  assign o[161] = t_9__862_ | 1'b0;
  assign o[162] = t_9__861_ | 1'b0;
  assign o[163] = t_9__860_ | 1'b0;
  assign o[164] = t_9__859_ | 1'b0;
  assign o[165] = t_9__858_ | 1'b0;
  assign o[166] = t_9__857_ | 1'b0;
  assign o[167] = t_9__856_ | 1'b0;
  assign o[168] = t_9__855_ | 1'b0;
  assign o[169] = t_9__854_ | 1'b0;
  assign o[170] = t_9__853_ | 1'b0;
  assign o[171] = t_9__852_ | 1'b0;
  assign o[172] = t_9__851_ | 1'b0;
  assign o[173] = t_9__850_ | 1'b0;
  assign o[174] = t_9__849_ | 1'b0;
  assign o[175] = t_9__848_ | 1'b0;
  assign o[176] = t_9__847_ | 1'b0;
  assign o[177] = t_9__846_ | 1'b0;
  assign o[178] = t_9__845_ | 1'b0;
  assign o[179] = t_9__844_ | 1'b0;
  assign o[180] = t_9__843_ | 1'b0;
  assign o[181] = t_9__842_ | 1'b0;
  assign o[182] = t_9__841_ | 1'b0;
  assign o[183] = t_9__840_ | 1'b0;
  assign o[184] = t_9__839_ | 1'b0;
  assign o[185] = t_9__838_ | 1'b0;
  assign o[186] = t_9__837_ | 1'b0;
  assign o[187] = t_9__836_ | 1'b0;
  assign o[188] = t_9__835_ | 1'b0;
  assign o[189] = t_9__834_ | 1'b0;
  assign o[190] = t_9__833_ | 1'b0;
  assign o[191] = t_9__832_ | 1'b0;
  assign o[192] = t_9__831_ | 1'b0;
  assign o[193] = t_9__830_ | 1'b0;
  assign o[194] = t_9__829_ | 1'b0;
  assign o[195] = t_9__828_ | 1'b0;
  assign o[196] = t_9__827_ | 1'b0;
  assign o[197] = t_9__826_ | 1'b0;
  assign o[198] = t_9__825_ | 1'b0;
  assign o[199] = t_9__824_ | 1'b0;
  assign o[200] = t_9__823_ | 1'b0;
  assign o[201] = t_9__822_ | 1'b0;
  assign o[202] = t_9__821_ | 1'b0;
  assign o[203] = t_9__820_ | 1'b0;
  assign o[204] = t_9__819_ | 1'b0;
  assign o[205] = t_9__818_ | 1'b0;
  assign o[206] = t_9__817_ | 1'b0;
  assign o[207] = t_9__816_ | 1'b0;
  assign o[208] = t_9__815_ | 1'b0;
  assign o[209] = t_9__814_ | 1'b0;
  assign o[210] = t_9__813_ | 1'b0;
  assign o[211] = t_9__812_ | 1'b0;
  assign o[212] = t_9__811_ | 1'b0;
  assign o[213] = t_9__810_ | 1'b0;
  assign o[214] = t_9__809_ | 1'b0;
  assign o[215] = t_9__808_ | 1'b0;
  assign o[216] = t_9__807_ | 1'b0;
  assign o[217] = t_9__806_ | 1'b0;
  assign o[218] = t_9__805_ | 1'b0;
  assign o[219] = t_9__804_ | 1'b0;
  assign o[220] = t_9__803_ | 1'b0;
  assign o[221] = t_9__802_ | 1'b0;
  assign o[222] = t_9__801_ | 1'b0;
  assign o[223] = t_9__800_ | 1'b0;
  assign o[224] = t_9__799_ | 1'b0;
  assign o[225] = t_9__798_ | 1'b0;
  assign o[226] = t_9__797_ | 1'b0;
  assign o[227] = t_9__796_ | 1'b0;
  assign o[228] = t_9__795_ | 1'b0;
  assign o[229] = t_9__794_ | 1'b0;
  assign o[230] = t_9__793_ | 1'b0;
  assign o[231] = t_9__792_ | 1'b0;
  assign o[232] = t_9__791_ | 1'b0;
  assign o[233] = t_9__790_ | 1'b0;
  assign o[234] = t_9__789_ | 1'b0;
  assign o[235] = t_9__788_ | 1'b0;
  assign o[236] = t_9__787_ | 1'b0;
  assign o[237] = t_9__786_ | 1'b0;
  assign o[238] = t_9__785_ | 1'b0;
  assign o[239] = t_9__784_ | 1'b0;
  assign o[240] = t_9__783_ | 1'b0;
  assign o[241] = t_9__782_ | 1'b0;
  assign o[242] = t_9__781_ | 1'b0;
  assign o[243] = t_9__780_ | 1'b0;
  assign o[244] = t_9__779_ | 1'b0;
  assign o[245] = t_9__778_ | 1'b0;
  assign o[246] = t_9__777_ | 1'b0;
  assign o[247] = t_9__776_ | 1'b0;
  assign o[248] = t_9__775_ | 1'b0;
  assign o[249] = t_9__774_ | 1'b0;
  assign o[250] = t_9__773_ | 1'b0;
  assign o[251] = t_9__772_ | 1'b0;
  assign o[252] = t_9__771_ | 1'b0;
  assign o[253] = t_9__770_ | 1'b0;
  assign o[254] = t_9__769_ | 1'b0;
  assign o[255] = t_9__768_ | 1'b0;
  assign o[256] = t_9__767_ | 1'b0;
  assign o[257] = t_9__766_ | 1'b0;
  assign o[258] = t_9__765_ | 1'b0;
  assign o[259] = t_9__764_ | 1'b0;
  assign o[260] = t_9__763_ | 1'b0;
  assign o[261] = t_9__762_ | 1'b0;
  assign o[262] = t_9__761_ | 1'b0;
  assign o[263] = t_9__760_ | 1'b0;
  assign o[264] = t_9__759_ | 1'b0;
  assign o[265] = t_9__758_ | 1'b0;
  assign o[266] = t_9__757_ | 1'b0;
  assign o[267] = t_9__756_ | 1'b0;
  assign o[268] = t_9__755_ | 1'b0;
  assign o[269] = t_9__754_ | 1'b0;
  assign o[270] = t_9__753_ | 1'b0;
  assign o[271] = t_9__752_ | 1'b0;
  assign o[272] = t_9__751_ | 1'b0;
  assign o[273] = t_9__750_ | 1'b0;
  assign o[274] = t_9__749_ | 1'b0;
  assign o[275] = t_9__748_ | 1'b0;
  assign o[276] = t_9__747_ | 1'b0;
  assign o[277] = t_9__746_ | 1'b0;
  assign o[278] = t_9__745_ | 1'b0;
  assign o[279] = t_9__744_ | 1'b0;
  assign o[280] = t_9__743_ | 1'b0;
  assign o[281] = t_9__742_ | 1'b0;
  assign o[282] = t_9__741_ | 1'b0;
  assign o[283] = t_9__740_ | 1'b0;
  assign o[284] = t_9__739_ | 1'b0;
  assign o[285] = t_9__738_ | 1'b0;
  assign o[286] = t_9__737_ | 1'b0;
  assign o[287] = t_9__736_ | 1'b0;
  assign o[288] = t_9__735_ | 1'b0;
  assign o[289] = t_9__734_ | 1'b0;
  assign o[290] = t_9__733_ | 1'b0;
  assign o[291] = t_9__732_ | 1'b0;
  assign o[292] = t_9__731_ | 1'b0;
  assign o[293] = t_9__730_ | 1'b0;
  assign o[294] = t_9__729_ | 1'b0;
  assign o[295] = t_9__728_ | 1'b0;
  assign o[296] = t_9__727_ | 1'b0;
  assign o[297] = t_9__726_ | 1'b0;
  assign o[298] = t_9__725_ | 1'b0;
  assign o[299] = t_9__724_ | 1'b0;
  assign o[300] = t_9__723_ | 1'b0;
  assign o[301] = t_9__722_ | 1'b0;
  assign o[302] = t_9__721_ | 1'b0;
  assign o[303] = t_9__720_ | 1'b0;
  assign o[304] = t_9__719_ | 1'b0;
  assign o[305] = t_9__718_ | 1'b0;
  assign o[306] = t_9__717_ | 1'b0;
  assign o[307] = t_9__716_ | 1'b0;
  assign o[308] = t_9__715_ | 1'b0;
  assign o[309] = t_9__714_ | 1'b0;
  assign o[310] = t_9__713_ | 1'b0;
  assign o[311] = t_9__712_ | 1'b0;
  assign o[312] = t_9__711_ | 1'b0;
  assign o[313] = t_9__710_ | 1'b0;
  assign o[314] = t_9__709_ | 1'b0;
  assign o[315] = t_9__708_ | 1'b0;
  assign o[316] = t_9__707_ | 1'b0;
  assign o[317] = t_9__706_ | 1'b0;
  assign o[318] = t_9__705_ | 1'b0;
  assign o[319] = t_9__704_ | 1'b0;
  assign o[320] = t_9__703_ | 1'b0;
  assign o[321] = t_9__702_ | 1'b0;
  assign o[322] = t_9__701_ | 1'b0;
  assign o[323] = t_9__700_ | 1'b0;
  assign o[324] = t_9__699_ | 1'b0;
  assign o[325] = t_9__698_ | 1'b0;
  assign o[326] = t_9__697_ | 1'b0;
  assign o[327] = t_9__696_ | 1'b0;
  assign o[328] = t_9__695_ | 1'b0;
  assign o[329] = t_9__694_ | 1'b0;
  assign o[330] = t_9__693_ | 1'b0;
  assign o[331] = t_9__692_ | 1'b0;
  assign o[332] = t_9__691_ | 1'b0;
  assign o[333] = t_9__690_ | 1'b0;
  assign o[334] = t_9__689_ | 1'b0;
  assign o[335] = t_9__688_ | 1'b0;
  assign o[336] = t_9__687_ | 1'b0;
  assign o[337] = t_9__686_ | 1'b0;
  assign o[338] = t_9__685_ | 1'b0;
  assign o[339] = t_9__684_ | 1'b0;
  assign o[340] = t_9__683_ | 1'b0;
  assign o[341] = t_9__682_ | 1'b0;
  assign o[342] = t_9__681_ | 1'b0;
  assign o[343] = t_9__680_ | 1'b0;
  assign o[344] = t_9__679_ | 1'b0;
  assign o[345] = t_9__678_ | 1'b0;
  assign o[346] = t_9__677_ | 1'b0;
  assign o[347] = t_9__676_ | 1'b0;
  assign o[348] = t_9__675_ | 1'b0;
  assign o[349] = t_9__674_ | 1'b0;
  assign o[350] = t_9__673_ | 1'b0;
  assign o[351] = t_9__672_ | 1'b0;
  assign o[352] = t_9__671_ | 1'b0;
  assign o[353] = t_9__670_ | 1'b0;
  assign o[354] = t_9__669_ | 1'b0;
  assign o[355] = t_9__668_ | 1'b0;
  assign o[356] = t_9__667_ | 1'b0;
  assign o[357] = t_9__666_ | 1'b0;
  assign o[358] = t_9__665_ | 1'b0;
  assign o[359] = t_9__664_ | 1'b0;
  assign o[360] = t_9__663_ | 1'b0;
  assign o[361] = t_9__662_ | 1'b0;
  assign o[362] = t_9__661_ | 1'b0;
  assign o[363] = t_9__660_ | 1'b0;
  assign o[364] = t_9__659_ | 1'b0;
  assign o[365] = t_9__658_ | 1'b0;
  assign o[366] = t_9__657_ | 1'b0;
  assign o[367] = t_9__656_ | 1'b0;
  assign o[368] = t_9__655_ | 1'b0;
  assign o[369] = t_9__654_ | 1'b0;
  assign o[370] = t_9__653_ | 1'b0;
  assign o[371] = t_9__652_ | 1'b0;
  assign o[372] = t_9__651_ | 1'b0;
  assign o[373] = t_9__650_ | 1'b0;
  assign o[374] = t_9__649_ | 1'b0;
  assign o[375] = t_9__648_ | 1'b0;
  assign o[376] = t_9__647_ | 1'b0;
  assign o[377] = t_9__646_ | 1'b0;
  assign o[378] = t_9__645_ | 1'b0;
  assign o[379] = t_9__644_ | 1'b0;
  assign o[380] = t_9__643_ | 1'b0;
  assign o[381] = t_9__642_ | 1'b0;
  assign o[382] = t_9__641_ | 1'b0;
  assign o[383] = t_9__640_ | 1'b0;
  assign o[384] = t_9__639_ | 1'b0;
  assign o[385] = t_9__638_ | 1'b0;
  assign o[386] = t_9__637_ | 1'b0;
  assign o[387] = t_9__636_ | 1'b0;
  assign o[388] = t_9__635_ | 1'b0;
  assign o[389] = t_9__634_ | 1'b0;
  assign o[390] = t_9__633_ | 1'b0;
  assign o[391] = t_9__632_ | 1'b0;
  assign o[392] = t_9__631_ | 1'b0;
  assign o[393] = t_9__630_ | 1'b0;
  assign o[394] = t_9__629_ | 1'b0;
  assign o[395] = t_9__628_ | 1'b0;
  assign o[396] = t_9__627_ | 1'b0;
  assign o[397] = t_9__626_ | 1'b0;
  assign o[398] = t_9__625_ | 1'b0;
  assign o[399] = t_9__624_ | 1'b0;
  assign o[400] = t_9__623_ | 1'b0;
  assign o[401] = t_9__622_ | 1'b0;
  assign o[402] = t_9__621_ | 1'b0;
  assign o[403] = t_9__620_ | 1'b0;
  assign o[404] = t_9__619_ | 1'b0;
  assign o[405] = t_9__618_ | 1'b0;
  assign o[406] = t_9__617_ | 1'b0;
  assign o[407] = t_9__616_ | 1'b0;
  assign o[408] = t_9__615_ | 1'b0;
  assign o[409] = t_9__614_ | 1'b0;
  assign o[410] = t_9__613_ | 1'b0;
  assign o[411] = t_9__612_ | 1'b0;
  assign o[412] = t_9__611_ | 1'b0;
  assign o[413] = t_9__610_ | 1'b0;
  assign o[414] = t_9__609_ | 1'b0;
  assign o[415] = t_9__608_ | 1'b0;
  assign o[416] = t_9__607_ | 1'b0;
  assign o[417] = t_9__606_ | 1'b0;
  assign o[418] = t_9__605_ | 1'b0;
  assign o[419] = t_9__604_ | 1'b0;
  assign o[420] = t_9__603_ | 1'b0;
  assign o[421] = t_9__602_ | 1'b0;
  assign o[422] = t_9__601_ | 1'b0;
  assign o[423] = t_9__600_ | 1'b0;
  assign o[424] = t_9__599_ | 1'b0;
  assign o[425] = t_9__598_ | 1'b0;
  assign o[426] = t_9__597_ | 1'b0;
  assign o[427] = t_9__596_ | 1'b0;
  assign o[428] = t_9__595_ | 1'b0;
  assign o[429] = t_9__594_ | 1'b0;
  assign o[430] = t_9__593_ | 1'b0;
  assign o[431] = t_9__592_ | 1'b0;
  assign o[432] = t_9__591_ | 1'b0;
  assign o[433] = t_9__590_ | 1'b0;
  assign o[434] = t_9__589_ | 1'b0;
  assign o[435] = t_9__588_ | 1'b0;
  assign o[436] = t_9__587_ | 1'b0;
  assign o[437] = t_9__586_ | 1'b0;
  assign o[438] = t_9__585_ | 1'b0;
  assign o[439] = t_9__584_ | 1'b0;
  assign o[440] = t_9__583_ | 1'b0;
  assign o[441] = t_9__582_ | 1'b0;
  assign o[442] = t_9__581_ | 1'b0;
  assign o[443] = t_9__580_ | 1'b0;
  assign o[444] = t_9__579_ | 1'b0;
  assign o[445] = t_9__578_ | 1'b0;
  assign o[446] = t_9__577_ | 1'b0;
  assign o[447] = t_9__576_ | 1'b0;
  assign o[448] = t_9__575_ | 1'b0;
  assign o[449] = t_9__574_ | 1'b0;
  assign o[450] = t_9__573_ | 1'b0;
  assign o[451] = t_9__572_ | 1'b0;
  assign o[452] = t_9__571_ | 1'b0;
  assign o[453] = t_9__570_ | 1'b0;
  assign o[454] = t_9__569_ | 1'b0;
  assign o[455] = t_9__568_ | 1'b0;
  assign o[456] = t_9__567_ | 1'b0;
  assign o[457] = t_9__566_ | 1'b0;
  assign o[458] = t_9__565_ | 1'b0;
  assign o[459] = t_9__564_ | 1'b0;
  assign o[460] = t_9__563_ | 1'b0;
  assign o[461] = t_9__562_ | 1'b0;
  assign o[462] = t_9__561_ | 1'b0;
  assign o[463] = t_9__560_ | 1'b0;
  assign o[464] = t_9__559_ | 1'b0;
  assign o[465] = t_9__558_ | 1'b0;
  assign o[466] = t_9__557_ | 1'b0;
  assign o[467] = t_9__556_ | 1'b0;
  assign o[468] = t_9__555_ | 1'b0;
  assign o[469] = t_9__554_ | 1'b0;
  assign o[470] = t_9__553_ | 1'b0;
  assign o[471] = t_9__552_ | 1'b0;
  assign o[472] = t_9__551_ | 1'b0;
  assign o[473] = t_9__550_ | 1'b0;
  assign o[474] = t_9__549_ | 1'b0;
  assign o[475] = t_9__548_ | 1'b0;
  assign o[476] = t_9__547_ | 1'b0;
  assign o[477] = t_9__546_ | 1'b0;
  assign o[478] = t_9__545_ | 1'b0;
  assign o[479] = t_9__544_ | 1'b0;
  assign o[480] = t_9__543_ | 1'b0;
  assign o[481] = t_9__542_ | 1'b0;
  assign o[482] = t_9__541_ | 1'b0;
  assign o[483] = t_9__540_ | 1'b0;
  assign o[484] = t_9__539_ | 1'b0;
  assign o[485] = t_9__538_ | 1'b0;
  assign o[486] = t_9__537_ | 1'b0;
  assign o[487] = t_9__536_ | 1'b0;
  assign o[488] = t_9__535_ | 1'b0;
  assign o[489] = t_9__534_ | 1'b0;
  assign o[490] = t_9__533_ | 1'b0;
  assign o[491] = t_9__532_ | 1'b0;
  assign o[492] = t_9__531_ | 1'b0;
  assign o[493] = t_9__530_ | 1'b0;
  assign o[494] = t_9__529_ | 1'b0;
  assign o[495] = t_9__528_ | 1'b0;
  assign o[496] = t_9__527_ | 1'b0;
  assign o[497] = t_9__526_ | 1'b0;
  assign o[498] = t_9__525_ | 1'b0;
  assign o[499] = t_9__524_ | 1'b0;
  assign o[500] = t_9__523_ | 1'b0;
  assign o[501] = t_9__522_ | 1'b0;
  assign o[502] = t_9__521_ | 1'b0;
  assign o[503] = t_9__520_ | 1'b0;
  assign o[504] = t_9__519_ | 1'b0;
  assign o[505] = t_9__518_ | 1'b0;
  assign o[506] = t_9__517_ | 1'b0;
  assign o[507] = t_9__516_ | 1'b0;
  assign o[508] = t_9__515_ | 1'b0;
  assign o[509] = t_9__514_ | 1'b0;
  assign o[510] = t_9__513_ | 1'b0;
  assign o[511] = t_9__512_ | 1'b0;
  assign o[512] = t_9__511_ | t_9__1023_;
  assign o[513] = t_9__510_ | t_9__1022_;
  assign o[514] = t_9__509_ | t_9__1021_;
  assign o[515] = t_9__508_ | t_9__1020_;
  assign o[516] = t_9__507_ | t_9__1019_;
  assign o[517] = t_9__506_ | t_9__1018_;
  assign o[518] = t_9__505_ | t_9__1017_;
  assign o[519] = t_9__504_ | t_9__1016_;
  assign o[520] = t_9__503_ | t_9__1015_;
  assign o[521] = t_9__502_ | t_9__1014_;
  assign o[522] = t_9__501_ | t_9__1013_;
  assign o[523] = t_9__500_ | t_9__1012_;
  assign o[524] = t_9__499_ | t_9__1011_;
  assign o[525] = t_9__498_ | t_9__1010_;
  assign o[526] = t_9__497_ | t_9__1009_;
  assign o[527] = t_9__496_ | t_9__1008_;
  assign o[528] = t_9__495_ | t_9__1007_;
  assign o[529] = t_9__494_ | t_9__1006_;
  assign o[530] = t_9__493_ | t_9__1005_;
  assign o[531] = t_9__492_ | t_9__1004_;
  assign o[532] = t_9__491_ | t_9__1003_;
  assign o[533] = t_9__490_ | t_9__1002_;
  assign o[534] = t_9__489_ | t_9__1001_;
  assign o[535] = t_9__488_ | t_9__1000_;
  assign o[536] = t_9__487_ | t_9__999_;
  assign o[537] = t_9__486_ | t_9__998_;
  assign o[538] = t_9__485_ | t_9__997_;
  assign o[539] = t_9__484_ | t_9__996_;
  assign o[540] = t_9__483_ | t_9__995_;
  assign o[541] = t_9__482_ | t_9__994_;
  assign o[542] = t_9__481_ | t_9__993_;
  assign o[543] = t_9__480_ | t_9__992_;
  assign o[544] = t_9__479_ | t_9__991_;
  assign o[545] = t_9__478_ | t_9__990_;
  assign o[546] = t_9__477_ | t_9__989_;
  assign o[547] = t_9__476_ | t_9__988_;
  assign o[548] = t_9__475_ | t_9__987_;
  assign o[549] = t_9__474_ | t_9__986_;
  assign o[550] = t_9__473_ | t_9__985_;
  assign o[551] = t_9__472_ | t_9__984_;
  assign o[552] = t_9__471_ | t_9__983_;
  assign o[553] = t_9__470_ | t_9__982_;
  assign o[554] = t_9__469_ | t_9__981_;
  assign o[555] = t_9__468_ | t_9__980_;
  assign o[556] = t_9__467_ | t_9__979_;
  assign o[557] = t_9__466_ | t_9__978_;
  assign o[558] = t_9__465_ | t_9__977_;
  assign o[559] = t_9__464_ | t_9__976_;
  assign o[560] = t_9__463_ | t_9__975_;
  assign o[561] = t_9__462_ | t_9__974_;
  assign o[562] = t_9__461_ | t_9__973_;
  assign o[563] = t_9__460_ | t_9__972_;
  assign o[564] = t_9__459_ | t_9__971_;
  assign o[565] = t_9__458_ | t_9__970_;
  assign o[566] = t_9__457_ | t_9__969_;
  assign o[567] = t_9__456_ | t_9__968_;
  assign o[568] = t_9__455_ | t_9__967_;
  assign o[569] = t_9__454_ | t_9__966_;
  assign o[570] = t_9__453_ | t_9__965_;
  assign o[571] = t_9__452_ | t_9__964_;
  assign o[572] = t_9__451_ | t_9__963_;
  assign o[573] = t_9__450_ | t_9__962_;
  assign o[574] = t_9__449_ | t_9__961_;
  assign o[575] = t_9__448_ | t_9__960_;
  assign o[576] = t_9__447_ | t_9__959_;
  assign o[577] = t_9__446_ | t_9__958_;
  assign o[578] = t_9__445_ | t_9__957_;
  assign o[579] = t_9__444_ | t_9__956_;
  assign o[580] = t_9__443_ | t_9__955_;
  assign o[581] = t_9__442_ | t_9__954_;
  assign o[582] = t_9__441_ | t_9__953_;
  assign o[583] = t_9__440_ | t_9__952_;
  assign o[584] = t_9__439_ | t_9__951_;
  assign o[585] = t_9__438_ | t_9__950_;
  assign o[586] = t_9__437_ | t_9__949_;
  assign o[587] = t_9__436_ | t_9__948_;
  assign o[588] = t_9__435_ | t_9__947_;
  assign o[589] = t_9__434_ | t_9__946_;
  assign o[590] = t_9__433_ | t_9__945_;
  assign o[591] = t_9__432_ | t_9__944_;
  assign o[592] = t_9__431_ | t_9__943_;
  assign o[593] = t_9__430_ | t_9__942_;
  assign o[594] = t_9__429_ | t_9__941_;
  assign o[595] = t_9__428_ | t_9__940_;
  assign o[596] = t_9__427_ | t_9__939_;
  assign o[597] = t_9__426_ | t_9__938_;
  assign o[598] = t_9__425_ | t_9__937_;
  assign o[599] = t_9__424_ | t_9__936_;
  assign o[600] = t_9__423_ | t_9__935_;
  assign o[601] = t_9__422_ | t_9__934_;
  assign o[602] = t_9__421_ | t_9__933_;
  assign o[603] = t_9__420_ | t_9__932_;
  assign o[604] = t_9__419_ | t_9__931_;
  assign o[605] = t_9__418_ | t_9__930_;
  assign o[606] = t_9__417_ | t_9__929_;
  assign o[607] = t_9__416_ | t_9__928_;
  assign o[608] = t_9__415_ | t_9__927_;
  assign o[609] = t_9__414_ | t_9__926_;
  assign o[610] = t_9__413_ | t_9__925_;
  assign o[611] = t_9__412_ | t_9__924_;
  assign o[612] = t_9__411_ | t_9__923_;
  assign o[613] = t_9__410_ | t_9__922_;
  assign o[614] = t_9__409_ | t_9__921_;
  assign o[615] = t_9__408_ | t_9__920_;
  assign o[616] = t_9__407_ | t_9__919_;
  assign o[617] = t_9__406_ | t_9__918_;
  assign o[618] = t_9__405_ | t_9__917_;
  assign o[619] = t_9__404_ | t_9__916_;
  assign o[620] = t_9__403_ | t_9__915_;
  assign o[621] = t_9__402_ | t_9__914_;
  assign o[622] = t_9__401_ | t_9__913_;
  assign o[623] = t_9__400_ | t_9__912_;
  assign o[624] = t_9__399_ | t_9__911_;
  assign o[625] = t_9__398_ | t_9__910_;
  assign o[626] = t_9__397_ | t_9__909_;
  assign o[627] = t_9__396_ | t_9__908_;
  assign o[628] = t_9__395_ | t_9__907_;
  assign o[629] = t_9__394_ | t_9__906_;
  assign o[630] = t_9__393_ | t_9__905_;
  assign o[631] = t_9__392_ | t_9__904_;
  assign o[632] = t_9__391_ | t_9__903_;
  assign o[633] = t_9__390_ | t_9__902_;
  assign o[634] = t_9__389_ | t_9__901_;
  assign o[635] = t_9__388_ | t_9__900_;
  assign o[636] = t_9__387_ | t_9__899_;
  assign o[637] = t_9__386_ | t_9__898_;
  assign o[638] = t_9__385_ | t_9__897_;
  assign o[639] = t_9__384_ | t_9__896_;
  assign o[640] = t_9__383_ | t_9__895_;
  assign o[641] = t_9__382_ | t_9__894_;
  assign o[642] = t_9__381_ | t_9__893_;
  assign o[643] = t_9__380_ | t_9__892_;
  assign o[644] = t_9__379_ | t_9__891_;
  assign o[645] = t_9__378_ | t_9__890_;
  assign o[646] = t_9__377_ | t_9__889_;
  assign o[647] = t_9__376_ | t_9__888_;
  assign o[648] = t_9__375_ | t_9__887_;
  assign o[649] = t_9__374_ | t_9__886_;
  assign o[650] = t_9__373_ | t_9__885_;
  assign o[651] = t_9__372_ | t_9__884_;
  assign o[652] = t_9__371_ | t_9__883_;
  assign o[653] = t_9__370_ | t_9__882_;
  assign o[654] = t_9__369_ | t_9__881_;
  assign o[655] = t_9__368_ | t_9__880_;
  assign o[656] = t_9__367_ | t_9__879_;
  assign o[657] = t_9__366_ | t_9__878_;
  assign o[658] = t_9__365_ | t_9__877_;
  assign o[659] = t_9__364_ | t_9__876_;
  assign o[660] = t_9__363_ | t_9__875_;
  assign o[661] = t_9__362_ | t_9__874_;
  assign o[662] = t_9__361_ | t_9__873_;
  assign o[663] = t_9__360_ | t_9__872_;
  assign o[664] = t_9__359_ | t_9__871_;
  assign o[665] = t_9__358_ | t_9__870_;
  assign o[666] = t_9__357_ | t_9__869_;
  assign o[667] = t_9__356_ | t_9__868_;
  assign o[668] = t_9__355_ | t_9__867_;
  assign o[669] = t_9__354_ | t_9__866_;
  assign o[670] = t_9__353_ | t_9__865_;
  assign o[671] = t_9__352_ | t_9__864_;
  assign o[672] = t_9__351_ | t_9__863_;
  assign o[673] = t_9__350_ | t_9__862_;
  assign o[674] = t_9__349_ | t_9__861_;
  assign o[675] = t_9__348_ | t_9__860_;
  assign o[676] = t_9__347_ | t_9__859_;
  assign o[677] = t_9__346_ | t_9__858_;
  assign o[678] = t_9__345_ | t_9__857_;
  assign o[679] = t_9__344_ | t_9__856_;
  assign o[680] = t_9__343_ | t_9__855_;
  assign o[681] = t_9__342_ | t_9__854_;
  assign o[682] = t_9__341_ | t_9__853_;
  assign o[683] = t_9__340_ | t_9__852_;
  assign o[684] = t_9__339_ | t_9__851_;
  assign o[685] = t_9__338_ | t_9__850_;
  assign o[686] = t_9__337_ | t_9__849_;
  assign o[687] = t_9__336_ | t_9__848_;
  assign o[688] = t_9__335_ | t_9__847_;
  assign o[689] = t_9__334_ | t_9__846_;
  assign o[690] = t_9__333_ | t_9__845_;
  assign o[691] = t_9__332_ | t_9__844_;
  assign o[692] = t_9__331_ | t_9__843_;
  assign o[693] = t_9__330_ | t_9__842_;
  assign o[694] = t_9__329_ | t_9__841_;
  assign o[695] = t_9__328_ | t_9__840_;
  assign o[696] = t_9__327_ | t_9__839_;
  assign o[697] = t_9__326_ | t_9__838_;
  assign o[698] = t_9__325_ | t_9__837_;
  assign o[699] = t_9__324_ | t_9__836_;
  assign o[700] = t_9__323_ | t_9__835_;
  assign o[701] = t_9__322_ | t_9__834_;
  assign o[702] = t_9__321_ | t_9__833_;
  assign o[703] = t_9__320_ | t_9__832_;
  assign o[704] = t_9__319_ | t_9__831_;
  assign o[705] = t_9__318_ | t_9__830_;
  assign o[706] = t_9__317_ | t_9__829_;
  assign o[707] = t_9__316_ | t_9__828_;
  assign o[708] = t_9__315_ | t_9__827_;
  assign o[709] = t_9__314_ | t_9__826_;
  assign o[710] = t_9__313_ | t_9__825_;
  assign o[711] = t_9__312_ | t_9__824_;
  assign o[712] = t_9__311_ | t_9__823_;
  assign o[713] = t_9__310_ | t_9__822_;
  assign o[714] = t_9__309_ | t_9__821_;
  assign o[715] = t_9__308_ | t_9__820_;
  assign o[716] = t_9__307_ | t_9__819_;
  assign o[717] = t_9__306_ | t_9__818_;
  assign o[718] = t_9__305_ | t_9__817_;
  assign o[719] = t_9__304_ | t_9__816_;
  assign o[720] = t_9__303_ | t_9__815_;
  assign o[721] = t_9__302_ | t_9__814_;
  assign o[722] = t_9__301_ | t_9__813_;
  assign o[723] = t_9__300_ | t_9__812_;
  assign o[724] = t_9__299_ | t_9__811_;
  assign o[725] = t_9__298_ | t_9__810_;
  assign o[726] = t_9__297_ | t_9__809_;
  assign o[727] = t_9__296_ | t_9__808_;
  assign o[728] = t_9__295_ | t_9__807_;
  assign o[729] = t_9__294_ | t_9__806_;
  assign o[730] = t_9__293_ | t_9__805_;
  assign o[731] = t_9__292_ | t_9__804_;
  assign o[732] = t_9__291_ | t_9__803_;
  assign o[733] = t_9__290_ | t_9__802_;
  assign o[734] = t_9__289_ | t_9__801_;
  assign o[735] = t_9__288_ | t_9__800_;
  assign o[736] = t_9__287_ | t_9__799_;
  assign o[737] = t_9__286_ | t_9__798_;
  assign o[738] = t_9__285_ | t_9__797_;
  assign o[739] = t_9__284_ | t_9__796_;
  assign o[740] = t_9__283_ | t_9__795_;
  assign o[741] = t_9__282_ | t_9__794_;
  assign o[742] = t_9__281_ | t_9__793_;
  assign o[743] = t_9__280_ | t_9__792_;
  assign o[744] = t_9__279_ | t_9__791_;
  assign o[745] = t_9__278_ | t_9__790_;
  assign o[746] = t_9__277_ | t_9__789_;
  assign o[747] = t_9__276_ | t_9__788_;
  assign o[748] = t_9__275_ | t_9__787_;
  assign o[749] = t_9__274_ | t_9__786_;
  assign o[750] = t_9__273_ | t_9__785_;
  assign o[751] = t_9__272_ | t_9__784_;
  assign o[752] = t_9__271_ | t_9__783_;
  assign o[753] = t_9__270_ | t_9__782_;
  assign o[754] = t_9__269_ | t_9__781_;
  assign o[755] = t_9__268_ | t_9__780_;
  assign o[756] = t_9__267_ | t_9__779_;
  assign o[757] = t_9__266_ | t_9__778_;
  assign o[758] = t_9__265_ | t_9__777_;
  assign o[759] = t_9__264_ | t_9__776_;
  assign o[760] = t_9__263_ | t_9__775_;
  assign o[761] = t_9__262_ | t_9__774_;
  assign o[762] = t_9__261_ | t_9__773_;
  assign o[763] = t_9__260_ | t_9__772_;
  assign o[764] = t_9__259_ | t_9__771_;
  assign o[765] = t_9__258_ | t_9__770_;
  assign o[766] = t_9__257_ | t_9__769_;
  assign o[767] = t_9__256_ | t_9__768_;
  assign o[768] = t_9__255_ | t_9__767_;
  assign o[769] = t_9__254_ | t_9__766_;
  assign o[770] = t_9__253_ | t_9__765_;
  assign o[771] = t_9__252_ | t_9__764_;
  assign o[772] = t_9__251_ | t_9__763_;
  assign o[773] = t_9__250_ | t_9__762_;
  assign o[774] = t_9__249_ | t_9__761_;
  assign o[775] = t_9__248_ | t_9__760_;
  assign o[776] = t_9__247_ | t_9__759_;
  assign o[777] = t_9__246_ | t_9__758_;
  assign o[778] = t_9__245_ | t_9__757_;
  assign o[779] = t_9__244_ | t_9__756_;
  assign o[780] = t_9__243_ | t_9__755_;
  assign o[781] = t_9__242_ | t_9__754_;
  assign o[782] = t_9__241_ | t_9__753_;
  assign o[783] = t_9__240_ | t_9__752_;
  assign o[784] = t_9__239_ | t_9__751_;
  assign o[785] = t_9__238_ | t_9__750_;
  assign o[786] = t_9__237_ | t_9__749_;
  assign o[787] = t_9__236_ | t_9__748_;
  assign o[788] = t_9__235_ | t_9__747_;
  assign o[789] = t_9__234_ | t_9__746_;
  assign o[790] = t_9__233_ | t_9__745_;
  assign o[791] = t_9__232_ | t_9__744_;
  assign o[792] = t_9__231_ | t_9__743_;
  assign o[793] = t_9__230_ | t_9__742_;
  assign o[794] = t_9__229_ | t_9__741_;
  assign o[795] = t_9__228_ | t_9__740_;
  assign o[796] = t_9__227_ | t_9__739_;
  assign o[797] = t_9__226_ | t_9__738_;
  assign o[798] = t_9__225_ | t_9__737_;
  assign o[799] = t_9__224_ | t_9__736_;
  assign o[800] = t_9__223_ | t_9__735_;
  assign o[801] = t_9__222_ | t_9__734_;
  assign o[802] = t_9__221_ | t_9__733_;
  assign o[803] = t_9__220_ | t_9__732_;
  assign o[804] = t_9__219_ | t_9__731_;
  assign o[805] = t_9__218_ | t_9__730_;
  assign o[806] = t_9__217_ | t_9__729_;
  assign o[807] = t_9__216_ | t_9__728_;
  assign o[808] = t_9__215_ | t_9__727_;
  assign o[809] = t_9__214_ | t_9__726_;
  assign o[810] = t_9__213_ | t_9__725_;
  assign o[811] = t_9__212_ | t_9__724_;
  assign o[812] = t_9__211_ | t_9__723_;
  assign o[813] = t_9__210_ | t_9__722_;
  assign o[814] = t_9__209_ | t_9__721_;
  assign o[815] = t_9__208_ | t_9__720_;
  assign o[816] = t_9__207_ | t_9__719_;
  assign o[817] = t_9__206_ | t_9__718_;
  assign o[818] = t_9__205_ | t_9__717_;
  assign o[819] = t_9__204_ | t_9__716_;
  assign o[820] = t_9__203_ | t_9__715_;
  assign o[821] = t_9__202_ | t_9__714_;
  assign o[822] = t_9__201_ | t_9__713_;
  assign o[823] = t_9__200_ | t_9__712_;
  assign o[824] = t_9__199_ | t_9__711_;
  assign o[825] = t_9__198_ | t_9__710_;
  assign o[826] = t_9__197_ | t_9__709_;
  assign o[827] = t_9__196_ | t_9__708_;
  assign o[828] = t_9__195_ | t_9__707_;
  assign o[829] = t_9__194_ | t_9__706_;
  assign o[830] = t_9__193_ | t_9__705_;
  assign o[831] = t_9__192_ | t_9__704_;
  assign o[832] = t_9__191_ | t_9__703_;
  assign o[833] = t_9__190_ | t_9__702_;
  assign o[834] = t_9__189_ | t_9__701_;
  assign o[835] = t_9__188_ | t_9__700_;
  assign o[836] = t_9__187_ | t_9__699_;
  assign o[837] = t_9__186_ | t_9__698_;
  assign o[838] = t_9__185_ | t_9__697_;
  assign o[839] = t_9__184_ | t_9__696_;
  assign o[840] = t_9__183_ | t_9__695_;
  assign o[841] = t_9__182_ | t_9__694_;
  assign o[842] = t_9__181_ | t_9__693_;
  assign o[843] = t_9__180_ | t_9__692_;
  assign o[844] = t_9__179_ | t_9__691_;
  assign o[845] = t_9__178_ | t_9__690_;
  assign o[846] = t_9__177_ | t_9__689_;
  assign o[847] = t_9__176_ | t_9__688_;
  assign o[848] = t_9__175_ | t_9__687_;
  assign o[849] = t_9__174_ | t_9__686_;
  assign o[850] = t_9__173_ | t_9__685_;
  assign o[851] = t_9__172_ | t_9__684_;
  assign o[852] = t_9__171_ | t_9__683_;
  assign o[853] = t_9__170_ | t_9__682_;
  assign o[854] = t_9__169_ | t_9__681_;
  assign o[855] = t_9__168_ | t_9__680_;
  assign o[856] = t_9__167_ | t_9__679_;
  assign o[857] = t_9__166_ | t_9__678_;
  assign o[858] = t_9__165_ | t_9__677_;
  assign o[859] = t_9__164_ | t_9__676_;
  assign o[860] = t_9__163_ | t_9__675_;
  assign o[861] = t_9__162_ | t_9__674_;
  assign o[862] = t_9__161_ | t_9__673_;
  assign o[863] = t_9__160_ | t_9__672_;
  assign o[864] = t_9__159_ | t_9__671_;
  assign o[865] = t_9__158_ | t_9__670_;
  assign o[866] = t_9__157_ | t_9__669_;
  assign o[867] = t_9__156_ | t_9__668_;
  assign o[868] = t_9__155_ | t_9__667_;
  assign o[869] = t_9__154_ | t_9__666_;
  assign o[870] = t_9__153_ | t_9__665_;
  assign o[871] = t_9__152_ | t_9__664_;
  assign o[872] = t_9__151_ | t_9__663_;
  assign o[873] = t_9__150_ | t_9__662_;
  assign o[874] = t_9__149_ | t_9__661_;
  assign o[875] = t_9__148_ | t_9__660_;
  assign o[876] = t_9__147_ | t_9__659_;
  assign o[877] = t_9__146_ | t_9__658_;
  assign o[878] = t_9__145_ | t_9__657_;
  assign o[879] = t_9__144_ | t_9__656_;
  assign o[880] = t_9__143_ | t_9__655_;
  assign o[881] = t_9__142_ | t_9__654_;
  assign o[882] = t_9__141_ | t_9__653_;
  assign o[883] = t_9__140_ | t_9__652_;
  assign o[884] = t_9__139_ | t_9__651_;
  assign o[885] = t_9__138_ | t_9__650_;
  assign o[886] = t_9__137_ | t_9__649_;
  assign o[887] = t_9__136_ | t_9__648_;
  assign o[888] = t_9__135_ | t_9__647_;
  assign o[889] = t_9__134_ | t_9__646_;
  assign o[890] = t_9__133_ | t_9__645_;
  assign o[891] = t_9__132_ | t_9__644_;
  assign o[892] = t_9__131_ | t_9__643_;
  assign o[893] = t_9__130_ | t_9__642_;
  assign o[894] = t_9__129_ | t_9__641_;
  assign o[895] = t_9__128_ | t_9__640_;
  assign o[896] = t_9__127_ | t_9__639_;
  assign o[897] = t_9__126_ | t_9__638_;
  assign o[898] = t_9__125_ | t_9__637_;
  assign o[899] = t_9__124_ | t_9__636_;
  assign o[900] = t_9__123_ | t_9__635_;
  assign o[901] = t_9__122_ | t_9__634_;
  assign o[902] = t_9__121_ | t_9__633_;
  assign o[903] = t_9__120_ | t_9__632_;
  assign o[904] = t_9__119_ | t_9__631_;
  assign o[905] = t_9__118_ | t_9__630_;
  assign o[906] = t_9__117_ | t_9__629_;
  assign o[907] = t_9__116_ | t_9__628_;
  assign o[908] = t_9__115_ | t_9__627_;
  assign o[909] = t_9__114_ | t_9__626_;
  assign o[910] = t_9__113_ | t_9__625_;
  assign o[911] = t_9__112_ | t_9__624_;
  assign o[912] = t_9__111_ | t_9__623_;
  assign o[913] = t_9__110_ | t_9__622_;
  assign o[914] = t_9__109_ | t_9__621_;
  assign o[915] = t_9__108_ | t_9__620_;
  assign o[916] = t_9__107_ | t_9__619_;
  assign o[917] = t_9__106_ | t_9__618_;
  assign o[918] = t_9__105_ | t_9__617_;
  assign o[919] = t_9__104_ | t_9__616_;
  assign o[920] = t_9__103_ | t_9__615_;
  assign o[921] = t_9__102_ | t_9__614_;
  assign o[922] = t_9__101_ | t_9__613_;
  assign o[923] = t_9__100_ | t_9__612_;
  assign o[924] = t_9__99_ | t_9__611_;
  assign o[925] = t_9__98_ | t_9__610_;
  assign o[926] = t_9__97_ | t_9__609_;
  assign o[927] = t_9__96_ | t_9__608_;
  assign o[928] = t_9__95_ | t_9__607_;
  assign o[929] = t_9__94_ | t_9__606_;
  assign o[930] = t_9__93_ | t_9__605_;
  assign o[931] = t_9__92_ | t_9__604_;
  assign o[932] = t_9__91_ | t_9__603_;
  assign o[933] = t_9__90_ | t_9__602_;
  assign o[934] = t_9__89_ | t_9__601_;
  assign o[935] = t_9__88_ | t_9__600_;
  assign o[936] = t_9__87_ | t_9__599_;
  assign o[937] = t_9__86_ | t_9__598_;
  assign o[938] = t_9__85_ | t_9__597_;
  assign o[939] = t_9__84_ | t_9__596_;
  assign o[940] = t_9__83_ | t_9__595_;
  assign o[941] = t_9__82_ | t_9__594_;
  assign o[942] = t_9__81_ | t_9__593_;
  assign o[943] = t_9__80_ | t_9__592_;
  assign o[944] = t_9__79_ | t_9__591_;
  assign o[945] = t_9__78_ | t_9__590_;
  assign o[946] = t_9__77_ | t_9__589_;
  assign o[947] = t_9__76_ | t_9__588_;
  assign o[948] = t_9__75_ | t_9__587_;
  assign o[949] = t_9__74_ | t_9__586_;
  assign o[950] = t_9__73_ | t_9__585_;
  assign o[951] = t_9__72_ | t_9__584_;
  assign o[952] = t_9__71_ | t_9__583_;
  assign o[953] = t_9__70_ | t_9__582_;
  assign o[954] = t_9__69_ | t_9__581_;
  assign o[955] = t_9__68_ | t_9__580_;
  assign o[956] = t_9__67_ | t_9__579_;
  assign o[957] = t_9__66_ | t_9__578_;
  assign o[958] = t_9__65_ | t_9__577_;
  assign o[959] = t_9__64_ | t_9__576_;
  assign o[960] = t_9__63_ | t_9__575_;
  assign o[961] = t_9__62_ | t_9__574_;
  assign o[962] = t_9__61_ | t_9__573_;
  assign o[963] = t_9__60_ | t_9__572_;
  assign o[964] = t_9__59_ | t_9__571_;
  assign o[965] = t_9__58_ | t_9__570_;
  assign o[966] = t_9__57_ | t_9__569_;
  assign o[967] = t_9__56_ | t_9__568_;
  assign o[968] = t_9__55_ | t_9__567_;
  assign o[969] = t_9__54_ | t_9__566_;
  assign o[970] = t_9__53_ | t_9__565_;
  assign o[971] = t_9__52_ | t_9__564_;
  assign o[972] = t_9__51_ | t_9__563_;
  assign o[973] = t_9__50_ | t_9__562_;
  assign o[974] = t_9__49_ | t_9__561_;
  assign o[975] = t_9__48_ | t_9__560_;
  assign o[976] = t_9__47_ | t_9__559_;
  assign o[977] = t_9__46_ | t_9__558_;
  assign o[978] = t_9__45_ | t_9__557_;
  assign o[979] = t_9__44_ | t_9__556_;
  assign o[980] = t_9__43_ | t_9__555_;
  assign o[981] = t_9__42_ | t_9__554_;
  assign o[982] = t_9__41_ | t_9__553_;
  assign o[983] = t_9__40_ | t_9__552_;
  assign o[984] = t_9__39_ | t_9__551_;
  assign o[985] = t_9__38_ | t_9__550_;
  assign o[986] = t_9__37_ | t_9__549_;
  assign o[987] = t_9__36_ | t_9__548_;
  assign o[988] = t_9__35_ | t_9__547_;
  assign o[989] = t_9__34_ | t_9__546_;
  assign o[990] = t_9__33_ | t_9__545_;
  assign o[991] = t_9__32_ | t_9__544_;
  assign o[992] = t_9__31_ | t_9__543_;
  assign o[993] = t_9__30_ | t_9__542_;
  assign o[994] = t_9__29_ | t_9__541_;
  assign o[995] = t_9__28_ | t_9__540_;
  assign o[996] = t_9__27_ | t_9__539_;
  assign o[997] = t_9__26_ | t_9__538_;
  assign o[998] = t_9__25_ | t_9__537_;
  assign o[999] = t_9__24_ | t_9__536_;
  assign o[1000] = t_9__23_ | t_9__535_;
  assign o[1001] = t_9__22_ | t_9__534_;
  assign o[1002] = t_9__21_ | t_9__533_;
  assign o[1003] = t_9__20_ | t_9__532_;
  assign o[1004] = t_9__19_ | t_9__531_;
  assign o[1005] = t_9__18_ | t_9__530_;
  assign o[1006] = t_9__17_ | t_9__529_;
  assign o[1007] = t_9__16_ | t_9__528_;
  assign o[1008] = t_9__15_ | t_9__527_;
  assign o[1009] = t_9__14_ | t_9__526_;
  assign o[1010] = t_9__13_ | t_9__525_;
  assign o[1011] = t_9__12_ | t_9__524_;
  assign o[1012] = t_9__11_ | t_9__523_;
  assign o[1013] = t_9__10_ | t_9__522_;
  assign o[1014] = t_9__9_ | t_9__521_;
  assign o[1015] = t_9__8_ | t_9__520_;
  assign o[1016] = t_9__7_ | t_9__519_;
  assign o[1017] = t_9__6_ | t_9__518_;
  assign o[1018] = t_9__5_ | t_9__517_;
  assign o[1019] = t_9__4_ | t_9__516_;
  assign o[1020] = t_9__3_ | t_9__515_;
  assign o[1021] = t_9__2_ | t_9__514_;
  assign o[1022] = t_9__1_ | t_9__513_;
  assign o[1023] = t_9__0_ | t_9__512_;

endmodule



module bsg_priority_encode_one_hot_out_width_p1024_lo_to_hi_p1
(
  i,
  o
);

  input [1023:0] i;
  output [1023:0] o;
  wire [1023:0] o;
  wire N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,N17,N18,N19,N20,N21,
  N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,N33,N34,N35,N36,N37,N38,N39,N40,N41,
  N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,N53,N54,N55,N56,N57,N58,N59,N60,N61,
  N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,N73,N74,N75,N76,N77,N78,N79,N80,N81,
  N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,N93,N94,N95,N96,N97,N98,N99,N100,N101,
  N102,N103,N104,N105,N106,N107,N108,N109,N110,N111,N112,N113,N114,N115,N116,N117,
  N118,N119,N120,N121,N122,N123,N124,N125,N126,N127,N128,N129,N130,N131,N132,N133,
  N134,N135,N136,N137,N138,N139,N140,N141,N142,N143,N144,N145,N146,N147,N148,N149,
  N150,N151,N152,N153,N154,N155,N156,N157,N158,N159,N160,N161,N162,N163,N164,N165,
  N166,N167,N168,N169,N170,N171,N172,N173,N174,N175,N176,N177,N178,N179,N180,N181,
  N182,N183,N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,N194,N195,N196,N197,
  N198,N199,N200,N201,N202,N203,N204,N205,N206,N207,N208,N209,N210,N211,N212,N213,
  N214,N215,N216,N217,N218,N219,N220,N221,N222,N223,N224,N225,N226,N227,N228,N229,
  N230,N231,N232,N233,N234,N235,N236,N237,N238,N239,N240,N241,N242,N243,N244,N245,
  N246,N247,N248,N249,N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,N260,N261,
  N262,N263,N264,N265,N266,N267,N268,N269,N270,N271,N272,N273,N274,N275,N276,N277,
  N278,N279,N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,N290,N291,N292,N293,
  N294,N295,N296,N297,N298,N299,N300,N301,N302,N303,N304,N305,N306,N307,N308,N309,
  N310,N311,N312,N313,N314,N315,N316,N317,N318,N319,N320,N321,N322,N323,N324,N325,
  N326,N327,N328,N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,N339,N340,N341,
  N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,N354,N355,N356,N357,
  N358,N359,N360,N361,N362,N363,N364,N365,N366,N367,N368,N369,N370,N371,N372,N373,
  N374,N375,N376,N377,N378,N379,N380,N381,N382,N383,N384,N385,N386,N387,N388,N389,
  N390,N391,N392,N393,N394,N395,N396,N397,N398,N399,N400,N401,N402,N403,N404,N405,
  N406,N407,N408,N409,N410,N411,N412,N413,N414,N415,N416,N417,N418,N419,N420,N421,
  N422,N423,N424,N425,N426,N427,N428,N429,N430,N431,N432,N433,N434,N435,N436,N437,
  N438,N439,N440,N441,N442,N443,N444,N445,N446,N447,N448,N449,N450,N451,N452,N453,
  N454,N455,N456,N457,N458,N459,N460,N461,N462,N463,N464,N465,N466,N467,N468,N469,
  N470,N471,N472,N473,N474,N475,N476,N477,N478,N479,N480,N481,N482,N483,N484,N485,
  N486,N487,N488,N489,N490,N491,N492,N493,N494,N495,N496,N497,N498,N499,N500,N501,
  N502,N503,N504,N505,N506,N507,N508,N509,N510,N511,N512,N513,N514,N515,N516,N517,
  N518,N519,N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,N530,N531,N532,N533,
  N534,N535,N536,N537,N538,N539,N540,N541,N542,N543,N544,N545,N546,N547,N548,N549,
  N550,N551,N552,N553,N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,N564,N565,
  N566,N567,N568,N569,N570,N571,N572,N573,N574,N575,N576,N577,N578,N579,N580,N581,
  N582,N583,N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,N594,N595,N596,N597,
  N598,N599,N600,N601,N602,N603,N604,N605,N606,N607,N608,N609,N610,N611,N612,N613,
  N614,N615,N616,N617,N618,N619,N620,N621,N622,N623,N624,N625,N626,N627,N628,N629,
  N630,N631,N632,N633,N634,N635,N636,N637,N638,N639,N640,N641,N642,N643,N644,N645,
  N646,N647,N648,N649,N650,N651,N652,N653,N654,N655,N656,N657,N658,N659,N660,N661,
  N662,N663,N664,N665,N666,N667,N668,N669,N670,N671,N672,N673,N674,N675,N676,N677,
  N678,N679,N680,N681,N682,N683,N684,N685,N686,N687,N688,N689,N690,N691,N692,N693,
  N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,N704,N705,N706,N707,N708,N709,
  N710,N711,N712,N713,N714,N715,N716,N717,N718,N719,N720,N721,N722,N723,N724,N725,
  N726,N727,N728,N729,N730,N731,N732,N733,N734,N735,N736,N737,N738,N739,N740,N741,
  N742,N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,N754,N755,N756,N757,
  N758,N759,N760,N761,N762,N763,N764,N765,N766,N767,N768,N769,N770,N771,N772,N773,
  N774,N775,N776,N777,N778,N779,N780,N781,N782,N783,N784,N785,N786,N787,N788,N789,
  N790,N791,N792,N793,N794,N795,N796,N797,N798,N799,N800,N801,N802,N803,N804,N805,
  N806,N807,N808,N809,N810,N811,N812,N813,N814,N815,N816,N817,N818,N819,N820,N821,
  N822,N823,N824,N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,N835,N836,N837,
  N838,N839,N840,N841,N842,N843,N844,N845,N846,N847,N848,N849,N850,N851,N852,N853,
  N854,N855,N856,N857,N858,N859,N860,N861,N862,N863,N864,N865,N866,N867,N868,N869,
  N870,N871,N872,N873,N874,N875,N876,N877,N878,N879,N880,N881,N882,N883,N884,N885,
  N886,N887,N888,N889,N890,N891,N892,N893,N894,N895,N896,N897,N898,N899,N900,N901,
  N902,N903,N904,N905,N906,N907,N908,N909,N910,N911,N912,N913,N914,N915,N916,N917,
  N918,N919,N920,N921,N922,N923,N924,N925,N926,N927,N928,N929,N930,N931,N932,N933,
  N934,N935,N936,N937,N938,N939,N940,N941,N942,N943,N944,N945,N946,N947,N948,N949,
  N950,N951,N952,N953,N954,N955,N956,N957,N958,N959,N960,N961,N962,N963,N964,N965,
  N966,N967,N968,N969,N970,N971,N972,N973,N974,N975,N976,N977,N978,N979,N980,N981,
  N982,N983,N984,N985,N986,N987,N988,N989,N990,N991,N992,N993,N994,N995,N996,N997,
  N998,N999,N1000,N1001,N1002,N1003,N1004,N1005,N1006,N1007,N1008,N1009,N1010,
  N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,N1019,N1020,N1021,N1022;
  wire [1023:1] scan_lo;

  bsg_scan_width_p1024_or_p1_lo_to_hi_p1
  genblk1_scan
  (
    .i(i),
    .o({ scan_lo, o[0:0] })
  );

  assign o[1023] = scan_lo[1023] & N0;
  assign N0 = ~scan_lo[1022];
  assign o[1022] = scan_lo[1022] & N1;
  assign N1 = ~scan_lo[1021];
  assign o[1021] = scan_lo[1021] & N2;
  assign N2 = ~scan_lo[1020];
  assign o[1020] = scan_lo[1020] & N3;
  assign N3 = ~scan_lo[1019];
  assign o[1019] = scan_lo[1019] & N4;
  assign N4 = ~scan_lo[1018];
  assign o[1018] = scan_lo[1018] & N5;
  assign N5 = ~scan_lo[1017];
  assign o[1017] = scan_lo[1017] & N6;
  assign N6 = ~scan_lo[1016];
  assign o[1016] = scan_lo[1016] & N7;
  assign N7 = ~scan_lo[1015];
  assign o[1015] = scan_lo[1015] & N8;
  assign N8 = ~scan_lo[1014];
  assign o[1014] = scan_lo[1014] & N9;
  assign N9 = ~scan_lo[1013];
  assign o[1013] = scan_lo[1013] & N10;
  assign N10 = ~scan_lo[1012];
  assign o[1012] = scan_lo[1012] & N11;
  assign N11 = ~scan_lo[1011];
  assign o[1011] = scan_lo[1011] & N12;
  assign N12 = ~scan_lo[1010];
  assign o[1010] = scan_lo[1010] & N13;
  assign N13 = ~scan_lo[1009];
  assign o[1009] = scan_lo[1009] & N14;
  assign N14 = ~scan_lo[1008];
  assign o[1008] = scan_lo[1008] & N15;
  assign N15 = ~scan_lo[1007];
  assign o[1007] = scan_lo[1007] & N16;
  assign N16 = ~scan_lo[1006];
  assign o[1006] = scan_lo[1006] & N17;
  assign N17 = ~scan_lo[1005];
  assign o[1005] = scan_lo[1005] & N18;
  assign N18 = ~scan_lo[1004];
  assign o[1004] = scan_lo[1004] & N19;
  assign N19 = ~scan_lo[1003];
  assign o[1003] = scan_lo[1003] & N20;
  assign N20 = ~scan_lo[1002];
  assign o[1002] = scan_lo[1002] & N21;
  assign N21 = ~scan_lo[1001];
  assign o[1001] = scan_lo[1001] & N22;
  assign N22 = ~scan_lo[1000];
  assign o[1000] = scan_lo[1000] & N23;
  assign N23 = ~scan_lo[999];
  assign o[999] = scan_lo[999] & N24;
  assign N24 = ~scan_lo[998];
  assign o[998] = scan_lo[998] & N25;
  assign N25 = ~scan_lo[997];
  assign o[997] = scan_lo[997] & N26;
  assign N26 = ~scan_lo[996];
  assign o[996] = scan_lo[996] & N27;
  assign N27 = ~scan_lo[995];
  assign o[995] = scan_lo[995] & N28;
  assign N28 = ~scan_lo[994];
  assign o[994] = scan_lo[994] & N29;
  assign N29 = ~scan_lo[993];
  assign o[993] = scan_lo[993] & N30;
  assign N30 = ~scan_lo[992];
  assign o[992] = scan_lo[992] & N31;
  assign N31 = ~scan_lo[991];
  assign o[991] = scan_lo[991] & N32;
  assign N32 = ~scan_lo[990];
  assign o[990] = scan_lo[990] & N33;
  assign N33 = ~scan_lo[989];
  assign o[989] = scan_lo[989] & N34;
  assign N34 = ~scan_lo[988];
  assign o[988] = scan_lo[988] & N35;
  assign N35 = ~scan_lo[987];
  assign o[987] = scan_lo[987] & N36;
  assign N36 = ~scan_lo[986];
  assign o[986] = scan_lo[986] & N37;
  assign N37 = ~scan_lo[985];
  assign o[985] = scan_lo[985] & N38;
  assign N38 = ~scan_lo[984];
  assign o[984] = scan_lo[984] & N39;
  assign N39 = ~scan_lo[983];
  assign o[983] = scan_lo[983] & N40;
  assign N40 = ~scan_lo[982];
  assign o[982] = scan_lo[982] & N41;
  assign N41 = ~scan_lo[981];
  assign o[981] = scan_lo[981] & N42;
  assign N42 = ~scan_lo[980];
  assign o[980] = scan_lo[980] & N43;
  assign N43 = ~scan_lo[979];
  assign o[979] = scan_lo[979] & N44;
  assign N44 = ~scan_lo[978];
  assign o[978] = scan_lo[978] & N45;
  assign N45 = ~scan_lo[977];
  assign o[977] = scan_lo[977] & N46;
  assign N46 = ~scan_lo[976];
  assign o[976] = scan_lo[976] & N47;
  assign N47 = ~scan_lo[975];
  assign o[975] = scan_lo[975] & N48;
  assign N48 = ~scan_lo[974];
  assign o[974] = scan_lo[974] & N49;
  assign N49 = ~scan_lo[973];
  assign o[973] = scan_lo[973] & N50;
  assign N50 = ~scan_lo[972];
  assign o[972] = scan_lo[972] & N51;
  assign N51 = ~scan_lo[971];
  assign o[971] = scan_lo[971] & N52;
  assign N52 = ~scan_lo[970];
  assign o[970] = scan_lo[970] & N53;
  assign N53 = ~scan_lo[969];
  assign o[969] = scan_lo[969] & N54;
  assign N54 = ~scan_lo[968];
  assign o[968] = scan_lo[968] & N55;
  assign N55 = ~scan_lo[967];
  assign o[967] = scan_lo[967] & N56;
  assign N56 = ~scan_lo[966];
  assign o[966] = scan_lo[966] & N57;
  assign N57 = ~scan_lo[965];
  assign o[965] = scan_lo[965] & N58;
  assign N58 = ~scan_lo[964];
  assign o[964] = scan_lo[964] & N59;
  assign N59 = ~scan_lo[963];
  assign o[963] = scan_lo[963] & N60;
  assign N60 = ~scan_lo[962];
  assign o[962] = scan_lo[962] & N61;
  assign N61 = ~scan_lo[961];
  assign o[961] = scan_lo[961] & N62;
  assign N62 = ~scan_lo[960];
  assign o[960] = scan_lo[960] & N63;
  assign N63 = ~scan_lo[959];
  assign o[959] = scan_lo[959] & N64;
  assign N64 = ~scan_lo[958];
  assign o[958] = scan_lo[958] & N65;
  assign N65 = ~scan_lo[957];
  assign o[957] = scan_lo[957] & N66;
  assign N66 = ~scan_lo[956];
  assign o[956] = scan_lo[956] & N67;
  assign N67 = ~scan_lo[955];
  assign o[955] = scan_lo[955] & N68;
  assign N68 = ~scan_lo[954];
  assign o[954] = scan_lo[954] & N69;
  assign N69 = ~scan_lo[953];
  assign o[953] = scan_lo[953] & N70;
  assign N70 = ~scan_lo[952];
  assign o[952] = scan_lo[952] & N71;
  assign N71 = ~scan_lo[951];
  assign o[951] = scan_lo[951] & N72;
  assign N72 = ~scan_lo[950];
  assign o[950] = scan_lo[950] & N73;
  assign N73 = ~scan_lo[949];
  assign o[949] = scan_lo[949] & N74;
  assign N74 = ~scan_lo[948];
  assign o[948] = scan_lo[948] & N75;
  assign N75 = ~scan_lo[947];
  assign o[947] = scan_lo[947] & N76;
  assign N76 = ~scan_lo[946];
  assign o[946] = scan_lo[946] & N77;
  assign N77 = ~scan_lo[945];
  assign o[945] = scan_lo[945] & N78;
  assign N78 = ~scan_lo[944];
  assign o[944] = scan_lo[944] & N79;
  assign N79 = ~scan_lo[943];
  assign o[943] = scan_lo[943] & N80;
  assign N80 = ~scan_lo[942];
  assign o[942] = scan_lo[942] & N81;
  assign N81 = ~scan_lo[941];
  assign o[941] = scan_lo[941] & N82;
  assign N82 = ~scan_lo[940];
  assign o[940] = scan_lo[940] & N83;
  assign N83 = ~scan_lo[939];
  assign o[939] = scan_lo[939] & N84;
  assign N84 = ~scan_lo[938];
  assign o[938] = scan_lo[938] & N85;
  assign N85 = ~scan_lo[937];
  assign o[937] = scan_lo[937] & N86;
  assign N86 = ~scan_lo[936];
  assign o[936] = scan_lo[936] & N87;
  assign N87 = ~scan_lo[935];
  assign o[935] = scan_lo[935] & N88;
  assign N88 = ~scan_lo[934];
  assign o[934] = scan_lo[934] & N89;
  assign N89 = ~scan_lo[933];
  assign o[933] = scan_lo[933] & N90;
  assign N90 = ~scan_lo[932];
  assign o[932] = scan_lo[932] & N91;
  assign N91 = ~scan_lo[931];
  assign o[931] = scan_lo[931] & N92;
  assign N92 = ~scan_lo[930];
  assign o[930] = scan_lo[930] & N93;
  assign N93 = ~scan_lo[929];
  assign o[929] = scan_lo[929] & N94;
  assign N94 = ~scan_lo[928];
  assign o[928] = scan_lo[928] & N95;
  assign N95 = ~scan_lo[927];
  assign o[927] = scan_lo[927] & N96;
  assign N96 = ~scan_lo[926];
  assign o[926] = scan_lo[926] & N97;
  assign N97 = ~scan_lo[925];
  assign o[925] = scan_lo[925] & N98;
  assign N98 = ~scan_lo[924];
  assign o[924] = scan_lo[924] & N99;
  assign N99 = ~scan_lo[923];
  assign o[923] = scan_lo[923] & N100;
  assign N100 = ~scan_lo[922];
  assign o[922] = scan_lo[922] & N101;
  assign N101 = ~scan_lo[921];
  assign o[921] = scan_lo[921] & N102;
  assign N102 = ~scan_lo[920];
  assign o[920] = scan_lo[920] & N103;
  assign N103 = ~scan_lo[919];
  assign o[919] = scan_lo[919] & N104;
  assign N104 = ~scan_lo[918];
  assign o[918] = scan_lo[918] & N105;
  assign N105 = ~scan_lo[917];
  assign o[917] = scan_lo[917] & N106;
  assign N106 = ~scan_lo[916];
  assign o[916] = scan_lo[916] & N107;
  assign N107 = ~scan_lo[915];
  assign o[915] = scan_lo[915] & N108;
  assign N108 = ~scan_lo[914];
  assign o[914] = scan_lo[914] & N109;
  assign N109 = ~scan_lo[913];
  assign o[913] = scan_lo[913] & N110;
  assign N110 = ~scan_lo[912];
  assign o[912] = scan_lo[912] & N111;
  assign N111 = ~scan_lo[911];
  assign o[911] = scan_lo[911] & N112;
  assign N112 = ~scan_lo[910];
  assign o[910] = scan_lo[910] & N113;
  assign N113 = ~scan_lo[909];
  assign o[909] = scan_lo[909] & N114;
  assign N114 = ~scan_lo[908];
  assign o[908] = scan_lo[908] & N115;
  assign N115 = ~scan_lo[907];
  assign o[907] = scan_lo[907] & N116;
  assign N116 = ~scan_lo[906];
  assign o[906] = scan_lo[906] & N117;
  assign N117 = ~scan_lo[905];
  assign o[905] = scan_lo[905] & N118;
  assign N118 = ~scan_lo[904];
  assign o[904] = scan_lo[904] & N119;
  assign N119 = ~scan_lo[903];
  assign o[903] = scan_lo[903] & N120;
  assign N120 = ~scan_lo[902];
  assign o[902] = scan_lo[902] & N121;
  assign N121 = ~scan_lo[901];
  assign o[901] = scan_lo[901] & N122;
  assign N122 = ~scan_lo[900];
  assign o[900] = scan_lo[900] & N123;
  assign N123 = ~scan_lo[899];
  assign o[899] = scan_lo[899] & N124;
  assign N124 = ~scan_lo[898];
  assign o[898] = scan_lo[898] & N125;
  assign N125 = ~scan_lo[897];
  assign o[897] = scan_lo[897] & N126;
  assign N126 = ~scan_lo[896];
  assign o[896] = scan_lo[896] & N127;
  assign N127 = ~scan_lo[895];
  assign o[895] = scan_lo[895] & N128;
  assign N128 = ~scan_lo[894];
  assign o[894] = scan_lo[894] & N129;
  assign N129 = ~scan_lo[893];
  assign o[893] = scan_lo[893] & N130;
  assign N130 = ~scan_lo[892];
  assign o[892] = scan_lo[892] & N131;
  assign N131 = ~scan_lo[891];
  assign o[891] = scan_lo[891] & N132;
  assign N132 = ~scan_lo[890];
  assign o[890] = scan_lo[890] & N133;
  assign N133 = ~scan_lo[889];
  assign o[889] = scan_lo[889] & N134;
  assign N134 = ~scan_lo[888];
  assign o[888] = scan_lo[888] & N135;
  assign N135 = ~scan_lo[887];
  assign o[887] = scan_lo[887] & N136;
  assign N136 = ~scan_lo[886];
  assign o[886] = scan_lo[886] & N137;
  assign N137 = ~scan_lo[885];
  assign o[885] = scan_lo[885] & N138;
  assign N138 = ~scan_lo[884];
  assign o[884] = scan_lo[884] & N139;
  assign N139 = ~scan_lo[883];
  assign o[883] = scan_lo[883] & N140;
  assign N140 = ~scan_lo[882];
  assign o[882] = scan_lo[882] & N141;
  assign N141 = ~scan_lo[881];
  assign o[881] = scan_lo[881] & N142;
  assign N142 = ~scan_lo[880];
  assign o[880] = scan_lo[880] & N143;
  assign N143 = ~scan_lo[879];
  assign o[879] = scan_lo[879] & N144;
  assign N144 = ~scan_lo[878];
  assign o[878] = scan_lo[878] & N145;
  assign N145 = ~scan_lo[877];
  assign o[877] = scan_lo[877] & N146;
  assign N146 = ~scan_lo[876];
  assign o[876] = scan_lo[876] & N147;
  assign N147 = ~scan_lo[875];
  assign o[875] = scan_lo[875] & N148;
  assign N148 = ~scan_lo[874];
  assign o[874] = scan_lo[874] & N149;
  assign N149 = ~scan_lo[873];
  assign o[873] = scan_lo[873] & N150;
  assign N150 = ~scan_lo[872];
  assign o[872] = scan_lo[872] & N151;
  assign N151 = ~scan_lo[871];
  assign o[871] = scan_lo[871] & N152;
  assign N152 = ~scan_lo[870];
  assign o[870] = scan_lo[870] & N153;
  assign N153 = ~scan_lo[869];
  assign o[869] = scan_lo[869] & N154;
  assign N154 = ~scan_lo[868];
  assign o[868] = scan_lo[868] & N155;
  assign N155 = ~scan_lo[867];
  assign o[867] = scan_lo[867] & N156;
  assign N156 = ~scan_lo[866];
  assign o[866] = scan_lo[866] & N157;
  assign N157 = ~scan_lo[865];
  assign o[865] = scan_lo[865] & N158;
  assign N158 = ~scan_lo[864];
  assign o[864] = scan_lo[864] & N159;
  assign N159 = ~scan_lo[863];
  assign o[863] = scan_lo[863] & N160;
  assign N160 = ~scan_lo[862];
  assign o[862] = scan_lo[862] & N161;
  assign N161 = ~scan_lo[861];
  assign o[861] = scan_lo[861] & N162;
  assign N162 = ~scan_lo[860];
  assign o[860] = scan_lo[860] & N163;
  assign N163 = ~scan_lo[859];
  assign o[859] = scan_lo[859] & N164;
  assign N164 = ~scan_lo[858];
  assign o[858] = scan_lo[858] & N165;
  assign N165 = ~scan_lo[857];
  assign o[857] = scan_lo[857] & N166;
  assign N166 = ~scan_lo[856];
  assign o[856] = scan_lo[856] & N167;
  assign N167 = ~scan_lo[855];
  assign o[855] = scan_lo[855] & N168;
  assign N168 = ~scan_lo[854];
  assign o[854] = scan_lo[854] & N169;
  assign N169 = ~scan_lo[853];
  assign o[853] = scan_lo[853] & N170;
  assign N170 = ~scan_lo[852];
  assign o[852] = scan_lo[852] & N171;
  assign N171 = ~scan_lo[851];
  assign o[851] = scan_lo[851] & N172;
  assign N172 = ~scan_lo[850];
  assign o[850] = scan_lo[850] & N173;
  assign N173 = ~scan_lo[849];
  assign o[849] = scan_lo[849] & N174;
  assign N174 = ~scan_lo[848];
  assign o[848] = scan_lo[848] & N175;
  assign N175 = ~scan_lo[847];
  assign o[847] = scan_lo[847] & N176;
  assign N176 = ~scan_lo[846];
  assign o[846] = scan_lo[846] & N177;
  assign N177 = ~scan_lo[845];
  assign o[845] = scan_lo[845] & N178;
  assign N178 = ~scan_lo[844];
  assign o[844] = scan_lo[844] & N179;
  assign N179 = ~scan_lo[843];
  assign o[843] = scan_lo[843] & N180;
  assign N180 = ~scan_lo[842];
  assign o[842] = scan_lo[842] & N181;
  assign N181 = ~scan_lo[841];
  assign o[841] = scan_lo[841] & N182;
  assign N182 = ~scan_lo[840];
  assign o[840] = scan_lo[840] & N183;
  assign N183 = ~scan_lo[839];
  assign o[839] = scan_lo[839] & N184;
  assign N184 = ~scan_lo[838];
  assign o[838] = scan_lo[838] & N185;
  assign N185 = ~scan_lo[837];
  assign o[837] = scan_lo[837] & N186;
  assign N186 = ~scan_lo[836];
  assign o[836] = scan_lo[836] & N187;
  assign N187 = ~scan_lo[835];
  assign o[835] = scan_lo[835] & N188;
  assign N188 = ~scan_lo[834];
  assign o[834] = scan_lo[834] & N189;
  assign N189 = ~scan_lo[833];
  assign o[833] = scan_lo[833] & N190;
  assign N190 = ~scan_lo[832];
  assign o[832] = scan_lo[832] & N191;
  assign N191 = ~scan_lo[831];
  assign o[831] = scan_lo[831] & N192;
  assign N192 = ~scan_lo[830];
  assign o[830] = scan_lo[830] & N193;
  assign N193 = ~scan_lo[829];
  assign o[829] = scan_lo[829] & N194;
  assign N194 = ~scan_lo[828];
  assign o[828] = scan_lo[828] & N195;
  assign N195 = ~scan_lo[827];
  assign o[827] = scan_lo[827] & N196;
  assign N196 = ~scan_lo[826];
  assign o[826] = scan_lo[826] & N197;
  assign N197 = ~scan_lo[825];
  assign o[825] = scan_lo[825] & N198;
  assign N198 = ~scan_lo[824];
  assign o[824] = scan_lo[824] & N199;
  assign N199 = ~scan_lo[823];
  assign o[823] = scan_lo[823] & N200;
  assign N200 = ~scan_lo[822];
  assign o[822] = scan_lo[822] & N201;
  assign N201 = ~scan_lo[821];
  assign o[821] = scan_lo[821] & N202;
  assign N202 = ~scan_lo[820];
  assign o[820] = scan_lo[820] & N203;
  assign N203 = ~scan_lo[819];
  assign o[819] = scan_lo[819] & N204;
  assign N204 = ~scan_lo[818];
  assign o[818] = scan_lo[818] & N205;
  assign N205 = ~scan_lo[817];
  assign o[817] = scan_lo[817] & N206;
  assign N206 = ~scan_lo[816];
  assign o[816] = scan_lo[816] & N207;
  assign N207 = ~scan_lo[815];
  assign o[815] = scan_lo[815] & N208;
  assign N208 = ~scan_lo[814];
  assign o[814] = scan_lo[814] & N209;
  assign N209 = ~scan_lo[813];
  assign o[813] = scan_lo[813] & N210;
  assign N210 = ~scan_lo[812];
  assign o[812] = scan_lo[812] & N211;
  assign N211 = ~scan_lo[811];
  assign o[811] = scan_lo[811] & N212;
  assign N212 = ~scan_lo[810];
  assign o[810] = scan_lo[810] & N213;
  assign N213 = ~scan_lo[809];
  assign o[809] = scan_lo[809] & N214;
  assign N214 = ~scan_lo[808];
  assign o[808] = scan_lo[808] & N215;
  assign N215 = ~scan_lo[807];
  assign o[807] = scan_lo[807] & N216;
  assign N216 = ~scan_lo[806];
  assign o[806] = scan_lo[806] & N217;
  assign N217 = ~scan_lo[805];
  assign o[805] = scan_lo[805] & N218;
  assign N218 = ~scan_lo[804];
  assign o[804] = scan_lo[804] & N219;
  assign N219 = ~scan_lo[803];
  assign o[803] = scan_lo[803] & N220;
  assign N220 = ~scan_lo[802];
  assign o[802] = scan_lo[802] & N221;
  assign N221 = ~scan_lo[801];
  assign o[801] = scan_lo[801] & N222;
  assign N222 = ~scan_lo[800];
  assign o[800] = scan_lo[800] & N223;
  assign N223 = ~scan_lo[799];
  assign o[799] = scan_lo[799] & N224;
  assign N224 = ~scan_lo[798];
  assign o[798] = scan_lo[798] & N225;
  assign N225 = ~scan_lo[797];
  assign o[797] = scan_lo[797] & N226;
  assign N226 = ~scan_lo[796];
  assign o[796] = scan_lo[796] & N227;
  assign N227 = ~scan_lo[795];
  assign o[795] = scan_lo[795] & N228;
  assign N228 = ~scan_lo[794];
  assign o[794] = scan_lo[794] & N229;
  assign N229 = ~scan_lo[793];
  assign o[793] = scan_lo[793] & N230;
  assign N230 = ~scan_lo[792];
  assign o[792] = scan_lo[792] & N231;
  assign N231 = ~scan_lo[791];
  assign o[791] = scan_lo[791] & N232;
  assign N232 = ~scan_lo[790];
  assign o[790] = scan_lo[790] & N233;
  assign N233 = ~scan_lo[789];
  assign o[789] = scan_lo[789] & N234;
  assign N234 = ~scan_lo[788];
  assign o[788] = scan_lo[788] & N235;
  assign N235 = ~scan_lo[787];
  assign o[787] = scan_lo[787] & N236;
  assign N236 = ~scan_lo[786];
  assign o[786] = scan_lo[786] & N237;
  assign N237 = ~scan_lo[785];
  assign o[785] = scan_lo[785] & N238;
  assign N238 = ~scan_lo[784];
  assign o[784] = scan_lo[784] & N239;
  assign N239 = ~scan_lo[783];
  assign o[783] = scan_lo[783] & N240;
  assign N240 = ~scan_lo[782];
  assign o[782] = scan_lo[782] & N241;
  assign N241 = ~scan_lo[781];
  assign o[781] = scan_lo[781] & N242;
  assign N242 = ~scan_lo[780];
  assign o[780] = scan_lo[780] & N243;
  assign N243 = ~scan_lo[779];
  assign o[779] = scan_lo[779] & N244;
  assign N244 = ~scan_lo[778];
  assign o[778] = scan_lo[778] & N245;
  assign N245 = ~scan_lo[777];
  assign o[777] = scan_lo[777] & N246;
  assign N246 = ~scan_lo[776];
  assign o[776] = scan_lo[776] & N247;
  assign N247 = ~scan_lo[775];
  assign o[775] = scan_lo[775] & N248;
  assign N248 = ~scan_lo[774];
  assign o[774] = scan_lo[774] & N249;
  assign N249 = ~scan_lo[773];
  assign o[773] = scan_lo[773] & N250;
  assign N250 = ~scan_lo[772];
  assign o[772] = scan_lo[772] & N251;
  assign N251 = ~scan_lo[771];
  assign o[771] = scan_lo[771] & N252;
  assign N252 = ~scan_lo[770];
  assign o[770] = scan_lo[770] & N253;
  assign N253 = ~scan_lo[769];
  assign o[769] = scan_lo[769] & N254;
  assign N254 = ~scan_lo[768];
  assign o[768] = scan_lo[768] & N255;
  assign N255 = ~scan_lo[767];
  assign o[767] = scan_lo[767] & N256;
  assign N256 = ~scan_lo[766];
  assign o[766] = scan_lo[766] & N257;
  assign N257 = ~scan_lo[765];
  assign o[765] = scan_lo[765] & N258;
  assign N258 = ~scan_lo[764];
  assign o[764] = scan_lo[764] & N259;
  assign N259 = ~scan_lo[763];
  assign o[763] = scan_lo[763] & N260;
  assign N260 = ~scan_lo[762];
  assign o[762] = scan_lo[762] & N261;
  assign N261 = ~scan_lo[761];
  assign o[761] = scan_lo[761] & N262;
  assign N262 = ~scan_lo[760];
  assign o[760] = scan_lo[760] & N263;
  assign N263 = ~scan_lo[759];
  assign o[759] = scan_lo[759] & N264;
  assign N264 = ~scan_lo[758];
  assign o[758] = scan_lo[758] & N265;
  assign N265 = ~scan_lo[757];
  assign o[757] = scan_lo[757] & N266;
  assign N266 = ~scan_lo[756];
  assign o[756] = scan_lo[756] & N267;
  assign N267 = ~scan_lo[755];
  assign o[755] = scan_lo[755] & N268;
  assign N268 = ~scan_lo[754];
  assign o[754] = scan_lo[754] & N269;
  assign N269 = ~scan_lo[753];
  assign o[753] = scan_lo[753] & N270;
  assign N270 = ~scan_lo[752];
  assign o[752] = scan_lo[752] & N271;
  assign N271 = ~scan_lo[751];
  assign o[751] = scan_lo[751] & N272;
  assign N272 = ~scan_lo[750];
  assign o[750] = scan_lo[750] & N273;
  assign N273 = ~scan_lo[749];
  assign o[749] = scan_lo[749] & N274;
  assign N274 = ~scan_lo[748];
  assign o[748] = scan_lo[748] & N275;
  assign N275 = ~scan_lo[747];
  assign o[747] = scan_lo[747] & N276;
  assign N276 = ~scan_lo[746];
  assign o[746] = scan_lo[746] & N277;
  assign N277 = ~scan_lo[745];
  assign o[745] = scan_lo[745] & N278;
  assign N278 = ~scan_lo[744];
  assign o[744] = scan_lo[744] & N279;
  assign N279 = ~scan_lo[743];
  assign o[743] = scan_lo[743] & N280;
  assign N280 = ~scan_lo[742];
  assign o[742] = scan_lo[742] & N281;
  assign N281 = ~scan_lo[741];
  assign o[741] = scan_lo[741] & N282;
  assign N282 = ~scan_lo[740];
  assign o[740] = scan_lo[740] & N283;
  assign N283 = ~scan_lo[739];
  assign o[739] = scan_lo[739] & N284;
  assign N284 = ~scan_lo[738];
  assign o[738] = scan_lo[738] & N285;
  assign N285 = ~scan_lo[737];
  assign o[737] = scan_lo[737] & N286;
  assign N286 = ~scan_lo[736];
  assign o[736] = scan_lo[736] & N287;
  assign N287 = ~scan_lo[735];
  assign o[735] = scan_lo[735] & N288;
  assign N288 = ~scan_lo[734];
  assign o[734] = scan_lo[734] & N289;
  assign N289 = ~scan_lo[733];
  assign o[733] = scan_lo[733] & N290;
  assign N290 = ~scan_lo[732];
  assign o[732] = scan_lo[732] & N291;
  assign N291 = ~scan_lo[731];
  assign o[731] = scan_lo[731] & N292;
  assign N292 = ~scan_lo[730];
  assign o[730] = scan_lo[730] & N293;
  assign N293 = ~scan_lo[729];
  assign o[729] = scan_lo[729] & N294;
  assign N294 = ~scan_lo[728];
  assign o[728] = scan_lo[728] & N295;
  assign N295 = ~scan_lo[727];
  assign o[727] = scan_lo[727] & N296;
  assign N296 = ~scan_lo[726];
  assign o[726] = scan_lo[726] & N297;
  assign N297 = ~scan_lo[725];
  assign o[725] = scan_lo[725] & N298;
  assign N298 = ~scan_lo[724];
  assign o[724] = scan_lo[724] & N299;
  assign N299 = ~scan_lo[723];
  assign o[723] = scan_lo[723] & N300;
  assign N300 = ~scan_lo[722];
  assign o[722] = scan_lo[722] & N301;
  assign N301 = ~scan_lo[721];
  assign o[721] = scan_lo[721] & N302;
  assign N302 = ~scan_lo[720];
  assign o[720] = scan_lo[720] & N303;
  assign N303 = ~scan_lo[719];
  assign o[719] = scan_lo[719] & N304;
  assign N304 = ~scan_lo[718];
  assign o[718] = scan_lo[718] & N305;
  assign N305 = ~scan_lo[717];
  assign o[717] = scan_lo[717] & N306;
  assign N306 = ~scan_lo[716];
  assign o[716] = scan_lo[716] & N307;
  assign N307 = ~scan_lo[715];
  assign o[715] = scan_lo[715] & N308;
  assign N308 = ~scan_lo[714];
  assign o[714] = scan_lo[714] & N309;
  assign N309 = ~scan_lo[713];
  assign o[713] = scan_lo[713] & N310;
  assign N310 = ~scan_lo[712];
  assign o[712] = scan_lo[712] & N311;
  assign N311 = ~scan_lo[711];
  assign o[711] = scan_lo[711] & N312;
  assign N312 = ~scan_lo[710];
  assign o[710] = scan_lo[710] & N313;
  assign N313 = ~scan_lo[709];
  assign o[709] = scan_lo[709] & N314;
  assign N314 = ~scan_lo[708];
  assign o[708] = scan_lo[708] & N315;
  assign N315 = ~scan_lo[707];
  assign o[707] = scan_lo[707] & N316;
  assign N316 = ~scan_lo[706];
  assign o[706] = scan_lo[706] & N317;
  assign N317 = ~scan_lo[705];
  assign o[705] = scan_lo[705] & N318;
  assign N318 = ~scan_lo[704];
  assign o[704] = scan_lo[704] & N319;
  assign N319 = ~scan_lo[703];
  assign o[703] = scan_lo[703] & N320;
  assign N320 = ~scan_lo[702];
  assign o[702] = scan_lo[702] & N321;
  assign N321 = ~scan_lo[701];
  assign o[701] = scan_lo[701] & N322;
  assign N322 = ~scan_lo[700];
  assign o[700] = scan_lo[700] & N323;
  assign N323 = ~scan_lo[699];
  assign o[699] = scan_lo[699] & N324;
  assign N324 = ~scan_lo[698];
  assign o[698] = scan_lo[698] & N325;
  assign N325 = ~scan_lo[697];
  assign o[697] = scan_lo[697] & N326;
  assign N326 = ~scan_lo[696];
  assign o[696] = scan_lo[696] & N327;
  assign N327 = ~scan_lo[695];
  assign o[695] = scan_lo[695] & N328;
  assign N328 = ~scan_lo[694];
  assign o[694] = scan_lo[694] & N329;
  assign N329 = ~scan_lo[693];
  assign o[693] = scan_lo[693] & N330;
  assign N330 = ~scan_lo[692];
  assign o[692] = scan_lo[692] & N331;
  assign N331 = ~scan_lo[691];
  assign o[691] = scan_lo[691] & N332;
  assign N332 = ~scan_lo[690];
  assign o[690] = scan_lo[690] & N333;
  assign N333 = ~scan_lo[689];
  assign o[689] = scan_lo[689] & N334;
  assign N334 = ~scan_lo[688];
  assign o[688] = scan_lo[688] & N335;
  assign N335 = ~scan_lo[687];
  assign o[687] = scan_lo[687] & N336;
  assign N336 = ~scan_lo[686];
  assign o[686] = scan_lo[686] & N337;
  assign N337 = ~scan_lo[685];
  assign o[685] = scan_lo[685] & N338;
  assign N338 = ~scan_lo[684];
  assign o[684] = scan_lo[684] & N339;
  assign N339 = ~scan_lo[683];
  assign o[683] = scan_lo[683] & N340;
  assign N340 = ~scan_lo[682];
  assign o[682] = scan_lo[682] & N341;
  assign N341 = ~scan_lo[681];
  assign o[681] = scan_lo[681] & N342;
  assign N342 = ~scan_lo[680];
  assign o[680] = scan_lo[680] & N343;
  assign N343 = ~scan_lo[679];
  assign o[679] = scan_lo[679] & N344;
  assign N344 = ~scan_lo[678];
  assign o[678] = scan_lo[678] & N345;
  assign N345 = ~scan_lo[677];
  assign o[677] = scan_lo[677] & N346;
  assign N346 = ~scan_lo[676];
  assign o[676] = scan_lo[676] & N347;
  assign N347 = ~scan_lo[675];
  assign o[675] = scan_lo[675] & N348;
  assign N348 = ~scan_lo[674];
  assign o[674] = scan_lo[674] & N349;
  assign N349 = ~scan_lo[673];
  assign o[673] = scan_lo[673] & N350;
  assign N350 = ~scan_lo[672];
  assign o[672] = scan_lo[672] & N351;
  assign N351 = ~scan_lo[671];
  assign o[671] = scan_lo[671] & N352;
  assign N352 = ~scan_lo[670];
  assign o[670] = scan_lo[670] & N353;
  assign N353 = ~scan_lo[669];
  assign o[669] = scan_lo[669] & N354;
  assign N354 = ~scan_lo[668];
  assign o[668] = scan_lo[668] & N355;
  assign N355 = ~scan_lo[667];
  assign o[667] = scan_lo[667] & N356;
  assign N356 = ~scan_lo[666];
  assign o[666] = scan_lo[666] & N357;
  assign N357 = ~scan_lo[665];
  assign o[665] = scan_lo[665] & N358;
  assign N358 = ~scan_lo[664];
  assign o[664] = scan_lo[664] & N359;
  assign N359 = ~scan_lo[663];
  assign o[663] = scan_lo[663] & N360;
  assign N360 = ~scan_lo[662];
  assign o[662] = scan_lo[662] & N361;
  assign N361 = ~scan_lo[661];
  assign o[661] = scan_lo[661] & N362;
  assign N362 = ~scan_lo[660];
  assign o[660] = scan_lo[660] & N363;
  assign N363 = ~scan_lo[659];
  assign o[659] = scan_lo[659] & N364;
  assign N364 = ~scan_lo[658];
  assign o[658] = scan_lo[658] & N365;
  assign N365 = ~scan_lo[657];
  assign o[657] = scan_lo[657] & N366;
  assign N366 = ~scan_lo[656];
  assign o[656] = scan_lo[656] & N367;
  assign N367 = ~scan_lo[655];
  assign o[655] = scan_lo[655] & N368;
  assign N368 = ~scan_lo[654];
  assign o[654] = scan_lo[654] & N369;
  assign N369 = ~scan_lo[653];
  assign o[653] = scan_lo[653] & N370;
  assign N370 = ~scan_lo[652];
  assign o[652] = scan_lo[652] & N371;
  assign N371 = ~scan_lo[651];
  assign o[651] = scan_lo[651] & N372;
  assign N372 = ~scan_lo[650];
  assign o[650] = scan_lo[650] & N373;
  assign N373 = ~scan_lo[649];
  assign o[649] = scan_lo[649] & N374;
  assign N374 = ~scan_lo[648];
  assign o[648] = scan_lo[648] & N375;
  assign N375 = ~scan_lo[647];
  assign o[647] = scan_lo[647] & N376;
  assign N376 = ~scan_lo[646];
  assign o[646] = scan_lo[646] & N377;
  assign N377 = ~scan_lo[645];
  assign o[645] = scan_lo[645] & N378;
  assign N378 = ~scan_lo[644];
  assign o[644] = scan_lo[644] & N379;
  assign N379 = ~scan_lo[643];
  assign o[643] = scan_lo[643] & N380;
  assign N380 = ~scan_lo[642];
  assign o[642] = scan_lo[642] & N381;
  assign N381 = ~scan_lo[641];
  assign o[641] = scan_lo[641] & N382;
  assign N382 = ~scan_lo[640];
  assign o[640] = scan_lo[640] & N383;
  assign N383 = ~scan_lo[639];
  assign o[639] = scan_lo[639] & N384;
  assign N384 = ~scan_lo[638];
  assign o[638] = scan_lo[638] & N385;
  assign N385 = ~scan_lo[637];
  assign o[637] = scan_lo[637] & N386;
  assign N386 = ~scan_lo[636];
  assign o[636] = scan_lo[636] & N387;
  assign N387 = ~scan_lo[635];
  assign o[635] = scan_lo[635] & N388;
  assign N388 = ~scan_lo[634];
  assign o[634] = scan_lo[634] & N389;
  assign N389 = ~scan_lo[633];
  assign o[633] = scan_lo[633] & N390;
  assign N390 = ~scan_lo[632];
  assign o[632] = scan_lo[632] & N391;
  assign N391 = ~scan_lo[631];
  assign o[631] = scan_lo[631] & N392;
  assign N392 = ~scan_lo[630];
  assign o[630] = scan_lo[630] & N393;
  assign N393 = ~scan_lo[629];
  assign o[629] = scan_lo[629] & N394;
  assign N394 = ~scan_lo[628];
  assign o[628] = scan_lo[628] & N395;
  assign N395 = ~scan_lo[627];
  assign o[627] = scan_lo[627] & N396;
  assign N396 = ~scan_lo[626];
  assign o[626] = scan_lo[626] & N397;
  assign N397 = ~scan_lo[625];
  assign o[625] = scan_lo[625] & N398;
  assign N398 = ~scan_lo[624];
  assign o[624] = scan_lo[624] & N399;
  assign N399 = ~scan_lo[623];
  assign o[623] = scan_lo[623] & N400;
  assign N400 = ~scan_lo[622];
  assign o[622] = scan_lo[622] & N401;
  assign N401 = ~scan_lo[621];
  assign o[621] = scan_lo[621] & N402;
  assign N402 = ~scan_lo[620];
  assign o[620] = scan_lo[620] & N403;
  assign N403 = ~scan_lo[619];
  assign o[619] = scan_lo[619] & N404;
  assign N404 = ~scan_lo[618];
  assign o[618] = scan_lo[618] & N405;
  assign N405 = ~scan_lo[617];
  assign o[617] = scan_lo[617] & N406;
  assign N406 = ~scan_lo[616];
  assign o[616] = scan_lo[616] & N407;
  assign N407 = ~scan_lo[615];
  assign o[615] = scan_lo[615] & N408;
  assign N408 = ~scan_lo[614];
  assign o[614] = scan_lo[614] & N409;
  assign N409 = ~scan_lo[613];
  assign o[613] = scan_lo[613] & N410;
  assign N410 = ~scan_lo[612];
  assign o[612] = scan_lo[612] & N411;
  assign N411 = ~scan_lo[611];
  assign o[611] = scan_lo[611] & N412;
  assign N412 = ~scan_lo[610];
  assign o[610] = scan_lo[610] & N413;
  assign N413 = ~scan_lo[609];
  assign o[609] = scan_lo[609] & N414;
  assign N414 = ~scan_lo[608];
  assign o[608] = scan_lo[608] & N415;
  assign N415 = ~scan_lo[607];
  assign o[607] = scan_lo[607] & N416;
  assign N416 = ~scan_lo[606];
  assign o[606] = scan_lo[606] & N417;
  assign N417 = ~scan_lo[605];
  assign o[605] = scan_lo[605] & N418;
  assign N418 = ~scan_lo[604];
  assign o[604] = scan_lo[604] & N419;
  assign N419 = ~scan_lo[603];
  assign o[603] = scan_lo[603] & N420;
  assign N420 = ~scan_lo[602];
  assign o[602] = scan_lo[602] & N421;
  assign N421 = ~scan_lo[601];
  assign o[601] = scan_lo[601] & N422;
  assign N422 = ~scan_lo[600];
  assign o[600] = scan_lo[600] & N423;
  assign N423 = ~scan_lo[599];
  assign o[599] = scan_lo[599] & N424;
  assign N424 = ~scan_lo[598];
  assign o[598] = scan_lo[598] & N425;
  assign N425 = ~scan_lo[597];
  assign o[597] = scan_lo[597] & N426;
  assign N426 = ~scan_lo[596];
  assign o[596] = scan_lo[596] & N427;
  assign N427 = ~scan_lo[595];
  assign o[595] = scan_lo[595] & N428;
  assign N428 = ~scan_lo[594];
  assign o[594] = scan_lo[594] & N429;
  assign N429 = ~scan_lo[593];
  assign o[593] = scan_lo[593] & N430;
  assign N430 = ~scan_lo[592];
  assign o[592] = scan_lo[592] & N431;
  assign N431 = ~scan_lo[591];
  assign o[591] = scan_lo[591] & N432;
  assign N432 = ~scan_lo[590];
  assign o[590] = scan_lo[590] & N433;
  assign N433 = ~scan_lo[589];
  assign o[589] = scan_lo[589] & N434;
  assign N434 = ~scan_lo[588];
  assign o[588] = scan_lo[588] & N435;
  assign N435 = ~scan_lo[587];
  assign o[587] = scan_lo[587] & N436;
  assign N436 = ~scan_lo[586];
  assign o[586] = scan_lo[586] & N437;
  assign N437 = ~scan_lo[585];
  assign o[585] = scan_lo[585] & N438;
  assign N438 = ~scan_lo[584];
  assign o[584] = scan_lo[584] & N439;
  assign N439 = ~scan_lo[583];
  assign o[583] = scan_lo[583] & N440;
  assign N440 = ~scan_lo[582];
  assign o[582] = scan_lo[582] & N441;
  assign N441 = ~scan_lo[581];
  assign o[581] = scan_lo[581] & N442;
  assign N442 = ~scan_lo[580];
  assign o[580] = scan_lo[580] & N443;
  assign N443 = ~scan_lo[579];
  assign o[579] = scan_lo[579] & N444;
  assign N444 = ~scan_lo[578];
  assign o[578] = scan_lo[578] & N445;
  assign N445 = ~scan_lo[577];
  assign o[577] = scan_lo[577] & N446;
  assign N446 = ~scan_lo[576];
  assign o[576] = scan_lo[576] & N447;
  assign N447 = ~scan_lo[575];
  assign o[575] = scan_lo[575] & N448;
  assign N448 = ~scan_lo[574];
  assign o[574] = scan_lo[574] & N449;
  assign N449 = ~scan_lo[573];
  assign o[573] = scan_lo[573] & N450;
  assign N450 = ~scan_lo[572];
  assign o[572] = scan_lo[572] & N451;
  assign N451 = ~scan_lo[571];
  assign o[571] = scan_lo[571] & N452;
  assign N452 = ~scan_lo[570];
  assign o[570] = scan_lo[570] & N453;
  assign N453 = ~scan_lo[569];
  assign o[569] = scan_lo[569] & N454;
  assign N454 = ~scan_lo[568];
  assign o[568] = scan_lo[568] & N455;
  assign N455 = ~scan_lo[567];
  assign o[567] = scan_lo[567] & N456;
  assign N456 = ~scan_lo[566];
  assign o[566] = scan_lo[566] & N457;
  assign N457 = ~scan_lo[565];
  assign o[565] = scan_lo[565] & N458;
  assign N458 = ~scan_lo[564];
  assign o[564] = scan_lo[564] & N459;
  assign N459 = ~scan_lo[563];
  assign o[563] = scan_lo[563] & N460;
  assign N460 = ~scan_lo[562];
  assign o[562] = scan_lo[562] & N461;
  assign N461 = ~scan_lo[561];
  assign o[561] = scan_lo[561] & N462;
  assign N462 = ~scan_lo[560];
  assign o[560] = scan_lo[560] & N463;
  assign N463 = ~scan_lo[559];
  assign o[559] = scan_lo[559] & N464;
  assign N464 = ~scan_lo[558];
  assign o[558] = scan_lo[558] & N465;
  assign N465 = ~scan_lo[557];
  assign o[557] = scan_lo[557] & N466;
  assign N466 = ~scan_lo[556];
  assign o[556] = scan_lo[556] & N467;
  assign N467 = ~scan_lo[555];
  assign o[555] = scan_lo[555] & N468;
  assign N468 = ~scan_lo[554];
  assign o[554] = scan_lo[554] & N469;
  assign N469 = ~scan_lo[553];
  assign o[553] = scan_lo[553] & N470;
  assign N470 = ~scan_lo[552];
  assign o[552] = scan_lo[552] & N471;
  assign N471 = ~scan_lo[551];
  assign o[551] = scan_lo[551] & N472;
  assign N472 = ~scan_lo[550];
  assign o[550] = scan_lo[550] & N473;
  assign N473 = ~scan_lo[549];
  assign o[549] = scan_lo[549] & N474;
  assign N474 = ~scan_lo[548];
  assign o[548] = scan_lo[548] & N475;
  assign N475 = ~scan_lo[547];
  assign o[547] = scan_lo[547] & N476;
  assign N476 = ~scan_lo[546];
  assign o[546] = scan_lo[546] & N477;
  assign N477 = ~scan_lo[545];
  assign o[545] = scan_lo[545] & N478;
  assign N478 = ~scan_lo[544];
  assign o[544] = scan_lo[544] & N479;
  assign N479 = ~scan_lo[543];
  assign o[543] = scan_lo[543] & N480;
  assign N480 = ~scan_lo[542];
  assign o[542] = scan_lo[542] & N481;
  assign N481 = ~scan_lo[541];
  assign o[541] = scan_lo[541] & N482;
  assign N482 = ~scan_lo[540];
  assign o[540] = scan_lo[540] & N483;
  assign N483 = ~scan_lo[539];
  assign o[539] = scan_lo[539] & N484;
  assign N484 = ~scan_lo[538];
  assign o[538] = scan_lo[538] & N485;
  assign N485 = ~scan_lo[537];
  assign o[537] = scan_lo[537] & N486;
  assign N486 = ~scan_lo[536];
  assign o[536] = scan_lo[536] & N487;
  assign N487 = ~scan_lo[535];
  assign o[535] = scan_lo[535] & N488;
  assign N488 = ~scan_lo[534];
  assign o[534] = scan_lo[534] & N489;
  assign N489 = ~scan_lo[533];
  assign o[533] = scan_lo[533] & N490;
  assign N490 = ~scan_lo[532];
  assign o[532] = scan_lo[532] & N491;
  assign N491 = ~scan_lo[531];
  assign o[531] = scan_lo[531] & N492;
  assign N492 = ~scan_lo[530];
  assign o[530] = scan_lo[530] & N493;
  assign N493 = ~scan_lo[529];
  assign o[529] = scan_lo[529] & N494;
  assign N494 = ~scan_lo[528];
  assign o[528] = scan_lo[528] & N495;
  assign N495 = ~scan_lo[527];
  assign o[527] = scan_lo[527] & N496;
  assign N496 = ~scan_lo[526];
  assign o[526] = scan_lo[526] & N497;
  assign N497 = ~scan_lo[525];
  assign o[525] = scan_lo[525] & N498;
  assign N498 = ~scan_lo[524];
  assign o[524] = scan_lo[524] & N499;
  assign N499 = ~scan_lo[523];
  assign o[523] = scan_lo[523] & N500;
  assign N500 = ~scan_lo[522];
  assign o[522] = scan_lo[522] & N501;
  assign N501 = ~scan_lo[521];
  assign o[521] = scan_lo[521] & N502;
  assign N502 = ~scan_lo[520];
  assign o[520] = scan_lo[520] & N503;
  assign N503 = ~scan_lo[519];
  assign o[519] = scan_lo[519] & N504;
  assign N504 = ~scan_lo[518];
  assign o[518] = scan_lo[518] & N505;
  assign N505 = ~scan_lo[517];
  assign o[517] = scan_lo[517] & N506;
  assign N506 = ~scan_lo[516];
  assign o[516] = scan_lo[516] & N507;
  assign N507 = ~scan_lo[515];
  assign o[515] = scan_lo[515] & N508;
  assign N508 = ~scan_lo[514];
  assign o[514] = scan_lo[514] & N509;
  assign N509 = ~scan_lo[513];
  assign o[513] = scan_lo[513] & N510;
  assign N510 = ~scan_lo[512];
  assign o[512] = scan_lo[512] & N511;
  assign N511 = ~scan_lo[511];
  assign o[511] = scan_lo[511] & N512;
  assign N512 = ~scan_lo[510];
  assign o[510] = scan_lo[510] & N513;
  assign N513 = ~scan_lo[509];
  assign o[509] = scan_lo[509] & N514;
  assign N514 = ~scan_lo[508];
  assign o[508] = scan_lo[508] & N515;
  assign N515 = ~scan_lo[507];
  assign o[507] = scan_lo[507] & N516;
  assign N516 = ~scan_lo[506];
  assign o[506] = scan_lo[506] & N517;
  assign N517 = ~scan_lo[505];
  assign o[505] = scan_lo[505] & N518;
  assign N518 = ~scan_lo[504];
  assign o[504] = scan_lo[504] & N519;
  assign N519 = ~scan_lo[503];
  assign o[503] = scan_lo[503] & N520;
  assign N520 = ~scan_lo[502];
  assign o[502] = scan_lo[502] & N521;
  assign N521 = ~scan_lo[501];
  assign o[501] = scan_lo[501] & N522;
  assign N522 = ~scan_lo[500];
  assign o[500] = scan_lo[500] & N523;
  assign N523 = ~scan_lo[499];
  assign o[499] = scan_lo[499] & N524;
  assign N524 = ~scan_lo[498];
  assign o[498] = scan_lo[498] & N525;
  assign N525 = ~scan_lo[497];
  assign o[497] = scan_lo[497] & N526;
  assign N526 = ~scan_lo[496];
  assign o[496] = scan_lo[496] & N527;
  assign N527 = ~scan_lo[495];
  assign o[495] = scan_lo[495] & N528;
  assign N528 = ~scan_lo[494];
  assign o[494] = scan_lo[494] & N529;
  assign N529 = ~scan_lo[493];
  assign o[493] = scan_lo[493] & N530;
  assign N530 = ~scan_lo[492];
  assign o[492] = scan_lo[492] & N531;
  assign N531 = ~scan_lo[491];
  assign o[491] = scan_lo[491] & N532;
  assign N532 = ~scan_lo[490];
  assign o[490] = scan_lo[490] & N533;
  assign N533 = ~scan_lo[489];
  assign o[489] = scan_lo[489] & N534;
  assign N534 = ~scan_lo[488];
  assign o[488] = scan_lo[488] & N535;
  assign N535 = ~scan_lo[487];
  assign o[487] = scan_lo[487] & N536;
  assign N536 = ~scan_lo[486];
  assign o[486] = scan_lo[486] & N537;
  assign N537 = ~scan_lo[485];
  assign o[485] = scan_lo[485] & N538;
  assign N538 = ~scan_lo[484];
  assign o[484] = scan_lo[484] & N539;
  assign N539 = ~scan_lo[483];
  assign o[483] = scan_lo[483] & N540;
  assign N540 = ~scan_lo[482];
  assign o[482] = scan_lo[482] & N541;
  assign N541 = ~scan_lo[481];
  assign o[481] = scan_lo[481] & N542;
  assign N542 = ~scan_lo[480];
  assign o[480] = scan_lo[480] & N543;
  assign N543 = ~scan_lo[479];
  assign o[479] = scan_lo[479] & N544;
  assign N544 = ~scan_lo[478];
  assign o[478] = scan_lo[478] & N545;
  assign N545 = ~scan_lo[477];
  assign o[477] = scan_lo[477] & N546;
  assign N546 = ~scan_lo[476];
  assign o[476] = scan_lo[476] & N547;
  assign N547 = ~scan_lo[475];
  assign o[475] = scan_lo[475] & N548;
  assign N548 = ~scan_lo[474];
  assign o[474] = scan_lo[474] & N549;
  assign N549 = ~scan_lo[473];
  assign o[473] = scan_lo[473] & N550;
  assign N550 = ~scan_lo[472];
  assign o[472] = scan_lo[472] & N551;
  assign N551 = ~scan_lo[471];
  assign o[471] = scan_lo[471] & N552;
  assign N552 = ~scan_lo[470];
  assign o[470] = scan_lo[470] & N553;
  assign N553 = ~scan_lo[469];
  assign o[469] = scan_lo[469] & N554;
  assign N554 = ~scan_lo[468];
  assign o[468] = scan_lo[468] & N555;
  assign N555 = ~scan_lo[467];
  assign o[467] = scan_lo[467] & N556;
  assign N556 = ~scan_lo[466];
  assign o[466] = scan_lo[466] & N557;
  assign N557 = ~scan_lo[465];
  assign o[465] = scan_lo[465] & N558;
  assign N558 = ~scan_lo[464];
  assign o[464] = scan_lo[464] & N559;
  assign N559 = ~scan_lo[463];
  assign o[463] = scan_lo[463] & N560;
  assign N560 = ~scan_lo[462];
  assign o[462] = scan_lo[462] & N561;
  assign N561 = ~scan_lo[461];
  assign o[461] = scan_lo[461] & N562;
  assign N562 = ~scan_lo[460];
  assign o[460] = scan_lo[460] & N563;
  assign N563 = ~scan_lo[459];
  assign o[459] = scan_lo[459] & N564;
  assign N564 = ~scan_lo[458];
  assign o[458] = scan_lo[458] & N565;
  assign N565 = ~scan_lo[457];
  assign o[457] = scan_lo[457] & N566;
  assign N566 = ~scan_lo[456];
  assign o[456] = scan_lo[456] & N567;
  assign N567 = ~scan_lo[455];
  assign o[455] = scan_lo[455] & N568;
  assign N568 = ~scan_lo[454];
  assign o[454] = scan_lo[454] & N569;
  assign N569 = ~scan_lo[453];
  assign o[453] = scan_lo[453] & N570;
  assign N570 = ~scan_lo[452];
  assign o[452] = scan_lo[452] & N571;
  assign N571 = ~scan_lo[451];
  assign o[451] = scan_lo[451] & N572;
  assign N572 = ~scan_lo[450];
  assign o[450] = scan_lo[450] & N573;
  assign N573 = ~scan_lo[449];
  assign o[449] = scan_lo[449] & N574;
  assign N574 = ~scan_lo[448];
  assign o[448] = scan_lo[448] & N575;
  assign N575 = ~scan_lo[447];
  assign o[447] = scan_lo[447] & N576;
  assign N576 = ~scan_lo[446];
  assign o[446] = scan_lo[446] & N577;
  assign N577 = ~scan_lo[445];
  assign o[445] = scan_lo[445] & N578;
  assign N578 = ~scan_lo[444];
  assign o[444] = scan_lo[444] & N579;
  assign N579 = ~scan_lo[443];
  assign o[443] = scan_lo[443] & N580;
  assign N580 = ~scan_lo[442];
  assign o[442] = scan_lo[442] & N581;
  assign N581 = ~scan_lo[441];
  assign o[441] = scan_lo[441] & N582;
  assign N582 = ~scan_lo[440];
  assign o[440] = scan_lo[440] & N583;
  assign N583 = ~scan_lo[439];
  assign o[439] = scan_lo[439] & N584;
  assign N584 = ~scan_lo[438];
  assign o[438] = scan_lo[438] & N585;
  assign N585 = ~scan_lo[437];
  assign o[437] = scan_lo[437] & N586;
  assign N586 = ~scan_lo[436];
  assign o[436] = scan_lo[436] & N587;
  assign N587 = ~scan_lo[435];
  assign o[435] = scan_lo[435] & N588;
  assign N588 = ~scan_lo[434];
  assign o[434] = scan_lo[434] & N589;
  assign N589 = ~scan_lo[433];
  assign o[433] = scan_lo[433] & N590;
  assign N590 = ~scan_lo[432];
  assign o[432] = scan_lo[432] & N591;
  assign N591 = ~scan_lo[431];
  assign o[431] = scan_lo[431] & N592;
  assign N592 = ~scan_lo[430];
  assign o[430] = scan_lo[430] & N593;
  assign N593 = ~scan_lo[429];
  assign o[429] = scan_lo[429] & N594;
  assign N594 = ~scan_lo[428];
  assign o[428] = scan_lo[428] & N595;
  assign N595 = ~scan_lo[427];
  assign o[427] = scan_lo[427] & N596;
  assign N596 = ~scan_lo[426];
  assign o[426] = scan_lo[426] & N597;
  assign N597 = ~scan_lo[425];
  assign o[425] = scan_lo[425] & N598;
  assign N598 = ~scan_lo[424];
  assign o[424] = scan_lo[424] & N599;
  assign N599 = ~scan_lo[423];
  assign o[423] = scan_lo[423] & N600;
  assign N600 = ~scan_lo[422];
  assign o[422] = scan_lo[422] & N601;
  assign N601 = ~scan_lo[421];
  assign o[421] = scan_lo[421] & N602;
  assign N602 = ~scan_lo[420];
  assign o[420] = scan_lo[420] & N603;
  assign N603 = ~scan_lo[419];
  assign o[419] = scan_lo[419] & N604;
  assign N604 = ~scan_lo[418];
  assign o[418] = scan_lo[418] & N605;
  assign N605 = ~scan_lo[417];
  assign o[417] = scan_lo[417] & N606;
  assign N606 = ~scan_lo[416];
  assign o[416] = scan_lo[416] & N607;
  assign N607 = ~scan_lo[415];
  assign o[415] = scan_lo[415] & N608;
  assign N608 = ~scan_lo[414];
  assign o[414] = scan_lo[414] & N609;
  assign N609 = ~scan_lo[413];
  assign o[413] = scan_lo[413] & N610;
  assign N610 = ~scan_lo[412];
  assign o[412] = scan_lo[412] & N611;
  assign N611 = ~scan_lo[411];
  assign o[411] = scan_lo[411] & N612;
  assign N612 = ~scan_lo[410];
  assign o[410] = scan_lo[410] & N613;
  assign N613 = ~scan_lo[409];
  assign o[409] = scan_lo[409] & N614;
  assign N614 = ~scan_lo[408];
  assign o[408] = scan_lo[408] & N615;
  assign N615 = ~scan_lo[407];
  assign o[407] = scan_lo[407] & N616;
  assign N616 = ~scan_lo[406];
  assign o[406] = scan_lo[406] & N617;
  assign N617 = ~scan_lo[405];
  assign o[405] = scan_lo[405] & N618;
  assign N618 = ~scan_lo[404];
  assign o[404] = scan_lo[404] & N619;
  assign N619 = ~scan_lo[403];
  assign o[403] = scan_lo[403] & N620;
  assign N620 = ~scan_lo[402];
  assign o[402] = scan_lo[402] & N621;
  assign N621 = ~scan_lo[401];
  assign o[401] = scan_lo[401] & N622;
  assign N622 = ~scan_lo[400];
  assign o[400] = scan_lo[400] & N623;
  assign N623 = ~scan_lo[399];
  assign o[399] = scan_lo[399] & N624;
  assign N624 = ~scan_lo[398];
  assign o[398] = scan_lo[398] & N625;
  assign N625 = ~scan_lo[397];
  assign o[397] = scan_lo[397] & N626;
  assign N626 = ~scan_lo[396];
  assign o[396] = scan_lo[396] & N627;
  assign N627 = ~scan_lo[395];
  assign o[395] = scan_lo[395] & N628;
  assign N628 = ~scan_lo[394];
  assign o[394] = scan_lo[394] & N629;
  assign N629 = ~scan_lo[393];
  assign o[393] = scan_lo[393] & N630;
  assign N630 = ~scan_lo[392];
  assign o[392] = scan_lo[392] & N631;
  assign N631 = ~scan_lo[391];
  assign o[391] = scan_lo[391] & N632;
  assign N632 = ~scan_lo[390];
  assign o[390] = scan_lo[390] & N633;
  assign N633 = ~scan_lo[389];
  assign o[389] = scan_lo[389] & N634;
  assign N634 = ~scan_lo[388];
  assign o[388] = scan_lo[388] & N635;
  assign N635 = ~scan_lo[387];
  assign o[387] = scan_lo[387] & N636;
  assign N636 = ~scan_lo[386];
  assign o[386] = scan_lo[386] & N637;
  assign N637 = ~scan_lo[385];
  assign o[385] = scan_lo[385] & N638;
  assign N638 = ~scan_lo[384];
  assign o[384] = scan_lo[384] & N639;
  assign N639 = ~scan_lo[383];
  assign o[383] = scan_lo[383] & N640;
  assign N640 = ~scan_lo[382];
  assign o[382] = scan_lo[382] & N641;
  assign N641 = ~scan_lo[381];
  assign o[381] = scan_lo[381] & N642;
  assign N642 = ~scan_lo[380];
  assign o[380] = scan_lo[380] & N643;
  assign N643 = ~scan_lo[379];
  assign o[379] = scan_lo[379] & N644;
  assign N644 = ~scan_lo[378];
  assign o[378] = scan_lo[378] & N645;
  assign N645 = ~scan_lo[377];
  assign o[377] = scan_lo[377] & N646;
  assign N646 = ~scan_lo[376];
  assign o[376] = scan_lo[376] & N647;
  assign N647 = ~scan_lo[375];
  assign o[375] = scan_lo[375] & N648;
  assign N648 = ~scan_lo[374];
  assign o[374] = scan_lo[374] & N649;
  assign N649 = ~scan_lo[373];
  assign o[373] = scan_lo[373] & N650;
  assign N650 = ~scan_lo[372];
  assign o[372] = scan_lo[372] & N651;
  assign N651 = ~scan_lo[371];
  assign o[371] = scan_lo[371] & N652;
  assign N652 = ~scan_lo[370];
  assign o[370] = scan_lo[370] & N653;
  assign N653 = ~scan_lo[369];
  assign o[369] = scan_lo[369] & N654;
  assign N654 = ~scan_lo[368];
  assign o[368] = scan_lo[368] & N655;
  assign N655 = ~scan_lo[367];
  assign o[367] = scan_lo[367] & N656;
  assign N656 = ~scan_lo[366];
  assign o[366] = scan_lo[366] & N657;
  assign N657 = ~scan_lo[365];
  assign o[365] = scan_lo[365] & N658;
  assign N658 = ~scan_lo[364];
  assign o[364] = scan_lo[364] & N659;
  assign N659 = ~scan_lo[363];
  assign o[363] = scan_lo[363] & N660;
  assign N660 = ~scan_lo[362];
  assign o[362] = scan_lo[362] & N661;
  assign N661 = ~scan_lo[361];
  assign o[361] = scan_lo[361] & N662;
  assign N662 = ~scan_lo[360];
  assign o[360] = scan_lo[360] & N663;
  assign N663 = ~scan_lo[359];
  assign o[359] = scan_lo[359] & N664;
  assign N664 = ~scan_lo[358];
  assign o[358] = scan_lo[358] & N665;
  assign N665 = ~scan_lo[357];
  assign o[357] = scan_lo[357] & N666;
  assign N666 = ~scan_lo[356];
  assign o[356] = scan_lo[356] & N667;
  assign N667 = ~scan_lo[355];
  assign o[355] = scan_lo[355] & N668;
  assign N668 = ~scan_lo[354];
  assign o[354] = scan_lo[354] & N669;
  assign N669 = ~scan_lo[353];
  assign o[353] = scan_lo[353] & N670;
  assign N670 = ~scan_lo[352];
  assign o[352] = scan_lo[352] & N671;
  assign N671 = ~scan_lo[351];
  assign o[351] = scan_lo[351] & N672;
  assign N672 = ~scan_lo[350];
  assign o[350] = scan_lo[350] & N673;
  assign N673 = ~scan_lo[349];
  assign o[349] = scan_lo[349] & N674;
  assign N674 = ~scan_lo[348];
  assign o[348] = scan_lo[348] & N675;
  assign N675 = ~scan_lo[347];
  assign o[347] = scan_lo[347] & N676;
  assign N676 = ~scan_lo[346];
  assign o[346] = scan_lo[346] & N677;
  assign N677 = ~scan_lo[345];
  assign o[345] = scan_lo[345] & N678;
  assign N678 = ~scan_lo[344];
  assign o[344] = scan_lo[344] & N679;
  assign N679 = ~scan_lo[343];
  assign o[343] = scan_lo[343] & N680;
  assign N680 = ~scan_lo[342];
  assign o[342] = scan_lo[342] & N681;
  assign N681 = ~scan_lo[341];
  assign o[341] = scan_lo[341] & N682;
  assign N682 = ~scan_lo[340];
  assign o[340] = scan_lo[340] & N683;
  assign N683 = ~scan_lo[339];
  assign o[339] = scan_lo[339] & N684;
  assign N684 = ~scan_lo[338];
  assign o[338] = scan_lo[338] & N685;
  assign N685 = ~scan_lo[337];
  assign o[337] = scan_lo[337] & N686;
  assign N686 = ~scan_lo[336];
  assign o[336] = scan_lo[336] & N687;
  assign N687 = ~scan_lo[335];
  assign o[335] = scan_lo[335] & N688;
  assign N688 = ~scan_lo[334];
  assign o[334] = scan_lo[334] & N689;
  assign N689 = ~scan_lo[333];
  assign o[333] = scan_lo[333] & N690;
  assign N690 = ~scan_lo[332];
  assign o[332] = scan_lo[332] & N691;
  assign N691 = ~scan_lo[331];
  assign o[331] = scan_lo[331] & N692;
  assign N692 = ~scan_lo[330];
  assign o[330] = scan_lo[330] & N693;
  assign N693 = ~scan_lo[329];
  assign o[329] = scan_lo[329] & N694;
  assign N694 = ~scan_lo[328];
  assign o[328] = scan_lo[328] & N695;
  assign N695 = ~scan_lo[327];
  assign o[327] = scan_lo[327] & N696;
  assign N696 = ~scan_lo[326];
  assign o[326] = scan_lo[326] & N697;
  assign N697 = ~scan_lo[325];
  assign o[325] = scan_lo[325] & N698;
  assign N698 = ~scan_lo[324];
  assign o[324] = scan_lo[324] & N699;
  assign N699 = ~scan_lo[323];
  assign o[323] = scan_lo[323] & N700;
  assign N700 = ~scan_lo[322];
  assign o[322] = scan_lo[322] & N701;
  assign N701 = ~scan_lo[321];
  assign o[321] = scan_lo[321] & N702;
  assign N702 = ~scan_lo[320];
  assign o[320] = scan_lo[320] & N703;
  assign N703 = ~scan_lo[319];
  assign o[319] = scan_lo[319] & N704;
  assign N704 = ~scan_lo[318];
  assign o[318] = scan_lo[318] & N705;
  assign N705 = ~scan_lo[317];
  assign o[317] = scan_lo[317] & N706;
  assign N706 = ~scan_lo[316];
  assign o[316] = scan_lo[316] & N707;
  assign N707 = ~scan_lo[315];
  assign o[315] = scan_lo[315] & N708;
  assign N708 = ~scan_lo[314];
  assign o[314] = scan_lo[314] & N709;
  assign N709 = ~scan_lo[313];
  assign o[313] = scan_lo[313] & N710;
  assign N710 = ~scan_lo[312];
  assign o[312] = scan_lo[312] & N711;
  assign N711 = ~scan_lo[311];
  assign o[311] = scan_lo[311] & N712;
  assign N712 = ~scan_lo[310];
  assign o[310] = scan_lo[310] & N713;
  assign N713 = ~scan_lo[309];
  assign o[309] = scan_lo[309] & N714;
  assign N714 = ~scan_lo[308];
  assign o[308] = scan_lo[308] & N715;
  assign N715 = ~scan_lo[307];
  assign o[307] = scan_lo[307] & N716;
  assign N716 = ~scan_lo[306];
  assign o[306] = scan_lo[306] & N717;
  assign N717 = ~scan_lo[305];
  assign o[305] = scan_lo[305] & N718;
  assign N718 = ~scan_lo[304];
  assign o[304] = scan_lo[304] & N719;
  assign N719 = ~scan_lo[303];
  assign o[303] = scan_lo[303] & N720;
  assign N720 = ~scan_lo[302];
  assign o[302] = scan_lo[302] & N721;
  assign N721 = ~scan_lo[301];
  assign o[301] = scan_lo[301] & N722;
  assign N722 = ~scan_lo[300];
  assign o[300] = scan_lo[300] & N723;
  assign N723 = ~scan_lo[299];
  assign o[299] = scan_lo[299] & N724;
  assign N724 = ~scan_lo[298];
  assign o[298] = scan_lo[298] & N725;
  assign N725 = ~scan_lo[297];
  assign o[297] = scan_lo[297] & N726;
  assign N726 = ~scan_lo[296];
  assign o[296] = scan_lo[296] & N727;
  assign N727 = ~scan_lo[295];
  assign o[295] = scan_lo[295] & N728;
  assign N728 = ~scan_lo[294];
  assign o[294] = scan_lo[294] & N729;
  assign N729 = ~scan_lo[293];
  assign o[293] = scan_lo[293] & N730;
  assign N730 = ~scan_lo[292];
  assign o[292] = scan_lo[292] & N731;
  assign N731 = ~scan_lo[291];
  assign o[291] = scan_lo[291] & N732;
  assign N732 = ~scan_lo[290];
  assign o[290] = scan_lo[290] & N733;
  assign N733 = ~scan_lo[289];
  assign o[289] = scan_lo[289] & N734;
  assign N734 = ~scan_lo[288];
  assign o[288] = scan_lo[288] & N735;
  assign N735 = ~scan_lo[287];
  assign o[287] = scan_lo[287] & N736;
  assign N736 = ~scan_lo[286];
  assign o[286] = scan_lo[286] & N737;
  assign N737 = ~scan_lo[285];
  assign o[285] = scan_lo[285] & N738;
  assign N738 = ~scan_lo[284];
  assign o[284] = scan_lo[284] & N739;
  assign N739 = ~scan_lo[283];
  assign o[283] = scan_lo[283] & N740;
  assign N740 = ~scan_lo[282];
  assign o[282] = scan_lo[282] & N741;
  assign N741 = ~scan_lo[281];
  assign o[281] = scan_lo[281] & N742;
  assign N742 = ~scan_lo[280];
  assign o[280] = scan_lo[280] & N743;
  assign N743 = ~scan_lo[279];
  assign o[279] = scan_lo[279] & N744;
  assign N744 = ~scan_lo[278];
  assign o[278] = scan_lo[278] & N745;
  assign N745 = ~scan_lo[277];
  assign o[277] = scan_lo[277] & N746;
  assign N746 = ~scan_lo[276];
  assign o[276] = scan_lo[276] & N747;
  assign N747 = ~scan_lo[275];
  assign o[275] = scan_lo[275] & N748;
  assign N748 = ~scan_lo[274];
  assign o[274] = scan_lo[274] & N749;
  assign N749 = ~scan_lo[273];
  assign o[273] = scan_lo[273] & N750;
  assign N750 = ~scan_lo[272];
  assign o[272] = scan_lo[272] & N751;
  assign N751 = ~scan_lo[271];
  assign o[271] = scan_lo[271] & N752;
  assign N752 = ~scan_lo[270];
  assign o[270] = scan_lo[270] & N753;
  assign N753 = ~scan_lo[269];
  assign o[269] = scan_lo[269] & N754;
  assign N754 = ~scan_lo[268];
  assign o[268] = scan_lo[268] & N755;
  assign N755 = ~scan_lo[267];
  assign o[267] = scan_lo[267] & N756;
  assign N756 = ~scan_lo[266];
  assign o[266] = scan_lo[266] & N757;
  assign N757 = ~scan_lo[265];
  assign o[265] = scan_lo[265] & N758;
  assign N758 = ~scan_lo[264];
  assign o[264] = scan_lo[264] & N759;
  assign N759 = ~scan_lo[263];
  assign o[263] = scan_lo[263] & N760;
  assign N760 = ~scan_lo[262];
  assign o[262] = scan_lo[262] & N761;
  assign N761 = ~scan_lo[261];
  assign o[261] = scan_lo[261] & N762;
  assign N762 = ~scan_lo[260];
  assign o[260] = scan_lo[260] & N763;
  assign N763 = ~scan_lo[259];
  assign o[259] = scan_lo[259] & N764;
  assign N764 = ~scan_lo[258];
  assign o[258] = scan_lo[258] & N765;
  assign N765 = ~scan_lo[257];
  assign o[257] = scan_lo[257] & N766;
  assign N766 = ~scan_lo[256];
  assign o[256] = scan_lo[256] & N767;
  assign N767 = ~scan_lo[255];
  assign o[255] = scan_lo[255] & N768;
  assign N768 = ~scan_lo[254];
  assign o[254] = scan_lo[254] & N769;
  assign N769 = ~scan_lo[253];
  assign o[253] = scan_lo[253] & N770;
  assign N770 = ~scan_lo[252];
  assign o[252] = scan_lo[252] & N771;
  assign N771 = ~scan_lo[251];
  assign o[251] = scan_lo[251] & N772;
  assign N772 = ~scan_lo[250];
  assign o[250] = scan_lo[250] & N773;
  assign N773 = ~scan_lo[249];
  assign o[249] = scan_lo[249] & N774;
  assign N774 = ~scan_lo[248];
  assign o[248] = scan_lo[248] & N775;
  assign N775 = ~scan_lo[247];
  assign o[247] = scan_lo[247] & N776;
  assign N776 = ~scan_lo[246];
  assign o[246] = scan_lo[246] & N777;
  assign N777 = ~scan_lo[245];
  assign o[245] = scan_lo[245] & N778;
  assign N778 = ~scan_lo[244];
  assign o[244] = scan_lo[244] & N779;
  assign N779 = ~scan_lo[243];
  assign o[243] = scan_lo[243] & N780;
  assign N780 = ~scan_lo[242];
  assign o[242] = scan_lo[242] & N781;
  assign N781 = ~scan_lo[241];
  assign o[241] = scan_lo[241] & N782;
  assign N782 = ~scan_lo[240];
  assign o[240] = scan_lo[240] & N783;
  assign N783 = ~scan_lo[239];
  assign o[239] = scan_lo[239] & N784;
  assign N784 = ~scan_lo[238];
  assign o[238] = scan_lo[238] & N785;
  assign N785 = ~scan_lo[237];
  assign o[237] = scan_lo[237] & N786;
  assign N786 = ~scan_lo[236];
  assign o[236] = scan_lo[236] & N787;
  assign N787 = ~scan_lo[235];
  assign o[235] = scan_lo[235] & N788;
  assign N788 = ~scan_lo[234];
  assign o[234] = scan_lo[234] & N789;
  assign N789 = ~scan_lo[233];
  assign o[233] = scan_lo[233] & N790;
  assign N790 = ~scan_lo[232];
  assign o[232] = scan_lo[232] & N791;
  assign N791 = ~scan_lo[231];
  assign o[231] = scan_lo[231] & N792;
  assign N792 = ~scan_lo[230];
  assign o[230] = scan_lo[230] & N793;
  assign N793 = ~scan_lo[229];
  assign o[229] = scan_lo[229] & N794;
  assign N794 = ~scan_lo[228];
  assign o[228] = scan_lo[228] & N795;
  assign N795 = ~scan_lo[227];
  assign o[227] = scan_lo[227] & N796;
  assign N796 = ~scan_lo[226];
  assign o[226] = scan_lo[226] & N797;
  assign N797 = ~scan_lo[225];
  assign o[225] = scan_lo[225] & N798;
  assign N798 = ~scan_lo[224];
  assign o[224] = scan_lo[224] & N799;
  assign N799 = ~scan_lo[223];
  assign o[223] = scan_lo[223] & N800;
  assign N800 = ~scan_lo[222];
  assign o[222] = scan_lo[222] & N801;
  assign N801 = ~scan_lo[221];
  assign o[221] = scan_lo[221] & N802;
  assign N802 = ~scan_lo[220];
  assign o[220] = scan_lo[220] & N803;
  assign N803 = ~scan_lo[219];
  assign o[219] = scan_lo[219] & N804;
  assign N804 = ~scan_lo[218];
  assign o[218] = scan_lo[218] & N805;
  assign N805 = ~scan_lo[217];
  assign o[217] = scan_lo[217] & N806;
  assign N806 = ~scan_lo[216];
  assign o[216] = scan_lo[216] & N807;
  assign N807 = ~scan_lo[215];
  assign o[215] = scan_lo[215] & N808;
  assign N808 = ~scan_lo[214];
  assign o[214] = scan_lo[214] & N809;
  assign N809 = ~scan_lo[213];
  assign o[213] = scan_lo[213] & N810;
  assign N810 = ~scan_lo[212];
  assign o[212] = scan_lo[212] & N811;
  assign N811 = ~scan_lo[211];
  assign o[211] = scan_lo[211] & N812;
  assign N812 = ~scan_lo[210];
  assign o[210] = scan_lo[210] & N813;
  assign N813 = ~scan_lo[209];
  assign o[209] = scan_lo[209] & N814;
  assign N814 = ~scan_lo[208];
  assign o[208] = scan_lo[208] & N815;
  assign N815 = ~scan_lo[207];
  assign o[207] = scan_lo[207] & N816;
  assign N816 = ~scan_lo[206];
  assign o[206] = scan_lo[206] & N817;
  assign N817 = ~scan_lo[205];
  assign o[205] = scan_lo[205] & N818;
  assign N818 = ~scan_lo[204];
  assign o[204] = scan_lo[204] & N819;
  assign N819 = ~scan_lo[203];
  assign o[203] = scan_lo[203] & N820;
  assign N820 = ~scan_lo[202];
  assign o[202] = scan_lo[202] & N821;
  assign N821 = ~scan_lo[201];
  assign o[201] = scan_lo[201] & N822;
  assign N822 = ~scan_lo[200];
  assign o[200] = scan_lo[200] & N823;
  assign N823 = ~scan_lo[199];
  assign o[199] = scan_lo[199] & N824;
  assign N824 = ~scan_lo[198];
  assign o[198] = scan_lo[198] & N825;
  assign N825 = ~scan_lo[197];
  assign o[197] = scan_lo[197] & N826;
  assign N826 = ~scan_lo[196];
  assign o[196] = scan_lo[196] & N827;
  assign N827 = ~scan_lo[195];
  assign o[195] = scan_lo[195] & N828;
  assign N828 = ~scan_lo[194];
  assign o[194] = scan_lo[194] & N829;
  assign N829 = ~scan_lo[193];
  assign o[193] = scan_lo[193] & N830;
  assign N830 = ~scan_lo[192];
  assign o[192] = scan_lo[192] & N831;
  assign N831 = ~scan_lo[191];
  assign o[191] = scan_lo[191] & N832;
  assign N832 = ~scan_lo[190];
  assign o[190] = scan_lo[190] & N833;
  assign N833 = ~scan_lo[189];
  assign o[189] = scan_lo[189] & N834;
  assign N834 = ~scan_lo[188];
  assign o[188] = scan_lo[188] & N835;
  assign N835 = ~scan_lo[187];
  assign o[187] = scan_lo[187] & N836;
  assign N836 = ~scan_lo[186];
  assign o[186] = scan_lo[186] & N837;
  assign N837 = ~scan_lo[185];
  assign o[185] = scan_lo[185] & N838;
  assign N838 = ~scan_lo[184];
  assign o[184] = scan_lo[184] & N839;
  assign N839 = ~scan_lo[183];
  assign o[183] = scan_lo[183] & N840;
  assign N840 = ~scan_lo[182];
  assign o[182] = scan_lo[182] & N841;
  assign N841 = ~scan_lo[181];
  assign o[181] = scan_lo[181] & N842;
  assign N842 = ~scan_lo[180];
  assign o[180] = scan_lo[180] & N843;
  assign N843 = ~scan_lo[179];
  assign o[179] = scan_lo[179] & N844;
  assign N844 = ~scan_lo[178];
  assign o[178] = scan_lo[178] & N845;
  assign N845 = ~scan_lo[177];
  assign o[177] = scan_lo[177] & N846;
  assign N846 = ~scan_lo[176];
  assign o[176] = scan_lo[176] & N847;
  assign N847 = ~scan_lo[175];
  assign o[175] = scan_lo[175] & N848;
  assign N848 = ~scan_lo[174];
  assign o[174] = scan_lo[174] & N849;
  assign N849 = ~scan_lo[173];
  assign o[173] = scan_lo[173] & N850;
  assign N850 = ~scan_lo[172];
  assign o[172] = scan_lo[172] & N851;
  assign N851 = ~scan_lo[171];
  assign o[171] = scan_lo[171] & N852;
  assign N852 = ~scan_lo[170];
  assign o[170] = scan_lo[170] & N853;
  assign N853 = ~scan_lo[169];
  assign o[169] = scan_lo[169] & N854;
  assign N854 = ~scan_lo[168];
  assign o[168] = scan_lo[168] & N855;
  assign N855 = ~scan_lo[167];
  assign o[167] = scan_lo[167] & N856;
  assign N856 = ~scan_lo[166];
  assign o[166] = scan_lo[166] & N857;
  assign N857 = ~scan_lo[165];
  assign o[165] = scan_lo[165] & N858;
  assign N858 = ~scan_lo[164];
  assign o[164] = scan_lo[164] & N859;
  assign N859 = ~scan_lo[163];
  assign o[163] = scan_lo[163] & N860;
  assign N860 = ~scan_lo[162];
  assign o[162] = scan_lo[162] & N861;
  assign N861 = ~scan_lo[161];
  assign o[161] = scan_lo[161] & N862;
  assign N862 = ~scan_lo[160];
  assign o[160] = scan_lo[160] & N863;
  assign N863 = ~scan_lo[159];
  assign o[159] = scan_lo[159] & N864;
  assign N864 = ~scan_lo[158];
  assign o[158] = scan_lo[158] & N865;
  assign N865 = ~scan_lo[157];
  assign o[157] = scan_lo[157] & N866;
  assign N866 = ~scan_lo[156];
  assign o[156] = scan_lo[156] & N867;
  assign N867 = ~scan_lo[155];
  assign o[155] = scan_lo[155] & N868;
  assign N868 = ~scan_lo[154];
  assign o[154] = scan_lo[154] & N869;
  assign N869 = ~scan_lo[153];
  assign o[153] = scan_lo[153] & N870;
  assign N870 = ~scan_lo[152];
  assign o[152] = scan_lo[152] & N871;
  assign N871 = ~scan_lo[151];
  assign o[151] = scan_lo[151] & N872;
  assign N872 = ~scan_lo[150];
  assign o[150] = scan_lo[150] & N873;
  assign N873 = ~scan_lo[149];
  assign o[149] = scan_lo[149] & N874;
  assign N874 = ~scan_lo[148];
  assign o[148] = scan_lo[148] & N875;
  assign N875 = ~scan_lo[147];
  assign o[147] = scan_lo[147] & N876;
  assign N876 = ~scan_lo[146];
  assign o[146] = scan_lo[146] & N877;
  assign N877 = ~scan_lo[145];
  assign o[145] = scan_lo[145] & N878;
  assign N878 = ~scan_lo[144];
  assign o[144] = scan_lo[144] & N879;
  assign N879 = ~scan_lo[143];
  assign o[143] = scan_lo[143] & N880;
  assign N880 = ~scan_lo[142];
  assign o[142] = scan_lo[142] & N881;
  assign N881 = ~scan_lo[141];
  assign o[141] = scan_lo[141] & N882;
  assign N882 = ~scan_lo[140];
  assign o[140] = scan_lo[140] & N883;
  assign N883 = ~scan_lo[139];
  assign o[139] = scan_lo[139] & N884;
  assign N884 = ~scan_lo[138];
  assign o[138] = scan_lo[138] & N885;
  assign N885 = ~scan_lo[137];
  assign o[137] = scan_lo[137] & N886;
  assign N886 = ~scan_lo[136];
  assign o[136] = scan_lo[136] & N887;
  assign N887 = ~scan_lo[135];
  assign o[135] = scan_lo[135] & N888;
  assign N888 = ~scan_lo[134];
  assign o[134] = scan_lo[134] & N889;
  assign N889 = ~scan_lo[133];
  assign o[133] = scan_lo[133] & N890;
  assign N890 = ~scan_lo[132];
  assign o[132] = scan_lo[132] & N891;
  assign N891 = ~scan_lo[131];
  assign o[131] = scan_lo[131] & N892;
  assign N892 = ~scan_lo[130];
  assign o[130] = scan_lo[130] & N893;
  assign N893 = ~scan_lo[129];
  assign o[129] = scan_lo[129] & N894;
  assign N894 = ~scan_lo[128];
  assign o[128] = scan_lo[128] & N895;
  assign N895 = ~scan_lo[127];
  assign o[127] = scan_lo[127] & N896;
  assign N896 = ~scan_lo[126];
  assign o[126] = scan_lo[126] & N897;
  assign N897 = ~scan_lo[125];
  assign o[125] = scan_lo[125] & N898;
  assign N898 = ~scan_lo[124];
  assign o[124] = scan_lo[124] & N899;
  assign N899 = ~scan_lo[123];
  assign o[123] = scan_lo[123] & N900;
  assign N900 = ~scan_lo[122];
  assign o[122] = scan_lo[122] & N901;
  assign N901 = ~scan_lo[121];
  assign o[121] = scan_lo[121] & N902;
  assign N902 = ~scan_lo[120];
  assign o[120] = scan_lo[120] & N903;
  assign N903 = ~scan_lo[119];
  assign o[119] = scan_lo[119] & N904;
  assign N904 = ~scan_lo[118];
  assign o[118] = scan_lo[118] & N905;
  assign N905 = ~scan_lo[117];
  assign o[117] = scan_lo[117] & N906;
  assign N906 = ~scan_lo[116];
  assign o[116] = scan_lo[116] & N907;
  assign N907 = ~scan_lo[115];
  assign o[115] = scan_lo[115] & N908;
  assign N908 = ~scan_lo[114];
  assign o[114] = scan_lo[114] & N909;
  assign N909 = ~scan_lo[113];
  assign o[113] = scan_lo[113] & N910;
  assign N910 = ~scan_lo[112];
  assign o[112] = scan_lo[112] & N911;
  assign N911 = ~scan_lo[111];
  assign o[111] = scan_lo[111] & N912;
  assign N912 = ~scan_lo[110];
  assign o[110] = scan_lo[110] & N913;
  assign N913 = ~scan_lo[109];
  assign o[109] = scan_lo[109] & N914;
  assign N914 = ~scan_lo[108];
  assign o[108] = scan_lo[108] & N915;
  assign N915 = ~scan_lo[107];
  assign o[107] = scan_lo[107] & N916;
  assign N916 = ~scan_lo[106];
  assign o[106] = scan_lo[106] & N917;
  assign N917 = ~scan_lo[105];
  assign o[105] = scan_lo[105] & N918;
  assign N918 = ~scan_lo[104];
  assign o[104] = scan_lo[104] & N919;
  assign N919 = ~scan_lo[103];
  assign o[103] = scan_lo[103] & N920;
  assign N920 = ~scan_lo[102];
  assign o[102] = scan_lo[102] & N921;
  assign N921 = ~scan_lo[101];
  assign o[101] = scan_lo[101] & N922;
  assign N922 = ~scan_lo[100];
  assign o[100] = scan_lo[100] & N923;
  assign N923 = ~scan_lo[99];
  assign o[99] = scan_lo[99] & N924;
  assign N924 = ~scan_lo[98];
  assign o[98] = scan_lo[98] & N925;
  assign N925 = ~scan_lo[97];
  assign o[97] = scan_lo[97] & N926;
  assign N926 = ~scan_lo[96];
  assign o[96] = scan_lo[96] & N927;
  assign N927 = ~scan_lo[95];
  assign o[95] = scan_lo[95] & N928;
  assign N928 = ~scan_lo[94];
  assign o[94] = scan_lo[94] & N929;
  assign N929 = ~scan_lo[93];
  assign o[93] = scan_lo[93] & N930;
  assign N930 = ~scan_lo[92];
  assign o[92] = scan_lo[92] & N931;
  assign N931 = ~scan_lo[91];
  assign o[91] = scan_lo[91] & N932;
  assign N932 = ~scan_lo[90];
  assign o[90] = scan_lo[90] & N933;
  assign N933 = ~scan_lo[89];
  assign o[89] = scan_lo[89] & N934;
  assign N934 = ~scan_lo[88];
  assign o[88] = scan_lo[88] & N935;
  assign N935 = ~scan_lo[87];
  assign o[87] = scan_lo[87] & N936;
  assign N936 = ~scan_lo[86];
  assign o[86] = scan_lo[86] & N937;
  assign N937 = ~scan_lo[85];
  assign o[85] = scan_lo[85] & N938;
  assign N938 = ~scan_lo[84];
  assign o[84] = scan_lo[84] & N939;
  assign N939 = ~scan_lo[83];
  assign o[83] = scan_lo[83] & N940;
  assign N940 = ~scan_lo[82];
  assign o[82] = scan_lo[82] & N941;
  assign N941 = ~scan_lo[81];
  assign o[81] = scan_lo[81] & N942;
  assign N942 = ~scan_lo[80];
  assign o[80] = scan_lo[80] & N943;
  assign N943 = ~scan_lo[79];
  assign o[79] = scan_lo[79] & N944;
  assign N944 = ~scan_lo[78];
  assign o[78] = scan_lo[78] & N945;
  assign N945 = ~scan_lo[77];
  assign o[77] = scan_lo[77] & N946;
  assign N946 = ~scan_lo[76];
  assign o[76] = scan_lo[76] & N947;
  assign N947 = ~scan_lo[75];
  assign o[75] = scan_lo[75] & N948;
  assign N948 = ~scan_lo[74];
  assign o[74] = scan_lo[74] & N949;
  assign N949 = ~scan_lo[73];
  assign o[73] = scan_lo[73] & N950;
  assign N950 = ~scan_lo[72];
  assign o[72] = scan_lo[72] & N951;
  assign N951 = ~scan_lo[71];
  assign o[71] = scan_lo[71] & N952;
  assign N952 = ~scan_lo[70];
  assign o[70] = scan_lo[70] & N953;
  assign N953 = ~scan_lo[69];
  assign o[69] = scan_lo[69] & N954;
  assign N954 = ~scan_lo[68];
  assign o[68] = scan_lo[68] & N955;
  assign N955 = ~scan_lo[67];
  assign o[67] = scan_lo[67] & N956;
  assign N956 = ~scan_lo[66];
  assign o[66] = scan_lo[66] & N957;
  assign N957 = ~scan_lo[65];
  assign o[65] = scan_lo[65] & N958;
  assign N958 = ~scan_lo[64];
  assign o[64] = scan_lo[64] & N959;
  assign N959 = ~scan_lo[63];
  assign o[63] = scan_lo[63] & N960;
  assign N960 = ~scan_lo[62];
  assign o[62] = scan_lo[62] & N961;
  assign N961 = ~scan_lo[61];
  assign o[61] = scan_lo[61] & N962;
  assign N962 = ~scan_lo[60];
  assign o[60] = scan_lo[60] & N963;
  assign N963 = ~scan_lo[59];
  assign o[59] = scan_lo[59] & N964;
  assign N964 = ~scan_lo[58];
  assign o[58] = scan_lo[58] & N965;
  assign N965 = ~scan_lo[57];
  assign o[57] = scan_lo[57] & N966;
  assign N966 = ~scan_lo[56];
  assign o[56] = scan_lo[56] & N967;
  assign N967 = ~scan_lo[55];
  assign o[55] = scan_lo[55] & N968;
  assign N968 = ~scan_lo[54];
  assign o[54] = scan_lo[54] & N969;
  assign N969 = ~scan_lo[53];
  assign o[53] = scan_lo[53] & N970;
  assign N970 = ~scan_lo[52];
  assign o[52] = scan_lo[52] & N971;
  assign N971 = ~scan_lo[51];
  assign o[51] = scan_lo[51] & N972;
  assign N972 = ~scan_lo[50];
  assign o[50] = scan_lo[50] & N973;
  assign N973 = ~scan_lo[49];
  assign o[49] = scan_lo[49] & N974;
  assign N974 = ~scan_lo[48];
  assign o[48] = scan_lo[48] & N975;
  assign N975 = ~scan_lo[47];
  assign o[47] = scan_lo[47] & N976;
  assign N976 = ~scan_lo[46];
  assign o[46] = scan_lo[46] & N977;
  assign N977 = ~scan_lo[45];
  assign o[45] = scan_lo[45] & N978;
  assign N978 = ~scan_lo[44];
  assign o[44] = scan_lo[44] & N979;
  assign N979 = ~scan_lo[43];
  assign o[43] = scan_lo[43] & N980;
  assign N980 = ~scan_lo[42];
  assign o[42] = scan_lo[42] & N981;
  assign N981 = ~scan_lo[41];
  assign o[41] = scan_lo[41] & N982;
  assign N982 = ~scan_lo[40];
  assign o[40] = scan_lo[40] & N983;
  assign N983 = ~scan_lo[39];
  assign o[39] = scan_lo[39] & N984;
  assign N984 = ~scan_lo[38];
  assign o[38] = scan_lo[38] & N985;
  assign N985 = ~scan_lo[37];
  assign o[37] = scan_lo[37] & N986;
  assign N986 = ~scan_lo[36];
  assign o[36] = scan_lo[36] & N987;
  assign N987 = ~scan_lo[35];
  assign o[35] = scan_lo[35] & N988;
  assign N988 = ~scan_lo[34];
  assign o[34] = scan_lo[34] & N989;
  assign N989 = ~scan_lo[33];
  assign o[33] = scan_lo[33] & N990;
  assign N990 = ~scan_lo[32];
  assign o[32] = scan_lo[32] & N991;
  assign N991 = ~scan_lo[31];
  assign o[31] = scan_lo[31] & N992;
  assign N992 = ~scan_lo[30];
  assign o[30] = scan_lo[30] & N993;
  assign N993 = ~scan_lo[29];
  assign o[29] = scan_lo[29] & N994;
  assign N994 = ~scan_lo[28];
  assign o[28] = scan_lo[28] & N995;
  assign N995 = ~scan_lo[27];
  assign o[27] = scan_lo[27] & N996;
  assign N996 = ~scan_lo[26];
  assign o[26] = scan_lo[26] & N997;
  assign N997 = ~scan_lo[25];
  assign o[25] = scan_lo[25] & N998;
  assign N998 = ~scan_lo[24];
  assign o[24] = scan_lo[24] & N999;
  assign N999 = ~scan_lo[23];
  assign o[23] = scan_lo[23] & N1000;
  assign N1000 = ~scan_lo[22];
  assign o[22] = scan_lo[22] & N1001;
  assign N1001 = ~scan_lo[21];
  assign o[21] = scan_lo[21] & N1002;
  assign N1002 = ~scan_lo[20];
  assign o[20] = scan_lo[20] & N1003;
  assign N1003 = ~scan_lo[19];
  assign o[19] = scan_lo[19] & N1004;
  assign N1004 = ~scan_lo[18];
  assign o[18] = scan_lo[18] & N1005;
  assign N1005 = ~scan_lo[17];
  assign o[17] = scan_lo[17] & N1006;
  assign N1006 = ~scan_lo[16];
  assign o[16] = scan_lo[16] & N1007;
  assign N1007 = ~scan_lo[15];
  assign o[15] = scan_lo[15] & N1008;
  assign N1008 = ~scan_lo[14];
  assign o[14] = scan_lo[14] & N1009;
  assign N1009 = ~scan_lo[13];
  assign o[13] = scan_lo[13] & N1010;
  assign N1010 = ~scan_lo[12];
  assign o[12] = scan_lo[12] & N1011;
  assign N1011 = ~scan_lo[11];
  assign o[11] = scan_lo[11] & N1012;
  assign N1012 = ~scan_lo[10];
  assign o[10] = scan_lo[10] & N1013;
  assign N1013 = ~scan_lo[9];
  assign o[9] = scan_lo[9] & N1014;
  assign N1014 = ~scan_lo[8];
  assign o[8] = scan_lo[8] & N1015;
  assign N1015 = ~scan_lo[7];
  assign o[7] = scan_lo[7] & N1016;
  assign N1016 = ~scan_lo[6];
  assign o[6] = scan_lo[6] & N1017;
  assign N1017 = ~scan_lo[5];
  assign o[5] = scan_lo[5] & N1018;
  assign N1018 = ~scan_lo[4];
  assign o[4] = scan_lo[4] & N1019;
  assign N1019 = ~scan_lo[3];
  assign o[3] = scan_lo[3] & N1020;
  assign N1020 = ~scan_lo[2];
  assign o[2] = scan_lo[2] & N1021;
  assign N1021 = ~scan_lo[1];
  assign o[1] = scan_lo[1] & N1022;
  assign N1022 = ~o[0];

endmodule



module bsg_encode_one_hot_width_p1
(
  i,
  addr_o,
  v_o
);

  input [0:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o;
  wire v_o;
  assign v_o = i[0];
  assign addr_o[0] = 1'b0;

endmodule



module bsg_encode_one_hot_width_p2
(
  i,
  addr_o,
  v_o
);

  input [1:0] i;
  output [0:0] addr_o;
  output v_o;
  wire [0:0] addr_o,aligned_vs;
  wire v_o;
  wire [1:0] aligned_addrs;

  bsg_encode_one_hot_width_p1
  aligned_left
  (
    .i(i[0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p1
  aligned_right
  (
    .i(i[1]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[0])
  );

  assign v_o = addr_o[0] | aligned_vs[0];

endmodule



module bsg_encode_one_hot_width_p4
(
  i,
  addr_o,
  v_o
);

  input [3:0] i;
  output [1:0] addr_o;
  output v_o;
  wire [1:0] addr_o,aligned_addrs;
  wire v_o;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p2
  aligned_left
  (
    .i(i[1:0]),
    .addr_o(aligned_addrs[0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p2
  aligned_right
  (
    .i(i[3:2]),
    .addr_o(aligned_addrs[1]),
    .v_o(addr_o[1])
  );

  assign v_o = addr_o[1] | aligned_vs[0];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[1];

endmodule



module bsg_encode_one_hot_width_p8
(
  i,
  addr_o,
  v_o
);

  input [7:0] i;
  output [2:0] addr_o;
  output v_o;
  wire [2:0] addr_o;
  wire v_o;
  wire [3:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p4
  aligned_left
  (
    .i(i[3:0]),
    .addr_o(aligned_addrs[1:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p4
  aligned_right
  (
    .i(i[7:4]),
    .addr_o(aligned_addrs[3:2]),
    .v_o(addr_o[2])
  );

  assign v_o = addr_o[2] | aligned_vs[0];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[3];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[2];

endmodule



module bsg_encode_one_hot_width_p16
(
  i,
  addr_o,
  v_o
);

  input [15:0] i;
  output [3:0] addr_o;
  output v_o;
  wire [3:0] addr_o;
  wire v_o;
  wire [5:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p8
  aligned_left
  (
    .i(i[7:0]),
    .addr_o(aligned_addrs[2:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p8
  aligned_right
  (
    .i(i[15:8]),
    .addr_o(aligned_addrs[5:3]),
    .v_o(addr_o[3])
  );

  assign v_o = addr_o[3] | aligned_vs[0];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[5];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[4];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[3];

endmodule



module bsg_encode_one_hot_width_p32
(
  i,
  addr_o,
  v_o
);

  input [31:0] i;
  output [4:0] addr_o;
  output v_o;
  wire [4:0] addr_o;
  wire v_o;
  wire [7:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p16
  aligned_left
  (
    .i(i[15:0]),
    .addr_o(aligned_addrs[3:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p16
  aligned_right
  (
    .i(i[31:16]),
    .addr_o(aligned_addrs[7:4]),
    .v_o(addr_o[4])
  );

  assign v_o = addr_o[4] | aligned_vs[0];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[7];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[6];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[5];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[4];

endmodule



module bsg_encode_one_hot_width_p64
(
  i,
  addr_o,
  v_o
);

  input [63:0] i;
  output [5:0] addr_o;
  output v_o;
  wire [5:0] addr_o;
  wire v_o;
  wire [9:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p32
  aligned_left
  (
    .i(i[31:0]),
    .addr_o(aligned_addrs[4:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p32
  aligned_right
  (
    .i(i[63:32]),
    .addr_o(aligned_addrs[9:5]),
    .v_o(addr_o[5])
  );

  assign v_o = addr_o[5] | aligned_vs[0];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[9];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[8];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[7];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[6];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[5];

endmodule



module bsg_encode_one_hot_width_p128
(
  i,
  addr_o,
  v_o
);

  input [127:0] i;
  output [6:0] addr_o;
  output v_o;
  wire [6:0] addr_o;
  wire v_o;
  wire [11:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p64
  aligned_left
  (
    .i(i[63:0]),
    .addr_o(aligned_addrs[5:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p64
  aligned_right
  (
    .i(i[127:64]),
    .addr_o(aligned_addrs[11:6]),
    .v_o(addr_o[6])
  );

  assign v_o = addr_o[6] | aligned_vs[0];
  assign addr_o[5] = aligned_addrs[5] | aligned_addrs[11];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[10];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[9];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[8];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[7];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[6];

endmodule



module bsg_encode_one_hot_width_p256
(
  i,
  addr_o,
  v_o
);

  input [255:0] i;
  output [7:0] addr_o;
  output v_o;
  wire [7:0] addr_o;
  wire v_o;
  wire [13:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p128
  aligned_left
  (
    .i(i[127:0]),
    .addr_o(aligned_addrs[6:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p128
  aligned_right
  (
    .i(i[255:128]),
    .addr_o(aligned_addrs[13:7]),
    .v_o(addr_o[7])
  );

  assign v_o = addr_o[7] | aligned_vs[0];
  assign addr_o[6] = aligned_addrs[6] | aligned_addrs[13];
  assign addr_o[5] = aligned_addrs[5] | aligned_addrs[12];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[11];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[10];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[9];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[8];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[7];

endmodule



module bsg_encode_one_hot_width_p512
(
  i,
  addr_o,
  v_o
);

  input [511:0] i;
  output [8:0] addr_o;
  output v_o;
  wire [8:0] addr_o;
  wire v_o;
  wire [15:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p256
  aligned_left
  (
    .i(i[255:0]),
    .addr_o(aligned_addrs[7:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p256
  aligned_right
  (
    .i(i[511:256]),
    .addr_o(aligned_addrs[15:8]),
    .v_o(addr_o[8])
  );

  assign v_o = addr_o[8] | aligned_vs[0];
  assign addr_o[7] = aligned_addrs[7] | aligned_addrs[15];
  assign addr_o[6] = aligned_addrs[6] | aligned_addrs[14];
  assign addr_o[5] = aligned_addrs[5] | aligned_addrs[13];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[12];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[11];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[10];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[9];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[8];

endmodule



module bsg_encode_one_hot_width_p1024_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [1023:0] i;
  output [9:0] addr_o;
  output v_o;
  wire [9:0] addr_o;
  wire v_o;
  wire [17:0] aligned_addrs;
  wire [0:0] aligned_vs;

  bsg_encode_one_hot_width_p512
  aligned_left
  (
    .i(i[511:0]),
    .addr_o(aligned_addrs[8:0]),
    .v_o(aligned_vs[0])
  );


  bsg_encode_one_hot_width_p512
  aligned_right
  (
    .i(i[1023:512]),
    .addr_o(aligned_addrs[17:9]),
    .v_o(addr_o[9])
  );

  assign v_o = addr_o[9] | aligned_vs[0];
  assign addr_o[8] = aligned_addrs[8] | aligned_addrs[17];
  assign addr_o[7] = aligned_addrs[7] | aligned_addrs[16];
  assign addr_o[6] = aligned_addrs[6] | aligned_addrs[15];
  assign addr_o[5] = aligned_addrs[5] | aligned_addrs[14];
  assign addr_o[4] = aligned_addrs[4] | aligned_addrs[13];
  assign addr_o[3] = aligned_addrs[3] | aligned_addrs[12];
  assign addr_o[2] = aligned_addrs[2] | aligned_addrs[11];
  assign addr_o[1] = aligned_addrs[1] | aligned_addrs[10];
  assign addr_o[0] = aligned_addrs[0] | aligned_addrs[9];

endmodule



module bsg_priority_encode_width_p1024_lo_to_hi_p1
(
  i,
  addr_o,
  v_o
);

  input [1023:0] i;
  output [9:0] addr_o;
  output v_o;
  wire [9:0] addr_o;
  wire v_o;
  wire [1023:0] enc_lo;

  bsg_priority_encode_one_hot_out_width_p1024_lo_to_hi_p1
  a
  (
    .i(i),
    .o(enc_lo)
  );


  bsg_encode_one_hot_width_p1024_lo_to_hi_p1
  b
  (
    .i(enc_lo),
    .addr_o(addr_o),
    .v_o(v_o)
  );


endmodule



module bsg_cam_1r1w
(
  clk_i,
  reset_i,
  en_i,
  w_v_i,
  w_set_not_clear_i,
  w_addr_i,
  w_data_i,
  r_v_i,
  r_data_i,
  r_v_o,
  r_addr_o,
  empty_v_o,
  empty_addr_o
);

  input [9:0] w_addr_i;
  input [31:0] w_data_i;
  input [31:0] r_data_i;
  output [9:0] r_addr_o;
  output [9:0] empty_addr_o;
  input clk_i;
  input reset_i;
  input en_i;
  input w_v_i;
  input w_set_not_clear_i;
  input r_v_i;
  output r_v_o;
  output empty_v_o;
  wire [9:0] r_addr_o,empty_addr_o;
  wire r_v_o,empty_v_o,N0,N1,N2,N3,N4,N5,N6,N7,N8,N9,N10,N11,N12,N13,N14,N15,N16,
  matched,empty_found,N17,N18,N19,N20,N21,N22,N23,N24,N25,N26,N27,N28,N29,N30,N31,N32,
  N33,N34,N35,N36,N37,N38,N39,N40,N41,N42,N43,N44,N45,N46,N47,N48,N49,N50,N51,N52,
  N53,N54,N55,N56,N57,N58,N59,N60,N61,N62,N63,N64,N65,N66,N67,N68,N69,N70,N71,N72,
  N73,N74,N75,N76,N77,N78,N79,N80,N81,N82,N83,N84,N85,N86,N87,N88,N89,N90,N91,N92,
  N93,N94,N95,N96,N97,N98,N99,N100,N101,N102,N103,N104,N105,N106,N107,N108,N109,
  N110,N111,N112,N113,N114,N115,N116,N117,N118,N119,N120,N121,N122,N123,N124,N125,
  N126,N127,N128,N129,N130,N131,N132,N133,N134,N135,N136,N137,N138,N139,N140,N141,
  N142,N143,N144,N145,N146,N147,N148,N149,N150,N151,N152,N153,N154,N155,N156,N157,
  N158,N159,N160,N161,N162,N163,N164,N165,N166,N167,N168,N169,N170,N171,N172,N173,
  N174,N175,N176,N177,N178,N179,N180,N181,N182,N183,N184,N185,N186,N187,N188,N189,
  N190,N191,N192,N193,N194,N195,N196,N197,N198,N199,N200,N201,N202,N203,N204,N205,
  N206,N207,N208,N209,N210,N211,N212,N213,N214,N215,N216,N217,N218,N219,N220,N221,
  N222,N223,N224,N225,N226,N227,N228,N229,N230,N231,N232,N233,N234,N235,N236,N237,
  N238,N239,N240,N241,N242,N243,N244,N245,N246,N247,N248,N249,N250,N251,N252,N253,
  N254,N255,N256,N257,N258,N259,N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
  N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,N280,N281,N282,N283,N284,N285,
  N286,N287,N288,N289,N290,N291,N292,N293,N294,N295,N296,N297,N298,N299,N300,N301,
  N302,N303,N304,N305,N306,N307,N308,N309,N310,N311,N312,N313,N314,N315,N316,N317,
  N318,N319,N320,N321,N322,N323,N324,N325,N326,N327,N328,N329,N330,N331,N332,N333,
  N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,N349,
  N350,N351,N352,N353,N354,N355,N356,N357,N358,N359,N360,N361,N362,N363,N364,N365,
  N366,N367,N368,N369,N370,N371,N372,N373,N374,N375,N376,N377,N378,N379,N380,N381,
  N382,N383,N384,N385,N386,N387,N388,N389,N390,N391,N392,N393,N394,N395,N396,N397,
  N398,N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,N409,N410,N411,N412,N413,
  N414,N415,N416,N417,N418,N419,N420,N421,N422,N423,N424,N425,N426,N427,N428,N429,
  N430,N431,N432,N433,N434,N435,N436,N437,N438,N439,N440,N441,N442,N443,N444,N445,
  N446,N447,N448,N449,N450,N451,N452,N453,N454,N455,N456,N457,N458,N459,N460,N461,
  N462,N463,N464,N465,N466,N467,N468,N469,N470,N471,N472,N473,N474,N475,N476,N477,
  N478,N479,N480,N481,N482,N483,N484,N485,N486,N487,N488,N489,N490,N491,N492,N493,
  N494,N495,N496,N497,N498,N499,N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
  N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,N520,N521,N522,N523,N524,N525,
  N526,N527,N528,N529,N530,N531,N532,N533,N534,N535,N536,N537,N538,N539,N540,N541,
  N542,N543,N544,N545,N546,N547,N548,N549,N550,N551,N552,N553,N554,N555,N556,N557,
  N558,N559,N560,N561,N562,N563,N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
  N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,N584,N585,N586,N587,N588,N589,
  N590,N591,N592,N593,N594,N595,N596,N597,N598,N599,N600,N601,N602,N603,N604,N605,
  N606,N607,N608,N609,N610,N611,N612,N613,N614,N615,N616,N617,N618,N619,N620,N621,
  N622,N623,N624,N625,N626,N627,N628,N629,N630,N631,N632,N633,N634,N635,N636,N637,
  N638,N639,N640,N641,N642,N643,N644,N645,N646,N647,N648,N649,N650,N651,N652,N653,
  N654,N655,N656,N657,N658,N659,N660,N661,N662,N663,N664,N665,N666,N667,N668,N669,
  N670,N671,N672,N673,N674,N675,N676,N677,N678,N679,N680,N681,N682,N683,N684,N685,
  N686,N687,N688,N689,N690,N691,N692,N693,N694,N695,N696,N697,N698,N699,N700,N701,
  N702,N703,N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,N714,N715,N716,N717,
  N718,N719,N720,N721,N722,N723,N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
  N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,N744,N745,N746,N747,N748,N749,
  N750,N751,N752,N753,N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,N764,N765,
  N766,N767,N768,N769,N770,N771,N772,N773,N774,N775,N776,N777,N778,N779,N780,N781,
  N782,N783,N784,N785,N786,N787,N788,N789,N790,N791,N792,N793,N794,N795,N796,N797,
  N798,N799,N800,N801,N802,N803,N804,N805,N806,N807,N808,N809,N810,N811,N812,N813,
  N814,N815,N816,N817,N818,N819,N820,N821,N822,N823,N824,N825,N826,N827,N828,N829,
  N830,N831,N832,N833,N834,N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,N845,
  N846,N847,N848,N849,N850,N851,N852,N853,N854,N855,N856,N857,N858,N859,N860,N861,
  N862,N863,N864,N865,N866,N867,N868,N869,N870,N871,N872,N873,N874,N875,N876,N877,
  N878,N879,N880,N881,N882,N883,N884,N885,N886,N887,N888,N889,N890,N891,N892,N893,
  N894,N895,N896,N897,N898,N899,N900,N901,N902,N903,N904,N905,N906,N907,N908,N909,
  N910,N911,N912,N913,N914,N915,N916,N917,N918,N919,N920,N921,N922,N923,N924,N925,
  N926,N927,N928,N929,N930,N931,N932,N933,N934,N935,N936,N937,N938,N939,N940,N941,
  N942,N943,N944,N945,N946,N947,N948,N949,N950,N951,N952,N953,N954,N955,N956,N957,
  N958,N959,N960,N961,N962,N963,N964,N965,N966,N967,N968,N969,N970,N971,N972,N973,
  N974,N975,N976,N977,N978,N979,N980,N981,N982,N983,N984,N985,N986,N987,N988,N989,
  N990,N991,N992,N993,N994,N995,N996,N997,N998,N999,N1000,N1001,N1002,N1003,N1004,
  N1005,N1006,N1007,N1008,N1009,N1010,N1011,N1012,N1013,N1014,N1015,N1016,N1017,N1018,
  N1019,N1020,N1021,N1022,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030,N1031,
  N1032,N1033,N1034,N1035,N1036,N1037,N1038,N1039,N1040,N1041,N1042,N1043,N1044,
  N1045,N1046,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054,N1055,N1056,N1057,N1058,
  N1059,N1060,N1061,N1062,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1071,
  N1072,N1073,N1074,N1075,N1076,N1077,N1078,N1079,N1080,N1081,N1082,N1083,N1084,
  N1085,N1086,N1087,N1088,N1089,N1090,N1091,N1092,N1093,N1094,N1095,N1096,N1097,N1098,
  N1099,N1100,N1101,N1102,N1103,N1104,N1105,N1106,N1107,N1108,N1109,N1110,N1111,
  N1112,N1113,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121,N1122,N1123,N1124,
  N1125,N1126,N1127,N1128,N1129,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137,N1138,
  N1139,N1140,N1141,N1142,N1143,N1144,N1145,N1146,N1147,N1148,N1149,N1150,N1151,
  N1152,N1153,N1154,N1155,N1156,N1157,N1158,N1159,N1160,N1161,N1162,N1163,N1164,
  N1165,N1166,N1167,N1168,N1169,N1170,N1171,N1172,N1173,N1174,N1175,N1176,N1177,N1178,
  N1179,N1180,N1181,N1182,N1183,N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1191,
  N1192,N1193,N1194,N1195,N1196,N1197,N1198,N1199,N1200,N1201,N1202,N1203,N1204,
  N1205,N1206,N1207,N1208,N1209,N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1217,N1218,
  N1219,N1220,N1221,N1222,N1223,N1224,N1225,N1226,N1227,N1228,N1229,N1230,N1231,
  N1232,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240,N1241,N1242,N1243,N1244,
  N1245,N1246,N1247,N1248,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256,N1257,N1258,
  N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266,N1267,N1268,N1269,N1270,N1271,
  N1272,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284,
  N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296,N1297,N1298,
  N1299,N1300,N1301,N1302,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310,N1311,
  N1312,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320,N1321,N1322,N1323,N1324,
  N1325,N1326,N1327,N1328,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336,N1337,N1338,
  N1339,N1340,N1341,N1342,N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,
  N1352,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362,N1363,N1364,
  N1365,N1366,N1367,N1368,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376,N1377,N1378,
  N1379,N1380,N1381,N1382,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390,N1391,
  N1392,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400,N1401,N1402,N1403,N1404,
  N1405,N1406,N1407,N1408,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416,N1417,N1418,
  N1419,N1420,N1421,N1422,N1423,N1424,N1425,N1426,N1427,N1428,N1429,N1430,N1431,
  N1432,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442,N1443,N1444,
  N1445,N1446,N1447,N1448,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1456,N1457,N1458,
  N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,
  N1472,N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484,
  N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496,N1497,N1498,
  N1499,N1500,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508,N1509,N1510,N1511,
  N1512,N1513,N1514,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523,N1524,
  N1525,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
  N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549,N1550,N1551,
  N1552,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563,N1564,
  N1565,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,N1577,N1578,
  N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,
  N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1601,N1602,N1603,N1604,
  N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1618,
  N1619,N1620,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630,N1631,
  N1632,N1633,N1634,N1635,N1636,N1637,N1638,N1639,N1640,N1641,N1642,N1643,N1644,
  N1645,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656,N1657,N1658,
  N1659,N1660,N1661,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670,N1671,
  N1672,N1673,N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1681,N1682,N1683,N1684,
  N1685,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694,N1695,N1696,N1697,N1698,
  N1699,N1700,N1701,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710,N1711,
  N1712,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720,N1721,N1722,N1723,N1724,
  N1725,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736,N1737,N1738,
  N1739,N1740,N1741,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750,N1751,
  N1752,N1753,N1754,N1755,N1756,N1757,N1758,N1759,N1760,N1761,N1762,N1763,N1764,
  N1765,N1766,N1767,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775,N1776,N1777,N1778,
  N1779,N1780,N1781,N1782,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791,
  N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,N1800,N1801,N1802,N1803,N1804,
  N1805,N1806,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814,N1815,N1816,N1817,N1818,
  N1819,N1820,N1821,N1822,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830,N1831,
  N1832,N1833,N1834,N1835,N1836,N1837,N1838,N1839,N1840,N1841,N1842,N1843,N1844,
  N1845,N1846,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,
  N1859,N1860,N1861,N1862,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870,N1871,
  N1872,N1873,N1874,N1875,N1876,N1877,N1878,N1879,N1880,N1881,N1882,N1883,N1884,
  N1885,N1886,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894,N1895,N1896,N1897,N1898,
  N1899,N1900,N1901,N1902,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910,N1911,
  N1912,N1913,N1914,N1915,N1916,N1917,N1918,N1919,N1920,N1921,N1922,N1923,N1924,
  N1925,N1926,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,N1937,N1938,
  N1939,N1940,N1941,N1942,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950,N1951,
  N1952,N1953,N1954,N1955,N1956,N1957,N1958,N1959,N1960,N1961,N1962,N1963,N1964,
  N1965,N1966,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974,N1975,N1976,N1977,N1978,
  N1979,N1980,N1981,N1982,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990,N1991,
  N1992,N1993,N1994,N1995,N1996,N1997,N1998,N1999,N2000,N2001,N2002,N2003,N2004,
  N2005,N2006,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014,N2015,N2016,N2017,N2018,
  N2019,N2020,N2021,N2022,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,
  N2032,N2033,N2034,N2035,N2036,N2037,N2038,N2039,N2040,N2041,N2042,N2043,N2044,
  N2045,N2046,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054,N2055,N2056,N2057,N2058,
  N2059,N2060,N2061,N2062,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070,N2071,
  N2072,N2073,N2074,N2075,N2076,N2077,N2078,N2079,N2080,N2081,N2082,N2083,N2084,
  N2085,N2086,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094,N2095,N2096,N2097,N2098,
  N2099,N2100,N2101,N2102,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110,N2111,
  N2112,N2113,N2114,N2115,N2116,N2117,N2118,N2119,N2120,N2121,N2122,N2123,N2124,
  N2125,N2126,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134,N2135,N2136,N2137,N2138,
  N2139,N2140,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150,N2151,
  N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161,N2162,N2163,N2164,
  N2165,N2166,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2178,
  N2179,N2180,N2181,N2182,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190,N2191,
  N2192,N2193,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204,
  N2205,N2206,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217,N2218,
  N2219,N2220,N2221,N2222,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230,N2231,
  N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243,N2244,
  N2245,N2246,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254,N2255,N2256,N2257,N2258,
  N2259,N2260,N2261,N2262,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270,N2271,
  N2272,N2273,N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2281,N2282,N2283,N2284,
  N2285,N2286,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298,
  N2299,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310,N2311,
  N2312,N2313,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321,N2322,N2323,N2324,
  N2325,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
  N2339,N2340,N2341,N2342,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350,N2351,
  N2352,N2353,N2354,N2355,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363,N2364,
  N2365,N2366,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374,N2375,N2376,N2377,N2378,
  N2379,N2380,N2381,N2382,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390,N2391,
  N2392,N2393,N2394,N2395,N2396,N2397,N2398,N2399,N2400,N2401,N2402,N2403,N2404,
  N2405,N2406,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418,
  N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430,N2431,
  N2432,N2433,N2434,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444,
  N2445,N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454,N2455,N2456,N2457,N2458,
  N2459,N2460,N2461,N2462,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470,N2471,
  N2472,N2473,N2474,N2475,N2476,N2477,N2478,N2479,N2480,N2481,N2482,N2483,N2484,
  N2485,N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494,N2495,N2496,N2497,N2498,
  N2499,N2500,N2501,N2502,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510,N2511,
  N2512,N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520,N2521,N2522,N2523,N2524,
  N2525,N2526,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537,N2538,
  N2539,N2540,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550,N2551,
  N2552,N2553,N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564,
  N2565,N2566,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574,N2575,N2576,N2577,N2578,
  N2579,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590,N2591,
  N2592,N2593,N2594,N2595,N2596,N2597,N2598,N2599,N2600,N2601,N2602,N2603,N2604,
  N2605,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616,N2617,N2618,
  N2619,N2620,N2621,N2622,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630,N2631,
  N2632,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640,N2641,N2642,N2643,N2644,
  N2645,N2646,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657,N2658,
  N2659,N2660,N2661,N2662,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670,N2671,
  N2672,N2673,N2674,N2675,N2676,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2684,
  N2685,N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694,N2695,N2696,N2697,N2698,
  N2699,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710,N2711,
  N2712,N2713,N2714,N2715,N2716,N2717,N2718,N2719,N2720,N2721,N2722,N2723,N2724,
  N2725,N2726,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
  N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750,N2751,
  N2752,N2753,N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761,N2762,N2763,N2764,
  N2765,N2766,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777,N2778,
  N2779,N2780,N2781,N2782,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790,N2791,
  N2792,N2793,N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801,N2802,N2803,N2804,
  N2805,N2806,N2807,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817,N2818,
  N2819,N2820,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828,N2829,N2830,N2831,
  N2832,N2833,N2834,N2835,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844,
  N2845,N2846,N2847,N2848,N2849,N2850,N2851,N2852,N2853,N2854,N2855,N2856,N2857,N2858,
  N2859,N2860,N2861,N2862,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870,N2871,
  N2872,N2873,N2874,N2875,N2876,N2877,N2878,N2879,N2880,N2881,N2882,N2883,N2884,
  N2885,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895,N2896,N2897,N2898,
  N2899,N2900,N2901,N2902,N2903,N2904,N2905,N2906,N2907,N2908,N2909,N2910,N2911,
  N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2922,N2923,N2924,
  N2925,N2926,N2927,N2928,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936,N2937,N2938,
  N2939,N2940,N2941,N2942,N2943,N2944,N2945,N2946,N2947,N2948,N2949,N2950,N2951,
  N2952,N2953,N2954,N2955,N2956,N2957,N2958,N2959,N2960,N2961,N2962,N2963,N2964,
  N2965,N2966,N2967,N2968,N2969,N2970,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978,
  N2979,N2980,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,
  N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3004,
  N3005,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013,N3014,N3015,N3016,N3017,N3018,
  N3019,N3020,N3021,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,
  N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,N3042,N3043,N3044,
  N3045,N3046,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054,N3055,N3056,N3057,N3058,
  N3059,N3060,N3061,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,
  N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,N3082,N3083,N3084,
  N3085,N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097,N3098,
  N3099,N3100,N3101,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,
  N3112,N3113,N3114,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122,N3123,N3124,
  N3125,N3126,N3127,N3128,N3129,N3130,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138,
  N3139,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147,N3148,N3149,N3150,N3151,
  N3152,N3153,N3154,N3155,N3156,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164,
  N3165,N3166,N3167,N3168,N3169,N3170,N3171,N3172,N3173,N3174,N3175,N3176,N3177,N3178,
  N3179,N3180,N3181,N3182,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190,N3191,
  N3192,N3193,N3194,N3195,N3196,N3197,N3198,N3199,N3200,N3201,N3202,N3203,N3204,
  N3205,N3206,N3207,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,
  N3219,N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231,
  N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240,N3241,N3242,N3243,N3244,
  N3245,N3246,N3247,N3248,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,
  N3259,N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,N3270,N3271,
  N3272,N3273,N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282,N3283,N3284,
  N3285,N3286,N3287,N3288,N3289,N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,
  N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,N3310,N3311,
  N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324,
  N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333,N3334,N3335,N3336,N3337,N3338,
  N3339,N3340,N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3348,N3349,N3350,N3351,
  N3352,N3353,N3354,N3355,N3356,N3357,N3358,N3359,N3360,N3361,N3362,N3363,N3364,
  N3365,N3366,N3367,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375,N3376,N3377,N3378,
  N3379,N3380,N3381,N3382,N3383,N3384,N3385,N3386,N3387,N3388,N3389,N3390,N3391,
  N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403,N3404,
  N3405,N3406,N3407,N3408,N3409,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417,N3418,
  N3419,N3420,N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428,N3429,N3430,N3431,
  N3432,N3433,N3434,N3435,N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443,N3444,
  N3445,N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458,
  N3459,N3460,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471,
  N3472,N3473,N3474,N3475,N3476,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484,
  N3485,N3486,N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3495,N3496,N3497,N3498,
  N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,N3509,N3510,N3511,
  N3512,N3513,N3514,N3515,N3516,N3517,N3518,N3519,N3520,N3521,N3522,N3523,N3524,
  N3525,N3526,N3527,N3528,N3529,N3530,N3531,N3532,N3533,N3534,N3535,N3536,N3537,N3538,
  N3539,N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,N3550,N3551,
  N3552,N3553,N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561,N3562,N3563,N3564,
  N3565,N3566,N3567,N3568,N3569,N3570,N3571,N3572,N3573,N3574,N3575,N3576,N3577,N3578,
  N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3591,
  N3592,N3593,N3594,N3595,N3596,N3597,N3598,N3599,N3600,N3601,N3602,N3603,N3604,
  N3605,N3606,N3607,N3608,N3609,N3610,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618,
  N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630,N3631,
  N3632,N3633,N3634,N3635,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,
  N3645,N3646,N3647,N3648,N3649,N3650,N3651,N3652,N3653,N3654,N3655,N3656,N3657,N3658,
  N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669,N3670,N3671,
  N3672,N3673,N3674,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682,N3683,N3684,
  N3685,N3686,N3687,N3688,N3689,N3690,N3691,N3692,N3693,N3694,N3695,N3696,N3697,N3698,
  N3699,N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707,N3708,N3709,N3710,N3711,
  N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,N3722,N3723,N3724,
  N3725,N3726,N3727,N3728,N3729,N3730,N3731,N3732,N3733,N3734,N3735,N3736,N3737,N3738,
  N3739,N3740,N3741,N3742,N3743,N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3751,
  N3752,N3753,N3754,N3755,N3756,N3757,N3758,N3759,N3760,N3761,N3762,N3763,N3764,
  N3765,N3766,N3767,N3768,N3769,N3770,N3771,N3772,N3773,N3774,N3775,N3776,N3777,N3778,
  N3779,N3780,N3781,N3782,N3783,N3784,N3785,N3786,N3787,N3788,N3789,N3790,N3791,
  N3792,N3793,N3794,N3795,N3796,N3797,N3798,N3799,N3800,N3801,N3802,N3803,N3804,
  N3805,N3806,N3807,N3808,N3809,N3810,N3811,N3812,N3813,N3814,N3815,N3816,N3817,N3818,
  N3819,N3820,N3821,N3822,N3823,N3824,N3825,N3826,N3827,N3828,N3829,N3830,N3831,
  N3832,N3833,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3841,N3842,N3843,N3844,
  N3845,N3846,N3847,N3848,N3849,N3850,N3851,N3852,N3853,N3854,N3855,N3856,N3857,N3858,
  N3859,N3860,N3861,N3862,N3863,N3864,N3865,N3866,N3867,N3868,N3869,N3870,N3871,
  N3872,N3873,N3874,N3875,N3876,N3877,N3878,N3879,N3880,N3881,N3882,N3883,N3884,
  N3885,N3886,N3887,N3888,N3889,N3890,N3891,N3892,N3893,N3894,N3895,N3896,N3897,N3898,
  N3899,N3900,N3901,N3902,N3903,N3904,N3905,N3906,N3907,N3908,N3909,N3910,N3911,
  N3912,N3913,N3914,N3915,N3916,N3917,N3918,N3919,N3920,N3921,N3922,N3923,N3924,
  N3925,N3926,N3927,N3928,N3929,N3930,N3931,N3932,N3933,N3934,N3935,N3936,N3937,N3938,
  N3939,N3940,N3941,N3942,N3943,N3944,N3945,N3946,N3947,N3948,N3949,N3950,N3951,
  N3952,N3953,N3954,N3955,N3956,N3957,N3958,N3959,N3960,N3961,N3962,N3963,N3964,
  N3965,N3966,N3967,N3968,N3969,N3970,N3971,N3972,N3973,N3974,N3975,N3976,N3977,N3978,
  N3979,N3980,N3981,N3982,N3983,N3984,N3985,N3986,N3987,N3988,N3989,N3990,N3991,
  N3992,N3993,N3994,N3995,N3996,N3997,N3998,N3999,N4000,N4001,N4002,N4003,N4004,
  N4005,N4006,N4007,N4008,N4009,N4010,N4011,N4012,N4013,N4014,N4015,N4016,N4017,N4018,
  N4019,N4020,N4021,N4022,N4023,N4024,N4025,N4026,N4027,N4028,N4029,N4030,N4031,
  N4032,N4033,N4034,N4035,N4036,N4037,N4038,N4039,N4040,N4041,N4042,N4043,N4044,
  N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,N4055,N4056,N4057,N4058,
  N4059,N4060,N4061,N4062,N4063,N4064,N4065,N4066,N4067,N4068,N4069,N4070,N4071,
  N4072,N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4081,N4082,N4083,N4084,
  N4085,N4086,N4087,N4088,N4089,N4090,N4091,N4092,N4093,N4094,N4095,N4096,N4097,N4098,
  N4099,N4100,N4101,N4102,N4103,N4104,N4105,N4106,N4107,N4108,N4109,N4110,N4111,
  N4112,N4113,N4114,N4115,N4116,N4117,N4118,N4119,N4120,N4121,N4122,N4123,N4124,
  N4125,N4126,N4127,N4128,N4129,N4130,N4131,N4132,N4133,N4134,N4135,N4136,N4137,N4138,
  N4139,N4140,N4141,N4142,N4143,N4144,N4145,N4146,N4147,N4148,N4149,N4150,N4151,
  N4152,N4153,N4154,N4155,N4156,N4157,N4158,N4159,N4160,N4161,N4162,N4163,N4164,
  N4165,N4166,N4167,N4168,N4169,N4170,N4171,N4172,N4173,N4174,N4175,N4176,N4177,N4178,
  N4179,N4180,N4181,N4182,N4183,N4184,N4185,N4186,N4187,N4188,N4189,N4190,N4191,
  N4192,N4193,N4194,N4195,N4196,N4197,N4198,N4199,N4200,N4201,N4202,N4203,N4204,
  N4205,N4206,N4207,N4208,N4209,N4210,N4211,N4212,N4213,N4214,N4215,N4216,N4217,N4218,
  N4219,N4220,N4221,N4222,N4223,N4224,N4225,N4226,N4227,N4228,N4229,N4230,N4231,
  N4232,N4233,N4234,N4235,N4236,N4237,N4238,N4239,N4240,N4241,N4242,N4243,N4244,
  N4245,N4246,N4247,N4248,N4249,N4250,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,
  N4259,N4260,N4261,N4262,N4263,N4264,N4265,N4266,N4267,N4268,N4269,N4270,N4271,
  N4272,N4273,N4274,N4275,N4276,N4277,N4278,N4279,N4280,N4281,N4282,N4283,N4284,
  N4285,N4286,N4287,N4288,N4289,N4290,N4291,N4292,N4293,N4294,N4295,N4296,N4297,N4298,
  N4299,N4300,N4301,N4302,N4303,N4304,N4305,N4306,N4307,N4308,N4309,N4310,N4311,
  N4312,N4313,N4314,N4315,N4316,N4317,N4318,N4319,N4320,N4321,N4322,N4323,N4324,
  N4325,N4326,N4327,N4328,N4329,N4330,N4331,N4332,N4333,N4334,N4335,N4336,N4337,N4338,
  N4339,N4340,N4341,N4342,N4343,N4344,N4345,N4346,N4347,N4348,N4349,N4350,N4351,
  N4352,N4353,N4354,N4355,N4356,N4357,N4358,N4359,N4360,N4361,N4362,N4363,N4364,
  N4365,N4366,N4367,N4368,N4369,N4370,N4371,N4372,N4373,N4374,N4375,N4376,N4377,N4378,
  N4379,N4380,N4381,N4382,N4383,N4384,N4385,N4386,N4387,N4388,N4389,N4390,N4391,
  N4392,N4393,N4394,N4395,N4396,N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404,
  N4405,N4406,N4407,N4408,N4409,N4410,N4411,N4412,N4413,N4414,N4415,N4416,N4417,N4418,
  N4419,N4420,N4421,N4422,N4423,N4424,N4425,N4426,N4427,N4428,N4429,N4430,N4431,
  N4432,N4433,N4434,N4435,N4436,N4437,N4438,N4439,N4440,N4441,N4442,N4443,N4444,
  N4445,N4446,N4447,N4448,N4449,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457,N4458,
  N4459,N4460,N4461,N4462,N4463,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4471,
  N4472,N4473,N4474,N4475,N4476,N4477,N4478,N4479,N4480,N4481,N4482,N4483,N4484,
  N4485,N4486,N4487,N4488,N4489,N4490,N4491,N4492,N4493,N4494,N4495,N4496,N4497,N4498,
  N4499,N4500,N4501,N4502,N4503,N4504,N4505,N4506,N4507,N4508,N4509,N4510,N4511,
  N4512,N4513,N4514,N4515,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523,N4524,
  N4525,N4526,N4527,N4528,N4529,N4530,N4531,N4532,N4533,N4534,N4535,N4536,N4537,N4538,
  N4539,N4540,N4541,N4542,N4543,N4544,N4545,N4546,N4547,N4548,N4549,N4550,N4551,
  N4552,N4553,N4554,N4555,N4556,N4557,N4558,N4559,N4560,N4561,N4562,N4563,N4564,
  N4565,N4566,N4567,N4568,N4569,N4570,N4571,N4572,N4573,N4574,N4575,N4576,N4577,N4578,
  N4579,N4580,N4581,N4582,N4583,N4584,N4585,N4586,N4587,N4588,N4589,N4590,N4591,
  N4592,N4593,N4594,N4595,N4596,N4597,N4598,N4599,N4600,N4601,N4602,N4603,N4604,
  N4605,N4606,N4607,N4608,N4609,N4610,N4611,N4612,N4613,N4614,N4615,N4616,N4617,N4618,
  N4619,N4620,N4621,N4622,N4623,N4624,N4625,N4626,N4627,N4628,N4629,N4630,N4631,
  N4632,N4633,N4634,N4635,N4636,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644,
  N4645,N4646,N4647,N4648,N4649,N4650,N4651,N4652,N4653,N4654,N4655,N4656,N4657,N4658,
  N4659,N4660,N4661,N4662,N4663,N4664,N4665,N4666,N4667,N4668,N4669,N4670,N4671,
  N4672,N4673,N4674,N4675,N4676,N4677,N4678,N4679,N4680,N4681,N4682,N4683,N4684,
  N4685,N4686,N4687,N4688,N4689,N4690,N4691,N4692,N4693,N4694,N4695,N4696,N4697,N4698,
  N4699,N4700,N4701,N4702,N4703,N4704,N4705,N4706,N4707,N4708,N4709,N4710,N4711,
  N4712,N4713,N4714,N4715,N4716,N4717,N4718,N4719,N4720,N4721,N4722,N4723,N4724,
  N4725,N4726,N4727,N4728,N4729,N4730,N4731,N4732,N4733,N4734,N4735,N4736,N4737,N4738,
  N4739,N4740,N4741,N4742,N4743,N4744,N4745,N4746,N4747,N4748,N4749,N4750,N4751,
  N4752,N4753,N4754,N4755,N4756,N4757,N4758,N4759,N4760,N4761,N4762,N4763,N4764,
  N4765,N4766,N4767,N4768,N4769,N4770,N4771,N4772,N4773,N4774,N4775,N4776,N4777,N4778,
  N4779,N4780,N4781,N4782,N4783,N4784,N4785,N4786,N4787,N4788,N4789,N4790,N4791,
  N4792,N4793,N4794,N4795,N4796,N4797,N4798,N4799,N4800,N4801,N4802,N4803,N4804,
  N4805,N4806,N4807,N4808,N4809,N4810,N4811,N4812,N4813,N4814,N4815,N4816,N4817,N4818,
  N4819,N4820,N4821,N4822,N4823,N4824,N4825,N4826,N4827,N4828,N4829,N4830,N4831,
  N4832,N4833,N4834,N4835,N4836,N4837,N4838,N4839,N4840,N4841,N4842,N4843,N4844,
  N4845,N4846,N4847,N4848,N4849,N4850,N4851,N4852,N4853,N4854,N4855,N4856,N4857,N4858,
  N4859,N4860,N4861,N4862,N4863,N4864,N4865,N4866,N4867,N4868,N4869,N4870,N4871,
  N4872,N4873,N4874,N4875,N4876,N4877,N4878,N4879,N4880,N4881,N4882,N4883,N4884,
  N4885,N4886,N4887,N4888,N4889,N4890,N4891,N4892,N4893,N4894,N4895,N4896,N4897,N4898,
  N4899,N4900,N4901,N4902,N4903,N4904,N4905,N4906,N4907,N4908,N4909,N4910,N4911,
  N4912,N4913,N4914,N4915,N4916,N4917,N4918,N4919,N4920,N4921,N4922,N4923,N4924,
  N4925,N4926,N4927,N4928,N4929,N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937,N4938,
  N4939,N4940,N4941,N4942,N4943,N4944,N4945,N4946,N4947,N4948,N4949,N4950,N4951,
  N4952,N4953,N4954,N4955,N4956,N4957,N4958,N4959,N4960,N4961,N4962,N4963,N4964,
  N4965,N4966,N4967,N4968,N4969,N4970,N4971,N4972,N4973,N4974,N4975,N4976,N4977,N4978,
  N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4986,N4987,N4988,N4989,N4990,N4991,
  N4992,N4993,N4994,N4995,N4996,N4997,N4998,N4999,N5000,N5001,N5002,N5003,N5004,
  N5005,N5006,N5007,N5008,N5009,N5010,N5011,N5012,N5013,N5014,N5015,N5016,N5017,N5018,
  N5019,N5020,N5021,N5022,N5023,N5024,N5025,N5026,N5027,N5028,N5029,N5030,N5031,
  N5032,N5033,N5034,N5035,N5036,N5037,N5038,N5039,N5040,N5041,N5042,N5043,N5044,
  N5045,N5046,N5047,N5048,N5049,N5050,N5051,N5052,N5053,N5054,N5055,N5056,N5057,N5058,
  N5059,N5060,N5061,N5062,N5063,N5064,N5065,N5066,N5067,N5068,N5069,N5070,N5071,
  N5072,N5073,N5074,N5075,N5076,N5077,N5078,N5079,N5080,N5081,N5082,N5083,N5084,
  N5085,N5086,N5087,N5088,N5089,N5090,N5091,N5092,N5093,N5094,N5095,N5096,N5097,N5098,
  N5099,N5100,N5101,N5102,N5103,N5104,N5105,N5106,N5107,N5108,N5109,N5110,N5111,
  N5112,N5113,N5114,N5115,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123,N5124,
  N5125,N5126,N5127,N5128,N5129,N5130,N5131,N5132,N5133,N5134,N5135,N5136,N5137,N5138,
  N5139,N5140,N5141,N5142,N5143,N5144,N5145,N5146,N5147,N5148,N5149,N5150,N5151,
  N5152,N5153,N5154,N5155,N5156,N5157,N5158,N5159,N5160,N5161,N5162,N5163,N5164,
  N5165,N5166,N5167,N5168,N5169,N5170,N5171,N5172,N5173,N5174,N5175,N5176,N5177,N5178,
  N5179,N5180,N5181,N5182,N5183,N5184,N5185,N5186,N5187,N5188,N5189,N5190,N5191,
  N5192,N5193,N5194,N5195,N5196,N5197,N5198,N5199,N5200,N5201,N5202,N5203,N5204,
  N5205,N5206,N5207,N5208,N5209,N5210,N5211,N5212,N5213,N5214,N5215,N5216,N5217,N5218,
  N5219,N5220,N5221,N5222,N5223,N5224,N5225,N5226,N5227,N5228,N5229,N5230,N5231,
  N5232,N5233,N5234,N5235,N5236,N5237,N5238,N5239,N5240,N5241,N5242,N5243,N5244,
  N5245,N5246,N5247,N5248,N5249,N5250,N5251,N5252,N5253,N5254,N5255,N5256,N5257,N5258,
  N5259,N5260,N5261,N5262,N5263,N5264,N5265,N5266,N5267,N5268,N5269,N5270,N5271,
  N5272,N5273,N5274,N5275,N5276,N5277,N5278,N5279,N5280,N5281,N5282,N5283,N5284,
  N5285,N5286,N5287,N5288,N5289,N5290,N5291,N5292,N5293,N5294,N5295,N5296,N5297,N5298,
  N5299,N5300,N5301,N5302,N5303,N5304,N5305,N5306,N5307,N5308,N5309,N5310,N5311,
  N5312,N5313,N5314,N5315,N5316,N5317,N5318,N5319,N5320,N5321,N5322,N5323,N5324,
  N5325,N5326,N5327,N5328,N5329,N5330,N5331,N5332,N5333,N5334,N5335,N5336,N5337,N5338,
  N5339,N5340,N5341,N5342,N5343,N5344,N5345,N5346,N5347,N5348,N5349,N5350,N5351,
  N5352,N5353,N5354,N5355,N5356,N5357,N5358,N5359,N5360,N5361,N5362,N5363,N5364,
  N5365,N5366,N5367,N5368,N5369,N5370,N5371,N5372,N5373,N5374,N5375,N5376,N5377,N5378,
  N5379,N5380,N5381,N5382,N5383,N5384,N5385,N5386,N5387,N5388,N5389,N5390,N5391,
  N5392,N5393,N5394,N5395,N5396,N5397,N5398,N5399,N5400,N5401,N5402,N5403,N5404,
  N5405,N5406,N5407,N5408,N5409,N5410,N5411,N5412,N5413,N5414,N5415,N5416,N5417,N5418,
  N5419,N5420,N5421,N5422,N5423,N5424,N5425,N5426,N5427,N5428,N5429,N5430,N5431,
  N5432,N5433,N5434,N5435,N5436,N5437,N5438,N5439,N5440,N5441,N5442,N5443,N5444,
  N5445,N5446,N5447,N5448,N5449,N5450,N5451,N5452,N5453,N5454,N5455,N5456,N5457,N5458,
  N5459,N5460,N5461,N5462,N5463,N5464,N5465,N5466,N5467,N5468,N5469,N5470,N5471,
  N5472,N5473,N5474,N5475,N5476,N5477,N5478,N5479,N5480,N5481,N5482,N5483,N5484,
  N5485,N5486,N5487,N5488,N5489,N5490,N5491,N5492,N5493,N5494,N5495,N5496,N5497,N5498,
  N5499,N5500,N5501,N5502,N5503,N5504,N5505,N5506,N5507,N5508,N5509,N5510,N5511,
  N5512,N5513,N5514,N5515,N5516,N5517,N5518,N5519,N5520,N5521,N5522,N5523,N5524,
  N5525,N5526,N5527,N5528,N5529,N5530,N5531,N5532,N5533,N5534,N5535,N5536,N5537,N5538,
  N5539,N5540,N5541,N5542,N5543,N5544,N5545,N5546,N5547,N5548,N5549,N5550,N5551,
  N5552,N5553,N5554,N5555,N5556,N5557,N5558,N5559,N5560,N5561,N5562,N5563,N5564,
  N5565,N5566,N5567,N5568,N5569,N5570,N5571,N5572,N5573,N5574,N5575,N5576,N5577,N5578,
  N5579,N5580,N5581,N5582,N5583,N5584,N5585,N5586,N5587,N5588,N5589,N5590,N5591,
  N5592,N5593,N5594,N5595,N5596,N5597,N5598,N5599,N5600,N5601,N5602,N5603,N5604,
  N5605,N5606,N5607,N5608,N5609,N5610,N5611,N5612,N5613,N5614,N5615,N5616,N5617,N5618,
  N5619,N5620,N5621,N5622,N5623,N5624,N5625,N5626,N5627,N5628,N5629,N5630,N5631,
  N5632,N5633,N5634,N5635,N5636,N5637,N5638,N5639,N5640,N5641,N5642,N5643,N5644,
  N5645,N5646,N5647,N5648,N5649,N5650,N5651,N5652,N5653,N5654,N5655,N5656,N5657,N5658,
  N5659,N5660,N5661,N5662,N5663,N5664,N5665,N5666,N5667,N5668,N5669,N5670,N5671,
  N5672,N5673,N5674,N5675,N5676,N5677,N5678,N5679,N5680,N5681,N5682,N5683,N5684,
  N5685,N5686,N5687,N5688,N5689,N5690,N5691,N5692,N5693,N5694,N5695,N5696,N5697,N5698,
  N5699,N5700,N5701,N5702,N5703,N5704,N5705,N5706,N5707,N5708,N5709,N5710,N5711,
  N5712,N5713,N5714,N5715,N5716,N5717,N5718,N5719,N5720,N5721,N5722,N5723,N5724,
  N5725,N5726,N5727,N5728,N5729,N5730,N5731,N5732,N5733,N5734,N5735,N5736,N5737,N5738,
  N5739,N5740,N5741,N5742,N5743,N5744,N5745,N5746,N5747,N5748,N5749,N5750,N5751,
  N5752,N5753,N5754,N5755,N5756,N5757,N5758,N5759,N5760,N5761,N5762,N5763,N5764,
  N5765,N5766,N5767,N5768,N5769,N5770,N5771,N5772,N5773,N5774,N5775,N5776,N5777,N5778,
  N5779,N5780,N5781,N5782,N5783,N5784,N5785,N5786,N5787,N5788,N5789,N5790,N5791,
  N5792,N5793,N5794,N5795,N5796,N5797,N5798,N5799,N5800,N5801,N5802,N5803,N5804,
  N5805,N5806,N5807,N5808,N5809,N5810,N5811,N5812,N5813,N5814,N5815,N5816,N5817,N5818,
  N5819,N5820,N5821,N5822,N5823,N5824,N5825,N5826,N5827,N5828,N5829,N5830,N5831,
  N5832,N5833,N5834,N5835,N5836,N5837,N5838,N5839,N5840,N5841,N5842,N5843,N5844,
  N5845,N5846,N5847,N5848,N5849,N5850,N5851,N5852,N5853,N5854,N5855,N5856,N5857,N5858,
  N5859,N5860,N5861,N5862,N5863,N5864,N5865,N5866,N5867,N5868,N5869,N5870,N5871,
  N5872,N5873,N5874,N5875,N5876,N5877,N5878,N5879,N5880,N5881,N5882,N5883,N5884,
  N5885,N5886,N5887,N5888,N5889,N5890,N5891,N5892,N5893,N5894,N5895,N5896,N5897,N5898,
  N5899,N5900,N5901,N5902,N5903,N5904,N5905,N5906,N5907,N5908,N5909,N5910,N5911,
  N5912,N5913,N5914,N5915,N5916,N5917,N5918,N5919,N5920,N5921,N5922,N5923,N5924,
  N5925,N5926,N5927,N5928,N5929,N5930,N5931,N5932,N5933,N5934,N5935,N5936,N5937,N5938,
  N5939,N5940,N5941,N5942,N5943,N5944,N5945,N5946,N5947,N5948,N5949,N5950,N5951,
  N5952,N5953,N5954,N5955,N5956,N5957,N5958,N5959,N5960,N5961,N5962,N5963,N5964,
  N5965,N5966,N5967,N5968,N5969,N5970,N5971,N5972,N5973,N5974,N5975,N5976,N5977,N5978,
  N5979,N5980,N5981,N5982,N5983,N5984,N5985,N5986,N5987,N5988,N5989,N5990,N5991,
  N5992,N5993,N5994,N5995,N5996,N5997,N5998,N5999,N6000,N6001,N6002,N6003,N6004,
  N6005,N6006,N6007,N6008,N6009,N6010,N6011,N6012,N6013,N6014,N6015,N6016,N6017,N6018,
  N6019,N6020,N6021,N6022,N6023,N6024,N6025,N6026,N6027,N6028,N6029,N6030,N6031,
  N6032,N6033,N6034,N6035,N6036,N6037,N6038,N6039,N6040,N6041,N6042,N6043,N6044,
  N6045,N6046,N6047,N6048,N6049,N6050,N6051,N6052,N6053,N6054,N6055,N6056,N6057,N6058,
  N6059,N6060,N6061,N6062,N6063,N6064,N6065,N6066,N6067,N6068,N6069,N6070,N6071,
  N6072,N6073,N6074,N6075,N6076,N6077,N6078,N6079,N6080,N6081,N6082,N6083,N6084,
  N6085,N6086,N6087,N6088,N6089,N6090,N6091,N6092,N6093,N6094,N6095,N6096,N6097,N6098,
  N6099,N6100,N6101,N6102,N6103,N6104,N6105,N6106,N6107,N6108,N6109,N6110,N6111,
  N6112,N6113,N6114,N6115,N6116,N6117,N6118,N6119,N6120,N6121,N6122,N6123,N6124,
  N6125,N6126,N6127,N6128,N6129,N6130,N6131,N6132,N6133,N6134,N6135,N6136,N6137,N6138,
  N6139,N6140,N6141,N6142,N6143,N6144,N6145,N6146,N6147,N6148,N6149,N6150,N6151,
  N6152,N6153,N6154,N6155,N6156,N6157,N6158,N6159,N6160,N6161,N6162,N6163,N6164,
  N6165,N6166,N6167,N6168,N6169,N6170,N6171,N6172,N6173,N6174,N6175,N6176,N6177,N6178,
  N6179,N6180,N6181,N6182,N6183,N6184,N6185,N6186,N6187,N6188,N6189,N6190,N6191,
  N6192,N6193,N6194,N6195,N6196,N6197,N6198,N6199,N6200,N6201,N6202,N6203,N6204,
  N6205,N6206,N6207,N6208,N6209,N6210,N6211,N6212,N6213,N6214,N6215,N6216,N6217,N6218,
  N6219,N6220,N6221,N6222,N6223,N6224,N6225,N6226,N6227,N6228,N6229,N6230,N6231,
  N6232,N6233,N6234,N6235,N6236,N6237,N6238,N6239,N6240,N6241,N6242,N6243,N6244,
  N6245,N6246,N6247,N6248,N6249,N6250,N6251,N6252,N6253,N6254,N6255,N6256,N6257,N6258,
  N6259,N6260,N6261,N6262,N6263,N6264,N6265,N6266,N6267,N6268,N6269,N6270,N6271,
  N6272,N6273,N6274,N6275,N6276,N6277,N6278,N6279,N6280,N6281,N6282,N6283,N6284,
  N6285,N6286,N6287,N6288,N6289,N6290,N6291,N6292,N6293,N6294,N6295,N6296,N6297,N6298,
  N6299,N6300,N6301,N6302,N6303,N6304,N6305,N6306,N6307,N6308,N6309,N6310,N6311,
  N6312,N6313,N6314,N6315,N6316,N6317,N6318,N6319,N6320,N6321,N6322,N6323,N6324,
  N6325,N6326,N6327,N6328,N6329,N6330,N6331,N6332,N6333,N6334,N6335,N6336,N6337,N6338,
  N6339,N6340,N6341,N6342,N6343,N6344,N6345,N6346,N6347,N6348,N6349,N6350,N6351,
  N6352,N6353,N6354,N6355,N6356,N6357,N6358,N6359,N6360,N6361,N6362,N6363,N6364,
  N6365,N6366,N6367,N6368,N6369,N6370,N6371,N6372,N6373,N6374,N6375,N6376,N6377,N6378,
  N6379,N6380,N6381,N6382,N6383,N6384,N6385,N6386,N6387,N6388,N6389,N6390,N6391,
  N6392,N6393,N6394,N6395,N6396,N6397,N6398,N6399,N6400,N6401,N6402,N6403,N6404,
  N6405,N6406,N6407,N6408,N6409,N6410,N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6418,
  N6419,N6420,N6421,N6422,N6423,N6424,N6425,N6426,N6427,N6428,N6429,N6430,N6431,
  N6432,N6433,N6434,N6435,N6436,N6437,N6438,N6439,N6440,N6441,N6442,N6443,N6444,
  N6445,N6446,N6447,N6448,N6449,N6450,N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458,
  N6459,N6460,N6461,N6462,N6463,N6464,N6465,N6466,N6467,N6468,N6469,N6470,N6471,
  N6472,N6473,N6474,N6475,N6476,N6477,N6478,N6479,N6480,N6481,N6482,N6483,N6484,
  N6485,N6486,N6487,N6488,N6489,N6490,N6491,N6492,N6493,N6494,N6495,N6496,N6497,N6498,
  N6499,N6500,N6501,N6502,N6503,N6504,N6505,N6506,N6507,N6508,N6509,N6510,N6511,
  N6512,N6513,N6514,N6515,N6516,N6517,N6518,N6519,N6520,N6521,N6522,N6523,N6524,
  N6525,N6526,N6527,N6528,N6529,N6530,N6531,N6532,N6533,N6534,N6535,N6536,N6537,N6538,
  N6539,N6540,N6541,N6542,N6543,N6544,N6545,N6546,N6547,N6548,N6549,N6550,N6551,
  N6552,N6553,N6554,N6555,N6556,N6557,N6558,N6559,N6560,N6561,N6562,N6563,N6564,
  N6565,N6566,N6567,N6568,N6569,N6570,N6571,N6572,N6573,N6574,N6575,N6576,N6577,N6578,
  N6579,N6580,N6581,N6582,N6583,N6584,N6585,N6586,N6587,N6588,N6589,N6590,N6591,
  N6592,N6593,N6594,N6595,N6596,N6597,N6598,N6599,N6600,N6601,N6602,N6603,N6604,
  N6605,N6606,N6607,N6608,N6609,N6610,N6611,N6612,N6613,N6614,N6615,N6616,N6617,N6618,
  N6619,N6620,N6621,N6622,N6623,N6624,N6625,N6626,N6627,N6628,N6629,N6630,N6631,
  N6632,N6633,N6634,N6635,N6636,N6637,N6638,N6639,N6640,N6641,N6642,N6643,N6644,
  N6645,N6646,N6647,N6648,N6649,N6650,N6651,N6652,N6653,N6654,N6655,N6656,N6657,N6658,
  N6659,N6660,N6661,N6662,N6663,N6664,N6665,N6666,N6667,N6668,N6669,N6670,N6671,
  N6672,N6673,N6674,N6675,N6676,N6677,N6678,N6679,N6680,N6681,N6682,N6683,N6684,
  N6685,N6686,N6687,N6688,N6689,N6690,N6691,N6692,N6693,N6694,N6695,N6696,N6697,N6698,
  N6699,N6700,N6701,N6702,N6703,N6704,N6705,N6706,N6707,N6708,N6709,N6710,N6711,
  N6712,N6713,N6714,N6715,N6716,N6717,N6718,N6719,N6720,N6721,N6722,N6723,N6724,
  N6725,N6726,N6727,N6728,N6729,N6730,N6731,N6732,N6733,N6734,N6735,N6736,N6737,N6738,
  N6739,N6740,N6741,N6742,N6743,N6744,N6745,N6746,N6747,N6748,N6749,N6750,N6751,
  N6752,N6753,N6754,N6755,N6756,N6757,N6758,N6759,N6760,N6761,N6762,N6763,N6764,
  N6765,N6766,N6767,N6768,N6769,N6770,N6771,N6772,N6773,N6774,N6775,N6776,N6777,N6778,
  N6779,N6780,N6781,N6782,N6783,N6784,N6785,N6786,N6787,N6788,N6789,N6790,N6791,
  N6792,N6793,N6794,N6795,N6796,N6797,N6798,N6799,N6800,N6801,N6802,N6803,N6804,
  N6805,N6806,N6807,N6808,N6809,N6810,N6811,N6812,N6813,N6814,N6815,N6816,N6817,N6818,
  N6819,N6820,N6821,N6822,N6823,N6824,N6825,N6826,N6827,N6828,N6829,N6830,N6831,
  N6832,N6833,N6834,N6835,N6836,N6837,N6838,N6839,N6840,N6841,N6842,N6843,N6844,
  N6845,N6846,N6847,N6848,N6849,N6850,N6851,N6852,N6853,N6854,N6855,N6856,N6857,N6858,
  N6859,N6860,N6861,N6862,N6863,N6864,N6865,N6866,N6867,N6868,N6869,N6870,N6871,
  N6872,N6873,N6874,N6875,N6876,N6877,N6878,N6879,N6880,N6881,N6882,N6883,N6884,
  N6885,N6886,N6887,N6888,N6889,N6890,N6891,N6892,N6893,N6894,N6895,N6896,N6897,N6898,
  N6899,N6900,N6901,N6902,N6903,N6904,N6905,N6906,N6907,N6908,N6909,N6910,N6911,
  N6912,N6913,N6914,N6915,N6916,N6917,N6918,N6919,N6920,N6921,N6922,N6923,N6924,
  N6925,N6926,N6927,N6928,N6929,N6930,N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6938,
  N6939,N6940,N6941,N6942,N6943,N6944,N6945,N6946,N6947,N6948,N6949,N6950,N6951,
  N6952,N6953,N6954,N6955,N6956,N6957,N6958,N6959,N6960,N6961,N6962,N6963,N6964,
  N6965,N6966,N6967,N6968,N6969,N6970,N6971,N6972,N6973,N6974,N6975,N6976,N6977,N6978,
  N6979,N6980,N6981,N6982,N6983,N6984,N6985,N6986,N6987,N6988,N6989,N6990,N6991,
  N6992,N6993,N6994,N6995,N6996,N6997,N6998,N6999,N7000,N7001,N7002,N7003,N7004,
  N7005,N7006,N7007,N7008,N7009,N7010,N7011,N7012,N7013,N7014,N7015,N7016,N7017,N7018,
  N7019,N7020,N7021,N7022,N7023,N7024,N7025,N7026,N7027,N7028,N7029,N7030,N7031,
  N7032,N7033,N7034,N7035,N7036,N7037,N7038,N7039,N7040,N7041,N7042,N7043,N7044,
  N7045,N7046,N7047,N7048,N7049,N7050,N7051,N7052,N7053,N7054,N7055,N7056,N7057,N7058,
  N7059,N7060,N7061,N7062,N7063,N7064,N7065,N7066,N7067,N7068,N7069,N7070,N7071,
  N7072,N7073,N7074,N7075,N7076,N7077,N7078,N7079,N7080,N7081,N7082,N7083,N7084,
  N7085,N7086,N7087,N7088,N7089,N7090,N7091,N7092,N7093,N7094,N7095,N7096,N7097,N7098,
  N7099,N7100,N7101,N7102,N7103,N7104,N7105,N7106,N7107,N7108,N7109,N7110,N7111,
  N7112,N7113,N7114,N7115,N7116,N7117,N7118,N7119,N7120,N7121,N7122,N7123,N7124,
  N7125,N7126,N7127,N7128,N7129,N7130,N7131,N7132,N7133,N7134,N7135,N7136,N7137,N7138,
  N7139,N7140,N7141,N7142,N7143,N7144,N7145,N7146,N7147,N7148,N7149,N7150,N7151,
  N7152,N7153,N7154,N7155,N7156,N7157,N7158,N7159,N7160,N7161,N7162,N7163,N7164,
  N7165,N7166,N7167,N7168,N7169,N7170,N7171,N7172,N7173,N7174,N7175,N7176,N7177,N7178,
  N7179,N7180,N7181,N7182,N7183,N7184,N7185,N7186,N7187,N7188,N7189,N7190,N7191,
  N7192,N7193,N7194,N7195,N7196,N7197,N7198,N7199,N7200,N7201,N7202,N7203,N7204,
  N7205,N7206,N7207,N7208,N7209,N7210,N7211,N7212,N7213,N7214,N7215,N7216,N7217,N7218,
  N7219,N7220,N7221,N7222,N7223,N7224,N7225,N7226,N7227,N7228,N7229,N7230,N7231,
  N7232,N7233,N7234,N7235,N7236,N7237,N7238,N7239,N7240,N7241,N7242,N7243,N7244,
  N7245,N7246,N7247,N7248,N7249,N7250,N7251,N7252,N7253,N7254,N7255,N7256,N7257,N7258,
  N7259,N7260,N7261,N7262,N7263,N7264,N7265,N7266,N7267,N7268,N7269,N7270,N7271,
  N7272,N7273,N7274,N7275,N7276,N7277,N7278,N7279,N7280,N7281,N7282,N7283,N7284,
  N7285,N7286,N7287,N7288,N7289,N7290,N7291,N7292,N7293,N7294,N7295,N7296,N7297,N7298,
  N7299,N7300,N7301,N7302,N7303,N7304,N7305,N7306,N7307,N7308,N7309,N7310,N7311,
  N7312,N7313,N7314,N7315,N7316,N7317,N7318,N7319,N7320,N7321,N7322,N7323,N7324,
  N7325,N7326,N7327,N7328,N7329,N7330,N7331,N7332,N7333,N7334,N7335,N7336,N7337,N7338,
  N7339,N7340,N7341,N7342,N7343,N7344,N7345,N7346,N7347,N7348,N7349,N7350,N7351,
  N7352,N7353,N7354,N7355,N7356,N7357,N7358,N7359,N7360,N7361,N7362,N7363,N7364,
  N7365,N7366,N7367,N7368,N7369,N7370,N7371,N7372,N7373,N7374,N7375,N7376,N7377,N7378,
  N7379,N7380,N7381,N7382,N7383,N7384,N7385,N7386,N7387,N7388,N7389,N7390,N7391,
  N7392,N7393,N7394,N7395,N7396,N7397,N7398,N7399,N7400,N7401,N7402,N7403,N7404,
  N7405,N7406,N7407,N7408,N7409,N7410,N7411,N7412,N7413,N7414,N7415,N7416,N7417,N7418,
  N7419,N7420,N7421,N7422,N7423,N7424,N7425,N7426,N7427,N7428,N7429,N7430,N7431,
  N7432,N7433,N7434,N7435,N7436,N7437,N7438,N7439,N7440,N7441,N7442,N7443,N7444,
  N7445,N7446,N7447,N7448,N7449,N7450,N7451,N7452,N7453,N7454,N7455,N7456,N7457,N7458,
  N7459,N7460,N7461,N7462,N7463,N7464,N7465,N7466,N7467,N7468,N7469,N7470,N7471,
  N7472,N7473,N7474,N7475,N7476,N7477,N7478,N7479,N7480,N7481,N7482,N7483,N7484,
  N7485,N7486,N7487,N7488,N7489,N7490,N7491,N7492,N7493,N7494,N7495,N7496,N7497,N7498,
  N7499,N7500,N7501,N7502,N7503,N7504,N7505,N7506,N7507,N7508,N7509,N7510,N7511,
  N7512,N7513,N7514,N7515,N7516,N7517,N7518,N7519,N7520,N7521,N7522,N7523,N7524,
  N7525,N7526,N7527,N7528,N7529,N7530,N7531,N7532,N7533,N7534,N7535,N7536,N7537,N7538,
  N7539,N7540,N7541,N7542,N7543,N7544,N7545,N7546,N7547,N7548,N7549,N7550,N7551,
  N7552,N7553,N7554,N7555,N7556,N7557,N7558,N7559,N7560,N7561,N7562,N7563,N7564,
  N7565,N7566,N7567,N7568,N7569,N7570,N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578,
  N7579,N7580,N7581,N7582,N7583,N7584,N7585,N7586,N7587,N7588,N7589,N7590,N7591,
  N7592,N7593,N7594,N7595,N7596,N7597,N7598,N7599,N7600,N7601,N7602,N7603,N7604,
  N7605,N7606,N7607,N7608,N7609,N7610,N7611,N7612,N7613,N7614,N7615,N7616,N7617,N7618,
  N7619,N7620,N7621,N7622,N7623,N7624,N7625,N7626,N7627,N7628,N7629,N7630,N7631,
  N7632,N7633,N7634,N7635,N7636,N7637,N7638,N7639,N7640,N7641,N7642,N7643,N7644,
  N7645,N7646,N7647,N7648,N7649,N7650,N7651,N7652,N7653,N7654,N7655,N7656,N7657,N7658,
  N7659,N7660,N7661,N7662,N7663,N7664,N7665,N7666,N7667,N7668,N7669,N7670,N7671,
  N7672,N7673,N7674,N7675,N7676,N7677,N7678,N7679,N7680,N7681,N7682,N7683,N7684,
  N7685,N7686,N7687,N7688,N7689,N7690,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698,
  N7699,N7700,N7701,N7702,N7703,N7704,N7705,N7706,N7707,N7708,N7709,N7710,N7711,
  N7712,N7713,N7714,N7715,N7716,N7717,N7718,N7719,N7720,N7721,N7722,N7723,N7724,
  N7725,N7726,N7727,N7728,N7729,N7730,N7731,N7732,N7733,N7734,N7735,N7736,N7737,N7738,
  N7739,N7740,N7741,N7742,N7743,N7744,N7745,N7746,N7747,N7748,N7749,N7750,N7751,
  N7752,N7753,N7754,N7755,N7756,N7757,N7758,N7759,N7760,N7761,N7762,N7763,N7764,
  N7765,N7766,N7767,N7768,N7769,N7770,N7771,N7772,N7773,N7774,N7775,N7776,N7777,N7778,
  N7779,N7780,N7781,N7782,N7783,N7784,N7785,N7786,N7787,N7788,N7789,N7790,N7791,
  N7792,N7793,N7794,N7795,N7796,N7797,N7798,N7799,N7800,N7801,N7802,N7803,N7804,
  N7805,N7806,N7807,N7808,N7809,N7810,N7811,N7812,N7813,N7814,N7815,N7816,N7817,N7818,
  N7819,N7820,N7821,N7822,N7823,N7824,N7825,N7826,N7827,N7828,N7829,N7830,N7831,
  N7832,N7833,N7834,N7835,N7836,N7837,N7838,N7839,N7840,N7841,N7842,N7843,N7844,
  N7845,N7846,N7847,N7848,N7849,N7850,N7851,N7852,N7853,N7854,N7855,N7856,N7857,N7858,
  N7859,N7860,N7861,N7862,N7863,N7864,N7865,N7866,N7867,N7868,N7869,N7870,N7871,
  N7872,N7873,N7874,N7875,N7876,N7877,N7878,N7879,N7880,N7881,N7882,N7883,N7884,
  N7885,N7886,N7887,N7888,N7889,N7890,N7891,N7892,N7893,N7894,N7895,N7896,N7897,N7898,
  N7899,N7900,N7901,N7902,N7903,N7904,N7905,N7906,N7907,N7908,N7909,N7910,N7911,
  N7912,N7913,N7914,N7915,N7916,N7917,N7918,N7919,N7920,N7921,N7922,N7923,N7924,
  N7925,N7926,N7927,N7928,N7929,N7930,N7931,N7932,N7933,N7934,N7935,N7936,N7937,N7938,
  N7939,N7940,N7941,N7942,N7943,N7944,N7945,N7946,N7947,N7948,N7949,N7950,N7951,
  N7952,N7953,N7954,N7955,N7956,N7957,N7958,N7959,N7960,N7961,N7962,N7963,N7964,
  N7965,N7966,N7967,N7968,N7969,N7970,N7971,N7972,N7973,N7974,N7975,N7976,N7977,N7978,
  N7979,N7980,N7981,N7982,N7983,N7984,N7985,N7986,N7987,N7988,N7989,N7990,N7991,
  N7992,N7993,N7994,N7995,N7996,N7997,N7998,N7999,N8000,N8001,N8002,N8003,N8004,
  N8005,N8006,N8007,N8008,N8009,N8010,N8011,N8012,N8013,N8014,N8015,N8016,N8017,N8018,
  N8019,N8020,N8021,N8022,N8023,N8024,N8025,N8026,N8027,N8028,N8029,N8030,N8031,
  N8032,N8033,N8034,N8035,N8036,N8037,N8038,N8039,N8040,N8041,N8042,N8043,N8044,
  N8045,N8046,N8047,N8048,N8049,N8050,N8051,N8052,N8053,N8054,N8055,N8056,N8057,N8058,
  N8059,N8060,N8061,N8062,N8063,N8064,N8065,N8066,N8067,N8068,N8069,N8070,N8071,
  N8072,N8073,N8074,N8075,N8076,N8077,N8078,N8079,N8080,N8081,N8082,N8083,N8084,
  N8085,N8086,N8087,N8088,N8089,N8090,N8091,N8092,N8093,N8094,N8095,N8096,N8097,N8098,
  N8099,N8100,N8101,N8102,N8103,N8104,N8105,N8106,N8107,N8108,N8109,N8110,N8111,
  N8112,N8113,N8114,N8115,N8116,N8117,N8118,N8119,N8120,N8121,N8122,N8123,N8124,
  N8125,N8126,N8127,N8128,N8129,N8130,N8131,N8132,N8133,N8134,N8135,N8136,N8137,N8138,
  N8139,N8140,N8141,N8142,N8143,N8144,N8145,N8146,N8147,N8148,N8149,N8150,N8151,
  N8152,N8153,N8154,N8155,N8156,N8157,N8158,N8159,N8160,N8161,N8162,N8163,N8164,
  N8165,N8166,N8167,N8168,N8169,N8170,N8171,N8172,N8173,N8174,N8175,N8176,N8177,N8178,
  N8179,N8180,N8181,N8182,N8183,N8184,N8185,N8186,N8187,N8188,N8189,N8190,N8191,
  N8192,N8193,N8194,N8195,N8196,N8197,N8198,N8199,N8200,N8201,N8202,N8203,N8204,
  N8205,N8206,N8207,N8208,N8209,N8210,N8211,N8212,N8213,N8214,N8215,N8216,N8217,N8218,
  N8219,N8220,N8221,N8222,N8223,N8224,N8225,N8226,N8227,N8228,N8229,N8230,N8231,
  N8232,N8233,N8234,N8235,N8236,N8237,N8238,N8239,N8240,N8241,N8242,N8243,N8244,
  N8245,N8246,N8247,N8248,N8249,N8250,N8251,N8252,N8253,N8254,N8255,N8256,N8257,N8258,
  N8259,N8260,N8261,N8262,N8263,N8264,N8265,N8266,N8267,N8268,N8269,N8270,N8271,
  N8272,N8273,N8274,N8275,N8276,N8277,N8278,N8279,N8280,N8281,N8282,N8283,N8284,
  N8285,N8286,N8287,N8288,N8289,N8290,N8291,N8292,N8293,N8294,N8295,N8296,N8297,N8298,
  N8299,N8300,N8301,N8302,N8303,N8304,N8305,N8306,N8307,N8308,N8309,N8310,N8311,
  N8312,N8313,N8314,N8315,N8316,N8317,N8318,N8319,N8320,N8321,N8322,N8323,N8324;
  wire [1023:0] match_array,empty_array;
  reg [32767:0] mem;
  reg [1023:0] valid;
  assign N3105 = mem[32767:32736] == r_data_i;
  assign N3106 = mem[32735:32704] == r_data_i;
  assign N3107 = mem[32703:32672] == r_data_i;
  assign N3108 = mem[32671:32640] == r_data_i;
  assign N3109 = mem[32639:32608] == r_data_i;
  assign N3110 = mem[32607:32576] == r_data_i;
  assign N3111 = mem[32575:32544] == r_data_i;
  assign N3112 = mem[32543:32512] == r_data_i;
  assign N3113 = mem[32511:32480] == r_data_i;
  assign N3114 = mem[32479:32448] == r_data_i;
  assign N3115 = mem[32447:32416] == r_data_i;
  assign N3116 = mem[32415:32384] == r_data_i;
  assign N3117 = mem[32383:32352] == r_data_i;
  assign N3118 = mem[32351:32320] == r_data_i;
  assign N3119 = mem[32319:32288] == r_data_i;
  assign N3120 = mem[32287:32256] == r_data_i;
  assign N3121 = mem[32255:32224] == r_data_i;
  assign N3122 = mem[32223:32192] == r_data_i;
  assign N3123 = mem[32191:32160] == r_data_i;
  assign N3124 = mem[32159:32128] == r_data_i;
  assign N3125 = mem[32127:32096] == r_data_i;
  assign N3126 = mem[32095:32064] == r_data_i;
  assign N3127 = mem[32063:32032] == r_data_i;
  assign N3128 = mem[32031:32000] == r_data_i;
  assign N3129 = mem[31999:31968] == r_data_i;
  assign N3130 = mem[31967:31936] == r_data_i;
  assign N3131 = mem[31935:31904] == r_data_i;
  assign N3132 = mem[31903:31872] == r_data_i;
  assign N3133 = mem[31871:31840] == r_data_i;
  assign N3134 = mem[31839:31808] == r_data_i;
  assign N3135 = mem[31807:31776] == r_data_i;
  assign N3136 = mem[31775:31744] == r_data_i;
  assign N3137 = mem[31743:31712] == r_data_i;
  assign N3138 = mem[31711:31680] == r_data_i;
  assign N3139 = mem[31679:31648] == r_data_i;
  assign N3140 = mem[31647:31616] == r_data_i;
  assign N3141 = mem[31615:31584] == r_data_i;
  assign N3142 = mem[31583:31552] == r_data_i;
  assign N3143 = mem[31551:31520] == r_data_i;
  assign N3144 = mem[31519:31488] == r_data_i;
  assign N3145 = mem[31487:31456] == r_data_i;
  assign N3146 = mem[31455:31424] == r_data_i;
  assign N3147 = mem[31423:31392] == r_data_i;
  assign N3148 = mem[31391:31360] == r_data_i;
  assign N3149 = mem[31359:31328] == r_data_i;
  assign N3150 = mem[31327:31296] == r_data_i;
  assign N3151 = mem[31295:31264] == r_data_i;
  assign N3152 = mem[31263:31232] == r_data_i;
  assign N3153 = mem[31231:31200] == r_data_i;
  assign N3154 = mem[31199:31168] == r_data_i;
  assign N3155 = mem[31167:31136] == r_data_i;
  assign N3156 = mem[31135:31104] == r_data_i;
  assign N3157 = mem[31103:31072] == r_data_i;
  assign N3158 = mem[31071:31040] == r_data_i;
  assign N3159 = mem[31039:31008] == r_data_i;
  assign N3160 = mem[31007:30976] == r_data_i;
  assign N3161 = mem[30975:30944] == r_data_i;
  assign N3162 = mem[30943:30912] == r_data_i;
  assign N3163 = mem[30911:30880] == r_data_i;
  assign N3164 = mem[30879:30848] == r_data_i;
  assign N3165 = mem[30847:30816] == r_data_i;
  assign N3166 = mem[30815:30784] == r_data_i;
  assign N3167 = mem[30783:30752] == r_data_i;
  assign N3168 = mem[30751:30720] == r_data_i;
  assign N3169 = mem[30719:30688] == r_data_i;
  assign N3170 = mem[30687:30656] == r_data_i;
  assign N3171 = mem[30655:30624] == r_data_i;
  assign N3172 = mem[30623:30592] == r_data_i;
  assign N3173 = mem[30591:30560] == r_data_i;
  assign N3174 = mem[30559:30528] == r_data_i;
  assign N3175 = mem[30527:30496] == r_data_i;
  assign N3176 = mem[30495:30464] == r_data_i;
  assign N3177 = mem[30463:30432] == r_data_i;
  assign N3178 = mem[30431:30400] == r_data_i;
  assign N3179 = mem[30399:30368] == r_data_i;
  assign N3180 = mem[30367:30336] == r_data_i;
  assign N3181 = mem[30335:30304] == r_data_i;
  assign N3182 = mem[30303:30272] == r_data_i;
  assign N3183 = mem[30271:30240] == r_data_i;
  assign N3184 = mem[30239:30208] == r_data_i;
  assign N3185 = mem[30207:30176] == r_data_i;
  assign N3186 = mem[30175:30144] == r_data_i;
  assign N3187 = mem[30143:30112] == r_data_i;
  assign N3188 = mem[30111:30080] == r_data_i;
  assign N3189 = mem[30079:30048] == r_data_i;
  assign N3190 = mem[30047:30016] == r_data_i;
  assign N3191 = mem[30015:29984] == r_data_i;
  assign N3192 = mem[29983:29952] == r_data_i;
  assign N3193 = mem[29951:29920] == r_data_i;
  assign N3194 = mem[29919:29888] == r_data_i;
  assign N3195 = mem[29887:29856] == r_data_i;
  assign N3196 = mem[29855:29824] == r_data_i;
  assign N3197 = mem[29823:29792] == r_data_i;
  assign N3198 = mem[29791:29760] == r_data_i;
  assign N3199 = mem[29759:29728] == r_data_i;
  assign N3200 = mem[29727:29696] == r_data_i;
  assign N3201 = mem[29695:29664] == r_data_i;
  assign N3202 = mem[29663:29632] == r_data_i;
  assign N3203 = mem[29631:29600] == r_data_i;
  assign N3204 = mem[29599:29568] == r_data_i;
  assign N3205 = mem[29567:29536] == r_data_i;
  assign N3206 = mem[29535:29504] == r_data_i;
  assign N3207 = mem[29503:29472] == r_data_i;
  assign N3208 = mem[29471:29440] == r_data_i;
  assign N3209 = mem[29439:29408] == r_data_i;
  assign N3210 = mem[29407:29376] == r_data_i;
  assign N3211 = mem[29375:29344] == r_data_i;
  assign N3212 = mem[29343:29312] == r_data_i;
  assign N3213 = mem[29311:29280] == r_data_i;
  assign N3214 = mem[29279:29248] == r_data_i;
  assign N3215 = mem[29247:29216] == r_data_i;
  assign N3216 = mem[29215:29184] == r_data_i;
  assign N3217 = mem[29183:29152] == r_data_i;
  assign N3218 = mem[29151:29120] == r_data_i;
  assign N3219 = mem[29119:29088] == r_data_i;
  assign N3220 = mem[29087:29056] == r_data_i;
  assign N3221 = mem[29055:29024] == r_data_i;
  assign N3222 = mem[29023:28992] == r_data_i;
  assign N3223 = mem[28991:28960] == r_data_i;
  assign N3224 = mem[28959:28928] == r_data_i;
  assign N3225 = mem[28927:28896] == r_data_i;
  assign N3226 = mem[28895:28864] == r_data_i;
  assign N3227 = mem[28863:28832] == r_data_i;
  assign N3228 = mem[28831:28800] == r_data_i;
  assign N3229 = mem[28799:28768] == r_data_i;
  assign N3230 = mem[28767:28736] == r_data_i;
  assign N3231 = mem[28735:28704] == r_data_i;
  assign N3232 = mem[28703:28672] == r_data_i;
  assign N3233 = mem[28671:28640] == r_data_i;
  assign N3234 = mem[28639:28608] == r_data_i;
  assign N3235 = mem[28607:28576] == r_data_i;
  assign N3236 = mem[28575:28544] == r_data_i;
  assign N3237 = mem[28543:28512] == r_data_i;
  assign N3238 = mem[28511:28480] == r_data_i;
  assign N3239 = mem[28479:28448] == r_data_i;
  assign N3240 = mem[28447:28416] == r_data_i;
  assign N3241 = mem[28415:28384] == r_data_i;
  assign N3242 = mem[28383:28352] == r_data_i;
  assign N3243 = mem[28351:28320] == r_data_i;
  assign N3244 = mem[28319:28288] == r_data_i;
  assign N3245 = mem[28287:28256] == r_data_i;
  assign N3246 = mem[28255:28224] == r_data_i;
  assign N3247 = mem[28223:28192] == r_data_i;
  assign N3248 = mem[28191:28160] == r_data_i;
  assign N3249 = mem[28159:28128] == r_data_i;
  assign N3250 = mem[28127:28096] == r_data_i;
  assign N3251 = mem[28095:28064] == r_data_i;
  assign N3252 = mem[28063:28032] == r_data_i;
  assign N3253 = mem[28031:28000] == r_data_i;
  assign N3254 = mem[27999:27968] == r_data_i;
  assign N3255 = mem[27967:27936] == r_data_i;
  assign N3256 = mem[27935:27904] == r_data_i;
  assign N3257 = mem[27903:27872] == r_data_i;
  assign N3258 = mem[27871:27840] == r_data_i;
  assign N3259 = mem[27839:27808] == r_data_i;
  assign N3260 = mem[27807:27776] == r_data_i;
  assign N3261 = mem[27775:27744] == r_data_i;
  assign N3262 = mem[27743:27712] == r_data_i;
  assign N3263 = mem[27711:27680] == r_data_i;
  assign N3264 = mem[27679:27648] == r_data_i;
  assign N3265 = mem[27647:27616] == r_data_i;
  assign N3266 = mem[27615:27584] == r_data_i;
  assign N3267 = mem[27583:27552] == r_data_i;
  assign N3268 = mem[27551:27520] == r_data_i;
  assign N3269 = mem[27519:27488] == r_data_i;
  assign N3270 = mem[27487:27456] == r_data_i;
  assign N3271 = mem[27455:27424] == r_data_i;
  assign N3272 = mem[27423:27392] == r_data_i;
  assign N3273 = mem[27391:27360] == r_data_i;
  assign N3274 = mem[27359:27328] == r_data_i;
  assign N3275 = mem[27327:27296] == r_data_i;
  assign N3276 = mem[27295:27264] == r_data_i;
  assign N3277 = mem[27263:27232] == r_data_i;
  assign N3278 = mem[27231:27200] == r_data_i;
  assign N3279 = mem[27199:27168] == r_data_i;
  assign N3280 = mem[27167:27136] == r_data_i;
  assign N3281 = mem[27135:27104] == r_data_i;
  assign N3282 = mem[27103:27072] == r_data_i;
  assign N3283 = mem[27071:27040] == r_data_i;
  assign N3284 = mem[27039:27008] == r_data_i;
  assign N3285 = mem[27007:26976] == r_data_i;
  assign N3286 = mem[26975:26944] == r_data_i;
  assign N3287 = mem[26943:26912] == r_data_i;
  assign N3288 = mem[26911:26880] == r_data_i;
  assign N3289 = mem[26879:26848] == r_data_i;
  assign N3290 = mem[26847:26816] == r_data_i;
  assign N3291 = mem[26815:26784] == r_data_i;
  assign N3292 = mem[26783:26752] == r_data_i;
  assign N3293 = mem[26751:26720] == r_data_i;
  assign N3294 = mem[26719:26688] == r_data_i;
  assign N3295 = mem[26687:26656] == r_data_i;
  assign N3296 = mem[26655:26624] == r_data_i;
  assign N3297 = mem[26623:26592] == r_data_i;
  assign N3298 = mem[26591:26560] == r_data_i;
  assign N3299 = mem[26559:26528] == r_data_i;
  assign N3300 = mem[26527:26496] == r_data_i;
  assign N3301 = mem[26495:26464] == r_data_i;
  assign N3302 = mem[26463:26432] == r_data_i;
  assign N3303 = mem[26431:26400] == r_data_i;
  assign N3304 = mem[26399:26368] == r_data_i;
  assign N3305 = mem[26367:26336] == r_data_i;
  assign N3306 = mem[26335:26304] == r_data_i;
  assign N3307 = mem[26303:26272] == r_data_i;
  assign N3308 = mem[26271:26240] == r_data_i;
  assign N3309 = mem[26239:26208] == r_data_i;
  assign N3310 = mem[26207:26176] == r_data_i;
  assign N3311 = mem[26175:26144] == r_data_i;
  assign N3312 = mem[26143:26112] == r_data_i;
  assign N3313 = mem[26111:26080] == r_data_i;
  assign N3314 = mem[26079:26048] == r_data_i;
  assign N3315 = mem[26047:26016] == r_data_i;
  assign N3316 = mem[26015:25984] == r_data_i;
  assign N3317 = mem[25983:25952] == r_data_i;
  assign N3318 = mem[25951:25920] == r_data_i;
  assign N3319 = mem[25919:25888] == r_data_i;
  assign N3320 = mem[25887:25856] == r_data_i;
  assign N3321 = mem[25855:25824] == r_data_i;
  assign N3322 = mem[25823:25792] == r_data_i;
  assign N3323 = mem[25791:25760] == r_data_i;
  assign N3324 = mem[25759:25728] == r_data_i;
  assign N3325 = mem[25727:25696] == r_data_i;
  assign N3326 = mem[25695:25664] == r_data_i;
  assign N3327 = mem[25663:25632] == r_data_i;
  assign N3328 = mem[25631:25600] == r_data_i;
  assign N3329 = mem[25599:25568] == r_data_i;
  assign N3330 = mem[25567:25536] == r_data_i;
  assign N3331 = mem[25535:25504] == r_data_i;
  assign N3332 = mem[25503:25472] == r_data_i;
  assign N3333 = mem[25471:25440] == r_data_i;
  assign N3334 = mem[25439:25408] == r_data_i;
  assign N3335 = mem[25407:25376] == r_data_i;
  assign N3336 = mem[25375:25344] == r_data_i;
  assign N3337 = mem[25343:25312] == r_data_i;
  assign N3338 = mem[25311:25280] == r_data_i;
  assign N3339 = mem[25279:25248] == r_data_i;
  assign N3340 = mem[25247:25216] == r_data_i;
  assign N3341 = mem[25215:25184] == r_data_i;
  assign N3342 = mem[25183:25152] == r_data_i;
  assign N3343 = mem[25151:25120] == r_data_i;
  assign N3344 = mem[25119:25088] == r_data_i;
  assign N3345 = mem[25087:25056] == r_data_i;
  assign N3346 = mem[25055:25024] == r_data_i;
  assign N3347 = mem[25023:24992] == r_data_i;
  assign N3348 = mem[24991:24960] == r_data_i;
  assign N3349 = mem[24959:24928] == r_data_i;
  assign N3350 = mem[24927:24896] == r_data_i;
  assign N3351 = mem[24895:24864] == r_data_i;
  assign N3352 = mem[24863:24832] == r_data_i;
  assign N3353 = mem[24831:24800] == r_data_i;
  assign N3354 = mem[24799:24768] == r_data_i;
  assign N3355 = mem[24767:24736] == r_data_i;
  assign N3356 = mem[24735:24704] == r_data_i;
  assign N3357 = mem[24703:24672] == r_data_i;
  assign N3358 = mem[24671:24640] == r_data_i;
  assign N3359 = mem[24639:24608] == r_data_i;
  assign N3360 = mem[24607:24576] == r_data_i;
  assign N3361 = mem[24575:24544] == r_data_i;
  assign N3362 = mem[24543:24512] == r_data_i;
  assign N3363 = mem[24511:24480] == r_data_i;
  assign N3364 = mem[24479:24448] == r_data_i;
  assign N3365 = mem[24447:24416] == r_data_i;
  assign N3366 = mem[24415:24384] == r_data_i;
  assign N3367 = mem[24383:24352] == r_data_i;
  assign N3368 = mem[24351:24320] == r_data_i;
  assign N3369 = mem[24319:24288] == r_data_i;
  assign N3370 = mem[24287:24256] == r_data_i;
  assign N3371 = mem[24255:24224] == r_data_i;
  assign N3372 = mem[24223:24192] == r_data_i;
  assign N3373 = mem[24191:24160] == r_data_i;
  assign N3374 = mem[24159:24128] == r_data_i;
  assign N3375 = mem[24127:24096] == r_data_i;
  assign N3376 = mem[24095:24064] == r_data_i;
  assign N3377 = mem[24063:24032] == r_data_i;
  assign N3378 = mem[24031:24000] == r_data_i;
  assign N3379 = mem[23999:23968] == r_data_i;
  assign N3380 = mem[23967:23936] == r_data_i;
  assign N3381 = mem[23935:23904] == r_data_i;
  assign N3382 = mem[23903:23872] == r_data_i;
  assign N3383 = mem[23871:23840] == r_data_i;
  assign N3384 = mem[23839:23808] == r_data_i;
  assign N3385 = mem[23807:23776] == r_data_i;
  assign N3386 = mem[23775:23744] == r_data_i;
  assign N3387 = mem[23743:23712] == r_data_i;
  assign N3388 = mem[23711:23680] == r_data_i;
  assign N3389 = mem[23679:23648] == r_data_i;
  assign N3390 = mem[23647:23616] == r_data_i;
  assign N3391 = mem[23615:23584] == r_data_i;
  assign N3392 = mem[23583:23552] == r_data_i;
  assign N3393 = mem[23551:23520] == r_data_i;
  assign N3394 = mem[23519:23488] == r_data_i;
  assign N3395 = mem[23487:23456] == r_data_i;
  assign N3396 = mem[23455:23424] == r_data_i;
  assign N3397 = mem[23423:23392] == r_data_i;
  assign N3398 = mem[23391:23360] == r_data_i;
  assign N3399 = mem[23359:23328] == r_data_i;
  assign N3400 = mem[23327:23296] == r_data_i;
  assign N3401 = mem[23295:23264] == r_data_i;
  assign N3402 = mem[23263:23232] == r_data_i;
  assign N3403 = mem[23231:23200] == r_data_i;
  assign N3404 = mem[23199:23168] == r_data_i;
  assign N3405 = mem[23167:23136] == r_data_i;
  assign N3406 = mem[23135:23104] == r_data_i;
  assign N3407 = mem[23103:23072] == r_data_i;
  assign N3408 = mem[23071:23040] == r_data_i;
  assign N3409 = mem[23039:23008] == r_data_i;
  assign N3410 = mem[23007:22976] == r_data_i;
  assign N3411 = mem[22975:22944] == r_data_i;
  assign N3412 = mem[22943:22912] == r_data_i;
  assign N3413 = mem[22911:22880] == r_data_i;
  assign N3414 = mem[22879:22848] == r_data_i;
  assign N3415 = mem[22847:22816] == r_data_i;
  assign N3416 = mem[22815:22784] == r_data_i;
  assign N3417 = mem[22783:22752] == r_data_i;
  assign N3418 = mem[22751:22720] == r_data_i;
  assign N3419 = mem[22719:22688] == r_data_i;
  assign N3420 = mem[22687:22656] == r_data_i;
  assign N3421 = mem[22655:22624] == r_data_i;
  assign N3422 = mem[22623:22592] == r_data_i;
  assign N3423 = mem[22591:22560] == r_data_i;
  assign N3424 = mem[22559:22528] == r_data_i;
  assign N3425 = mem[22527:22496] == r_data_i;
  assign N3426 = mem[22495:22464] == r_data_i;
  assign N3427 = mem[22463:22432] == r_data_i;
  assign N3428 = mem[22431:22400] == r_data_i;
  assign N3429 = mem[22399:22368] == r_data_i;
  assign N3430 = mem[22367:22336] == r_data_i;
  assign N3431 = mem[22335:22304] == r_data_i;
  assign N3432 = mem[22303:22272] == r_data_i;
  assign N3433 = mem[22271:22240] == r_data_i;
  assign N3434 = mem[22239:22208] == r_data_i;
  assign N3435 = mem[22207:22176] == r_data_i;
  assign N3436 = mem[22175:22144] == r_data_i;
  assign N3437 = mem[22143:22112] == r_data_i;
  assign N3438 = mem[22111:22080] == r_data_i;
  assign N3439 = mem[22079:22048] == r_data_i;
  assign N3440 = mem[22047:22016] == r_data_i;
  assign N3441 = mem[22015:21984] == r_data_i;
  assign N3442 = mem[21983:21952] == r_data_i;
  assign N3443 = mem[21951:21920] == r_data_i;
  assign N3444 = mem[21919:21888] == r_data_i;
  assign N3445 = mem[21887:21856] == r_data_i;
  assign N3446 = mem[21855:21824] == r_data_i;
  assign N3447 = mem[21823:21792] == r_data_i;
  assign N3448 = mem[21791:21760] == r_data_i;
  assign N3449 = mem[21759:21728] == r_data_i;
  assign N3450 = mem[21727:21696] == r_data_i;
  assign N3451 = mem[21695:21664] == r_data_i;
  assign N3452 = mem[21663:21632] == r_data_i;
  assign N3453 = mem[21631:21600] == r_data_i;
  assign N3454 = mem[21599:21568] == r_data_i;
  assign N3455 = mem[21567:21536] == r_data_i;
  assign N3456 = mem[21535:21504] == r_data_i;
  assign N3457 = mem[21503:21472] == r_data_i;
  assign N3458 = mem[21471:21440] == r_data_i;
  assign N3459 = mem[21439:21408] == r_data_i;
  assign N3460 = mem[21407:21376] == r_data_i;
  assign N3461 = mem[21375:21344] == r_data_i;
  assign N3462 = mem[21343:21312] == r_data_i;
  assign N3463 = mem[21311:21280] == r_data_i;
  assign N3464 = mem[21279:21248] == r_data_i;
  assign N3465 = mem[21247:21216] == r_data_i;
  assign N3466 = mem[21215:21184] == r_data_i;
  assign N3467 = mem[21183:21152] == r_data_i;
  assign N3468 = mem[21151:21120] == r_data_i;
  assign N3469 = mem[21119:21088] == r_data_i;
  assign N3470 = mem[21087:21056] == r_data_i;
  assign N3471 = mem[21055:21024] == r_data_i;
  assign N3472 = mem[21023:20992] == r_data_i;
  assign N3473 = mem[20991:20960] == r_data_i;
  assign N3474 = mem[20959:20928] == r_data_i;
  assign N3475 = mem[20927:20896] == r_data_i;
  assign N3476 = mem[20895:20864] == r_data_i;
  assign N3477 = mem[20863:20832] == r_data_i;
  assign N3478 = mem[20831:20800] == r_data_i;
  assign N3479 = mem[20799:20768] == r_data_i;
  assign N3480 = mem[20767:20736] == r_data_i;
  assign N3481 = mem[20735:20704] == r_data_i;
  assign N3482 = mem[20703:20672] == r_data_i;
  assign N3483 = mem[20671:20640] == r_data_i;
  assign N3484 = mem[20639:20608] == r_data_i;
  assign N3485 = mem[20607:20576] == r_data_i;
  assign N3486 = mem[20575:20544] == r_data_i;
  assign N3487 = mem[20543:20512] == r_data_i;
  assign N3488 = mem[20511:20480] == r_data_i;
  assign N3489 = mem[20479:20448] == r_data_i;
  assign N3490 = mem[20447:20416] == r_data_i;
  assign N3491 = mem[20415:20384] == r_data_i;
  assign N3492 = mem[20383:20352] == r_data_i;
  assign N3493 = mem[20351:20320] == r_data_i;
  assign N3494 = mem[20319:20288] == r_data_i;
  assign N3495 = mem[20287:20256] == r_data_i;
  assign N3496 = mem[20255:20224] == r_data_i;
  assign N3497 = mem[20223:20192] == r_data_i;
  assign N3498 = mem[20191:20160] == r_data_i;
  assign N3499 = mem[20159:20128] == r_data_i;
  assign N3500 = mem[20127:20096] == r_data_i;
  assign N3501 = mem[20095:20064] == r_data_i;
  assign N3502 = mem[20063:20032] == r_data_i;
  assign N3503 = mem[20031:20000] == r_data_i;
  assign N3504 = mem[19999:19968] == r_data_i;
  assign N3505 = mem[19967:19936] == r_data_i;
  assign N3506 = mem[19935:19904] == r_data_i;
  assign N3507 = mem[19903:19872] == r_data_i;
  assign N3508 = mem[19871:19840] == r_data_i;
  assign N3509 = mem[19839:19808] == r_data_i;
  assign N3510 = mem[19807:19776] == r_data_i;
  assign N3511 = mem[19775:19744] == r_data_i;
  assign N3512 = mem[19743:19712] == r_data_i;
  assign N3513 = mem[19711:19680] == r_data_i;
  assign N3514 = mem[19679:19648] == r_data_i;
  assign N3515 = mem[19647:19616] == r_data_i;
  assign N3516 = mem[19615:19584] == r_data_i;
  assign N3517 = mem[19583:19552] == r_data_i;
  assign N3518 = mem[19551:19520] == r_data_i;
  assign N3519 = mem[19519:19488] == r_data_i;
  assign N3520 = mem[19487:19456] == r_data_i;
  assign N3521 = mem[19455:19424] == r_data_i;
  assign N3522 = mem[19423:19392] == r_data_i;
  assign N3523 = mem[19391:19360] == r_data_i;
  assign N3524 = mem[19359:19328] == r_data_i;
  assign N3525 = mem[19327:19296] == r_data_i;
  assign N3526 = mem[19295:19264] == r_data_i;
  assign N3527 = mem[19263:19232] == r_data_i;
  assign N3528 = mem[19231:19200] == r_data_i;
  assign N3529 = mem[19199:19168] == r_data_i;
  assign N3530 = mem[19167:19136] == r_data_i;
  assign N3531 = mem[19135:19104] == r_data_i;
  assign N3532 = mem[19103:19072] == r_data_i;
  assign N3533 = mem[19071:19040] == r_data_i;
  assign N3534 = mem[19039:19008] == r_data_i;
  assign N3535 = mem[19007:18976] == r_data_i;
  assign N3536 = mem[18975:18944] == r_data_i;
  assign N3537 = mem[18943:18912] == r_data_i;
  assign N3538 = mem[18911:18880] == r_data_i;
  assign N3539 = mem[18879:18848] == r_data_i;
  assign N3540 = mem[18847:18816] == r_data_i;
  assign N3541 = mem[18815:18784] == r_data_i;
  assign N3542 = mem[18783:18752] == r_data_i;
  assign N3543 = mem[18751:18720] == r_data_i;
  assign N3544 = mem[18719:18688] == r_data_i;
  assign N3545 = mem[18687:18656] == r_data_i;
  assign N3546 = mem[18655:18624] == r_data_i;
  assign N3547 = mem[18623:18592] == r_data_i;
  assign N3548 = mem[18591:18560] == r_data_i;
  assign N3549 = mem[18559:18528] == r_data_i;
  assign N3550 = mem[18527:18496] == r_data_i;
  assign N3551 = mem[18495:18464] == r_data_i;
  assign N3552 = mem[18463:18432] == r_data_i;
  assign N3553 = mem[18431:18400] == r_data_i;
  assign N3554 = mem[18399:18368] == r_data_i;
  assign N3555 = mem[18367:18336] == r_data_i;
  assign N3556 = mem[18335:18304] == r_data_i;
  assign N3557 = mem[18303:18272] == r_data_i;
  assign N3558 = mem[18271:18240] == r_data_i;
  assign N3559 = mem[18239:18208] == r_data_i;
  assign N3560 = mem[18207:18176] == r_data_i;
  assign N3561 = mem[18175:18144] == r_data_i;
  assign N3562 = mem[18143:18112] == r_data_i;
  assign N3563 = mem[18111:18080] == r_data_i;
  assign N3564 = mem[18079:18048] == r_data_i;
  assign N3565 = mem[18047:18016] == r_data_i;
  assign N3566 = mem[18015:17984] == r_data_i;
  assign N3567 = mem[17983:17952] == r_data_i;
  assign N3568 = mem[17951:17920] == r_data_i;
  assign N3569 = mem[17919:17888] == r_data_i;
  assign N3570 = mem[17887:17856] == r_data_i;
  assign N3571 = mem[17855:17824] == r_data_i;
  assign N3572 = mem[17823:17792] == r_data_i;
  assign N3573 = mem[17791:17760] == r_data_i;
  assign N3574 = mem[17759:17728] == r_data_i;
  assign N3575 = mem[17727:17696] == r_data_i;
  assign N3576 = mem[17695:17664] == r_data_i;
  assign N3577 = mem[17663:17632] == r_data_i;
  assign N3578 = mem[17631:17600] == r_data_i;
  assign N3579 = mem[17599:17568] == r_data_i;
  assign N3580 = mem[17567:17536] == r_data_i;
  assign N3581 = mem[17535:17504] == r_data_i;
  assign N3582 = mem[17503:17472] == r_data_i;
  assign N3583 = mem[17471:17440] == r_data_i;
  assign N3584 = mem[17439:17408] == r_data_i;
  assign N3585 = mem[17407:17376] == r_data_i;
  assign N3586 = mem[17375:17344] == r_data_i;
  assign N3587 = mem[17343:17312] == r_data_i;
  assign N3588 = mem[17311:17280] == r_data_i;
  assign N3589 = mem[17279:17248] == r_data_i;
  assign N3590 = mem[17247:17216] == r_data_i;
  assign N3591 = mem[17215:17184] == r_data_i;
  assign N3592 = mem[17183:17152] == r_data_i;
  assign N3593 = mem[17151:17120] == r_data_i;
  assign N3594 = mem[17119:17088] == r_data_i;
  assign N3595 = mem[17087:17056] == r_data_i;
  assign N3596 = mem[17055:17024] == r_data_i;
  assign N3597 = mem[17023:16992] == r_data_i;
  assign N3598 = mem[16991:16960] == r_data_i;
  assign N3599 = mem[16959:16928] == r_data_i;
  assign N3600 = mem[16927:16896] == r_data_i;
  assign N3601 = mem[16895:16864] == r_data_i;
  assign N3602 = mem[16863:16832] == r_data_i;
  assign N3603 = mem[16831:16800] == r_data_i;
  assign N3604 = mem[16799:16768] == r_data_i;
  assign N3605 = mem[16767:16736] == r_data_i;
  assign N3606 = mem[16735:16704] == r_data_i;
  assign N3607 = mem[16703:16672] == r_data_i;
  assign N3608 = mem[16671:16640] == r_data_i;
  assign N3609 = mem[16639:16608] == r_data_i;
  assign N3610 = mem[16607:16576] == r_data_i;
  assign N3611 = mem[16575:16544] == r_data_i;
  assign N3612 = mem[16543:16512] == r_data_i;
  assign N3613 = mem[16511:16480] == r_data_i;
  assign N3614 = mem[16479:16448] == r_data_i;
  assign N3615 = mem[16447:16416] == r_data_i;
  assign N3616 = mem[16415:16384] == r_data_i;
  assign N3617 = mem[16383:16352] == r_data_i;
  assign N3618 = mem[16351:16320] == r_data_i;
  assign N3619 = mem[16319:16288] == r_data_i;
  assign N3620 = mem[16287:16256] == r_data_i;
  assign N3621 = mem[16255:16224] == r_data_i;
  assign N3622 = mem[16223:16192] == r_data_i;
  assign N3623 = mem[16191:16160] == r_data_i;
  assign N3624 = mem[16159:16128] == r_data_i;
  assign N3625 = mem[16127:16096] == r_data_i;
  assign N3626 = mem[16095:16064] == r_data_i;
  assign N3627 = mem[16063:16032] == r_data_i;
  assign N3628 = mem[16031:16000] == r_data_i;
  assign N3629 = mem[15999:15968] == r_data_i;
  assign N3630 = mem[15967:15936] == r_data_i;
  assign N3631 = mem[15935:15904] == r_data_i;
  assign N3632 = mem[15903:15872] == r_data_i;
  assign N3633 = mem[15871:15840] == r_data_i;
  assign N3634 = mem[15839:15808] == r_data_i;
  assign N3635 = mem[15807:15776] == r_data_i;
  assign N3636 = mem[15775:15744] == r_data_i;
  assign N3637 = mem[15743:15712] == r_data_i;
  assign N3638 = mem[15711:15680] == r_data_i;
  assign N3639 = mem[15679:15648] == r_data_i;
  assign N3640 = mem[15647:15616] == r_data_i;
  assign N3641 = mem[15615:15584] == r_data_i;
  assign N3642 = mem[15583:15552] == r_data_i;
  assign N3643 = mem[15551:15520] == r_data_i;
  assign N3644 = mem[15519:15488] == r_data_i;
  assign N3645 = mem[15487:15456] == r_data_i;
  assign N3646 = mem[15455:15424] == r_data_i;
  assign N3647 = mem[15423:15392] == r_data_i;
  assign N3648 = mem[15391:15360] == r_data_i;
  assign N3649 = mem[15359:15328] == r_data_i;
  assign N3650 = mem[15327:15296] == r_data_i;
  assign N3651 = mem[15295:15264] == r_data_i;
  assign N3652 = mem[15263:15232] == r_data_i;
  assign N3653 = mem[15231:15200] == r_data_i;
  assign N3654 = mem[15199:15168] == r_data_i;
  assign N3655 = mem[15167:15136] == r_data_i;
  assign N3656 = mem[15135:15104] == r_data_i;
  assign N3657 = mem[15103:15072] == r_data_i;
  assign N3658 = mem[15071:15040] == r_data_i;
  assign N3659 = mem[15039:15008] == r_data_i;
  assign N3660 = mem[15007:14976] == r_data_i;
  assign N3661 = mem[14975:14944] == r_data_i;
  assign N3662 = mem[14943:14912] == r_data_i;
  assign N3663 = mem[14911:14880] == r_data_i;
  assign N3664 = mem[14879:14848] == r_data_i;
  assign N3665 = mem[14847:14816] == r_data_i;
  assign N3666 = mem[14815:14784] == r_data_i;
  assign N3667 = mem[14783:14752] == r_data_i;
  assign N3668 = mem[14751:14720] == r_data_i;
  assign N3669 = mem[14719:14688] == r_data_i;
  assign N3670 = mem[14687:14656] == r_data_i;
  assign N3671 = mem[14655:14624] == r_data_i;
  assign N3672 = mem[14623:14592] == r_data_i;
  assign N3673 = mem[14591:14560] == r_data_i;
  assign N3674 = mem[14559:14528] == r_data_i;
  assign N3675 = mem[14527:14496] == r_data_i;
  assign N3676 = mem[14495:14464] == r_data_i;
  assign N3677 = mem[14463:14432] == r_data_i;
  assign N3678 = mem[14431:14400] == r_data_i;
  assign N3679 = mem[14399:14368] == r_data_i;
  assign N3680 = mem[14367:14336] == r_data_i;
  assign N3681 = mem[14335:14304] == r_data_i;
  assign N3682 = mem[14303:14272] == r_data_i;
  assign N3683 = mem[14271:14240] == r_data_i;
  assign N3684 = mem[14239:14208] == r_data_i;
  assign N3685 = mem[14207:14176] == r_data_i;
  assign N3686 = mem[14175:14144] == r_data_i;
  assign N3687 = mem[14143:14112] == r_data_i;
  assign N3688 = mem[14111:14080] == r_data_i;
  assign N3689 = mem[14079:14048] == r_data_i;
  assign N3690 = mem[14047:14016] == r_data_i;
  assign N3691 = mem[14015:13984] == r_data_i;
  assign N3692 = mem[13983:13952] == r_data_i;
  assign N3693 = mem[13951:13920] == r_data_i;
  assign N3694 = mem[13919:13888] == r_data_i;
  assign N3695 = mem[13887:13856] == r_data_i;
  assign N3696 = mem[13855:13824] == r_data_i;
  assign N3697 = mem[13823:13792] == r_data_i;
  assign N3698 = mem[13791:13760] == r_data_i;
  assign N3699 = mem[13759:13728] == r_data_i;
  assign N3700 = mem[13727:13696] == r_data_i;
  assign N3701 = mem[13695:13664] == r_data_i;
  assign N3702 = mem[13663:13632] == r_data_i;
  assign N3703 = mem[13631:13600] == r_data_i;
  assign N3704 = mem[13599:13568] == r_data_i;
  assign N3705 = mem[13567:13536] == r_data_i;
  assign N3706 = mem[13535:13504] == r_data_i;
  assign N3707 = mem[13503:13472] == r_data_i;
  assign N3708 = mem[13471:13440] == r_data_i;
  assign N3709 = mem[13439:13408] == r_data_i;
  assign N3710 = mem[13407:13376] == r_data_i;
  assign N3711 = mem[13375:13344] == r_data_i;
  assign N3712 = mem[13343:13312] == r_data_i;
  assign N3713 = mem[13311:13280] == r_data_i;
  assign N3714 = mem[13279:13248] == r_data_i;
  assign N3715 = mem[13247:13216] == r_data_i;
  assign N3716 = mem[13215:13184] == r_data_i;
  assign N3717 = mem[13183:13152] == r_data_i;
  assign N3718 = mem[13151:13120] == r_data_i;
  assign N3719 = mem[13119:13088] == r_data_i;
  assign N3720 = mem[13087:13056] == r_data_i;
  assign N3721 = mem[13055:13024] == r_data_i;
  assign N3722 = mem[13023:12992] == r_data_i;
  assign N3723 = mem[12991:12960] == r_data_i;
  assign N3724 = mem[12959:12928] == r_data_i;
  assign N3725 = mem[12927:12896] == r_data_i;
  assign N3726 = mem[12895:12864] == r_data_i;
  assign N3727 = mem[12863:12832] == r_data_i;
  assign N3728 = mem[12831:12800] == r_data_i;
  assign N3729 = mem[12799:12768] == r_data_i;
  assign N3730 = mem[12767:12736] == r_data_i;
  assign N3731 = mem[12735:12704] == r_data_i;
  assign N3732 = mem[12703:12672] == r_data_i;
  assign N3733 = mem[12671:12640] == r_data_i;
  assign N3734 = mem[12639:12608] == r_data_i;
  assign N3735 = mem[12607:12576] == r_data_i;
  assign N3736 = mem[12575:12544] == r_data_i;
  assign N3737 = mem[12543:12512] == r_data_i;
  assign N3738 = mem[12511:12480] == r_data_i;
  assign N3739 = mem[12479:12448] == r_data_i;
  assign N3740 = mem[12447:12416] == r_data_i;
  assign N3741 = mem[12415:12384] == r_data_i;
  assign N3742 = mem[12383:12352] == r_data_i;
  assign N3743 = mem[12351:12320] == r_data_i;
  assign N3744 = mem[12319:12288] == r_data_i;
  assign N3745 = mem[12287:12256] == r_data_i;
  assign N3746 = mem[12255:12224] == r_data_i;
  assign N3747 = mem[12223:12192] == r_data_i;
  assign N3748 = mem[12191:12160] == r_data_i;
  assign N3749 = mem[12159:12128] == r_data_i;
  assign N3750 = mem[12127:12096] == r_data_i;
  assign N3751 = mem[12095:12064] == r_data_i;
  assign N3752 = mem[12063:12032] == r_data_i;
  assign N3753 = mem[12031:12000] == r_data_i;
  assign N3754 = mem[11999:11968] == r_data_i;
  assign N3755 = mem[11967:11936] == r_data_i;
  assign N3756 = mem[11935:11904] == r_data_i;
  assign N3757 = mem[11903:11872] == r_data_i;
  assign N3758 = mem[11871:11840] == r_data_i;
  assign N3759 = mem[11839:11808] == r_data_i;
  assign N3760 = mem[11807:11776] == r_data_i;
  assign N3761 = mem[11775:11744] == r_data_i;
  assign N3762 = mem[11743:11712] == r_data_i;
  assign N3763 = mem[11711:11680] == r_data_i;
  assign N3764 = mem[11679:11648] == r_data_i;
  assign N3765 = mem[11647:11616] == r_data_i;
  assign N3766 = mem[11615:11584] == r_data_i;
  assign N3767 = mem[11583:11552] == r_data_i;
  assign N3768 = mem[11551:11520] == r_data_i;
  assign N3769 = mem[11519:11488] == r_data_i;
  assign N3770 = mem[11487:11456] == r_data_i;
  assign N3771 = mem[11455:11424] == r_data_i;
  assign N3772 = mem[11423:11392] == r_data_i;
  assign N3773 = mem[11391:11360] == r_data_i;
  assign N3774 = mem[11359:11328] == r_data_i;
  assign N3775 = mem[11327:11296] == r_data_i;
  assign N3776 = mem[11295:11264] == r_data_i;
  assign N3777 = mem[11263:11232] == r_data_i;
  assign N3778 = mem[11231:11200] == r_data_i;
  assign N3779 = mem[11199:11168] == r_data_i;
  assign N3780 = mem[11167:11136] == r_data_i;
  assign N3781 = mem[11135:11104] == r_data_i;
  assign N3782 = mem[11103:11072] == r_data_i;
  assign N3783 = mem[11071:11040] == r_data_i;
  assign N3784 = mem[11039:11008] == r_data_i;
  assign N3785 = mem[11007:10976] == r_data_i;
  assign N3786 = mem[10975:10944] == r_data_i;
  assign N3787 = mem[10943:10912] == r_data_i;
  assign N3788 = mem[10911:10880] == r_data_i;
  assign N3789 = mem[10879:10848] == r_data_i;
  assign N3790 = mem[10847:10816] == r_data_i;
  assign N3791 = mem[10815:10784] == r_data_i;
  assign N3792 = mem[10783:10752] == r_data_i;
  assign N3793 = mem[10751:10720] == r_data_i;
  assign N3794 = mem[10719:10688] == r_data_i;
  assign N3795 = mem[10687:10656] == r_data_i;
  assign N3796 = mem[10655:10624] == r_data_i;
  assign N3797 = mem[10623:10592] == r_data_i;
  assign N3798 = mem[10591:10560] == r_data_i;
  assign N3799 = mem[10559:10528] == r_data_i;
  assign N3800 = mem[10527:10496] == r_data_i;
  assign N3801 = mem[10495:10464] == r_data_i;
  assign N3802 = mem[10463:10432] == r_data_i;
  assign N3803 = mem[10431:10400] == r_data_i;
  assign N3804 = mem[10399:10368] == r_data_i;
  assign N3805 = mem[10367:10336] == r_data_i;
  assign N3806 = mem[10335:10304] == r_data_i;
  assign N3807 = mem[10303:10272] == r_data_i;
  assign N3808 = mem[10271:10240] == r_data_i;
  assign N3809 = mem[10239:10208] == r_data_i;
  assign N3810 = mem[10207:10176] == r_data_i;
  assign N3811 = mem[10175:10144] == r_data_i;
  assign N3812 = mem[10143:10112] == r_data_i;
  assign N3813 = mem[10111:10080] == r_data_i;
  assign N3814 = mem[10079:10048] == r_data_i;
  assign N3815 = mem[10047:10016] == r_data_i;
  assign N3816 = mem[10015:9984] == r_data_i;
  assign N3817 = mem[9983:9952] == r_data_i;
  assign N3818 = mem[9951:9920] == r_data_i;
  assign N3819 = mem[9919:9888] == r_data_i;
  assign N3820 = mem[9887:9856] == r_data_i;
  assign N3821 = mem[9855:9824] == r_data_i;
  assign N3822 = mem[9823:9792] == r_data_i;
  assign N3823 = mem[9791:9760] == r_data_i;
  assign N3824 = mem[9759:9728] == r_data_i;
  assign N3825 = mem[9727:9696] == r_data_i;
  assign N3826 = mem[9695:9664] == r_data_i;
  assign N3827 = mem[9663:9632] == r_data_i;
  assign N3828 = mem[9631:9600] == r_data_i;
  assign N3829 = mem[9599:9568] == r_data_i;
  assign N3830 = mem[9567:9536] == r_data_i;
  assign N3831 = mem[9535:9504] == r_data_i;
  assign N3832 = mem[9503:9472] == r_data_i;
  assign N3833 = mem[9471:9440] == r_data_i;
  assign N3834 = mem[9439:9408] == r_data_i;
  assign N3835 = mem[9407:9376] == r_data_i;
  assign N3836 = mem[9375:9344] == r_data_i;
  assign N3837 = mem[9343:9312] == r_data_i;
  assign N3838 = mem[9311:9280] == r_data_i;
  assign N3839 = mem[9279:9248] == r_data_i;
  assign N3840 = mem[9247:9216] == r_data_i;
  assign N3841 = mem[9215:9184] == r_data_i;
  assign N3842 = mem[9183:9152] == r_data_i;
  assign N3843 = mem[9151:9120] == r_data_i;
  assign N3844 = mem[9119:9088] == r_data_i;
  assign N3845 = mem[9087:9056] == r_data_i;
  assign N3846 = mem[9055:9024] == r_data_i;
  assign N3847 = mem[9023:8992] == r_data_i;
  assign N3848 = mem[8991:8960] == r_data_i;
  assign N3849 = mem[8959:8928] == r_data_i;
  assign N3850 = mem[8927:8896] == r_data_i;
  assign N3851 = mem[8895:8864] == r_data_i;
  assign N3852 = mem[8863:8832] == r_data_i;
  assign N3853 = mem[8831:8800] == r_data_i;
  assign N3854 = mem[8799:8768] == r_data_i;
  assign N3855 = mem[8767:8736] == r_data_i;
  assign N3856 = mem[8735:8704] == r_data_i;
  assign N3857 = mem[8703:8672] == r_data_i;
  assign N3858 = mem[8671:8640] == r_data_i;
  assign N3859 = mem[8639:8608] == r_data_i;
  assign N3860 = mem[8607:8576] == r_data_i;
  assign N3861 = mem[8575:8544] == r_data_i;
  assign N3862 = mem[8543:8512] == r_data_i;
  assign N3863 = mem[8511:8480] == r_data_i;
  assign N3864 = mem[8479:8448] == r_data_i;
  assign N3865 = mem[8447:8416] == r_data_i;
  assign N3866 = mem[8415:8384] == r_data_i;
  assign N3867 = mem[8383:8352] == r_data_i;
  assign N3868 = mem[8351:8320] == r_data_i;
  assign N3869 = mem[8319:8288] == r_data_i;
  assign N3870 = mem[8287:8256] == r_data_i;
  assign N3871 = mem[8255:8224] == r_data_i;
  assign N3872 = mem[8223:8192] == r_data_i;
  assign N3873 = mem[8191:8160] == r_data_i;
  assign N3874 = mem[8159:8128] == r_data_i;
  assign N3875 = mem[8127:8096] == r_data_i;
  assign N3876 = mem[8095:8064] == r_data_i;
  assign N3877 = mem[8063:8032] == r_data_i;
  assign N3878 = mem[8031:8000] == r_data_i;
  assign N3879 = mem[7999:7968] == r_data_i;
  assign N3880 = mem[7967:7936] == r_data_i;
  assign N3881 = mem[7935:7904] == r_data_i;
  assign N3882 = mem[7903:7872] == r_data_i;
  assign N3883 = mem[7871:7840] == r_data_i;
  assign N3884 = mem[7839:7808] == r_data_i;
  assign N3885 = mem[7807:7776] == r_data_i;
  assign N3886 = mem[7775:7744] == r_data_i;
  assign N3887 = mem[7743:7712] == r_data_i;
  assign N3888 = mem[7711:7680] == r_data_i;
  assign N3889 = mem[7679:7648] == r_data_i;
  assign N3890 = mem[7647:7616] == r_data_i;
  assign N3891 = mem[7615:7584] == r_data_i;
  assign N3892 = mem[7583:7552] == r_data_i;
  assign N3893 = mem[7551:7520] == r_data_i;
  assign N3894 = mem[7519:7488] == r_data_i;
  assign N3895 = mem[7487:7456] == r_data_i;
  assign N3896 = mem[7455:7424] == r_data_i;
  assign N3897 = mem[7423:7392] == r_data_i;
  assign N3898 = mem[7391:7360] == r_data_i;
  assign N3899 = mem[7359:7328] == r_data_i;
  assign N3900 = mem[7327:7296] == r_data_i;
  assign N3901 = mem[7295:7264] == r_data_i;
  assign N3902 = mem[7263:7232] == r_data_i;
  assign N3903 = mem[7231:7200] == r_data_i;
  assign N3904 = mem[7199:7168] == r_data_i;
  assign N3905 = mem[7167:7136] == r_data_i;
  assign N3906 = mem[7135:7104] == r_data_i;
  assign N3907 = mem[7103:7072] == r_data_i;
  assign N3908 = mem[7071:7040] == r_data_i;
  assign N3909 = mem[7039:7008] == r_data_i;
  assign N3910 = mem[7007:6976] == r_data_i;
  assign N3911 = mem[6975:6944] == r_data_i;
  assign N3912 = mem[6943:6912] == r_data_i;
  assign N3913 = mem[6911:6880] == r_data_i;
  assign N3914 = mem[6879:6848] == r_data_i;
  assign N3915 = mem[6847:6816] == r_data_i;
  assign N3916 = mem[6815:6784] == r_data_i;
  assign N3917 = mem[6783:6752] == r_data_i;
  assign N3918 = mem[6751:6720] == r_data_i;
  assign N3919 = mem[6719:6688] == r_data_i;
  assign N3920 = mem[6687:6656] == r_data_i;
  assign N3921 = mem[6655:6624] == r_data_i;
  assign N3922 = mem[6623:6592] == r_data_i;
  assign N3923 = mem[6591:6560] == r_data_i;
  assign N3924 = mem[6559:6528] == r_data_i;
  assign N3925 = mem[6527:6496] == r_data_i;
  assign N3926 = mem[6495:6464] == r_data_i;
  assign N3927 = mem[6463:6432] == r_data_i;
  assign N3928 = mem[6431:6400] == r_data_i;
  assign N3929 = mem[6399:6368] == r_data_i;
  assign N3930 = mem[6367:6336] == r_data_i;
  assign N3931 = mem[6335:6304] == r_data_i;
  assign N3932 = mem[6303:6272] == r_data_i;
  assign N3933 = mem[6271:6240] == r_data_i;
  assign N3934 = mem[6239:6208] == r_data_i;
  assign N3935 = mem[6207:6176] == r_data_i;
  assign N3936 = mem[6175:6144] == r_data_i;
  assign N3937 = mem[6143:6112] == r_data_i;
  assign N3938 = mem[6111:6080] == r_data_i;
  assign N3939 = mem[6079:6048] == r_data_i;
  assign N3940 = mem[6047:6016] == r_data_i;
  assign N3941 = mem[6015:5984] == r_data_i;
  assign N3942 = mem[5983:5952] == r_data_i;
  assign N3943 = mem[5951:5920] == r_data_i;
  assign N3944 = mem[5919:5888] == r_data_i;
  assign N3945 = mem[5887:5856] == r_data_i;
  assign N3946 = mem[5855:5824] == r_data_i;
  assign N3947 = mem[5823:5792] == r_data_i;
  assign N3948 = mem[5791:5760] == r_data_i;
  assign N3949 = mem[5759:5728] == r_data_i;
  assign N3950 = mem[5727:5696] == r_data_i;
  assign N3951 = mem[5695:5664] == r_data_i;
  assign N3952 = mem[5663:5632] == r_data_i;
  assign N3953 = mem[5631:5600] == r_data_i;
  assign N3954 = mem[5599:5568] == r_data_i;
  assign N3955 = mem[5567:5536] == r_data_i;
  assign N3956 = mem[5535:5504] == r_data_i;
  assign N3957 = mem[5503:5472] == r_data_i;
  assign N3958 = mem[5471:5440] == r_data_i;
  assign N3959 = mem[5439:5408] == r_data_i;
  assign N3960 = mem[5407:5376] == r_data_i;
  assign N3961 = mem[5375:5344] == r_data_i;
  assign N3962 = mem[5343:5312] == r_data_i;
  assign N3963 = mem[5311:5280] == r_data_i;
  assign N3964 = mem[5279:5248] == r_data_i;
  assign N3965 = mem[5247:5216] == r_data_i;
  assign N3966 = mem[5215:5184] == r_data_i;
  assign N3967 = mem[5183:5152] == r_data_i;
  assign N3968 = mem[5151:5120] == r_data_i;
  assign N3969 = mem[5119:5088] == r_data_i;
  assign N3970 = mem[5087:5056] == r_data_i;
  assign N3971 = mem[5055:5024] == r_data_i;
  assign N3972 = mem[5023:4992] == r_data_i;
  assign N3973 = mem[4991:4960] == r_data_i;
  assign N3974 = mem[4959:4928] == r_data_i;
  assign N3975 = mem[4927:4896] == r_data_i;
  assign N3976 = mem[4895:4864] == r_data_i;
  assign N3977 = mem[4863:4832] == r_data_i;
  assign N3978 = mem[4831:4800] == r_data_i;
  assign N3979 = mem[4799:4768] == r_data_i;
  assign N3980 = mem[4767:4736] == r_data_i;
  assign N3981 = mem[4735:4704] == r_data_i;
  assign N3982 = mem[4703:4672] == r_data_i;
  assign N3983 = mem[4671:4640] == r_data_i;
  assign N3984 = mem[4639:4608] == r_data_i;
  assign N3985 = mem[4607:4576] == r_data_i;
  assign N3986 = mem[4575:4544] == r_data_i;
  assign N3987 = mem[4543:4512] == r_data_i;
  assign N3988 = mem[4511:4480] == r_data_i;
  assign N3989 = mem[4479:4448] == r_data_i;
  assign N3990 = mem[4447:4416] == r_data_i;
  assign N3991 = mem[4415:4384] == r_data_i;
  assign N3992 = mem[4383:4352] == r_data_i;
  assign N3993 = mem[4351:4320] == r_data_i;
  assign N3994 = mem[4319:4288] == r_data_i;
  assign N3995 = mem[4287:4256] == r_data_i;
  assign N3996 = mem[4255:4224] == r_data_i;
  assign N3997 = mem[4223:4192] == r_data_i;
  assign N3998 = mem[4191:4160] == r_data_i;
  assign N3999 = mem[4159:4128] == r_data_i;
  assign N4000 = mem[4127:4096] == r_data_i;
  assign N4001 = mem[4095:4064] == r_data_i;
  assign N4002 = mem[4063:4032] == r_data_i;
  assign N4003 = mem[4031:4000] == r_data_i;
  assign N4004 = mem[3999:3968] == r_data_i;
  assign N4005 = mem[3967:3936] == r_data_i;
  assign N4006 = mem[3935:3904] == r_data_i;
  assign N4007 = mem[3903:3872] == r_data_i;
  assign N4008 = mem[3871:3840] == r_data_i;
  assign N4009 = mem[3839:3808] == r_data_i;
  assign N4010 = mem[3807:3776] == r_data_i;
  assign N4011 = mem[3775:3744] == r_data_i;
  assign N4012 = mem[3743:3712] == r_data_i;
  assign N4013 = mem[3711:3680] == r_data_i;
  assign N4014 = mem[3679:3648] == r_data_i;
  assign N4015 = mem[3647:3616] == r_data_i;
  assign N4016 = mem[3615:3584] == r_data_i;
  assign N4017 = mem[3583:3552] == r_data_i;
  assign N4018 = mem[3551:3520] == r_data_i;
  assign N4019 = mem[3519:3488] == r_data_i;
  assign N4020 = mem[3487:3456] == r_data_i;
  assign N4021 = mem[3455:3424] == r_data_i;
  assign N4022 = mem[3423:3392] == r_data_i;
  assign N4023 = mem[3391:3360] == r_data_i;
  assign N4024 = mem[3359:3328] == r_data_i;
  assign N4025 = mem[3327:3296] == r_data_i;
  assign N4026 = mem[3295:3264] == r_data_i;
  assign N4027 = mem[3263:3232] == r_data_i;
  assign N4028 = mem[3231:3200] == r_data_i;
  assign N4029 = mem[3199:3168] == r_data_i;
  assign N4030 = mem[3167:3136] == r_data_i;
  assign N4031 = mem[3135:3104] == r_data_i;
  assign N4032 = mem[3103:3072] == r_data_i;
  assign N4033 = mem[3071:3040] == r_data_i;
  assign N4034 = mem[3039:3008] == r_data_i;
  assign N4035 = mem[3007:2976] == r_data_i;
  assign N4036 = mem[2975:2944] == r_data_i;
  assign N4037 = mem[2943:2912] == r_data_i;
  assign N4038 = mem[2911:2880] == r_data_i;
  assign N4039 = mem[2879:2848] == r_data_i;
  assign N4040 = mem[2847:2816] == r_data_i;
  assign N4041 = mem[2815:2784] == r_data_i;
  assign N4042 = mem[2783:2752] == r_data_i;
  assign N4043 = mem[2751:2720] == r_data_i;
  assign N4044 = mem[2719:2688] == r_data_i;
  assign N4045 = mem[2687:2656] == r_data_i;
  assign N4046 = mem[2655:2624] == r_data_i;
  assign N4047 = mem[2623:2592] == r_data_i;
  assign N4048 = mem[2591:2560] == r_data_i;
  assign N4049 = mem[2559:2528] == r_data_i;
  assign N4050 = mem[2527:2496] == r_data_i;
  assign N4051 = mem[2495:2464] == r_data_i;
  assign N4052 = mem[2463:2432] == r_data_i;
  assign N4053 = mem[2431:2400] == r_data_i;
  assign N4054 = mem[2399:2368] == r_data_i;
  assign N4055 = mem[2367:2336] == r_data_i;
  assign N4056 = mem[2335:2304] == r_data_i;
  assign N4057 = mem[2303:2272] == r_data_i;
  assign N4058 = mem[2271:2240] == r_data_i;
  assign N4059 = mem[2239:2208] == r_data_i;
  assign N4060 = mem[2207:2176] == r_data_i;
  assign N4061 = mem[2175:2144] == r_data_i;
  assign N4062 = mem[2143:2112] == r_data_i;
  assign N4063 = mem[2111:2080] == r_data_i;
  assign N4064 = mem[2079:2048] == r_data_i;
  assign N4065 = mem[2047:2016] == r_data_i;
  assign N4066 = mem[2015:1984] == r_data_i;
  assign N4067 = mem[1983:1952] == r_data_i;
  assign N4068 = mem[1951:1920] == r_data_i;
  assign N4069 = mem[1919:1888] == r_data_i;
  assign N4070 = mem[1887:1856] == r_data_i;
  assign N4071 = mem[1855:1824] == r_data_i;
  assign N4072 = mem[1823:1792] == r_data_i;
  assign N4073 = mem[1791:1760] == r_data_i;
  assign N4074 = mem[1759:1728] == r_data_i;
  assign N4075 = mem[1727:1696] == r_data_i;
  assign N4076 = mem[1695:1664] == r_data_i;
  assign N4077 = mem[1663:1632] == r_data_i;
  assign N4078 = mem[1631:1600] == r_data_i;
  assign N4079 = mem[1599:1568] == r_data_i;
  assign N4080 = mem[1567:1536] == r_data_i;
  assign N4081 = mem[1535:1504] == r_data_i;
  assign N4082 = mem[1503:1472] == r_data_i;
  assign N4083 = mem[1471:1440] == r_data_i;
  assign N4084 = mem[1439:1408] == r_data_i;
  assign N4085 = mem[1407:1376] == r_data_i;
  assign N4086 = mem[1375:1344] == r_data_i;
  assign N4087 = mem[1343:1312] == r_data_i;
  assign N4088 = mem[1311:1280] == r_data_i;
  assign N4089 = mem[1279:1248] == r_data_i;
  assign N4090 = mem[1247:1216] == r_data_i;
  assign N4091 = mem[1215:1184] == r_data_i;
  assign N4092 = mem[1183:1152] == r_data_i;
  assign N4093 = mem[1151:1120] == r_data_i;
  assign N4094 = mem[1119:1088] == r_data_i;
  assign N4095 = mem[1087:1056] == r_data_i;
  assign N4096 = mem[1055:1024] == r_data_i;
  assign N4097 = mem[1023:992] == r_data_i;
  assign N4098 = mem[991:960] == r_data_i;
  assign N4099 = mem[959:928] == r_data_i;
  assign N4100 = mem[927:896] == r_data_i;
  assign N4101 = mem[895:864] == r_data_i;
  assign N4102 = mem[863:832] == r_data_i;
  assign N4103 = mem[831:800] == r_data_i;
  assign N4104 = mem[799:768] == r_data_i;
  assign N4105 = mem[767:736] == r_data_i;
  assign N4106 = mem[735:704] == r_data_i;
  assign N4107 = mem[703:672] == r_data_i;
  assign N4108 = mem[671:640] == r_data_i;
  assign N4109 = mem[639:608] == r_data_i;
  assign N4110 = mem[607:576] == r_data_i;
  assign N4111 = mem[575:544] == r_data_i;
  assign N4112 = mem[543:512] == r_data_i;
  assign N4113 = mem[511:480] == r_data_i;
  assign N4114 = mem[479:448] == r_data_i;
  assign N4115 = mem[447:416] == r_data_i;
  assign N4116 = mem[415:384] == r_data_i;
  assign N4117 = mem[383:352] == r_data_i;
  assign N4118 = mem[351:320] == r_data_i;
  assign N4119 = mem[319:288] == r_data_i;
  assign N4120 = mem[287:256] == r_data_i;
  assign N4121 = mem[255:224] == r_data_i;
  assign N4122 = mem[223:192] == r_data_i;
  assign N4123 = mem[191:160] == r_data_i;
  assign N4124 = mem[159:128] == r_data_i;
  assign N4125 = mem[127:96] == r_data_i;
  assign N4126 = mem[95:64] == r_data_i;
  assign N4127 = mem[63:32] == r_data_i;
  assign N4128 = mem[31:0] == r_data_i;

  bsg_priority_encode_width_p1024_lo_to_hi_p1
  fi3_pe
  (
    .i(match_array),
    .addr_o(r_addr_o),
    .v_o(matched)
  );


  bsg_priority_encode_width_p1024_lo_to_hi_p1
  fi5_epe
  (
    .i(empty_array),
    .addr_o(empty_addr_o),
    .v_o(empty_found)
  );

  assign N4129 = w_addr_i[8] & w_addr_i[9];
  assign N4130 = N0 & w_addr_i[9];
  assign N0 = ~w_addr_i[8];
  assign N4131 = w_addr_i[8] & N1;
  assign N1 = ~w_addr_i[9];
  assign N4132 = N2 & N3;
  assign N2 = ~w_addr_i[8];
  assign N3 = ~w_addr_i[9];
  assign N4133 = ~w_addr_i[7];
  assign N4134 = w_addr_i[5] & w_addr_i[6];
  assign N4135 = N4 & w_addr_i[6];
  assign N4 = ~w_addr_i[5];
  assign N4136 = w_addr_i[5] & N5;
  assign N5 = ~w_addr_i[6];
  assign N4137 = N6 & N7;
  assign N6 = ~w_addr_i[5];
  assign N7 = ~w_addr_i[6];
  assign N4138 = w_addr_i[7] & N4134;
  assign N4139 = w_addr_i[7] & N4135;
  assign N4140 = w_addr_i[7] & N4136;
  assign N4141 = w_addr_i[7] & N4137;
  assign N4142 = N4133 & N4134;
  assign N4143 = N4133 & N4135;
  assign N4144 = N4133 & N4136;
  assign N4145 = N4133 & N4137;
  assign N4146 = N4129 & N4138;
  assign N4147 = N4129 & N4139;
  assign N4148 = N4129 & N4140;
  assign N4149 = N4129 & N4141;
  assign N4150 = N4129 & N4142;
  assign N4151 = N4129 & N4143;
  assign N4152 = N4129 & N4144;
  assign N4153 = N4129 & N4145;
  assign N4154 = N4130 & N4138;
  assign N4155 = N4130 & N4139;
  assign N4156 = N4130 & N4140;
  assign N4157 = N4130 & N4141;
  assign N4158 = N4130 & N4142;
  assign N4159 = N4130 & N4143;
  assign N4160 = N4130 & N4144;
  assign N4161 = N4130 & N4145;
  assign N4162 = N4131 & N4138;
  assign N4163 = N4131 & N4139;
  assign N4164 = N4131 & N4140;
  assign N4165 = N4131 & N4141;
  assign N4166 = N4131 & N4142;
  assign N4167 = N4131 & N4143;
  assign N4168 = N4131 & N4144;
  assign N4169 = N4131 & N4145;
  assign N4170 = N4132 & N4138;
  assign N4171 = N4132 & N4139;
  assign N4172 = N4132 & N4140;
  assign N4173 = N4132 & N4141;
  assign N4174 = N4132 & N4142;
  assign N4175 = N4132 & N4143;
  assign N4176 = N4132 & N4144;
  assign N4177 = N4132 & N4145;
  assign N4178 = w_addr_i[3] & w_addr_i[4];
  assign N4179 = N8 & w_addr_i[4];
  assign N8 = ~w_addr_i[3];
  assign N4180 = w_addr_i[3] & N9;
  assign N9 = ~w_addr_i[4];
  assign N4181 = N10 & N11;
  assign N10 = ~w_addr_i[3];
  assign N11 = ~w_addr_i[4];
  assign N4182 = ~w_addr_i[2];
  assign N4183 = w_addr_i[0] & w_addr_i[1];
  assign N4184 = N12 & w_addr_i[1];
  assign N12 = ~w_addr_i[0];
  assign N4185 = w_addr_i[0] & N13;
  assign N13 = ~w_addr_i[1];
  assign N4186 = N14 & N15;
  assign N14 = ~w_addr_i[0];
  assign N15 = ~w_addr_i[1];
  assign N4187 = w_addr_i[2] & N4183;
  assign N4188 = w_addr_i[2] & N4184;
  assign N4189 = w_addr_i[2] & N4185;
  assign N4190 = w_addr_i[2] & N4186;
  assign N4191 = N4182 & N4183;
  assign N4192 = N4182 & N4184;
  assign N4193 = N4182 & N4185;
  assign N4194 = N4182 & N4186;
  assign N4195 = N4178 & N4187;
  assign N4196 = N4178 & N4188;
  assign N4197 = N4178 & N4189;
  assign N4198 = N4178 & N4190;
  assign N4199 = N4178 & N4191;
  assign N4200 = N4178 & N4192;
  assign N4201 = N4178 & N4193;
  assign N4202 = N4178 & N4194;
  assign N4203 = N4179 & N4187;
  assign N4204 = N4179 & N4188;
  assign N4205 = N4179 & N4189;
  assign N4206 = N4179 & N4190;
  assign N4207 = N4179 & N4191;
  assign N4208 = N4179 & N4192;
  assign N4209 = N4179 & N4193;
  assign N4210 = N4179 & N4194;
  assign N4211 = N4180 & N4187;
  assign N4212 = N4180 & N4188;
  assign N4213 = N4180 & N4189;
  assign N4214 = N4180 & N4190;
  assign N4215 = N4180 & N4191;
  assign N4216 = N4180 & N4192;
  assign N4217 = N4180 & N4193;
  assign N4218 = N4180 & N4194;
  assign N4219 = N4181 & N4187;
  assign N4220 = N4181 & N4188;
  assign N4221 = N4181 & N4189;
  assign N4222 = N4181 & N4190;
  assign N4223 = N4181 & N4191;
  assign N4224 = N4181 & N4192;
  assign N4225 = N4181 & N4193;
  assign N4226 = N4181 & N4194;
  assign N1043 = N4146 & N4195;
  assign N1042 = N4146 & N4196;
  assign N1041 = N4146 & N4197;
  assign N1040 = N4146 & N4198;
  assign N1039 = N4146 & N4199;
  assign N1038 = N4146 & N4200;
  assign N1037 = N4146 & N4201;
  assign N1036 = N4146 & N4202;
  assign N1035 = N4146 & N4203;
  assign N1034 = N4146 & N4204;
  assign N1033 = N4146 & N4205;
  assign N1032 = N4146 & N4206;
  assign N1031 = N4146 & N4207;
  assign N1030 = N4146 & N4208;
  assign N1029 = N4146 & N4209;
  assign N1028 = N4146 & N4210;
  assign N1027 = N4146 & N4211;
  assign N1026 = N4146 & N4212;
  assign N1025 = N4146 & N4213;
  assign N1024 = N4146 & N4214;
  assign N1023 = N4146 & N4215;
  assign N1022 = N4146 & N4216;
  assign N1021 = N4146 & N4217;
  assign N1020 = N4146 & N4218;
  assign N1019 = N4146 & N4219;
  assign N1018 = N4146 & N4220;
  assign N1017 = N4146 & N4221;
  assign N1016 = N4146 & N4222;
  assign N1015 = N4146 & N4223;
  assign N1014 = N4146 & N4224;
  assign N1013 = N4146 & N4225;
  assign N1012 = N4146 & N4226;
  assign N1011 = N4147 & N4195;
  assign N1010 = N4147 & N4196;
  assign N1009 = N4147 & N4197;
  assign N1008 = N4147 & N4198;
  assign N1007 = N4147 & N4199;
  assign N1006 = N4147 & N4200;
  assign N1005 = N4147 & N4201;
  assign N1004 = N4147 & N4202;
  assign N1003 = N4147 & N4203;
  assign N1002 = N4147 & N4204;
  assign N1001 = N4147 & N4205;
  assign N1000 = N4147 & N4206;
  assign N999 = N4147 & N4207;
  assign N998 = N4147 & N4208;
  assign N997 = N4147 & N4209;
  assign N996 = N4147 & N4210;
  assign N995 = N4147 & N4211;
  assign N994 = N4147 & N4212;
  assign N993 = N4147 & N4213;
  assign N992 = N4147 & N4214;
  assign N991 = N4147 & N4215;
  assign N990 = N4147 & N4216;
  assign N989 = N4147 & N4217;
  assign N988 = N4147 & N4218;
  assign N987 = N4147 & N4219;
  assign N986 = N4147 & N4220;
  assign N985 = N4147 & N4221;
  assign N984 = N4147 & N4222;
  assign N983 = N4147 & N4223;
  assign N982 = N4147 & N4224;
  assign N981 = N4147 & N4225;
  assign N980 = N4147 & N4226;
  assign N979 = N4148 & N4195;
  assign N978 = N4148 & N4196;
  assign N977 = N4148 & N4197;
  assign N976 = N4148 & N4198;
  assign N975 = N4148 & N4199;
  assign N974 = N4148 & N4200;
  assign N973 = N4148 & N4201;
  assign N972 = N4148 & N4202;
  assign N971 = N4148 & N4203;
  assign N970 = N4148 & N4204;
  assign N969 = N4148 & N4205;
  assign N968 = N4148 & N4206;
  assign N967 = N4148 & N4207;
  assign N966 = N4148 & N4208;
  assign N965 = N4148 & N4209;
  assign N964 = N4148 & N4210;
  assign N963 = N4148 & N4211;
  assign N962 = N4148 & N4212;
  assign N961 = N4148 & N4213;
  assign N960 = N4148 & N4214;
  assign N959 = N4148 & N4215;
  assign N958 = N4148 & N4216;
  assign N957 = N4148 & N4217;
  assign N956 = N4148 & N4218;
  assign N955 = N4148 & N4219;
  assign N954 = N4148 & N4220;
  assign N953 = N4148 & N4221;
  assign N952 = N4148 & N4222;
  assign N951 = N4148 & N4223;
  assign N950 = N4148 & N4224;
  assign N949 = N4148 & N4225;
  assign N948 = N4148 & N4226;
  assign N947 = N4149 & N4195;
  assign N946 = N4149 & N4196;
  assign N945 = N4149 & N4197;
  assign N944 = N4149 & N4198;
  assign N943 = N4149 & N4199;
  assign N942 = N4149 & N4200;
  assign N941 = N4149 & N4201;
  assign N940 = N4149 & N4202;
  assign N939 = N4149 & N4203;
  assign N938 = N4149 & N4204;
  assign N937 = N4149 & N4205;
  assign N936 = N4149 & N4206;
  assign N935 = N4149 & N4207;
  assign N934 = N4149 & N4208;
  assign N933 = N4149 & N4209;
  assign N932 = N4149 & N4210;
  assign N931 = N4149 & N4211;
  assign N930 = N4149 & N4212;
  assign N929 = N4149 & N4213;
  assign N928 = N4149 & N4214;
  assign N927 = N4149 & N4215;
  assign N926 = N4149 & N4216;
  assign N925 = N4149 & N4217;
  assign N924 = N4149 & N4218;
  assign N923 = N4149 & N4219;
  assign N922 = N4149 & N4220;
  assign N921 = N4149 & N4221;
  assign N920 = N4149 & N4222;
  assign N919 = N4149 & N4223;
  assign N918 = N4149 & N4224;
  assign N917 = N4149 & N4225;
  assign N916 = N4149 & N4226;
  assign N915 = N4150 & N4195;
  assign N914 = N4150 & N4196;
  assign N913 = N4150 & N4197;
  assign N912 = N4150 & N4198;
  assign N911 = N4150 & N4199;
  assign N910 = N4150 & N4200;
  assign N909 = N4150 & N4201;
  assign N908 = N4150 & N4202;
  assign N907 = N4150 & N4203;
  assign N906 = N4150 & N4204;
  assign N905 = N4150 & N4205;
  assign N904 = N4150 & N4206;
  assign N903 = N4150 & N4207;
  assign N902 = N4150 & N4208;
  assign N901 = N4150 & N4209;
  assign N900 = N4150 & N4210;
  assign N899 = N4150 & N4211;
  assign N898 = N4150 & N4212;
  assign N897 = N4150 & N4213;
  assign N896 = N4150 & N4214;
  assign N895 = N4150 & N4215;
  assign N894 = N4150 & N4216;
  assign N893 = N4150 & N4217;
  assign N892 = N4150 & N4218;
  assign N891 = N4150 & N4219;
  assign N890 = N4150 & N4220;
  assign N889 = N4150 & N4221;
  assign N888 = N4150 & N4222;
  assign N887 = N4150 & N4223;
  assign N886 = N4150 & N4224;
  assign N885 = N4150 & N4225;
  assign N884 = N4150 & N4226;
  assign N883 = N4151 & N4195;
  assign N882 = N4151 & N4196;
  assign N881 = N4151 & N4197;
  assign N880 = N4151 & N4198;
  assign N879 = N4151 & N4199;
  assign N878 = N4151 & N4200;
  assign N877 = N4151 & N4201;
  assign N876 = N4151 & N4202;
  assign N875 = N4151 & N4203;
  assign N874 = N4151 & N4204;
  assign N873 = N4151 & N4205;
  assign N872 = N4151 & N4206;
  assign N871 = N4151 & N4207;
  assign N870 = N4151 & N4208;
  assign N869 = N4151 & N4209;
  assign N868 = N4151 & N4210;
  assign N867 = N4151 & N4211;
  assign N866 = N4151 & N4212;
  assign N865 = N4151 & N4213;
  assign N864 = N4151 & N4214;
  assign N863 = N4151 & N4215;
  assign N862 = N4151 & N4216;
  assign N861 = N4151 & N4217;
  assign N860 = N4151 & N4218;
  assign N859 = N4151 & N4219;
  assign N858 = N4151 & N4220;
  assign N857 = N4151 & N4221;
  assign N856 = N4151 & N4222;
  assign N855 = N4151 & N4223;
  assign N854 = N4151 & N4224;
  assign N853 = N4151 & N4225;
  assign N852 = N4151 & N4226;
  assign N851 = N4152 & N4195;
  assign N850 = N4152 & N4196;
  assign N849 = N4152 & N4197;
  assign N848 = N4152 & N4198;
  assign N847 = N4152 & N4199;
  assign N846 = N4152 & N4200;
  assign N845 = N4152 & N4201;
  assign N844 = N4152 & N4202;
  assign N843 = N4152 & N4203;
  assign N842 = N4152 & N4204;
  assign N841 = N4152 & N4205;
  assign N840 = N4152 & N4206;
  assign N839 = N4152 & N4207;
  assign N838 = N4152 & N4208;
  assign N837 = N4152 & N4209;
  assign N836 = N4152 & N4210;
  assign N835 = N4152 & N4211;
  assign N834 = N4152 & N4212;
  assign N833 = N4152 & N4213;
  assign N832 = N4152 & N4214;
  assign N831 = N4152 & N4215;
  assign N830 = N4152 & N4216;
  assign N829 = N4152 & N4217;
  assign N828 = N4152 & N4218;
  assign N827 = N4152 & N4219;
  assign N826 = N4152 & N4220;
  assign N825 = N4152 & N4221;
  assign N824 = N4152 & N4222;
  assign N823 = N4152 & N4223;
  assign N822 = N4152 & N4224;
  assign N821 = N4152 & N4225;
  assign N820 = N4152 & N4226;
  assign N819 = N4153 & N4195;
  assign N818 = N4153 & N4196;
  assign N817 = N4153 & N4197;
  assign N816 = N4153 & N4198;
  assign N815 = N4153 & N4199;
  assign N814 = N4153 & N4200;
  assign N813 = N4153 & N4201;
  assign N812 = N4153 & N4202;
  assign N811 = N4153 & N4203;
  assign N810 = N4153 & N4204;
  assign N809 = N4153 & N4205;
  assign N808 = N4153 & N4206;
  assign N807 = N4153 & N4207;
  assign N806 = N4153 & N4208;
  assign N805 = N4153 & N4209;
  assign N804 = N4153 & N4210;
  assign N803 = N4153 & N4211;
  assign N802 = N4153 & N4212;
  assign N801 = N4153 & N4213;
  assign N800 = N4153 & N4214;
  assign N799 = N4153 & N4215;
  assign N798 = N4153 & N4216;
  assign N797 = N4153 & N4217;
  assign N796 = N4153 & N4218;
  assign N795 = N4153 & N4219;
  assign N794 = N4153 & N4220;
  assign N793 = N4153 & N4221;
  assign N792 = N4153 & N4222;
  assign N791 = N4153 & N4223;
  assign N790 = N4153 & N4224;
  assign N789 = N4153 & N4225;
  assign N788 = N4153 & N4226;
  assign N787 = N4154 & N4195;
  assign N786 = N4154 & N4196;
  assign N785 = N4154 & N4197;
  assign N784 = N4154 & N4198;
  assign N783 = N4154 & N4199;
  assign N782 = N4154 & N4200;
  assign N781 = N4154 & N4201;
  assign N780 = N4154 & N4202;
  assign N779 = N4154 & N4203;
  assign N778 = N4154 & N4204;
  assign N777 = N4154 & N4205;
  assign N776 = N4154 & N4206;
  assign N775 = N4154 & N4207;
  assign N774 = N4154 & N4208;
  assign N773 = N4154 & N4209;
  assign N772 = N4154 & N4210;
  assign N771 = N4154 & N4211;
  assign N770 = N4154 & N4212;
  assign N769 = N4154 & N4213;
  assign N768 = N4154 & N4214;
  assign N767 = N4154 & N4215;
  assign N766 = N4154 & N4216;
  assign N765 = N4154 & N4217;
  assign N764 = N4154 & N4218;
  assign N763 = N4154 & N4219;
  assign N762 = N4154 & N4220;
  assign N761 = N4154 & N4221;
  assign N760 = N4154 & N4222;
  assign N759 = N4154 & N4223;
  assign N758 = N4154 & N4224;
  assign N757 = N4154 & N4225;
  assign N756 = N4154 & N4226;
  assign N755 = N4155 & N4195;
  assign N754 = N4155 & N4196;
  assign N753 = N4155 & N4197;
  assign N752 = N4155 & N4198;
  assign N751 = N4155 & N4199;
  assign N750 = N4155 & N4200;
  assign N749 = N4155 & N4201;
  assign N748 = N4155 & N4202;
  assign N747 = N4155 & N4203;
  assign N746 = N4155 & N4204;
  assign N745 = N4155 & N4205;
  assign N744 = N4155 & N4206;
  assign N743 = N4155 & N4207;
  assign N742 = N4155 & N4208;
  assign N741 = N4155 & N4209;
  assign N740 = N4155 & N4210;
  assign N739 = N4155 & N4211;
  assign N738 = N4155 & N4212;
  assign N737 = N4155 & N4213;
  assign N736 = N4155 & N4214;
  assign N735 = N4155 & N4215;
  assign N734 = N4155 & N4216;
  assign N733 = N4155 & N4217;
  assign N732 = N4155 & N4218;
  assign N731 = N4155 & N4219;
  assign N730 = N4155 & N4220;
  assign N729 = N4155 & N4221;
  assign N728 = N4155 & N4222;
  assign N727 = N4155 & N4223;
  assign N726 = N4155 & N4224;
  assign N725 = N4155 & N4225;
  assign N724 = N4155 & N4226;
  assign N723 = N4156 & N4195;
  assign N722 = N4156 & N4196;
  assign N721 = N4156 & N4197;
  assign N720 = N4156 & N4198;
  assign N719 = N4156 & N4199;
  assign N718 = N4156 & N4200;
  assign N717 = N4156 & N4201;
  assign N716 = N4156 & N4202;
  assign N715 = N4156 & N4203;
  assign N714 = N4156 & N4204;
  assign N713 = N4156 & N4205;
  assign N712 = N4156 & N4206;
  assign N711 = N4156 & N4207;
  assign N710 = N4156 & N4208;
  assign N709 = N4156 & N4209;
  assign N708 = N4156 & N4210;
  assign N707 = N4156 & N4211;
  assign N706 = N4156 & N4212;
  assign N705 = N4156 & N4213;
  assign N704 = N4156 & N4214;
  assign N703 = N4156 & N4215;
  assign N702 = N4156 & N4216;
  assign N701 = N4156 & N4217;
  assign N700 = N4156 & N4218;
  assign N699 = N4156 & N4219;
  assign N698 = N4156 & N4220;
  assign N697 = N4156 & N4221;
  assign N696 = N4156 & N4222;
  assign N695 = N4156 & N4223;
  assign N694 = N4156 & N4224;
  assign N693 = N4156 & N4225;
  assign N692 = N4156 & N4226;
  assign N691 = N4157 & N4195;
  assign N690 = N4157 & N4196;
  assign N689 = N4157 & N4197;
  assign N688 = N4157 & N4198;
  assign N687 = N4157 & N4199;
  assign N686 = N4157 & N4200;
  assign N685 = N4157 & N4201;
  assign N684 = N4157 & N4202;
  assign N683 = N4157 & N4203;
  assign N682 = N4157 & N4204;
  assign N681 = N4157 & N4205;
  assign N680 = N4157 & N4206;
  assign N679 = N4157 & N4207;
  assign N678 = N4157 & N4208;
  assign N677 = N4157 & N4209;
  assign N676 = N4157 & N4210;
  assign N675 = N4157 & N4211;
  assign N674 = N4157 & N4212;
  assign N673 = N4157 & N4213;
  assign N672 = N4157 & N4214;
  assign N671 = N4157 & N4215;
  assign N670 = N4157 & N4216;
  assign N669 = N4157 & N4217;
  assign N668 = N4157 & N4218;
  assign N667 = N4157 & N4219;
  assign N666 = N4157 & N4220;
  assign N665 = N4157 & N4221;
  assign N664 = N4157 & N4222;
  assign N663 = N4157 & N4223;
  assign N662 = N4157 & N4224;
  assign N661 = N4157 & N4225;
  assign N660 = N4157 & N4226;
  assign N659 = N4158 & N4195;
  assign N658 = N4158 & N4196;
  assign N657 = N4158 & N4197;
  assign N656 = N4158 & N4198;
  assign N655 = N4158 & N4199;
  assign N654 = N4158 & N4200;
  assign N653 = N4158 & N4201;
  assign N652 = N4158 & N4202;
  assign N651 = N4158 & N4203;
  assign N650 = N4158 & N4204;
  assign N649 = N4158 & N4205;
  assign N648 = N4158 & N4206;
  assign N647 = N4158 & N4207;
  assign N646 = N4158 & N4208;
  assign N645 = N4158 & N4209;
  assign N644 = N4158 & N4210;
  assign N643 = N4158 & N4211;
  assign N642 = N4158 & N4212;
  assign N641 = N4158 & N4213;
  assign N640 = N4158 & N4214;
  assign N639 = N4158 & N4215;
  assign N638 = N4158 & N4216;
  assign N637 = N4158 & N4217;
  assign N636 = N4158 & N4218;
  assign N635 = N4158 & N4219;
  assign N634 = N4158 & N4220;
  assign N633 = N4158 & N4221;
  assign N632 = N4158 & N4222;
  assign N631 = N4158 & N4223;
  assign N630 = N4158 & N4224;
  assign N629 = N4158 & N4225;
  assign N628 = N4158 & N4226;
  assign N627 = N4159 & N4195;
  assign N626 = N4159 & N4196;
  assign N625 = N4159 & N4197;
  assign N624 = N4159 & N4198;
  assign N623 = N4159 & N4199;
  assign N622 = N4159 & N4200;
  assign N621 = N4159 & N4201;
  assign N620 = N4159 & N4202;
  assign N619 = N4159 & N4203;
  assign N618 = N4159 & N4204;
  assign N617 = N4159 & N4205;
  assign N616 = N4159 & N4206;
  assign N615 = N4159 & N4207;
  assign N614 = N4159 & N4208;
  assign N613 = N4159 & N4209;
  assign N612 = N4159 & N4210;
  assign N611 = N4159 & N4211;
  assign N610 = N4159 & N4212;
  assign N609 = N4159 & N4213;
  assign N608 = N4159 & N4214;
  assign N607 = N4159 & N4215;
  assign N606 = N4159 & N4216;
  assign N605 = N4159 & N4217;
  assign N604 = N4159 & N4218;
  assign N603 = N4159 & N4219;
  assign N602 = N4159 & N4220;
  assign N601 = N4159 & N4221;
  assign N600 = N4159 & N4222;
  assign N599 = N4159 & N4223;
  assign N598 = N4159 & N4224;
  assign N597 = N4159 & N4225;
  assign N596 = N4159 & N4226;
  assign N595 = N4160 & N4195;
  assign N594 = N4160 & N4196;
  assign N593 = N4160 & N4197;
  assign N592 = N4160 & N4198;
  assign N591 = N4160 & N4199;
  assign N590 = N4160 & N4200;
  assign N589 = N4160 & N4201;
  assign N588 = N4160 & N4202;
  assign N587 = N4160 & N4203;
  assign N586 = N4160 & N4204;
  assign N585 = N4160 & N4205;
  assign N584 = N4160 & N4206;
  assign N583 = N4160 & N4207;
  assign N582 = N4160 & N4208;
  assign N581 = N4160 & N4209;
  assign N580 = N4160 & N4210;
  assign N579 = N4160 & N4211;
  assign N578 = N4160 & N4212;
  assign N577 = N4160 & N4213;
  assign N576 = N4160 & N4214;
  assign N575 = N4160 & N4215;
  assign N574 = N4160 & N4216;
  assign N573 = N4160 & N4217;
  assign N572 = N4160 & N4218;
  assign N571 = N4160 & N4219;
  assign N570 = N4160 & N4220;
  assign N569 = N4160 & N4221;
  assign N568 = N4160 & N4222;
  assign N567 = N4160 & N4223;
  assign N566 = N4160 & N4224;
  assign N565 = N4160 & N4225;
  assign N564 = N4160 & N4226;
  assign N563 = N4161 & N4195;
  assign N562 = N4161 & N4196;
  assign N561 = N4161 & N4197;
  assign N560 = N4161 & N4198;
  assign N559 = N4161 & N4199;
  assign N558 = N4161 & N4200;
  assign N557 = N4161 & N4201;
  assign N556 = N4161 & N4202;
  assign N555 = N4161 & N4203;
  assign N554 = N4161 & N4204;
  assign N553 = N4161 & N4205;
  assign N552 = N4161 & N4206;
  assign N551 = N4161 & N4207;
  assign N550 = N4161 & N4208;
  assign N549 = N4161 & N4209;
  assign N548 = N4161 & N4210;
  assign N547 = N4161 & N4211;
  assign N546 = N4161 & N4212;
  assign N545 = N4161 & N4213;
  assign N544 = N4161 & N4214;
  assign N543 = N4161 & N4215;
  assign N542 = N4161 & N4216;
  assign N541 = N4161 & N4217;
  assign N540 = N4161 & N4218;
  assign N539 = N4161 & N4219;
  assign N538 = N4161 & N4220;
  assign N537 = N4161 & N4221;
  assign N536 = N4161 & N4222;
  assign N535 = N4161 & N4223;
  assign N534 = N4161 & N4224;
  assign N533 = N4161 & N4225;
  assign N532 = N4161 & N4226;
  assign N531 = N4162 & N4195;
  assign N530 = N4162 & N4196;
  assign N529 = N4162 & N4197;
  assign N528 = N4162 & N4198;
  assign N527 = N4162 & N4199;
  assign N526 = N4162 & N4200;
  assign N525 = N4162 & N4201;
  assign N524 = N4162 & N4202;
  assign N523 = N4162 & N4203;
  assign N522 = N4162 & N4204;
  assign N521 = N4162 & N4205;
  assign N520 = N4162 & N4206;
  assign N519 = N4162 & N4207;
  assign N518 = N4162 & N4208;
  assign N517 = N4162 & N4209;
  assign N516 = N4162 & N4210;
  assign N515 = N4162 & N4211;
  assign N514 = N4162 & N4212;
  assign N513 = N4162 & N4213;
  assign N512 = N4162 & N4214;
  assign N511 = N4162 & N4215;
  assign N510 = N4162 & N4216;
  assign N509 = N4162 & N4217;
  assign N508 = N4162 & N4218;
  assign N507 = N4162 & N4219;
  assign N506 = N4162 & N4220;
  assign N505 = N4162 & N4221;
  assign N504 = N4162 & N4222;
  assign N503 = N4162 & N4223;
  assign N502 = N4162 & N4224;
  assign N501 = N4162 & N4225;
  assign N500 = N4162 & N4226;
  assign N499 = N4163 & N4195;
  assign N498 = N4163 & N4196;
  assign N497 = N4163 & N4197;
  assign N496 = N4163 & N4198;
  assign N495 = N4163 & N4199;
  assign N494 = N4163 & N4200;
  assign N493 = N4163 & N4201;
  assign N492 = N4163 & N4202;
  assign N491 = N4163 & N4203;
  assign N490 = N4163 & N4204;
  assign N489 = N4163 & N4205;
  assign N488 = N4163 & N4206;
  assign N487 = N4163 & N4207;
  assign N486 = N4163 & N4208;
  assign N485 = N4163 & N4209;
  assign N484 = N4163 & N4210;
  assign N483 = N4163 & N4211;
  assign N482 = N4163 & N4212;
  assign N481 = N4163 & N4213;
  assign N480 = N4163 & N4214;
  assign N479 = N4163 & N4215;
  assign N478 = N4163 & N4216;
  assign N477 = N4163 & N4217;
  assign N476 = N4163 & N4218;
  assign N475 = N4163 & N4219;
  assign N474 = N4163 & N4220;
  assign N473 = N4163 & N4221;
  assign N472 = N4163 & N4222;
  assign N471 = N4163 & N4223;
  assign N470 = N4163 & N4224;
  assign N469 = N4163 & N4225;
  assign N468 = N4163 & N4226;
  assign N467 = N4164 & N4195;
  assign N466 = N4164 & N4196;
  assign N465 = N4164 & N4197;
  assign N464 = N4164 & N4198;
  assign N463 = N4164 & N4199;
  assign N462 = N4164 & N4200;
  assign N461 = N4164 & N4201;
  assign N460 = N4164 & N4202;
  assign N459 = N4164 & N4203;
  assign N458 = N4164 & N4204;
  assign N457 = N4164 & N4205;
  assign N456 = N4164 & N4206;
  assign N455 = N4164 & N4207;
  assign N454 = N4164 & N4208;
  assign N453 = N4164 & N4209;
  assign N452 = N4164 & N4210;
  assign N451 = N4164 & N4211;
  assign N450 = N4164 & N4212;
  assign N449 = N4164 & N4213;
  assign N448 = N4164 & N4214;
  assign N447 = N4164 & N4215;
  assign N446 = N4164 & N4216;
  assign N445 = N4164 & N4217;
  assign N444 = N4164 & N4218;
  assign N443 = N4164 & N4219;
  assign N442 = N4164 & N4220;
  assign N441 = N4164 & N4221;
  assign N440 = N4164 & N4222;
  assign N439 = N4164 & N4223;
  assign N438 = N4164 & N4224;
  assign N437 = N4164 & N4225;
  assign N436 = N4164 & N4226;
  assign N435 = N4165 & N4195;
  assign N434 = N4165 & N4196;
  assign N433 = N4165 & N4197;
  assign N432 = N4165 & N4198;
  assign N431 = N4165 & N4199;
  assign N430 = N4165 & N4200;
  assign N429 = N4165 & N4201;
  assign N428 = N4165 & N4202;
  assign N427 = N4165 & N4203;
  assign N426 = N4165 & N4204;
  assign N425 = N4165 & N4205;
  assign N424 = N4165 & N4206;
  assign N423 = N4165 & N4207;
  assign N422 = N4165 & N4208;
  assign N421 = N4165 & N4209;
  assign N420 = N4165 & N4210;
  assign N419 = N4165 & N4211;
  assign N418 = N4165 & N4212;
  assign N417 = N4165 & N4213;
  assign N416 = N4165 & N4214;
  assign N415 = N4165 & N4215;
  assign N414 = N4165 & N4216;
  assign N413 = N4165 & N4217;
  assign N412 = N4165 & N4218;
  assign N411 = N4165 & N4219;
  assign N410 = N4165 & N4220;
  assign N409 = N4165 & N4221;
  assign N408 = N4165 & N4222;
  assign N407 = N4165 & N4223;
  assign N406 = N4165 & N4224;
  assign N405 = N4165 & N4225;
  assign N404 = N4165 & N4226;
  assign N403 = N4166 & N4195;
  assign N402 = N4166 & N4196;
  assign N401 = N4166 & N4197;
  assign N400 = N4166 & N4198;
  assign N399 = N4166 & N4199;
  assign N398 = N4166 & N4200;
  assign N397 = N4166 & N4201;
  assign N396 = N4166 & N4202;
  assign N395 = N4166 & N4203;
  assign N394 = N4166 & N4204;
  assign N393 = N4166 & N4205;
  assign N392 = N4166 & N4206;
  assign N391 = N4166 & N4207;
  assign N390 = N4166 & N4208;
  assign N389 = N4166 & N4209;
  assign N388 = N4166 & N4210;
  assign N387 = N4166 & N4211;
  assign N386 = N4166 & N4212;
  assign N385 = N4166 & N4213;
  assign N384 = N4166 & N4214;
  assign N383 = N4166 & N4215;
  assign N382 = N4166 & N4216;
  assign N381 = N4166 & N4217;
  assign N380 = N4166 & N4218;
  assign N379 = N4166 & N4219;
  assign N378 = N4166 & N4220;
  assign N377 = N4166 & N4221;
  assign N376 = N4166 & N4222;
  assign N375 = N4166 & N4223;
  assign N374 = N4166 & N4224;
  assign N373 = N4166 & N4225;
  assign N372 = N4166 & N4226;
  assign N371 = N4167 & N4195;
  assign N370 = N4167 & N4196;
  assign N369 = N4167 & N4197;
  assign N368 = N4167 & N4198;
  assign N367 = N4167 & N4199;
  assign N366 = N4167 & N4200;
  assign N365 = N4167 & N4201;
  assign N364 = N4167 & N4202;
  assign N363 = N4167 & N4203;
  assign N362 = N4167 & N4204;
  assign N361 = N4167 & N4205;
  assign N360 = N4167 & N4206;
  assign N359 = N4167 & N4207;
  assign N358 = N4167 & N4208;
  assign N357 = N4167 & N4209;
  assign N356 = N4167 & N4210;
  assign N355 = N4167 & N4211;
  assign N354 = N4167 & N4212;
  assign N353 = N4167 & N4213;
  assign N352 = N4167 & N4214;
  assign N351 = N4167 & N4215;
  assign N350 = N4167 & N4216;
  assign N349 = N4167 & N4217;
  assign N348 = N4167 & N4218;
  assign N347 = N4167 & N4219;
  assign N346 = N4167 & N4220;
  assign N345 = N4167 & N4221;
  assign N344 = N4167 & N4222;
  assign N343 = N4167 & N4223;
  assign N342 = N4167 & N4224;
  assign N341 = N4167 & N4225;
  assign N340 = N4167 & N4226;
  assign N339 = N4168 & N4195;
  assign N338 = N4168 & N4196;
  assign N337 = N4168 & N4197;
  assign N336 = N4168 & N4198;
  assign N335 = N4168 & N4199;
  assign N334 = N4168 & N4200;
  assign N333 = N4168 & N4201;
  assign N332 = N4168 & N4202;
  assign N331 = N4168 & N4203;
  assign N330 = N4168 & N4204;
  assign N329 = N4168 & N4205;
  assign N328 = N4168 & N4206;
  assign N327 = N4168 & N4207;
  assign N326 = N4168 & N4208;
  assign N325 = N4168 & N4209;
  assign N324 = N4168 & N4210;
  assign N323 = N4168 & N4211;
  assign N322 = N4168 & N4212;
  assign N321 = N4168 & N4213;
  assign N320 = N4168 & N4214;
  assign N319 = N4168 & N4215;
  assign N318 = N4168 & N4216;
  assign N317 = N4168 & N4217;
  assign N316 = N4168 & N4218;
  assign N315 = N4168 & N4219;
  assign N314 = N4168 & N4220;
  assign N313 = N4168 & N4221;
  assign N312 = N4168 & N4222;
  assign N311 = N4168 & N4223;
  assign N310 = N4168 & N4224;
  assign N309 = N4168 & N4225;
  assign N308 = N4168 & N4226;
  assign N307 = N4169 & N4195;
  assign N306 = N4169 & N4196;
  assign N305 = N4169 & N4197;
  assign N304 = N4169 & N4198;
  assign N303 = N4169 & N4199;
  assign N302 = N4169 & N4200;
  assign N301 = N4169 & N4201;
  assign N300 = N4169 & N4202;
  assign N299 = N4169 & N4203;
  assign N298 = N4169 & N4204;
  assign N297 = N4169 & N4205;
  assign N296 = N4169 & N4206;
  assign N295 = N4169 & N4207;
  assign N294 = N4169 & N4208;
  assign N293 = N4169 & N4209;
  assign N292 = N4169 & N4210;
  assign N291 = N4169 & N4211;
  assign N290 = N4169 & N4212;
  assign N289 = N4169 & N4213;
  assign N288 = N4169 & N4214;
  assign N287 = N4169 & N4215;
  assign N286 = N4169 & N4216;
  assign N285 = N4169 & N4217;
  assign N284 = N4169 & N4218;
  assign N283 = N4169 & N4219;
  assign N282 = N4169 & N4220;
  assign N281 = N4169 & N4221;
  assign N280 = N4169 & N4222;
  assign N279 = N4169 & N4223;
  assign N278 = N4169 & N4224;
  assign N277 = N4169 & N4225;
  assign N276 = N4169 & N4226;
  assign N275 = N4170 & N4195;
  assign N274 = N4170 & N4196;
  assign N273 = N4170 & N4197;
  assign N272 = N4170 & N4198;
  assign N271 = N4170 & N4199;
  assign N270 = N4170 & N4200;
  assign N269 = N4170 & N4201;
  assign N268 = N4170 & N4202;
  assign N267 = N4170 & N4203;
  assign N266 = N4170 & N4204;
  assign N265 = N4170 & N4205;
  assign N264 = N4170 & N4206;
  assign N263 = N4170 & N4207;
  assign N262 = N4170 & N4208;
  assign N261 = N4170 & N4209;
  assign N260 = N4170 & N4210;
  assign N259 = N4170 & N4211;
  assign N258 = N4170 & N4212;
  assign N257 = N4170 & N4213;
  assign N256 = N4170 & N4214;
  assign N255 = N4170 & N4215;
  assign N254 = N4170 & N4216;
  assign N253 = N4170 & N4217;
  assign N252 = N4170 & N4218;
  assign N251 = N4170 & N4219;
  assign N250 = N4170 & N4220;
  assign N249 = N4170 & N4221;
  assign N248 = N4170 & N4222;
  assign N247 = N4170 & N4223;
  assign N246 = N4170 & N4224;
  assign N245 = N4170 & N4225;
  assign N244 = N4170 & N4226;
  assign N243 = N4171 & N4195;
  assign N242 = N4171 & N4196;
  assign N241 = N4171 & N4197;
  assign N240 = N4171 & N4198;
  assign N239 = N4171 & N4199;
  assign N238 = N4171 & N4200;
  assign N237 = N4171 & N4201;
  assign N236 = N4171 & N4202;
  assign N235 = N4171 & N4203;
  assign N234 = N4171 & N4204;
  assign N233 = N4171 & N4205;
  assign N232 = N4171 & N4206;
  assign N231 = N4171 & N4207;
  assign N230 = N4171 & N4208;
  assign N229 = N4171 & N4209;
  assign N228 = N4171 & N4210;
  assign N227 = N4171 & N4211;
  assign N226 = N4171 & N4212;
  assign N225 = N4171 & N4213;
  assign N224 = N4171 & N4214;
  assign N223 = N4171 & N4215;
  assign N222 = N4171 & N4216;
  assign N221 = N4171 & N4217;
  assign N220 = N4171 & N4218;
  assign N219 = N4171 & N4219;
  assign N218 = N4171 & N4220;
  assign N217 = N4171 & N4221;
  assign N216 = N4171 & N4222;
  assign N215 = N4171 & N4223;
  assign N214 = N4171 & N4224;
  assign N213 = N4171 & N4225;
  assign N212 = N4171 & N4226;
  assign N211 = N4172 & N4195;
  assign N210 = N4172 & N4196;
  assign N209 = N4172 & N4197;
  assign N208 = N4172 & N4198;
  assign N207 = N4172 & N4199;
  assign N206 = N4172 & N4200;
  assign N205 = N4172 & N4201;
  assign N204 = N4172 & N4202;
  assign N203 = N4172 & N4203;
  assign N202 = N4172 & N4204;
  assign N201 = N4172 & N4205;
  assign N200 = N4172 & N4206;
  assign N199 = N4172 & N4207;
  assign N198 = N4172 & N4208;
  assign N197 = N4172 & N4209;
  assign N196 = N4172 & N4210;
  assign N195 = N4172 & N4211;
  assign N194 = N4172 & N4212;
  assign N193 = N4172 & N4213;
  assign N192 = N4172 & N4214;
  assign N191 = N4172 & N4215;
  assign N190 = N4172 & N4216;
  assign N189 = N4172 & N4217;
  assign N188 = N4172 & N4218;
  assign N187 = N4172 & N4219;
  assign N186 = N4172 & N4220;
  assign N185 = N4172 & N4221;
  assign N184 = N4172 & N4222;
  assign N183 = N4172 & N4223;
  assign N182 = N4172 & N4224;
  assign N181 = N4172 & N4225;
  assign N180 = N4172 & N4226;
  assign N179 = N4173 & N4195;
  assign N178 = N4173 & N4196;
  assign N177 = N4173 & N4197;
  assign N176 = N4173 & N4198;
  assign N175 = N4173 & N4199;
  assign N174 = N4173 & N4200;
  assign N173 = N4173 & N4201;
  assign N172 = N4173 & N4202;
  assign N171 = N4173 & N4203;
  assign N170 = N4173 & N4204;
  assign N169 = N4173 & N4205;
  assign N168 = N4173 & N4206;
  assign N167 = N4173 & N4207;
  assign N166 = N4173 & N4208;
  assign N165 = N4173 & N4209;
  assign N164 = N4173 & N4210;
  assign N163 = N4173 & N4211;
  assign N162 = N4173 & N4212;
  assign N161 = N4173 & N4213;
  assign N160 = N4173 & N4214;
  assign N159 = N4173 & N4215;
  assign N158 = N4173 & N4216;
  assign N157 = N4173 & N4217;
  assign N156 = N4173 & N4218;
  assign N155 = N4173 & N4219;
  assign N154 = N4173 & N4220;
  assign N153 = N4173 & N4221;
  assign N152 = N4173 & N4222;
  assign N151 = N4173 & N4223;
  assign N150 = N4173 & N4224;
  assign N149 = N4173 & N4225;
  assign N148 = N4173 & N4226;
  assign N147 = N4174 & N4195;
  assign N146 = N4174 & N4196;
  assign N145 = N4174 & N4197;
  assign N144 = N4174 & N4198;
  assign N143 = N4174 & N4199;
  assign N142 = N4174 & N4200;
  assign N141 = N4174 & N4201;
  assign N140 = N4174 & N4202;
  assign N139 = N4174 & N4203;
  assign N138 = N4174 & N4204;
  assign N137 = N4174 & N4205;
  assign N136 = N4174 & N4206;
  assign N135 = N4174 & N4207;
  assign N134 = N4174 & N4208;
  assign N133 = N4174 & N4209;
  assign N132 = N4174 & N4210;
  assign N131 = N4174 & N4211;
  assign N130 = N4174 & N4212;
  assign N129 = N4174 & N4213;
  assign N128 = N4174 & N4214;
  assign N127 = N4174 & N4215;
  assign N126 = N4174 & N4216;
  assign N125 = N4174 & N4217;
  assign N124 = N4174 & N4218;
  assign N123 = N4174 & N4219;
  assign N122 = N4174 & N4220;
  assign N121 = N4174 & N4221;
  assign N120 = N4174 & N4222;
  assign N119 = N4174 & N4223;
  assign N118 = N4174 & N4224;
  assign N117 = N4174 & N4225;
  assign N116 = N4174 & N4226;
  assign N115 = N4175 & N4195;
  assign N114 = N4175 & N4196;
  assign N113 = N4175 & N4197;
  assign N112 = N4175 & N4198;
  assign N111 = N4175 & N4199;
  assign N110 = N4175 & N4200;
  assign N109 = N4175 & N4201;
  assign N108 = N4175 & N4202;
  assign N107 = N4175 & N4203;
  assign N106 = N4175 & N4204;
  assign N105 = N4175 & N4205;
  assign N104 = N4175 & N4206;
  assign N103 = N4175 & N4207;
  assign N102 = N4175 & N4208;
  assign N101 = N4175 & N4209;
  assign N100 = N4175 & N4210;
  assign N99 = N4175 & N4211;
  assign N98 = N4175 & N4212;
  assign N97 = N4175 & N4213;
  assign N96 = N4175 & N4214;
  assign N95 = N4175 & N4215;
  assign N94 = N4175 & N4216;
  assign N93 = N4175 & N4217;
  assign N92 = N4175 & N4218;
  assign N91 = N4175 & N4219;
  assign N90 = N4175 & N4220;
  assign N89 = N4175 & N4221;
  assign N88 = N4175 & N4222;
  assign N87 = N4175 & N4223;
  assign N86 = N4175 & N4224;
  assign N85 = N4175 & N4225;
  assign N84 = N4175 & N4226;
  assign N83 = N4176 & N4195;
  assign N82 = N4176 & N4196;
  assign N81 = N4176 & N4197;
  assign N80 = N4176 & N4198;
  assign N79 = N4176 & N4199;
  assign N78 = N4176 & N4200;
  assign N77 = N4176 & N4201;
  assign N76 = N4176 & N4202;
  assign N75 = N4176 & N4203;
  assign N74 = N4176 & N4204;
  assign N73 = N4176 & N4205;
  assign N72 = N4176 & N4206;
  assign N71 = N4176 & N4207;
  assign N70 = N4176 & N4208;
  assign N69 = N4176 & N4209;
  assign N68 = N4176 & N4210;
  assign N67 = N4176 & N4211;
  assign N66 = N4176 & N4212;
  assign N65 = N4176 & N4213;
  assign N64 = N4176 & N4214;
  assign N63 = N4176 & N4215;
  assign N62 = N4176 & N4216;
  assign N61 = N4176 & N4217;
  assign N60 = N4176 & N4218;
  assign N59 = N4176 & N4219;
  assign N58 = N4176 & N4220;
  assign N57 = N4176 & N4221;
  assign N56 = N4176 & N4222;
  assign N55 = N4176 & N4223;
  assign N54 = N4176 & N4224;
  assign N53 = N4176 & N4225;
  assign N52 = N4176 & N4226;
  assign N51 = N4177 & N4195;
  assign N50 = N4177 & N4196;
  assign N49 = N4177 & N4197;
  assign N48 = N4177 & N4198;
  assign N47 = N4177 & N4199;
  assign N46 = N4177 & N4200;
  assign N45 = N4177 & N4201;
  assign N44 = N4177 & N4202;
  assign N43 = N4177 & N4203;
  assign N42 = N4177 & N4204;
  assign N41 = N4177 & N4205;
  assign N40 = N4177 & N4206;
  assign N39 = N4177 & N4207;
  assign N38 = N4177 & N4208;
  assign N37 = N4177 & N4209;
  assign N36 = N4177 & N4210;
  assign N35 = N4177 & N4211;
  assign N34 = N4177 & N4212;
  assign N33 = N4177 & N4213;
  assign N32 = N4177 & N4214;
  assign N31 = N4177 & N4215;
  assign N30 = N4177 & N4216;
  assign N29 = N4177 & N4217;
  assign N28 = N4177 & N4218;
  assign N27 = N4177 & N4219;
  assign N26 = N4177 & N4220;
  assign N25 = N4177 & N4221;
  assign N24 = N4177 & N4222;
  assign N23 = N4177 & N4223;
  assign N22 = N4177 & N4224;
  assign N21 = N4177 & N4225;
  assign N20 = N4177 & N4226;
  assign { N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2071, N2070, N2069, N2068, N2067, N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057, N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047, N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037, N2036, N2035, N2034, N2033, N2032, N2031, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987, N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977, N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967, N1966, N1965, N1964, N1963, N1962, N1961, N1960, N1959, N1958, N1957, N1956, N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946, N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N1930, N1929, N1928, N1927, N1926, N1925, N1924, N1923, N1922, N1921, N1920, N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, N1899, N1898, N1897, N1896, N1895, N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886, N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876, N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866, N1865, N1864, N1863, N1862, N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N1830, N1829, N1828, N1827, N1826, N1825, N1824, N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814, N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804, N1803, N1802, N1801, N1800, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, N1790, N1789, N1788, N1787, N1786, N1785, N1784, N1783, N1782, N1781, N1780, N1779, N1778, N1777, N1776, N1775, N1774, N1773, N1772, N1771, N1770, N1769, N1768, N1767, N1766, N1765, N1764, N1763, N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735, N1734, N1733, N1732, N1731, N1730, N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722, N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712, N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702, N1701, N1700, N1699, N1698, N1697, N1696, N1695, N1694, N1693, N1692, N1691, N1690, N1689, N1688, N1687, N1686, N1685, N1684, N1683, N1682, N1681, N1680, N1679, N1678, N1677, N1676, N1675, N1674, N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, N1660, N1659, N1658, N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648, N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638, N1637, N1636, N1635, N1634, N1633, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624, N1623, N1622, N1621, N1620, N1619, N1618, N1617, N1616, N1615, N1614, N1613, N1612, N1611, N1610, N1609, N1608, N1607, N1606, N1605, N1604, N1603, N1602, N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1594, N1593, N1592, N1591, N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581, N1580, N1579, N1578, N1577, N1576, N1575, N1574, N1573, N1572, N1571, N1570, N1569, N1568, N1567, N1566, N1565, N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555, N1554, N1553, N1552, N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532, N1531, N1530, N1529, N1528, N1527, N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517, N1516, N1515, N1514, N1513, N1512, N1511, N1510, N1509, N1508, N1507, N1506, N1505, N1504, N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494, N1493, N1492, N1491, N1490, N1489, N1488, N1487, N1486, N1485, N1484, N1483, N1482, N1481, N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471, N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461, N1460, N1459, N1458, N1457, N1456, N1455, N1454, N1453, N1452, N1451, N1450, N1449, N1448, N1447, N1446, N1445, N1444, N1443, N1442, N1441, N1440, N1439, N1438, N1437, N1436, N1435, N1434, N1433, N1432, N1431, N1430, N1429, N1428, N1427, N1426, N1425, N1424, N1423, N1422, N1421, N1420, N1419, N1418, N1417, N1416, N1415, N1414, N1413, N1412, N1411, N1410, N1409, N1408, N1407, N1406, N1405, N1404, N1403, N1402, N1401, N1400, N1399, N1398, N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1388, N1387, N1386, N1385, N1384, N1383, N1382, N1381, N1380, N1379, N1378, N1377, N1376, N1375, N1374, N1373, N1372, N1371, N1370, N1369, N1368, N1367, N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, N1356, N1355, N1354, N1353, N1352, N1351, N1350, N1349, N1348, N1347, N1346, N1345, N1344, N1343, N1342, N1341, N1340, N1339, N1338, N1337, N1336, N1335, N1334, N1333, N1332, N1331, N1330, N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N1320, N1319, N1318, N1317, N1316, N1315, N1314, N1313, N1312, N1311, N1310, N1309, N1308, N1307, N1306, N1305, N1304, N1303, N1302, N1301, N1300, N1299, N1298, N1297, N1296, N1295, N1294, N1293, N1292, N1291, N1290, N1289, N1288, N1287, N1286, N1285, N1284, N1283, N1282, N1281, N1280, N1279, N1278, N1277, N1276, N1275, N1274, N1273, N1272, N1271, N1270, N1269, N1268, N1267, N1266, N1265, N1264, N1263, N1262, N1261, N1260, N1259, N1258, N1257, N1256, N1255, N1254, N1253, N1252, N1251, N1250, N1249, N1248, N1247, N1246, N1245, N1244, N1243, N1242, N1241, N1240, N1239, N1238, N1237, N1236, N1235, N1234, N1233, N1232, N1231, N1230, N1229, N1228, N1227, N1226, N1225, N1224, N1223, N1222, N1221, N1220, N1219, N1218, N1217, N1216, N1215, N1214, N1213, N1212, N1211, N1210, N1209, N1208, N1207, N1206, N1205, N1204, N1203, N1202, N1201, N1200, N1199, N1198, N1197, N1196, N1195, N1194, N1193, N1192, N1191, N1190, N1189, N1188, N1187, N1186, N1185, N1184, N1183, N1182, N1181, N1180, N1179, N1178, N1177, N1176, N1175, N1174, N1173, N1172, N1171, N1170, N1169, N1168, N1167, N1166, N1165, N1164, N1163, N1162, N1161, N1160, N1159, N1158, N1157, N1156, N1155, N1154, N1153, N1152, N1151, N1150, N1149, N1148, N1147, N1146, N1145, N1144, N1143, N1142, N1141, N1140, N1139, N1138, N1137, N1136, N1135, N1134, N1133, N1132, N1131, N1130, N1129, N1128, N1127, N1126, N1125, N1124, N1123, N1122, N1121, N1120, N1119, N1118, N1117, N1116, N1115, N1114, N1113, N1112, N1111, N1110, N1109, N1108, N1107, N1106, N1105, N1104, N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1064, N1062, N1060, N1058, N1056, N1054, N1052, N1050, N1048, N1046, N1044 } = (N16)? { 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3104)? { N1043, N1042, N1041, N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, N1002, N1001, N1000, N999, N998, N997, N996, N995, N994, N993, N992, N991, N990, N989, N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, N940, N939, N938, N937, N936, N935, N934, N933, N932, N931, N930, N929, N928, N927, N926, N925, N924, N923, N922, N921, N920, N919, N918, N917, N916, N915, N914, N913, N912, N911, N910, N909, N908, N907, N906, N905, N904, N903, N902, N901, N900, N899, N898, N897, N896, N895, N894, N893, N892, N891, N890, N889, N888, N887, N886, N885, N884, N883, N882, N881, N880, N879, N878, N877, N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, N864, N863, N862, N861, N860, N859, N858, N857, N856, N855, N854, N853, N852, N851, N850, N849, N848, N847, N846, N845, N844, N843, N842, N841, N840, N839, N838, N837, N836, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N805, N804, N803, N802, N801, N800, N799, N798, N797, N796, N795, N794, N793, N792, N791, N790, N789, N788, N787, N786, N785, N784, N783, N782, N781, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, N527, N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, N514, N513, N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, N265, N264, N263, N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign N16 = reset_i;
  assign { N1065, N1063, N1061, N1059, N1057, N1055, N1053, N1051, N1049, N1047, N1045 } = (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                           (N3104)? { w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i, w_set_not_clear_i } : 1'b0;
  assign { N3102, N3101, N3100, N3099, N3098, N3097, N3096, N3095, N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081, N3080, N3079, N3078, N3077, N3076, N3075, N3074, N3073, N3072, N3071, N3070, N3069, N3068, N3067, N3066, N3065, N3064, N3063, N3062, N3061, N3060, N3059, N3058, N3057, N3056, N3055, N3054, N3053, N3052, N3051, N3050, N3049, N3048, N3047, N3046, N3045, N3044, N3043, N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, N3023, N3022, N3021, N3020, N3019, N3018, N3017, N3016, N3015, N3014, N3013, N3012, N3011, N3010, N3009, N3008, N3007, N3006, N3005, N3004, N3003, N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989, N2988, N2987, N2986, N2985, N2984, N2983, N2982, N2981, N2980, N2979, N2978, N2977, N2976, N2975, N2974, N2973, N2972, N2971, N2970, N2969, N2968, N2967, N2966, N2965, N2964, N2963, N2962, N2961, N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, N2940, N2939, N2938, N2937, N2936, N2935, N2934, N2933, N2932, N2931, N2930, N2929, N2928, N2927, N2926, N2925, N2924, N2923, N2922, N2921, N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907, N2906, N2905, N2904, N2903, N2902, N2901, N2900, N2899, N2898, N2897, N2896, N2895, N2894, N2893, N2892, N2891, N2890, N2889, N2888, N2887, N2886, N2885, N2884, N2883, N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, N2848, N2847, N2846, N2845, N2844, N2843, N2842, N2841, N2840, N2839, N2838, N2837, N2836, N2835, N2834, N2833, N2832, N2831, N2830, N2829, N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815, N2814, N2813, N2812, N2811, N2810, N2809, N2808, N2807, N2806, N2805, N2804, N2803, N2802, N2801, N2800, N2799, N2798, N2797, N2796, N2795, N2794, N2793, N2792, N2791, N2790, N2789, N2788, N2787, N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, N2766, N2765, N2764, N2763, N2762, N2761, N2760, N2759, N2758, N2757, N2756, N2755, N2754, N2753, N2752, N2751, N2750, N2749, N2748, N2747, N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733, N2732, N2731, N2730, N2729, N2728, N2727, N2726, N2725, N2724, N2723, N2722, N2721, N2720, N2719, N2718, N2717, N2716, N2715, N2714, N2713, N2712, N2711, N2710, N2709, N2708, N2707, N2706, N2705, N2704, N2703, N2702, N2701, N2700, N2699, N2698, N2697, N2696, N2695, N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661, N2660, N2659, N2658, N2657, N2656, N2655, N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641, N2640, N2639, N2638, N2637, N2636, N2635, N2634, N2633, N2632, N2631, N2630, N2629, N2628, N2627, N2626, N2625, N2624, N2623, N2622, N2621, N2620, N2619, N2618, N2617, N2616, N2615, N2614, N2613, N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, N2592, N2591, N2590, N2589, N2588, N2587, N2586, N2585, N2584, N2583, N2582, N2581, N2580, N2579, N2578, N2577, N2576, N2575, N2574, N2573, N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559, N2558, N2557, N2556, N2555, N2554, N2553, N2552, N2551, N2550, N2549, N2548, N2547, N2546, N2545, N2544, N2543, N2542, N2541, N2540, N2539, N2538, N2537, N2536, N2535, N2534, N2533, N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515, N2514, N2513, N2512, N2511, N2510, N2509, N2508, N2507, N2506, N2505, N2504, N2503, N2502, N2501, N2500, N2499, N2498, N2497, N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463, N2462, N2461, N2460, N2459, N2458, N2457, N2456, N2455, N2454, N2453, N2452, N2451, N2450, N2449, N2448, N2447, N2446, N2445, N2444, N2443, N2442, N2441, N2440, N2439, N2438, N2437, N2436, N2435, N2434, N2433, N2432, N2431, N2430, N2429, N2428, N2427, N2426, N2425, N2424, N2423, N2422, N2421, N2420, N2419, N2418, N2417, N2416, N2415, N2414, N2413, N2412, N2411, N2410, N2409, N2408, N2407, N2406, N2405, N2404, N2403, N2402, N2401, N2400, N2399, N2398, N2397, N2396, N2395, N2394, N2393, N2392, N2391, N2390, N2389, N2388, N2387, N2386, N2385, N2384, N2383, N2382, N2381, N2380, N2379, N2378, N2377, N2376, N2375, N2374, N2373, N2372, N2371, N2370, N2369, N2368, N2367, N2366, N2365, N2364, N2363, N2362, N2361, N2360, N2359, N2358, N2357, N2356, N2355, N2354, N2353, N2352, N2351, N2350, N2349, N2348, N2347, N2346, N2345, N2344, N2343, N2342, N2341, N2340, N2339, N2338, N2337, N2336, N2335, N2334, N2333, N2332, N2331, N2330, N2329, N2328, N2327, N2326, N2325, N2324, N2323, N2322, N2321, N2320, N2319, N2318, N2317, N2316, N2315, N2314, N2313, N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, N2275, N2274, N2273, N2272, N2271, N2270, N2269, N2268, N2267, N2266, N2265, N2264, N2263, N2262, N2261, N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243, N2242, N2241, N2240, N2239, N2238, N2237, N2236, N2235, N2234, N2233, N2232, N2231, N2230, N2229, N2228, N2227, N2226, N2225, N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197, N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2188, N2187, N2186, N2185, N2184, N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2145, N2144, N2143, N2142, N2141, N2140, N2139, N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129, N2128, N2127, N2126, N2125, N2124, N2123, N2122, N2121, N2120, N2119, N2118, N2117, N2116, N2115, N2114, N2113, N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081, N2080, N2079 } = (N16)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N3104)? { N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043 } : 
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              (N19)? { 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0 } : 1'b0;
  assign r_v_o = N4227 & matched;
  assign N4227 = en_i & r_v_i;
  assign empty_v_o = en_i & empty_found;
  assign N17 = en_i & w_v_i;
  assign N18 = N17 | reset_i;
  assign N19 = ~N18;
  assign N3103 = ~reset_i;
  assign N3104 = N17 & N3103;
  assign match_array[0] = N4230 & valid[0];
  assign N4230 = N4229 & N3105;
  assign N4229 = N4228 & en_i;
  assign N4228 = ~reset_i;
  assign empty_array[0] = N4231 & N4232;
  assign N4231 = N4228 & en_i;
  assign N4232 = ~valid[0];
  assign match_array[1] = N4234 & valid[1];
  assign N4234 = N4233 & N3106;
  assign N4233 = N4228 & en_i;
  assign empty_array[1] = N4235 & N4236;
  assign N4235 = N4228 & en_i;
  assign N4236 = ~valid[1];
  assign match_array[2] = N4238 & valid[2];
  assign N4238 = N4237 & N3107;
  assign N4237 = N4228 & en_i;
  assign empty_array[2] = N4239 & N4240;
  assign N4239 = N4228 & en_i;
  assign N4240 = ~valid[2];
  assign match_array[3] = N4242 & valid[3];
  assign N4242 = N4241 & N3108;
  assign N4241 = N4228 & en_i;
  assign empty_array[3] = N4243 & N4244;
  assign N4243 = N4228 & en_i;
  assign N4244 = ~valid[3];
  assign match_array[4] = N4246 & valid[4];
  assign N4246 = N4245 & N3109;
  assign N4245 = N4228 & en_i;
  assign empty_array[4] = N4247 & N4248;
  assign N4247 = N4228 & en_i;
  assign N4248 = ~valid[4];
  assign match_array[5] = N4250 & valid[5];
  assign N4250 = N4249 & N3110;
  assign N4249 = N4228 & en_i;
  assign empty_array[5] = N4251 & N4252;
  assign N4251 = N4228 & en_i;
  assign N4252 = ~valid[5];
  assign match_array[6] = N4254 & valid[6];
  assign N4254 = N4253 & N3111;
  assign N4253 = N4228 & en_i;
  assign empty_array[6] = N4255 & N4256;
  assign N4255 = N4228 & en_i;
  assign N4256 = ~valid[6];
  assign match_array[7] = N4258 & valid[7];
  assign N4258 = N4257 & N3112;
  assign N4257 = N4228 & en_i;
  assign empty_array[7] = N4259 & N4260;
  assign N4259 = N4228 & en_i;
  assign N4260 = ~valid[7];
  assign match_array[8] = N4262 & valid[8];
  assign N4262 = N4261 & N3113;
  assign N4261 = N4228 & en_i;
  assign empty_array[8] = N4263 & N4264;
  assign N4263 = N4228 & en_i;
  assign N4264 = ~valid[8];
  assign match_array[9] = N4266 & valid[9];
  assign N4266 = N4265 & N3114;
  assign N4265 = N4228 & en_i;
  assign empty_array[9] = N4267 & N4268;
  assign N4267 = N4228 & en_i;
  assign N4268 = ~valid[9];
  assign match_array[10] = N4270 & valid[10];
  assign N4270 = N4269 & N3115;
  assign N4269 = N4228 & en_i;
  assign empty_array[10] = N4271 & N4272;
  assign N4271 = N4228 & en_i;
  assign N4272 = ~valid[10];
  assign match_array[11] = N4274 & valid[11];
  assign N4274 = N4273 & N3116;
  assign N4273 = N4228 & en_i;
  assign empty_array[11] = N4275 & N4276;
  assign N4275 = N4228 & en_i;
  assign N4276 = ~valid[11];
  assign match_array[12] = N4278 & valid[12];
  assign N4278 = N4277 & N3117;
  assign N4277 = N4228 & en_i;
  assign empty_array[12] = N4279 & N4280;
  assign N4279 = N4228 & en_i;
  assign N4280 = ~valid[12];
  assign match_array[13] = N4282 & valid[13];
  assign N4282 = N4281 & N3118;
  assign N4281 = N4228 & en_i;
  assign empty_array[13] = N4283 & N4284;
  assign N4283 = N4228 & en_i;
  assign N4284 = ~valid[13];
  assign match_array[14] = N4286 & valid[14];
  assign N4286 = N4285 & N3119;
  assign N4285 = N4228 & en_i;
  assign empty_array[14] = N4287 & N4288;
  assign N4287 = N4228 & en_i;
  assign N4288 = ~valid[14];
  assign match_array[15] = N4290 & valid[15];
  assign N4290 = N4289 & N3120;
  assign N4289 = N4228 & en_i;
  assign empty_array[15] = N4291 & N4292;
  assign N4291 = N4228 & en_i;
  assign N4292 = ~valid[15];
  assign match_array[16] = N4294 & valid[16];
  assign N4294 = N4293 & N3121;
  assign N4293 = N4228 & en_i;
  assign empty_array[16] = N4295 & N4296;
  assign N4295 = N4228 & en_i;
  assign N4296 = ~valid[16];
  assign match_array[17] = N4298 & valid[17];
  assign N4298 = N4297 & N3122;
  assign N4297 = N4228 & en_i;
  assign empty_array[17] = N4299 & N4300;
  assign N4299 = N4228 & en_i;
  assign N4300 = ~valid[17];
  assign match_array[18] = N4302 & valid[18];
  assign N4302 = N4301 & N3123;
  assign N4301 = N4228 & en_i;
  assign empty_array[18] = N4303 & N4304;
  assign N4303 = N4228 & en_i;
  assign N4304 = ~valid[18];
  assign match_array[19] = N4306 & valid[19];
  assign N4306 = N4305 & N3124;
  assign N4305 = N4228 & en_i;
  assign empty_array[19] = N4307 & N4308;
  assign N4307 = N4228 & en_i;
  assign N4308 = ~valid[19];
  assign match_array[20] = N4310 & valid[20];
  assign N4310 = N4309 & N3125;
  assign N4309 = N4228 & en_i;
  assign empty_array[20] = N4311 & N4312;
  assign N4311 = N4228 & en_i;
  assign N4312 = ~valid[20];
  assign match_array[21] = N4314 & valid[21];
  assign N4314 = N4313 & N3126;
  assign N4313 = N4228 & en_i;
  assign empty_array[21] = N4315 & N4316;
  assign N4315 = N4228 & en_i;
  assign N4316 = ~valid[21];
  assign match_array[22] = N4318 & valid[22];
  assign N4318 = N4317 & N3127;
  assign N4317 = N4228 & en_i;
  assign empty_array[22] = N4319 & N4320;
  assign N4319 = N4228 & en_i;
  assign N4320 = ~valid[22];
  assign match_array[23] = N4322 & valid[23];
  assign N4322 = N4321 & N3128;
  assign N4321 = N4228 & en_i;
  assign empty_array[23] = N4323 & N4324;
  assign N4323 = N4228 & en_i;
  assign N4324 = ~valid[23];
  assign match_array[24] = N4326 & valid[24];
  assign N4326 = N4325 & N3129;
  assign N4325 = N4228 & en_i;
  assign empty_array[24] = N4327 & N4328;
  assign N4327 = N4228 & en_i;
  assign N4328 = ~valid[24];
  assign match_array[25] = N4330 & valid[25];
  assign N4330 = N4329 & N3130;
  assign N4329 = N4228 & en_i;
  assign empty_array[25] = N4331 & N4332;
  assign N4331 = N4228 & en_i;
  assign N4332 = ~valid[25];
  assign match_array[26] = N4334 & valid[26];
  assign N4334 = N4333 & N3131;
  assign N4333 = N4228 & en_i;
  assign empty_array[26] = N4335 & N4336;
  assign N4335 = N4228 & en_i;
  assign N4336 = ~valid[26];
  assign match_array[27] = N4338 & valid[27];
  assign N4338 = N4337 & N3132;
  assign N4337 = N4228 & en_i;
  assign empty_array[27] = N4339 & N4340;
  assign N4339 = N4228 & en_i;
  assign N4340 = ~valid[27];
  assign match_array[28] = N4342 & valid[28];
  assign N4342 = N4341 & N3133;
  assign N4341 = N4228 & en_i;
  assign empty_array[28] = N4343 & N4344;
  assign N4343 = N4228 & en_i;
  assign N4344 = ~valid[28];
  assign match_array[29] = N4346 & valid[29];
  assign N4346 = N4345 & N3134;
  assign N4345 = N4228 & en_i;
  assign empty_array[29] = N4347 & N4348;
  assign N4347 = N4228 & en_i;
  assign N4348 = ~valid[29];
  assign match_array[30] = N4350 & valid[30];
  assign N4350 = N4349 & N3135;
  assign N4349 = N4228 & en_i;
  assign empty_array[30] = N4351 & N4352;
  assign N4351 = N4228 & en_i;
  assign N4352 = ~valid[30];
  assign match_array[31] = N4354 & valid[31];
  assign N4354 = N4353 & N3136;
  assign N4353 = N4228 & en_i;
  assign empty_array[31] = N4355 & N4356;
  assign N4355 = N4228 & en_i;
  assign N4356 = ~valid[31];
  assign match_array[32] = N4358 & valid[32];
  assign N4358 = N4357 & N3137;
  assign N4357 = N4228 & en_i;
  assign empty_array[32] = N4359 & N4360;
  assign N4359 = N4228 & en_i;
  assign N4360 = ~valid[32];
  assign match_array[33] = N4362 & valid[33];
  assign N4362 = N4361 & N3138;
  assign N4361 = N4228 & en_i;
  assign empty_array[33] = N4363 & N4364;
  assign N4363 = N4228 & en_i;
  assign N4364 = ~valid[33];
  assign match_array[34] = N4366 & valid[34];
  assign N4366 = N4365 & N3139;
  assign N4365 = N4228 & en_i;
  assign empty_array[34] = N4367 & N4368;
  assign N4367 = N4228 & en_i;
  assign N4368 = ~valid[34];
  assign match_array[35] = N4370 & valid[35];
  assign N4370 = N4369 & N3140;
  assign N4369 = N4228 & en_i;
  assign empty_array[35] = N4371 & N4372;
  assign N4371 = N4228 & en_i;
  assign N4372 = ~valid[35];
  assign match_array[36] = N4374 & valid[36];
  assign N4374 = N4373 & N3141;
  assign N4373 = N4228 & en_i;
  assign empty_array[36] = N4375 & N4376;
  assign N4375 = N4228 & en_i;
  assign N4376 = ~valid[36];
  assign match_array[37] = N4378 & valid[37];
  assign N4378 = N4377 & N3142;
  assign N4377 = N4228 & en_i;
  assign empty_array[37] = N4379 & N4380;
  assign N4379 = N4228 & en_i;
  assign N4380 = ~valid[37];
  assign match_array[38] = N4382 & valid[38];
  assign N4382 = N4381 & N3143;
  assign N4381 = N4228 & en_i;
  assign empty_array[38] = N4383 & N4384;
  assign N4383 = N4228 & en_i;
  assign N4384 = ~valid[38];
  assign match_array[39] = N4386 & valid[39];
  assign N4386 = N4385 & N3144;
  assign N4385 = N4228 & en_i;
  assign empty_array[39] = N4387 & N4388;
  assign N4387 = N4228 & en_i;
  assign N4388 = ~valid[39];
  assign match_array[40] = N4390 & valid[40];
  assign N4390 = N4389 & N3145;
  assign N4389 = N4228 & en_i;
  assign empty_array[40] = N4391 & N4392;
  assign N4391 = N4228 & en_i;
  assign N4392 = ~valid[40];
  assign match_array[41] = N4394 & valid[41];
  assign N4394 = N4393 & N3146;
  assign N4393 = N4228 & en_i;
  assign empty_array[41] = N4395 & N4396;
  assign N4395 = N4228 & en_i;
  assign N4396 = ~valid[41];
  assign match_array[42] = N4398 & valid[42];
  assign N4398 = N4397 & N3147;
  assign N4397 = N4228 & en_i;
  assign empty_array[42] = N4399 & N4400;
  assign N4399 = N4228 & en_i;
  assign N4400 = ~valid[42];
  assign match_array[43] = N4402 & valid[43];
  assign N4402 = N4401 & N3148;
  assign N4401 = N4228 & en_i;
  assign empty_array[43] = N4403 & N4404;
  assign N4403 = N4228 & en_i;
  assign N4404 = ~valid[43];
  assign match_array[44] = N4406 & valid[44];
  assign N4406 = N4405 & N3149;
  assign N4405 = N4228 & en_i;
  assign empty_array[44] = N4407 & N4408;
  assign N4407 = N4228 & en_i;
  assign N4408 = ~valid[44];
  assign match_array[45] = N4410 & valid[45];
  assign N4410 = N4409 & N3150;
  assign N4409 = N4228 & en_i;
  assign empty_array[45] = N4411 & N4412;
  assign N4411 = N4228 & en_i;
  assign N4412 = ~valid[45];
  assign match_array[46] = N4414 & valid[46];
  assign N4414 = N4413 & N3151;
  assign N4413 = N4228 & en_i;
  assign empty_array[46] = N4415 & N4416;
  assign N4415 = N4228 & en_i;
  assign N4416 = ~valid[46];
  assign match_array[47] = N4418 & valid[47];
  assign N4418 = N4417 & N3152;
  assign N4417 = N4228 & en_i;
  assign empty_array[47] = N4419 & N4420;
  assign N4419 = N4228 & en_i;
  assign N4420 = ~valid[47];
  assign match_array[48] = N4422 & valid[48];
  assign N4422 = N4421 & N3153;
  assign N4421 = N4228 & en_i;
  assign empty_array[48] = N4423 & N4424;
  assign N4423 = N4228 & en_i;
  assign N4424 = ~valid[48];
  assign match_array[49] = N4426 & valid[49];
  assign N4426 = N4425 & N3154;
  assign N4425 = N4228 & en_i;
  assign empty_array[49] = N4427 & N4428;
  assign N4427 = N4228 & en_i;
  assign N4428 = ~valid[49];
  assign match_array[50] = N4430 & valid[50];
  assign N4430 = N4429 & N3155;
  assign N4429 = N4228 & en_i;
  assign empty_array[50] = N4431 & N4432;
  assign N4431 = N4228 & en_i;
  assign N4432 = ~valid[50];
  assign match_array[51] = N4434 & valid[51];
  assign N4434 = N4433 & N3156;
  assign N4433 = N4228 & en_i;
  assign empty_array[51] = N4435 & N4436;
  assign N4435 = N4228 & en_i;
  assign N4436 = ~valid[51];
  assign match_array[52] = N4438 & valid[52];
  assign N4438 = N4437 & N3157;
  assign N4437 = N4228 & en_i;
  assign empty_array[52] = N4439 & N4440;
  assign N4439 = N4228 & en_i;
  assign N4440 = ~valid[52];
  assign match_array[53] = N4442 & valid[53];
  assign N4442 = N4441 & N3158;
  assign N4441 = N4228 & en_i;
  assign empty_array[53] = N4443 & N4444;
  assign N4443 = N4228 & en_i;
  assign N4444 = ~valid[53];
  assign match_array[54] = N4446 & valid[54];
  assign N4446 = N4445 & N3159;
  assign N4445 = N4228 & en_i;
  assign empty_array[54] = N4447 & N4448;
  assign N4447 = N4228 & en_i;
  assign N4448 = ~valid[54];
  assign match_array[55] = N4450 & valid[55];
  assign N4450 = N4449 & N3160;
  assign N4449 = N4228 & en_i;
  assign empty_array[55] = N4451 & N4452;
  assign N4451 = N4228 & en_i;
  assign N4452 = ~valid[55];
  assign match_array[56] = N4454 & valid[56];
  assign N4454 = N4453 & N3161;
  assign N4453 = N4228 & en_i;
  assign empty_array[56] = N4455 & N4456;
  assign N4455 = N4228 & en_i;
  assign N4456 = ~valid[56];
  assign match_array[57] = N4458 & valid[57];
  assign N4458 = N4457 & N3162;
  assign N4457 = N4228 & en_i;
  assign empty_array[57] = N4459 & N4460;
  assign N4459 = N4228 & en_i;
  assign N4460 = ~valid[57];
  assign match_array[58] = N4462 & valid[58];
  assign N4462 = N4461 & N3163;
  assign N4461 = N4228 & en_i;
  assign empty_array[58] = N4463 & N4464;
  assign N4463 = N4228 & en_i;
  assign N4464 = ~valid[58];
  assign match_array[59] = N4466 & valid[59];
  assign N4466 = N4465 & N3164;
  assign N4465 = N4228 & en_i;
  assign empty_array[59] = N4467 & N4468;
  assign N4467 = N4228 & en_i;
  assign N4468 = ~valid[59];
  assign match_array[60] = N4470 & valid[60];
  assign N4470 = N4469 & N3165;
  assign N4469 = N4228 & en_i;
  assign empty_array[60] = N4471 & N4472;
  assign N4471 = N4228 & en_i;
  assign N4472 = ~valid[60];
  assign match_array[61] = N4474 & valid[61];
  assign N4474 = N4473 & N3166;
  assign N4473 = N4228 & en_i;
  assign empty_array[61] = N4475 & N4476;
  assign N4475 = N4228 & en_i;
  assign N4476 = ~valid[61];
  assign match_array[62] = N4478 & valid[62];
  assign N4478 = N4477 & N3167;
  assign N4477 = N4228 & en_i;
  assign empty_array[62] = N4479 & N4480;
  assign N4479 = N4228 & en_i;
  assign N4480 = ~valid[62];
  assign match_array[63] = N4482 & valid[63];
  assign N4482 = N4481 & N3168;
  assign N4481 = N4228 & en_i;
  assign empty_array[63] = N4483 & N4484;
  assign N4483 = N4228 & en_i;
  assign N4484 = ~valid[63];
  assign match_array[64] = N4486 & valid[64];
  assign N4486 = N4485 & N3169;
  assign N4485 = N4228 & en_i;
  assign empty_array[64] = N4487 & N4488;
  assign N4487 = N4228 & en_i;
  assign N4488 = ~valid[64];
  assign match_array[65] = N4490 & valid[65];
  assign N4490 = N4489 & N3170;
  assign N4489 = N4228 & en_i;
  assign empty_array[65] = N4491 & N4492;
  assign N4491 = N4228 & en_i;
  assign N4492 = ~valid[65];
  assign match_array[66] = N4494 & valid[66];
  assign N4494 = N4493 & N3171;
  assign N4493 = N4228 & en_i;
  assign empty_array[66] = N4495 & N4496;
  assign N4495 = N4228 & en_i;
  assign N4496 = ~valid[66];
  assign match_array[67] = N4498 & valid[67];
  assign N4498 = N4497 & N3172;
  assign N4497 = N4228 & en_i;
  assign empty_array[67] = N4499 & N4500;
  assign N4499 = N4228 & en_i;
  assign N4500 = ~valid[67];
  assign match_array[68] = N4502 & valid[68];
  assign N4502 = N4501 & N3173;
  assign N4501 = N4228 & en_i;
  assign empty_array[68] = N4503 & N4504;
  assign N4503 = N4228 & en_i;
  assign N4504 = ~valid[68];
  assign match_array[69] = N4506 & valid[69];
  assign N4506 = N4505 & N3174;
  assign N4505 = N4228 & en_i;
  assign empty_array[69] = N4507 & N4508;
  assign N4507 = N4228 & en_i;
  assign N4508 = ~valid[69];
  assign match_array[70] = N4510 & valid[70];
  assign N4510 = N4509 & N3175;
  assign N4509 = N4228 & en_i;
  assign empty_array[70] = N4511 & N4512;
  assign N4511 = N4228 & en_i;
  assign N4512 = ~valid[70];
  assign match_array[71] = N4514 & valid[71];
  assign N4514 = N4513 & N3176;
  assign N4513 = N4228 & en_i;
  assign empty_array[71] = N4515 & N4516;
  assign N4515 = N4228 & en_i;
  assign N4516 = ~valid[71];
  assign match_array[72] = N4518 & valid[72];
  assign N4518 = N4517 & N3177;
  assign N4517 = N4228 & en_i;
  assign empty_array[72] = N4519 & N4520;
  assign N4519 = N4228 & en_i;
  assign N4520 = ~valid[72];
  assign match_array[73] = N4522 & valid[73];
  assign N4522 = N4521 & N3178;
  assign N4521 = N4228 & en_i;
  assign empty_array[73] = N4523 & N4524;
  assign N4523 = N4228 & en_i;
  assign N4524 = ~valid[73];
  assign match_array[74] = N4526 & valid[74];
  assign N4526 = N4525 & N3179;
  assign N4525 = N4228 & en_i;
  assign empty_array[74] = N4527 & N4528;
  assign N4527 = N4228 & en_i;
  assign N4528 = ~valid[74];
  assign match_array[75] = N4530 & valid[75];
  assign N4530 = N4529 & N3180;
  assign N4529 = N4228 & en_i;
  assign empty_array[75] = N4531 & N4532;
  assign N4531 = N4228 & en_i;
  assign N4532 = ~valid[75];
  assign match_array[76] = N4534 & valid[76];
  assign N4534 = N4533 & N3181;
  assign N4533 = N4228 & en_i;
  assign empty_array[76] = N4535 & N4536;
  assign N4535 = N4228 & en_i;
  assign N4536 = ~valid[76];
  assign match_array[77] = N4538 & valid[77];
  assign N4538 = N4537 & N3182;
  assign N4537 = N4228 & en_i;
  assign empty_array[77] = N4539 & N4540;
  assign N4539 = N4228 & en_i;
  assign N4540 = ~valid[77];
  assign match_array[78] = N4542 & valid[78];
  assign N4542 = N4541 & N3183;
  assign N4541 = N4228 & en_i;
  assign empty_array[78] = N4543 & N4544;
  assign N4543 = N4228 & en_i;
  assign N4544 = ~valid[78];
  assign match_array[79] = N4546 & valid[79];
  assign N4546 = N4545 & N3184;
  assign N4545 = N4228 & en_i;
  assign empty_array[79] = N4547 & N4548;
  assign N4547 = N4228 & en_i;
  assign N4548 = ~valid[79];
  assign match_array[80] = N4550 & valid[80];
  assign N4550 = N4549 & N3185;
  assign N4549 = N4228 & en_i;
  assign empty_array[80] = N4551 & N4552;
  assign N4551 = N4228 & en_i;
  assign N4552 = ~valid[80];
  assign match_array[81] = N4554 & valid[81];
  assign N4554 = N4553 & N3186;
  assign N4553 = N4228 & en_i;
  assign empty_array[81] = N4555 & N4556;
  assign N4555 = N4228 & en_i;
  assign N4556 = ~valid[81];
  assign match_array[82] = N4558 & valid[82];
  assign N4558 = N4557 & N3187;
  assign N4557 = N4228 & en_i;
  assign empty_array[82] = N4559 & N4560;
  assign N4559 = N4228 & en_i;
  assign N4560 = ~valid[82];
  assign match_array[83] = N4562 & valid[83];
  assign N4562 = N4561 & N3188;
  assign N4561 = N4228 & en_i;
  assign empty_array[83] = N4563 & N4564;
  assign N4563 = N4228 & en_i;
  assign N4564 = ~valid[83];
  assign match_array[84] = N4566 & valid[84];
  assign N4566 = N4565 & N3189;
  assign N4565 = N4228 & en_i;
  assign empty_array[84] = N4567 & N4568;
  assign N4567 = N4228 & en_i;
  assign N4568 = ~valid[84];
  assign match_array[85] = N4570 & valid[85];
  assign N4570 = N4569 & N3190;
  assign N4569 = N4228 & en_i;
  assign empty_array[85] = N4571 & N4572;
  assign N4571 = N4228 & en_i;
  assign N4572 = ~valid[85];
  assign match_array[86] = N4574 & valid[86];
  assign N4574 = N4573 & N3191;
  assign N4573 = N4228 & en_i;
  assign empty_array[86] = N4575 & N4576;
  assign N4575 = N4228 & en_i;
  assign N4576 = ~valid[86];
  assign match_array[87] = N4578 & valid[87];
  assign N4578 = N4577 & N3192;
  assign N4577 = N4228 & en_i;
  assign empty_array[87] = N4579 & N4580;
  assign N4579 = N4228 & en_i;
  assign N4580 = ~valid[87];
  assign match_array[88] = N4582 & valid[88];
  assign N4582 = N4581 & N3193;
  assign N4581 = N4228 & en_i;
  assign empty_array[88] = N4583 & N4584;
  assign N4583 = N4228 & en_i;
  assign N4584 = ~valid[88];
  assign match_array[89] = N4586 & valid[89];
  assign N4586 = N4585 & N3194;
  assign N4585 = N4228 & en_i;
  assign empty_array[89] = N4587 & N4588;
  assign N4587 = N4228 & en_i;
  assign N4588 = ~valid[89];
  assign match_array[90] = N4590 & valid[90];
  assign N4590 = N4589 & N3195;
  assign N4589 = N4228 & en_i;
  assign empty_array[90] = N4591 & N4592;
  assign N4591 = N4228 & en_i;
  assign N4592 = ~valid[90];
  assign match_array[91] = N4594 & valid[91];
  assign N4594 = N4593 & N3196;
  assign N4593 = N4228 & en_i;
  assign empty_array[91] = N4595 & N4596;
  assign N4595 = N4228 & en_i;
  assign N4596 = ~valid[91];
  assign match_array[92] = N4598 & valid[92];
  assign N4598 = N4597 & N3197;
  assign N4597 = N4228 & en_i;
  assign empty_array[92] = N4599 & N4600;
  assign N4599 = N4228 & en_i;
  assign N4600 = ~valid[92];
  assign match_array[93] = N4602 & valid[93];
  assign N4602 = N4601 & N3198;
  assign N4601 = N4228 & en_i;
  assign empty_array[93] = N4603 & N4604;
  assign N4603 = N4228 & en_i;
  assign N4604 = ~valid[93];
  assign match_array[94] = N4606 & valid[94];
  assign N4606 = N4605 & N3199;
  assign N4605 = N4228 & en_i;
  assign empty_array[94] = N4607 & N4608;
  assign N4607 = N4228 & en_i;
  assign N4608 = ~valid[94];
  assign match_array[95] = N4610 & valid[95];
  assign N4610 = N4609 & N3200;
  assign N4609 = N4228 & en_i;
  assign empty_array[95] = N4611 & N4612;
  assign N4611 = N4228 & en_i;
  assign N4612 = ~valid[95];
  assign match_array[96] = N4614 & valid[96];
  assign N4614 = N4613 & N3201;
  assign N4613 = N4228 & en_i;
  assign empty_array[96] = N4615 & N4616;
  assign N4615 = N4228 & en_i;
  assign N4616 = ~valid[96];
  assign match_array[97] = N4618 & valid[97];
  assign N4618 = N4617 & N3202;
  assign N4617 = N4228 & en_i;
  assign empty_array[97] = N4619 & N4620;
  assign N4619 = N4228 & en_i;
  assign N4620 = ~valid[97];
  assign match_array[98] = N4622 & valid[98];
  assign N4622 = N4621 & N3203;
  assign N4621 = N4228 & en_i;
  assign empty_array[98] = N4623 & N4624;
  assign N4623 = N4228 & en_i;
  assign N4624 = ~valid[98];
  assign match_array[99] = N4626 & valid[99];
  assign N4626 = N4625 & N3204;
  assign N4625 = N4228 & en_i;
  assign empty_array[99] = N4627 & N4628;
  assign N4627 = N4228 & en_i;
  assign N4628 = ~valid[99];
  assign match_array[100] = N4630 & valid[100];
  assign N4630 = N4629 & N3205;
  assign N4629 = N4228 & en_i;
  assign empty_array[100] = N4631 & N4632;
  assign N4631 = N4228 & en_i;
  assign N4632 = ~valid[100];
  assign match_array[101] = N4634 & valid[101];
  assign N4634 = N4633 & N3206;
  assign N4633 = N4228 & en_i;
  assign empty_array[101] = N4635 & N4636;
  assign N4635 = N4228 & en_i;
  assign N4636 = ~valid[101];
  assign match_array[102] = N4638 & valid[102];
  assign N4638 = N4637 & N3207;
  assign N4637 = N4228 & en_i;
  assign empty_array[102] = N4639 & N4640;
  assign N4639 = N4228 & en_i;
  assign N4640 = ~valid[102];
  assign match_array[103] = N4642 & valid[103];
  assign N4642 = N4641 & N3208;
  assign N4641 = N4228 & en_i;
  assign empty_array[103] = N4643 & N4644;
  assign N4643 = N4228 & en_i;
  assign N4644 = ~valid[103];
  assign match_array[104] = N4646 & valid[104];
  assign N4646 = N4645 & N3209;
  assign N4645 = N4228 & en_i;
  assign empty_array[104] = N4647 & N4648;
  assign N4647 = N4228 & en_i;
  assign N4648 = ~valid[104];
  assign match_array[105] = N4650 & valid[105];
  assign N4650 = N4649 & N3210;
  assign N4649 = N4228 & en_i;
  assign empty_array[105] = N4651 & N4652;
  assign N4651 = N4228 & en_i;
  assign N4652 = ~valid[105];
  assign match_array[106] = N4654 & valid[106];
  assign N4654 = N4653 & N3211;
  assign N4653 = N4228 & en_i;
  assign empty_array[106] = N4655 & N4656;
  assign N4655 = N4228 & en_i;
  assign N4656 = ~valid[106];
  assign match_array[107] = N4658 & valid[107];
  assign N4658 = N4657 & N3212;
  assign N4657 = N4228 & en_i;
  assign empty_array[107] = N4659 & N4660;
  assign N4659 = N4228 & en_i;
  assign N4660 = ~valid[107];
  assign match_array[108] = N4662 & valid[108];
  assign N4662 = N4661 & N3213;
  assign N4661 = N4228 & en_i;
  assign empty_array[108] = N4663 & N4664;
  assign N4663 = N4228 & en_i;
  assign N4664 = ~valid[108];
  assign match_array[109] = N4666 & valid[109];
  assign N4666 = N4665 & N3214;
  assign N4665 = N4228 & en_i;
  assign empty_array[109] = N4667 & N4668;
  assign N4667 = N4228 & en_i;
  assign N4668 = ~valid[109];
  assign match_array[110] = N4670 & valid[110];
  assign N4670 = N4669 & N3215;
  assign N4669 = N4228 & en_i;
  assign empty_array[110] = N4671 & N4672;
  assign N4671 = N4228 & en_i;
  assign N4672 = ~valid[110];
  assign match_array[111] = N4674 & valid[111];
  assign N4674 = N4673 & N3216;
  assign N4673 = N4228 & en_i;
  assign empty_array[111] = N4675 & N4676;
  assign N4675 = N4228 & en_i;
  assign N4676 = ~valid[111];
  assign match_array[112] = N4678 & valid[112];
  assign N4678 = N4677 & N3217;
  assign N4677 = N4228 & en_i;
  assign empty_array[112] = N4679 & N4680;
  assign N4679 = N4228 & en_i;
  assign N4680 = ~valid[112];
  assign match_array[113] = N4682 & valid[113];
  assign N4682 = N4681 & N3218;
  assign N4681 = N4228 & en_i;
  assign empty_array[113] = N4683 & N4684;
  assign N4683 = N4228 & en_i;
  assign N4684 = ~valid[113];
  assign match_array[114] = N4686 & valid[114];
  assign N4686 = N4685 & N3219;
  assign N4685 = N4228 & en_i;
  assign empty_array[114] = N4687 & N4688;
  assign N4687 = N4228 & en_i;
  assign N4688 = ~valid[114];
  assign match_array[115] = N4690 & valid[115];
  assign N4690 = N4689 & N3220;
  assign N4689 = N4228 & en_i;
  assign empty_array[115] = N4691 & N4692;
  assign N4691 = N4228 & en_i;
  assign N4692 = ~valid[115];
  assign match_array[116] = N4694 & valid[116];
  assign N4694 = N4693 & N3221;
  assign N4693 = N4228 & en_i;
  assign empty_array[116] = N4695 & N4696;
  assign N4695 = N4228 & en_i;
  assign N4696 = ~valid[116];
  assign match_array[117] = N4698 & valid[117];
  assign N4698 = N4697 & N3222;
  assign N4697 = N4228 & en_i;
  assign empty_array[117] = N4699 & N4700;
  assign N4699 = N4228 & en_i;
  assign N4700 = ~valid[117];
  assign match_array[118] = N4702 & valid[118];
  assign N4702 = N4701 & N3223;
  assign N4701 = N4228 & en_i;
  assign empty_array[118] = N4703 & N4704;
  assign N4703 = N4228 & en_i;
  assign N4704 = ~valid[118];
  assign match_array[119] = N4706 & valid[119];
  assign N4706 = N4705 & N3224;
  assign N4705 = N4228 & en_i;
  assign empty_array[119] = N4707 & N4708;
  assign N4707 = N4228 & en_i;
  assign N4708 = ~valid[119];
  assign match_array[120] = N4710 & valid[120];
  assign N4710 = N4709 & N3225;
  assign N4709 = N4228 & en_i;
  assign empty_array[120] = N4711 & N4712;
  assign N4711 = N4228 & en_i;
  assign N4712 = ~valid[120];
  assign match_array[121] = N4714 & valid[121];
  assign N4714 = N4713 & N3226;
  assign N4713 = N4228 & en_i;
  assign empty_array[121] = N4715 & N4716;
  assign N4715 = N4228 & en_i;
  assign N4716 = ~valid[121];
  assign match_array[122] = N4718 & valid[122];
  assign N4718 = N4717 & N3227;
  assign N4717 = N4228 & en_i;
  assign empty_array[122] = N4719 & N4720;
  assign N4719 = N4228 & en_i;
  assign N4720 = ~valid[122];
  assign match_array[123] = N4722 & valid[123];
  assign N4722 = N4721 & N3228;
  assign N4721 = N4228 & en_i;
  assign empty_array[123] = N4723 & N4724;
  assign N4723 = N4228 & en_i;
  assign N4724 = ~valid[123];
  assign match_array[124] = N4726 & valid[124];
  assign N4726 = N4725 & N3229;
  assign N4725 = N4228 & en_i;
  assign empty_array[124] = N4727 & N4728;
  assign N4727 = N4228 & en_i;
  assign N4728 = ~valid[124];
  assign match_array[125] = N4730 & valid[125];
  assign N4730 = N4729 & N3230;
  assign N4729 = N4228 & en_i;
  assign empty_array[125] = N4731 & N4732;
  assign N4731 = N4228 & en_i;
  assign N4732 = ~valid[125];
  assign match_array[126] = N4734 & valid[126];
  assign N4734 = N4733 & N3231;
  assign N4733 = N4228 & en_i;
  assign empty_array[126] = N4735 & N4736;
  assign N4735 = N4228 & en_i;
  assign N4736 = ~valid[126];
  assign match_array[127] = N4738 & valid[127];
  assign N4738 = N4737 & N3232;
  assign N4737 = N4228 & en_i;
  assign empty_array[127] = N4739 & N4740;
  assign N4739 = N4228 & en_i;
  assign N4740 = ~valid[127];
  assign match_array[128] = N4742 & valid[128];
  assign N4742 = N4741 & N3233;
  assign N4741 = N4228 & en_i;
  assign empty_array[128] = N4743 & N4744;
  assign N4743 = N4228 & en_i;
  assign N4744 = ~valid[128];
  assign match_array[129] = N4746 & valid[129];
  assign N4746 = N4745 & N3234;
  assign N4745 = N4228 & en_i;
  assign empty_array[129] = N4747 & N4748;
  assign N4747 = N4228 & en_i;
  assign N4748 = ~valid[129];
  assign match_array[130] = N4750 & valid[130];
  assign N4750 = N4749 & N3235;
  assign N4749 = N4228 & en_i;
  assign empty_array[130] = N4751 & N4752;
  assign N4751 = N4228 & en_i;
  assign N4752 = ~valid[130];
  assign match_array[131] = N4754 & valid[131];
  assign N4754 = N4753 & N3236;
  assign N4753 = N4228 & en_i;
  assign empty_array[131] = N4755 & N4756;
  assign N4755 = N4228 & en_i;
  assign N4756 = ~valid[131];
  assign match_array[132] = N4758 & valid[132];
  assign N4758 = N4757 & N3237;
  assign N4757 = N4228 & en_i;
  assign empty_array[132] = N4759 & N4760;
  assign N4759 = N4228 & en_i;
  assign N4760 = ~valid[132];
  assign match_array[133] = N4762 & valid[133];
  assign N4762 = N4761 & N3238;
  assign N4761 = N4228 & en_i;
  assign empty_array[133] = N4763 & N4764;
  assign N4763 = N4228 & en_i;
  assign N4764 = ~valid[133];
  assign match_array[134] = N4766 & valid[134];
  assign N4766 = N4765 & N3239;
  assign N4765 = N4228 & en_i;
  assign empty_array[134] = N4767 & N4768;
  assign N4767 = N4228 & en_i;
  assign N4768 = ~valid[134];
  assign match_array[135] = N4770 & valid[135];
  assign N4770 = N4769 & N3240;
  assign N4769 = N4228 & en_i;
  assign empty_array[135] = N4771 & N4772;
  assign N4771 = N4228 & en_i;
  assign N4772 = ~valid[135];
  assign match_array[136] = N4774 & valid[136];
  assign N4774 = N4773 & N3241;
  assign N4773 = N4228 & en_i;
  assign empty_array[136] = N4775 & N4776;
  assign N4775 = N4228 & en_i;
  assign N4776 = ~valid[136];
  assign match_array[137] = N4778 & valid[137];
  assign N4778 = N4777 & N3242;
  assign N4777 = N4228 & en_i;
  assign empty_array[137] = N4779 & N4780;
  assign N4779 = N4228 & en_i;
  assign N4780 = ~valid[137];
  assign match_array[138] = N4782 & valid[138];
  assign N4782 = N4781 & N3243;
  assign N4781 = N4228 & en_i;
  assign empty_array[138] = N4783 & N4784;
  assign N4783 = N4228 & en_i;
  assign N4784 = ~valid[138];
  assign match_array[139] = N4786 & valid[139];
  assign N4786 = N4785 & N3244;
  assign N4785 = N4228 & en_i;
  assign empty_array[139] = N4787 & N4788;
  assign N4787 = N4228 & en_i;
  assign N4788 = ~valid[139];
  assign match_array[140] = N4790 & valid[140];
  assign N4790 = N4789 & N3245;
  assign N4789 = N4228 & en_i;
  assign empty_array[140] = N4791 & N4792;
  assign N4791 = N4228 & en_i;
  assign N4792 = ~valid[140];
  assign match_array[141] = N4794 & valid[141];
  assign N4794 = N4793 & N3246;
  assign N4793 = N4228 & en_i;
  assign empty_array[141] = N4795 & N4796;
  assign N4795 = N4228 & en_i;
  assign N4796 = ~valid[141];
  assign match_array[142] = N4798 & valid[142];
  assign N4798 = N4797 & N3247;
  assign N4797 = N4228 & en_i;
  assign empty_array[142] = N4799 & N4800;
  assign N4799 = N4228 & en_i;
  assign N4800 = ~valid[142];
  assign match_array[143] = N4802 & valid[143];
  assign N4802 = N4801 & N3248;
  assign N4801 = N4228 & en_i;
  assign empty_array[143] = N4803 & N4804;
  assign N4803 = N4228 & en_i;
  assign N4804 = ~valid[143];
  assign match_array[144] = N4806 & valid[144];
  assign N4806 = N4805 & N3249;
  assign N4805 = N4228 & en_i;
  assign empty_array[144] = N4807 & N4808;
  assign N4807 = N4228 & en_i;
  assign N4808 = ~valid[144];
  assign match_array[145] = N4810 & valid[145];
  assign N4810 = N4809 & N3250;
  assign N4809 = N4228 & en_i;
  assign empty_array[145] = N4811 & N4812;
  assign N4811 = N4228 & en_i;
  assign N4812 = ~valid[145];
  assign match_array[146] = N4814 & valid[146];
  assign N4814 = N4813 & N3251;
  assign N4813 = N4228 & en_i;
  assign empty_array[146] = N4815 & N4816;
  assign N4815 = N4228 & en_i;
  assign N4816 = ~valid[146];
  assign match_array[147] = N4818 & valid[147];
  assign N4818 = N4817 & N3252;
  assign N4817 = N4228 & en_i;
  assign empty_array[147] = N4819 & N4820;
  assign N4819 = N4228 & en_i;
  assign N4820 = ~valid[147];
  assign match_array[148] = N4822 & valid[148];
  assign N4822 = N4821 & N3253;
  assign N4821 = N4228 & en_i;
  assign empty_array[148] = N4823 & N4824;
  assign N4823 = N4228 & en_i;
  assign N4824 = ~valid[148];
  assign match_array[149] = N4826 & valid[149];
  assign N4826 = N4825 & N3254;
  assign N4825 = N4228 & en_i;
  assign empty_array[149] = N4827 & N4828;
  assign N4827 = N4228 & en_i;
  assign N4828 = ~valid[149];
  assign match_array[150] = N4830 & valid[150];
  assign N4830 = N4829 & N3255;
  assign N4829 = N4228 & en_i;
  assign empty_array[150] = N4831 & N4832;
  assign N4831 = N4228 & en_i;
  assign N4832 = ~valid[150];
  assign match_array[151] = N4834 & valid[151];
  assign N4834 = N4833 & N3256;
  assign N4833 = N4228 & en_i;
  assign empty_array[151] = N4835 & N4836;
  assign N4835 = N4228 & en_i;
  assign N4836 = ~valid[151];
  assign match_array[152] = N4838 & valid[152];
  assign N4838 = N4837 & N3257;
  assign N4837 = N4228 & en_i;
  assign empty_array[152] = N4839 & N4840;
  assign N4839 = N4228 & en_i;
  assign N4840 = ~valid[152];
  assign match_array[153] = N4842 & valid[153];
  assign N4842 = N4841 & N3258;
  assign N4841 = N4228 & en_i;
  assign empty_array[153] = N4843 & N4844;
  assign N4843 = N4228 & en_i;
  assign N4844 = ~valid[153];
  assign match_array[154] = N4846 & valid[154];
  assign N4846 = N4845 & N3259;
  assign N4845 = N4228 & en_i;
  assign empty_array[154] = N4847 & N4848;
  assign N4847 = N4228 & en_i;
  assign N4848 = ~valid[154];
  assign match_array[155] = N4850 & valid[155];
  assign N4850 = N4849 & N3260;
  assign N4849 = N4228 & en_i;
  assign empty_array[155] = N4851 & N4852;
  assign N4851 = N4228 & en_i;
  assign N4852 = ~valid[155];
  assign match_array[156] = N4854 & valid[156];
  assign N4854 = N4853 & N3261;
  assign N4853 = N4228 & en_i;
  assign empty_array[156] = N4855 & N4856;
  assign N4855 = N4228 & en_i;
  assign N4856 = ~valid[156];
  assign match_array[157] = N4858 & valid[157];
  assign N4858 = N4857 & N3262;
  assign N4857 = N4228 & en_i;
  assign empty_array[157] = N4859 & N4860;
  assign N4859 = N4228 & en_i;
  assign N4860 = ~valid[157];
  assign match_array[158] = N4862 & valid[158];
  assign N4862 = N4861 & N3263;
  assign N4861 = N4228 & en_i;
  assign empty_array[158] = N4863 & N4864;
  assign N4863 = N4228 & en_i;
  assign N4864 = ~valid[158];
  assign match_array[159] = N4866 & valid[159];
  assign N4866 = N4865 & N3264;
  assign N4865 = N4228 & en_i;
  assign empty_array[159] = N4867 & N4868;
  assign N4867 = N4228 & en_i;
  assign N4868 = ~valid[159];
  assign match_array[160] = N4870 & valid[160];
  assign N4870 = N4869 & N3265;
  assign N4869 = N4228 & en_i;
  assign empty_array[160] = N4871 & N4872;
  assign N4871 = N4228 & en_i;
  assign N4872 = ~valid[160];
  assign match_array[161] = N4874 & valid[161];
  assign N4874 = N4873 & N3266;
  assign N4873 = N4228 & en_i;
  assign empty_array[161] = N4875 & N4876;
  assign N4875 = N4228 & en_i;
  assign N4876 = ~valid[161];
  assign match_array[162] = N4878 & valid[162];
  assign N4878 = N4877 & N3267;
  assign N4877 = N4228 & en_i;
  assign empty_array[162] = N4879 & N4880;
  assign N4879 = N4228 & en_i;
  assign N4880 = ~valid[162];
  assign match_array[163] = N4882 & valid[163];
  assign N4882 = N4881 & N3268;
  assign N4881 = N4228 & en_i;
  assign empty_array[163] = N4883 & N4884;
  assign N4883 = N4228 & en_i;
  assign N4884 = ~valid[163];
  assign match_array[164] = N4886 & valid[164];
  assign N4886 = N4885 & N3269;
  assign N4885 = N4228 & en_i;
  assign empty_array[164] = N4887 & N4888;
  assign N4887 = N4228 & en_i;
  assign N4888 = ~valid[164];
  assign match_array[165] = N4890 & valid[165];
  assign N4890 = N4889 & N3270;
  assign N4889 = N4228 & en_i;
  assign empty_array[165] = N4891 & N4892;
  assign N4891 = N4228 & en_i;
  assign N4892 = ~valid[165];
  assign match_array[166] = N4894 & valid[166];
  assign N4894 = N4893 & N3271;
  assign N4893 = N4228 & en_i;
  assign empty_array[166] = N4895 & N4896;
  assign N4895 = N4228 & en_i;
  assign N4896 = ~valid[166];
  assign match_array[167] = N4898 & valid[167];
  assign N4898 = N4897 & N3272;
  assign N4897 = N4228 & en_i;
  assign empty_array[167] = N4899 & N4900;
  assign N4899 = N4228 & en_i;
  assign N4900 = ~valid[167];
  assign match_array[168] = N4902 & valid[168];
  assign N4902 = N4901 & N3273;
  assign N4901 = N4228 & en_i;
  assign empty_array[168] = N4903 & N4904;
  assign N4903 = N4228 & en_i;
  assign N4904 = ~valid[168];
  assign match_array[169] = N4906 & valid[169];
  assign N4906 = N4905 & N3274;
  assign N4905 = N4228 & en_i;
  assign empty_array[169] = N4907 & N4908;
  assign N4907 = N4228 & en_i;
  assign N4908 = ~valid[169];
  assign match_array[170] = N4910 & valid[170];
  assign N4910 = N4909 & N3275;
  assign N4909 = N4228 & en_i;
  assign empty_array[170] = N4911 & N4912;
  assign N4911 = N4228 & en_i;
  assign N4912 = ~valid[170];
  assign match_array[171] = N4914 & valid[171];
  assign N4914 = N4913 & N3276;
  assign N4913 = N4228 & en_i;
  assign empty_array[171] = N4915 & N4916;
  assign N4915 = N4228 & en_i;
  assign N4916 = ~valid[171];
  assign match_array[172] = N4918 & valid[172];
  assign N4918 = N4917 & N3277;
  assign N4917 = N4228 & en_i;
  assign empty_array[172] = N4919 & N4920;
  assign N4919 = N4228 & en_i;
  assign N4920 = ~valid[172];
  assign match_array[173] = N4922 & valid[173];
  assign N4922 = N4921 & N3278;
  assign N4921 = N4228 & en_i;
  assign empty_array[173] = N4923 & N4924;
  assign N4923 = N4228 & en_i;
  assign N4924 = ~valid[173];
  assign match_array[174] = N4926 & valid[174];
  assign N4926 = N4925 & N3279;
  assign N4925 = N4228 & en_i;
  assign empty_array[174] = N4927 & N4928;
  assign N4927 = N4228 & en_i;
  assign N4928 = ~valid[174];
  assign match_array[175] = N4930 & valid[175];
  assign N4930 = N4929 & N3280;
  assign N4929 = N4228 & en_i;
  assign empty_array[175] = N4931 & N4932;
  assign N4931 = N4228 & en_i;
  assign N4932 = ~valid[175];
  assign match_array[176] = N4934 & valid[176];
  assign N4934 = N4933 & N3281;
  assign N4933 = N4228 & en_i;
  assign empty_array[176] = N4935 & N4936;
  assign N4935 = N4228 & en_i;
  assign N4936 = ~valid[176];
  assign match_array[177] = N4938 & valid[177];
  assign N4938 = N4937 & N3282;
  assign N4937 = N4228 & en_i;
  assign empty_array[177] = N4939 & N4940;
  assign N4939 = N4228 & en_i;
  assign N4940 = ~valid[177];
  assign match_array[178] = N4942 & valid[178];
  assign N4942 = N4941 & N3283;
  assign N4941 = N4228 & en_i;
  assign empty_array[178] = N4943 & N4944;
  assign N4943 = N4228 & en_i;
  assign N4944 = ~valid[178];
  assign match_array[179] = N4946 & valid[179];
  assign N4946 = N4945 & N3284;
  assign N4945 = N4228 & en_i;
  assign empty_array[179] = N4947 & N4948;
  assign N4947 = N4228 & en_i;
  assign N4948 = ~valid[179];
  assign match_array[180] = N4950 & valid[180];
  assign N4950 = N4949 & N3285;
  assign N4949 = N4228 & en_i;
  assign empty_array[180] = N4951 & N4952;
  assign N4951 = N4228 & en_i;
  assign N4952 = ~valid[180];
  assign match_array[181] = N4954 & valid[181];
  assign N4954 = N4953 & N3286;
  assign N4953 = N4228 & en_i;
  assign empty_array[181] = N4955 & N4956;
  assign N4955 = N4228 & en_i;
  assign N4956 = ~valid[181];
  assign match_array[182] = N4958 & valid[182];
  assign N4958 = N4957 & N3287;
  assign N4957 = N4228 & en_i;
  assign empty_array[182] = N4959 & N4960;
  assign N4959 = N4228 & en_i;
  assign N4960 = ~valid[182];
  assign match_array[183] = N4962 & valid[183];
  assign N4962 = N4961 & N3288;
  assign N4961 = N4228 & en_i;
  assign empty_array[183] = N4963 & N4964;
  assign N4963 = N4228 & en_i;
  assign N4964 = ~valid[183];
  assign match_array[184] = N4966 & valid[184];
  assign N4966 = N4965 & N3289;
  assign N4965 = N4228 & en_i;
  assign empty_array[184] = N4967 & N4968;
  assign N4967 = N4228 & en_i;
  assign N4968 = ~valid[184];
  assign match_array[185] = N4970 & valid[185];
  assign N4970 = N4969 & N3290;
  assign N4969 = N4228 & en_i;
  assign empty_array[185] = N4971 & N4972;
  assign N4971 = N4228 & en_i;
  assign N4972 = ~valid[185];
  assign match_array[186] = N4974 & valid[186];
  assign N4974 = N4973 & N3291;
  assign N4973 = N4228 & en_i;
  assign empty_array[186] = N4975 & N4976;
  assign N4975 = N4228 & en_i;
  assign N4976 = ~valid[186];
  assign match_array[187] = N4978 & valid[187];
  assign N4978 = N4977 & N3292;
  assign N4977 = N4228 & en_i;
  assign empty_array[187] = N4979 & N4980;
  assign N4979 = N4228 & en_i;
  assign N4980 = ~valid[187];
  assign match_array[188] = N4982 & valid[188];
  assign N4982 = N4981 & N3293;
  assign N4981 = N4228 & en_i;
  assign empty_array[188] = N4983 & N4984;
  assign N4983 = N4228 & en_i;
  assign N4984 = ~valid[188];
  assign match_array[189] = N4986 & valid[189];
  assign N4986 = N4985 & N3294;
  assign N4985 = N4228 & en_i;
  assign empty_array[189] = N4987 & N4988;
  assign N4987 = N4228 & en_i;
  assign N4988 = ~valid[189];
  assign match_array[190] = N4990 & valid[190];
  assign N4990 = N4989 & N3295;
  assign N4989 = N4228 & en_i;
  assign empty_array[190] = N4991 & N4992;
  assign N4991 = N4228 & en_i;
  assign N4992 = ~valid[190];
  assign match_array[191] = N4994 & valid[191];
  assign N4994 = N4993 & N3296;
  assign N4993 = N4228 & en_i;
  assign empty_array[191] = N4995 & N4996;
  assign N4995 = N4228 & en_i;
  assign N4996 = ~valid[191];
  assign match_array[192] = N4998 & valid[192];
  assign N4998 = N4997 & N3297;
  assign N4997 = N4228 & en_i;
  assign empty_array[192] = N4999 & N5000;
  assign N4999 = N4228 & en_i;
  assign N5000 = ~valid[192];
  assign match_array[193] = N5002 & valid[193];
  assign N5002 = N5001 & N3298;
  assign N5001 = N4228 & en_i;
  assign empty_array[193] = N5003 & N5004;
  assign N5003 = N4228 & en_i;
  assign N5004 = ~valid[193];
  assign match_array[194] = N5006 & valid[194];
  assign N5006 = N5005 & N3299;
  assign N5005 = N4228 & en_i;
  assign empty_array[194] = N5007 & N5008;
  assign N5007 = N4228 & en_i;
  assign N5008 = ~valid[194];
  assign match_array[195] = N5010 & valid[195];
  assign N5010 = N5009 & N3300;
  assign N5009 = N4228 & en_i;
  assign empty_array[195] = N5011 & N5012;
  assign N5011 = N4228 & en_i;
  assign N5012 = ~valid[195];
  assign match_array[196] = N5014 & valid[196];
  assign N5014 = N5013 & N3301;
  assign N5013 = N4228 & en_i;
  assign empty_array[196] = N5015 & N5016;
  assign N5015 = N4228 & en_i;
  assign N5016 = ~valid[196];
  assign match_array[197] = N5018 & valid[197];
  assign N5018 = N5017 & N3302;
  assign N5017 = N4228 & en_i;
  assign empty_array[197] = N5019 & N5020;
  assign N5019 = N4228 & en_i;
  assign N5020 = ~valid[197];
  assign match_array[198] = N5022 & valid[198];
  assign N5022 = N5021 & N3303;
  assign N5021 = N4228 & en_i;
  assign empty_array[198] = N5023 & N5024;
  assign N5023 = N4228 & en_i;
  assign N5024 = ~valid[198];
  assign match_array[199] = N5026 & valid[199];
  assign N5026 = N5025 & N3304;
  assign N5025 = N4228 & en_i;
  assign empty_array[199] = N5027 & N5028;
  assign N5027 = N4228 & en_i;
  assign N5028 = ~valid[199];
  assign match_array[200] = N5030 & valid[200];
  assign N5030 = N5029 & N3305;
  assign N5029 = N4228 & en_i;
  assign empty_array[200] = N5031 & N5032;
  assign N5031 = N4228 & en_i;
  assign N5032 = ~valid[200];
  assign match_array[201] = N5034 & valid[201];
  assign N5034 = N5033 & N3306;
  assign N5033 = N4228 & en_i;
  assign empty_array[201] = N5035 & N5036;
  assign N5035 = N4228 & en_i;
  assign N5036 = ~valid[201];
  assign match_array[202] = N5038 & valid[202];
  assign N5038 = N5037 & N3307;
  assign N5037 = N4228 & en_i;
  assign empty_array[202] = N5039 & N5040;
  assign N5039 = N4228 & en_i;
  assign N5040 = ~valid[202];
  assign match_array[203] = N5042 & valid[203];
  assign N5042 = N5041 & N3308;
  assign N5041 = N4228 & en_i;
  assign empty_array[203] = N5043 & N5044;
  assign N5043 = N4228 & en_i;
  assign N5044 = ~valid[203];
  assign match_array[204] = N5046 & valid[204];
  assign N5046 = N5045 & N3309;
  assign N5045 = N4228 & en_i;
  assign empty_array[204] = N5047 & N5048;
  assign N5047 = N4228 & en_i;
  assign N5048 = ~valid[204];
  assign match_array[205] = N5050 & valid[205];
  assign N5050 = N5049 & N3310;
  assign N5049 = N4228 & en_i;
  assign empty_array[205] = N5051 & N5052;
  assign N5051 = N4228 & en_i;
  assign N5052 = ~valid[205];
  assign match_array[206] = N5054 & valid[206];
  assign N5054 = N5053 & N3311;
  assign N5053 = N4228 & en_i;
  assign empty_array[206] = N5055 & N5056;
  assign N5055 = N4228 & en_i;
  assign N5056 = ~valid[206];
  assign match_array[207] = N5058 & valid[207];
  assign N5058 = N5057 & N3312;
  assign N5057 = N4228 & en_i;
  assign empty_array[207] = N5059 & N5060;
  assign N5059 = N4228 & en_i;
  assign N5060 = ~valid[207];
  assign match_array[208] = N5062 & valid[208];
  assign N5062 = N5061 & N3313;
  assign N5061 = N4228 & en_i;
  assign empty_array[208] = N5063 & N5064;
  assign N5063 = N4228 & en_i;
  assign N5064 = ~valid[208];
  assign match_array[209] = N5066 & valid[209];
  assign N5066 = N5065 & N3314;
  assign N5065 = N4228 & en_i;
  assign empty_array[209] = N5067 & N5068;
  assign N5067 = N4228 & en_i;
  assign N5068 = ~valid[209];
  assign match_array[210] = N5070 & valid[210];
  assign N5070 = N5069 & N3315;
  assign N5069 = N4228 & en_i;
  assign empty_array[210] = N5071 & N5072;
  assign N5071 = N4228 & en_i;
  assign N5072 = ~valid[210];
  assign match_array[211] = N5074 & valid[211];
  assign N5074 = N5073 & N3316;
  assign N5073 = N4228 & en_i;
  assign empty_array[211] = N5075 & N5076;
  assign N5075 = N4228 & en_i;
  assign N5076 = ~valid[211];
  assign match_array[212] = N5078 & valid[212];
  assign N5078 = N5077 & N3317;
  assign N5077 = N4228 & en_i;
  assign empty_array[212] = N5079 & N5080;
  assign N5079 = N4228 & en_i;
  assign N5080 = ~valid[212];
  assign match_array[213] = N5082 & valid[213];
  assign N5082 = N5081 & N3318;
  assign N5081 = N4228 & en_i;
  assign empty_array[213] = N5083 & N5084;
  assign N5083 = N4228 & en_i;
  assign N5084 = ~valid[213];
  assign match_array[214] = N5086 & valid[214];
  assign N5086 = N5085 & N3319;
  assign N5085 = N4228 & en_i;
  assign empty_array[214] = N5087 & N5088;
  assign N5087 = N4228 & en_i;
  assign N5088 = ~valid[214];
  assign match_array[215] = N5090 & valid[215];
  assign N5090 = N5089 & N3320;
  assign N5089 = N4228 & en_i;
  assign empty_array[215] = N5091 & N5092;
  assign N5091 = N4228 & en_i;
  assign N5092 = ~valid[215];
  assign match_array[216] = N5094 & valid[216];
  assign N5094 = N5093 & N3321;
  assign N5093 = N4228 & en_i;
  assign empty_array[216] = N5095 & N5096;
  assign N5095 = N4228 & en_i;
  assign N5096 = ~valid[216];
  assign match_array[217] = N5098 & valid[217];
  assign N5098 = N5097 & N3322;
  assign N5097 = N4228 & en_i;
  assign empty_array[217] = N5099 & N5100;
  assign N5099 = N4228 & en_i;
  assign N5100 = ~valid[217];
  assign match_array[218] = N5102 & valid[218];
  assign N5102 = N5101 & N3323;
  assign N5101 = N4228 & en_i;
  assign empty_array[218] = N5103 & N5104;
  assign N5103 = N4228 & en_i;
  assign N5104 = ~valid[218];
  assign match_array[219] = N5106 & valid[219];
  assign N5106 = N5105 & N3324;
  assign N5105 = N4228 & en_i;
  assign empty_array[219] = N5107 & N5108;
  assign N5107 = N4228 & en_i;
  assign N5108 = ~valid[219];
  assign match_array[220] = N5110 & valid[220];
  assign N5110 = N5109 & N3325;
  assign N5109 = N4228 & en_i;
  assign empty_array[220] = N5111 & N5112;
  assign N5111 = N4228 & en_i;
  assign N5112 = ~valid[220];
  assign match_array[221] = N5114 & valid[221];
  assign N5114 = N5113 & N3326;
  assign N5113 = N4228 & en_i;
  assign empty_array[221] = N5115 & N5116;
  assign N5115 = N4228 & en_i;
  assign N5116 = ~valid[221];
  assign match_array[222] = N5118 & valid[222];
  assign N5118 = N5117 & N3327;
  assign N5117 = N4228 & en_i;
  assign empty_array[222] = N5119 & N5120;
  assign N5119 = N4228 & en_i;
  assign N5120 = ~valid[222];
  assign match_array[223] = N5122 & valid[223];
  assign N5122 = N5121 & N3328;
  assign N5121 = N4228 & en_i;
  assign empty_array[223] = N5123 & N5124;
  assign N5123 = N4228 & en_i;
  assign N5124 = ~valid[223];
  assign match_array[224] = N5126 & valid[224];
  assign N5126 = N5125 & N3329;
  assign N5125 = N4228 & en_i;
  assign empty_array[224] = N5127 & N5128;
  assign N5127 = N4228 & en_i;
  assign N5128 = ~valid[224];
  assign match_array[225] = N5130 & valid[225];
  assign N5130 = N5129 & N3330;
  assign N5129 = N4228 & en_i;
  assign empty_array[225] = N5131 & N5132;
  assign N5131 = N4228 & en_i;
  assign N5132 = ~valid[225];
  assign match_array[226] = N5134 & valid[226];
  assign N5134 = N5133 & N3331;
  assign N5133 = N4228 & en_i;
  assign empty_array[226] = N5135 & N5136;
  assign N5135 = N4228 & en_i;
  assign N5136 = ~valid[226];
  assign match_array[227] = N5138 & valid[227];
  assign N5138 = N5137 & N3332;
  assign N5137 = N4228 & en_i;
  assign empty_array[227] = N5139 & N5140;
  assign N5139 = N4228 & en_i;
  assign N5140 = ~valid[227];
  assign match_array[228] = N5142 & valid[228];
  assign N5142 = N5141 & N3333;
  assign N5141 = N4228 & en_i;
  assign empty_array[228] = N5143 & N5144;
  assign N5143 = N4228 & en_i;
  assign N5144 = ~valid[228];
  assign match_array[229] = N5146 & valid[229];
  assign N5146 = N5145 & N3334;
  assign N5145 = N4228 & en_i;
  assign empty_array[229] = N5147 & N5148;
  assign N5147 = N4228 & en_i;
  assign N5148 = ~valid[229];
  assign match_array[230] = N5150 & valid[230];
  assign N5150 = N5149 & N3335;
  assign N5149 = N4228 & en_i;
  assign empty_array[230] = N5151 & N5152;
  assign N5151 = N4228 & en_i;
  assign N5152 = ~valid[230];
  assign match_array[231] = N5154 & valid[231];
  assign N5154 = N5153 & N3336;
  assign N5153 = N4228 & en_i;
  assign empty_array[231] = N5155 & N5156;
  assign N5155 = N4228 & en_i;
  assign N5156 = ~valid[231];
  assign match_array[232] = N5158 & valid[232];
  assign N5158 = N5157 & N3337;
  assign N5157 = N4228 & en_i;
  assign empty_array[232] = N5159 & N5160;
  assign N5159 = N4228 & en_i;
  assign N5160 = ~valid[232];
  assign match_array[233] = N5162 & valid[233];
  assign N5162 = N5161 & N3338;
  assign N5161 = N4228 & en_i;
  assign empty_array[233] = N5163 & N5164;
  assign N5163 = N4228 & en_i;
  assign N5164 = ~valid[233];
  assign match_array[234] = N5166 & valid[234];
  assign N5166 = N5165 & N3339;
  assign N5165 = N4228 & en_i;
  assign empty_array[234] = N5167 & N5168;
  assign N5167 = N4228 & en_i;
  assign N5168 = ~valid[234];
  assign match_array[235] = N5170 & valid[235];
  assign N5170 = N5169 & N3340;
  assign N5169 = N4228 & en_i;
  assign empty_array[235] = N5171 & N5172;
  assign N5171 = N4228 & en_i;
  assign N5172 = ~valid[235];
  assign match_array[236] = N5174 & valid[236];
  assign N5174 = N5173 & N3341;
  assign N5173 = N4228 & en_i;
  assign empty_array[236] = N5175 & N5176;
  assign N5175 = N4228 & en_i;
  assign N5176 = ~valid[236];
  assign match_array[237] = N5178 & valid[237];
  assign N5178 = N5177 & N3342;
  assign N5177 = N4228 & en_i;
  assign empty_array[237] = N5179 & N5180;
  assign N5179 = N4228 & en_i;
  assign N5180 = ~valid[237];
  assign match_array[238] = N5182 & valid[238];
  assign N5182 = N5181 & N3343;
  assign N5181 = N4228 & en_i;
  assign empty_array[238] = N5183 & N5184;
  assign N5183 = N4228 & en_i;
  assign N5184 = ~valid[238];
  assign match_array[239] = N5186 & valid[239];
  assign N5186 = N5185 & N3344;
  assign N5185 = N4228 & en_i;
  assign empty_array[239] = N5187 & N5188;
  assign N5187 = N4228 & en_i;
  assign N5188 = ~valid[239];
  assign match_array[240] = N5190 & valid[240];
  assign N5190 = N5189 & N3345;
  assign N5189 = N4228 & en_i;
  assign empty_array[240] = N5191 & N5192;
  assign N5191 = N4228 & en_i;
  assign N5192 = ~valid[240];
  assign match_array[241] = N5194 & valid[241];
  assign N5194 = N5193 & N3346;
  assign N5193 = N4228 & en_i;
  assign empty_array[241] = N5195 & N5196;
  assign N5195 = N4228 & en_i;
  assign N5196 = ~valid[241];
  assign match_array[242] = N5198 & valid[242];
  assign N5198 = N5197 & N3347;
  assign N5197 = N4228 & en_i;
  assign empty_array[242] = N5199 & N5200;
  assign N5199 = N4228 & en_i;
  assign N5200 = ~valid[242];
  assign match_array[243] = N5202 & valid[243];
  assign N5202 = N5201 & N3348;
  assign N5201 = N4228 & en_i;
  assign empty_array[243] = N5203 & N5204;
  assign N5203 = N4228 & en_i;
  assign N5204 = ~valid[243];
  assign match_array[244] = N5206 & valid[244];
  assign N5206 = N5205 & N3349;
  assign N5205 = N4228 & en_i;
  assign empty_array[244] = N5207 & N5208;
  assign N5207 = N4228 & en_i;
  assign N5208 = ~valid[244];
  assign match_array[245] = N5210 & valid[245];
  assign N5210 = N5209 & N3350;
  assign N5209 = N4228 & en_i;
  assign empty_array[245] = N5211 & N5212;
  assign N5211 = N4228 & en_i;
  assign N5212 = ~valid[245];
  assign match_array[246] = N5214 & valid[246];
  assign N5214 = N5213 & N3351;
  assign N5213 = N4228 & en_i;
  assign empty_array[246] = N5215 & N5216;
  assign N5215 = N4228 & en_i;
  assign N5216 = ~valid[246];
  assign match_array[247] = N5218 & valid[247];
  assign N5218 = N5217 & N3352;
  assign N5217 = N4228 & en_i;
  assign empty_array[247] = N5219 & N5220;
  assign N5219 = N4228 & en_i;
  assign N5220 = ~valid[247];
  assign match_array[248] = N5222 & valid[248];
  assign N5222 = N5221 & N3353;
  assign N5221 = N4228 & en_i;
  assign empty_array[248] = N5223 & N5224;
  assign N5223 = N4228 & en_i;
  assign N5224 = ~valid[248];
  assign match_array[249] = N5226 & valid[249];
  assign N5226 = N5225 & N3354;
  assign N5225 = N4228 & en_i;
  assign empty_array[249] = N5227 & N5228;
  assign N5227 = N4228 & en_i;
  assign N5228 = ~valid[249];
  assign match_array[250] = N5230 & valid[250];
  assign N5230 = N5229 & N3355;
  assign N5229 = N4228 & en_i;
  assign empty_array[250] = N5231 & N5232;
  assign N5231 = N4228 & en_i;
  assign N5232 = ~valid[250];
  assign match_array[251] = N5234 & valid[251];
  assign N5234 = N5233 & N3356;
  assign N5233 = N4228 & en_i;
  assign empty_array[251] = N5235 & N5236;
  assign N5235 = N4228 & en_i;
  assign N5236 = ~valid[251];
  assign match_array[252] = N5238 & valid[252];
  assign N5238 = N5237 & N3357;
  assign N5237 = N4228 & en_i;
  assign empty_array[252] = N5239 & N5240;
  assign N5239 = N4228 & en_i;
  assign N5240 = ~valid[252];
  assign match_array[253] = N5242 & valid[253];
  assign N5242 = N5241 & N3358;
  assign N5241 = N4228 & en_i;
  assign empty_array[253] = N5243 & N5244;
  assign N5243 = N4228 & en_i;
  assign N5244 = ~valid[253];
  assign match_array[254] = N5246 & valid[254];
  assign N5246 = N5245 & N3359;
  assign N5245 = N4228 & en_i;
  assign empty_array[254] = N5247 & N5248;
  assign N5247 = N4228 & en_i;
  assign N5248 = ~valid[254];
  assign match_array[255] = N5250 & valid[255];
  assign N5250 = N5249 & N3360;
  assign N5249 = N4228 & en_i;
  assign empty_array[255] = N5251 & N5252;
  assign N5251 = N4228 & en_i;
  assign N5252 = ~valid[255];
  assign match_array[256] = N5254 & valid[256];
  assign N5254 = N5253 & N3361;
  assign N5253 = N4228 & en_i;
  assign empty_array[256] = N5255 & N5256;
  assign N5255 = N4228 & en_i;
  assign N5256 = ~valid[256];
  assign match_array[257] = N5258 & valid[257];
  assign N5258 = N5257 & N3362;
  assign N5257 = N4228 & en_i;
  assign empty_array[257] = N5259 & N5260;
  assign N5259 = N4228 & en_i;
  assign N5260 = ~valid[257];
  assign match_array[258] = N5262 & valid[258];
  assign N5262 = N5261 & N3363;
  assign N5261 = N4228 & en_i;
  assign empty_array[258] = N5263 & N5264;
  assign N5263 = N4228 & en_i;
  assign N5264 = ~valid[258];
  assign match_array[259] = N5266 & valid[259];
  assign N5266 = N5265 & N3364;
  assign N5265 = N4228 & en_i;
  assign empty_array[259] = N5267 & N5268;
  assign N5267 = N4228 & en_i;
  assign N5268 = ~valid[259];
  assign match_array[260] = N5270 & valid[260];
  assign N5270 = N5269 & N3365;
  assign N5269 = N4228 & en_i;
  assign empty_array[260] = N5271 & N5272;
  assign N5271 = N4228 & en_i;
  assign N5272 = ~valid[260];
  assign match_array[261] = N5274 & valid[261];
  assign N5274 = N5273 & N3366;
  assign N5273 = N4228 & en_i;
  assign empty_array[261] = N5275 & N5276;
  assign N5275 = N4228 & en_i;
  assign N5276 = ~valid[261];
  assign match_array[262] = N5278 & valid[262];
  assign N5278 = N5277 & N3367;
  assign N5277 = N4228 & en_i;
  assign empty_array[262] = N5279 & N5280;
  assign N5279 = N4228 & en_i;
  assign N5280 = ~valid[262];
  assign match_array[263] = N5282 & valid[263];
  assign N5282 = N5281 & N3368;
  assign N5281 = N4228 & en_i;
  assign empty_array[263] = N5283 & N5284;
  assign N5283 = N4228 & en_i;
  assign N5284 = ~valid[263];
  assign match_array[264] = N5286 & valid[264];
  assign N5286 = N5285 & N3369;
  assign N5285 = N4228 & en_i;
  assign empty_array[264] = N5287 & N5288;
  assign N5287 = N4228 & en_i;
  assign N5288 = ~valid[264];
  assign match_array[265] = N5290 & valid[265];
  assign N5290 = N5289 & N3370;
  assign N5289 = N4228 & en_i;
  assign empty_array[265] = N5291 & N5292;
  assign N5291 = N4228 & en_i;
  assign N5292 = ~valid[265];
  assign match_array[266] = N5294 & valid[266];
  assign N5294 = N5293 & N3371;
  assign N5293 = N4228 & en_i;
  assign empty_array[266] = N5295 & N5296;
  assign N5295 = N4228 & en_i;
  assign N5296 = ~valid[266];
  assign match_array[267] = N5298 & valid[267];
  assign N5298 = N5297 & N3372;
  assign N5297 = N4228 & en_i;
  assign empty_array[267] = N5299 & N5300;
  assign N5299 = N4228 & en_i;
  assign N5300 = ~valid[267];
  assign match_array[268] = N5302 & valid[268];
  assign N5302 = N5301 & N3373;
  assign N5301 = N4228 & en_i;
  assign empty_array[268] = N5303 & N5304;
  assign N5303 = N4228 & en_i;
  assign N5304 = ~valid[268];
  assign match_array[269] = N5306 & valid[269];
  assign N5306 = N5305 & N3374;
  assign N5305 = N4228 & en_i;
  assign empty_array[269] = N5307 & N5308;
  assign N5307 = N4228 & en_i;
  assign N5308 = ~valid[269];
  assign match_array[270] = N5310 & valid[270];
  assign N5310 = N5309 & N3375;
  assign N5309 = N4228 & en_i;
  assign empty_array[270] = N5311 & N5312;
  assign N5311 = N4228 & en_i;
  assign N5312 = ~valid[270];
  assign match_array[271] = N5314 & valid[271];
  assign N5314 = N5313 & N3376;
  assign N5313 = N4228 & en_i;
  assign empty_array[271] = N5315 & N5316;
  assign N5315 = N4228 & en_i;
  assign N5316 = ~valid[271];
  assign match_array[272] = N5318 & valid[272];
  assign N5318 = N5317 & N3377;
  assign N5317 = N4228 & en_i;
  assign empty_array[272] = N5319 & N5320;
  assign N5319 = N4228 & en_i;
  assign N5320 = ~valid[272];
  assign match_array[273] = N5322 & valid[273];
  assign N5322 = N5321 & N3378;
  assign N5321 = N4228 & en_i;
  assign empty_array[273] = N5323 & N5324;
  assign N5323 = N4228 & en_i;
  assign N5324 = ~valid[273];
  assign match_array[274] = N5326 & valid[274];
  assign N5326 = N5325 & N3379;
  assign N5325 = N4228 & en_i;
  assign empty_array[274] = N5327 & N5328;
  assign N5327 = N4228 & en_i;
  assign N5328 = ~valid[274];
  assign match_array[275] = N5330 & valid[275];
  assign N5330 = N5329 & N3380;
  assign N5329 = N4228 & en_i;
  assign empty_array[275] = N5331 & N5332;
  assign N5331 = N4228 & en_i;
  assign N5332 = ~valid[275];
  assign match_array[276] = N5334 & valid[276];
  assign N5334 = N5333 & N3381;
  assign N5333 = N4228 & en_i;
  assign empty_array[276] = N5335 & N5336;
  assign N5335 = N4228 & en_i;
  assign N5336 = ~valid[276];
  assign match_array[277] = N5338 & valid[277];
  assign N5338 = N5337 & N3382;
  assign N5337 = N4228 & en_i;
  assign empty_array[277] = N5339 & N5340;
  assign N5339 = N4228 & en_i;
  assign N5340 = ~valid[277];
  assign match_array[278] = N5342 & valid[278];
  assign N5342 = N5341 & N3383;
  assign N5341 = N4228 & en_i;
  assign empty_array[278] = N5343 & N5344;
  assign N5343 = N4228 & en_i;
  assign N5344 = ~valid[278];
  assign match_array[279] = N5346 & valid[279];
  assign N5346 = N5345 & N3384;
  assign N5345 = N4228 & en_i;
  assign empty_array[279] = N5347 & N5348;
  assign N5347 = N4228 & en_i;
  assign N5348 = ~valid[279];
  assign match_array[280] = N5350 & valid[280];
  assign N5350 = N5349 & N3385;
  assign N5349 = N4228 & en_i;
  assign empty_array[280] = N5351 & N5352;
  assign N5351 = N4228 & en_i;
  assign N5352 = ~valid[280];
  assign match_array[281] = N5354 & valid[281];
  assign N5354 = N5353 & N3386;
  assign N5353 = N4228 & en_i;
  assign empty_array[281] = N5355 & N5356;
  assign N5355 = N4228 & en_i;
  assign N5356 = ~valid[281];
  assign match_array[282] = N5358 & valid[282];
  assign N5358 = N5357 & N3387;
  assign N5357 = N4228 & en_i;
  assign empty_array[282] = N5359 & N5360;
  assign N5359 = N4228 & en_i;
  assign N5360 = ~valid[282];
  assign match_array[283] = N5362 & valid[283];
  assign N5362 = N5361 & N3388;
  assign N5361 = N4228 & en_i;
  assign empty_array[283] = N5363 & N5364;
  assign N5363 = N4228 & en_i;
  assign N5364 = ~valid[283];
  assign match_array[284] = N5366 & valid[284];
  assign N5366 = N5365 & N3389;
  assign N5365 = N4228 & en_i;
  assign empty_array[284] = N5367 & N5368;
  assign N5367 = N4228 & en_i;
  assign N5368 = ~valid[284];
  assign match_array[285] = N5370 & valid[285];
  assign N5370 = N5369 & N3390;
  assign N5369 = N4228 & en_i;
  assign empty_array[285] = N5371 & N5372;
  assign N5371 = N4228 & en_i;
  assign N5372 = ~valid[285];
  assign match_array[286] = N5374 & valid[286];
  assign N5374 = N5373 & N3391;
  assign N5373 = N4228 & en_i;
  assign empty_array[286] = N5375 & N5376;
  assign N5375 = N4228 & en_i;
  assign N5376 = ~valid[286];
  assign match_array[287] = N5378 & valid[287];
  assign N5378 = N5377 & N3392;
  assign N5377 = N4228 & en_i;
  assign empty_array[287] = N5379 & N5380;
  assign N5379 = N4228 & en_i;
  assign N5380 = ~valid[287];
  assign match_array[288] = N5382 & valid[288];
  assign N5382 = N5381 & N3393;
  assign N5381 = N4228 & en_i;
  assign empty_array[288] = N5383 & N5384;
  assign N5383 = N4228 & en_i;
  assign N5384 = ~valid[288];
  assign match_array[289] = N5386 & valid[289];
  assign N5386 = N5385 & N3394;
  assign N5385 = N4228 & en_i;
  assign empty_array[289] = N5387 & N5388;
  assign N5387 = N4228 & en_i;
  assign N5388 = ~valid[289];
  assign match_array[290] = N5390 & valid[290];
  assign N5390 = N5389 & N3395;
  assign N5389 = N4228 & en_i;
  assign empty_array[290] = N5391 & N5392;
  assign N5391 = N4228 & en_i;
  assign N5392 = ~valid[290];
  assign match_array[291] = N5394 & valid[291];
  assign N5394 = N5393 & N3396;
  assign N5393 = N4228 & en_i;
  assign empty_array[291] = N5395 & N5396;
  assign N5395 = N4228 & en_i;
  assign N5396 = ~valid[291];
  assign match_array[292] = N5398 & valid[292];
  assign N5398 = N5397 & N3397;
  assign N5397 = N4228 & en_i;
  assign empty_array[292] = N5399 & N5400;
  assign N5399 = N4228 & en_i;
  assign N5400 = ~valid[292];
  assign match_array[293] = N5402 & valid[293];
  assign N5402 = N5401 & N3398;
  assign N5401 = N4228 & en_i;
  assign empty_array[293] = N5403 & N5404;
  assign N5403 = N4228 & en_i;
  assign N5404 = ~valid[293];
  assign match_array[294] = N5406 & valid[294];
  assign N5406 = N5405 & N3399;
  assign N5405 = N4228 & en_i;
  assign empty_array[294] = N5407 & N5408;
  assign N5407 = N4228 & en_i;
  assign N5408 = ~valid[294];
  assign match_array[295] = N5410 & valid[295];
  assign N5410 = N5409 & N3400;
  assign N5409 = N4228 & en_i;
  assign empty_array[295] = N5411 & N5412;
  assign N5411 = N4228 & en_i;
  assign N5412 = ~valid[295];
  assign match_array[296] = N5414 & valid[296];
  assign N5414 = N5413 & N3401;
  assign N5413 = N4228 & en_i;
  assign empty_array[296] = N5415 & N5416;
  assign N5415 = N4228 & en_i;
  assign N5416 = ~valid[296];
  assign match_array[297] = N5418 & valid[297];
  assign N5418 = N5417 & N3402;
  assign N5417 = N4228 & en_i;
  assign empty_array[297] = N5419 & N5420;
  assign N5419 = N4228 & en_i;
  assign N5420 = ~valid[297];
  assign match_array[298] = N5422 & valid[298];
  assign N5422 = N5421 & N3403;
  assign N5421 = N4228 & en_i;
  assign empty_array[298] = N5423 & N5424;
  assign N5423 = N4228 & en_i;
  assign N5424 = ~valid[298];
  assign match_array[299] = N5426 & valid[299];
  assign N5426 = N5425 & N3404;
  assign N5425 = N4228 & en_i;
  assign empty_array[299] = N5427 & N5428;
  assign N5427 = N4228 & en_i;
  assign N5428 = ~valid[299];
  assign match_array[300] = N5430 & valid[300];
  assign N5430 = N5429 & N3405;
  assign N5429 = N4228 & en_i;
  assign empty_array[300] = N5431 & N5432;
  assign N5431 = N4228 & en_i;
  assign N5432 = ~valid[300];
  assign match_array[301] = N5434 & valid[301];
  assign N5434 = N5433 & N3406;
  assign N5433 = N4228 & en_i;
  assign empty_array[301] = N5435 & N5436;
  assign N5435 = N4228 & en_i;
  assign N5436 = ~valid[301];
  assign match_array[302] = N5438 & valid[302];
  assign N5438 = N5437 & N3407;
  assign N5437 = N4228 & en_i;
  assign empty_array[302] = N5439 & N5440;
  assign N5439 = N4228 & en_i;
  assign N5440 = ~valid[302];
  assign match_array[303] = N5442 & valid[303];
  assign N5442 = N5441 & N3408;
  assign N5441 = N4228 & en_i;
  assign empty_array[303] = N5443 & N5444;
  assign N5443 = N4228 & en_i;
  assign N5444 = ~valid[303];
  assign match_array[304] = N5446 & valid[304];
  assign N5446 = N5445 & N3409;
  assign N5445 = N4228 & en_i;
  assign empty_array[304] = N5447 & N5448;
  assign N5447 = N4228 & en_i;
  assign N5448 = ~valid[304];
  assign match_array[305] = N5450 & valid[305];
  assign N5450 = N5449 & N3410;
  assign N5449 = N4228 & en_i;
  assign empty_array[305] = N5451 & N5452;
  assign N5451 = N4228 & en_i;
  assign N5452 = ~valid[305];
  assign match_array[306] = N5454 & valid[306];
  assign N5454 = N5453 & N3411;
  assign N5453 = N4228 & en_i;
  assign empty_array[306] = N5455 & N5456;
  assign N5455 = N4228 & en_i;
  assign N5456 = ~valid[306];
  assign match_array[307] = N5458 & valid[307];
  assign N5458 = N5457 & N3412;
  assign N5457 = N4228 & en_i;
  assign empty_array[307] = N5459 & N5460;
  assign N5459 = N4228 & en_i;
  assign N5460 = ~valid[307];
  assign match_array[308] = N5462 & valid[308];
  assign N5462 = N5461 & N3413;
  assign N5461 = N4228 & en_i;
  assign empty_array[308] = N5463 & N5464;
  assign N5463 = N4228 & en_i;
  assign N5464 = ~valid[308];
  assign match_array[309] = N5466 & valid[309];
  assign N5466 = N5465 & N3414;
  assign N5465 = N4228 & en_i;
  assign empty_array[309] = N5467 & N5468;
  assign N5467 = N4228 & en_i;
  assign N5468 = ~valid[309];
  assign match_array[310] = N5470 & valid[310];
  assign N5470 = N5469 & N3415;
  assign N5469 = N4228 & en_i;
  assign empty_array[310] = N5471 & N5472;
  assign N5471 = N4228 & en_i;
  assign N5472 = ~valid[310];
  assign match_array[311] = N5474 & valid[311];
  assign N5474 = N5473 & N3416;
  assign N5473 = N4228 & en_i;
  assign empty_array[311] = N5475 & N5476;
  assign N5475 = N4228 & en_i;
  assign N5476 = ~valid[311];
  assign match_array[312] = N5478 & valid[312];
  assign N5478 = N5477 & N3417;
  assign N5477 = N4228 & en_i;
  assign empty_array[312] = N5479 & N5480;
  assign N5479 = N4228 & en_i;
  assign N5480 = ~valid[312];
  assign match_array[313] = N5482 & valid[313];
  assign N5482 = N5481 & N3418;
  assign N5481 = N4228 & en_i;
  assign empty_array[313] = N5483 & N5484;
  assign N5483 = N4228 & en_i;
  assign N5484 = ~valid[313];
  assign match_array[314] = N5486 & valid[314];
  assign N5486 = N5485 & N3419;
  assign N5485 = N4228 & en_i;
  assign empty_array[314] = N5487 & N5488;
  assign N5487 = N4228 & en_i;
  assign N5488 = ~valid[314];
  assign match_array[315] = N5490 & valid[315];
  assign N5490 = N5489 & N3420;
  assign N5489 = N4228 & en_i;
  assign empty_array[315] = N5491 & N5492;
  assign N5491 = N4228 & en_i;
  assign N5492 = ~valid[315];
  assign match_array[316] = N5494 & valid[316];
  assign N5494 = N5493 & N3421;
  assign N5493 = N4228 & en_i;
  assign empty_array[316] = N5495 & N5496;
  assign N5495 = N4228 & en_i;
  assign N5496 = ~valid[316];
  assign match_array[317] = N5498 & valid[317];
  assign N5498 = N5497 & N3422;
  assign N5497 = N4228 & en_i;
  assign empty_array[317] = N5499 & N5500;
  assign N5499 = N4228 & en_i;
  assign N5500 = ~valid[317];
  assign match_array[318] = N5502 & valid[318];
  assign N5502 = N5501 & N3423;
  assign N5501 = N4228 & en_i;
  assign empty_array[318] = N5503 & N5504;
  assign N5503 = N4228 & en_i;
  assign N5504 = ~valid[318];
  assign match_array[319] = N5506 & valid[319];
  assign N5506 = N5505 & N3424;
  assign N5505 = N4228 & en_i;
  assign empty_array[319] = N5507 & N5508;
  assign N5507 = N4228 & en_i;
  assign N5508 = ~valid[319];
  assign match_array[320] = N5510 & valid[320];
  assign N5510 = N5509 & N3425;
  assign N5509 = N4228 & en_i;
  assign empty_array[320] = N5511 & N5512;
  assign N5511 = N4228 & en_i;
  assign N5512 = ~valid[320];
  assign match_array[321] = N5514 & valid[321];
  assign N5514 = N5513 & N3426;
  assign N5513 = N4228 & en_i;
  assign empty_array[321] = N5515 & N5516;
  assign N5515 = N4228 & en_i;
  assign N5516 = ~valid[321];
  assign match_array[322] = N5518 & valid[322];
  assign N5518 = N5517 & N3427;
  assign N5517 = N4228 & en_i;
  assign empty_array[322] = N5519 & N5520;
  assign N5519 = N4228 & en_i;
  assign N5520 = ~valid[322];
  assign match_array[323] = N5522 & valid[323];
  assign N5522 = N5521 & N3428;
  assign N5521 = N4228 & en_i;
  assign empty_array[323] = N5523 & N5524;
  assign N5523 = N4228 & en_i;
  assign N5524 = ~valid[323];
  assign match_array[324] = N5526 & valid[324];
  assign N5526 = N5525 & N3429;
  assign N5525 = N4228 & en_i;
  assign empty_array[324] = N5527 & N5528;
  assign N5527 = N4228 & en_i;
  assign N5528 = ~valid[324];
  assign match_array[325] = N5530 & valid[325];
  assign N5530 = N5529 & N3430;
  assign N5529 = N4228 & en_i;
  assign empty_array[325] = N5531 & N5532;
  assign N5531 = N4228 & en_i;
  assign N5532 = ~valid[325];
  assign match_array[326] = N5534 & valid[326];
  assign N5534 = N5533 & N3431;
  assign N5533 = N4228 & en_i;
  assign empty_array[326] = N5535 & N5536;
  assign N5535 = N4228 & en_i;
  assign N5536 = ~valid[326];
  assign match_array[327] = N5538 & valid[327];
  assign N5538 = N5537 & N3432;
  assign N5537 = N4228 & en_i;
  assign empty_array[327] = N5539 & N5540;
  assign N5539 = N4228 & en_i;
  assign N5540 = ~valid[327];
  assign match_array[328] = N5542 & valid[328];
  assign N5542 = N5541 & N3433;
  assign N5541 = N4228 & en_i;
  assign empty_array[328] = N5543 & N5544;
  assign N5543 = N4228 & en_i;
  assign N5544 = ~valid[328];
  assign match_array[329] = N5546 & valid[329];
  assign N5546 = N5545 & N3434;
  assign N5545 = N4228 & en_i;
  assign empty_array[329] = N5547 & N5548;
  assign N5547 = N4228 & en_i;
  assign N5548 = ~valid[329];
  assign match_array[330] = N5550 & valid[330];
  assign N5550 = N5549 & N3435;
  assign N5549 = N4228 & en_i;
  assign empty_array[330] = N5551 & N5552;
  assign N5551 = N4228 & en_i;
  assign N5552 = ~valid[330];
  assign match_array[331] = N5554 & valid[331];
  assign N5554 = N5553 & N3436;
  assign N5553 = N4228 & en_i;
  assign empty_array[331] = N5555 & N5556;
  assign N5555 = N4228 & en_i;
  assign N5556 = ~valid[331];
  assign match_array[332] = N5558 & valid[332];
  assign N5558 = N5557 & N3437;
  assign N5557 = N4228 & en_i;
  assign empty_array[332] = N5559 & N5560;
  assign N5559 = N4228 & en_i;
  assign N5560 = ~valid[332];
  assign match_array[333] = N5562 & valid[333];
  assign N5562 = N5561 & N3438;
  assign N5561 = N4228 & en_i;
  assign empty_array[333] = N5563 & N5564;
  assign N5563 = N4228 & en_i;
  assign N5564 = ~valid[333];
  assign match_array[334] = N5566 & valid[334];
  assign N5566 = N5565 & N3439;
  assign N5565 = N4228 & en_i;
  assign empty_array[334] = N5567 & N5568;
  assign N5567 = N4228 & en_i;
  assign N5568 = ~valid[334];
  assign match_array[335] = N5570 & valid[335];
  assign N5570 = N5569 & N3440;
  assign N5569 = N4228 & en_i;
  assign empty_array[335] = N5571 & N5572;
  assign N5571 = N4228 & en_i;
  assign N5572 = ~valid[335];
  assign match_array[336] = N5574 & valid[336];
  assign N5574 = N5573 & N3441;
  assign N5573 = N4228 & en_i;
  assign empty_array[336] = N5575 & N5576;
  assign N5575 = N4228 & en_i;
  assign N5576 = ~valid[336];
  assign match_array[337] = N5578 & valid[337];
  assign N5578 = N5577 & N3442;
  assign N5577 = N4228 & en_i;
  assign empty_array[337] = N5579 & N5580;
  assign N5579 = N4228 & en_i;
  assign N5580 = ~valid[337];
  assign match_array[338] = N5582 & valid[338];
  assign N5582 = N5581 & N3443;
  assign N5581 = N4228 & en_i;
  assign empty_array[338] = N5583 & N5584;
  assign N5583 = N4228 & en_i;
  assign N5584 = ~valid[338];
  assign match_array[339] = N5586 & valid[339];
  assign N5586 = N5585 & N3444;
  assign N5585 = N4228 & en_i;
  assign empty_array[339] = N5587 & N5588;
  assign N5587 = N4228 & en_i;
  assign N5588 = ~valid[339];
  assign match_array[340] = N5590 & valid[340];
  assign N5590 = N5589 & N3445;
  assign N5589 = N4228 & en_i;
  assign empty_array[340] = N5591 & N5592;
  assign N5591 = N4228 & en_i;
  assign N5592 = ~valid[340];
  assign match_array[341] = N5594 & valid[341];
  assign N5594 = N5593 & N3446;
  assign N5593 = N4228 & en_i;
  assign empty_array[341] = N5595 & N5596;
  assign N5595 = N4228 & en_i;
  assign N5596 = ~valid[341];
  assign match_array[342] = N5598 & valid[342];
  assign N5598 = N5597 & N3447;
  assign N5597 = N4228 & en_i;
  assign empty_array[342] = N5599 & N5600;
  assign N5599 = N4228 & en_i;
  assign N5600 = ~valid[342];
  assign match_array[343] = N5602 & valid[343];
  assign N5602 = N5601 & N3448;
  assign N5601 = N4228 & en_i;
  assign empty_array[343] = N5603 & N5604;
  assign N5603 = N4228 & en_i;
  assign N5604 = ~valid[343];
  assign match_array[344] = N5606 & valid[344];
  assign N5606 = N5605 & N3449;
  assign N5605 = N4228 & en_i;
  assign empty_array[344] = N5607 & N5608;
  assign N5607 = N4228 & en_i;
  assign N5608 = ~valid[344];
  assign match_array[345] = N5610 & valid[345];
  assign N5610 = N5609 & N3450;
  assign N5609 = N4228 & en_i;
  assign empty_array[345] = N5611 & N5612;
  assign N5611 = N4228 & en_i;
  assign N5612 = ~valid[345];
  assign match_array[346] = N5614 & valid[346];
  assign N5614 = N5613 & N3451;
  assign N5613 = N4228 & en_i;
  assign empty_array[346] = N5615 & N5616;
  assign N5615 = N4228 & en_i;
  assign N5616 = ~valid[346];
  assign match_array[347] = N5618 & valid[347];
  assign N5618 = N5617 & N3452;
  assign N5617 = N4228 & en_i;
  assign empty_array[347] = N5619 & N5620;
  assign N5619 = N4228 & en_i;
  assign N5620 = ~valid[347];
  assign match_array[348] = N5622 & valid[348];
  assign N5622 = N5621 & N3453;
  assign N5621 = N4228 & en_i;
  assign empty_array[348] = N5623 & N5624;
  assign N5623 = N4228 & en_i;
  assign N5624 = ~valid[348];
  assign match_array[349] = N5626 & valid[349];
  assign N5626 = N5625 & N3454;
  assign N5625 = N4228 & en_i;
  assign empty_array[349] = N5627 & N5628;
  assign N5627 = N4228 & en_i;
  assign N5628 = ~valid[349];
  assign match_array[350] = N5630 & valid[350];
  assign N5630 = N5629 & N3455;
  assign N5629 = N4228 & en_i;
  assign empty_array[350] = N5631 & N5632;
  assign N5631 = N4228 & en_i;
  assign N5632 = ~valid[350];
  assign match_array[351] = N5634 & valid[351];
  assign N5634 = N5633 & N3456;
  assign N5633 = N4228 & en_i;
  assign empty_array[351] = N5635 & N5636;
  assign N5635 = N4228 & en_i;
  assign N5636 = ~valid[351];
  assign match_array[352] = N5638 & valid[352];
  assign N5638 = N5637 & N3457;
  assign N5637 = N4228 & en_i;
  assign empty_array[352] = N5639 & N5640;
  assign N5639 = N4228 & en_i;
  assign N5640 = ~valid[352];
  assign match_array[353] = N5642 & valid[353];
  assign N5642 = N5641 & N3458;
  assign N5641 = N4228 & en_i;
  assign empty_array[353] = N5643 & N5644;
  assign N5643 = N4228 & en_i;
  assign N5644 = ~valid[353];
  assign match_array[354] = N5646 & valid[354];
  assign N5646 = N5645 & N3459;
  assign N5645 = N4228 & en_i;
  assign empty_array[354] = N5647 & N5648;
  assign N5647 = N4228 & en_i;
  assign N5648 = ~valid[354];
  assign match_array[355] = N5650 & valid[355];
  assign N5650 = N5649 & N3460;
  assign N5649 = N4228 & en_i;
  assign empty_array[355] = N5651 & N5652;
  assign N5651 = N4228 & en_i;
  assign N5652 = ~valid[355];
  assign match_array[356] = N5654 & valid[356];
  assign N5654 = N5653 & N3461;
  assign N5653 = N4228 & en_i;
  assign empty_array[356] = N5655 & N5656;
  assign N5655 = N4228 & en_i;
  assign N5656 = ~valid[356];
  assign match_array[357] = N5658 & valid[357];
  assign N5658 = N5657 & N3462;
  assign N5657 = N4228 & en_i;
  assign empty_array[357] = N5659 & N5660;
  assign N5659 = N4228 & en_i;
  assign N5660 = ~valid[357];
  assign match_array[358] = N5662 & valid[358];
  assign N5662 = N5661 & N3463;
  assign N5661 = N4228 & en_i;
  assign empty_array[358] = N5663 & N5664;
  assign N5663 = N4228 & en_i;
  assign N5664 = ~valid[358];
  assign match_array[359] = N5666 & valid[359];
  assign N5666 = N5665 & N3464;
  assign N5665 = N4228 & en_i;
  assign empty_array[359] = N5667 & N5668;
  assign N5667 = N4228 & en_i;
  assign N5668 = ~valid[359];
  assign match_array[360] = N5670 & valid[360];
  assign N5670 = N5669 & N3465;
  assign N5669 = N4228 & en_i;
  assign empty_array[360] = N5671 & N5672;
  assign N5671 = N4228 & en_i;
  assign N5672 = ~valid[360];
  assign match_array[361] = N5674 & valid[361];
  assign N5674 = N5673 & N3466;
  assign N5673 = N4228 & en_i;
  assign empty_array[361] = N5675 & N5676;
  assign N5675 = N4228 & en_i;
  assign N5676 = ~valid[361];
  assign match_array[362] = N5678 & valid[362];
  assign N5678 = N5677 & N3467;
  assign N5677 = N4228 & en_i;
  assign empty_array[362] = N5679 & N5680;
  assign N5679 = N4228 & en_i;
  assign N5680 = ~valid[362];
  assign match_array[363] = N5682 & valid[363];
  assign N5682 = N5681 & N3468;
  assign N5681 = N4228 & en_i;
  assign empty_array[363] = N5683 & N5684;
  assign N5683 = N4228 & en_i;
  assign N5684 = ~valid[363];
  assign match_array[364] = N5686 & valid[364];
  assign N5686 = N5685 & N3469;
  assign N5685 = N4228 & en_i;
  assign empty_array[364] = N5687 & N5688;
  assign N5687 = N4228 & en_i;
  assign N5688 = ~valid[364];
  assign match_array[365] = N5690 & valid[365];
  assign N5690 = N5689 & N3470;
  assign N5689 = N4228 & en_i;
  assign empty_array[365] = N5691 & N5692;
  assign N5691 = N4228 & en_i;
  assign N5692 = ~valid[365];
  assign match_array[366] = N5694 & valid[366];
  assign N5694 = N5693 & N3471;
  assign N5693 = N4228 & en_i;
  assign empty_array[366] = N5695 & N5696;
  assign N5695 = N4228 & en_i;
  assign N5696 = ~valid[366];
  assign match_array[367] = N5698 & valid[367];
  assign N5698 = N5697 & N3472;
  assign N5697 = N4228 & en_i;
  assign empty_array[367] = N5699 & N5700;
  assign N5699 = N4228 & en_i;
  assign N5700 = ~valid[367];
  assign match_array[368] = N5702 & valid[368];
  assign N5702 = N5701 & N3473;
  assign N5701 = N4228 & en_i;
  assign empty_array[368] = N5703 & N5704;
  assign N5703 = N4228 & en_i;
  assign N5704 = ~valid[368];
  assign match_array[369] = N5706 & valid[369];
  assign N5706 = N5705 & N3474;
  assign N5705 = N4228 & en_i;
  assign empty_array[369] = N5707 & N5708;
  assign N5707 = N4228 & en_i;
  assign N5708 = ~valid[369];
  assign match_array[370] = N5710 & valid[370];
  assign N5710 = N5709 & N3475;
  assign N5709 = N4228 & en_i;
  assign empty_array[370] = N5711 & N5712;
  assign N5711 = N4228 & en_i;
  assign N5712 = ~valid[370];
  assign match_array[371] = N5714 & valid[371];
  assign N5714 = N5713 & N3476;
  assign N5713 = N4228 & en_i;
  assign empty_array[371] = N5715 & N5716;
  assign N5715 = N4228 & en_i;
  assign N5716 = ~valid[371];
  assign match_array[372] = N5718 & valid[372];
  assign N5718 = N5717 & N3477;
  assign N5717 = N4228 & en_i;
  assign empty_array[372] = N5719 & N5720;
  assign N5719 = N4228 & en_i;
  assign N5720 = ~valid[372];
  assign match_array[373] = N5722 & valid[373];
  assign N5722 = N5721 & N3478;
  assign N5721 = N4228 & en_i;
  assign empty_array[373] = N5723 & N5724;
  assign N5723 = N4228 & en_i;
  assign N5724 = ~valid[373];
  assign match_array[374] = N5726 & valid[374];
  assign N5726 = N5725 & N3479;
  assign N5725 = N4228 & en_i;
  assign empty_array[374] = N5727 & N5728;
  assign N5727 = N4228 & en_i;
  assign N5728 = ~valid[374];
  assign match_array[375] = N5730 & valid[375];
  assign N5730 = N5729 & N3480;
  assign N5729 = N4228 & en_i;
  assign empty_array[375] = N5731 & N5732;
  assign N5731 = N4228 & en_i;
  assign N5732 = ~valid[375];
  assign match_array[376] = N5734 & valid[376];
  assign N5734 = N5733 & N3481;
  assign N5733 = N4228 & en_i;
  assign empty_array[376] = N5735 & N5736;
  assign N5735 = N4228 & en_i;
  assign N5736 = ~valid[376];
  assign match_array[377] = N5738 & valid[377];
  assign N5738 = N5737 & N3482;
  assign N5737 = N4228 & en_i;
  assign empty_array[377] = N5739 & N5740;
  assign N5739 = N4228 & en_i;
  assign N5740 = ~valid[377];
  assign match_array[378] = N5742 & valid[378];
  assign N5742 = N5741 & N3483;
  assign N5741 = N4228 & en_i;
  assign empty_array[378] = N5743 & N5744;
  assign N5743 = N4228 & en_i;
  assign N5744 = ~valid[378];
  assign match_array[379] = N5746 & valid[379];
  assign N5746 = N5745 & N3484;
  assign N5745 = N4228 & en_i;
  assign empty_array[379] = N5747 & N5748;
  assign N5747 = N4228 & en_i;
  assign N5748 = ~valid[379];
  assign match_array[380] = N5750 & valid[380];
  assign N5750 = N5749 & N3485;
  assign N5749 = N4228 & en_i;
  assign empty_array[380] = N5751 & N5752;
  assign N5751 = N4228 & en_i;
  assign N5752 = ~valid[380];
  assign match_array[381] = N5754 & valid[381];
  assign N5754 = N5753 & N3486;
  assign N5753 = N4228 & en_i;
  assign empty_array[381] = N5755 & N5756;
  assign N5755 = N4228 & en_i;
  assign N5756 = ~valid[381];
  assign match_array[382] = N5758 & valid[382];
  assign N5758 = N5757 & N3487;
  assign N5757 = N4228 & en_i;
  assign empty_array[382] = N5759 & N5760;
  assign N5759 = N4228 & en_i;
  assign N5760 = ~valid[382];
  assign match_array[383] = N5762 & valid[383];
  assign N5762 = N5761 & N3488;
  assign N5761 = N4228 & en_i;
  assign empty_array[383] = N5763 & N5764;
  assign N5763 = N4228 & en_i;
  assign N5764 = ~valid[383];
  assign match_array[384] = N5766 & valid[384];
  assign N5766 = N5765 & N3489;
  assign N5765 = N4228 & en_i;
  assign empty_array[384] = N5767 & N5768;
  assign N5767 = N4228 & en_i;
  assign N5768 = ~valid[384];
  assign match_array[385] = N5770 & valid[385];
  assign N5770 = N5769 & N3490;
  assign N5769 = N4228 & en_i;
  assign empty_array[385] = N5771 & N5772;
  assign N5771 = N4228 & en_i;
  assign N5772 = ~valid[385];
  assign match_array[386] = N5774 & valid[386];
  assign N5774 = N5773 & N3491;
  assign N5773 = N4228 & en_i;
  assign empty_array[386] = N5775 & N5776;
  assign N5775 = N4228 & en_i;
  assign N5776 = ~valid[386];
  assign match_array[387] = N5778 & valid[387];
  assign N5778 = N5777 & N3492;
  assign N5777 = N4228 & en_i;
  assign empty_array[387] = N5779 & N5780;
  assign N5779 = N4228 & en_i;
  assign N5780 = ~valid[387];
  assign match_array[388] = N5782 & valid[388];
  assign N5782 = N5781 & N3493;
  assign N5781 = N4228 & en_i;
  assign empty_array[388] = N5783 & N5784;
  assign N5783 = N4228 & en_i;
  assign N5784 = ~valid[388];
  assign match_array[389] = N5786 & valid[389];
  assign N5786 = N5785 & N3494;
  assign N5785 = N4228 & en_i;
  assign empty_array[389] = N5787 & N5788;
  assign N5787 = N4228 & en_i;
  assign N5788 = ~valid[389];
  assign match_array[390] = N5790 & valid[390];
  assign N5790 = N5789 & N3495;
  assign N5789 = N4228 & en_i;
  assign empty_array[390] = N5791 & N5792;
  assign N5791 = N4228 & en_i;
  assign N5792 = ~valid[390];
  assign match_array[391] = N5794 & valid[391];
  assign N5794 = N5793 & N3496;
  assign N5793 = N4228 & en_i;
  assign empty_array[391] = N5795 & N5796;
  assign N5795 = N4228 & en_i;
  assign N5796 = ~valid[391];
  assign match_array[392] = N5798 & valid[392];
  assign N5798 = N5797 & N3497;
  assign N5797 = N4228 & en_i;
  assign empty_array[392] = N5799 & N5800;
  assign N5799 = N4228 & en_i;
  assign N5800 = ~valid[392];
  assign match_array[393] = N5802 & valid[393];
  assign N5802 = N5801 & N3498;
  assign N5801 = N4228 & en_i;
  assign empty_array[393] = N5803 & N5804;
  assign N5803 = N4228 & en_i;
  assign N5804 = ~valid[393];
  assign match_array[394] = N5806 & valid[394];
  assign N5806 = N5805 & N3499;
  assign N5805 = N4228 & en_i;
  assign empty_array[394] = N5807 & N5808;
  assign N5807 = N4228 & en_i;
  assign N5808 = ~valid[394];
  assign match_array[395] = N5810 & valid[395];
  assign N5810 = N5809 & N3500;
  assign N5809 = N4228 & en_i;
  assign empty_array[395] = N5811 & N5812;
  assign N5811 = N4228 & en_i;
  assign N5812 = ~valid[395];
  assign match_array[396] = N5814 & valid[396];
  assign N5814 = N5813 & N3501;
  assign N5813 = N4228 & en_i;
  assign empty_array[396] = N5815 & N5816;
  assign N5815 = N4228 & en_i;
  assign N5816 = ~valid[396];
  assign match_array[397] = N5818 & valid[397];
  assign N5818 = N5817 & N3502;
  assign N5817 = N4228 & en_i;
  assign empty_array[397] = N5819 & N5820;
  assign N5819 = N4228 & en_i;
  assign N5820 = ~valid[397];
  assign match_array[398] = N5822 & valid[398];
  assign N5822 = N5821 & N3503;
  assign N5821 = N4228 & en_i;
  assign empty_array[398] = N5823 & N5824;
  assign N5823 = N4228 & en_i;
  assign N5824 = ~valid[398];
  assign match_array[399] = N5826 & valid[399];
  assign N5826 = N5825 & N3504;
  assign N5825 = N4228 & en_i;
  assign empty_array[399] = N5827 & N5828;
  assign N5827 = N4228 & en_i;
  assign N5828 = ~valid[399];
  assign match_array[400] = N5830 & valid[400];
  assign N5830 = N5829 & N3505;
  assign N5829 = N4228 & en_i;
  assign empty_array[400] = N5831 & N5832;
  assign N5831 = N4228 & en_i;
  assign N5832 = ~valid[400];
  assign match_array[401] = N5834 & valid[401];
  assign N5834 = N5833 & N3506;
  assign N5833 = N4228 & en_i;
  assign empty_array[401] = N5835 & N5836;
  assign N5835 = N4228 & en_i;
  assign N5836 = ~valid[401];
  assign match_array[402] = N5838 & valid[402];
  assign N5838 = N5837 & N3507;
  assign N5837 = N4228 & en_i;
  assign empty_array[402] = N5839 & N5840;
  assign N5839 = N4228 & en_i;
  assign N5840 = ~valid[402];
  assign match_array[403] = N5842 & valid[403];
  assign N5842 = N5841 & N3508;
  assign N5841 = N4228 & en_i;
  assign empty_array[403] = N5843 & N5844;
  assign N5843 = N4228 & en_i;
  assign N5844 = ~valid[403];
  assign match_array[404] = N5846 & valid[404];
  assign N5846 = N5845 & N3509;
  assign N5845 = N4228 & en_i;
  assign empty_array[404] = N5847 & N5848;
  assign N5847 = N4228 & en_i;
  assign N5848 = ~valid[404];
  assign match_array[405] = N5850 & valid[405];
  assign N5850 = N5849 & N3510;
  assign N5849 = N4228 & en_i;
  assign empty_array[405] = N5851 & N5852;
  assign N5851 = N4228 & en_i;
  assign N5852 = ~valid[405];
  assign match_array[406] = N5854 & valid[406];
  assign N5854 = N5853 & N3511;
  assign N5853 = N4228 & en_i;
  assign empty_array[406] = N5855 & N5856;
  assign N5855 = N4228 & en_i;
  assign N5856 = ~valid[406];
  assign match_array[407] = N5858 & valid[407];
  assign N5858 = N5857 & N3512;
  assign N5857 = N4228 & en_i;
  assign empty_array[407] = N5859 & N5860;
  assign N5859 = N4228 & en_i;
  assign N5860 = ~valid[407];
  assign match_array[408] = N5862 & valid[408];
  assign N5862 = N5861 & N3513;
  assign N5861 = N4228 & en_i;
  assign empty_array[408] = N5863 & N5864;
  assign N5863 = N4228 & en_i;
  assign N5864 = ~valid[408];
  assign match_array[409] = N5866 & valid[409];
  assign N5866 = N5865 & N3514;
  assign N5865 = N4228 & en_i;
  assign empty_array[409] = N5867 & N5868;
  assign N5867 = N4228 & en_i;
  assign N5868 = ~valid[409];
  assign match_array[410] = N5870 & valid[410];
  assign N5870 = N5869 & N3515;
  assign N5869 = N4228 & en_i;
  assign empty_array[410] = N5871 & N5872;
  assign N5871 = N4228 & en_i;
  assign N5872 = ~valid[410];
  assign match_array[411] = N5874 & valid[411];
  assign N5874 = N5873 & N3516;
  assign N5873 = N4228 & en_i;
  assign empty_array[411] = N5875 & N5876;
  assign N5875 = N4228 & en_i;
  assign N5876 = ~valid[411];
  assign match_array[412] = N5878 & valid[412];
  assign N5878 = N5877 & N3517;
  assign N5877 = N4228 & en_i;
  assign empty_array[412] = N5879 & N5880;
  assign N5879 = N4228 & en_i;
  assign N5880 = ~valid[412];
  assign match_array[413] = N5882 & valid[413];
  assign N5882 = N5881 & N3518;
  assign N5881 = N4228 & en_i;
  assign empty_array[413] = N5883 & N5884;
  assign N5883 = N4228 & en_i;
  assign N5884 = ~valid[413];
  assign match_array[414] = N5886 & valid[414];
  assign N5886 = N5885 & N3519;
  assign N5885 = N4228 & en_i;
  assign empty_array[414] = N5887 & N5888;
  assign N5887 = N4228 & en_i;
  assign N5888 = ~valid[414];
  assign match_array[415] = N5890 & valid[415];
  assign N5890 = N5889 & N3520;
  assign N5889 = N4228 & en_i;
  assign empty_array[415] = N5891 & N5892;
  assign N5891 = N4228 & en_i;
  assign N5892 = ~valid[415];
  assign match_array[416] = N5894 & valid[416];
  assign N5894 = N5893 & N3521;
  assign N5893 = N4228 & en_i;
  assign empty_array[416] = N5895 & N5896;
  assign N5895 = N4228 & en_i;
  assign N5896 = ~valid[416];
  assign match_array[417] = N5898 & valid[417];
  assign N5898 = N5897 & N3522;
  assign N5897 = N4228 & en_i;
  assign empty_array[417] = N5899 & N5900;
  assign N5899 = N4228 & en_i;
  assign N5900 = ~valid[417];
  assign match_array[418] = N5902 & valid[418];
  assign N5902 = N5901 & N3523;
  assign N5901 = N4228 & en_i;
  assign empty_array[418] = N5903 & N5904;
  assign N5903 = N4228 & en_i;
  assign N5904 = ~valid[418];
  assign match_array[419] = N5906 & valid[419];
  assign N5906 = N5905 & N3524;
  assign N5905 = N4228 & en_i;
  assign empty_array[419] = N5907 & N5908;
  assign N5907 = N4228 & en_i;
  assign N5908 = ~valid[419];
  assign match_array[420] = N5910 & valid[420];
  assign N5910 = N5909 & N3525;
  assign N5909 = N4228 & en_i;
  assign empty_array[420] = N5911 & N5912;
  assign N5911 = N4228 & en_i;
  assign N5912 = ~valid[420];
  assign match_array[421] = N5914 & valid[421];
  assign N5914 = N5913 & N3526;
  assign N5913 = N4228 & en_i;
  assign empty_array[421] = N5915 & N5916;
  assign N5915 = N4228 & en_i;
  assign N5916 = ~valid[421];
  assign match_array[422] = N5918 & valid[422];
  assign N5918 = N5917 & N3527;
  assign N5917 = N4228 & en_i;
  assign empty_array[422] = N5919 & N5920;
  assign N5919 = N4228 & en_i;
  assign N5920 = ~valid[422];
  assign match_array[423] = N5922 & valid[423];
  assign N5922 = N5921 & N3528;
  assign N5921 = N4228 & en_i;
  assign empty_array[423] = N5923 & N5924;
  assign N5923 = N4228 & en_i;
  assign N5924 = ~valid[423];
  assign match_array[424] = N5926 & valid[424];
  assign N5926 = N5925 & N3529;
  assign N5925 = N4228 & en_i;
  assign empty_array[424] = N5927 & N5928;
  assign N5927 = N4228 & en_i;
  assign N5928 = ~valid[424];
  assign match_array[425] = N5930 & valid[425];
  assign N5930 = N5929 & N3530;
  assign N5929 = N4228 & en_i;
  assign empty_array[425] = N5931 & N5932;
  assign N5931 = N4228 & en_i;
  assign N5932 = ~valid[425];
  assign match_array[426] = N5934 & valid[426];
  assign N5934 = N5933 & N3531;
  assign N5933 = N4228 & en_i;
  assign empty_array[426] = N5935 & N5936;
  assign N5935 = N4228 & en_i;
  assign N5936 = ~valid[426];
  assign match_array[427] = N5938 & valid[427];
  assign N5938 = N5937 & N3532;
  assign N5937 = N4228 & en_i;
  assign empty_array[427] = N5939 & N5940;
  assign N5939 = N4228 & en_i;
  assign N5940 = ~valid[427];
  assign match_array[428] = N5942 & valid[428];
  assign N5942 = N5941 & N3533;
  assign N5941 = N4228 & en_i;
  assign empty_array[428] = N5943 & N5944;
  assign N5943 = N4228 & en_i;
  assign N5944 = ~valid[428];
  assign match_array[429] = N5946 & valid[429];
  assign N5946 = N5945 & N3534;
  assign N5945 = N4228 & en_i;
  assign empty_array[429] = N5947 & N5948;
  assign N5947 = N4228 & en_i;
  assign N5948 = ~valid[429];
  assign match_array[430] = N5950 & valid[430];
  assign N5950 = N5949 & N3535;
  assign N5949 = N4228 & en_i;
  assign empty_array[430] = N5951 & N5952;
  assign N5951 = N4228 & en_i;
  assign N5952 = ~valid[430];
  assign match_array[431] = N5954 & valid[431];
  assign N5954 = N5953 & N3536;
  assign N5953 = N4228 & en_i;
  assign empty_array[431] = N5955 & N5956;
  assign N5955 = N4228 & en_i;
  assign N5956 = ~valid[431];
  assign match_array[432] = N5958 & valid[432];
  assign N5958 = N5957 & N3537;
  assign N5957 = N4228 & en_i;
  assign empty_array[432] = N5959 & N5960;
  assign N5959 = N4228 & en_i;
  assign N5960 = ~valid[432];
  assign match_array[433] = N5962 & valid[433];
  assign N5962 = N5961 & N3538;
  assign N5961 = N4228 & en_i;
  assign empty_array[433] = N5963 & N5964;
  assign N5963 = N4228 & en_i;
  assign N5964 = ~valid[433];
  assign match_array[434] = N5966 & valid[434];
  assign N5966 = N5965 & N3539;
  assign N5965 = N4228 & en_i;
  assign empty_array[434] = N5967 & N5968;
  assign N5967 = N4228 & en_i;
  assign N5968 = ~valid[434];
  assign match_array[435] = N5970 & valid[435];
  assign N5970 = N5969 & N3540;
  assign N5969 = N4228 & en_i;
  assign empty_array[435] = N5971 & N5972;
  assign N5971 = N4228 & en_i;
  assign N5972 = ~valid[435];
  assign match_array[436] = N5974 & valid[436];
  assign N5974 = N5973 & N3541;
  assign N5973 = N4228 & en_i;
  assign empty_array[436] = N5975 & N5976;
  assign N5975 = N4228 & en_i;
  assign N5976 = ~valid[436];
  assign match_array[437] = N5978 & valid[437];
  assign N5978 = N5977 & N3542;
  assign N5977 = N4228 & en_i;
  assign empty_array[437] = N5979 & N5980;
  assign N5979 = N4228 & en_i;
  assign N5980 = ~valid[437];
  assign match_array[438] = N5982 & valid[438];
  assign N5982 = N5981 & N3543;
  assign N5981 = N4228 & en_i;
  assign empty_array[438] = N5983 & N5984;
  assign N5983 = N4228 & en_i;
  assign N5984 = ~valid[438];
  assign match_array[439] = N5986 & valid[439];
  assign N5986 = N5985 & N3544;
  assign N5985 = N4228 & en_i;
  assign empty_array[439] = N5987 & N5988;
  assign N5987 = N4228 & en_i;
  assign N5988 = ~valid[439];
  assign match_array[440] = N5990 & valid[440];
  assign N5990 = N5989 & N3545;
  assign N5989 = N4228 & en_i;
  assign empty_array[440] = N5991 & N5992;
  assign N5991 = N4228 & en_i;
  assign N5992 = ~valid[440];
  assign match_array[441] = N5994 & valid[441];
  assign N5994 = N5993 & N3546;
  assign N5993 = N4228 & en_i;
  assign empty_array[441] = N5995 & N5996;
  assign N5995 = N4228 & en_i;
  assign N5996 = ~valid[441];
  assign match_array[442] = N5998 & valid[442];
  assign N5998 = N5997 & N3547;
  assign N5997 = N4228 & en_i;
  assign empty_array[442] = N5999 & N6000;
  assign N5999 = N4228 & en_i;
  assign N6000 = ~valid[442];
  assign match_array[443] = N6002 & valid[443];
  assign N6002 = N6001 & N3548;
  assign N6001 = N4228 & en_i;
  assign empty_array[443] = N6003 & N6004;
  assign N6003 = N4228 & en_i;
  assign N6004 = ~valid[443];
  assign match_array[444] = N6006 & valid[444];
  assign N6006 = N6005 & N3549;
  assign N6005 = N4228 & en_i;
  assign empty_array[444] = N6007 & N6008;
  assign N6007 = N4228 & en_i;
  assign N6008 = ~valid[444];
  assign match_array[445] = N6010 & valid[445];
  assign N6010 = N6009 & N3550;
  assign N6009 = N4228 & en_i;
  assign empty_array[445] = N6011 & N6012;
  assign N6011 = N4228 & en_i;
  assign N6012 = ~valid[445];
  assign match_array[446] = N6014 & valid[446];
  assign N6014 = N6013 & N3551;
  assign N6013 = N4228 & en_i;
  assign empty_array[446] = N6015 & N6016;
  assign N6015 = N4228 & en_i;
  assign N6016 = ~valid[446];
  assign match_array[447] = N6018 & valid[447];
  assign N6018 = N6017 & N3552;
  assign N6017 = N4228 & en_i;
  assign empty_array[447] = N6019 & N6020;
  assign N6019 = N4228 & en_i;
  assign N6020 = ~valid[447];
  assign match_array[448] = N6022 & valid[448];
  assign N6022 = N6021 & N3553;
  assign N6021 = N4228 & en_i;
  assign empty_array[448] = N6023 & N6024;
  assign N6023 = N4228 & en_i;
  assign N6024 = ~valid[448];
  assign match_array[449] = N6026 & valid[449];
  assign N6026 = N6025 & N3554;
  assign N6025 = N4228 & en_i;
  assign empty_array[449] = N6027 & N6028;
  assign N6027 = N4228 & en_i;
  assign N6028 = ~valid[449];
  assign match_array[450] = N6030 & valid[450];
  assign N6030 = N6029 & N3555;
  assign N6029 = N4228 & en_i;
  assign empty_array[450] = N6031 & N6032;
  assign N6031 = N4228 & en_i;
  assign N6032 = ~valid[450];
  assign match_array[451] = N6034 & valid[451];
  assign N6034 = N6033 & N3556;
  assign N6033 = N4228 & en_i;
  assign empty_array[451] = N6035 & N6036;
  assign N6035 = N4228 & en_i;
  assign N6036 = ~valid[451];
  assign match_array[452] = N6038 & valid[452];
  assign N6038 = N6037 & N3557;
  assign N6037 = N4228 & en_i;
  assign empty_array[452] = N6039 & N6040;
  assign N6039 = N4228 & en_i;
  assign N6040 = ~valid[452];
  assign match_array[453] = N6042 & valid[453];
  assign N6042 = N6041 & N3558;
  assign N6041 = N4228 & en_i;
  assign empty_array[453] = N6043 & N6044;
  assign N6043 = N4228 & en_i;
  assign N6044 = ~valid[453];
  assign match_array[454] = N6046 & valid[454];
  assign N6046 = N6045 & N3559;
  assign N6045 = N4228 & en_i;
  assign empty_array[454] = N6047 & N6048;
  assign N6047 = N4228 & en_i;
  assign N6048 = ~valid[454];
  assign match_array[455] = N6050 & valid[455];
  assign N6050 = N6049 & N3560;
  assign N6049 = N4228 & en_i;
  assign empty_array[455] = N6051 & N6052;
  assign N6051 = N4228 & en_i;
  assign N6052 = ~valid[455];
  assign match_array[456] = N6054 & valid[456];
  assign N6054 = N6053 & N3561;
  assign N6053 = N4228 & en_i;
  assign empty_array[456] = N6055 & N6056;
  assign N6055 = N4228 & en_i;
  assign N6056 = ~valid[456];
  assign match_array[457] = N6058 & valid[457];
  assign N6058 = N6057 & N3562;
  assign N6057 = N4228 & en_i;
  assign empty_array[457] = N6059 & N6060;
  assign N6059 = N4228 & en_i;
  assign N6060 = ~valid[457];
  assign match_array[458] = N6062 & valid[458];
  assign N6062 = N6061 & N3563;
  assign N6061 = N4228 & en_i;
  assign empty_array[458] = N6063 & N6064;
  assign N6063 = N4228 & en_i;
  assign N6064 = ~valid[458];
  assign match_array[459] = N6066 & valid[459];
  assign N6066 = N6065 & N3564;
  assign N6065 = N4228 & en_i;
  assign empty_array[459] = N6067 & N6068;
  assign N6067 = N4228 & en_i;
  assign N6068 = ~valid[459];
  assign match_array[460] = N6070 & valid[460];
  assign N6070 = N6069 & N3565;
  assign N6069 = N4228 & en_i;
  assign empty_array[460] = N6071 & N6072;
  assign N6071 = N4228 & en_i;
  assign N6072 = ~valid[460];
  assign match_array[461] = N6074 & valid[461];
  assign N6074 = N6073 & N3566;
  assign N6073 = N4228 & en_i;
  assign empty_array[461] = N6075 & N6076;
  assign N6075 = N4228 & en_i;
  assign N6076 = ~valid[461];
  assign match_array[462] = N6078 & valid[462];
  assign N6078 = N6077 & N3567;
  assign N6077 = N4228 & en_i;
  assign empty_array[462] = N6079 & N6080;
  assign N6079 = N4228 & en_i;
  assign N6080 = ~valid[462];
  assign match_array[463] = N6082 & valid[463];
  assign N6082 = N6081 & N3568;
  assign N6081 = N4228 & en_i;
  assign empty_array[463] = N6083 & N6084;
  assign N6083 = N4228 & en_i;
  assign N6084 = ~valid[463];
  assign match_array[464] = N6086 & valid[464];
  assign N6086 = N6085 & N3569;
  assign N6085 = N4228 & en_i;
  assign empty_array[464] = N6087 & N6088;
  assign N6087 = N4228 & en_i;
  assign N6088 = ~valid[464];
  assign match_array[465] = N6090 & valid[465];
  assign N6090 = N6089 & N3570;
  assign N6089 = N4228 & en_i;
  assign empty_array[465] = N6091 & N6092;
  assign N6091 = N4228 & en_i;
  assign N6092 = ~valid[465];
  assign match_array[466] = N6094 & valid[466];
  assign N6094 = N6093 & N3571;
  assign N6093 = N4228 & en_i;
  assign empty_array[466] = N6095 & N6096;
  assign N6095 = N4228 & en_i;
  assign N6096 = ~valid[466];
  assign match_array[467] = N6098 & valid[467];
  assign N6098 = N6097 & N3572;
  assign N6097 = N4228 & en_i;
  assign empty_array[467] = N6099 & N6100;
  assign N6099 = N4228 & en_i;
  assign N6100 = ~valid[467];
  assign match_array[468] = N6102 & valid[468];
  assign N6102 = N6101 & N3573;
  assign N6101 = N4228 & en_i;
  assign empty_array[468] = N6103 & N6104;
  assign N6103 = N4228 & en_i;
  assign N6104 = ~valid[468];
  assign match_array[469] = N6106 & valid[469];
  assign N6106 = N6105 & N3574;
  assign N6105 = N4228 & en_i;
  assign empty_array[469] = N6107 & N6108;
  assign N6107 = N4228 & en_i;
  assign N6108 = ~valid[469];
  assign match_array[470] = N6110 & valid[470];
  assign N6110 = N6109 & N3575;
  assign N6109 = N4228 & en_i;
  assign empty_array[470] = N6111 & N6112;
  assign N6111 = N4228 & en_i;
  assign N6112 = ~valid[470];
  assign match_array[471] = N6114 & valid[471];
  assign N6114 = N6113 & N3576;
  assign N6113 = N4228 & en_i;
  assign empty_array[471] = N6115 & N6116;
  assign N6115 = N4228 & en_i;
  assign N6116 = ~valid[471];
  assign match_array[472] = N6118 & valid[472];
  assign N6118 = N6117 & N3577;
  assign N6117 = N4228 & en_i;
  assign empty_array[472] = N6119 & N6120;
  assign N6119 = N4228 & en_i;
  assign N6120 = ~valid[472];
  assign match_array[473] = N6122 & valid[473];
  assign N6122 = N6121 & N3578;
  assign N6121 = N4228 & en_i;
  assign empty_array[473] = N6123 & N6124;
  assign N6123 = N4228 & en_i;
  assign N6124 = ~valid[473];
  assign match_array[474] = N6126 & valid[474];
  assign N6126 = N6125 & N3579;
  assign N6125 = N4228 & en_i;
  assign empty_array[474] = N6127 & N6128;
  assign N6127 = N4228 & en_i;
  assign N6128 = ~valid[474];
  assign match_array[475] = N6130 & valid[475];
  assign N6130 = N6129 & N3580;
  assign N6129 = N4228 & en_i;
  assign empty_array[475] = N6131 & N6132;
  assign N6131 = N4228 & en_i;
  assign N6132 = ~valid[475];
  assign match_array[476] = N6134 & valid[476];
  assign N6134 = N6133 & N3581;
  assign N6133 = N4228 & en_i;
  assign empty_array[476] = N6135 & N6136;
  assign N6135 = N4228 & en_i;
  assign N6136 = ~valid[476];
  assign match_array[477] = N6138 & valid[477];
  assign N6138 = N6137 & N3582;
  assign N6137 = N4228 & en_i;
  assign empty_array[477] = N6139 & N6140;
  assign N6139 = N4228 & en_i;
  assign N6140 = ~valid[477];
  assign match_array[478] = N6142 & valid[478];
  assign N6142 = N6141 & N3583;
  assign N6141 = N4228 & en_i;
  assign empty_array[478] = N6143 & N6144;
  assign N6143 = N4228 & en_i;
  assign N6144 = ~valid[478];
  assign match_array[479] = N6146 & valid[479];
  assign N6146 = N6145 & N3584;
  assign N6145 = N4228 & en_i;
  assign empty_array[479] = N6147 & N6148;
  assign N6147 = N4228 & en_i;
  assign N6148 = ~valid[479];
  assign match_array[480] = N6150 & valid[480];
  assign N6150 = N6149 & N3585;
  assign N6149 = N4228 & en_i;
  assign empty_array[480] = N6151 & N6152;
  assign N6151 = N4228 & en_i;
  assign N6152 = ~valid[480];
  assign match_array[481] = N6154 & valid[481];
  assign N6154 = N6153 & N3586;
  assign N6153 = N4228 & en_i;
  assign empty_array[481] = N6155 & N6156;
  assign N6155 = N4228 & en_i;
  assign N6156 = ~valid[481];
  assign match_array[482] = N6158 & valid[482];
  assign N6158 = N6157 & N3587;
  assign N6157 = N4228 & en_i;
  assign empty_array[482] = N6159 & N6160;
  assign N6159 = N4228 & en_i;
  assign N6160 = ~valid[482];
  assign match_array[483] = N6162 & valid[483];
  assign N6162 = N6161 & N3588;
  assign N6161 = N4228 & en_i;
  assign empty_array[483] = N6163 & N6164;
  assign N6163 = N4228 & en_i;
  assign N6164 = ~valid[483];
  assign match_array[484] = N6166 & valid[484];
  assign N6166 = N6165 & N3589;
  assign N6165 = N4228 & en_i;
  assign empty_array[484] = N6167 & N6168;
  assign N6167 = N4228 & en_i;
  assign N6168 = ~valid[484];
  assign match_array[485] = N6170 & valid[485];
  assign N6170 = N6169 & N3590;
  assign N6169 = N4228 & en_i;
  assign empty_array[485] = N6171 & N6172;
  assign N6171 = N4228 & en_i;
  assign N6172 = ~valid[485];
  assign match_array[486] = N6174 & valid[486];
  assign N6174 = N6173 & N3591;
  assign N6173 = N4228 & en_i;
  assign empty_array[486] = N6175 & N6176;
  assign N6175 = N4228 & en_i;
  assign N6176 = ~valid[486];
  assign match_array[487] = N6178 & valid[487];
  assign N6178 = N6177 & N3592;
  assign N6177 = N4228 & en_i;
  assign empty_array[487] = N6179 & N6180;
  assign N6179 = N4228 & en_i;
  assign N6180 = ~valid[487];
  assign match_array[488] = N6182 & valid[488];
  assign N6182 = N6181 & N3593;
  assign N6181 = N4228 & en_i;
  assign empty_array[488] = N6183 & N6184;
  assign N6183 = N4228 & en_i;
  assign N6184 = ~valid[488];
  assign match_array[489] = N6186 & valid[489];
  assign N6186 = N6185 & N3594;
  assign N6185 = N4228 & en_i;
  assign empty_array[489] = N6187 & N6188;
  assign N6187 = N4228 & en_i;
  assign N6188 = ~valid[489];
  assign match_array[490] = N6190 & valid[490];
  assign N6190 = N6189 & N3595;
  assign N6189 = N4228 & en_i;
  assign empty_array[490] = N6191 & N6192;
  assign N6191 = N4228 & en_i;
  assign N6192 = ~valid[490];
  assign match_array[491] = N6194 & valid[491];
  assign N6194 = N6193 & N3596;
  assign N6193 = N4228 & en_i;
  assign empty_array[491] = N6195 & N6196;
  assign N6195 = N4228 & en_i;
  assign N6196 = ~valid[491];
  assign match_array[492] = N6198 & valid[492];
  assign N6198 = N6197 & N3597;
  assign N6197 = N4228 & en_i;
  assign empty_array[492] = N6199 & N6200;
  assign N6199 = N4228 & en_i;
  assign N6200 = ~valid[492];
  assign match_array[493] = N6202 & valid[493];
  assign N6202 = N6201 & N3598;
  assign N6201 = N4228 & en_i;
  assign empty_array[493] = N6203 & N6204;
  assign N6203 = N4228 & en_i;
  assign N6204 = ~valid[493];
  assign match_array[494] = N6206 & valid[494];
  assign N6206 = N6205 & N3599;
  assign N6205 = N4228 & en_i;
  assign empty_array[494] = N6207 & N6208;
  assign N6207 = N4228 & en_i;
  assign N6208 = ~valid[494];
  assign match_array[495] = N6210 & valid[495];
  assign N6210 = N6209 & N3600;
  assign N6209 = N4228 & en_i;
  assign empty_array[495] = N6211 & N6212;
  assign N6211 = N4228 & en_i;
  assign N6212 = ~valid[495];
  assign match_array[496] = N6214 & valid[496];
  assign N6214 = N6213 & N3601;
  assign N6213 = N4228 & en_i;
  assign empty_array[496] = N6215 & N6216;
  assign N6215 = N4228 & en_i;
  assign N6216 = ~valid[496];
  assign match_array[497] = N6218 & valid[497];
  assign N6218 = N6217 & N3602;
  assign N6217 = N4228 & en_i;
  assign empty_array[497] = N6219 & N6220;
  assign N6219 = N4228 & en_i;
  assign N6220 = ~valid[497];
  assign match_array[498] = N6222 & valid[498];
  assign N6222 = N6221 & N3603;
  assign N6221 = N4228 & en_i;
  assign empty_array[498] = N6223 & N6224;
  assign N6223 = N4228 & en_i;
  assign N6224 = ~valid[498];
  assign match_array[499] = N6226 & valid[499];
  assign N6226 = N6225 & N3604;
  assign N6225 = N4228 & en_i;
  assign empty_array[499] = N6227 & N6228;
  assign N6227 = N4228 & en_i;
  assign N6228 = ~valid[499];
  assign match_array[500] = N6230 & valid[500];
  assign N6230 = N6229 & N3605;
  assign N6229 = N4228 & en_i;
  assign empty_array[500] = N6231 & N6232;
  assign N6231 = N4228 & en_i;
  assign N6232 = ~valid[500];
  assign match_array[501] = N6234 & valid[501];
  assign N6234 = N6233 & N3606;
  assign N6233 = N4228 & en_i;
  assign empty_array[501] = N6235 & N6236;
  assign N6235 = N4228 & en_i;
  assign N6236 = ~valid[501];
  assign match_array[502] = N6238 & valid[502];
  assign N6238 = N6237 & N3607;
  assign N6237 = N4228 & en_i;
  assign empty_array[502] = N6239 & N6240;
  assign N6239 = N4228 & en_i;
  assign N6240 = ~valid[502];
  assign match_array[503] = N6242 & valid[503];
  assign N6242 = N6241 & N3608;
  assign N6241 = N4228 & en_i;
  assign empty_array[503] = N6243 & N6244;
  assign N6243 = N4228 & en_i;
  assign N6244 = ~valid[503];
  assign match_array[504] = N6246 & valid[504];
  assign N6246 = N6245 & N3609;
  assign N6245 = N4228 & en_i;
  assign empty_array[504] = N6247 & N6248;
  assign N6247 = N4228 & en_i;
  assign N6248 = ~valid[504];
  assign match_array[505] = N6250 & valid[505];
  assign N6250 = N6249 & N3610;
  assign N6249 = N4228 & en_i;
  assign empty_array[505] = N6251 & N6252;
  assign N6251 = N4228 & en_i;
  assign N6252 = ~valid[505];
  assign match_array[506] = N6254 & valid[506];
  assign N6254 = N6253 & N3611;
  assign N6253 = N4228 & en_i;
  assign empty_array[506] = N6255 & N6256;
  assign N6255 = N4228 & en_i;
  assign N6256 = ~valid[506];
  assign match_array[507] = N6258 & valid[507];
  assign N6258 = N6257 & N3612;
  assign N6257 = N4228 & en_i;
  assign empty_array[507] = N6259 & N6260;
  assign N6259 = N4228 & en_i;
  assign N6260 = ~valid[507];
  assign match_array[508] = N6262 & valid[508];
  assign N6262 = N6261 & N3613;
  assign N6261 = N4228 & en_i;
  assign empty_array[508] = N6263 & N6264;
  assign N6263 = N4228 & en_i;
  assign N6264 = ~valid[508];
  assign match_array[509] = N6266 & valid[509];
  assign N6266 = N6265 & N3614;
  assign N6265 = N4228 & en_i;
  assign empty_array[509] = N6267 & N6268;
  assign N6267 = N4228 & en_i;
  assign N6268 = ~valid[509];
  assign match_array[510] = N6270 & valid[510];
  assign N6270 = N6269 & N3615;
  assign N6269 = N4228 & en_i;
  assign empty_array[510] = N6271 & N6272;
  assign N6271 = N4228 & en_i;
  assign N6272 = ~valid[510];
  assign match_array[511] = N6274 & valid[511];
  assign N6274 = N6273 & N3616;
  assign N6273 = N4228 & en_i;
  assign empty_array[511] = N6275 & N6276;
  assign N6275 = N4228 & en_i;
  assign N6276 = ~valid[511];
  assign match_array[512] = N6278 & valid[512];
  assign N6278 = N6277 & N3617;
  assign N6277 = N4228 & en_i;
  assign empty_array[512] = N6279 & N6280;
  assign N6279 = N4228 & en_i;
  assign N6280 = ~valid[512];
  assign match_array[513] = N6282 & valid[513];
  assign N6282 = N6281 & N3618;
  assign N6281 = N4228 & en_i;
  assign empty_array[513] = N6283 & N6284;
  assign N6283 = N4228 & en_i;
  assign N6284 = ~valid[513];
  assign match_array[514] = N6286 & valid[514];
  assign N6286 = N6285 & N3619;
  assign N6285 = N4228 & en_i;
  assign empty_array[514] = N6287 & N6288;
  assign N6287 = N4228 & en_i;
  assign N6288 = ~valid[514];
  assign match_array[515] = N6290 & valid[515];
  assign N6290 = N6289 & N3620;
  assign N6289 = N4228 & en_i;
  assign empty_array[515] = N6291 & N6292;
  assign N6291 = N4228 & en_i;
  assign N6292 = ~valid[515];
  assign match_array[516] = N6294 & valid[516];
  assign N6294 = N6293 & N3621;
  assign N6293 = N4228 & en_i;
  assign empty_array[516] = N6295 & N6296;
  assign N6295 = N4228 & en_i;
  assign N6296 = ~valid[516];
  assign match_array[517] = N6298 & valid[517];
  assign N6298 = N6297 & N3622;
  assign N6297 = N4228 & en_i;
  assign empty_array[517] = N6299 & N6300;
  assign N6299 = N4228 & en_i;
  assign N6300 = ~valid[517];
  assign match_array[518] = N6302 & valid[518];
  assign N6302 = N6301 & N3623;
  assign N6301 = N4228 & en_i;
  assign empty_array[518] = N6303 & N6304;
  assign N6303 = N4228 & en_i;
  assign N6304 = ~valid[518];
  assign match_array[519] = N6306 & valid[519];
  assign N6306 = N6305 & N3624;
  assign N6305 = N4228 & en_i;
  assign empty_array[519] = N6307 & N6308;
  assign N6307 = N4228 & en_i;
  assign N6308 = ~valid[519];
  assign match_array[520] = N6310 & valid[520];
  assign N6310 = N6309 & N3625;
  assign N6309 = N4228 & en_i;
  assign empty_array[520] = N6311 & N6312;
  assign N6311 = N4228 & en_i;
  assign N6312 = ~valid[520];
  assign match_array[521] = N6314 & valid[521];
  assign N6314 = N6313 & N3626;
  assign N6313 = N4228 & en_i;
  assign empty_array[521] = N6315 & N6316;
  assign N6315 = N4228 & en_i;
  assign N6316 = ~valid[521];
  assign match_array[522] = N6318 & valid[522];
  assign N6318 = N6317 & N3627;
  assign N6317 = N4228 & en_i;
  assign empty_array[522] = N6319 & N6320;
  assign N6319 = N4228 & en_i;
  assign N6320 = ~valid[522];
  assign match_array[523] = N6322 & valid[523];
  assign N6322 = N6321 & N3628;
  assign N6321 = N4228 & en_i;
  assign empty_array[523] = N6323 & N6324;
  assign N6323 = N4228 & en_i;
  assign N6324 = ~valid[523];
  assign match_array[524] = N6326 & valid[524];
  assign N6326 = N6325 & N3629;
  assign N6325 = N4228 & en_i;
  assign empty_array[524] = N6327 & N6328;
  assign N6327 = N4228 & en_i;
  assign N6328 = ~valid[524];
  assign match_array[525] = N6330 & valid[525];
  assign N6330 = N6329 & N3630;
  assign N6329 = N4228 & en_i;
  assign empty_array[525] = N6331 & N6332;
  assign N6331 = N4228 & en_i;
  assign N6332 = ~valid[525];
  assign match_array[526] = N6334 & valid[526];
  assign N6334 = N6333 & N3631;
  assign N6333 = N4228 & en_i;
  assign empty_array[526] = N6335 & N6336;
  assign N6335 = N4228 & en_i;
  assign N6336 = ~valid[526];
  assign match_array[527] = N6338 & valid[527];
  assign N6338 = N6337 & N3632;
  assign N6337 = N4228 & en_i;
  assign empty_array[527] = N6339 & N6340;
  assign N6339 = N4228 & en_i;
  assign N6340 = ~valid[527];
  assign match_array[528] = N6342 & valid[528];
  assign N6342 = N6341 & N3633;
  assign N6341 = N4228 & en_i;
  assign empty_array[528] = N6343 & N6344;
  assign N6343 = N4228 & en_i;
  assign N6344 = ~valid[528];
  assign match_array[529] = N6346 & valid[529];
  assign N6346 = N6345 & N3634;
  assign N6345 = N4228 & en_i;
  assign empty_array[529] = N6347 & N6348;
  assign N6347 = N4228 & en_i;
  assign N6348 = ~valid[529];
  assign match_array[530] = N6350 & valid[530];
  assign N6350 = N6349 & N3635;
  assign N6349 = N4228 & en_i;
  assign empty_array[530] = N6351 & N6352;
  assign N6351 = N4228 & en_i;
  assign N6352 = ~valid[530];
  assign match_array[531] = N6354 & valid[531];
  assign N6354 = N6353 & N3636;
  assign N6353 = N4228 & en_i;
  assign empty_array[531] = N6355 & N6356;
  assign N6355 = N4228 & en_i;
  assign N6356 = ~valid[531];
  assign match_array[532] = N6358 & valid[532];
  assign N6358 = N6357 & N3637;
  assign N6357 = N4228 & en_i;
  assign empty_array[532] = N6359 & N6360;
  assign N6359 = N4228 & en_i;
  assign N6360 = ~valid[532];
  assign match_array[533] = N6362 & valid[533];
  assign N6362 = N6361 & N3638;
  assign N6361 = N4228 & en_i;
  assign empty_array[533] = N6363 & N6364;
  assign N6363 = N4228 & en_i;
  assign N6364 = ~valid[533];
  assign match_array[534] = N6366 & valid[534];
  assign N6366 = N6365 & N3639;
  assign N6365 = N4228 & en_i;
  assign empty_array[534] = N6367 & N6368;
  assign N6367 = N4228 & en_i;
  assign N6368 = ~valid[534];
  assign match_array[535] = N6370 & valid[535];
  assign N6370 = N6369 & N3640;
  assign N6369 = N4228 & en_i;
  assign empty_array[535] = N6371 & N6372;
  assign N6371 = N4228 & en_i;
  assign N6372 = ~valid[535];
  assign match_array[536] = N6374 & valid[536];
  assign N6374 = N6373 & N3641;
  assign N6373 = N4228 & en_i;
  assign empty_array[536] = N6375 & N6376;
  assign N6375 = N4228 & en_i;
  assign N6376 = ~valid[536];
  assign match_array[537] = N6378 & valid[537];
  assign N6378 = N6377 & N3642;
  assign N6377 = N4228 & en_i;
  assign empty_array[537] = N6379 & N6380;
  assign N6379 = N4228 & en_i;
  assign N6380 = ~valid[537];
  assign match_array[538] = N6382 & valid[538];
  assign N6382 = N6381 & N3643;
  assign N6381 = N4228 & en_i;
  assign empty_array[538] = N6383 & N6384;
  assign N6383 = N4228 & en_i;
  assign N6384 = ~valid[538];
  assign match_array[539] = N6386 & valid[539];
  assign N6386 = N6385 & N3644;
  assign N6385 = N4228 & en_i;
  assign empty_array[539] = N6387 & N6388;
  assign N6387 = N4228 & en_i;
  assign N6388 = ~valid[539];
  assign match_array[540] = N6390 & valid[540];
  assign N6390 = N6389 & N3645;
  assign N6389 = N4228 & en_i;
  assign empty_array[540] = N6391 & N6392;
  assign N6391 = N4228 & en_i;
  assign N6392 = ~valid[540];
  assign match_array[541] = N6394 & valid[541];
  assign N6394 = N6393 & N3646;
  assign N6393 = N4228 & en_i;
  assign empty_array[541] = N6395 & N6396;
  assign N6395 = N4228 & en_i;
  assign N6396 = ~valid[541];
  assign match_array[542] = N6398 & valid[542];
  assign N6398 = N6397 & N3647;
  assign N6397 = N4228 & en_i;
  assign empty_array[542] = N6399 & N6400;
  assign N6399 = N4228 & en_i;
  assign N6400 = ~valid[542];
  assign match_array[543] = N6402 & valid[543];
  assign N6402 = N6401 & N3648;
  assign N6401 = N4228 & en_i;
  assign empty_array[543] = N6403 & N6404;
  assign N6403 = N4228 & en_i;
  assign N6404 = ~valid[543];
  assign match_array[544] = N6406 & valid[544];
  assign N6406 = N6405 & N3649;
  assign N6405 = N4228 & en_i;
  assign empty_array[544] = N6407 & N6408;
  assign N6407 = N4228 & en_i;
  assign N6408 = ~valid[544];
  assign match_array[545] = N6410 & valid[545];
  assign N6410 = N6409 & N3650;
  assign N6409 = N4228 & en_i;
  assign empty_array[545] = N6411 & N6412;
  assign N6411 = N4228 & en_i;
  assign N6412 = ~valid[545];
  assign match_array[546] = N6414 & valid[546];
  assign N6414 = N6413 & N3651;
  assign N6413 = N4228 & en_i;
  assign empty_array[546] = N6415 & N6416;
  assign N6415 = N4228 & en_i;
  assign N6416 = ~valid[546];
  assign match_array[547] = N6418 & valid[547];
  assign N6418 = N6417 & N3652;
  assign N6417 = N4228 & en_i;
  assign empty_array[547] = N6419 & N6420;
  assign N6419 = N4228 & en_i;
  assign N6420 = ~valid[547];
  assign match_array[548] = N6422 & valid[548];
  assign N6422 = N6421 & N3653;
  assign N6421 = N4228 & en_i;
  assign empty_array[548] = N6423 & N6424;
  assign N6423 = N4228 & en_i;
  assign N6424 = ~valid[548];
  assign match_array[549] = N6426 & valid[549];
  assign N6426 = N6425 & N3654;
  assign N6425 = N4228 & en_i;
  assign empty_array[549] = N6427 & N6428;
  assign N6427 = N4228 & en_i;
  assign N6428 = ~valid[549];
  assign match_array[550] = N6430 & valid[550];
  assign N6430 = N6429 & N3655;
  assign N6429 = N4228 & en_i;
  assign empty_array[550] = N6431 & N6432;
  assign N6431 = N4228 & en_i;
  assign N6432 = ~valid[550];
  assign match_array[551] = N6434 & valid[551];
  assign N6434 = N6433 & N3656;
  assign N6433 = N4228 & en_i;
  assign empty_array[551] = N6435 & N6436;
  assign N6435 = N4228 & en_i;
  assign N6436 = ~valid[551];
  assign match_array[552] = N6438 & valid[552];
  assign N6438 = N6437 & N3657;
  assign N6437 = N4228 & en_i;
  assign empty_array[552] = N6439 & N6440;
  assign N6439 = N4228 & en_i;
  assign N6440 = ~valid[552];
  assign match_array[553] = N6442 & valid[553];
  assign N6442 = N6441 & N3658;
  assign N6441 = N4228 & en_i;
  assign empty_array[553] = N6443 & N6444;
  assign N6443 = N4228 & en_i;
  assign N6444 = ~valid[553];
  assign match_array[554] = N6446 & valid[554];
  assign N6446 = N6445 & N3659;
  assign N6445 = N4228 & en_i;
  assign empty_array[554] = N6447 & N6448;
  assign N6447 = N4228 & en_i;
  assign N6448 = ~valid[554];
  assign match_array[555] = N6450 & valid[555];
  assign N6450 = N6449 & N3660;
  assign N6449 = N4228 & en_i;
  assign empty_array[555] = N6451 & N6452;
  assign N6451 = N4228 & en_i;
  assign N6452 = ~valid[555];
  assign match_array[556] = N6454 & valid[556];
  assign N6454 = N6453 & N3661;
  assign N6453 = N4228 & en_i;
  assign empty_array[556] = N6455 & N6456;
  assign N6455 = N4228 & en_i;
  assign N6456 = ~valid[556];
  assign match_array[557] = N6458 & valid[557];
  assign N6458 = N6457 & N3662;
  assign N6457 = N4228 & en_i;
  assign empty_array[557] = N6459 & N6460;
  assign N6459 = N4228 & en_i;
  assign N6460 = ~valid[557];
  assign match_array[558] = N6462 & valid[558];
  assign N6462 = N6461 & N3663;
  assign N6461 = N4228 & en_i;
  assign empty_array[558] = N6463 & N6464;
  assign N6463 = N4228 & en_i;
  assign N6464 = ~valid[558];
  assign match_array[559] = N6466 & valid[559];
  assign N6466 = N6465 & N3664;
  assign N6465 = N4228 & en_i;
  assign empty_array[559] = N6467 & N6468;
  assign N6467 = N4228 & en_i;
  assign N6468 = ~valid[559];
  assign match_array[560] = N6470 & valid[560];
  assign N6470 = N6469 & N3665;
  assign N6469 = N4228 & en_i;
  assign empty_array[560] = N6471 & N6472;
  assign N6471 = N4228 & en_i;
  assign N6472 = ~valid[560];
  assign match_array[561] = N6474 & valid[561];
  assign N6474 = N6473 & N3666;
  assign N6473 = N4228 & en_i;
  assign empty_array[561] = N6475 & N6476;
  assign N6475 = N4228 & en_i;
  assign N6476 = ~valid[561];
  assign match_array[562] = N6478 & valid[562];
  assign N6478 = N6477 & N3667;
  assign N6477 = N4228 & en_i;
  assign empty_array[562] = N6479 & N6480;
  assign N6479 = N4228 & en_i;
  assign N6480 = ~valid[562];
  assign match_array[563] = N6482 & valid[563];
  assign N6482 = N6481 & N3668;
  assign N6481 = N4228 & en_i;
  assign empty_array[563] = N6483 & N6484;
  assign N6483 = N4228 & en_i;
  assign N6484 = ~valid[563];
  assign match_array[564] = N6486 & valid[564];
  assign N6486 = N6485 & N3669;
  assign N6485 = N4228 & en_i;
  assign empty_array[564] = N6487 & N6488;
  assign N6487 = N4228 & en_i;
  assign N6488 = ~valid[564];
  assign match_array[565] = N6490 & valid[565];
  assign N6490 = N6489 & N3670;
  assign N6489 = N4228 & en_i;
  assign empty_array[565] = N6491 & N6492;
  assign N6491 = N4228 & en_i;
  assign N6492 = ~valid[565];
  assign match_array[566] = N6494 & valid[566];
  assign N6494 = N6493 & N3671;
  assign N6493 = N4228 & en_i;
  assign empty_array[566] = N6495 & N6496;
  assign N6495 = N4228 & en_i;
  assign N6496 = ~valid[566];
  assign match_array[567] = N6498 & valid[567];
  assign N6498 = N6497 & N3672;
  assign N6497 = N4228 & en_i;
  assign empty_array[567] = N6499 & N6500;
  assign N6499 = N4228 & en_i;
  assign N6500 = ~valid[567];
  assign match_array[568] = N6502 & valid[568];
  assign N6502 = N6501 & N3673;
  assign N6501 = N4228 & en_i;
  assign empty_array[568] = N6503 & N6504;
  assign N6503 = N4228 & en_i;
  assign N6504 = ~valid[568];
  assign match_array[569] = N6506 & valid[569];
  assign N6506 = N6505 & N3674;
  assign N6505 = N4228 & en_i;
  assign empty_array[569] = N6507 & N6508;
  assign N6507 = N4228 & en_i;
  assign N6508 = ~valid[569];
  assign match_array[570] = N6510 & valid[570];
  assign N6510 = N6509 & N3675;
  assign N6509 = N4228 & en_i;
  assign empty_array[570] = N6511 & N6512;
  assign N6511 = N4228 & en_i;
  assign N6512 = ~valid[570];
  assign match_array[571] = N6514 & valid[571];
  assign N6514 = N6513 & N3676;
  assign N6513 = N4228 & en_i;
  assign empty_array[571] = N6515 & N6516;
  assign N6515 = N4228 & en_i;
  assign N6516 = ~valid[571];
  assign match_array[572] = N6518 & valid[572];
  assign N6518 = N6517 & N3677;
  assign N6517 = N4228 & en_i;
  assign empty_array[572] = N6519 & N6520;
  assign N6519 = N4228 & en_i;
  assign N6520 = ~valid[572];
  assign match_array[573] = N6522 & valid[573];
  assign N6522 = N6521 & N3678;
  assign N6521 = N4228 & en_i;
  assign empty_array[573] = N6523 & N6524;
  assign N6523 = N4228 & en_i;
  assign N6524 = ~valid[573];
  assign match_array[574] = N6526 & valid[574];
  assign N6526 = N6525 & N3679;
  assign N6525 = N4228 & en_i;
  assign empty_array[574] = N6527 & N6528;
  assign N6527 = N4228 & en_i;
  assign N6528 = ~valid[574];
  assign match_array[575] = N6530 & valid[575];
  assign N6530 = N6529 & N3680;
  assign N6529 = N4228 & en_i;
  assign empty_array[575] = N6531 & N6532;
  assign N6531 = N4228 & en_i;
  assign N6532 = ~valid[575];
  assign match_array[576] = N6534 & valid[576];
  assign N6534 = N6533 & N3681;
  assign N6533 = N4228 & en_i;
  assign empty_array[576] = N6535 & N6536;
  assign N6535 = N4228 & en_i;
  assign N6536 = ~valid[576];
  assign match_array[577] = N6538 & valid[577];
  assign N6538 = N6537 & N3682;
  assign N6537 = N4228 & en_i;
  assign empty_array[577] = N6539 & N6540;
  assign N6539 = N4228 & en_i;
  assign N6540 = ~valid[577];
  assign match_array[578] = N6542 & valid[578];
  assign N6542 = N6541 & N3683;
  assign N6541 = N4228 & en_i;
  assign empty_array[578] = N6543 & N6544;
  assign N6543 = N4228 & en_i;
  assign N6544 = ~valid[578];
  assign match_array[579] = N6546 & valid[579];
  assign N6546 = N6545 & N3684;
  assign N6545 = N4228 & en_i;
  assign empty_array[579] = N6547 & N6548;
  assign N6547 = N4228 & en_i;
  assign N6548 = ~valid[579];
  assign match_array[580] = N6550 & valid[580];
  assign N6550 = N6549 & N3685;
  assign N6549 = N4228 & en_i;
  assign empty_array[580] = N6551 & N6552;
  assign N6551 = N4228 & en_i;
  assign N6552 = ~valid[580];
  assign match_array[581] = N6554 & valid[581];
  assign N6554 = N6553 & N3686;
  assign N6553 = N4228 & en_i;
  assign empty_array[581] = N6555 & N6556;
  assign N6555 = N4228 & en_i;
  assign N6556 = ~valid[581];
  assign match_array[582] = N6558 & valid[582];
  assign N6558 = N6557 & N3687;
  assign N6557 = N4228 & en_i;
  assign empty_array[582] = N6559 & N6560;
  assign N6559 = N4228 & en_i;
  assign N6560 = ~valid[582];
  assign match_array[583] = N6562 & valid[583];
  assign N6562 = N6561 & N3688;
  assign N6561 = N4228 & en_i;
  assign empty_array[583] = N6563 & N6564;
  assign N6563 = N4228 & en_i;
  assign N6564 = ~valid[583];
  assign match_array[584] = N6566 & valid[584];
  assign N6566 = N6565 & N3689;
  assign N6565 = N4228 & en_i;
  assign empty_array[584] = N6567 & N6568;
  assign N6567 = N4228 & en_i;
  assign N6568 = ~valid[584];
  assign match_array[585] = N6570 & valid[585];
  assign N6570 = N6569 & N3690;
  assign N6569 = N4228 & en_i;
  assign empty_array[585] = N6571 & N6572;
  assign N6571 = N4228 & en_i;
  assign N6572 = ~valid[585];
  assign match_array[586] = N6574 & valid[586];
  assign N6574 = N6573 & N3691;
  assign N6573 = N4228 & en_i;
  assign empty_array[586] = N6575 & N6576;
  assign N6575 = N4228 & en_i;
  assign N6576 = ~valid[586];
  assign match_array[587] = N6578 & valid[587];
  assign N6578 = N6577 & N3692;
  assign N6577 = N4228 & en_i;
  assign empty_array[587] = N6579 & N6580;
  assign N6579 = N4228 & en_i;
  assign N6580 = ~valid[587];
  assign match_array[588] = N6582 & valid[588];
  assign N6582 = N6581 & N3693;
  assign N6581 = N4228 & en_i;
  assign empty_array[588] = N6583 & N6584;
  assign N6583 = N4228 & en_i;
  assign N6584 = ~valid[588];
  assign match_array[589] = N6586 & valid[589];
  assign N6586 = N6585 & N3694;
  assign N6585 = N4228 & en_i;
  assign empty_array[589] = N6587 & N6588;
  assign N6587 = N4228 & en_i;
  assign N6588 = ~valid[589];
  assign match_array[590] = N6590 & valid[590];
  assign N6590 = N6589 & N3695;
  assign N6589 = N4228 & en_i;
  assign empty_array[590] = N6591 & N6592;
  assign N6591 = N4228 & en_i;
  assign N6592 = ~valid[590];
  assign match_array[591] = N6594 & valid[591];
  assign N6594 = N6593 & N3696;
  assign N6593 = N4228 & en_i;
  assign empty_array[591] = N6595 & N6596;
  assign N6595 = N4228 & en_i;
  assign N6596 = ~valid[591];
  assign match_array[592] = N6598 & valid[592];
  assign N6598 = N6597 & N3697;
  assign N6597 = N4228 & en_i;
  assign empty_array[592] = N6599 & N6600;
  assign N6599 = N4228 & en_i;
  assign N6600 = ~valid[592];
  assign match_array[593] = N6602 & valid[593];
  assign N6602 = N6601 & N3698;
  assign N6601 = N4228 & en_i;
  assign empty_array[593] = N6603 & N6604;
  assign N6603 = N4228 & en_i;
  assign N6604 = ~valid[593];
  assign match_array[594] = N6606 & valid[594];
  assign N6606 = N6605 & N3699;
  assign N6605 = N4228 & en_i;
  assign empty_array[594] = N6607 & N6608;
  assign N6607 = N4228 & en_i;
  assign N6608 = ~valid[594];
  assign match_array[595] = N6610 & valid[595];
  assign N6610 = N6609 & N3700;
  assign N6609 = N4228 & en_i;
  assign empty_array[595] = N6611 & N6612;
  assign N6611 = N4228 & en_i;
  assign N6612 = ~valid[595];
  assign match_array[596] = N6614 & valid[596];
  assign N6614 = N6613 & N3701;
  assign N6613 = N4228 & en_i;
  assign empty_array[596] = N6615 & N6616;
  assign N6615 = N4228 & en_i;
  assign N6616 = ~valid[596];
  assign match_array[597] = N6618 & valid[597];
  assign N6618 = N6617 & N3702;
  assign N6617 = N4228 & en_i;
  assign empty_array[597] = N6619 & N6620;
  assign N6619 = N4228 & en_i;
  assign N6620 = ~valid[597];
  assign match_array[598] = N6622 & valid[598];
  assign N6622 = N6621 & N3703;
  assign N6621 = N4228 & en_i;
  assign empty_array[598] = N6623 & N6624;
  assign N6623 = N4228 & en_i;
  assign N6624 = ~valid[598];
  assign match_array[599] = N6626 & valid[599];
  assign N6626 = N6625 & N3704;
  assign N6625 = N4228 & en_i;
  assign empty_array[599] = N6627 & N6628;
  assign N6627 = N4228 & en_i;
  assign N6628 = ~valid[599];
  assign match_array[600] = N6630 & valid[600];
  assign N6630 = N6629 & N3705;
  assign N6629 = N4228 & en_i;
  assign empty_array[600] = N6631 & N6632;
  assign N6631 = N4228 & en_i;
  assign N6632 = ~valid[600];
  assign match_array[601] = N6634 & valid[601];
  assign N6634 = N6633 & N3706;
  assign N6633 = N4228 & en_i;
  assign empty_array[601] = N6635 & N6636;
  assign N6635 = N4228 & en_i;
  assign N6636 = ~valid[601];
  assign match_array[602] = N6638 & valid[602];
  assign N6638 = N6637 & N3707;
  assign N6637 = N4228 & en_i;
  assign empty_array[602] = N6639 & N6640;
  assign N6639 = N4228 & en_i;
  assign N6640 = ~valid[602];
  assign match_array[603] = N6642 & valid[603];
  assign N6642 = N6641 & N3708;
  assign N6641 = N4228 & en_i;
  assign empty_array[603] = N6643 & N6644;
  assign N6643 = N4228 & en_i;
  assign N6644 = ~valid[603];
  assign match_array[604] = N6646 & valid[604];
  assign N6646 = N6645 & N3709;
  assign N6645 = N4228 & en_i;
  assign empty_array[604] = N6647 & N6648;
  assign N6647 = N4228 & en_i;
  assign N6648 = ~valid[604];
  assign match_array[605] = N6650 & valid[605];
  assign N6650 = N6649 & N3710;
  assign N6649 = N4228 & en_i;
  assign empty_array[605] = N6651 & N6652;
  assign N6651 = N4228 & en_i;
  assign N6652 = ~valid[605];
  assign match_array[606] = N6654 & valid[606];
  assign N6654 = N6653 & N3711;
  assign N6653 = N4228 & en_i;
  assign empty_array[606] = N6655 & N6656;
  assign N6655 = N4228 & en_i;
  assign N6656 = ~valid[606];
  assign match_array[607] = N6658 & valid[607];
  assign N6658 = N6657 & N3712;
  assign N6657 = N4228 & en_i;
  assign empty_array[607] = N6659 & N6660;
  assign N6659 = N4228 & en_i;
  assign N6660 = ~valid[607];
  assign match_array[608] = N6662 & valid[608];
  assign N6662 = N6661 & N3713;
  assign N6661 = N4228 & en_i;
  assign empty_array[608] = N6663 & N6664;
  assign N6663 = N4228 & en_i;
  assign N6664 = ~valid[608];
  assign match_array[609] = N6666 & valid[609];
  assign N6666 = N6665 & N3714;
  assign N6665 = N4228 & en_i;
  assign empty_array[609] = N6667 & N6668;
  assign N6667 = N4228 & en_i;
  assign N6668 = ~valid[609];
  assign match_array[610] = N6670 & valid[610];
  assign N6670 = N6669 & N3715;
  assign N6669 = N4228 & en_i;
  assign empty_array[610] = N6671 & N6672;
  assign N6671 = N4228 & en_i;
  assign N6672 = ~valid[610];
  assign match_array[611] = N6674 & valid[611];
  assign N6674 = N6673 & N3716;
  assign N6673 = N4228 & en_i;
  assign empty_array[611] = N6675 & N6676;
  assign N6675 = N4228 & en_i;
  assign N6676 = ~valid[611];
  assign match_array[612] = N6678 & valid[612];
  assign N6678 = N6677 & N3717;
  assign N6677 = N4228 & en_i;
  assign empty_array[612] = N6679 & N6680;
  assign N6679 = N4228 & en_i;
  assign N6680 = ~valid[612];
  assign match_array[613] = N6682 & valid[613];
  assign N6682 = N6681 & N3718;
  assign N6681 = N4228 & en_i;
  assign empty_array[613] = N6683 & N6684;
  assign N6683 = N4228 & en_i;
  assign N6684 = ~valid[613];
  assign match_array[614] = N6686 & valid[614];
  assign N6686 = N6685 & N3719;
  assign N6685 = N4228 & en_i;
  assign empty_array[614] = N6687 & N6688;
  assign N6687 = N4228 & en_i;
  assign N6688 = ~valid[614];
  assign match_array[615] = N6690 & valid[615];
  assign N6690 = N6689 & N3720;
  assign N6689 = N4228 & en_i;
  assign empty_array[615] = N6691 & N6692;
  assign N6691 = N4228 & en_i;
  assign N6692 = ~valid[615];
  assign match_array[616] = N6694 & valid[616];
  assign N6694 = N6693 & N3721;
  assign N6693 = N4228 & en_i;
  assign empty_array[616] = N6695 & N6696;
  assign N6695 = N4228 & en_i;
  assign N6696 = ~valid[616];
  assign match_array[617] = N6698 & valid[617];
  assign N6698 = N6697 & N3722;
  assign N6697 = N4228 & en_i;
  assign empty_array[617] = N6699 & N6700;
  assign N6699 = N4228 & en_i;
  assign N6700 = ~valid[617];
  assign match_array[618] = N6702 & valid[618];
  assign N6702 = N6701 & N3723;
  assign N6701 = N4228 & en_i;
  assign empty_array[618] = N6703 & N6704;
  assign N6703 = N4228 & en_i;
  assign N6704 = ~valid[618];
  assign match_array[619] = N6706 & valid[619];
  assign N6706 = N6705 & N3724;
  assign N6705 = N4228 & en_i;
  assign empty_array[619] = N6707 & N6708;
  assign N6707 = N4228 & en_i;
  assign N6708 = ~valid[619];
  assign match_array[620] = N6710 & valid[620];
  assign N6710 = N6709 & N3725;
  assign N6709 = N4228 & en_i;
  assign empty_array[620] = N6711 & N6712;
  assign N6711 = N4228 & en_i;
  assign N6712 = ~valid[620];
  assign match_array[621] = N6714 & valid[621];
  assign N6714 = N6713 & N3726;
  assign N6713 = N4228 & en_i;
  assign empty_array[621] = N6715 & N6716;
  assign N6715 = N4228 & en_i;
  assign N6716 = ~valid[621];
  assign match_array[622] = N6718 & valid[622];
  assign N6718 = N6717 & N3727;
  assign N6717 = N4228 & en_i;
  assign empty_array[622] = N6719 & N6720;
  assign N6719 = N4228 & en_i;
  assign N6720 = ~valid[622];
  assign match_array[623] = N6722 & valid[623];
  assign N6722 = N6721 & N3728;
  assign N6721 = N4228 & en_i;
  assign empty_array[623] = N6723 & N6724;
  assign N6723 = N4228 & en_i;
  assign N6724 = ~valid[623];
  assign match_array[624] = N6726 & valid[624];
  assign N6726 = N6725 & N3729;
  assign N6725 = N4228 & en_i;
  assign empty_array[624] = N6727 & N6728;
  assign N6727 = N4228 & en_i;
  assign N6728 = ~valid[624];
  assign match_array[625] = N6730 & valid[625];
  assign N6730 = N6729 & N3730;
  assign N6729 = N4228 & en_i;
  assign empty_array[625] = N6731 & N6732;
  assign N6731 = N4228 & en_i;
  assign N6732 = ~valid[625];
  assign match_array[626] = N6734 & valid[626];
  assign N6734 = N6733 & N3731;
  assign N6733 = N4228 & en_i;
  assign empty_array[626] = N6735 & N6736;
  assign N6735 = N4228 & en_i;
  assign N6736 = ~valid[626];
  assign match_array[627] = N6738 & valid[627];
  assign N6738 = N6737 & N3732;
  assign N6737 = N4228 & en_i;
  assign empty_array[627] = N6739 & N6740;
  assign N6739 = N4228 & en_i;
  assign N6740 = ~valid[627];
  assign match_array[628] = N6742 & valid[628];
  assign N6742 = N6741 & N3733;
  assign N6741 = N4228 & en_i;
  assign empty_array[628] = N6743 & N6744;
  assign N6743 = N4228 & en_i;
  assign N6744 = ~valid[628];
  assign match_array[629] = N6746 & valid[629];
  assign N6746 = N6745 & N3734;
  assign N6745 = N4228 & en_i;
  assign empty_array[629] = N6747 & N6748;
  assign N6747 = N4228 & en_i;
  assign N6748 = ~valid[629];
  assign match_array[630] = N6750 & valid[630];
  assign N6750 = N6749 & N3735;
  assign N6749 = N4228 & en_i;
  assign empty_array[630] = N6751 & N6752;
  assign N6751 = N4228 & en_i;
  assign N6752 = ~valid[630];
  assign match_array[631] = N6754 & valid[631];
  assign N6754 = N6753 & N3736;
  assign N6753 = N4228 & en_i;
  assign empty_array[631] = N6755 & N6756;
  assign N6755 = N4228 & en_i;
  assign N6756 = ~valid[631];
  assign match_array[632] = N6758 & valid[632];
  assign N6758 = N6757 & N3737;
  assign N6757 = N4228 & en_i;
  assign empty_array[632] = N6759 & N6760;
  assign N6759 = N4228 & en_i;
  assign N6760 = ~valid[632];
  assign match_array[633] = N6762 & valid[633];
  assign N6762 = N6761 & N3738;
  assign N6761 = N4228 & en_i;
  assign empty_array[633] = N6763 & N6764;
  assign N6763 = N4228 & en_i;
  assign N6764 = ~valid[633];
  assign match_array[634] = N6766 & valid[634];
  assign N6766 = N6765 & N3739;
  assign N6765 = N4228 & en_i;
  assign empty_array[634] = N6767 & N6768;
  assign N6767 = N4228 & en_i;
  assign N6768 = ~valid[634];
  assign match_array[635] = N6770 & valid[635];
  assign N6770 = N6769 & N3740;
  assign N6769 = N4228 & en_i;
  assign empty_array[635] = N6771 & N6772;
  assign N6771 = N4228 & en_i;
  assign N6772 = ~valid[635];
  assign match_array[636] = N6774 & valid[636];
  assign N6774 = N6773 & N3741;
  assign N6773 = N4228 & en_i;
  assign empty_array[636] = N6775 & N6776;
  assign N6775 = N4228 & en_i;
  assign N6776 = ~valid[636];
  assign match_array[637] = N6778 & valid[637];
  assign N6778 = N6777 & N3742;
  assign N6777 = N4228 & en_i;
  assign empty_array[637] = N6779 & N6780;
  assign N6779 = N4228 & en_i;
  assign N6780 = ~valid[637];
  assign match_array[638] = N6782 & valid[638];
  assign N6782 = N6781 & N3743;
  assign N6781 = N4228 & en_i;
  assign empty_array[638] = N6783 & N6784;
  assign N6783 = N4228 & en_i;
  assign N6784 = ~valid[638];
  assign match_array[639] = N6786 & valid[639];
  assign N6786 = N6785 & N3744;
  assign N6785 = N4228 & en_i;
  assign empty_array[639] = N6787 & N6788;
  assign N6787 = N4228 & en_i;
  assign N6788 = ~valid[639];
  assign match_array[640] = N6790 & valid[640];
  assign N6790 = N6789 & N3745;
  assign N6789 = N4228 & en_i;
  assign empty_array[640] = N6791 & N6792;
  assign N6791 = N4228 & en_i;
  assign N6792 = ~valid[640];
  assign match_array[641] = N6794 & valid[641];
  assign N6794 = N6793 & N3746;
  assign N6793 = N4228 & en_i;
  assign empty_array[641] = N6795 & N6796;
  assign N6795 = N4228 & en_i;
  assign N6796 = ~valid[641];
  assign match_array[642] = N6798 & valid[642];
  assign N6798 = N6797 & N3747;
  assign N6797 = N4228 & en_i;
  assign empty_array[642] = N6799 & N6800;
  assign N6799 = N4228 & en_i;
  assign N6800 = ~valid[642];
  assign match_array[643] = N6802 & valid[643];
  assign N6802 = N6801 & N3748;
  assign N6801 = N4228 & en_i;
  assign empty_array[643] = N6803 & N6804;
  assign N6803 = N4228 & en_i;
  assign N6804 = ~valid[643];
  assign match_array[644] = N6806 & valid[644];
  assign N6806 = N6805 & N3749;
  assign N6805 = N4228 & en_i;
  assign empty_array[644] = N6807 & N6808;
  assign N6807 = N4228 & en_i;
  assign N6808 = ~valid[644];
  assign match_array[645] = N6810 & valid[645];
  assign N6810 = N6809 & N3750;
  assign N6809 = N4228 & en_i;
  assign empty_array[645] = N6811 & N6812;
  assign N6811 = N4228 & en_i;
  assign N6812 = ~valid[645];
  assign match_array[646] = N6814 & valid[646];
  assign N6814 = N6813 & N3751;
  assign N6813 = N4228 & en_i;
  assign empty_array[646] = N6815 & N6816;
  assign N6815 = N4228 & en_i;
  assign N6816 = ~valid[646];
  assign match_array[647] = N6818 & valid[647];
  assign N6818 = N6817 & N3752;
  assign N6817 = N4228 & en_i;
  assign empty_array[647] = N6819 & N6820;
  assign N6819 = N4228 & en_i;
  assign N6820 = ~valid[647];
  assign match_array[648] = N6822 & valid[648];
  assign N6822 = N6821 & N3753;
  assign N6821 = N4228 & en_i;
  assign empty_array[648] = N6823 & N6824;
  assign N6823 = N4228 & en_i;
  assign N6824 = ~valid[648];
  assign match_array[649] = N6826 & valid[649];
  assign N6826 = N6825 & N3754;
  assign N6825 = N4228 & en_i;
  assign empty_array[649] = N6827 & N6828;
  assign N6827 = N4228 & en_i;
  assign N6828 = ~valid[649];
  assign match_array[650] = N6830 & valid[650];
  assign N6830 = N6829 & N3755;
  assign N6829 = N4228 & en_i;
  assign empty_array[650] = N6831 & N6832;
  assign N6831 = N4228 & en_i;
  assign N6832 = ~valid[650];
  assign match_array[651] = N6834 & valid[651];
  assign N6834 = N6833 & N3756;
  assign N6833 = N4228 & en_i;
  assign empty_array[651] = N6835 & N6836;
  assign N6835 = N4228 & en_i;
  assign N6836 = ~valid[651];
  assign match_array[652] = N6838 & valid[652];
  assign N6838 = N6837 & N3757;
  assign N6837 = N4228 & en_i;
  assign empty_array[652] = N6839 & N6840;
  assign N6839 = N4228 & en_i;
  assign N6840 = ~valid[652];
  assign match_array[653] = N6842 & valid[653];
  assign N6842 = N6841 & N3758;
  assign N6841 = N4228 & en_i;
  assign empty_array[653] = N6843 & N6844;
  assign N6843 = N4228 & en_i;
  assign N6844 = ~valid[653];
  assign match_array[654] = N6846 & valid[654];
  assign N6846 = N6845 & N3759;
  assign N6845 = N4228 & en_i;
  assign empty_array[654] = N6847 & N6848;
  assign N6847 = N4228 & en_i;
  assign N6848 = ~valid[654];
  assign match_array[655] = N6850 & valid[655];
  assign N6850 = N6849 & N3760;
  assign N6849 = N4228 & en_i;
  assign empty_array[655] = N6851 & N6852;
  assign N6851 = N4228 & en_i;
  assign N6852 = ~valid[655];
  assign match_array[656] = N6854 & valid[656];
  assign N6854 = N6853 & N3761;
  assign N6853 = N4228 & en_i;
  assign empty_array[656] = N6855 & N6856;
  assign N6855 = N4228 & en_i;
  assign N6856 = ~valid[656];
  assign match_array[657] = N6858 & valid[657];
  assign N6858 = N6857 & N3762;
  assign N6857 = N4228 & en_i;
  assign empty_array[657] = N6859 & N6860;
  assign N6859 = N4228 & en_i;
  assign N6860 = ~valid[657];
  assign match_array[658] = N6862 & valid[658];
  assign N6862 = N6861 & N3763;
  assign N6861 = N4228 & en_i;
  assign empty_array[658] = N6863 & N6864;
  assign N6863 = N4228 & en_i;
  assign N6864 = ~valid[658];
  assign match_array[659] = N6866 & valid[659];
  assign N6866 = N6865 & N3764;
  assign N6865 = N4228 & en_i;
  assign empty_array[659] = N6867 & N6868;
  assign N6867 = N4228 & en_i;
  assign N6868 = ~valid[659];
  assign match_array[660] = N6870 & valid[660];
  assign N6870 = N6869 & N3765;
  assign N6869 = N4228 & en_i;
  assign empty_array[660] = N6871 & N6872;
  assign N6871 = N4228 & en_i;
  assign N6872 = ~valid[660];
  assign match_array[661] = N6874 & valid[661];
  assign N6874 = N6873 & N3766;
  assign N6873 = N4228 & en_i;
  assign empty_array[661] = N6875 & N6876;
  assign N6875 = N4228 & en_i;
  assign N6876 = ~valid[661];
  assign match_array[662] = N6878 & valid[662];
  assign N6878 = N6877 & N3767;
  assign N6877 = N4228 & en_i;
  assign empty_array[662] = N6879 & N6880;
  assign N6879 = N4228 & en_i;
  assign N6880 = ~valid[662];
  assign match_array[663] = N6882 & valid[663];
  assign N6882 = N6881 & N3768;
  assign N6881 = N4228 & en_i;
  assign empty_array[663] = N6883 & N6884;
  assign N6883 = N4228 & en_i;
  assign N6884 = ~valid[663];
  assign match_array[664] = N6886 & valid[664];
  assign N6886 = N6885 & N3769;
  assign N6885 = N4228 & en_i;
  assign empty_array[664] = N6887 & N6888;
  assign N6887 = N4228 & en_i;
  assign N6888 = ~valid[664];
  assign match_array[665] = N6890 & valid[665];
  assign N6890 = N6889 & N3770;
  assign N6889 = N4228 & en_i;
  assign empty_array[665] = N6891 & N6892;
  assign N6891 = N4228 & en_i;
  assign N6892 = ~valid[665];
  assign match_array[666] = N6894 & valid[666];
  assign N6894 = N6893 & N3771;
  assign N6893 = N4228 & en_i;
  assign empty_array[666] = N6895 & N6896;
  assign N6895 = N4228 & en_i;
  assign N6896 = ~valid[666];
  assign match_array[667] = N6898 & valid[667];
  assign N6898 = N6897 & N3772;
  assign N6897 = N4228 & en_i;
  assign empty_array[667] = N6899 & N6900;
  assign N6899 = N4228 & en_i;
  assign N6900 = ~valid[667];
  assign match_array[668] = N6902 & valid[668];
  assign N6902 = N6901 & N3773;
  assign N6901 = N4228 & en_i;
  assign empty_array[668] = N6903 & N6904;
  assign N6903 = N4228 & en_i;
  assign N6904 = ~valid[668];
  assign match_array[669] = N6906 & valid[669];
  assign N6906 = N6905 & N3774;
  assign N6905 = N4228 & en_i;
  assign empty_array[669] = N6907 & N6908;
  assign N6907 = N4228 & en_i;
  assign N6908 = ~valid[669];
  assign match_array[670] = N6910 & valid[670];
  assign N6910 = N6909 & N3775;
  assign N6909 = N4228 & en_i;
  assign empty_array[670] = N6911 & N6912;
  assign N6911 = N4228 & en_i;
  assign N6912 = ~valid[670];
  assign match_array[671] = N6914 & valid[671];
  assign N6914 = N6913 & N3776;
  assign N6913 = N4228 & en_i;
  assign empty_array[671] = N6915 & N6916;
  assign N6915 = N4228 & en_i;
  assign N6916 = ~valid[671];
  assign match_array[672] = N6918 & valid[672];
  assign N6918 = N6917 & N3777;
  assign N6917 = N4228 & en_i;
  assign empty_array[672] = N6919 & N6920;
  assign N6919 = N4228 & en_i;
  assign N6920 = ~valid[672];
  assign match_array[673] = N6922 & valid[673];
  assign N6922 = N6921 & N3778;
  assign N6921 = N4228 & en_i;
  assign empty_array[673] = N6923 & N6924;
  assign N6923 = N4228 & en_i;
  assign N6924 = ~valid[673];
  assign match_array[674] = N6926 & valid[674];
  assign N6926 = N6925 & N3779;
  assign N6925 = N4228 & en_i;
  assign empty_array[674] = N6927 & N6928;
  assign N6927 = N4228 & en_i;
  assign N6928 = ~valid[674];
  assign match_array[675] = N6930 & valid[675];
  assign N6930 = N6929 & N3780;
  assign N6929 = N4228 & en_i;
  assign empty_array[675] = N6931 & N6932;
  assign N6931 = N4228 & en_i;
  assign N6932 = ~valid[675];
  assign match_array[676] = N6934 & valid[676];
  assign N6934 = N6933 & N3781;
  assign N6933 = N4228 & en_i;
  assign empty_array[676] = N6935 & N6936;
  assign N6935 = N4228 & en_i;
  assign N6936 = ~valid[676];
  assign match_array[677] = N6938 & valid[677];
  assign N6938 = N6937 & N3782;
  assign N6937 = N4228 & en_i;
  assign empty_array[677] = N6939 & N6940;
  assign N6939 = N4228 & en_i;
  assign N6940 = ~valid[677];
  assign match_array[678] = N6942 & valid[678];
  assign N6942 = N6941 & N3783;
  assign N6941 = N4228 & en_i;
  assign empty_array[678] = N6943 & N6944;
  assign N6943 = N4228 & en_i;
  assign N6944 = ~valid[678];
  assign match_array[679] = N6946 & valid[679];
  assign N6946 = N6945 & N3784;
  assign N6945 = N4228 & en_i;
  assign empty_array[679] = N6947 & N6948;
  assign N6947 = N4228 & en_i;
  assign N6948 = ~valid[679];
  assign match_array[680] = N6950 & valid[680];
  assign N6950 = N6949 & N3785;
  assign N6949 = N4228 & en_i;
  assign empty_array[680] = N6951 & N6952;
  assign N6951 = N4228 & en_i;
  assign N6952 = ~valid[680];
  assign match_array[681] = N6954 & valid[681];
  assign N6954 = N6953 & N3786;
  assign N6953 = N4228 & en_i;
  assign empty_array[681] = N6955 & N6956;
  assign N6955 = N4228 & en_i;
  assign N6956 = ~valid[681];
  assign match_array[682] = N6958 & valid[682];
  assign N6958 = N6957 & N3787;
  assign N6957 = N4228 & en_i;
  assign empty_array[682] = N6959 & N6960;
  assign N6959 = N4228 & en_i;
  assign N6960 = ~valid[682];
  assign match_array[683] = N6962 & valid[683];
  assign N6962 = N6961 & N3788;
  assign N6961 = N4228 & en_i;
  assign empty_array[683] = N6963 & N6964;
  assign N6963 = N4228 & en_i;
  assign N6964 = ~valid[683];
  assign match_array[684] = N6966 & valid[684];
  assign N6966 = N6965 & N3789;
  assign N6965 = N4228 & en_i;
  assign empty_array[684] = N6967 & N6968;
  assign N6967 = N4228 & en_i;
  assign N6968 = ~valid[684];
  assign match_array[685] = N6970 & valid[685];
  assign N6970 = N6969 & N3790;
  assign N6969 = N4228 & en_i;
  assign empty_array[685] = N6971 & N6972;
  assign N6971 = N4228 & en_i;
  assign N6972 = ~valid[685];
  assign match_array[686] = N6974 & valid[686];
  assign N6974 = N6973 & N3791;
  assign N6973 = N4228 & en_i;
  assign empty_array[686] = N6975 & N6976;
  assign N6975 = N4228 & en_i;
  assign N6976 = ~valid[686];
  assign match_array[687] = N6978 & valid[687];
  assign N6978 = N6977 & N3792;
  assign N6977 = N4228 & en_i;
  assign empty_array[687] = N6979 & N6980;
  assign N6979 = N4228 & en_i;
  assign N6980 = ~valid[687];
  assign match_array[688] = N6982 & valid[688];
  assign N6982 = N6981 & N3793;
  assign N6981 = N4228 & en_i;
  assign empty_array[688] = N6983 & N6984;
  assign N6983 = N4228 & en_i;
  assign N6984 = ~valid[688];
  assign match_array[689] = N6986 & valid[689];
  assign N6986 = N6985 & N3794;
  assign N6985 = N4228 & en_i;
  assign empty_array[689] = N6987 & N6988;
  assign N6987 = N4228 & en_i;
  assign N6988 = ~valid[689];
  assign match_array[690] = N6990 & valid[690];
  assign N6990 = N6989 & N3795;
  assign N6989 = N4228 & en_i;
  assign empty_array[690] = N6991 & N6992;
  assign N6991 = N4228 & en_i;
  assign N6992 = ~valid[690];
  assign match_array[691] = N6994 & valid[691];
  assign N6994 = N6993 & N3796;
  assign N6993 = N4228 & en_i;
  assign empty_array[691] = N6995 & N6996;
  assign N6995 = N4228 & en_i;
  assign N6996 = ~valid[691];
  assign match_array[692] = N6998 & valid[692];
  assign N6998 = N6997 & N3797;
  assign N6997 = N4228 & en_i;
  assign empty_array[692] = N6999 & N7000;
  assign N6999 = N4228 & en_i;
  assign N7000 = ~valid[692];
  assign match_array[693] = N7002 & valid[693];
  assign N7002 = N7001 & N3798;
  assign N7001 = N4228 & en_i;
  assign empty_array[693] = N7003 & N7004;
  assign N7003 = N4228 & en_i;
  assign N7004 = ~valid[693];
  assign match_array[694] = N7006 & valid[694];
  assign N7006 = N7005 & N3799;
  assign N7005 = N4228 & en_i;
  assign empty_array[694] = N7007 & N7008;
  assign N7007 = N4228 & en_i;
  assign N7008 = ~valid[694];
  assign match_array[695] = N7010 & valid[695];
  assign N7010 = N7009 & N3800;
  assign N7009 = N4228 & en_i;
  assign empty_array[695] = N7011 & N7012;
  assign N7011 = N4228 & en_i;
  assign N7012 = ~valid[695];
  assign match_array[696] = N7014 & valid[696];
  assign N7014 = N7013 & N3801;
  assign N7013 = N4228 & en_i;
  assign empty_array[696] = N7015 & N7016;
  assign N7015 = N4228 & en_i;
  assign N7016 = ~valid[696];
  assign match_array[697] = N7018 & valid[697];
  assign N7018 = N7017 & N3802;
  assign N7017 = N4228 & en_i;
  assign empty_array[697] = N7019 & N7020;
  assign N7019 = N4228 & en_i;
  assign N7020 = ~valid[697];
  assign match_array[698] = N7022 & valid[698];
  assign N7022 = N7021 & N3803;
  assign N7021 = N4228 & en_i;
  assign empty_array[698] = N7023 & N7024;
  assign N7023 = N4228 & en_i;
  assign N7024 = ~valid[698];
  assign match_array[699] = N7026 & valid[699];
  assign N7026 = N7025 & N3804;
  assign N7025 = N4228 & en_i;
  assign empty_array[699] = N7027 & N7028;
  assign N7027 = N4228 & en_i;
  assign N7028 = ~valid[699];
  assign match_array[700] = N7030 & valid[700];
  assign N7030 = N7029 & N3805;
  assign N7029 = N4228 & en_i;
  assign empty_array[700] = N7031 & N7032;
  assign N7031 = N4228 & en_i;
  assign N7032 = ~valid[700];
  assign match_array[701] = N7034 & valid[701];
  assign N7034 = N7033 & N3806;
  assign N7033 = N4228 & en_i;
  assign empty_array[701] = N7035 & N7036;
  assign N7035 = N4228 & en_i;
  assign N7036 = ~valid[701];
  assign match_array[702] = N7038 & valid[702];
  assign N7038 = N7037 & N3807;
  assign N7037 = N4228 & en_i;
  assign empty_array[702] = N7039 & N7040;
  assign N7039 = N4228 & en_i;
  assign N7040 = ~valid[702];
  assign match_array[703] = N7042 & valid[703];
  assign N7042 = N7041 & N3808;
  assign N7041 = N4228 & en_i;
  assign empty_array[703] = N7043 & N7044;
  assign N7043 = N4228 & en_i;
  assign N7044 = ~valid[703];
  assign match_array[704] = N7046 & valid[704];
  assign N7046 = N7045 & N3809;
  assign N7045 = N4228 & en_i;
  assign empty_array[704] = N7047 & N7048;
  assign N7047 = N4228 & en_i;
  assign N7048 = ~valid[704];
  assign match_array[705] = N7050 & valid[705];
  assign N7050 = N7049 & N3810;
  assign N7049 = N4228 & en_i;
  assign empty_array[705] = N7051 & N7052;
  assign N7051 = N4228 & en_i;
  assign N7052 = ~valid[705];
  assign match_array[706] = N7054 & valid[706];
  assign N7054 = N7053 & N3811;
  assign N7053 = N4228 & en_i;
  assign empty_array[706] = N7055 & N7056;
  assign N7055 = N4228 & en_i;
  assign N7056 = ~valid[706];
  assign match_array[707] = N7058 & valid[707];
  assign N7058 = N7057 & N3812;
  assign N7057 = N4228 & en_i;
  assign empty_array[707] = N7059 & N7060;
  assign N7059 = N4228 & en_i;
  assign N7060 = ~valid[707];
  assign match_array[708] = N7062 & valid[708];
  assign N7062 = N7061 & N3813;
  assign N7061 = N4228 & en_i;
  assign empty_array[708] = N7063 & N7064;
  assign N7063 = N4228 & en_i;
  assign N7064 = ~valid[708];
  assign match_array[709] = N7066 & valid[709];
  assign N7066 = N7065 & N3814;
  assign N7065 = N4228 & en_i;
  assign empty_array[709] = N7067 & N7068;
  assign N7067 = N4228 & en_i;
  assign N7068 = ~valid[709];
  assign match_array[710] = N7070 & valid[710];
  assign N7070 = N7069 & N3815;
  assign N7069 = N4228 & en_i;
  assign empty_array[710] = N7071 & N7072;
  assign N7071 = N4228 & en_i;
  assign N7072 = ~valid[710];
  assign match_array[711] = N7074 & valid[711];
  assign N7074 = N7073 & N3816;
  assign N7073 = N4228 & en_i;
  assign empty_array[711] = N7075 & N7076;
  assign N7075 = N4228 & en_i;
  assign N7076 = ~valid[711];
  assign match_array[712] = N7078 & valid[712];
  assign N7078 = N7077 & N3817;
  assign N7077 = N4228 & en_i;
  assign empty_array[712] = N7079 & N7080;
  assign N7079 = N4228 & en_i;
  assign N7080 = ~valid[712];
  assign match_array[713] = N7082 & valid[713];
  assign N7082 = N7081 & N3818;
  assign N7081 = N4228 & en_i;
  assign empty_array[713] = N7083 & N7084;
  assign N7083 = N4228 & en_i;
  assign N7084 = ~valid[713];
  assign match_array[714] = N7086 & valid[714];
  assign N7086 = N7085 & N3819;
  assign N7085 = N4228 & en_i;
  assign empty_array[714] = N7087 & N7088;
  assign N7087 = N4228 & en_i;
  assign N7088 = ~valid[714];
  assign match_array[715] = N7090 & valid[715];
  assign N7090 = N7089 & N3820;
  assign N7089 = N4228 & en_i;
  assign empty_array[715] = N7091 & N7092;
  assign N7091 = N4228 & en_i;
  assign N7092 = ~valid[715];
  assign match_array[716] = N7094 & valid[716];
  assign N7094 = N7093 & N3821;
  assign N7093 = N4228 & en_i;
  assign empty_array[716] = N7095 & N7096;
  assign N7095 = N4228 & en_i;
  assign N7096 = ~valid[716];
  assign match_array[717] = N7098 & valid[717];
  assign N7098 = N7097 & N3822;
  assign N7097 = N4228 & en_i;
  assign empty_array[717] = N7099 & N7100;
  assign N7099 = N4228 & en_i;
  assign N7100 = ~valid[717];
  assign match_array[718] = N7102 & valid[718];
  assign N7102 = N7101 & N3823;
  assign N7101 = N4228 & en_i;
  assign empty_array[718] = N7103 & N7104;
  assign N7103 = N4228 & en_i;
  assign N7104 = ~valid[718];
  assign match_array[719] = N7106 & valid[719];
  assign N7106 = N7105 & N3824;
  assign N7105 = N4228 & en_i;
  assign empty_array[719] = N7107 & N7108;
  assign N7107 = N4228 & en_i;
  assign N7108 = ~valid[719];
  assign match_array[720] = N7110 & valid[720];
  assign N7110 = N7109 & N3825;
  assign N7109 = N4228 & en_i;
  assign empty_array[720] = N7111 & N7112;
  assign N7111 = N4228 & en_i;
  assign N7112 = ~valid[720];
  assign match_array[721] = N7114 & valid[721];
  assign N7114 = N7113 & N3826;
  assign N7113 = N4228 & en_i;
  assign empty_array[721] = N7115 & N7116;
  assign N7115 = N4228 & en_i;
  assign N7116 = ~valid[721];
  assign match_array[722] = N7118 & valid[722];
  assign N7118 = N7117 & N3827;
  assign N7117 = N4228 & en_i;
  assign empty_array[722] = N7119 & N7120;
  assign N7119 = N4228 & en_i;
  assign N7120 = ~valid[722];
  assign match_array[723] = N7122 & valid[723];
  assign N7122 = N7121 & N3828;
  assign N7121 = N4228 & en_i;
  assign empty_array[723] = N7123 & N7124;
  assign N7123 = N4228 & en_i;
  assign N7124 = ~valid[723];
  assign match_array[724] = N7126 & valid[724];
  assign N7126 = N7125 & N3829;
  assign N7125 = N4228 & en_i;
  assign empty_array[724] = N7127 & N7128;
  assign N7127 = N4228 & en_i;
  assign N7128 = ~valid[724];
  assign match_array[725] = N7130 & valid[725];
  assign N7130 = N7129 & N3830;
  assign N7129 = N4228 & en_i;
  assign empty_array[725] = N7131 & N7132;
  assign N7131 = N4228 & en_i;
  assign N7132 = ~valid[725];
  assign match_array[726] = N7134 & valid[726];
  assign N7134 = N7133 & N3831;
  assign N7133 = N4228 & en_i;
  assign empty_array[726] = N7135 & N7136;
  assign N7135 = N4228 & en_i;
  assign N7136 = ~valid[726];
  assign match_array[727] = N7138 & valid[727];
  assign N7138 = N7137 & N3832;
  assign N7137 = N4228 & en_i;
  assign empty_array[727] = N7139 & N7140;
  assign N7139 = N4228 & en_i;
  assign N7140 = ~valid[727];
  assign match_array[728] = N7142 & valid[728];
  assign N7142 = N7141 & N3833;
  assign N7141 = N4228 & en_i;
  assign empty_array[728] = N7143 & N7144;
  assign N7143 = N4228 & en_i;
  assign N7144 = ~valid[728];
  assign match_array[729] = N7146 & valid[729];
  assign N7146 = N7145 & N3834;
  assign N7145 = N4228 & en_i;
  assign empty_array[729] = N7147 & N7148;
  assign N7147 = N4228 & en_i;
  assign N7148 = ~valid[729];
  assign match_array[730] = N7150 & valid[730];
  assign N7150 = N7149 & N3835;
  assign N7149 = N4228 & en_i;
  assign empty_array[730] = N7151 & N7152;
  assign N7151 = N4228 & en_i;
  assign N7152 = ~valid[730];
  assign match_array[731] = N7154 & valid[731];
  assign N7154 = N7153 & N3836;
  assign N7153 = N4228 & en_i;
  assign empty_array[731] = N7155 & N7156;
  assign N7155 = N4228 & en_i;
  assign N7156 = ~valid[731];
  assign match_array[732] = N7158 & valid[732];
  assign N7158 = N7157 & N3837;
  assign N7157 = N4228 & en_i;
  assign empty_array[732] = N7159 & N7160;
  assign N7159 = N4228 & en_i;
  assign N7160 = ~valid[732];
  assign match_array[733] = N7162 & valid[733];
  assign N7162 = N7161 & N3838;
  assign N7161 = N4228 & en_i;
  assign empty_array[733] = N7163 & N7164;
  assign N7163 = N4228 & en_i;
  assign N7164 = ~valid[733];
  assign match_array[734] = N7166 & valid[734];
  assign N7166 = N7165 & N3839;
  assign N7165 = N4228 & en_i;
  assign empty_array[734] = N7167 & N7168;
  assign N7167 = N4228 & en_i;
  assign N7168 = ~valid[734];
  assign match_array[735] = N7170 & valid[735];
  assign N7170 = N7169 & N3840;
  assign N7169 = N4228 & en_i;
  assign empty_array[735] = N7171 & N7172;
  assign N7171 = N4228 & en_i;
  assign N7172 = ~valid[735];
  assign match_array[736] = N7174 & valid[736];
  assign N7174 = N7173 & N3841;
  assign N7173 = N4228 & en_i;
  assign empty_array[736] = N7175 & N7176;
  assign N7175 = N4228 & en_i;
  assign N7176 = ~valid[736];
  assign match_array[737] = N7178 & valid[737];
  assign N7178 = N7177 & N3842;
  assign N7177 = N4228 & en_i;
  assign empty_array[737] = N7179 & N7180;
  assign N7179 = N4228 & en_i;
  assign N7180 = ~valid[737];
  assign match_array[738] = N7182 & valid[738];
  assign N7182 = N7181 & N3843;
  assign N7181 = N4228 & en_i;
  assign empty_array[738] = N7183 & N7184;
  assign N7183 = N4228 & en_i;
  assign N7184 = ~valid[738];
  assign match_array[739] = N7186 & valid[739];
  assign N7186 = N7185 & N3844;
  assign N7185 = N4228 & en_i;
  assign empty_array[739] = N7187 & N7188;
  assign N7187 = N4228 & en_i;
  assign N7188 = ~valid[739];
  assign match_array[740] = N7190 & valid[740];
  assign N7190 = N7189 & N3845;
  assign N7189 = N4228 & en_i;
  assign empty_array[740] = N7191 & N7192;
  assign N7191 = N4228 & en_i;
  assign N7192 = ~valid[740];
  assign match_array[741] = N7194 & valid[741];
  assign N7194 = N7193 & N3846;
  assign N7193 = N4228 & en_i;
  assign empty_array[741] = N7195 & N7196;
  assign N7195 = N4228 & en_i;
  assign N7196 = ~valid[741];
  assign match_array[742] = N7198 & valid[742];
  assign N7198 = N7197 & N3847;
  assign N7197 = N4228 & en_i;
  assign empty_array[742] = N7199 & N7200;
  assign N7199 = N4228 & en_i;
  assign N7200 = ~valid[742];
  assign match_array[743] = N7202 & valid[743];
  assign N7202 = N7201 & N3848;
  assign N7201 = N4228 & en_i;
  assign empty_array[743] = N7203 & N7204;
  assign N7203 = N4228 & en_i;
  assign N7204 = ~valid[743];
  assign match_array[744] = N7206 & valid[744];
  assign N7206 = N7205 & N3849;
  assign N7205 = N4228 & en_i;
  assign empty_array[744] = N7207 & N7208;
  assign N7207 = N4228 & en_i;
  assign N7208 = ~valid[744];
  assign match_array[745] = N7210 & valid[745];
  assign N7210 = N7209 & N3850;
  assign N7209 = N4228 & en_i;
  assign empty_array[745] = N7211 & N7212;
  assign N7211 = N4228 & en_i;
  assign N7212 = ~valid[745];
  assign match_array[746] = N7214 & valid[746];
  assign N7214 = N7213 & N3851;
  assign N7213 = N4228 & en_i;
  assign empty_array[746] = N7215 & N7216;
  assign N7215 = N4228 & en_i;
  assign N7216 = ~valid[746];
  assign match_array[747] = N7218 & valid[747];
  assign N7218 = N7217 & N3852;
  assign N7217 = N4228 & en_i;
  assign empty_array[747] = N7219 & N7220;
  assign N7219 = N4228 & en_i;
  assign N7220 = ~valid[747];
  assign match_array[748] = N7222 & valid[748];
  assign N7222 = N7221 & N3853;
  assign N7221 = N4228 & en_i;
  assign empty_array[748] = N7223 & N7224;
  assign N7223 = N4228 & en_i;
  assign N7224 = ~valid[748];
  assign match_array[749] = N7226 & valid[749];
  assign N7226 = N7225 & N3854;
  assign N7225 = N4228 & en_i;
  assign empty_array[749] = N7227 & N7228;
  assign N7227 = N4228 & en_i;
  assign N7228 = ~valid[749];
  assign match_array[750] = N7230 & valid[750];
  assign N7230 = N7229 & N3855;
  assign N7229 = N4228 & en_i;
  assign empty_array[750] = N7231 & N7232;
  assign N7231 = N4228 & en_i;
  assign N7232 = ~valid[750];
  assign match_array[751] = N7234 & valid[751];
  assign N7234 = N7233 & N3856;
  assign N7233 = N4228 & en_i;
  assign empty_array[751] = N7235 & N7236;
  assign N7235 = N4228 & en_i;
  assign N7236 = ~valid[751];
  assign match_array[752] = N7238 & valid[752];
  assign N7238 = N7237 & N3857;
  assign N7237 = N4228 & en_i;
  assign empty_array[752] = N7239 & N7240;
  assign N7239 = N4228 & en_i;
  assign N7240 = ~valid[752];
  assign match_array[753] = N7242 & valid[753];
  assign N7242 = N7241 & N3858;
  assign N7241 = N4228 & en_i;
  assign empty_array[753] = N7243 & N7244;
  assign N7243 = N4228 & en_i;
  assign N7244 = ~valid[753];
  assign match_array[754] = N7246 & valid[754];
  assign N7246 = N7245 & N3859;
  assign N7245 = N4228 & en_i;
  assign empty_array[754] = N7247 & N7248;
  assign N7247 = N4228 & en_i;
  assign N7248 = ~valid[754];
  assign match_array[755] = N7250 & valid[755];
  assign N7250 = N7249 & N3860;
  assign N7249 = N4228 & en_i;
  assign empty_array[755] = N7251 & N7252;
  assign N7251 = N4228 & en_i;
  assign N7252 = ~valid[755];
  assign match_array[756] = N7254 & valid[756];
  assign N7254 = N7253 & N3861;
  assign N7253 = N4228 & en_i;
  assign empty_array[756] = N7255 & N7256;
  assign N7255 = N4228 & en_i;
  assign N7256 = ~valid[756];
  assign match_array[757] = N7258 & valid[757];
  assign N7258 = N7257 & N3862;
  assign N7257 = N4228 & en_i;
  assign empty_array[757] = N7259 & N7260;
  assign N7259 = N4228 & en_i;
  assign N7260 = ~valid[757];
  assign match_array[758] = N7262 & valid[758];
  assign N7262 = N7261 & N3863;
  assign N7261 = N4228 & en_i;
  assign empty_array[758] = N7263 & N7264;
  assign N7263 = N4228 & en_i;
  assign N7264 = ~valid[758];
  assign match_array[759] = N7266 & valid[759];
  assign N7266 = N7265 & N3864;
  assign N7265 = N4228 & en_i;
  assign empty_array[759] = N7267 & N7268;
  assign N7267 = N4228 & en_i;
  assign N7268 = ~valid[759];
  assign match_array[760] = N7270 & valid[760];
  assign N7270 = N7269 & N3865;
  assign N7269 = N4228 & en_i;
  assign empty_array[760] = N7271 & N7272;
  assign N7271 = N4228 & en_i;
  assign N7272 = ~valid[760];
  assign match_array[761] = N7274 & valid[761];
  assign N7274 = N7273 & N3866;
  assign N7273 = N4228 & en_i;
  assign empty_array[761] = N7275 & N7276;
  assign N7275 = N4228 & en_i;
  assign N7276 = ~valid[761];
  assign match_array[762] = N7278 & valid[762];
  assign N7278 = N7277 & N3867;
  assign N7277 = N4228 & en_i;
  assign empty_array[762] = N7279 & N7280;
  assign N7279 = N4228 & en_i;
  assign N7280 = ~valid[762];
  assign match_array[763] = N7282 & valid[763];
  assign N7282 = N7281 & N3868;
  assign N7281 = N4228 & en_i;
  assign empty_array[763] = N7283 & N7284;
  assign N7283 = N4228 & en_i;
  assign N7284 = ~valid[763];
  assign match_array[764] = N7286 & valid[764];
  assign N7286 = N7285 & N3869;
  assign N7285 = N4228 & en_i;
  assign empty_array[764] = N7287 & N7288;
  assign N7287 = N4228 & en_i;
  assign N7288 = ~valid[764];
  assign match_array[765] = N7290 & valid[765];
  assign N7290 = N7289 & N3870;
  assign N7289 = N4228 & en_i;
  assign empty_array[765] = N7291 & N7292;
  assign N7291 = N4228 & en_i;
  assign N7292 = ~valid[765];
  assign match_array[766] = N7294 & valid[766];
  assign N7294 = N7293 & N3871;
  assign N7293 = N4228 & en_i;
  assign empty_array[766] = N7295 & N7296;
  assign N7295 = N4228 & en_i;
  assign N7296 = ~valid[766];
  assign match_array[767] = N7298 & valid[767];
  assign N7298 = N7297 & N3872;
  assign N7297 = N4228 & en_i;
  assign empty_array[767] = N7299 & N7300;
  assign N7299 = N4228 & en_i;
  assign N7300 = ~valid[767];
  assign match_array[768] = N7302 & valid[768];
  assign N7302 = N7301 & N3873;
  assign N7301 = N4228 & en_i;
  assign empty_array[768] = N7303 & N7304;
  assign N7303 = N4228 & en_i;
  assign N7304 = ~valid[768];
  assign match_array[769] = N7306 & valid[769];
  assign N7306 = N7305 & N3874;
  assign N7305 = N4228 & en_i;
  assign empty_array[769] = N7307 & N7308;
  assign N7307 = N4228 & en_i;
  assign N7308 = ~valid[769];
  assign match_array[770] = N7310 & valid[770];
  assign N7310 = N7309 & N3875;
  assign N7309 = N4228 & en_i;
  assign empty_array[770] = N7311 & N7312;
  assign N7311 = N4228 & en_i;
  assign N7312 = ~valid[770];
  assign match_array[771] = N7314 & valid[771];
  assign N7314 = N7313 & N3876;
  assign N7313 = N4228 & en_i;
  assign empty_array[771] = N7315 & N7316;
  assign N7315 = N4228 & en_i;
  assign N7316 = ~valid[771];
  assign match_array[772] = N7318 & valid[772];
  assign N7318 = N7317 & N3877;
  assign N7317 = N4228 & en_i;
  assign empty_array[772] = N7319 & N7320;
  assign N7319 = N4228 & en_i;
  assign N7320 = ~valid[772];
  assign match_array[773] = N7322 & valid[773];
  assign N7322 = N7321 & N3878;
  assign N7321 = N4228 & en_i;
  assign empty_array[773] = N7323 & N7324;
  assign N7323 = N4228 & en_i;
  assign N7324 = ~valid[773];
  assign match_array[774] = N7326 & valid[774];
  assign N7326 = N7325 & N3879;
  assign N7325 = N4228 & en_i;
  assign empty_array[774] = N7327 & N7328;
  assign N7327 = N4228 & en_i;
  assign N7328 = ~valid[774];
  assign match_array[775] = N7330 & valid[775];
  assign N7330 = N7329 & N3880;
  assign N7329 = N4228 & en_i;
  assign empty_array[775] = N7331 & N7332;
  assign N7331 = N4228 & en_i;
  assign N7332 = ~valid[775];
  assign match_array[776] = N7334 & valid[776];
  assign N7334 = N7333 & N3881;
  assign N7333 = N4228 & en_i;
  assign empty_array[776] = N7335 & N7336;
  assign N7335 = N4228 & en_i;
  assign N7336 = ~valid[776];
  assign match_array[777] = N7338 & valid[777];
  assign N7338 = N7337 & N3882;
  assign N7337 = N4228 & en_i;
  assign empty_array[777] = N7339 & N7340;
  assign N7339 = N4228 & en_i;
  assign N7340 = ~valid[777];
  assign match_array[778] = N7342 & valid[778];
  assign N7342 = N7341 & N3883;
  assign N7341 = N4228 & en_i;
  assign empty_array[778] = N7343 & N7344;
  assign N7343 = N4228 & en_i;
  assign N7344 = ~valid[778];
  assign match_array[779] = N7346 & valid[779];
  assign N7346 = N7345 & N3884;
  assign N7345 = N4228 & en_i;
  assign empty_array[779] = N7347 & N7348;
  assign N7347 = N4228 & en_i;
  assign N7348 = ~valid[779];
  assign match_array[780] = N7350 & valid[780];
  assign N7350 = N7349 & N3885;
  assign N7349 = N4228 & en_i;
  assign empty_array[780] = N7351 & N7352;
  assign N7351 = N4228 & en_i;
  assign N7352 = ~valid[780];
  assign match_array[781] = N7354 & valid[781];
  assign N7354 = N7353 & N3886;
  assign N7353 = N4228 & en_i;
  assign empty_array[781] = N7355 & N7356;
  assign N7355 = N4228 & en_i;
  assign N7356 = ~valid[781];
  assign match_array[782] = N7358 & valid[782];
  assign N7358 = N7357 & N3887;
  assign N7357 = N4228 & en_i;
  assign empty_array[782] = N7359 & N7360;
  assign N7359 = N4228 & en_i;
  assign N7360 = ~valid[782];
  assign match_array[783] = N7362 & valid[783];
  assign N7362 = N7361 & N3888;
  assign N7361 = N4228 & en_i;
  assign empty_array[783] = N7363 & N7364;
  assign N7363 = N4228 & en_i;
  assign N7364 = ~valid[783];
  assign match_array[784] = N7366 & valid[784];
  assign N7366 = N7365 & N3889;
  assign N7365 = N4228 & en_i;
  assign empty_array[784] = N7367 & N7368;
  assign N7367 = N4228 & en_i;
  assign N7368 = ~valid[784];
  assign match_array[785] = N7370 & valid[785];
  assign N7370 = N7369 & N3890;
  assign N7369 = N4228 & en_i;
  assign empty_array[785] = N7371 & N7372;
  assign N7371 = N4228 & en_i;
  assign N7372 = ~valid[785];
  assign match_array[786] = N7374 & valid[786];
  assign N7374 = N7373 & N3891;
  assign N7373 = N4228 & en_i;
  assign empty_array[786] = N7375 & N7376;
  assign N7375 = N4228 & en_i;
  assign N7376 = ~valid[786];
  assign match_array[787] = N7378 & valid[787];
  assign N7378 = N7377 & N3892;
  assign N7377 = N4228 & en_i;
  assign empty_array[787] = N7379 & N7380;
  assign N7379 = N4228 & en_i;
  assign N7380 = ~valid[787];
  assign match_array[788] = N7382 & valid[788];
  assign N7382 = N7381 & N3893;
  assign N7381 = N4228 & en_i;
  assign empty_array[788] = N7383 & N7384;
  assign N7383 = N4228 & en_i;
  assign N7384 = ~valid[788];
  assign match_array[789] = N7386 & valid[789];
  assign N7386 = N7385 & N3894;
  assign N7385 = N4228 & en_i;
  assign empty_array[789] = N7387 & N7388;
  assign N7387 = N4228 & en_i;
  assign N7388 = ~valid[789];
  assign match_array[790] = N7390 & valid[790];
  assign N7390 = N7389 & N3895;
  assign N7389 = N4228 & en_i;
  assign empty_array[790] = N7391 & N7392;
  assign N7391 = N4228 & en_i;
  assign N7392 = ~valid[790];
  assign match_array[791] = N7394 & valid[791];
  assign N7394 = N7393 & N3896;
  assign N7393 = N4228 & en_i;
  assign empty_array[791] = N7395 & N7396;
  assign N7395 = N4228 & en_i;
  assign N7396 = ~valid[791];
  assign match_array[792] = N7398 & valid[792];
  assign N7398 = N7397 & N3897;
  assign N7397 = N4228 & en_i;
  assign empty_array[792] = N7399 & N7400;
  assign N7399 = N4228 & en_i;
  assign N7400 = ~valid[792];
  assign match_array[793] = N7402 & valid[793];
  assign N7402 = N7401 & N3898;
  assign N7401 = N4228 & en_i;
  assign empty_array[793] = N7403 & N7404;
  assign N7403 = N4228 & en_i;
  assign N7404 = ~valid[793];
  assign match_array[794] = N7406 & valid[794];
  assign N7406 = N7405 & N3899;
  assign N7405 = N4228 & en_i;
  assign empty_array[794] = N7407 & N7408;
  assign N7407 = N4228 & en_i;
  assign N7408 = ~valid[794];
  assign match_array[795] = N7410 & valid[795];
  assign N7410 = N7409 & N3900;
  assign N7409 = N4228 & en_i;
  assign empty_array[795] = N7411 & N7412;
  assign N7411 = N4228 & en_i;
  assign N7412 = ~valid[795];
  assign match_array[796] = N7414 & valid[796];
  assign N7414 = N7413 & N3901;
  assign N7413 = N4228 & en_i;
  assign empty_array[796] = N7415 & N7416;
  assign N7415 = N4228 & en_i;
  assign N7416 = ~valid[796];
  assign match_array[797] = N7418 & valid[797];
  assign N7418 = N7417 & N3902;
  assign N7417 = N4228 & en_i;
  assign empty_array[797] = N7419 & N7420;
  assign N7419 = N4228 & en_i;
  assign N7420 = ~valid[797];
  assign match_array[798] = N7422 & valid[798];
  assign N7422 = N7421 & N3903;
  assign N7421 = N4228 & en_i;
  assign empty_array[798] = N7423 & N7424;
  assign N7423 = N4228 & en_i;
  assign N7424 = ~valid[798];
  assign match_array[799] = N7426 & valid[799];
  assign N7426 = N7425 & N3904;
  assign N7425 = N4228 & en_i;
  assign empty_array[799] = N7427 & N7428;
  assign N7427 = N4228 & en_i;
  assign N7428 = ~valid[799];
  assign match_array[800] = N7430 & valid[800];
  assign N7430 = N7429 & N3905;
  assign N7429 = N4228 & en_i;
  assign empty_array[800] = N7431 & N7432;
  assign N7431 = N4228 & en_i;
  assign N7432 = ~valid[800];
  assign match_array[801] = N7434 & valid[801];
  assign N7434 = N7433 & N3906;
  assign N7433 = N4228 & en_i;
  assign empty_array[801] = N7435 & N7436;
  assign N7435 = N4228 & en_i;
  assign N7436 = ~valid[801];
  assign match_array[802] = N7438 & valid[802];
  assign N7438 = N7437 & N3907;
  assign N7437 = N4228 & en_i;
  assign empty_array[802] = N7439 & N7440;
  assign N7439 = N4228 & en_i;
  assign N7440 = ~valid[802];
  assign match_array[803] = N7442 & valid[803];
  assign N7442 = N7441 & N3908;
  assign N7441 = N4228 & en_i;
  assign empty_array[803] = N7443 & N7444;
  assign N7443 = N4228 & en_i;
  assign N7444 = ~valid[803];
  assign match_array[804] = N7446 & valid[804];
  assign N7446 = N7445 & N3909;
  assign N7445 = N4228 & en_i;
  assign empty_array[804] = N7447 & N7448;
  assign N7447 = N4228 & en_i;
  assign N7448 = ~valid[804];
  assign match_array[805] = N7450 & valid[805];
  assign N7450 = N7449 & N3910;
  assign N7449 = N4228 & en_i;
  assign empty_array[805] = N7451 & N7452;
  assign N7451 = N4228 & en_i;
  assign N7452 = ~valid[805];
  assign match_array[806] = N7454 & valid[806];
  assign N7454 = N7453 & N3911;
  assign N7453 = N4228 & en_i;
  assign empty_array[806] = N7455 & N7456;
  assign N7455 = N4228 & en_i;
  assign N7456 = ~valid[806];
  assign match_array[807] = N7458 & valid[807];
  assign N7458 = N7457 & N3912;
  assign N7457 = N4228 & en_i;
  assign empty_array[807] = N7459 & N7460;
  assign N7459 = N4228 & en_i;
  assign N7460 = ~valid[807];
  assign match_array[808] = N7462 & valid[808];
  assign N7462 = N7461 & N3913;
  assign N7461 = N4228 & en_i;
  assign empty_array[808] = N7463 & N7464;
  assign N7463 = N4228 & en_i;
  assign N7464 = ~valid[808];
  assign match_array[809] = N7466 & valid[809];
  assign N7466 = N7465 & N3914;
  assign N7465 = N4228 & en_i;
  assign empty_array[809] = N7467 & N7468;
  assign N7467 = N4228 & en_i;
  assign N7468 = ~valid[809];
  assign match_array[810] = N7470 & valid[810];
  assign N7470 = N7469 & N3915;
  assign N7469 = N4228 & en_i;
  assign empty_array[810] = N7471 & N7472;
  assign N7471 = N4228 & en_i;
  assign N7472 = ~valid[810];
  assign match_array[811] = N7474 & valid[811];
  assign N7474 = N7473 & N3916;
  assign N7473 = N4228 & en_i;
  assign empty_array[811] = N7475 & N7476;
  assign N7475 = N4228 & en_i;
  assign N7476 = ~valid[811];
  assign match_array[812] = N7478 & valid[812];
  assign N7478 = N7477 & N3917;
  assign N7477 = N4228 & en_i;
  assign empty_array[812] = N7479 & N7480;
  assign N7479 = N4228 & en_i;
  assign N7480 = ~valid[812];
  assign match_array[813] = N7482 & valid[813];
  assign N7482 = N7481 & N3918;
  assign N7481 = N4228 & en_i;
  assign empty_array[813] = N7483 & N7484;
  assign N7483 = N4228 & en_i;
  assign N7484 = ~valid[813];
  assign match_array[814] = N7486 & valid[814];
  assign N7486 = N7485 & N3919;
  assign N7485 = N4228 & en_i;
  assign empty_array[814] = N7487 & N7488;
  assign N7487 = N4228 & en_i;
  assign N7488 = ~valid[814];
  assign match_array[815] = N7490 & valid[815];
  assign N7490 = N7489 & N3920;
  assign N7489 = N4228 & en_i;
  assign empty_array[815] = N7491 & N7492;
  assign N7491 = N4228 & en_i;
  assign N7492 = ~valid[815];
  assign match_array[816] = N7494 & valid[816];
  assign N7494 = N7493 & N3921;
  assign N7493 = N4228 & en_i;
  assign empty_array[816] = N7495 & N7496;
  assign N7495 = N4228 & en_i;
  assign N7496 = ~valid[816];
  assign match_array[817] = N7498 & valid[817];
  assign N7498 = N7497 & N3922;
  assign N7497 = N4228 & en_i;
  assign empty_array[817] = N7499 & N7500;
  assign N7499 = N4228 & en_i;
  assign N7500 = ~valid[817];
  assign match_array[818] = N7502 & valid[818];
  assign N7502 = N7501 & N3923;
  assign N7501 = N4228 & en_i;
  assign empty_array[818] = N7503 & N7504;
  assign N7503 = N4228 & en_i;
  assign N7504 = ~valid[818];
  assign match_array[819] = N7506 & valid[819];
  assign N7506 = N7505 & N3924;
  assign N7505 = N4228 & en_i;
  assign empty_array[819] = N7507 & N7508;
  assign N7507 = N4228 & en_i;
  assign N7508 = ~valid[819];
  assign match_array[820] = N7510 & valid[820];
  assign N7510 = N7509 & N3925;
  assign N7509 = N4228 & en_i;
  assign empty_array[820] = N7511 & N7512;
  assign N7511 = N4228 & en_i;
  assign N7512 = ~valid[820];
  assign match_array[821] = N7514 & valid[821];
  assign N7514 = N7513 & N3926;
  assign N7513 = N4228 & en_i;
  assign empty_array[821] = N7515 & N7516;
  assign N7515 = N4228 & en_i;
  assign N7516 = ~valid[821];
  assign match_array[822] = N7518 & valid[822];
  assign N7518 = N7517 & N3927;
  assign N7517 = N4228 & en_i;
  assign empty_array[822] = N7519 & N7520;
  assign N7519 = N4228 & en_i;
  assign N7520 = ~valid[822];
  assign match_array[823] = N7522 & valid[823];
  assign N7522 = N7521 & N3928;
  assign N7521 = N4228 & en_i;
  assign empty_array[823] = N7523 & N7524;
  assign N7523 = N4228 & en_i;
  assign N7524 = ~valid[823];
  assign match_array[824] = N7526 & valid[824];
  assign N7526 = N7525 & N3929;
  assign N7525 = N4228 & en_i;
  assign empty_array[824] = N7527 & N7528;
  assign N7527 = N4228 & en_i;
  assign N7528 = ~valid[824];
  assign match_array[825] = N7530 & valid[825];
  assign N7530 = N7529 & N3930;
  assign N7529 = N4228 & en_i;
  assign empty_array[825] = N7531 & N7532;
  assign N7531 = N4228 & en_i;
  assign N7532 = ~valid[825];
  assign match_array[826] = N7534 & valid[826];
  assign N7534 = N7533 & N3931;
  assign N7533 = N4228 & en_i;
  assign empty_array[826] = N7535 & N7536;
  assign N7535 = N4228 & en_i;
  assign N7536 = ~valid[826];
  assign match_array[827] = N7538 & valid[827];
  assign N7538 = N7537 & N3932;
  assign N7537 = N4228 & en_i;
  assign empty_array[827] = N7539 & N7540;
  assign N7539 = N4228 & en_i;
  assign N7540 = ~valid[827];
  assign match_array[828] = N7542 & valid[828];
  assign N7542 = N7541 & N3933;
  assign N7541 = N4228 & en_i;
  assign empty_array[828] = N7543 & N7544;
  assign N7543 = N4228 & en_i;
  assign N7544 = ~valid[828];
  assign match_array[829] = N7546 & valid[829];
  assign N7546 = N7545 & N3934;
  assign N7545 = N4228 & en_i;
  assign empty_array[829] = N7547 & N7548;
  assign N7547 = N4228 & en_i;
  assign N7548 = ~valid[829];
  assign match_array[830] = N7550 & valid[830];
  assign N7550 = N7549 & N3935;
  assign N7549 = N4228 & en_i;
  assign empty_array[830] = N7551 & N7552;
  assign N7551 = N4228 & en_i;
  assign N7552 = ~valid[830];
  assign match_array[831] = N7554 & valid[831];
  assign N7554 = N7553 & N3936;
  assign N7553 = N4228 & en_i;
  assign empty_array[831] = N7555 & N7556;
  assign N7555 = N4228 & en_i;
  assign N7556 = ~valid[831];
  assign match_array[832] = N7558 & valid[832];
  assign N7558 = N7557 & N3937;
  assign N7557 = N4228 & en_i;
  assign empty_array[832] = N7559 & N7560;
  assign N7559 = N4228 & en_i;
  assign N7560 = ~valid[832];
  assign match_array[833] = N7562 & valid[833];
  assign N7562 = N7561 & N3938;
  assign N7561 = N4228 & en_i;
  assign empty_array[833] = N7563 & N7564;
  assign N7563 = N4228 & en_i;
  assign N7564 = ~valid[833];
  assign match_array[834] = N7566 & valid[834];
  assign N7566 = N7565 & N3939;
  assign N7565 = N4228 & en_i;
  assign empty_array[834] = N7567 & N7568;
  assign N7567 = N4228 & en_i;
  assign N7568 = ~valid[834];
  assign match_array[835] = N7570 & valid[835];
  assign N7570 = N7569 & N3940;
  assign N7569 = N4228 & en_i;
  assign empty_array[835] = N7571 & N7572;
  assign N7571 = N4228 & en_i;
  assign N7572 = ~valid[835];
  assign match_array[836] = N7574 & valid[836];
  assign N7574 = N7573 & N3941;
  assign N7573 = N4228 & en_i;
  assign empty_array[836] = N7575 & N7576;
  assign N7575 = N4228 & en_i;
  assign N7576 = ~valid[836];
  assign match_array[837] = N7578 & valid[837];
  assign N7578 = N7577 & N3942;
  assign N7577 = N4228 & en_i;
  assign empty_array[837] = N7579 & N7580;
  assign N7579 = N4228 & en_i;
  assign N7580 = ~valid[837];
  assign match_array[838] = N7582 & valid[838];
  assign N7582 = N7581 & N3943;
  assign N7581 = N4228 & en_i;
  assign empty_array[838] = N7583 & N7584;
  assign N7583 = N4228 & en_i;
  assign N7584 = ~valid[838];
  assign match_array[839] = N7586 & valid[839];
  assign N7586 = N7585 & N3944;
  assign N7585 = N4228 & en_i;
  assign empty_array[839] = N7587 & N7588;
  assign N7587 = N4228 & en_i;
  assign N7588 = ~valid[839];
  assign match_array[840] = N7590 & valid[840];
  assign N7590 = N7589 & N3945;
  assign N7589 = N4228 & en_i;
  assign empty_array[840] = N7591 & N7592;
  assign N7591 = N4228 & en_i;
  assign N7592 = ~valid[840];
  assign match_array[841] = N7594 & valid[841];
  assign N7594 = N7593 & N3946;
  assign N7593 = N4228 & en_i;
  assign empty_array[841] = N7595 & N7596;
  assign N7595 = N4228 & en_i;
  assign N7596 = ~valid[841];
  assign match_array[842] = N7598 & valid[842];
  assign N7598 = N7597 & N3947;
  assign N7597 = N4228 & en_i;
  assign empty_array[842] = N7599 & N7600;
  assign N7599 = N4228 & en_i;
  assign N7600 = ~valid[842];
  assign match_array[843] = N7602 & valid[843];
  assign N7602 = N7601 & N3948;
  assign N7601 = N4228 & en_i;
  assign empty_array[843] = N7603 & N7604;
  assign N7603 = N4228 & en_i;
  assign N7604 = ~valid[843];
  assign match_array[844] = N7606 & valid[844];
  assign N7606 = N7605 & N3949;
  assign N7605 = N4228 & en_i;
  assign empty_array[844] = N7607 & N7608;
  assign N7607 = N4228 & en_i;
  assign N7608 = ~valid[844];
  assign match_array[845] = N7610 & valid[845];
  assign N7610 = N7609 & N3950;
  assign N7609 = N4228 & en_i;
  assign empty_array[845] = N7611 & N7612;
  assign N7611 = N4228 & en_i;
  assign N7612 = ~valid[845];
  assign match_array[846] = N7614 & valid[846];
  assign N7614 = N7613 & N3951;
  assign N7613 = N4228 & en_i;
  assign empty_array[846] = N7615 & N7616;
  assign N7615 = N4228 & en_i;
  assign N7616 = ~valid[846];
  assign match_array[847] = N7618 & valid[847];
  assign N7618 = N7617 & N3952;
  assign N7617 = N4228 & en_i;
  assign empty_array[847] = N7619 & N7620;
  assign N7619 = N4228 & en_i;
  assign N7620 = ~valid[847];
  assign match_array[848] = N7622 & valid[848];
  assign N7622 = N7621 & N3953;
  assign N7621 = N4228 & en_i;
  assign empty_array[848] = N7623 & N7624;
  assign N7623 = N4228 & en_i;
  assign N7624 = ~valid[848];
  assign match_array[849] = N7626 & valid[849];
  assign N7626 = N7625 & N3954;
  assign N7625 = N4228 & en_i;
  assign empty_array[849] = N7627 & N7628;
  assign N7627 = N4228 & en_i;
  assign N7628 = ~valid[849];
  assign match_array[850] = N7630 & valid[850];
  assign N7630 = N7629 & N3955;
  assign N7629 = N4228 & en_i;
  assign empty_array[850] = N7631 & N7632;
  assign N7631 = N4228 & en_i;
  assign N7632 = ~valid[850];
  assign match_array[851] = N7634 & valid[851];
  assign N7634 = N7633 & N3956;
  assign N7633 = N4228 & en_i;
  assign empty_array[851] = N7635 & N7636;
  assign N7635 = N4228 & en_i;
  assign N7636 = ~valid[851];
  assign match_array[852] = N7638 & valid[852];
  assign N7638 = N7637 & N3957;
  assign N7637 = N4228 & en_i;
  assign empty_array[852] = N7639 & N7640;
  assign N7639 = N4228 & en_i;
  assign N7640 = ~valid[852];
  assign match_array[853] = N7642 & valid[853];
  assign N7642 = N7641 & N3958;
  assign N7641 = N4228 & en_i;
  assign empty_array[853] = N7643 & N7644;
  assign N7643 = N4228 & en_i;
  assign N7644 = ~valid[853];
  assign match_array[854] = N7646 & valid[854];
  assign N7646 = N7645 & N3959;
  assign N7645 = N4228 & en_i;
  assign empty_array[854] = N7647 & N7648;
  assign N7647 = N4228 & en_i;
  assign N7648 = ~valid[854];
  assign match_array[855] = N7650 & valid[855];
  assign N7650 = N7649 & N3960;
  assign N7649 = N4228 & en_i;
  assign empty_array[855] = N7651 & N7652;
  assign N7651 = N4228 & en_i;
  assign N7652 = ~valid[855];
  assign match_array[856] = N7654 & valid[856];
  assign N7654 = N7653 & N3961;
  assign N7653 = N4228 & en_i;
  assign empty_array[856] = N7655 & N7656;
  assign N7655 = N4228 & en_i;
  assign N7656 = ~valid[856];
  assign match_array[857] = N7658 & valid[857];
  assign N7658 = N7657 & N3962;
  assign N7657 = N4228 & en_i;
  assign empty_array[857] = N7659 & N7660;
  assign N7659 = N4228 & en_i;
  assign N7660 = ~valid[857];
  assign match_array[858] = N7662 & valid[858];
  assign N7662 = N7661 & N3963;
  assign N7661 = N4228 & en_i;
  assign empty_array[858] = N7663 & N7664;
  assign N7663 = N4228 & en_i;
  assign N7664 = ~valid[858];
  assign match_array[859] = N7666 & valid[859];
  assign N7666 = N7665 & N3964;
  assign N7665 = N4228 & en_i;
  assign empty_array[859] = N7667 & N7668;
  assign N7667 = N4228 & en_i;
  assign N7668 = ~valid[859];
  assign match_array[860] = N7670 & valid[860];
  assign N7670 = N7669 & N3965;
  assign N7669 = N4228 & en_i;
  assign empty_array[860] = N7671 & N7672;
  assign N7671 = N4228 & en_i;
  assign N7672 = ~valid[860];
  assign match_array[861] = N7674 & valid[861];
  assign N7674 = N7673 & N3966;
  assign N7673 = N4228 & en_i;
  assign empty_array[861] = N7675 & N7676;
  assign N7675 = N4228 & en_i;
  assign N7676 = ~valid[861];
  assign match_array[862] = N7678 & valid[862];
  assign N7678 = N7677 & N3967;
  assign N7677 = N4228 & en_i;
  assign empty_array[862] = N7679 & N7680;
  assign N7679 = N4228 & en_i;
  assign N7680 = ~valid[862];
  assign match_array[863] = N7682 & valid[863];
  assign N7682 = N7681 & N3968;
  assign N7681 = N4228 & en_i;
  assign empty_array[863] = N7683 & N7684;
  assign N7683 = N4228 & en_i;
  assign N7684 = ~valid[863];
  assign match_array[864] = N7686 & valid[864];
  assign N7686 = N7685 & N3969;
  assign N7685 = N4228 & en_i;
  assign empty_array[864] = N7687 & N7688;
  assign N7687 = N4228 & en_i;
  assign N7688 = ~valid[864];
  assign match_array[865] = N7690 & valid[865];
  assign N7690 = N7689 & N3970;
  assign N7689 = N4228 & en_i;
  assign empty_array[865] = N7691 & N7692;
  assign N7691 = N4228 & en_i;
  assign N7692 = ~valid[865];
  assign match_array[866] = N7694 & valid[866];
  assign N7694 = N7693 & N3971;
  assign N7693 = N4228 & en_i;
  assign empty_array[866] = N7695 & N7696;
  assign N7695 = N4228 & en_i;
  assign N7696 = ~valid[866];
  assign match_array[867] = N7698 & valid[867];
  assign N7698 = N7697 & N3972;
  assign N7697 = N4228 & en_i;
  assign empty_array[867] = N7699 & N7700;
  assign N7699 = N4228 & en_i;
  assign N7700 = ~valid[867];
  assign match_array[868] = N7702 & valid[868];
  assign N7702 = N7701 & N3973;
  assign N7701 = N4228 & en_i;
  assign empty_array[868] = N7703 & N7704;
  assign N7703 = N4228 & en_i;
  assign N7704 = ~valid[868];
  assign match_array[869] = N7706 & valid[869];
  assign N7706 = N7705 & N3974;
  assign N7705 = N4228 & en_i;
  assign empty_array[869] = N7707 & N7708;
  assign N7707 = N4228 & en_i;
  assign N7708 = ~valid[869];
  assign match_array[870] = N7710 & valid[870];
  assign N7710 = N7709 & N3975;
  assign N7709 = N4228 & en_i;
  assign empty_array[870] = N7711 & N7712;
  assign N7711 = N4228 & en_i;
  assign N7712 = ~valid[870];
  assign match_array[871] = N7714 & valid[871];
  assign N7714 = N7713 & N3976;
  assign N7713 = N4228 & en_i;
  assign empty_array[871] = N7715 & N7716;
  assign N7715 = N4228 & en_i;
  assign N7716 = ~valid[871];
  assign match_array[872] = N7718 & valid[872];
  assign N7718 = N7717 & N3977;
  assign N7717 = N4228 & en_i;
  assign empty_array[872] = N7719 & N7720;
  assign N7719 = N4228 & en_i;
  assign N7720 = ~valid[872];
  assign match_array[873] = N7722 & valid[873];
  assign N7722 = N7721 & N3978;
  assign N7721 = N4228 & en_i;
  assign empty_array[873] = N7723 & N7724;
  assign N7723 = N4228 & en_i;
  assign N7724 = ~valid[873];
  assign match_array[874] = N7726 & valid[874];
  assign N7726 = N7725 & N3979;
  assign N7725 = N4228 & en_i;
  assign empty_array[874] = N7727 & N7728;
  assign N7727 = N4228 & en_i;
  assign N7728 = ~valid[874];
  assign match_array[875] = N7730 & valid[875];
  assign N7730 = N7729 & N3980;
  assign N7729 = N4228 & en_i;
  assign empty_array[875] = N7731 & N7732;
  assign N7731 = N4228 & en_i;
  assign N7732 = ~valid[875];
  assign match_array[876] = N7734 & valid[876];
  assign N7734 = N7733 & N3981;
  assign N7733 = N4228 & en_i;
  assign empty_array[876] = N7735 & N7736;
  assign N7735 = N4228 & en_i;
  assign N7736 = ~valid[876];
  assign match_array[877] = N7738 & valid[877];
  assign N7738 = N7737 & N3982;
  assign N7737 = N4228 & en_i;
  assign empty_array[877] = N7739 & N7740;
  assign N7739 = N4228 & en_i;
  assign N7740 = ~valid[877];
  assign match_array[878] = N7742 & valid[878];
  assign N7742 = N7741 & N3983;
  assign N7741 = N4228 & en_i;
  assign empty_array[878] = N7743 & N7744;
  assign N7743 = N4228 & en_i;
  assign N7744 = ~valid[878];
  assign match_array[879] = N7746 & valid[879];
  assign N7746 = N7745 & N3984;
  assign N7745 = N4228 & en_i;
  assign empty_array[879] = N7747 & N7748;
  assign N7747 = N4228 & en_i;
  assign N7748 = ~valid[879];
  assign match_array[880] = N7750 & valid[880];
  assign N7750 = N7749 & N3985;
  assign N7749 = N4228 & en_i;
  assign empty_array[880] = N7751 & N7752;
  assign N7751 = N4228 & en_i;
  assign N7752 = ~valid[880];
  assign match_array[881] = N7754 & valid[881];
  assign N7754 = N7753 & N3986;
  assign N7753 = N4228 & en_i;
  assign empty_array[881] = N7755 & N7756;
  assign N7755 = N4228 & en_i;
  assign N7756 = ~valid[881];
  assign match_array[882] = N7758 & valid[882];
  assign N7758 = N7757 & N3987;
  assign N7757 = N4228 & en_i;
  assign empty_array[882] = N7759 & N7760;
  assign N7759 = N4228 & en_i;
  assign N7760 = ~valid[882];
  assign match_array[883] = N7762 & valid[883];
  assign N7762 = N7761 & N3988;
  assign N7761 = N4228 & en_i;
  assign empty_array[883] = N7763 & N7764;
  assign N7763 = N4228 & en_i;
  assign N7764 = ~valid[883];
  assign match_array[884] = N7766 & valid[884];
  assign N7766 = N7765 & N3989;
  assign N7765 = N4228 & en_i;
  assign empty_array[884] = N7767 & N7768;
  assign N7767 = N4228 & en_i;
  assign N7768 = ~valid[884];
  assign match_array[885] = N7770 & valid[885];
  assign N7770 = N7769 & N3990;
  assign N7769 = N4228 & en_i;
  assign empty_array[885] = N7771 & N7772;
  assign N7771 = N4228 & en_i;
  assign N7772 = ~valid[885];
  assign match_array[886] = N7774 & valid[886];
  assign N7774 = N7773 & N3991;
  assign N7773 = N4228 & en_i;
  assign empty_array[886] = N7775 & N7776;
  assign N7775 = N4228 & en_i;
  assign N7776 = ~valid[886];
  assign match_array[887] = N7778 & valid[887];
  assign N7778 = N7777 & N3992;
  assign N7777 = N4228 & en_i;
  assign empty_array[887] = N7779 & N7780;
  assign N7779 = N4228 & en_i;
  assign N7780 = ~valid[887];
  assign match_array[888] = N7782 & valid[888];
  assign N7782 = N7781 & N3993;
  assign N7781 = N4228 & en_i;
  assign empty_array[888] = N7783 & N7784;
  assign N7783 = N4228 & en_i;
  assign N7784 = ~valid[888];
  assign match_array[889] = N7786 & valid[889];
  assign N7786 = N7785 & N3994;
  assign N7785 = N4228 & en_i;
  assign empty_array[889] = N7787 & N7788;
  assign N7787 = N4228 & en_i;
  assign N7788 = ~valid[889];
  assign match_array[890] = N7790 & valid[890];
  assign N7790 = N7789 & N3995;
  assign N7789 = N4228 & en_i;
  assign empty_array[890] = N7791 & N7792;
  assign N7791 = N4228 & en_i;
  assign N7792 = ~valid[890];
  assign match_array[891] = N7794 & valid[891];
  assign N7794 = N7793 & N3996;
  assign N7793 = N4228 & en_i;
  assign empty_array[891] = N7795 & N7796;
  assign N7795 = N4228 & en_i;
  assign N7796 = ~valid[891];
  assign match_array[892] = N7798 & valid[892];
  assign N7798 = N7797 & N3997;
  assign N7797 = N4228 & en_i;
  assign empty_array[892] = N7799 & N7800;
  assign N7799 = N4228 & en_i;
  assign N7800 = ~valid[892];
  assign match_array[893] = N7802 & valid[893];
  assign N7802 = N7801 & N3998;
  assign N7801 = N4228 & en_i;
  assign empty_array[893] = N7803 & N7804;
  assign N7803 = N4228 & en_i;
  assign N7804 = ~valid[893];
  assign match_array[894] = N7806 & valid[894];
  assign N7806 = N7805 & N3999;
  assign N7805 = N4228 & en_i;
  assign empty_array[894] = N7807 & N7808;
  assign N7807 = N4228 & en_i;
  assign N7808 = ~valid[894];
  assign match_array[895] = N7810 & valid[895];
  assign N7810 = N7809 & N4000;
  assign N7809 = N4228 & en_i;
  assign empty_array[895] = N7811 & N7812;
  assign N7811 = N4228 & en_i;
  assign N7812 = ~valid[895];
  assign match_array[896] = N7814 & valid[896];
  assign N7814 = N7813 & N4001;
  assign N7813 = N4228 & en_i;
  assign empty_array[896] = N7815 & N7816;
  assign N7815 = N4228 & en_i;
  assign N7816 = ~valid[896];
  assign match_array[897] = N7818 & valid[897];
  assign N7818 = N7817 & N4002;
  assign N7817 = N4228 & en_i;
  assign empty_array[897] = N7819 & N7820;
  assign N7819 = N4228 & en_i;
  assign N7820 = ~valid[897];
  assign match_array[898] = N7822 & valid[898];
  assign N7822 = N7821 & N4003;
  assign N7821 = N4228 & en_i;
  assign empty_array[898] = N7823 & N7824;
  assign N7823 = N4228 & en_i;
  assign N7824 = ~valid[898];
  assign match_array[899] = N7826 & valid[899];
  assign N7826 = N7825 & N4004;
  assign N7825 = N4228 & en_i;
  assign empty_array[899] = N7827 & N7828;
  assign N7827 = N4228 & en_i;
  assign N7828 = ~valid[899];
  assign match_array[900] = N7830 & valid[900];
  assign N7830 = N7829 & N4005;
  assign N7829 = N4228 & en_i;
  assign empty_array[900] = N7831 & N7832;
  assign N7831 = N4228 & en_i;
  assign N7832 = ~valid[900];
  assign match_array[901] = N7834 & valid[901];
  assign N7834 = N7833 & N4006;
  assign N7833 = N4228 & en_i;
  assign empty_array[901] = N7835 & N7836;
  assign N7835 = N4228 & en_i;
  assign N7836 = ~valid[901];
  assign match_array[902] = N7838 & valid[902];
  assign N7838 = N7837 & N4007;
  assign N7837 = N4228 & en_i;
  assign empty_array[902] = N7839 & N7840;
  assign N7839 = N4228 & en_i;
  assign N7840 = ~valid[902];
  assign match_array[903] = N7842 & valid[903];
  assign N7842 = N7841 & N4008;
  assign N7841 = N4228 & en_i;
  assign empty_array[903] = N7843 & N7844;
  assign N7843 = N4228 & en_i;
  assign N7844 = ~valid[903];
  assign match_array[904] = N7846 & valid[904];
  assign N7846 = N7845 & N4009;
  assign N7845 = N4228 & en_i;
  assign empty_array[904] = N7847 & N7848;
  assign N7847 = N4228 & en_i;
  assign N7848 = ~valid[904];
  assign match_array[905] = N7850 & valid[905];
  assign N7850 = N7849 & N4010;
  assign N7849 = N4228 & en_i;
  assign empty_array[905] = N7851 & N7852;
  assign N7851 = N4228 & en_i;
  assign N7852 = ~valid[905];
  assign match_array[906] = N7854 & valid[906];
  assign N7854 = N7853 & N4011;
  assign N7853 = N4228 & en_i;
  assign empty_array[906] = N7855 & N7856;
  assign N7855 = N4228 & en_i;
  assign N7856 = ~valid[906];
  assign match_array[907] = N7858 & valid[907];
  assign N7858 = N7857 & N4012;
  assign N7857 = N4228 & en_i;
  assign empty_array[907] = N7859 & N7860;
  assign N7859 = N4228 & en_i;
  assign N7860 = ~valid[907];
  assign match_array[908] = N7862 & valid[908];
  assign N7862 = N7861 & N4013;
  assign N7861 = N4228 & en_i;
  assign empty_array[908] = N7863 & N7864;
  assign N7863 = N4228 & en_i;
  assign N7864 = ~valid[908];
  assign match_array[909] = N7866 & valid[909];
  assign N7866 = N7865 & N4014;
  assign N7865 = N4228 & en_i;
  assign empty_array[909] = N7867 & N7868;
  assign N7867 = N4228 & en_i;
  assign N7868 = ~valid[909];
  assign match_array[910] = N7870 & valid[910];
  assign N7870 = N7869 & N4015;
  assign N7869 = N4228 & en_i;
  assign empty_array[910] = N7871 & N7872;
  assign N7871 = N4228 & en_i;
  assign N7872 = ~valid[910];
  assign match_array[911] = N7874 & valid[911];
  assign N7874 = N7873 & N4016;
  assign N7873 = N4228 & en_i;
  assign empty_array[911] = N7875 & N7876;
  assign N7875 = N4228 & en_i;
  assign N7876 = ~valid[911];
  assign match_array[912] = N7878 & valid[912];
  assign N7878 = N7877 & N4017;
  assign N7877 = N4228 & en_i;
  assign empty_array[912] = N7879 & N7880;
  assign N7879 = N4228 & en_i;
  assign N7880 = ~valid[912];
  assign match_array[913] = N7882 & valid[913];
  assign N7882 = N7881 & N4018;
  assign N7881 = N4228 & en_i;
  assign empty_array[913] = N7883 & N7884;
  assign N7883 = N4228 & en_i;
  assign N7884 = ~valid[913];
  assign match_array[914] = N7886 & valid[914];
  assign N7886 = N7885 & N4019;
  assign N7885 = N4228 & en_i;
  assign empty_array[914] = N7887 & N7888;
  assign N7887 = N4228 & en_i;
  assign N7888 = ~valid[914];
  assign match_array[915] = N7890 & valid[915];
  assign N7890 = N7889 & N4020;
  assign N7889 = N4228 & en_i;
  assign empty_array[915] = N7891 & N7892;
  assign N7891 = N4228 & en_i;
  assign N7892 = ~valid[915];
  assign match_array[916] = N7894 & valid[916];
  assign N7894 = N7893 & N4021;
  assign N7893 = N4228 & en_i;
  assign empty_array[916] = N7895 & N7896;
  assign N7895 = N4228 & en_i;
  assign N7896 = ~valid[916];
  assign match_array[917] = N7898 & valid[917];
  assign N7898 = N7897 & N4022;
  assign N7897 = N4228 & en_i;
  assign empty_array[917] = N7899 & N7900;
  assign N7899 = N4228 & en_i;
  assign N7900 = ~valid[917];
  assign match_array[918] = N7902 & valid[918];
  assign N7902 = N7901 & N4023;
  assign N7901 = N4228 & en_i;
  assign empty_array[918] = N7903 & N7904;
  assign N7903 = N4228 & en_i;
  assign N7904 = ~valid[918];
  assign match_array[919] = N7906 & valid[919];
  assign N7906 = N7905 & N4024;
  assign N7905 = N4228 & en_i;
  assign empty_array[919] = N7907 & N7908;
  assign N7907 = N4228 & en_i;
  assign N7908 = ~valid[919];
  assign match_array[920] = N7910 & valid[920];
  assign N7910 = N7909 & N4025;
  assign N7909 = N4228 & en_i;
  assign empty_array[920] = N7911 & N7912;
  assign N7911 = N4228 & en_i;
  assign N7912 = ~valid[920];
  assign match_array[921] = N7914 & valid[921];
  assign N7914 = N7913 & N4026;
  assign N7913 = N4228 & en_i;
  assign empty_array[921] = N7915 & N7916;
  assign N7915 = N4228 & en_i;
  assign N7916 = ~valid[921];
  assign match_array[922] = N7918 & valid[922];
  assign N7918 = N7917 & N4027;
  assign N7917 = N4228 & en_i;
  assign empty_array[922] = N7919 & N7920;
  assign N7919 = N4228 & en_i;
  assign N7920 = ~valid[922];
  assign match_array[923] = N7922 & valid[923];
  assign N7922 = N7921 & N4028;
  assign N7921 = N4228 & en_i;
  assign empty_array[923] = N7923 & N7924;
  assign N7923 = N4228 & en_i;
  assign N7924 = ~valid[923];
  assign match_array[924] = N7926 & valid[924];
  assign N7926 = N7925 & N4029;
  assign N7925 = N4228 & en_i;
  assign empty_array[924] = N7927 & N7928;
  assign N7927 = N4228 & en_i;
  assign N7928 = ~valid[924];
  assign match_array[925] = N7930 & valid[925];
  assign N7930 = N7929 & N4030;
  assign N7929 = N4228 & en_i;
  assign empty_array[925] = N7931 & N7932;
  assign N7931 = N4228 & en_i;
  assign N7932 = ~valid[925];
  assign match_array[926] = N7934 & valid[926];
  assign N7934 = N7933 & N4031;
  assign N7933 = N4228 & en_i;
  assign empty_array[926] = N7935 & N7936;
  assign N7935 = N4228 & en_i;
  assign N7936 = ~valid[926];
  assign match_array[927] = N7938 & valid[927];
  assign N7938 = N7937 & N4032;
  assign N7937 = N4228 & en_i;
  assign empty_array[927] = N7939 & N7940;
  assign N7939 = N4228 & en_i;
  assign N7940 = ~valid[927];
  assign match_array[928] = N7942 & valid[928];
  assign N7942 = N7941 & N4033;
  assign N7941 = N4228 & en_i;
  assign empty_array[928] = N7943 & N7944;
  assign N7943 = N4228 & en_i;
  assign N7944 = ~valid[928];
  assign match_array[929] = N7946 & valid[929];
  assign N7946 = N7945 & N4034;
  assign N7945 = N4228 & en_i;
  assign empty_array[929] = N7947 & N7948;
  assign N7947 = N4228 & en_i;
  assign N7948 = ~valid[929];
  assign match_array[930] = N7950 & valid[930];
  assign N7950 = N7949 & N4035;
  assign N7949 = N4228 & en_i;
  assign empty_array[930] = N7951 & N7952;
  assign N7951 = N4228 & en_i;
  assign N7952 = ~valid[930];
  assign match_array[931] = N7954 & valid[931];
  assign N7954 = N7953 & N4036;
  assign N7953 = N4228 & en_i;
  assign empty_array[931] = N7955 & N7956;
  assign N7955 = N4228 & en_i;
  assign N7956 = ~valid[931];
  assign match_array[932] = N7958 & valid[932];
  assign N7958 = N7957 & N4037;
  assign N7957 = N4228 & en_i;
  assign empty_array[932] = N7959 & N7960;
  assign N7959 = N4228 & en_i;
  assign N7960 = ~valid[932];
  assign match_array[933] = N7962 & valid[933];
  assign N7962 = N7961 & N4038;
  assign N7961 = N4228 & en_i;
  assign empty_array[933] = N7963 & N7964;
  assign N7963 = N4228 & en_i;
  assign N7964 = ~valid[933];
  assign match_array[934] = N7966 & valid[934];
  assign N7966 = N7965 & N4039;
  assign N7965 = N4228 & en_i;
  assign empty_array[934] = N7967 & N7968;
  assign N7967 = N4228 & en_i;
  assign N7968 = ~valid[934];
  assign match_array[935] = N7970 & valid[935];
  assign N7970 = N7969 & N4040;
  assign N7969 = N4228 & en_i;
  assign empty_array[935] = N7971 & N7972;
  assign N7971 = N4228 & en_i;
  assign N7972 = ~valid[935];
  assign match_array[936] = N7974 & valid[936];
  assign N7974 = N7973 & N4041;
  assign N7973 = N4228 & en_i;
  assign empty_array[936] = N7975 & N7976;
  assign N7975 = N4228 & en_i;
  assign N7976 = ~valid[936];
  assign match_array[937] = N7978 & valid[937];
  assign N7978 = N7977 & N4042;
  assign N7977 = N4228 & en_i;
  assign empty_array[937] = N7979 & N7980;
  assign N7979 = N4228 & en_i;
  assign N7980 = ~valid[937];
  assign match_array[938] = N7982 & valid[938];
  assign N7982 = N7981 & N4043;
  assign N7981 = N4228 & en_i;
  assign empty_array[938] = N7983 & N7984;
  assign N7983 = N4228 & en_i;
  assign N7984 = ~valid[938];
  assign match_array[939] = N7986 & valid[939];
  assign N7986 = N7985 & N4044;
  assign N7985 = N4228 & en_i;
  assign empty_array[939] = N7987 & N7988;
  assign N7987 = N4228 & en_i;
  assign N7988 = ~valid[939];
  assign match_array[940] = N7990 & valid[940];
  assign N7990 = N7989 & N4045;
  assign N7989 = N4228 & en_i;
  assign empty_array[940] = N7991 & N7992;
  assign N7991 = N4228 & en_i;
  assign N7992 = ~valid[940];
  assign match_array[941] = N7994 & valid[941];
  assign N7994 = N7993 & N4046;
  assign N7993 = N4228 & en_i;
  assign empty_array[941] = N7995 & N7996;
  assign N7995 = N4228 & en_i;
  assign N7996 = ~valid[941];
  assign match_array[942] = N7998 & valid[942];
  assign N7998 = N7997 & N4047;
  assign N7997 = N4228 & en_i;
  assign empty_array[942] = N7999 & N8000;
  assign N7999 = N4228 & en_i;
  assign N8000 = ~valid[942];
  assign match_array[943] = N8002 & valid[943];
  assign N8002 = N8001 & N4048;
  assign N8001 = N4228 & en_i;
  assign empty_array[943] = N8003 & N8004;
  assign N8003 = N4228 & en_i;
  assign N8004 = ~valid[943];
  assign match_array[944] = N8006 & valid[944];
  assign N8006 = N8005 & N4049;
  assign N8005 = N4228 & en_i;
  assign empty_array[944] = N8007 & N8008;
  assign N8007 = N4228 & en_i;
  assign N8008 = ~valid[944];
  assign match_array[945] = N8010 & valid[945];
  assign N8010 = N8009 & N4050;
  assign N8009 = N4228 & en_i;
  assign empty_array[945] = N8011 & N8012;
  assign N8011 = N4228 & en_i;
  assign N8012 = ~valid[945];
  assign match_array[946] = N8014 & valid[946];
  assign N8014 = N8013 & N4051;
  assign N8013 = N4228 & en_i;
  assign empty_array[946] = N8015 & N8016;
  assign N8015 = N4228 & en_i;
  assign N8016 = ~valid[946];
  assign match_array[947] = N8018 & valid[947];
  assign N8018 = N8017 & N4052;
  assign N8017 = N4228 & en_i;
  assign empty_array[947] = N8019 & N8020;
  assign N8019 = N4228 & en_i;
  assign N8020 = ~valid[947];
  assign match_array[948] = N8022 & valid[948];
  assign N8022 = N8021 & N4053;
  assign N8021 = N4228 & en_i;
  assign empty_array[948] = N8023 & N8024;
  assign N8023 = N4228 & en_i;
  assign N8024 = ~valid[948];
  assign match_array[949] = N8026 & valid[949];
  assign N8026 = N8025 & N4054;
  assign N8025 = N4228 & en_i;
  assign empty_array[949] = N8027 & N8028;
  assign N8027 = N4228 & en_i;
  assign N8028 = ~valid[949];
  assign match_array[950] = N8030 & valid[950];
  assign N8030 = N8029 & N4055;
  assign N8029 = N4228 & en_i;
  assign empty_array[950] = N8031 & N8032;
  assign N8031 = N4228 & en_i;
  assign N8032 = ~valid[950];
  assign match_array[951] = N8034 & valid[951];
  assign N8034 = N8033 & N4056;
  assign N8033 = N4228 & en_i;
  assign empty_array[951] = N8035 & N8036;
  assign N8035 = N4228 & en_i;
  assign N8036 = ~valid[951];
  assign match_array[952] = N8038 & valid[952];
  assign N8038 = N8037 & N4057;
  assign N8037 = N4228 & en_i;
  assign empty_array[952] = N8039 & N8040;
  assign N8039 = N4228 & en_i;
  assign N8040 = ~valid[952];
  assign match_array[953] = N8042 & valid[953];
  assign N8042 = N8041 & N4058;
  assign N8041 = N4228 & en_i;
  assign empty_array[953] = N8043 & N8044;
  assign N8043 = N4228 & en_i;
  assign N8044 = ~valid[953];
  assign match_array[954] = N8046 & valid[954];
  assign N8046 = N8045 & N4059;
  assign N8045 = N4228 & en_i;
  assign empty_array[954] = N8047 & N8048;
  assign N8047 = N4228 & en_i;
  assign N8048 = ~valid[954];
  assign match_array[955] = N8050 & valid[955];
  assign N8050 = N8049 & N4060;
  assign N8049 = N4228 & en_i;
  assign empty_array[955] = N8051 & N8052;
  assign N8051 = N4228 & en_i;
  assign N8052 = ~valid[955];
  assign match_array[956] = N8054 & valid[956];
  assign N8054 = N8053 & N4061;
  assign N8053 = N4228 & en_i;
  assign empty_array[956] = N8055 & N8056;
  assign N8055 = N4228 & en_i;
  assign N8056 = ~valid[956];
  assign match_array[957] = N8058 & valid[957];
  assign N8058 = N8057 & N4062;
  assign N8057 = N4228 & en_i;
  assign empty_array[957] = N8059 & N8060;
  assign N8059 = N4228 & en_i;
  assign N8060 = ~valid[957];
  assign match_array[958] = N8062 & valid[958];
  assign N8062 = N8061 & N4063;
  assign N8061 = N4228 & en_i;
  assign empty_array[958] = N8063 & N8064;
  assign N8063 = N4228 & en_i;
  assign N8064 = ~valid[958];
  assign match_array[959] = N8066 & valid[959];
  assign N8066 = N8065 & N4064;
  assign N8065 = N4228 & en_i;
  assign empty_array[959] = N8067 & N8068;
  assign N8067 = N4228 & en_i;
  assign N8068 = ~valid[959];
  assign match_array[960] = N8070 & valid[960];
  assign N8070 = N8069 & N4065;
  assign N8069 = N4228 & en_i;
  assign empty_array[960] = N8071 & N8072;
  assign N8071 = N4228 & en_i;
  assign N8072 = ~valid[960];
  assign match_array[961] = N8074 & valid[961];
  assign N8074 = N8073 & N4066;
  assign N8073 = N4228 & en_i;
  assign empty_array[961] = N8075 & N8076;
  assign N8075 = N4228 & en_i;
  assign N8076 = ~valid[961];
  assign match_array[962] = N8078 & valid[962];
  assign N8078 = N8077 & N4067;
  assign N8077 = N4228 & en_i;
  assign empty_array[962] = N8079 & N8080;
  assign N8079 = N4228 & en_i;
  assign N8080 = ~valid[962];
  assign match_array[963] = N8082 & valid[963];
  assign N8082 = N8081 & N4068;
  assign N8081 = N4228 & en_i;
  assign empty_array[963] = N8083 & N8084;
  assign N8083 = N4228 & en_i;
  assign N8084 = ~valid[963];
  assign match_array[964] = N8086 & valid[964];
  assign N8086 = N8085 & N4069;
  assign N8085 = N4228 & en_i;
  assign empty_array[964] = N8087 & N8088;
  assign N8087 = N4228 & en_i;
  assign N8088 = ~valid[964];
  assign match_array[965] = N8090 & valid[965];
  assign N8090 = N8089 & N4070;
  assign N8089 = N4228 & en_i;
  assign empty_array[965] = N8091 & N8092;
  assign N8091 = N4228 & en_i;
  assign N8092 = ~valid[965];
  assign match_array[966] = N8094 & valid[966];
  assign N8094 = N8093 & N4071;
  assign N8093 = N4228 & en_i;
  assign empty_array[966] = N8095 & N8096;
  assign N8095 = N4228 & en_i;
  assign N8096 = ~valid[966];
  assign match_array[967] = N8098 & valid[967];
  assign N8098 = N8097 & N4072;
  assign N8097 = N4228 & en_i;
  assign empty_array[967] = N8099 & N8100;
  assign N8099 = N4228 & en_i;
  assign N8100 = ~valid[967];
  assign match_array[968] = N8102 & valid[968];
  assign N8102 = N8101 & N4073;
  assign N8101 = N4228 & en_i;
  assign empty_array[968] = N8103 & N8104;
  assign N8103 = N4228 & en_i;
  assign N8104 = ~valid[968];
  assign match_array[969] = N8106 & valid[969];
  assign N8106 = N8105 & N4074;
  assign N8105 = N4228 & en_i;
  assign empty_array[969] = N8107 & N8108;
  assign N8107 = N4228 & en_i;
  assign N8108 = ~valid[969];
  assign match_array[970] = N8110 & valid[970];
  assign N8110 = N8109 & N4075;
  assign N8109 = N4228 & en_i;
  assign empty_array[970] = N8111 & N8112;
  assign N8111 = N4228 & en_i;
  assign N8112 = ~valid[970];
  assign match_array[971] = N8114 & valid[971];
  assign N8114 = N8113 & N4076;
  assign N8113 = N4228 & en_i;
  assign empty_array[971] = N8115 & N8116;
  assign N8115 = N4228 & en_i;
  assign N8116 = ~valid[971];
  assign match_array[972] = N8118 & valid[972];
  assign N8118 = N8117 & N4077;
  assign N8117 = N4228 & en_i;
  assign empty_array[972] = N8119 & N8120;
  assign N8119 = N4228 & en_i;
  assign N8120 = ~valid[972];
  assign match_array[973] = N8122 & valid[973];
  assign N8122 = N8121 & N4078;
  assign N8121 = N4228 & en_i;
  assign empty_array[973] = N8123 & N8124;
  assign N8123 = N4228 & en_i;
  assign N8124 = ~valid[973];
  assign match_array[974] = N8126 & valid[974];
  assign N8126 = N8125 & N4079;
  assign N8125 = N4228 & en_i;
  assign empty_array[974] = N8127 & N8128;
  assign N8127 = N4228 & en_i;
  assign N8128 = ~valid[974];
  assign match_array[975] = N8130 & valid[975];
  assign N8130 = N8129 & N4080;
  assign N8129 = N4228 & en_i;
  assign empty_array[975] = N8131 & N8132;
  assign N8131 = N4228 & en_i;
  assign N8132 = ~valid[975];
  assign match_array[976] = N8134 & valid[976];
  assign N8134 = N8133 & N4081;
  assign N8133 = N4228 & en_i;
  assign empty_array[976] = N8135 & N8136;
  assign N8135 = N4228 & en_i;
  assign N8136 = ~valid[976];
  assign match_array[977] = N8138 & valid[977];
  assign N8138 = N8137 & N4082;
  assign N8137 = N4228 & en_i;
  assign empty_array[977] = N8139 & N8140;
  assign N8139 = N4228 & en_i;
  assign N8140 = ~valid[977];
  assign match_array[978] = N8142 & valid[978];
  assign N8142 = N8141 & N4083;
  assign N8141 = N4228 & en_i;
  assign empty_array[978] = N8143 & N8144;
  assign N8143 = N4228 & en_i;
  assign N8144 = ~valid[978];
  assign match_array[979] = N8146 & valid[979];
  assign N8146 = N8145 & N4084;
  assign N8145 = N4228 & en_i;
  assign empty_array[979] = N8147 & N8148;
  assign N8147 = N4228 & en_i;
  assign N8148 = ~valid[979];
  assign match_array[980] = N8150 & valid[980];
  assign N8150 = N8149 & N4085;
  assign N8149 = N4228 & en_i;
  assign empty_array[980] = N8151 & N8152;
  assign N8151 = N4228 & en_i;
  assign N8152 = ~valid[980];
  assign match_array[981] = N8154 & valid[981];
  assign N8154 = N8153 & N4086;
  assign N8153 = N4228 & en_i;
  assign empty_array[981] = N8155 & N8156;
  assign N8155 = N4228 & en_i;
  assign N8156 = ~valid[981];
  assign match_array[982] = N8158 & valid[982];
  assign N8158 = N8157 & N4087;
  assign N8157 = N4228 & en_i;
  assign empty_array[982] = N8159 & N8160;
  assign N8159 = N4228 & en_i;
  assign N8160 = ~valid[982];
  assign match_array[983] = N8162 & valid[983];
  assign N8162 = N8161 & N4088;
  assign N8161 = N4228 & en_i;
  assign empty_array[983] = N8163 & N8164;
  assign N8163 = N4228 & en_i;
  assign N8164 = ~valid[983];
  assign match_array[984] = N8166 & valid[984];
  assign N8166 = N8165 & N4089;
  assign N8165 = N4228 & en_i;
  assign empty_array[984] = N8167 & N8168;
  assign N8167 = N4228 & en_i;
  assign N8168 = ~valid[984];
  assign match_array[985] = N8170 & valid[985];
  assign N8170 = N8169 & N4090;
  assign N8169 = N4228 & en_i;
  assign empty_array[985] = N8171 & N8172;
  assign N8171 = N4228 & en_i;
  assign N8172 = ~valid[985];
  assign match_array[986] = N8174 & valid[986];
  assign N8174 = N8173 & N4091;
  assign N8173 = N4228 & en_i;
  assign empty_array[986] = N8175 & N8176;
  assign N8175 = N4228 & en_i;
  assign N8176 = ~valid[986];
  assign match_array[987] = N8178 & valid[987];
  assign N8178 = N8177 & N4092;
  assign N8177 = N4228 & en_i;
  assign empty_array[987] = N8179 & N8180;
  assign N8179 = N4228 & en_i;
  assign N8180 = ~valid[987];
  assign match_array[988] = N8182 & valid[988];
  assign N8182 = N8181 & N4093;
  assign N8181 = N4228 & en_i;
  assign empty_array[988] = N8183 & N8184;
  assign N8183 = N4228 & en_i;
  assign N8184 = ~valid[988];
  assign match_array[989] = N8186 & valid[989];
  assign N8186 = N8185 & N4094;
  assign N8185 = N4228 & en_i;
  assign empty_array[989] = N8187 & N8188;
  assign N8187 = N4228 & en_i;
  assign N8188 = ~valid[989];
  assign match_array[990] = N8190 & valid[990];
  assign N8190 = N8189 & N4095;
  assign N8189 = N4228 & en_i;
  assign empty_array[990] = N8191 & N8192;
  assign N8191 = N4228 & en_i;
  assign N8192 = ~valid[990];
  assign match_array[991] = N8194 & valid[991];
  assign N8194 = N8193 & N4096;
  assign N8193 = N4228 & en_i;
  assign empty_array[991] = N8195 & N8196;
  assign N8195 = N4228 & en_i;
  assign N8196 = ~valid[991];
  assign match_array[992] = N8198 & valid[992];
  assign N8198 = N8197 & N4097;
  assign N8197 = N4228 & en_i;
  assign empty_array[992] = N8199 & N8200;
  assign N8199 = N4228 & en_i;
  assign N8200 = ~valid[992];
  assign match_array[993] = N8202 & valid[993];
  assign N8202 = N8201 & N4098;
  assign N8201 = N4228 & en_i;
  assign empty_array[993] = N8203 & N8204;
  assign N8203 = N4228 & en_i;
  assign N8204 = ~valid[993];
  assign match_array[994] = N8206 & valid[994];
  assign N8206 = N8205 & N4099;
  assign N8205 = N4228 & en_i;
  assign empty_array[994] = N8207 & N8208;
  assign N8207 = N4228 & en_i;
  assign N8208 = ~valid[994];
  assign match_array[995] = N8210 & valid[995];
  assign N8210 = N8209 & N4100;
  assign N8209 = N4228 & en_i;
  assign empty_array[995] = N8211 & N8212;
  assign N8211 = N4228 & en_i;
  assign N8212 = ~valid[995];
  assign match_array[996] = N8214 & valid[996];
  assign N8214 = N8213 & N4101;
  assign N8213 = N4228 & en_i;
  assign empty_array[996] = N8215 & N8216;
  assign N8215 = N4228 & en_i;
  assign N8216 = ~valid[996];
  assign match_array[997] = N8218 & valid[997];
  assign N8218 = N8217 & N4102;
  assign N8217 = N4228 & en_i;
  assign empty_array[997] = N8219 & N8220;
  assign N8219 = N4228 & en_i;
  assign N8220 = ~valid[997];
  assign match_array[998] = N8222 & valid[998];
  assign N8222 = N8221 & N4103;
  assign N8221 = N4228 & en_i;
  assign empty_array[998] = N8223 & N8224;
  assign N8223 = N4228 & en_i;
  assign N8224 = ~valid[998];
  assign match_array[999] = N8226 & valid[999];
  assign N8226 = N8225 & N4104;
  assign N8225 = N4228 & en_i;
  assign empty_array[999] = N8227 & N8228;
  assign N8227 = N4228 & en_i;
  assign N8228 = ~valid[999];
  assign match_array[1000] = N8230 & valid[1000];
  assign N8230 = N8229 & N4105;
  assign N8229 = N4228 & en_i;
  assign empty_array[1000] = N8231 & N8232;
  assign N8231 = N4228 & en_i;
  assign N8232 = ~valid[1000];
  assign match_array[1001] = N8234 & valid[1001];
  assign N8234 = N8233 & N4106;
  assign N8233 = N4228 & en_i;
  assign empty_array[1001] = N8235 & N8236;
  assign N8235 = N4228 & en_i;
  assign N8236 = ~valid[1001];
  assign match_array[1002] = N8238 & valid[1002];
  assign N8238 = N8237 & N4107;
  assign N8237 = N4228 & en_i;
  assign empty_array[1002] = N8239 & N8240;
  assign N8239 = N4228 & en_i;
  assign N8240 = ~valid[1002];
  assign match_array[1003] = N8242 & valid[1003];
  assign N8242 = N8241 & N4108;
  assign N8241 = N4228 & en_i;
  assign empty_array[1003] = N8243 & N8244;
  assign N8243 = N4228 & en_i;
  assign N8244 = ~valid[1003];
  assign match_array[1004] = N8246 & valid[1004];
  assign N8246 = N8245 & N4109;
  assign N8245 = N4228 & en_i;
  assign empty_array[1004] = N8247 & N8248;
  assign N8247 = N4228 & en_i;
  assign N8248 = ~valid[1004];
  assign match_array[1005] = N8250 & valid[1005];
  assign N8250 = N8249 & N4110;
  assign N8249 = N4228 & en_i;
  assign empty_array[1005] = N8251 & N8252;
  assign N8251 = N4228 & en_i;
  assign N8252 = ~valid[1005];
  assign match_array[1006] = N8254 & valid[1006];
  assign N8254 = N8253 & N4111;
  assign N8253 = N4228 & en_i;
  assign empty_array[1006] = N8255 & N8256;
  assign N8255 = N4228 & en_i;
  assign N8256 = ~valid[1006];
  assign match_array[1007] = N8258 & valid[1007];
  assign N8258 = N8257 & N4112;
  assign N8257 = N4228 & en_i;
  assign empty_array[1007] = N8259 & N8260;
  assign N8259 = N4228 & en_i;
  assign N8260 = ~valid[1007];
  assign match_array[1008] = N8262 & valid[1008];
  assign N8262 = N8261 & N4113;
  assign N8261 = N4228 & en_i;
  assign empty_array[1008] = N8263 & N8264;
  assign N8263 = N4228 & en_i;
  assign N8264 = ~valid[1008];
  assign match_array[1009] = N8266 & valid[1009];
  assign N8266 = N8265 & N4114;
  assign N8265 = N4228 & en_i;
  assign empty_array[1009] = N8267 & N8268;
  assign N8267 = N4228 & en_i;
  assign N8268 = ~valid[1009];
  assign match_array[1010] = N8270 & valid[1010];
  assign N8270 = N8269 & N4115;
  assign N8269 = N4228 & en_i;
  assign empty_array[1010] = N8271 & N8272;
  assign N8271 = N4228 & en_i;
  assign N8272 = ~valid[1010];
  assign match_array[1011] = N8274 & valid[1011];
  assign N8274 = N8273 & N4116;
  assign N8273 = N4228 & en_i;
  assign empty_array[1011] = N8275 & N8276;
  assign N8275 = N4228 & en_i;
  assign N8276 = ~valid[1011];
  assign match_array[1012] = N8278 & valid[1012];
  assign N8278 = N8277 & N4117;
  assign N8277 = N4228 & en_i;
  assign empty_array[1012] = N8279 & N8280;
  assign N8279 = N4228 & en_i;
  assign N8280 = ~valid[1012];
  assign match_array[1013] = N8282 & valid[1013];
  assign N8282 = N8281 & N4118;
  assign N8281 = N4228 & en_i;
  assign empty_array[1013] = N8283 & N8284;
  assign N8283 = N4228 & en_i;
  assign N8284 = ~valid[1013];
  assign match_array[1014] = N8286 & valid[1014];
  assign N8286 = N8285 & N4119;
  assign N8285 = N4228 & en_i;
  assign empty_array[1014] = N8287 & N8288;
  assign N8287 = N4228 & en_i;
  assign N8288 = ~valid[1014];
  assign match_array[1015] = N8290 & valid[1015];
  assign N8290 = N8289 & N4120;
  assign N8289 = N4228 & en_i;
  assign empty_array[1015] = N8291 & N8292;
  assign N8291 = N4228 & en_i;
  assign N8292 = ~valid[1015];
  assign match_array[1016] = N8294 & valid[1016];
  assign N8294 = N8293 & N4121;
  assign N8293 = N4228 & en_i;
  assign empty_array[1016] = N8295 & N8296;
  assign N8295 = N4228 & en_i;
  assign N8296 = ~valid[1016];
  assign match_array[1017] = N8298 & valid[1017];
  assign N8298 = N8297 & N4122;
  assign N8297 = N4228 & en_i;
  assign empty_array[1017] = N8299 & N8300;
  assign N8299 = N4228 & en_i;
  assign N8300 = ~valid[1017];
  assign match_array[1018] = N8302 & valid[1018];
  assign N8302 = N8301 & N4123;
  assign N8301 = N4228 & en_i;
  assign empty_array[1018] = N8303 & N8304;
  assign N8303 = N4228 & en_i;
  assign N8304 = ~valid[1018];
  assign match_array[1019] = N8306 & valid[1019];
  assign N8306 = N8305 & N4124;
  assign N8305 = N4228 & en_i;
  assign empty_array[1019] = N8307 & N8308;
  assign N8307 = N4228 & en_i;
  assign N8308 = ~valid[1019];
  assign match_array[1020] = N8310 & valid[1020];
  assign N8310 = N8309 & N4125;
  assign N8309 = N4228 & en_i;
  assign empty_array[1020] = N8311 & N8312;
  assign N8311 = N4228 & en_i;
  assign N8312 = ~valid[1020];
  assign match_array[1021] = N8314 & valid[1021];
  assign N8314 = N8313 & N4126;
  assign N8313 = N4228 & en_i;
  assign empty_array[1021] = N8315 & N8316;
  assign N8315 = N4228 & en_i;
  assign N8316 = ~valid[1021];
  assign match_array[1022] = N8318 & valid[1022];
  assign N8318 = N8317 & N4127;
  assign N8317 = N4228 & en_i;
  assign empty_array[1022] = N8319 & N8320;
  assign N8319 = N4228 & en_i;
  assign N8320 = ~valid[1022];
  assign match_array[1023] = N8322 & valid[1023];
  assign N8322 = N8321 & N4128;
  assign N8321 = N4228 & en_i;
  assign empty_array[1023] = N8323 & N8324;
  assign N8323 = N4228 & en_i;
  assign N8324 = ~valid[1023];

  always @(posedge clk_i) begin
    if(N3102) begin
      { mem[32767:32736] } <= { w_data_i[31:0] };
    end 
    if(N3101) begin
      { mem[32735:32704] } <= { w_data_i[31:0] };
    end 
    if(N3100) begin
      { mem[32703:32672] } <= { w_data_i[31:0] };
    end 
    if(N3099) begin
      { mem[32671:32640] } <= { w_data_i[31:0] };
    end 
    if(N3098) begin
      { mem[32639:32608] } <= { w_data_i[31:0] };
    end 
    if(N3097) begin
      { mem[32607:32576] } <= { w_data_i[31:0] };
    end 
    if(N3096) begin
      { mem[32575:32544] } <= { w_data_i[31:0] };
    end 
    if(N3095) begin
      { mem[32543:32512] } <= { w_data_i[31:0] };
    end 
    if(N3094) begin
      { mem[32511:32480] } <= { w_data_i[31:0] };
    end 
    if(N3093) begin
      { mem[32479:32448] } <= { w_data_i[31:0] };
    end 
    if(N3092) begin
      { mem[32447:32416] } <= { w_data_i[31:0] };
    end 
    if(N3091) begin
      { mem[32415:32384] } <= { w_data_i[31:0] };
    end 
    if(N3090) begin
      { mem[32383:32352] } <= { w_data_i[31:0] };
    end 
    if(N3089) begin
      { mem[32351:32320] } <= { w_data_i[31:0] };
    end 
    if(N3088) begin
      { mem[32319:32288] } <= { w_data_i[31:0] };
    end 
    if(N3087) begin
      { mem[32287:32256] } <= { w_data_i[31:0] };
    end 
    if(N3086) begin
      { mem[32255:32224] } <= { w_data_i[31:0] };
    end 
    if(N3085) begin
      { mem[32223:32192] } <= { w_data_i[31:0] };
    end 
    if(N3084) begin
      { mem[32191:32160] } <= { w_data_i[31:0] };
    end 
    if(N3083) begin
      { mem[32159:32128] } <= { w_data_i[31:0] };
    end 
    if(N3082) begin
      { mem[32127:32096] } <= { w_data_i[31:0] };
    end 
    if(N3081) begin
      { mem[32095:32064] } <= { w_data_i[31:0] };
    end 
    if(N3080) begin
      { mem[32063:32032] } <= { w_data_i[31:0] };
    end 
    if(N3079) begin
      { mem[32031:32000] } <= { w_data_i[31:0] };
    end 
    if(N3078) begin
      { mem[31999:31968] } <= { w_data_i[31:0] };
    end 
    if(N3077) begin
      { mem[31967:31936] } <= { w_data_i[31:0] };
    end 
    if(N3076) begin
      { mem[31935:31904] } <= { w_data_i[31:0] };
    end 
    if(N3075) begin
      { mem[31903:31872] } <= { w_data_i[31:0] };
    end 
    if(N3074) begin
      { mem[31871:31840] } <= { w_data_i[31:0] };
    end 
    if(N3073) begin
      { mem[31839:31808] } <= { w_data_i[31:0] };
    end 
    if(N3072) begin
      { mem[31807:31776] } <= { w_data_i[31:0] };
    end 
    if(N3071) begin
      { mem[31775:31744] } <= { w_data_i[31:0] };
    end 
    if(N3070) begin
      { mem[31743:31712] } <= { w_data_i[31:0] };
    end 
    if(N3069) begin
      { mem[31711:31680] } <= { w_data_i[31:0] };
    end 
    if(N3068) begin
      { mem[31679:31648] } <= { w_data_i[31:0] };
    end 
    if(N3067) begin
      { mem[31647:31616] } <= { w_data_i[31:0] };
    end 
    if(N3066) begin
      { mem[31615:31584] } <= { w_data_i[31:0] };
    end 
    if(N3065) begin
      { mem[31583:31552] } <= { w_data_i[31:0] };
    end 
    if(N3064) begin
      { mem[31551:31520] } <= { w_data_i[31:0] };
    end 
    if(N3063) begin
      { mem[31519:31488] } <= { w_data_i[31:0] };
    end 
    if(N3062) begin
      { mem[31487:31456] } <= { w_data_i[31:0] };
    end 
    if(N3061) begin
      { mem[31455:31424] } <= { w_data_i[31:0] };
    end 
    if(N3060) begin
      { mem[31423:31392] } <= { w_data_i[31:0] };
    end 
    if(N3059) begin
      { mem[31391:31360] } <= { w_data_i[31:0] };
    end 
    if(N3058) begin
      { mem[31359:31328] } <= { w_data_i[31:0] };
    end 
    if(N3057) begin
      { mem[31327:31296] } <= { w_data_i[31:0] };
    end 
    if(N3056) begin
      { mem[31295:31264] } <= { w_data_i[31:0] };
    end 
    if(N3055) begin
      { mem[31263:31232] } <= { w_data_i[31:0] };
    end 
    if(N3054) begin
      { mem[31231:31200] } <= { w_data_i[31:0] };
    end 
    if(N3053) begin
      { mem[31199:31168] } <= { w_data_i[31:0] };
    end 
    if(N3052) begin
      { mem[31167:31136] } <= { w_data_i[31:0] };
    end 
    if(N3051) begin
      { mem[31135:31104] } <= { w_data_i[31:0] };
    end 
    if(N3050) begin
      { mem[31103:31072] } <= { w_data_i[31:0] };
    end 
    if(N3049) begin
      { mem[31071:31040] } <= { w_data_i[31:0] };
    end 
    if(N3048) begin
      { mem[31039:31008] } <= { w_data_i[31:0] };
    end 
    if(N3047) begin
      { mem[31007:30976] } <= { w_data_i[31:0] };
    end 
    if(N3046) begin
      { mem[30975:30944] } <= { w_data_i[31:0] };
    end 
    if(N3045) begin
      { mem[30943:30912] } <= { w_data_i[31:0] };
    end 
    if(N3044) begin
      { mem[30911:30880] } <= { w_data_i[31:0] };
    end 
    if(N3043) begin
      { mem[30879:30848] } <= { w_data_i[31:0] };
    end 
    if(N3042) begin
      { mem[30847:30816] } <= { w_data_i[31:0] };
    end 
    if(N3041) begin
      { mem[30815:30784] } <= { w_data_i[31:0] };
    end 
    if(N3040) begin
      { mem[30783:30752] } <= { w_data_i[31:0] };
    end 
    if(N3039) begin
      { mem[30751:30720] } <= { w_data_i[31:0] };
    end 
    if(N3038) begin
      { mem[30719:30688] } <= { w_data_i[31:0] };
    end 
    if(N3037) begin
      { mem[30687:30656] } <= { w_data_i[31:0] };
    end 
    if(N3036) begin
      { mem[30655:30624] } <= { w_data_i[31:0] };
    end 
    if(N3035) begin
      { mem[30623:30592] } <= { w_data_i[31:0] };
    end 
    if(N3034) begin
      { mem[30591:30560] } <= { w_data_i[31:0] };
    end 
    if(N3033) begin
      { mem[30559:30528] } <= { w_data_i[31:0] };
    end 
    if(N3032) begin
      { mem[30527:30496] } <= { w_data_i[31:0] };
    end 
    if(N3031) begin
      { mem[30495:30464] } <= { w_data_i[31:0] };
    end 
    if(N3030) begin
      { mem[30463:30432] } <= { w_data_i[31:0] };
    end 
    if(N3029) begin
      { mem[30431:30400] } <= { w_data_i[31:0] };
    end 
    if(N3028) begin
      { mem[30399:30368] } <= { w_data_i[31:0] };
    end 
    if(N3027) begin
      { mem[30367:30336] } <= { w_data_i[31:0] };
    end 
    if(N3026) begin
      { mem[30335:30304] } <= { w_data_i[31:0] };
    end 
    if(N3025) begin
      { mem[30303:30272] } <= { w_data_i[31:0] };
    end 
    if(N3024) begin
      { mem[30271:30240] } <= { w_data_i[31:0] };
    end 
    if(N3023) begin
      { mem[30239:30208] } <= { w_data_i[31:0] };
    end 
    if(N3022) begin
      { mem[30207:30176] } <= { w_data_i[31:0] };
    end 
    if(N3021) begin
      { mem[30175:30144] } <= { w_data_i[31:0] };
    end 
    if(N3020) begin
      { mem[30143:30112] } <= { w_data_i[31:0] };
    end 
    if(N3019) begin
      { mem[30111:30080] } <= { w_data_i[31:0] };
    end 
    if(N3018) begin
      { mem[30079:30048] } <= { w_data_i[31:0] };
    end 
    if(N3017) begin
      { mem[30047:30016] } <= { w_data_i[31:0] };
    end 
    if(N3016) begin
      { mem[30015:29984] } <= { w_data_i[31:0] };
    end 
    if(N3015) begin
      { mem[29983:29952] } <= { w_data_i[31:0] };
    end 
    if(N3014) begin
      { mem[29951:29920] } <= { w_data_i[31:0] };
    end 
    if(N3013) begin
      { mem[29919:29888] } <= { w_data_i[31:0] };
    end 
    if(N3012) begin
      { mem[29887:29856] } <= { w_data_i[31:0] };
    end 
    if(N3011) begin
      { mem[29855:29824] } <= { w_data_i[31:0] };
    end 
    if(N3010) begin
      { mem[29823:29792] } <= { w_data_i[31:0] };
    end 
    if(N3009) begin
      { mem[29791:29760] } <= { w_data_i[31:0] };
    end 
    if(N3008) begin
      { mem[29759:29728] } <= { w_data_i[31:0] };
    end 
    if(N3007) begin
      { mem[29727:29696] } <= { w_data_i[31:0] };
    end 
    if(N3006) begin
      { mem[29695:29664] } <= { w_data_i[31:0] };
    end 
    if(N3005) begin
      { mem[29663:29632] } <= { w_data_i[31:0] };
    end 
    if(N3004) begin
      { mem[29631:29600] } <= { w_data_i[31:0] };
    end 
    if(N3003) begin
      { mem[29599:29568] } <= { w_data_i[31:0] };
    end 
    if(N3002) begin
      { mem[29567:29536] } <= { w_data_i[31:0] };
    end 
    if(N3001) begin
      { mem[29535:29504] } <= { w_data_i[31:0] };
    end 
    if(N3000) begin
      { mem[29503:29472] } <= { w_data_i[31:0] };
    end 
    if(N2999) begin
      { mem[29471:29440] } <= { w_data_i[31:0] };
    end 
    if(N2998) begin
      { mem[29439:29408] } <= { w_data_i[31:0] };
    end 
    if(N2997) begin
      { mem[29407:29376] } <= { w_data_i[31:0] };
    end 
    if(N2996) begin
      { mem[29375:29344] } <= { w_data_i[31:0] };
    end 
    if(N2995) begin
      { mem[29343:29312] } <= { w_data_i[31:0] };
    end 
    if(N2994) begin
      { mem[29311:29280] } <= { w_data_i[31:0] };
    end 
    if(N2993) begin
      { mem[29279:29248] } <= { w_data_i[31:0] };
    end 
    if(N2992) begin
      { mem[29247:29216] } <= { w_data_i[31:0] };
    end 
    if(N2991) begin
      { mem[29215:29184] } <= { w_data_i[31:0] };
    end 
    if(N2990) begin
      { mem[29183:29152] } <= { w_data_i[31:0] };
    end 
    if(N2989) begin
      { mem[29151:29120] } <= { w_data_i[31:0] };
    end 
    if(N2988) begin
      { mem[29119:29088] } <= { w_data_i[31:0] };
    end 
    if(N2987) begin
      { mem[29087:29056] } <= { w_data_i[31:0] };
    end 
    if(N2986) begin
      { mem[29055:29024] } <= { w_data_i[31:0] };
    end 
    if(N2985) begin
      { mem[29023:28992] } <= { w_data_i[31:0] };
    end 
    if(N2984) begin
      { mem[28991:28960] } <= { w_data_i[31:0] };
    end 
    if(N2983) begin
      { mem[28959:28928] } <= { w_data_i[31:0] };
    end 
    if(N2982) begin
      { mem[28927:28896] } <= { w_data_i[31:0] };
    end 
    if(N2981) begin
      { mem[28895:28864] } <= { w_data_i[31:0] };
    end 
    if(N2980) begin
      { mem[28863:28832] } <= { w_data_i[31:0] };
    end 
    if(N2979) begin
      { mem[28831:28800] } <= { w_data_i[31:0] };
    end 
    if(N2978) begin
      { mem[28799:28768] } <= { w_data_i[31:0] };
    end 
    if(N2977) begin
      { mem[28767:28736] } <= { w_data_i[31:0] };
    end 
    if(N2976) begin
      { mem[28735:28704] } <= { w_data_i[31:0] };
    end 
    if(N2975) begin
      { mem[28703:28672] } <= { w_data_i[31:0] };
    end 
    if(N2974) begin
      { mem[28671:28640] } <= { w_data_i[31:0] };
    end 
    if(N2973) begin
      { mem[28639:28608] } <= { w_data_i[31:0] };
    end 
    if(N2972) begin
      { mem[28607:28576] } <= { w_data_i[31:0] };
    end 
    if(N2971) begin
      { mem[28575:28544] } <= { w_data_i[31:0] };
    end 
    if(N2970) begin
      { mem[28543:28512] } <= { w_data_i[31:0] };
    end 
    if(N2969) begin
      { mem[28511:28480] } <= { w_data_i[31:0] };
    end 
    if(N2968) begin
      { mem[28479:28448] } <= { w_data_i[31:0] };
    end 
    if(N2967) begin
      { mem[28447:28416] } <= { w_data_i[31:0] };
    end 
    if(N2966) begin
      { mem[28415:28384] } <= { w_data_i[31:0] };
    end 
    if(N2965) begin
      { mem[28383:28352] } <= { w_data_i[31:0] };
    end 
    if(N2964) begin
      { mem[28351:28320] } <= { w_data_i[31:0] };
    end 
    if(N2963) begin
      { mem[28319:28288] } <= { w_data_i[31:0] };
    end 
    if(N2962) begin
      { mem[28287:28256] } <= { w_data_i[31:0] };
    end 
    if(N2961) begin
      { mem[28255:28224] } <= { w_data_i[31:0] };
    end 
    if(N2960) begin
      { mem[28223:28192] } <= { w_data_i[31:0] };
    end 
    if(N2959) begin
      { mem[28191:28160] } <= { w_data_i[31:0] };
    end 
    if(N2958) begin
      { mem[28159:28128] } <= { w_data_i[31:0] };
    end 
    if(N2957) begin
      { mem[28127:28096] } <= { w_data_i[31:0] };
    end 
    if(N2956) begin
      { mem[28095:28064] } <= { w_data_i[31:0] };
    end 
    if(N2955) begin
      { mem[28063:28032] } <= { w_data_i[31:0] };
    end 
    if(N2954) begin
      { mem[28031:28000] } <= { w_data_i[31:0] };
    end 
    if(N2953) begin
      { mem[27999:27968] } <= { w_data_i[31:0] };
    end 
    if(N2952) begin
      { mem[27967:27936] } <= { w_data_i[31:0] };
    end 
    if(N2951) begin
      { mem[27935:27904] } <= { w_data_i[31:0] };
    end 
    if(N2950) begin
      { mem[27903:27872] } <= { w_data_i[31:0] };
    end 
    if(N2949) begin
      { mem[27871:27840] } <= { w_data_i[31:0] };
    end 
    if(N2948) begin
      { mem[27839:27808] } <= { w_data_i[31:0] };
    end 
    if(N2947) begin
      { mem[27807:27776] } <= { w_data_i[31:0] };
    end 
    if(N2946) begin
      { mem[27775:27744] } <= { w_data_i[31:0] };
    end 
    if(N2945) begin
      { mem[27743:27712] } <= { w_data_i[31:0] };
    end 
    if(N2944) begin
      { mem[27711:27680] } <= { w_data_i[31:0] };
    end 
    if(N2943) begin
      { mem[27679:27648] } <= { w_data_i[31:0] };
    end 
    if(N2942) begin
      { mem[27647:27616] } <= { w_data_i[31:0] };
    end 
    if(N2941) begin
      { mem[27615:27584] } <= { w_data_i[31:0] };
    end 
    if(N2940) begin
      { mem[27583:27552] } <= { w_data_i[31:0] };
    end 
    if(N2939) begin
      { mem[27551:27520] } <= { w_data_i[31:0] };
    end 
    if(N2938) begin
      { mem[27519:27488] } <= { w_data_i[31:0] };
    end 
    if(N2937) begin
      { mem[27487:27456] } <= { w_data_i[31:0] };
    end 
    if(N2936) begin
      { mem[27455:27424] } <= { w_data_i[31:0] };
    end 
    if(N2935) begin
      { mem[27423:27392] } <= { w_data_i[31:0] };
    end 
    if(N2934) begin
      { mem[27391:27360] } <= { w_data_i[31:0] };
    end 
    if(N2933) begin
      { mem[27359:27328] } <= { w_data_i[31:0] };
    end 
    if(N2932) begin
      { mem[27327:27296] } <= { w_data_i[31:0] };
    end 
    if(N2931) begin
      { mem[27295:27264] } <= { w_data_i[31:0] };
    end 
    if(N2930) begin
      { mem[27263:27232] } <= { w_data_i[31:0] };
    end 
    if(N2929) begin
      { mem[27231:27200] } <= { w_data_i[31:0] };
    end 
    if(N2928) begin
      { mem[27199:27168] } <= { w_data_i[31:0] };
    end 
    if(N2927) begin
      { mem[27167:27136] } <= { w_data_i[31:0] };
    end 
    if(N2926) begin
      { mem[27135:27104] } <= { w_data_i[31:0] };
    end 
    if(N2925) begin
      { mem[27103:27072] } <= { w_data_i[31:0] };
    end 
    if(N2924) begin
      { mem[27071:27040] } <= { w_data_i[31:0] };
    end 
    if(N2923) begin
      { mem[27039:27008] } <= { w_data_i[31:0] };
    end 
    if(N2922) begin
      { mem[27007:26976] } <= { w_data_i[31:0] };
    end 
    if(N2921) begin
      { mem[26975:26944] } <= { w_data_i[31:0] };
    end 
    if(N2920) begin
      { mem[26943:26912] } <= { w_data_i[31:0] };
    end 
    if(N2919) begin
      { mem[26911:26880] } <= { w_data_i[31:0] };
    end 
    if(N2918) begin
      { mem[26879:26848] } <= { w_data_i[31:0] };
    end 
    if(N2917) begin
      { mem[26847:26816] } <= { w_data_i[31:0] };
    end 
    if(N2916) begin
      { mem[26815:26784] } <= { w_data_i[31:0] };
    end 
    if(N2915) begin
      { mem[26783:26752] } <= { w_data_i[31:0] };
    end 
    if(N2914) begin
      { mem[26751:26720] } <= { w_data_i[31:0] };
    end 
    if(N2913) begin
      { mem[26719:26688] } <= { w_data_i[31:0] };
    end 
    if(N2912) begin
      { mem[26687:26656] } <= { w_data_i[31:0] };
    end 
    if(N2911) begin
      { mem[26655:26624] } <= { w_data_i[31:0] };
    end 
    if(N2910) begin
      { mem[26623:26592] } <= { w_data_i[31:0] };
    end 
    if(N2909) begin
      { mem[26591:26560] } <= { w_data_i[31:0] };
    end 
    if(N2908) begin
      { mem[26559:26528] } <= { w_data_i[31:0] };
    end 
    if(N2907) begin
      { mem[26527:26496] } <= { w_data_i[31:0] };
    end 
    if(N2906) begin
      { mem[26495:26464] } <= { w_data_i[31:0] };
    end 
    if(N2905) begin
      { mem[26463:26432] } <= { w_data_i[31:0] };
    end 
    if(N2904) begin
      { mem[26431:26400] } <= { w_data_i[31:0] };
    end 
    if(N2903) begin
      { mem[26399:26368] } <= { w_data_i[31:0] };
    end 
    if(N2902) begin
      { mem[26367:26336] } <= { w_data_i[31:0] };
    end 
    if(N2901) begin
      { mem[26335:26304] } <= { w_data_i[31:0] };
    end 
    if(N2900) begin
      { mem[26303:26272] } <= { w_data_i[31:0] };
    end 
    if(N2899) begin
      { mem[26271:26240] } <= { w_data_i[31:0] };
    end 
    if(N2898) begin
      { mem[26239:26208] } <= { w_data_i[31:0] };
    end 
    if(N2897) begin
      { mem[26207:26176] } <= { w_data_i[31:0] };
    end 
    if(N2896) begin
      { mem[26175:26144] } <= { w_data_i[31:0] };
    end 
    if(N2895) begin
      { mem[26143:26112] } <= { w_data_i[31:0] };
    end 
    if(N2894) begin
      { mem[26111:26080] } <= { w_data_i[31:0] };
    end 
    if(N2893) begin
      { mem[26079:26048] } <= { w_data_i[31:0] };
    end 
    if(N2892) begin
      { mem[26047:26016] } <= { w_data_i[31:0] };
    end 
    if(N2891) begin
      { mem[26015:25984] } <= { w_data_i[31:0] };
    end 
    if(N2890) begin
      { mem[25983:25952] } <= { w_data_i[31:0] };
    end 
    if(N2889) begin
      { mem[25951:25920] } <= { w_data_i[31:0] };
    end 
    if(N2888) begin
      { mem[25919:25888] } <= { w_data_i[31:0] };
    end 
    if(N2887) begin
      { mem[25887:25856] } <= { w_data_i[31:0] };
    end 
    if(N2886) begin
      { mem[25855:25824] } <= { w_data_i[31:0] };
    end 
    if(N2885) begin
      { mem[25823:25792] } <= { w_data_i[31:0] };
    end 
    if(N2884) begin
      { mem[25791:25760] } <= { w_data_i[31:0] };
    end 
    if(N2883) begin
      { mem[25759:25728] } <= { w_data_i[31:0] };
    end 
    if(N2882) begin
      { mem[25727:25696] } <= { w_data_i[31:0] };
    end 
    if(N2881) begin
      { mem[25695:25664] } <= { w_data_i[31:0] };
    end 
    if(N2880) begin
      { mem[25663:25632] } <= { w_data_i[31:0] };
    end 
    if(N2879) begin
      { mem[25631:25600] } <= { w_data_i[31:0] };
    end 
    if(N2878) begin
      { mem[25599:25568] } <= { w_data_i[31:0] };
    end 
    if(N2877) begin
      { mem[25567:25536] } <= { w_data_i[31:0] };
    end 
    if(N2876) begin
      { mem[25535:25504] } <= { w_data_i[31:0] };
    end 
    if(N2875) begin
      { mem[25503:25472] } <= { w_data_i[31:0] };
    end 
    if(N2874) begin
      { mem[25471:25440] } <= { w_data_i[31:0] };
    end 
    if(N2873) begin
      { mem[25439:25408] } <= { w_data_i[31:0] };
    end 
    if(N2872) begin
      { mem[25407:25376] } <= { w_data_i[31:0] };
    end 
    if(N2871) begin
      { mem[25375:25344] } <= { w_data_i[31:0] };
    end 
    if(N2870) begin
      { mem[25343:25312] } <= { w_data_i[31:0] };
    end 
    if(N2869) begin
      { mem[25311:25280] } <= { w_data_i[31:0] };
    end 
    if(N2868) begin
      { mem[25279:25248] } <= { w_data_i[31:0] };
    end 
    if(N2867) begin
      { mem[25247:25216] } <= { w_data_i[31:0] };
    end 
    if(N2866) begin
      { mem[25215:25184] } <= { w_data_i[31:0] };
    end 
    if(N2865) begin
      { mem[25183:25152] } <= { w_data_i[31:0] };
    end 
    if(N2864) begin
      { mem[25151:25120] } <= { w_data_i[31:0] };
    end 
    if(N2863) begin
      { mem[25119:25088] } <= { w_data_i[31:0] };
    end 
    if(N2862) begin
      { mem[25087:25056] } <= { w_data_i[31:0] };
    end 
    if(N2861) begin
      { mem[25055:25024] } <= { w_data_i[31:0] };
    end 
    if(N2860) begin
      { mem[25023:24992] } <= { w_data_i[31:0] };
    end 
    if(N2859) begin
      { mem[24991:24960] } <= { w_data_i[31:0] };
    end 
    if(N2858) begin
      { mem[24959:24928] } <= { w_data_i[31:0] };
    end 
    if(N2857) begin
      { mem[24927:24896] } <= { w_data_i[31:0] };
    end 
    if(N2856) begin
      { mem[24895:24864] } <= { w_data_i[31:0] };
    end 
    if(N2855) begin
      { mem[24863:24832] } <= { w_data_i[31:0] };
    end 
    if(N2854) begin
      { mem[24831:24800] } <= { w_data_i[31:0] };
    end 
    if(N2853) begin
      { mem[24799:24768] } <= { w_data_i[31:0] };
    end 
    if(N2852) begin
      { mem[24767:24736] } <= { w_data_i[31:0] };
    end 
    if(N2851) begin
      { mem[24735:24704] } <= { w_data_i[31:0] };
    end 
    if(N2850) begin
      { mem[24703:24672] } <= { w_data_i[31:0] };
    end 
    if(N2849) begin
      { mem[24671:24640] } <= { w_data_i[31:0] };
    end 
    if(N2848) begin
      { mem[24639:24608] } <= { w_data_i[31:0] };
    end 
    if(N2847) begin
      { mem[24607:24576] } <= { w_data_i[31:0] };
    end 
    if(N2846) begin
      { mem[24575:24544] } <= { w_data_i[31:0] };
    end 
    if(N2845) begin
      { mem[24543:24512] } <= { w_data_i[31:0] };
    end 
    if(N2844) begin
      { mem[24511:24480] } <= { w_data_i[31:0] };
    end 
    if(N2843) begin
      { mem[24479:24448] } <= { w_data_i[31:0] };
    end 
    if(N2842) begin
      { mem[24447:24416] } <= { w_data_i[31:0] };
    end 
    if(N2841) begin
      { mem[24415:24384] } <= { w_data_i[31:0] };
    end 
    if(N2840) begin
      { mem[24383:24352] } <= { w_data_i[31:0] };
    end 
    if(N2839) begin
      { mem[24351:24320] } <= { w_data_i[31:0] };
    end 
    if(N2838) begin
      { mem[24319:24288] } <= { w_data_i[31:0] };
    end 
    if(N2837) begin
      { mem[24287:24256] } <= { w_data_i[31:0] };
    end 
    if(N2836) begin
      { mem[24255:24224] } <= { w_data_i[31:0] };
    end 
    if(N2835) begin
      { mem[24223:24192] } <= { w_data_i[31:0] };
    end 
    if(N2834) begin
      { mem[24191:24160] } <= { w_data_i[31:0] };
    end 
    if(N2833) begin
      { mem[24159:24128] } <= { w_data_i[31:0] };
    end 
    if(N2832) begin
      { mem[24127:24096] } <= { w_data_i[31:0] };
    end 
    if(N2831) begin
      { mem[24095:24064] } <= { w_data_i[31:0] };
    end 
    if(N2830) begin
      { mem[24063:24032] } <= { w_data_i[31:0] };
    end 
    if(N2829) begin
      { mem[24031:24000] } <= { w_data_i[31:0] };
    end 
    if(N2828) begin
      { mem[23999:23968] } <= { w_data_i[31:0] };
    end 
    if(N2827) begin
      { mem[23967:23936] } <= { w_data_i[31:0] };
    end 
    if(N2826) begin
      { mem[23935:23904] } <= { w_data_i[31:0] };
    end 
    if(N2825) begin
      { mem[23903:23872] } <= { w_data_i[31:0] };
    end 
    if(N2824) begin
      { mem[23871:23840] } <= { w_data_i[31:0] };
    end 
    if(N2823) begin
      { mem[23839:23808] } <= { w_data_i[31:0] };
    end 
    if(N2822) begin
      { mem[23807:23776] } <= { w_data_i[31:0] };
    end 
    if(N2821) begin
      { mem[23775:23744] } <= { w_data_i[31:0] };
    end 
    if(N2820) begin
      { mem[23743:23712] } <= { w_data_i[31:0] };
    end 
    if(N2819) begin
      { mem[23711:23680] } <= { w_data_i[31:0] };
    end 
    if(N2818) begin
      { mem[23679:23648] } <= { w_data_i[31:0] };
    end 
    if(N2817) begin
      { mem[23647:23616] } <= { w_data_i[31:0] };
    end 
    if(N2816) begin
      { mem[23615:23584] } <= { w_data_i[31:0] };
    end 
    if(N2815) begin
      { mem[23583:23552] } <= { w_data_i[31:0] };
    end 
    if(N2814) begin
      { mem[23551:23520] } <= { w_data_i[31:0] };
    end 
    if(N2813) begin
      { mem[23519:23488] } <= { w_data_i[31:0] };
    end 
    if(N2812) begin
      { mem[23487:23456] } <= { w_data_i[31:0] };
    end 
    if(N2811) begin
      { mem[23455:23424] } <= { w_data_i[31:0] };
    end 
    if(N2810) begin
      { mem[23423:23392] } <= { w_data_i[31:0] };
    end 
    if(N2809) begin
      { mem[23391:23360] } <= { w_data_i[31:0] };
    end 
    if(N2808) begin
      { mem[23359:23328] } <= { w_data_i[31:0] };
    end 
    if(N2807) begin
      { mem[23327:23296] } <= { w_data_i[31:0] };
    end 
    if(N2806) begin
      { mem[23295:23264] } <= { w_data_i[31:0] };
    end 
    if(N2805) begin
      { mem[23263:23232] } <= { w_data_i[31:0] };
    end 
    if(N2804) begin
      { mem[23231:23200] } <= { w_data_i[31:0] };
    end 
    if(N2803) begin
      { mem[23199:23168] } <= { w_data_i[31:0] };
    end 
    if(N2802) begin
      { mem[23167:23136] } <= { w_data_i[31:0] };
    end 
    if(N2801) begin
      { mem[23135:23104] } <= { w_data_i[31:0] };
    end 
    if(N2800) begin
      { mem[23103:23072] } <= { w_data_i[31:0] };
    end 
    if(N2799) begin
      { mem[23071:23040] } <= { w_data_i[31:0] };
    end 
    if(N2798) begin
      { mem[23039:23008] } <= { w_data_i[31:0] };
    end 
    if(N2797) begin
      { mem[23007:22976] } <= { w_data_i[31:0] };
    end 
    if(N2796) begin
      { mem[22975:22944] } <= { w_data_i[31:0] };
    end 
    if(N2795) begin
      { mem[22943:22912] } <= { w_data_i[31:0] };
    end 
    if(N2794) begin
      { mem[22911:22880] } <= { w_data_i[31:0] };
    end 
    if(N2793) begin
      { mem[22879:22848] } <= { w_data_i[31:0] };
    end 
    if(N2792) begin
      { mem[22847:22816] } <= { w_data_i[31:0] };
    end 
    if(N2791) begin
      { mem[22815:22784] } <= { w_data_i[31:0] };
    end 
    if(N2790) begin
      { mem[22783:22752] } <= { w_data_i[31:0] };
    end 
    if(N2789) begin
      { mem[22751:22720] } <= { w_data_i[31:0] };
    end 
    if(N2788) begin
      { mem[22719:22688] } <= { w_data_i[31:0] };
    end 
    if(N2787) begin
      { mem[22687:22656] } <= { w_data_i[31:0] };
    end 
    if(N2786) begin
      { mem[22655:22624] } <= { w_data_i[31:0] };
    end 
    if(N2785) begin
      { mem[22623:22592] } <= { w_data_i[31:0] };
    end 
    if(N2784) begin
      { mem[22591:22560] } <= { w_data_i[31:0] };
    end 
    if(N2783) begin
      { mem[22559:22528] } <= { w_data_i[31:0] };
    end 
    if(N2782) begin
      { mem[22527:22496] } <= { w_data_i[31:0] };
    end 
    if(N2781) begin
      { mem[22495:22464] } <= { w_data_i[31:0] };
    end 
    if(N2780) begin
      { mem[22463:22432] } <= { w_data_i[31:0] };
    end 
    if(N2779) begin
      { mem[22431:22400] } <= { w_data_i[31:0] };
    end 
    if(N2778) begin
      { mem[22399:22368] } <= { w_data_i[31:0] };
    end 
    if(N2777) begin
      { mem[22367:22336] } <= { w_data_i[31:0] };
    end 
    if(N2776) begin
      { mem[22335:22304] } <= { w_data_i[31:0] };
    end 
    if(N2775) begin
      { mem[22303:22272] } <= { w_data_i[31:0] };
    end 
    if(N2774) begin
      { mem[22271:22240] } <= { w_data_i[31:0] };
    end 
    if(N2773) begin
      { mem[22239:22208] } <= { w_data_i[31:0] };
    end 
    if(N2772) begin
      { mem[22207:22176] } <= { w_data_i[31:0] };
    end 
    if(N2771) begin
      { mem[22175:22144] } <= { w_data_i[31:0] };
    end 
    if(N2770) begin
      { mem[22143:22112] } <= { w_data_i[31:0] };
    end 
    if(N2769) begin
      { mem[22111:22080] } <= { w_data_i[31:0] };
    end 
    if(N2768) begin
      { mem[22079:22048] } <= { w_data_i[31:0] };
    end 
    if(N2767) begin
      { mem[22047:22016] } <= { w_data_i[31:0] };
    end 
    if(N2766) begin
      { mem[22015:21984] } <= { w_data_i[31:0] };
    end 
    if(N2765) begin
      { mem[21983:21952] } <= { w_data_i[31:0] };
    end 
    if(N2764) begin
      { mem[21951:21920] } <= { w_data_i[31:0] };
    end 
    if(N2763) begin
      { mem[21919:21888] } <= { w_data_i[31:0] };
    end 
    if(N2762) begin
      { mem[21887:21856] } <= { w_data_i[31:0] };
    end 
    if(N2761) begin
      { mem[21855:21824] } <= { w_data_i[31:0] };
    end 
    if(N2760) begin
      { mem[21823:21792] } <= { w_data_i[31:0] };
    end 
    if(N2759) begin
      { mem[21791:21760] } <= { w_data_i[31:0] };
    end 
    if(N2758) begin
      { mem[21759:21728] } <= { w_data_i[31:0] };
    end 
    if(N2757) begin
      { mem[21727:21696] } <= { w_data_i[31:0] };
    end 
    if(N2756) begin
      { mem[21695:21664] } <= { w_data_i[31:0] };
    end 
    if(N2755) begin
      { mem[21663:21632] } <= { w_data_i[31:0] };
    end 
    if(N2754) begin
      { mem[21631:21600] } <= { w_data_i[31:0] };
    end 
    if(N2753) begin
      { mem[21599:21568] } <= { w_data_i[31:0] };
    end 
    if(N2752) begin
      { mem[21567:21536] } <= { w_data_i[31:0] };
    end 
    if(N2751) begin
      { mem[21535:21504] } <= { w_data_i[31:0] };
    end 
    if(N2750) begin
      { mem[21503:21472] } <= { w_data_i[31:0] };
    end 
    if(N2749) begin
      { mem[21471:21440] } <= { w_data_i[31:0] };
    end 
    if(N2748) begin
      { mem[21439:21408] } <= { w_data_i[31:0] };
    end 
    if(N2747) begin
      { mem[21407:21376] } <= { w_data_i[31:0] };
    end 
    if(N2746) begin
      { mem[21375:21344] } <= { w_data_i[31:0] };
    end 
    if(N2745) begin
      { mem[21343:21312] } <= { w_data_i[31:0] };
    end 
    if(N2744) begin
      { mem[21311:21280] } <= { w_data_i[31:0] };
    end 
    if(N2743) begin
      { mem[21279:21248] } <= { w_data_i[31:0] };
    end 
    if(N2742) begin
      { mem[21247:21216] } <= { w_data_i[31:0] };
    end 
    if(N2741) begin
      { mem[21215:21184] } <= { w_data_i[31:0] };
    end 
    if(N2740) begin
      { mem[21183:21152] } <= { w_data_i[31:0] };
    end 
    if(N2739) begin
      { mem[21151:21120] } <= { w_data_i[31:0] };
    end 
    if(N2738) begin
      { mem[21119:21088] } <= { w_data_i[31:0] };
    end 
    if(N2737) begin
      { mem[21087:21056] } <= { w_data_i[31:0] };
    end 
    if(N2736) begin
      { mem[21055:21024] } <= { w_data_i[31:0] };
    end 
    if(N2735) begin
      { mem[21023:20992] } <= { w_data_i[31:0] };
    end 
    if(N2734) begin
      { mem[20991:20960] } <= { w_data_i[31:0] };
    end 
    if(N2733) begin
      { mem[20959:20928] } <= { w_data_i[31:0] };
    end 
    if(N2732) begin
      { mem[20927:20896] } <= { w_data_i[31:0] };
    end 
    if(N2731) begin
      { mem[20895:20864] } <= { w_data_i[31:0] };
    end 
    if(N2730) begin
      { mem[20863:20832] } <= { w_data_i[31:0] };
    end 
    if(N2729) begin
      { mem[20831:20800] } <= { w_data_i[31:0] };
    end 
    if(N2728) begin
      { mem[20799:20768] } <= { w_data_i[31:0] };
    end 
    if(N2727) begin
      { mem[20767:20736] } <= { w_data_i[31:0] };
    end 
    if(N2726) begin
      { mem[20735:20704] } <= { w_data_i[31:0] };
    end 
    if(N2725) begin
      { mem[20703:20672] } <= { w_data_i[31:0] };
    end 
    if(N2724) begin
      { mem[20671:20640] } <= { w_data_i[31:0] };
    end 
    if(N2723) begin
      { mem[20639:20608] } <= { w_data_i[31:0] };
    end 
    if(N2722) begin
      { mem[20607:20576] } <= { w_data_i[31:0] };
    end 
    if(N2721) begin
      { mem[20575:20544] } <= { w_data_i[31:0] };
    end 
    if(N2720) begin
      { mem[20543:20512] } <= { w_data_i[31:0] };
    end 
    if(N2719) begin
      { mem[20511:20480] } <= { w_data_i[31:0] };
    end 
    if(N2718) begin
      { mem[20479:20448] } <= { w_data_i[31:0] };
    end 
    if(N2717) begin
      { mem[20447:20416] } <= { w_data_i[31:0] };
    end 
    if(N2716) begin
      { mem[20415:20384] } <= { w_data_i[31:0] };
    end 
    if(N2715) begin
      { mem[20383:20352] } <= { w_data_i[31:0] };
    end 
    if(N2714) begin
      { mem[20351:20320] } <= { w_data_i[31:0] };
    end 
    if(N2713) begin
      { mem[20319:20288] } <= { w_data_i[31:0] };
    end 
    if(N2712) begin
      { mem[20287:20256] } <= { w_data_i[31:0] };
    end 
    if(N2711) begin
      { mem[20255:20224] } <= { w_data_i[31:0] };
    end 
    if(N2710) begin
      { mem[20223:20192] } <= { w_data_i[31:0] };
    end 
    if(N2709) begin
      { mem[20191:20160] } <= { w_data_i[31:0] };
    end 
    if(N2708) begin
      { mem[20159:20128] } <= { w_data_i[31:0] };
    end 
    if(N2707) begin
      { mem[20127:20096] } <= { w_data_i[31:0] };
    end 
    if(N2706) begin
      { mem[20095:20064] } <= { w_data_i[31:0] };
    end 
    if(N2705) begin
      { mem[20063:20032] } <= { w_data_i[31:0] };
    end 
    if(N2704) begin
      { mem[20031:20000] } <= { w_data_i[31:0] };
    end 
    if(N2703) begin
      { mem[19999:19968] } <= { w_data_i[31:0] };
    end 
    if(N2702) begin
      { mem[19967:19936] } <= { w_data_i[31:0] };
    end 
    if(N2701) begin
      { mem[19935:19904] } <= { w_data_i[31:0] };
    end 
    if(N2700) begin
      { mem[19903:19872] } <= { w_data_i[31:0] };
    end 
    if(N2699) begin
      { mem[19871:19840] } <= { w_data_i[31:0] };
    end 
    if(N2698) begin
      { mem[19839:19808] } <= { w_data_i[31:0] };
    end 
    if(N2697) begin
      { mem[19807:19776] } <= { w_data_i[31:0] };
    end 
    if(N2696) begin
      { mem[19775:19744] } <= { w_data_i[31:0] };
    end 
    if(N2695) begin
      { mem[19743:19712] } <= { w_data_i[31:0] };
    end 
    if(N2694) begin
      { mem[19711:19680] } <= { w_data_i[31:0] };
    end 
    if(N2693) begin
      { mem[19679:19648] } <= { w_data_i[31:0] };
    end 
    if(N2692) begin
      { mem[19647:19616] } <= { w_data_i[31:0] };
    end 
    if(N2691) begin
      { mem[19615:19584] } <= { w_data_i[31:0] };
    end 
    if(N2690) begin
      { mem[19583:19552] } <= { w_data_i[31:0] };
    end 
    if(N2689) begin
      { mem[19551:19520] } <= { w_data_i[31:0] };
    end 
    if(N2688) begin
      { mem[19519:19488] } <= { w_data_i[31:0] };
    end 
    if(N2687) begin
      { mem[19487:19456] } <= { w_data_i[31:0] };
    end 
    if(N2686) begin
      { mem[19455:19424] } <= { w_data_i[31:0] };
    end 
    if(N2685) begin
      { mem[19423:19392] } <= { w_data_i[31:0] };
    end 
    if(N2684) begin
      { mem[19391:19360] } <= { w_data_i[31:0] };
    end 
    if(N2683) begin
      { mem[19359:19328] } <= { w_data_i[31:0] };
    end 
    if(N2682) begin
      { mem[19327:19296] } <= { w_data_i[31:0] };
    end 
    if(N2681) begin
      { mem[19295:19264] } <= { w_data_i[31:0] };
    end 
    if(N2680) begin
      { mem[19263:19232] } <= { w_data_i[31:0] };
    end 
    if(N2679) begin
      { mem[19231:19200] } <= { w_data_i[31:0] };
    end 
    if(N2678) begin
      { mem[19199:19168] } <= { w_data_i[31:0] };
    end 
    if(N2677) begin
      { mem[19167:19136] } <= { w_data_i[31:0] };
    end 
    if(N2676) begin
      { mem[19135:19104] } <= { w_data_i[31:0] };
    end 
    if(N2675) begin
      { mem[19103:19072] } <= { w_data_i[31:0] };
    end 
    if(N2674) begin
      { mem[19071:19040] } <= { w_data_i[31:0] };
    end 
    if(N2673) begin
      { mem[19039:19008] } <= { w_data_i[31:0] };
    end 
    if(N2672) begin
      { mem[19007:18976] } <= { w_data_i[31:0] };
    end 
    if(N2671) begin
      { mem[18975:18944] } <= { w_data_i[31:0] };
    end 
    if(N2670) begin
      { mem[18943:18912] } <= { w_data_i[31:0] };
    end 
    if(N2669) begin
      { mem[18911:18880] } <= { w_data_i[31:0] };
    end 
    if(N2668) begin
      { mem[18879:18848] } <= { w_data_i[31:0] };
    end 
    if(N2667) begin
      { mem[18847:18816] } <= { w_data_i[31:0] };
    end 
    if(N2666) begin
      { mem[18815:18784] } <= { w_data_i[31:0] };
    end 
    if(N2665) begin
      { mem[18783:18752] } <= { w_data_i[31:0] };
    end 
    if(N2664) begin
      { mem[18751:18720] } <= { w_data_i[31:0] };
    end 
    if(N2663) begin
      { mem[18719:18688] } <= { w_data_i[31:0] };
    end 
    if(N2662) begin
      { mem[18687:18656] } <= { w_data_i[31:0] };
    end 
    if(N2661) begin
      { mem[18655:18624] } <= { w_data_i[31:0] };
    end 
    if(N2660) begin
      { mem[18623:18592] } <= { w_data_i[31:0] };
    end 
    if(N2659) begin
      { mem[18591:18560] } <= { w_data_i[31:0] };
    end 
    if(N2658) begin
      { mem[18559:18528] } <= { w_data_i[31:0] };
    end 
    if(N2657) begin
      { mem[18527:18496] } <= { w_data_i[31:0] };
    end 
    if(N2656) begin
      { mem[18495:18464] } <= { w_data_i[31:0] };
    end 
    if(N2655) begin
      { mem[18463:18432] } <= { w_data_i[31:0] };
    end 
    if(N2654) begin
      { mem[18431:18400] } <= { w_data_i[31:0] };
    end 
    if(N2653) begin
      { mem[18399:18368] } <= { w_data_i[31:0] };
    end 
    if(N2652) begin
      { mem[18367:18336] } <= { w_data_i[31:0] };
    end 
    if(N2651) begin
      { mem[18335:18304] } <= { w_data_i[31:0] };
    end 
    if(N2650) begin
      { mem[18303:18272] } <= { w_data_i[31:0] };
    end 
    if(N2649) begin
      { mem[18271:18240] } <= { w_data_i[31:0] };
    end 
    if(N2648) begin
      { mem[18239:18208] } <= { w_data_i[31:0] };
    end 
    if(N2647) begin
      { mem[18207:18176] } <= { w_data_i[31:0] };
    end 
    if(N2646) begin
      { mem[18175:18144] } <= { w_data_i[31:0] };
    end 
    if(N2645) begin
      { mem[18143:18112] } <= { w_data_i[31:0] };
    end 
    if(N2644) begin
      { mem[18111:18080] } <= { w_data_i[31:0] };
    end 
    if(N2643) begin
      { mem[18079:18048] } <= { w_data_i[31:0] };
    end 
    if(N2642) begin
      { mem[18047:18016] } <= { w_data_i[31:0] };
    end 
    if(N2641) begin
      { mem[18015:17984] } <= { w_data_i[31:0] };
    end 
    if(N2640) begin
      { mem[17983:17952] } <= { w_data_i[31:0] };
    end 
    if(N2639) begin
      { mem[17951:17920] } <= { w_data_i[31:0] };
    end 
    if(N2638) begin
      { mem[17919:17888] } <= { w_data_i[31:0] };
    end 
    if(N2637) begin
      { mem[17887:17856] } <= { w_data_i[31:0] };
    end 
    if(N2636) begin
      { mem[17855:17824] } <= { w_data_i[31:0] };
    end 
    if(N2635) begin
      { mem[17823:17792] } <= { w_data_i[31:0] };
    end 
    if(N2634) begin
      { mem[17791:17760] } <= { w_data_i[31:0] };
    end 
    if(N2633) begin
      { mem[17759:17728] } <= { w_data_i[31:0] };
    end 
    if(N2632) begin
      { mem[17727:17696] } <= { w_data_i[31:0] };
    end 
    if(N2631) begin
      { mem[17695:17664] } <= { w_data_i[31:0] };
    end 
    if(N2630) begin
      { mem[17663:17632] } <= { w_data_i[31:0] };
    end 
    if(N2629) begin
      { mem[17631:17600] } <= { w_data_i[31:0] };
    end 
    if(N2628) begin
      { mem[17599:17568] } <= { w_data_i[31:0] };
    end 
    if(N2627) begin
      { mem[17567:17536] } <= { w_data_i[31:0] };
    end 
    if(N2626) begin
      { mem[17535:17504] } <= { w_data_i[31:0] };
    end 
    if(N2625) begin
      { mem[17503:17472] } <= { w_data_i[31:0] };
    end 
    if(N2624) begin
      { mem[17471:17440] } <= { w_data_i[31:0] };
    end 
    if(N2623) begin
      { mem[17439:17408] } <= { w_data_i[31:0] };
    end 
    if(N2622) begin
      { mem[17407:17376] } <= { w_data_i[31:0] };
    end 
    if(N2621) begin
      { mem[17375:17344] } <= { w_data_i[31:0] };
    end 
    if(N2620) begin
      { mem[17343:17312] } <= { w_data_i[31:0] };
    end 
    if(N2619) begin
      { mem[17311:17280] } <= { w_data_i[31:0] };
    end 
    if(N2618) begin
      { mem[17279:17248] } <= { w_data_i[31:0] };
    end 
    if(N2617) begin
      { mem[17247:17216] } <= { w_data_i[31:0] };
    end 
    if(N2616) begin
      { mem[17215:17184] } <= { w_data_i[31:0] };
    end 
    if(N2615) begin
      { mem[17183:17152] } <= { w_data_i[31:0] };
    end 
    if(N2614) begin
      { mem[17151:17120] } <= { w_data_i[31:0] };
    end 
    if(N2613) begin
      { mem[17119:17088] } <= { w_data_i[31:0] };
    end 
    if(N2612) begin
      { mem[17087:17056] } <= { w_data_i[31:0] };
    end 
    if(N2611) begin
      { mem[17055:17024] } <= { w_data_i[31:0] };
    end 
    if(N2610) begin
      { mem[17023:16992] } <= { w_data_i[31:0] };
    end 
    if(N2609) begin
      { mem[16991:16960] } <= { w_data_i[31:0] };
    end 
    if(N2608) begin
      { mem[16959:16928] } <= { w_data_i[31:0] };
    end 
    if(N2607) begin
      { mem[16927:16896] } <= { w_data_i[31:0] };
    end 
    if(N2606) begin
      { mem[16895:16864] } <= { w_data_i[31:0] };
    end 
    if(N2605) begin
      { mem[16863:16832] } <= { w_data_i[31:0] };
    end 
    if(N2604) begin
      { mem[16831:16800] } <= { w_data_i[31:0] };
    end 
    if(N2603) begin
      { mem[16799:16768] } <= { w_data_i[31:0] };
    end 
    if(N2602) begin
      { mem[16767:16736] } <= { w_data_i[31:0] };
    end 
    if(N2601) begin
      { mem[16735:16704] } <= { w_data_i[31:0] };
    end 
    if(N2600) begin
      { mem[16703:16672] } <= { w_data_i[31:0] };
    end 
    if(N2599) begin
      { mem[16671:16640] } <= { w_data_i[31:0] };
    end 
    if(N2598) begin
      { mem[16639:16608] } <= { w_data_i[31:0] };
    end 
    if(N2597) begin
      { mem[16607:16576] } <= { w_data_i[31:0] };
    end 
    if(N2596) begin
      { mem[16575:16544] } <= { w_data_i[31:0] };
    end 
    if(N2595) begin
      { mem[16543:16512] } <= { w_data_i[31:0] };
    end 
    if(N2594) begin
      { mem[16511:16480] } <= { w_data_i[31:0] };
    end 
    if(N2593) begin
      { mem[16479:16448] } <= { w_data_i[31:0] };
    end 
    if(N2592) begin
      { mem[16447:16416] } <= { w_data_i[31:0] };
    end 
    if(N2591) begin
      { mem[16415:16384] } <= { w_data_i[31:0] };
    end 
    if(N2590) begin
      { mem[16383:16352] } <= { w_data_i[31:0] };
    end 
    if(N2589) begin
      { mem[16351:16320] } <= { w_data_i[31:0] };
    end 
    if(N2588) begin
      { mem[16319:16288] } <= { w_data_i[31:0] };
    end 
    if(N2587) begin
      { mem[16287:16256] } <= { w_data_i[31:0] };
    end 
    if(N2586) begin
      { mem[16255:16224] } <= { w_data_i[31:0] };
    end 
    if(N2585) begin
      { mem[16223:16192] } <= { w_data_i[31:0] };
    end 
    if(N2584) begin
      { mem[16191:16160] } <= { w_data_i[31:0] };
    end 
    if(N2583) begin
      { mem[16159:16128] } <= { w_data_i[31:0] };
    end 
    if(N2582) begin
      { mem[16127:16096] } <= { w_data_i[31:0] };
    end 
    if(N2581) begin
      { mem[16095:16064] } <= { w_data_i[31:0] };
    end 
    if(N2580) begin
      { mem[16063:16032] } <= { w_data_i[31:0] };
    end 
    if(N2579) begin
      { mem[16031:16000] } <= { w_data_i[31:0] };
    end 
    if(N2578) begin
      { mem[15999:15968] } <= { w_data_i[31:0] };
    end 
    if(N2577) begin
      { mem[15967:15936] } <= { w_data_i[31:0] };
    end 
    if(N2576) begin
      { mem[15935:15904] } <= { w_data_i[31:0] };
    end 
    if(N2575) begin
      { mem[15903:15872] } <= { w_data_i[31:0] };
    end 
    if(N2574) begin
      { mem[15871:15840] } <= { w_data_i[31:0] };
    end 
    if(N2573) begin
      { mem[15839:15808] } <= { w_data_i[31:0] };
    end 
    if(N2572) begin
      { mem[15807:15776] } <= { w_data_i[31:0] };
    end 
    if(N2571) begin
      { mem[15775:15744] } <= { w_data_i[31:0] };
    end 
    if(N2570) begin
      { mem[15743:15712] } <= { w_data_i[31:0] };
    end 
    if(N2569) begin
      { mem[15711:15680] } <= { w_data_i[31:0] };
    end 
    if(N2568) begin
      { mem[15679:15648] } <= { w_data_i[31:0] };
    end 
    if(N2567) begin
      { mem[15647:15616] } <= { w_data_i[31:0] };
    end 
    if(N2566) begin
      { mem[15615:15584] } <= { w_data_i[31:0] };
    end 
    if(N2565) begin
      { mem[15583:15552] } <= { w_data_i[31:0] };
    end 
    if(N2564) begin
      { mem[15551:15520] } <= { w_data_i[31:0] };
    end 
    if(N2563) begin
      { mem[15519:15488] } <= { w_data_i[31:0] };
    end 
    if(N2562) begin
      { mem[15487:15456] } <= { w_data_i[31:0] };
    end 
    if(N2561) begin
      { mem[15455:15424] } <= { w_data_i[31:0] };
    end 
    if(N2560) begin
      { mem[15423:15392] } <= { w_data_i[31:0] };
    end 
    if(N2559) begin
      { mem[15391:15360] } <= { w_data_i[31:0] };
    end 
    if(N2558) begin
      { mem[15359:15328] } <= { w_data_i[31:0] };
    end 
    if(N2557) begin
      { mem[15327:15296] } <= { w_data_i[31:0] };
    end 
    if(N2556) begin
      { mem[15295:15264] } <= { w_data_i[31:0] };
    end 
    if(N2555) begin
      { mem[15263:15232] } <= { w_data_i[31:0] };
    end 
    if(N2554) begin
      { mem[15231:15200] } <= { w_data_i[31:0] };
    end 
    if(N2553) begin
      { mem[15199:15168] } <= { w_data_i[31:0] };
    end 
    if(N2552) begin
      { mem[15167:15136] } <= { w_data_i[31:0] };
    end 
    if(N2551) begin
      { mem[15135:15104] } <= { w_data_i[31:0] };
    end 
    if(N2550) begin
      { mem[15103:15072] } <= { w_data_i[31:0] };
    end 
    if(N2549) begin
      { mem[15071:15040] } <= { w_data_i[31:0] };
    end 
    if(N2548) begin
      { mem[15039:15008] } <= { w_data_i[31:0] };
    end 
    if(N2547) begin
      { mem[15007:14976] } <= { w_data_i[31:0] };
    end 
    if(N2546) begin
      { mem[14975:14944] } <= { w_data_i[31:0] };
    end 
    if(N2545) begin
      { mem[14943:14912] } <= { w_data_i[31:0] };
    end 
    if(N2544) begin
      { mem[14911:14880] } <= { w_data_i[31:0] };
    end 
    if(N2543) begin
      { mem[14879:14848] } <= { w_data_i[31:0] };
    end 
    if(N2542) begin
      { mem[14847:14816] } <= { w_data_i[31:0] };
    end 
    if(N2541) begin
      { mem[14815:14784] } <= { w_data_i[31:0] };
    end 
    if(N2540) begin
      { mem[14783:14752] } <= { w_data_i[31:0] };
    end 
    if(N2539) begin
      { mem[14751:14720] } <= { w_data_i[31:0] };
    end 
    if(N2538) begin
      { mem[14719:14688] } <= { w_data_i[31:0] };
    end 
    if(N2537) begin
      { mem[14687:14656] } <= { w_data_i[31:0] };
    end 
    if(N2536) begin
      { mem[14655:14624] } <= { w_data_i[31:0] };
    end 
    if(N2535) begin
      { mem[14623:14592] } <= { w_data_i[31:0] };
    end 
    if(N2534) begin
      { mem[14591:14560] } <= { w_data_i[31:0] };
    end 
    if(N2533) begin
      { mem[14559:14528] } <= { w_data_i[31:0] };
    end 
    if(N2532) begin
      { mem[14527:14496] } <= { w_data_i[31:0] };
    end 
    if(N2531) begin
      { mem[14495:14464] } <= { w_data_i[31:0] };
    end 
    if(N2530) begin
      { mem[14463:14432] } <= { w_data_i[31:0] };
    end 
    if(N2529) begin
      { mem[14431:14400] } <= { w_data_i[31:0] };
    end 
    if(N2528) begin
      { mem[14399:14368] } <= { w_data_i[31:0] };
    end 
    if(N2527) begin
      { mem[14367:14336] } <= { w_data_i[31:0] };
    end 
    if(N2526) begin
      { mem[14335:14304] } <= { w_data_i[31:0] };
    end 
    if(N2525) begin
      { mem[14303:14272] } <= { w_data_i[31:0] };
    end 
    if(N2524) begin
      { mem[14271:14240] } <= { w_data_i[31:0] };
    end 
    if(N2523) begin
      { mem[14239:14208] } <= { w_data_i[31:0] };
    end 
    if(N2522) begin
      { mem[14207:14176] } <= { w_data_i[31:0] };
    end 
    if(N2521) begin
      { mem[14175:14144] } <= { w_data_i[31:0] };
    end 
    if(N2520) begin
      { mem[14143:14112] } <= { w_data_i[31:0] };
    end 
    if(N2519) begin
      { mem[14111:14080] } <= { w_data_i[31:0] };
    end 
    if(N2518) begin
      { mem[14079:14048] } <= { w_data_i[31:0] };
    end 
    if(N2517) begin
      { mem[14047:14016] } <= { w_data_i[31:0] };
    end 
    if(N2516) begin
      { mem[14015:13984] } <= { w_data_i[31:0] };
    end 
    if(N2515) begin
      { mem[13983:13952] } <= { w_data_i[31:0] };
    end 
    if(N2514) begin
      { mem[13951:13920] } <= { w_data_i[31:0] };
    end 
    if(N2513) begin
      { mem[13919:13888] } <= { w_data_i[31:0] };
    end 
    if(N2512) begin
      { mem[13887:13856] } <= { w_data_i[31:0] };
    end 
    if(N2511) begin
      { mem[13855:13824] } <= { w_data_i[31:0] };
    end 
    if(N2510) begin
      { mem[13823:13792] } <= { w_data_i[31:0] };
    end 
    if(N2509) begin
      { mem[13791:13760] } <= { w_data_i[31:0] };
    end 
    if(N2508) begin
      { mem[13759:13728] } <= { w_data_i[31:0] };
    end 
    if(N2507) begin
      { mem[13727:13696] } <= { w_data_i[31:0] };
    end 
    if(N2506) begin
      { mem[13695:13664] } <= { w_data_i[31:0] };
    end 
    if(N2505) begin
      { mem[13663:13632] } <= { w_data_i[31:0] };
    end 
    if(N2504) begin
      { mem[13631:13600] } <= { w_data_i[31:0] };
    end 
    if(N2503) begin
      { mem[13599:13568] } <= { w_data_i[31:0] };
    end 
    if(N2502) begin
      { mem[13567:13536] } <= { w_data_i[31:0] };
    end 
    if(N2501) begin
      { mem[13535:13504] } <= { w_data_i[31:0] };
    end 
    if(N2500) begin
      { mem[13503:13472] } <= { w_data_i[31:0] };
    end 
    if(N2499) begin
      { mem[13471:13440] } <= { w_data_i[31:0] };
    end 
    if(N2498) begin
      { mem[13439:13408] } <= { w_data_i[31:0] };
    end 
    if(N2497) begin
      { mem[13407:13376] } <= { w_data_i[31:0] };
    end 
    if(N2496) begin
      { mem[13375:13344] } <= { w_data_i[31:0] };
    end 
    if(N2495) begin
      { mem[13343:13312] } <= { w_data_i[31:0] };
    end 
    if(N2494) begin
      { mem[13311:13280] } <= { w_data_i[31:0] };
    end 
    if(N2493) begin
      { mem[13279:13248] } <= { w_data_i[31:0] };
    end 
    if(N2492) begin
      { mem[13247:13216] } <= { w_data_i[31:0] };
    end 
    if(N2491) begin
      { mem[13215:13184] } <= { w_data_i[31:0] };
    end 
    if(N2490) begin
      { mem[13183:13152] } <= { w_data_i[31:0] };
    end 
    if(N2489) begin
      { mem[13151:13120] } <= { w_data_i[31:0] };
    end 
    if(N2488) begin
      { mem[13119:13088] } <= { w_data_i[31:0] };
    end 
    if(N2487) begin
      { mem[13087:13056] } <= { w_data_i[31:0] };
    end 
    if(N2486) begin
      { mem[13055:13024] } <= { w_data_i[31:0] };
    end 
    if(N2485) begin
      { mem[13023:12992] } <= { w_data_i[31:0] };
    end 
    if(N2484) begin
      { mem[12991:12960] } <= { w_data_i[31:0] };
    end 
    if(N2483) begin
      { mem[12959:12928] } <= { w_data_i[31:0] };
    end 
    if(N2482) begin
      { mem[12927:12896] } <= { w_data_i[31:0] };
    end 
    if(N2481) begin
      { mem[12895:12864] } <= { w_data_i[31:0] };
    end 
    if(N2480) begin
      { mem[12863:12832] } <= { w_data_i[31:0] };
    end 
    if(N2479) begin
      { mem[12831:12800] } <= { w_data_i[31:0] };
    end 
    if(N2478) begin
      { mem[12799:12768] } <= { w_data_i[31:0] };
    end 
    if(N2477) begin
      { mem[12767:12736] } <= { w_data_i[31:0] };
    end 
    if(N2476) begin
      { mem[12735:12704] } <= { w_data_i[31:0] };
    end 
    if(N2475) begin
      { mem[12703:12672] } <= { w_data_i[31:0] };
    end 
    if(N2474) begin
      { mem[12671:12640] } <= { w_data_i[31:0] };
    end 
    if(N2473) begin
      { mem[12639:12608] } <= { w_data_i[31:0] };
    end 
    if(N2472) begin
      { mem[12607:12576] } <= { w_data_i[31:0] };
    end 
    if(N2471) begin
      { mem[12575:12544] } <= { w_data_i[31:0] };
    end 
    if(N2470) begin
      { mem[12543:12512] } <= { w_data_i[31:0] };
    end 
    if(N2469) begin
      { mem[12511:12480] } <= { w_data_i[31:0] };
    end 
    if(N2468) begin
      { mem[12479:12448] } <= { w_data_i[31:0] };
    end 
    if(N2467) begin
      { mem[12447:12416] } <= { w_data_i[31:0] };
    end 
    if(N2466) begin
      { mem[12415:12384] } <= { w_data_i[31:0] };
    end 
    if(N2465) begin
      { mem[12383:12352] } <= { w_data_i[31:0] };
    end 
    if(N2464) begin
      { mem[12351:12320] } <= { w_data_i[31:0] };
    end 
    if(N2463) begin
      { mem[12319:12288] } <= { w_data_i[31:0] };
    end 
    if(N2462) begin
      { mem[12287:12256] } <= { w_data_i[31:0] };
    end 
    if(N2461) begin
      { mem[12255:12224] } <= { w_data_i[31:0] };
    end 
    if(N2460) begin
      { mem[12223:12192] } <= { w_data_i[31:0] };
    end 
    if(N2459) begin
      { mem[12191:12160] } <= { w_data_i[31:0] };
    end 
    if(N2458) begin
      { mem[12159:12128] } <= { w_data_i[31:0] };
    end 
    if(N2457) begin
      { mem[12127:12096] } <= { w_data_i[31:0] };
    end 
    if(N2456) begin
      { mem[12095:12064] } <= { w_data_i[31:0] };
    end 
    if(N2455) begin
      { mem[12063:12032] } <= { w_data_i[31:0] };
    end 
    if(N2454) begin
      { mem[12031:12000] } <= { w_data_i[31:0] };
    end 
    if(N2453) begin
      { mem[11999:11968] } <= { w_data_i[31:0] };
    end 
    if(N2452) begin
      { mem[11967:11936] } <= { w_data_i[31:0] };
    end 
    if(N2451) begin
      { mem[11935:11904] } <= { w_data_i[31:0] };
    end 
    if(N2450) begin
      { mem[11903:11872] } <= { w_data_i[31:0] };
    end 
    if(N2449) begin
      { mem[11871:11840] } <= { w_data_i[31:0] };
    end 
    if(N2448) begin
      { mem[11839:11808] } <= { w_data_i[31:0] };
    end 
    if(N2447) begin
      { mem[11807:11776] } <= { w_data_i[31:0] };
    end 
    if(N2446) begin
      { mem[11775:11744] } <= { w_data_i[31:0] };
    end 
    if(N2445) begin
      { mem[11743:11712] } <= { w_data_i[31:0] };
    end 
    if(N2444) begin
      { mem[11711:11680] } <= { w_data_i[31:0] };
    end 
    if(N2443) begin
      { mem[11679:11648] } <= { w_data_i[31:0] };
    end 
    if(N2442) begin
      { mem[11647:11616] } <= { w_data_i[31:0] };
    end 
    if(N2441) begin
      { mem[11615:11584] } <= { w_data_i[31:0] };
    end 
    if(N2440) begin
      { mem[11583:11552] } <= { w_data_i[31:0] };
    end 
    if(N2439) begin
      { mem[11551:11520] } <= { w_data_i[31:0] };
    end 
    if(N2438) begin
      { mem[11519:11488] } <= { w_data_i[31:0] };
    end 
    if(N2437) begin
      { mem[11487:11456] } <= { w_data_i[31:0] };
    end 
    if(N2436) begin
      { mem[11455:11424] } <= { w_data_i[31:0] };
    end 
    if(N2435) begin
      { mem[11423:11392] } <= { w_data_i[31:0] };
    end 
    if(N2434) begin
      { mem[11391:11360] } <= { w_data_i[31:0] };
    end 
    if(N2433) begin
      { mem[11359:11328] } <= { w_data_i[31:0] };
    end 
    if(N2432) begin
      { mem[11327:11296] } <= { w_data_i[31:0] };
    end 
    if(N2431) begin
      { mem[11295:11264] } <= { w_data_i[31:0] };
    end 
    if(N2430) begin
      { mem[11263:11232] } <= { w_data_i[31:0] };
    end 
    if(N2429) begin
      { mem[11231:11200] } <= { w_data_i[31:0] };
    end 
    if(N2428) begin
      { mem[11199:11168] } <= { w_data_i[31:0] };
    end 
    if(N2427) begin
      { mem[11167:11136] } <= { w_data_i[31:0] };
    end 
    if(N2426) begin
      { mem[11135:11104] } <= { w_data_i[31:0] };
    end 
    if(N2425) begin
      { mem[11103:11072] } <= { w_data_i[31:0] };
    end 
    if(N2424) begin
      { mem[11071:11040] } <= { w_data_i[31:0] };
    end 
    if(N2423) begin
      { mem[11039:11008] } <= { w_data_i[31:0] };
    end 
    if(N2422) begin
      { mem[11007:10976] } <= { w_data_i[31:0] };
    end 
    if(N2421) begin
      { mem[10975:10944] } <= { w_data_i[31:0] };
    end 
    if(N2420) begin
      { mem[10943:10912] } <= { w_data_i[31:0] };
    end 
    if(N2419) begin
      { mem[10911:10880] } <= { w_data_i[31:0] };
    end 
    if(N2418) begin
      { mem[10879:10848] } <= { w_data_i[31:0] };
    end 
    if(N2417) begin
      { mem[10847:10816] } <= { w_data_i[31:0] };
    end 
    if(N2416) begin
      { mem[10815:10784] } <= { w_data_i[31:0] };
    end 
    if(N2415) begin
      { mem[10783:10752] } <= { w_data_i[31:0] };
    end 
    if(N2414) begin
      { mem[10751:10720] } <= { w_data_i[31:0] };
    end 
    if(N2413) begin
      { mem[10719:10688] } <= { w_data_i[31:0] };
    end 
    if(N2412) begin
      { mem[10687:10656] } <= { w_data_i[31:0] };
    end 
    if(N2411) begin
      { mem[10655:10624] } <= { w_data_i[31:0] };
    end 
    if(N2410) begin
      { mem[10623:10592] } <= { w_data_i[31:0] };
    end 
    if(N2409) begin
      { mem[10591:10560] } <= { w_data_i[31:0] };
    end 
    if(N2408) begin
      { mem[10559:10528] } <= { w_data_i[31:0] };
    end 
    if(N2407) begin
      { mem[10527:10496] } <= { w_data_i[31:0] };
    end 
    if(N2406) begin
      { mem[10495:10464] } <= { w_data_i[31:0] };
    end 
    if(N2405) begin
      { mem[10463:10432] } <= { w_data_i[31:0] };
    end 
    if(N2404) begin
      { mem[10431:10400] } <= { w_data_i[31:0] };
    end 
    if(N2403) begin
      { mem[10399:10368] } <= { w_data_i[31:0] };
    end 
    if(N2402) begin
      { mem[10367:10336] } <= { w_data_i[31:0] };
    end 
    if(N2401) begin
      { mem[10335:10304] } <= { w_data_i[31:0] };
    end 
    if(N2400) begin
      { mem[10303:10272] } <= { w_data_i[31:0] };
    end 
    if(N2399) begin
      { mem[10271:10240] } <= { w_data_i[31:0] };
    end 
    if(N2398) begin
      { mem[10239:10208] } <= { w_data_i[31:0] };
    end 
    if(N2397) begin
      { mem[10207:10176] } <= { w_data_i[31:0] };
    end 
    if(N2396) begin
      { mem[10175:10144] } <= { w_data_i[31:0] };
    end 
    if(N2395) begin
      { mem[10143:10112] } <= { w_data_i[31:0] };
    end 
    if(N2394) begin
      { mem[10111:10080] } <= { w_data_i[31:0] };
    end 
    if(N2393) begin
      { mem[10079:10048] } <= { w_data_i[31:0] };
    end 
    if(N2392) begin
      { mem[10047:10016] } <= { w_data_i[31:0] };
    end 
    if(N2391) begin
      { mem[10015:9984] } <= { w_data_i[31:0] };
    end 
    if(N2390) begin
      { mem[9983:9952] } <= { w_data_i[31:0] };
    end 
    if(N2389) begin
      { mem[9951:9920] } <= { w_data_i[31:0] };
    end 
    if(N2388) begin
      { mem[9919:9888] } <= { w_data_i[31:0] };
    end 
    if(N2387) begin
      { mem[9887:9856] } <= { w_data_i[31:0] };
    end 
    if(N2386) begin
      { mem[9855:9824] } <= { w_data_i[31:0] };
    end 
    if(N2385) begin
      { mem[9823:9792] } <= { w_data_i[31:0] };
    end 
    if(N2384) begin
      { mem[9791:9760] } <= { w_data_i[31:0] };
    end 
    if(N2383) begin
      { mem[9759:9728] } <= { w_data_i[31:0] };
    end 
    if(N2382) begin
      { mem[9727:9696] } <= { w_data_i[31:0] };
    end 
    if(N2381) begin
      { mem[9695:9664] } <= { w_data_i[31:0] };
    end 
    if(N2380) begin
      { mem[9663:9632] } <= { w_data_i[31:0] };
    end 
    if(N2379) begin
      { mem[9631:9600] } <= { w_data_i[31:0] };
    end 
    if(N2378) begin
      { mem[9599:9568] } <= { w_data_i[31:0] };
    end 
    if(N2377) begin
      { mem[9567:9536] } <= { w_data_i[31:0] };
    end 
    if(N2376) begin
      { mem[9535:9504] } <= { w_data_i[31:0] };
    end 
    if(N2375) begin
      { mem[9503:9472] } <= { w_data_i[31:0] };
    end 
    if(N2374) begin
      { mem[9471:9440] } <= { w_data_i[31:0] };
    end 
    if(N2373) begin
      { mem[9439:9408] } <= { w_data_i[31:0] };
    end 
    if(N2372) begin
      { mem[9407:9376] } <= { w_data_i[31:0] };
    end 
    if(N2371) begin
      { mem[9375:9344] } <= { w_data_i[31:0] };
    end 
    if(N2370) begin
      { mem[9343:9312] } <= { w_data_i[31:0] };
    end 
    if(N2369) begin
      { mem[9311:9280] } <= { w_data_i[31:0] };
    end 
    if(N2368) begin
      { mem[9279:9248] } <= { w_data_i[31:0] };
    end 
    if(N2367) begin
      { mem[9247:9216] } <= { w_data_i[31:0] };
    end 
    if(N2366) begin
      { mem[9215:9184] } <= { w_data_i[31:0] };
    end 
    if(N2365) begin
      { mem[9183:9152] } <= { w_data_i[31:0] };
    end 
    if(N2364) begin
      { mem[9151:9120] } <= { w_data_i[31:0] };
    end 
    if(N2363) begin
      { mem[9119:9088] } <= { w_data_i[31:0] };
    end 
    if(N2362) begin
      { mem[9087:9056] } <= { w_data_i[31:0] };
    end 
    if(N2361) begin
      { mem[9055:9024] } <= { w_data_i[31:0] };
    end 
    if(N2360) begin
      { mem[9023:8992] } <= { w_data_i[31:0] };
    end 
    if(N2359) begin
      { mem[8991:8960] } <= { w_data_i[31:0] };
    end 
    if(N2358) begin
      { mem[8959:8928] } <= { w_data_i[31:0] };
    end 
    if(N2357) begin
      { mem[8927:8896] } <= { w_data_i[31:0] };
    end 
    if(N2356) begin
      { mem[8895:8864] } <= { w_data_i[31:0] };
    end 
    if(N2355) begin
      { mem[8863:8832] } <= { w_data_i[31:0] };
    end 
    if(N2354) begin
      { mem[8831:8800] } <= { w_data_i[31:0] };
    end 
    if(N2353) begin
      { mem[8799:8768] } <= { w_data_i[31:0] };
    end 
    if(N2352) begin
      { mem[8767:8736] } <= { w_data_i[31:0] };
    end 
    if(N2351) begin
      { mem[8735:8704] } <= { w_data_i[31:0] };
    end 
    if(N2350) begin
      { mem[8703:8672] } <= { w_data_i[31:0] };
    end 
    if(N2349) begin
      { mem[8671:8640] } <= { w_data_i[31:0] };
    end 
    if(N2348) begin
      { mem[8639:8608] } <= { w_data_i[31:0] };
    end 
    if(N2347) begin
      { mem[8607:8576] } <= { w_data_i[31:0] };
    end 
    if(N2346) begin
      { mem[8575:8544] } <= { w_data_i[31:0] };
    end 
    if(N2345) begin
      { mem[8543:8512] } <= { w_data_i[31:0] };
    end 
    if(N2344) begin
      { mem[8511:8480] } <= { w_data_i[31:0] };
    end 
    if(N2343) begin
      { mem[8479:8448] } <= { w_data_i[31:0] };
    end 
    if(N2342) begin
      { mem[8447:8416] } <= { w_data_i[31:0] };
    end 
    if(N2341) begin
      { mem[8415:8384] } <= { w_data_i[31:0] };
    end 
    if(N2340) begin
      { mem[8383:8352] } <= { w_data_i[31:0] };
    end 
    if(N2339) begin
      { mem[8351:8320] } <= { w_data_i[31:0] };
    end 
    if(N2338) begin
      { mem[8319:8288] } <= { w_data_i[31:0] };
    end 
    if(N2337) begin
      { mem[8287:8256] } <= { w_data_i[31:0] };
    end 
    if(N2336) begin
      { mem[8255:8224] } <= { w_data_i[31:0] };
    end 
    if(N2335) begin
      { mem[8223:8192] } <= { w_data_i[31:0] };
    end 
    if(N2334) begin
      { mem[8191:8160] } <= { w_data_i[31:0] };
    end 
    if(N2333) begin
      { mem[8159:8128] } <= { w_data_i[31:0] };
    end 
    if(N2332) begin
      { mem[8127:8096] } <= { w_data_i[31:0] };
    end 
    if(N2331) begin
      { mem[8095:8064] } <= { w_data_i[31:0] };
    end 
    if(N2330) begin
      { mem[8063:8032] } <= { w_data_i[31:0] };
    end 
    if(N2329) begin
      { mem[8031:8000] } <= { w_data_i[31:0] };
    end 
    if(N2328) begin
      { mem[7999:7968] } <= { w_data_i[31:0] };
    end 
    if(N2327) begin
      { mem[7967:7936] } <= { w_data_i[31:0] };
    end 
    if(N2326) begin
      { mem[7935:7904] } <= { w_data_i[31:0] };
    end 
    if(N2325) begin
      { mem[7903:7872] } <= { w_data_i[31:0] };
    end 
    if(N2324) begin
      { mem[7871:7840] } <= { w_data_i[31:0] };
    end 
    if(N2323) begin
      { mem[7839:7808] } <= { w_data_i[31:0] };
    end 
    if(N2322) begin
      { mem[7807:7776] } <= { w_data_i[31:0] };
    end 
    if(N2321) begin
      { mem[7775:7744] } <= { w_data_i[31:0] };
    end 
    if(N2320) begin
      { mem[7743:7712] } <= { w_data_i[31:0] };
    end 
    if(N2319) begin
      { mem[7711:7680] } <= { w_data_i[31:0] };
    end 
    if(N2318) begin
      { mem[7679:7648] } <= { w_data_i[31:0] };
    end 
    if(N2317) begin
      { mem[7647:7616] } <= { w_data_i[31:0] };
    end 
    if(N2316) begin
      { mem[7615:7584] } <= { w_data_i[31:0] };
    end 
    if(N2315) begin
      { mem[7583:7552] } <= { w_data_i[31:0] };
    end 
    if(N2314) begin
      { mem[7551:7520] } <= { w_data_i[31:0] };
    end 
    if(N2313) begin
      { mem[7519:7488] } <= { w_data_i[31:0] };
    end 
    if(N2312) begin
      { mem[7487:7456] } <= { w_data_i[31:0] };
    end 
    if(N2311) begin
      { mem[7455:7424] } <= { w_data_i[31:0] };
    end 
    if(N2310) begin
      { mem[7423:7392] } <= { w_data_i[31:0] };
    end 
    if(N2309) begin
      { mem[7391:7360] } <= { w_data_i[31:0] };
    end 
    if(N2308) begin
      { mem[7359:7328] } <= { w_data_i[31:0] };
    end 
    if(N2307) begin
      { mem[7327:7296] } <= { w_data_i[31:0] };
    end 
    if(N2306) begin
      { mem[7295:7264] } <= { w_data_i[31:0] };
    end 
    if(N2305) begin
      { mem[7263:7232] } <= { w_data_i[31:0] };
    end 
    if(N2304) begin
      { mem[7231:7200] } <= { w_data_i[31:0] };
    end 
    if(N2303) begin
      { mem[7199:7168] } <= { w_data_i[31:0] };
    end 
    if(N2302) begin
      { mem[7167:7136] } <= { w_data_i[31:0] };
    end 
    if(N2301) begin
      { mem[7135:7104] } <= { w_data_i[31:0] };
    end 
    if(N2300) begin
      { mem[7103:7072] } <= { w_data_i[31:0] };
    end 
    if(N2299) begin
      { mem[7071:7040] } <= { w_data_i[31:0] };
    end 
    if(N2298) begin
      { mem[7039:7008] } <= { w_data_i[31:0] };
    end 
    if(N2297) begin
      { mem[7007:6976] } <= { w_data_i[31:0] };
    end 
    if(N2296) begin
      { mem[6975:6944] } <= { w_data_i[31:0] };
    end 
    if(N2295) begin
      { mem[6943:6912] } <= { w_data_i[31:0] };
    end 
    if(N2294) begin
      { mem[6911:6880] } <= { w_data_i[31:0] };
    end 
    if(N2293) begin
      { mem[6879:6848] } <= { w_data_i[31:0] };
    end 
    if(N2292) begin
      { mem[6847:6816] } <= { w_data_i[31:0] };
    end 
    if(N2291) begin
      { mem[6815:6784] } <= { w_data_i[31:0] };
    end 
    if(N2290) begin
      { mem[6783:6752] } <= { w_data_i[31:0] };
    end 
    if(N2289) begin
      { mem[6751:6720] } <= { w_data_i[31:0] };
    end 
    if(N2288) begin
      { mem[6719:6688] } <= { w_data_i[31:0] };
    end 
    if(N2287) begin
      { mem[6687:6656] } <= { w_data_i[31:0] };
    end 
    if(N2286) begin
      { mem[6655:6624] } <= { w_data_i[31:0] };
    end 
    if(N2285) begin
      { mem[6623:6592] } <= { w_data_i[31:0] };
    end 
    if(N2284) begin
      { mem[6591:6560] } <= { w_data_i[31:0] };
    end 
    if(N2283) begin
      { mem[6559:6528] } <= { w_data_i[31:0] };
    end 
    if(N2282) begin
      { mem[6527:6496] } <= { w_data_i[31:0] };
    end 
    if(N2281) begin
      { mem[6495:6464] } <= { w_data_i[31:0] };
    end 
    if(N2280) begin
      { mem[6463:6432] } <= { w_data_i[31:0] };
    end 
    if(N2279) begin
      { mem[6431:6400] } <= { w_data_i[31:0] };
    end 
    if(N2278) begin
      { mem[6399:6368] } <= { w_data_i[31:0] };
    end 
    if(N2277) begin
      { mem[6367:6336] } <= { w_data_i[31:0] };
    end 
    if(N2276) begin
      { mem[6335:6304] } <= { w_data_i[31:0] };
    end 
    if(N2275) begin
      { mem[6303:6272] } <= { w_data_i[31:0] };
    end 
    if(N2274) begin
      { mem[6271:6240] } <= { w_data_i[31:0] };
    end 
    if(N2273) begin
      { mem[6239:6208] } <= { w_data_i[31:0] };
    end 
    if(N2272) begin
      { mem[6207:6176] } <= { w_data_i[31:0] };
    end 
    if(N2271) begin
      { mem[6175:6144] } <= { w_data_i[31:0] };
    end 
    if(N2270) begin
      { mem[6143:6112] } <= { w_data_i[31:0] };
    end 
    if(N2269) begin
      { mem[6111:6080] } <= { w_data_i[31:0] };
    end 
    if(N2268) begin
      { mem[6079:6048] } <= { w_data_i[31:0] };
    end 
    if(N2267) begin
      { mem[6047:6016] } <= { w_data_i[31:0] };
    end 
    if(N2266) begin
      { mem[6015:5984] } <= { w_data_i[31:0] };
    end 
    if(N2265) begin
      { mem[5983:5952] } <= { w_data_i[31:0] };
    end 
    if(N2264) begin
      { mem[5951:5920] } <= { w_data_i[31:0] };
    end 
    if(N2263) begin
      { mem[5919:5888] } <= { w_data_i[31:0] };
    end 
    if(N2262) begin
      { mem[5887:5856] } <= { w_data_i[31:0] };
    end 
    if(N2261) begin
      { mem[5855:5824] } <= { w_data_i[31:0] };
    end 
    if(N2260) begin
      { mem[5823:5792] } <= { w_data_i[31:0] };
    end 
    if(N2259) begin
      { mem[5791:5760] } <= { w_data_i[31:0] };
    end 
    if(N2258) begin
      { mem[5759:5728] } <= { w_data_i[31:0] };
    end 
    if(N2257) begin
      { mem[5727:5696] } <= { w_data_i[31:0] };
    end 
    if(N2256) begin
      { mem[5695:5664] } <= { w_data_i[31:0] };
    end 
    if(N2255) begin
      { mem[5663:5632] } <= { w_data_i[31:0] };
    end 
    if(N2254) begin
      { mem[5631:5600] } <= { w_data_i[31:0] };
    end 
    if(N2253) begin
      { mem[5599:5568] } <= { w_data_i[31:0] };
    end 
    if(N2252) begin
      { mem[5567:5536] } <= { w_data_i[31:0] };
    end 
    if(N2251) begin
      { mem[5535:5504] } <= { w_data_i[31:0] };
    end 
    if(N2250) begin
      { mem[5503:5472] } <= { w_data_i[31:0] };
    end 
    if(N2249) begin
      { mem[5471:5440] } <= { w_data_i[31:0] };
    end 
    if(N2248) begin
      { mem[5439:5408] } <= { w_data_i[31:0] };
    end 
    if(N2247) begin
      { mem[5407:5376] } <= { w_data_i[31:0] };
    end 
    if(N2246) begin
      { mem[5375:5344] } <= { w_data_i[31:0] };
    end 
    if(N2245) begin
      { mem[5343:5312] } <= { w_data_i[31:0] };
    end 
    if(N2244) begin
      { mem[5311:5280] } <= { w_data_i[31:0] };
    end 
    if(N2243) begin
      { mem[5279:5248] } <= { w_data_i[31:0] };
    end 
    if(N2242) begin
      { mem[5247:5216] } <= { w_data_i[31:0] };
    end 
    if(N2241) begin
      { mem[5215:5184] } <= { w_data_i[31:0] };
    end 
    if(N2240) begin
      { mem[5183:5152] } <= { w_data_i[31:0] };
    end 
    if(N2239) begin
      { mem[5151:5120] } <= { w_data_i[31:0] };
    end 
    if(N2238) begin
      { mem[5119:5088] } <= { w_data_i[31:0] };
    end 
    if(N2237) begin
      { mem[5087:5056] } <= { w_data_i[31:0] };
    end 
    if(N2236) begin
      { mem[5055:5024] } <= { w_data_i[31:0] };
    end 
    if(N2235) begin
      { mem[5023:4992] } <= { w_data_i[31:0] };
    end 
    if(N2234) begin
      { mem[4991:4960] } <= { w_data_i[31:0] };
    end 
    if(N2233) begin
      { mem[4959:4928] } <= { w_data_i[31:0] };
    end 
    if(N2232) begin
      { mem[4927:4896] } <= { w_data_i[31:0] };
    end 
    if(N2231) begin
      { mem[4895:4864] } <= { w_data_i[31:0] };
    end 
    if(N2230) begin
      { mem[4863:4832] } <= { w_data_i[31:0] };
    end 
    if(N2229) begin
      { mem[4831:4800] } <= { w_data_i[31:0] };
    end 
    if(N2228) begin
      { mem[4799:4768] } <= { w_data_i[31:0] };
    end 
    if(N2227) begin
      { mem[4767:4736] } <= { w_data_i[31:0] };
    end 
    if(N2226) begin
      { mem[4735:4704] } <= { w_data_i[31:0] };
    end 
    if(N2225) begin
      { mem[4703:4672] } <= { w_data_i[31:0] };
    end 
    if(N2224) begin
      { mem[4671:4640] } <= { w_data_i[31:0] };
    end 
    if(N2223) begin
      { mem[4639:4608] } <= { w_data_i[31:0] };
    end 
    if(N2222) begin
      { mem[4607:4576] } <= { w_data_i[31:0] };
    end 
    if(N2221) begin
      { mem[4575:4544] } <= { w_data_i[31:0] };
    end 
    if(N2220) begin
      { mem[4543:4512] } <= { w_data_i[31:0] };
    end 
    if(N2219) begin
      { mem[4511:4480] } <= { w_data_i[31:0] };
    end 
    if(N2218) begin
      { mem[4479:4448] } <= { w_data_i[31:0] };
    end 
    if(N2217) begin
      { mem[4447:4416] } <= { w_data_i[31:0] };
    end 
    if(N2216) begin
      { mem[4415:4384] } <= { w_data_i[31:0] };
    end 
    if(N2215) begin
      { mem[4383:4352] } <= { w_data_i[31:0] };
    end 
    if(N2214) begin
      { mem[4351:4320] } <= { w_data_i[31:0] };
    end 
    if(N2213) begin
      { mem[4319:4288] } <= { w_data_i[31:0] };
    end 
    if(N2212) begin
      { mem[4287:4256] } <= { w_data_i[31:0] };
    end 
    if(N2211) begin
      { mem[4255:4224] } <= { w_data_i[31:0] };
    end 
    if(N2210) begin
      { mem[4223:4192] } <= { w_data_i[31:0] };
    end 
    if(N2209) begin
      { mem[4191:4160] } <= { w_data_i[31:0] };
    end 
    if(N2208) begin
      { mem[4159:4128] } <= { w_data_i[31:0] };
    end 
    if(N2207) begin
      { mem[4127:4096] } <= { w_data_i[31:0] };
    end 
    if(N2206) begin
      { mem[4095:4064] } <= { w_data_i[31:0] };
    end 
    if(N2205) begin
      { mem[4063:4032] } <= { w_data_i[31:0] };
    end 
    if(N2204) begin
      { mem[4031:4000] } <= { w_data_i[31:0] };
    end 
    if(N2203) begin
      { mem[3999:3968] } <= { w_data_i[31:0] };
    end 
    if(N2202) begin
      { mem[3967:3936] } <= { w_data_i[31:0] };
    end 
    if(N2201) begin
      { mem[3935:3904] } <= { w_data_i[31:0] };
    end 
    if(N2200) begin
      { mem[3903:3872] } <= { w_data_i[31:0] };
    end 
    if(N2199) begin
      { mem[3871:3840] } <= { w_data_i[31:0] };
    end 
    if(N2198) begin
      { mem[3839:3808] } <= { w_data_i[31:0] };
    end 
    if(N2197) begin
      { mem[3807:3776] } <= { w_data_i[31:0] };
    end 
    if(N2196) begin
      { mem[3775:3744] } <= { w_data_i[31:0] };
    end 
    if(N2195) begin
      { mem[3743:3712] } <= { w_data_i[31:0] };
    end 
    if(N2194) begin
      { mem[3711:3680] } <= { w_data_i[31:0] };
    end 
    if(N2193) begin
      { mem[3679:3648] } <= { w_data_i[31:0] };
    end 
    if(N2192) begin
      { mem[3647:3616] } <= { w_data_i[31:0] };
    end 
    if(N2191) begin
      { mem[3615:3584] } <= { w_data_i[31:0] };
    end 
    if(N2190) begin
      { mem[3583:3552] } <= { w_data_i[31:0] };
    end 
    if(N2189) begin
      { mem[3551:3520] } <= { w_data_i[31:0] };
    end 
    if(N2188) begin
      { mem[3519:3488] } <= { w_data_i[31:0] };
    end 
    if(N2187) begin
      { mem[3487:3456] } <= { w_data_i[31:0] };
    end 
    if(N2186) begin
      { mem[3455:3424] } <= { w_data_i[31:0] };
    end 
    if(N2185) begin
      { mem[3423:3392] } <= { w_data_i[31:0] };
    end 
    if(N2184) begin
      { mem[3391:3360] } <= { w_data_i[31:0] };
    end 
    if(N2183) begin
      { mem[3359:3328] } <= { w_data_i[31:0] };
    end 
    if(N2182) begin
      { mem[3327:3296] } <= { w_data_i[31:0] };
    end 
    if(N2181) begin
      { mem[3295:3264] } <= { w_data_i[31:0] };
    end 
    if(N2180) begin
      { mem[3263:3232] } <= { w_data_i[31:0] };
    end 
    if(N2179) begin
      { mem[3231:3200] } <= { w_data_i[31:0] };
    end 
    if(N2178) begin
      { mem[3199:3168] } <= { w_data_i[31:0] };
    end 
    if(N2177) begin
      { mem[3167:3136] } <= { w_data_i[31:0] };
    end 
    if(N2176) begin
      { mem[3135:3104] } <= { w_data_i[31:0] };
    end 
    if(N2175) begin
      { mem[3103:3072] } <= { w_data_i[31:0] };
    end 
    if(N2174) begin
      { mem[3071:3040] } <= { w_data_i[31:0] };
    end 
    if(N2173) begin
      { mem[3039:3008] } <= { w_data_i[31:0] };
    end 
    if(N2172) begin
      { mem[3007:2976] } <= { w_data_i[31:0] };
    end 
    if(N2171) begin
      { mem[2975:2944] } <= { w_data_i[31:0] };
    end 
    if(N2170) begin
      { mem[2943:2912] } <= { w_data_i[31:0] };
    end 
    if(N2169) begin
      { mem[2911:2880] } <= { w_data_i[31:0] };
    end 
    if(N2168) begin
      { mem[2879:2848] } <= { w_data_i[31:0] };
    end 
    if(N2167) begin
      { mem[2847:2816] } <= { w_data_i[31:0] };
    end 
    if(N2166) begin
      { mem[2815:2784] } <= { w_data_i[31:0] };
    end 
    if(N2165) begin
      { mem[2783:2752] } <= { w_data_i[31:0] };
    end 
    if(N2164) begin
      { mem[2751:2720] } <= { w_data_i[31:0] };
    end 
    if(N2163) begin
      { mem[2719:2688] } <= { w_data_i[31:0] };
    end 
    if(N2162) begin
      { mem[2687:2656] } <= { w_data_i[31:0] };
    end 
    if(N2161) begin
      { mem[2655:2624] } <= { w_data_i[31:0] };
    end 
    if(N2160) begin
      { mem[2623:2592] } <= { w_data_i[31:0] };
    end 
    if(N2159) begin
      { mem[2591:2560] } <= { w_data_i[31:0] };
    end 
    if(N2158) begin
      { mem[2559:2528] } <= { w_data_i[31:0] };
    end 
    if(N2157) begin
      { mem[2527:2496] } <= { w_data_i[31:0] };
    end 
    if(N2156) begin
      { mem[2495:2464] } <= { w_data_i[31:0] };
    end 
    if(N2155) begin
      { mem[2463:2432] } <= { w_data_i[31:0] };
    end 
    if(N2154) begin
      { mem[2431:2400] } <= { w_data_i[31:0] };
    end 
    if(N2153) begin
      { mem[2399:2368] } <= { w_data_i[31:0] };
    end 
    if(N2152) begin
      { mem[2367:2336] } <= { w_data_i[31:0] };
    end 
    if(N2151) begin
      { mem[2335:2304] } <= { w_data_i[31:0] };
    end 
    if(N2150) begin
      { mem[2303:2272] } <= { w_data_i[31:0] };
    end 
    if(N2149) begin
      { mem[2271:2240] } <= { w_data_i[31:0] };
    end 
    if(N2148) begin
      { mem[2239:2208] } <= { w_data_i[31:0] };
    end 
    if(N2147) begin
      { mem[2207:2176] } <= { w_data_i[31:0] };
    end 
    if(N2146) begin
      { mem[2175:2144] } <= { w_data_i[31:0] };
    end 
    if(N2145) begin
      { mem[2143:2112] } <= { w_data_i[31:0] };
    end 
    if(N2144) begin
      { mem[2111:2080] } <= { w_data_i[31:0] };
    end 
    if(N2143) begin
      { mem[2079:2048] } <= { w_data_i[31:0] };
    end 
    if(N2142) begin
      { mem[2047:2016] } <= { w_data_i[31:0] };
    end 
    if(N2141) begin
      { mem[2015:1984] } <= { w_data_i[31:0] };
    end 
    if(N2140) begin
      { mem[1983:1952] } <= { w_data_i[31:0] };
    end 
    if(N2139) begin
      { mem[1951:1920] } <= { w_data_i[31:0] };
    end 
    if(N2138) begin
      { mem[1919:1888] } <= { w_data_i[31:0] };
    end 
    if(N2137) begin
      { mem[1887:1856] } <= { w_data_i[31:0] };
    end 
    if(N2136) begin
      { mem[1855:1824] } <= { w_data_i[31:0] };
    end 
    if(N2135) begin
      { mem[1823:1792] } <= { w_data_i[31:0] };
    end 
    if(N2134) begin
      { mem[1791:1760] } <= { w_data_i[31:0] };
    end 
    if(N2133) begin
      { mem[1759:1728] } <= { w_data_i[31:0] };
    end 
    if(N2132) begin
      { mem[1727:1696] } <= { w_data_i[31:0] };
    end 
    if(N2131) begin
      { mem[1695:1664] } <= { w_data_i[31:0] };
    end 
    if(N2130) begin
      { mem[1663:1632] } <= { w_data_i[31:0] };
    end 
    if(N2129) begin
      { mem[1631:1600] } <= { w_data_i[31:0] };
    end 
    if(N2128) begin
      { mem[1599:1568] } <= { w_data_i[31:0] };
    end 
    if(N2127) begin
      { mem[1567:1536] } <= { w_data_i[31:0] };
    end 
    if(N2126) begin
      { mem[1535:1504] } <= { w_data_i[31:0] };
    end 
    if(N2125) begin
      { mem[1503:1472] } <= { w_data_i[31:0] };
    end 
    if(N2124) begin
      { mem[1471:1440] } <= { w_data_i[31:0] };
    end 
    if(N2123) begin
      { mem[1439:1408] } <= { w_data_i[31:0] };
    end 
    if(N2122) begin
      { mem[1407:1376] } <= { w_data_i[31:0] };
    end 
    if(N2121) begin
      { mem[1375:1344] } <= { w_data_i[31:0] };
    end 
    if(N2120) begin
      { mem[1343:1312] } <= { w_data_i[31:0] };
    end 
    if(N2119) begin
      { mem[1311:1280] } <= { w_data_i[31:0] };
    end 
    if(N2118) begin
      { mem[1279:1248] } <= { w_data_i[31:0] };
    end 
    if(N2117) begin
      { mem[1247:1216] } <= { w_data_i[31:0] };
    end 
    if(N2116) begin
      { mem[1215:1184] } <= { w_data_i[31:0] };
    end 
    if(N2115) begin
      { mem[1183:1152] } <= { w_data_i[31:0] };
    end 
    if(N2114) begin
      { mem[1151:1120] } <= { w_data_i[31:0] };
    end 
    if(N2113) begin
      { mem[1119:1088] } <= { w_data_i[31:0] };
    end 
    if(N2112) begin
      { mem[1087:1056] } <= { w_data_i[31:0] };
    end 
    if(N2111) begin
      { mem[1055:1024] } <= { w_data_i[31:0] };
    end 
    if(N2110) begin
      { mem[1023:992] } <= { w_data_i[31:0] };
    end 
    if(N2109) begin
      { mem[991:960] } <= { w_data_i[31:0] };
    end 
    if(N2108) begin
      { mem[959:928] } <= { w_data_i[31:0] };
    end 
    if(N2107) begin
      { mem[927:896] } <= { w_data_i[31:0] };
    end 
    if(N2106) begin
      { mem[895:864] } <= { w_data_i[31:0] };
    end 
    if(N2105) begin
      { mem[863:832] } <= { w_data_i[31:0] };
    end 
    if(N2104) begin
      { mem[831:800] } <= { w_data_i[31:0] };
    end 
    if(N2103) begin
      { mem[799:768] } <= { w_data_i[31:0] };
    end 
    if(N2102) begin
      { mem[767:736] } <= { w_data_i[31:0] };
    end 
    if(N2101) begin
      { mem[735:704] } <= { w_data_i[31:0] };
    end 
    if(N2100) begin
      { mem[703:672] } <= { w_data_i[31:0] };
    end 
    if(N2099) begin
      { mem[671:640] } <= { w_data_i[31:0] };
    end 
    if(N2098) begin
      { mem[639:608] } <= { w_data_i[31:0] };
    end 
    if(N2097) begin
      { mem[607:576] } <= { w_data_i[31:0] };
    end 
    if(N2096) begin
      { mem[575:544] } <= { w_data_i[31:0] };
    end 
    if(N2095) begin
      { mem[543:512] } <= { w_data_i[31:0] };
    end 
    if(N2094) begin
      { mem[511:480] } <= { w_data_i[31:0] };
    end 
    if(N2093) begin
      { mem[479:448] } <= { w_data_i[31:0] };
    end 
    if(N2092) begin
      { mem[447:416] } <= { w_data_i[31:0] };
    end 
    if(N2091) begin
      { mem[415:384] } <= { w_data_i[31:0] };
    end 
    if(N2090) begin
      { mem[383:352] } <= { w_data_i[31:0] };
    end 
    if(N2089) begin
      { mem[351:320] } <= { w_data_i[31:0] };
    end 
    if(N2088) begin
      { mem[319:288] } <= { w_data_i[31:0] };
    end 
    if(N2087) begin
      { mem[287:256] } <= { w_data_i[31:0] };
    end 
    if(N2086) begin
      { mem[255:224] } <= { w_data_i[31:0] };
    end 
    if(N2085) begin
      { mem[223:192] } <= { w_data_i[31:0] };
    end 
    if(N2084) begin
      { mem[191:160] } <= { w_data_i[31:0] };
    end 
    if(N2083) begin
      { mem[159:128] } <= { w_data_i[31:0] };
    end 
    if(N2082) begin
      { mem[127:96] } <= { w_data_i[31:0] };
    end 
    if(N2081) begin
      { mem[95:64] } <= { w_data_i[31:0] };
    end 
    if(N2080) begin
      { mem[63:32] } <= { w_data_i[31:0] };
    end 
    if(N2079) begin
      { mem[31:0] } <= { w_data_i[31:0] };
    end 
    if(N2078) begin
      { valid[1023:1023] } <= { N1045 };
    end 
    if(N2077) begin
      { valid[1022:1022] } <= { N1045 };
    end 
    if(N2076) begin
      { valid[1021:1021] } <= { N1045 };
    end 
    if(N2075) begin
      { valid[1020:1020] } <= { N1045 };
    end 
    if(N2074) begin
      { valid[1019:1019] } <= { N1045 };
    end 
    if(N2073) begin
      { valid[1018:1018] } <= { N1045 };
    end 
    if(N2072) begin
      { valid[1017:1017] } <= { N1045 };
    end 
    if(N2071) begin
      { valid[1016:1016] } <= { N1045 };
    end 
    if(N2070) begin
      { valid[1015:1015] } <= { N1045 };
    end 
    if(N2069) begin
      { valid[1014:1014] } <= { N1045 };
    end 
    if(N2068) begin
      { valid[1013:1013] } <= { N1045 };
    end 
    if(N2067) begin
      { valid[1012:1012] } <= { N1045 };
    end 
    if(N2066) begin
      { valid[1011:1011] } <= { N1045 };
    end 
    if(N2065) begin
      { valid[1010:1010] } <= { N1045 };
    end 
    if(N2064) begin
      { valid[1009:1009] } <= { N1045 };
    end 
    if(N2063) begin
      { valid[1008:1008] } <= { N1045 };
    end 
    if(N2062) begin
      { valid[1007:1007] } <= { N1045 };
    end 
    if(N2061) begin
      { valid[1006:1006] } <= { N1045 };
    end 
    if(N2060) begin
      { valid[1005:1005] } <= { N1045 };
    end 
    if(N2059) begin
      { valid[1004:1004] } <= { N1045 };
    end 
    if(N2058) begin
      { valid[1003:1003] } <= { N1045 };
    end 
    if(N2057) begin
      { valid[1002:1002] } <= { N1045 };
    end 
    if(N2056) begin
      { valid[1001:1001] } <= { N1045 };
    end 
    if(N2055) begin
      { valid[1000:1000] } <= { N1045 };
    end 
    if(N2054) begin
      { valid[999:999] } <= { N1045 };
    end 
    if(N2053) begin
      { valid[998:998] } <= { N1045 };
    end 
    if(N2052) begin
      { valid[997:997] } <= { N1045 };
    end 
    if(N2051) begin
      { valid[996:996] } <= { N1045 };
    end 
    if(N2050) begin
      { valid[995:995] } <= { N1045 };
    end 
    if(N2049) begin
      { valid[994:994] } <= { N1045 };
    end 
    if(N2048) begin
      { valid[993:993] } <= { N1045 };
    end 
    if(N2047) begin
      { valid[992:992] } <= { N1045 };
    end 
    if(N2046) begin
      { valid[991:991] } <= { N1045 };
    end 
    if(N2045) begin
      { valid[990:990] } <= { N1045 };
    end 
    if(N2044) begin
      { valid[989:989] } <= { N1045 };
    end 
    if(N2043) begin
      { valid[988:988] } <= { N1045 };
    end 
    if(N2042) begin
      { valid[987:987] } <= { N1045 };
    end 
    if(N2041) begin
      { valid[986:986] } <= { N1045 };
    end 
    if(N2040) begin
      { valid[985:985] } <= { N1045 };
    end 
    if(N2039) begin
      { valid[984:984] } <= { N1045 };
    end 
    if(N2038) begin
      { valid[983:983] } <= { N1045 };
    end 
    if(N2037) begin
      { valid[982:982] } <= { N1045 };
    end 
    if(N2036) begin
      { valid[981:981] } <= { N1045 };
    end 
    if(N2035) begin
      { valid[980:980] } <= { N1045 };
    end 
    if(N2034) begin
      { valid[979:979] } <= { N1045 };
    end 
    if(N2033) begin
      { valid[978:978] } <= { N1045 };
    end 
    if(N2032) begin
      { valid[977:977] } <= { N1045 };
    end 
    if(N2031) begin
      { valid[976:976] } <= { N1045 };
    end 
    if(N2030) begin
      { valid[975:975] } <= { N1045 };
    end 
    if(N2029) begin
      { valid[974:974] } <= { N1045 };
    end 
    if(N2028) begin
      { valid[973:973] } <= { N1045 };
    end 
    if(N2027) begin
      { valid[972:972] } <= { N1045 };
    end 
    if(N2026) begin
      { valid[971:971] } <= { N1045 };
    end 
    if(N2025) begin
      { valid[970:970] } <= { N1045 };
    end 
    if(N2024) begin
      { valid[969:969] } <= { N1045 };
    end 
    if(N2023) begin
      { valid[968:968] } <= { N1045 };
    end 
    if(N2022) begin
      { valid[967:967] } <= { N1045 };
    end 
    if(N2021) begin
      { valid[966:966] } <= { N1045 };
    end 
    if(N2020) begin
      { valid[965:965] } <= { N1045 };
    end 
    if(N2019) begin
      { valid[964:964] } <= { N1045 };
    end 
    if(N2018) begin
      { valid[963:963] } <= { N1045 };
    end 
    if(N2017) begin
      { valid[962:962] } <= { N1045 };
    end 
    if(N2016) begin
      { valid[961:961] } <= { N1045 };
    end 
    if(N2015) begin
      { valid[960:960] } <= { N1045 };
    end 
    if(N2014) begin
      { valid[959:959] } <= { N1045 };
    end 
    if(N2013) begin
      { valid[958:958] } <= { N1045 };
    end 
    if(N2012) begin
      { valid[957:957] } <= { N1045 };
    end 
    if(N2011) begin
      { valid[956:956] } <= { N1045 };
    end 
    if(N2010) begin
      { valid[955:955] } <= { N1045 };
    end 
    if(N2009) begin
      { valid[954:954] } <= { N1045 };
    end 
    if(N2008) begin
      { valid[953:953] } <= { N1045 };
    end 
    if(N2007) begin
      { valid[952:952] } <= { N1045 };
    end 
    if(N2006) begin
      { valid[951:951] } <= { N1045 };
    end 
    if(N2005) begin
      { valid[950:950] } <= { N1045 };
    end 
    if(N2004) begin
      { valid[949:949] } <= { N1045 };
    end 
    if(N2003) begin
      { valid[948:948] } <= { N1045 };
    end 
    if(N2002) begin
      { valid[947:947] } <= { N1045 };
    end 
    if(N2001) begin
      { valid[946:946] } <= { N1045 };
    end 
    if(N2000) begin
      { valid[945:945] } <= { N1045 };
    end 
    if(N1999) begin
      { valid[944:944] } <= { N1045 };
    end 
    if(N1998) begin
      { valid[943:943] } <= { N1045 };
    end 
    if(N1997) begin
      { valid[942:942] } <= { N1045 };
    end 
    if(N1996) begin
      { valid[941:941] } <= { N1045 };
    end 
    if(N1995) begin
      { valid[940:940] } <= { N1045 };
    end 
    if(N1994) begin
      { valid[939:939] } <= { N1045 };
    end 
    if(N1993) begin
      { valid[938:938] } <= { N1045 };
    end 
    if(N1992) begin
      { valid[937:937] } <= { N1045 };
    end 
    if(N1991) begin
      { valid[936:936] } <= { N1045 };
    end 
    if(N1990) begin
      { valid[935:935] } <= { N1045 };
    end 
    if(N1989) begin
      { valid[934:934] } <= { N1045 };
    end 
    if(N1988) begin
      { valid[933:933] } <= { N1045 };
    end 
    if(N1987) begin
      { valid[932:932] } <= { N1045 };
    end 
    if(N1986) begin
      { valid[931:931] } <= { N1045 };
    end 
    if(N1985) begin
      { valid[930:930] } <= { N1045 };
    end 
    if(N1984) begin
      { valid[929:929] } <= { N1045 };
    end 
    if(N1983) begin
      { valid[928:928] } <= { N1045 };
    end 
    if(N1982) begin
      { valid[927:927] } <= { N1045 };
    end 
    if(N1981) begin
      { valid[926:926] } <= { N1045 };
    end 
    if(N1980) begin
      { valid[925:925] } <= { N1045 };
    end 
    if(N1979) begin
      { valid[924:924] } <= { N1047 };
    end 
    if(N1978) begin
      { valid[923:923] } <= { N1047 };
    end 
    if(N1977) begin
      { valid[922:922] } <= { N1047 };
    end 
    if(N1976) begin
      { valid[921:921] } <= { N1047 };
    end 
    if(N1975) begin
      { valid[920:920] } <= { N1047 };
    end 
    if(N1974) begin
      { valid[919:919] } <= { N1047 };
    end 
    if(N1973) begin
      { valid[918:918] } <= { N1047 };
    end 
    if(N1972) begin
      { valid[917:917] } <= { N1047 };
    end 
    if(N1971) begin
      { valid[916:916] } <= { N1047 };
    end 
    if(N1970) begin
      { valid[915:915] } <= { N1047 };
    end 
    if(N1969) begin
      { valid[914:914] } <= { N1047 };
    end 
    if(N1968) begin
      { valid[913:913] } <= { N1047 };
    end 
    if(N1967) begin
      { valid[912:912] } <= { N1047 };
    end 
    if(N1966) begin
      { valid[911:911] } <= { N1047 };
    end 
    if(N1965) begin
      { valid[910:910] } <= { N1047 };
    end 
    if(N1964) begin
      { valid[909:909] } <= { N1047 };
    end 
    if(N1963) begin
      { valid[908:908] } <= { N1047 };
    end 
    if(N1962) begin
      { valid[907:907] } <= { N1047 };
    end 
    if(N1961) begin
      { valid[906:906] } <= { N1047 };
    end 
    if(N1960) begin
      { valid[905:905] } <= { N1047 };
    end 
    if(N1959) begin
      { valid[904:904] } <= { N1047 };
    end 
    if(N1958) begin
      { valid[903:903] } <= { N1047 };
    end 
    if(N1957) begin
      { valid[902:902] } <= { N1047 };
    end 
    if(N1956) begin
      { valid[901:901] } <= { N1047 };
    end 
    if(N1955) begin
      { valid[900:900] } <= { N1047 };
    end 
    if(N1954) begin
      { valid[899:899] } <= { N1047 };
    end 
    if(N1953) begin
      { valid[898:898] } <= { N1047 };
    end 
    if(N1952) begin
      { valid[897:897] } <= { N1047 };
    end 
    if(N1951) begin
      { valid[896:896] } <= { N1047 };
    end 
    if(N1950) begin
      { valid[895:895] } <= { N1047 };
    end 
    if(N1949) begin
      { valid[894:894] } <= { N1047 };
    end 
    if(N1948) begin
      { valid[893:893] } <= { N1047 };
    end 
    if(N1947) begin
      { valid[892:892] } <= { N1047 };
    end 
    if(N1946) begin
      { valid[891:891] } <= { N1047 };
    end 
    if(N1945) begin
      { valid[890:890] } <= { N1047 };
    end 
    if(N1944) begin
      { valid[889:889] } <= { N1047 };
    end 
    if(N1943) begin
      { valid[888:888] } <= { N1047 };
    end 
    if(N1942) begin
      { valid[887:887] } <= { N1047 };
    end 
    if(N1941) begin
      { valid[886:886] } <= { N1047 };
    end 
    if(N1940) begin
      { valid[885:885] } <= { N1047 };
    end 
    if(N1939) begin
      { valid[884:884] } <= { N1047 };
    end 
    if(N1938) begin
      { valid[883:883] } <= { N1047 };
    end 
    if(N1937) begin
      { valid[882:882] } <= { N1047 };
    end 
    if(N1936) begin
      { valid[881:881] } <= { N1047 };
    end 
    if(N1935) begin
      { valid[880:880] } <= { N1047 };
    end 
    if(N1934) begin
      { valid[879:879] } <= { N1047 };
    end 
    if(N1933) begin
      { valid[878:878] } <= { N1047 };
    end 
    if(N1932) begin
      { valid[877:877] } <= { N1047 };
    end 
    if(N1931) begin
      { valid[876:876] } <= { N1047 };
    end 
    if(N1930) begin
      { valid[875:875] } <= { N1047 };
    end 
    if(N1929) begin
      { valid[874:874] } <= { N1047 };
    end 
    if(N1928) begin
      { valid[873:873] } <= { N1047 };
    end 
    if(N1927) begin
      { valid[872:872] } <= { N1047 };
    end 
    if(N1926) begin
      { valid[871:871] } <= { N1047 };
    end 
    if(N1925) begin
      { valid[870:870] } <= { N1047 };
    end 
    if(N1924) begin
      { valid[869:869] } <= { N1047 };
    end 
    if(N1923) begin
      { valid[868:868] } <= { N1047 };
    end 
    if(N1922) begin
      { valid[867:867] } <= { N1047 };
    end 
    if(N1921) begin
      { valid[866:866] } <= { N1047 };
    end 
    if(N1920) begin
      { valid[865:865] } <= { N1047 };
    end 
    if(N1919) begin
      { valid[864:864] } <= { N1047 };
    end 
    if(N1918) begin
      { valid[863:863] } <= { N1047 };
    end 
    if(N1917) begin
      { valid[862:862] } <= { N1047 };
    end 
    if(N1916) begin
      { valid[861:861] } <= { N1047 };
    end 
    if(N1915) begin
      { valid[860:860] } <= { N1047 };
    end 
    if(N1914) begin
      { valid[859:859] } <= { N1047 };
    end 
    if(N1913) begin
      { valid[858:858] } <= { N1047 };
    end 
    if(N1912) begin
      { valid[857:857] } <= { N1047 };
    end 
    if(N1911) begin
      { valid[856:856] } <= { N1047 };
    end 
    if(N1910) begin
      { valid[855:855] } <= { N1047 };
    end 
    if(N1909) begin
      { valid[854:854] } <= { N1047 };
    end 
    if(N1908) begin
      { valid[853:853] } <= { N1047 };
    end 
    if(N1907) begin
      { valid[852:852] } <= { N1047 };
    end 
    if(N1906) begin
      { valid[851:851] } <= { N1047 };
    end 
    if(N1905) begin
      { valid[850:850] } <= { N1047 };
    end 
    if(N1904) begin
      { valid[849:849] } <= { N1047 };
    end 
    if(N1903) begin
      { valid[848:848] } <= { N1047 };
    end 
    if(N1902) begin
      { valid[847:847] } <= { N1047 };
    end 
    if(N1901) begin
      { valid[846:846] } <= { N1047 };
    end 
    if(N1900) begin
      { valid[845:845] } <= { N1047 };
    end 
    if(N1899) begin
      { valid[844:844] } <= { N1047 };
    end 
    if(N1898) begin
      { valid[843:843] } <= { N1047 };
    end 
    if(N1897) begin
      { valid[842:842] } <= { N1047 };
    end 
    if(N1896) begin
      { valid[841:841] } <= { N1047 };
    end 
    if(N1895) begin
      { valid[840:840] } <= { N1047 };
    end 
    if(N1894) begin
      { valid[839:839] } <= { N1047 };
    end 
    if(N1893) begin
      { valid[838:838] } <= { N1047 };
    end 
    if(N1892) begin
      { valid[837:837] } <= { N1047 };
    end 
    if(N1891) begin
      { valid[836:836] } <= { N1047 };
    end 
    if(N1890) begin
      { valid[835:835] } <= { N1047 };
    end 
    if(N1889) begin
      { valid[834:834] } <= { N1047 };
    end 
    if(N1888) begin
      { valid[833:833] } <= { N1047 };
    end 
    if(N1887) begin
      { valid[832:832] } <= { N1047 };
    end 
    if(N1886) begin
      { valid[831:831] } <= { N1047 };
    end 
    if(N1885) begin
      { valid[830:830] } <= { N1047 };
    end 
    if(N1884) begin
      { valid[829:829] } <= { N1047 };
    end 
    if(N1883) begin
      { valid[828:828] } <= { N1047 };
    end 
    if(N1882) begin
      { valid[827:827] } <= { N1047 };
    end 
    if(N1881) begin
      { valid[826:826] } <= { N1047 };
    end 
    if(N1880) begin
      { valid[825:825] } <= { N1049 };
    end 
    if(N1879) begin
      { valid[824:824] } <= { N1049 };
    end 
    if(N1878) begin
      { valid[823:823] } <= { N1049 };
    end 
    if(N1877) begin
      { valid[822:822] } <= { N1049 };
    end 
    if(N1876) begin
      { valid[821:821] } <= { N1049 };
    end 
    if(N1875) begin
      { valid[820:820] } <= { N1049 };
    end 
    if(N1874) begin
      { valid[819:819] } <= { N1049 };
    end 
    if(N1873) begin
      { valid[818:818] } <= { N1049 };
    end 
    if(N1872) begin
      { valid[817:817] } <= { N1049 };
    end 
    if(N1871) begin
      { valid[816:816] } <= { N1049 };
    end 
    if(N1870) begin
      { valid[815:815] } <= { N1049 };
    end 
    if(N1869) begin
      { valid[814:814] } <= { N1049 };
    end 
    if(N1868) begin
      { valid[813:813] } <= { N1049 };
    end 
    if(N1867) begin
      { valid[812:812] } <= { N1049 };
    end 
    if(N1866) begin
      { valid[811:811] } <= { N1049 };
    end 
    if(N1865) begin
      { valid[810:810] } <= { N1049 };
    end 
    if(N1864) begin
      { valid[809:809] } <= { N1049 };
    end 
    if(N1863) begin
      { valid[808:808] } <= { N1049 };
    end 
    if(N1862) begin
      { valid[807:807] } <= { N1049 };
    end 
    if(N1861) begin
      { valid[806:806] } <= { N1049 };
    end 
    if(N1860) begin
      { valid[805:805] } <= { N1049 };
    end 
    if(N1859) begin
      { valid[804:804] } <= { N1049 };
    end 
    if(N1858) begin
      { valid[803:803] } <= { N1049 };
    end 
    if(N1857) begin
      { valid[802:802] } <= { N1049 };
    end 
    if(N1856) begin
      { valid[801:801] } <= { N1049 };
    end 
    if(N1855) begin
      { valid[800:800] } <= { N1049 };
    end 
    if(N1854) begin
      { valid[799:799] } <= { N1049 };
    end 
    if(N1853) begin
      { valid[798:798] } <= { N1049 };
    end 
    if(N1852) begin
      { valid[797:797] } <= { N1049 };
    end 
    if(N1851) begin
      { valid[796:796] } <= { N1049 };
    end 
    if(N1850) begin
      { valid[795:795] } <= { N1049 };
    end 
    if(N1849) begin
      { valid[794:794] } <= { N1049 };
    end 
    if(N1848) begin
      { valid[793:793] } <= { N1049 };
    end 
    if(N1847) begin
      { valid[792:792] } <= { N1049 };
    end 
    if(N1846) begin
      { valid[791:791] } <= { N1049 };
    end 
    if(N1845) begin
      { valid[790:790] } <= { N1049 };
    end 
    if(N1844) begin
      { valid[789:789] } <= { N1049 };
    end 
    if(N1843) begin
      { valid[788:788] } <= { N1049 };
    end 
    if(N1842) begin
      { valid[787:787] } <= { N1049 };
    end 
    if(N1841) begin
      { valid[786:786] } <= { N1049 };
    end 
    if(N1840) begin
      { valid[785:785] } <= { N1049 };
    end 
    if(N1839) begin
      { valid[784:784] } <= { N1049 };
    end 
    if(N1838) begin
      { valid[783:783] } <= { N1049 };
    end 
    if(N1837) begin
      { valid[782:782] } <= { N1049 };
    end 
    if(N1836) begin
      { valid[781:781] } <= { N1049 };
    end 
    if(N1835) begin
      { valid[780:780] } <= { N1049 };
    end 
    if(N1834) begin
      { valid[779:779] } <= { N1049 };
    end 
    if(N1833) begin
      { valid[778:778] } <= { N1049 };
    end 
    if(N1832) begin
      { valid[777:777] } <= { N1049 };
    end 
    if(N1831) begin
      { valid[776:776] } <= { N1049 };
    end 
    if(N1830) begin
      { valid[775:775] } <= { N1049 };
    end 
    if(N1829) begin
      { valid[774:774] } <= { N1049 };
    end 
    if(N1828) begin
      { valid[773:773] } <= { N1049 };
    end 
    if(N1827) begin
      { valid[772:772] } <= { N1049 };
    end 
    if(N1826) begin
      { valid[771:771] } <= { N1049 };
    end 
    if(N1825) begin
      { valid[770:770] } <= { N1049 };
    end 
    if(N1824) begin
      { valid[769:769] } <= { N1049 };
    end 
    if(N1823) begin
      { valid[768:768] } <= { N1049 };
    end 
    if(N1822) begin
      { valid[767:767] } <= { N1049 };
    end 
    if(N1821) begin
      { valid[766:766] } <= { N1049 };
    end 
    if(N1820) begin
      { valid[765:765] } <= { N1049 };
    end 
    if(N1819) begin
      { valid[764:764] } <= { N1049 };
    end 
    if(N1818) begin
      { valid[763:763] } <= { N1049 };
    end 
    if(N1817) begin
      { valid[762:762] } <= { N1049 };
    end 
    if(N1816) begin
      { valid[761:761] } <= { N1049 };
    end 
    if(N1815) begin
      { valid[760:760] } <= { N1049 };
    end 
    if(N1814) begin
      { valid[759:759] } <= { N1049 };
    end 
    if(N1813) begin
      { valid[758:758] } <= { N1049 };
    end 
    if(N1812) begin
      { valid[757:757] } <= { N1049 };
    end 
    if(N1811) begin
      { valid[756:756] } <= { N1049 };
    end 
    if(N1810) begin
      { valid[755:755] } <= { N1049 };
    end 
    if(N1809) begin
      { valid[754:754] } <= { N1049 };
    end 
    if(N1808) begin
      { valid[753:753] } <= { N1049 };
    end 
    if(N1807) begin
      { valid[752:752] } <= { N1049 };
    end 
    if(N1806) begin
      { valid[751:751] } <= { N1049 };
    end 
    if(N1805) begin
      { valid[750:750] } <= { N1049 };
    end 
    if(N1804) begin
      { valid[749:749] } <= { N1049 };
    end 
    if(N1803) begin
      { valid[748:748] } <= { N1049 };
    end 
    if(N1802) begin
      { valid[747:747] } <= { N1049 };
    end 
    if(N1801) begin
      { valid[746:746] } <= { N1049 };
    end 
    if(N1800) begin
      { valid[745:745] } <= { N1049 };
    end 
    if(N1799) begin
      { valid[744:744] } <= { N1049 };
    end 
    if(N1798) begin
      { valid[743:743] } <= { N1049 };
    end 
    if(N1797) begin
      { valid[742:742] } <= { N1049 };
    end 
    if(N1796) begin
      { valid[741:741] } <= { N1049 };
    end 
    if(N1795) begin
      { valid[740:740] } <= { N1049 };
    end 
    if(N1794) begin
      { valid[739:739] } <= { N1049 };
    end 
    if(N1793) begin
      { valid[738:738] } <= { N1049 };
    end 
    if(N1792) begin
      { valid[737:737] } <= { N1049 };
    end 
    if(N1791) begin
      { valid[736:736] } <= { N1049 };
    end 
    if(N1790) begin
      { valid[735:735] } <= { N1049 };
    end 
    if(N1789) begin
      { valid[734:734] } <= { N1049 };
    end 
    if(N1788) begin
      { valid[733:733] } <= { N1049 };
    end 
    if(N1787) begin
      { valid[732:732] } <= { N1049 };
    end 
    if(N1786) begin
      { valid[731:731] } <= { N1049 };
    end 
    if(N1785) begin
      { valid[730:730] } <= { N1049 };
    end 
    if(N1784) begin
      { valid[729:729] } <= { N1049 };
    end 
    if(N1783) begin
      { valid[728:728] } <= { N1049 };
    end 
    if(N1782) begin
      { valid[727:727] } <= { N1049 };
    end 
    if(N1781) begin
      { valid[726:726] } <= { N1051 };
    end 
    if(N1780) begin
      { valid[725:725] } <= { N1051 };
    end 
    if(N1779) begin
      { valid[724:724] } <= { N1051 };
    end 
    if(N1778) begin
      { valid[723:723] } <= { N1051 };
    end 
    if(N1777) begin
      { valid[722:722] } <= { N1051 };
    end 
    if(N1776) begin
      { valid[721:721] } <= { N1051 };
    end 
    if(N1775) begin
      { valid[720:720] } <= { N1051 };
    end 
    if(N1774) begin
      { valid[719:719] } <= { N1051 };
    end 
    if(N1773) begin
      { valid[718:718] } <= { N1051 };
    end 
    if(N1772) begin
      { valid[717:717] } <= { N1051 };
    end 
    if(N1771) begin
      { valid[716:716] } <= { N1051 };
    end 
    if(N1770) begin
      { valid[715:715] } <= { N1051 };
    end 
    if(N1769) begin
      { valid[714:714] } <= { N1051 };
    end 
    if(N1768) begin
      { valid[713:713] } <= { N1051 };
    end 
    if(N1767) begin
      { valid[712:712] } <= { N1051 };
    end 
    if(N1766) begin
      { valid[711:711] } <= { N1051 };
    end 
    if(N1765) begin
      { valid[710:710] } <= { N1051 };
    end 
    if(N1764) begin
      { valid[709:709] } <= { N1051 };
    end 
    if(N1763) begin
      { valid[708:708] } <= { N1051 };
    end 
    if(N1762) begin
      { valid[707:707] } <= { N1051 };
    end 
    if(N1761) begin
      { valid[706:706] } <= { N1051 };
    end 
    if(N1760) begin
      { valid[705:705] } <= { N1051 };
    end 
    if(N1759) begin
      { valid[704:704] } <= { N1051 };
    end 
    if(N1758) begin
      { valid[703:703] } <= { N1051 };
    end 
    if(N1757) begin
      { valid[702:702] } <= { N1051 };
    end 
    if(N1756) begin
      { valid[701:701] } <= { N1051 };
    end 
    if(N1755) begin
      { valid[700:700] } <= { N1051 };
    end 
    if(N1754) begin
      { valid[699:699] } <= { N1051 };
    end 
    if(N1753) begin
      { valid[698:698] } <= { N1051 };
    end 
    if(N1752) begin
      { valid[697:697] } <= { N1051 };
    end 
    if(N1751) begin
      { valid[696:696] } <= { N1051 };
    end 
    if(N1750) begin
      { valid[695:695] } <= { N1051 };
    end 
    if(N1749) begin
      { valid[694:694] } <= { N1051 };
    end 
    if(N1748) begin
      { valid[693:693] } <= { N1051 };
    end 
    if(N1747) begin
      { valid[692:692] } <= { N1051 };
    end 
    if(N1746) begin
      { valid[691:691] } <= { N1051 };
    end 
    if(N1745) begin
      { valid[690:690] } <= { N1051 };
    end 
    if(N1744) begin
      { valid[689:689] } <= { N1051 };
    end 
    if(N1743) begin
      { valid[688:688] } <= { N1051 };
    end 
    if(N1742) begin
      { valid[687:687] } <= { N1051 };
    end 
    if(N1741) begin
      { valid[686:686] } <= { N1051 };
    end 
    if(N1740) begin
      { valid[685:685] } <= { N1051 };
    end 
    if(N1739) begin
      { valid[684:684] } <= { N1051 };
    end 
    if(N1738) begin
      { valid[683:683] } <= { N1051 };
    end 
    if(N1737) begin
      { valid[682:682] } <= { N1051 };
    end 
    if(N1736) begin
      { valid[681:681] } <= { N1051 };
    end 
    if(N1735) begin
      { valid[680:680] } <= { N1051 };
    end 
    if(N1734) begin
      { valid[679:679] } <= { N1051 };
    end 
    if(N1733) begin
      { valid[678:678] } <= { N1051 };
    end 
    if(N1732) begin
      { valid[677:677] } <= { N1051 };
    end 
    if(N1731) begin
      { valid[676:676] } <= { N1051 };
    end 
    if(N1730) begin
      { valid[675:675] } <= { N1051 };
    end 
    if(N1729) begin
      { valid[674:674] } <= { N1051 };
    end 
    if(N1728) begin
      { valid[673:673] } <= { N1051 };
    end 
    if(N1727) begin
      { valid[672:672] } <= { N1051 };
    end 
    if(N1726) begin
      { valid[671:671] } <= { N1051 };
    end 
    if(N1725) begin
      { valid[670:670] } <= { N1051 };
    end 
    if(N1724) begin
      { valid[669:669] } <= { N1051 };
    end 
    if(N1723) begin
      { valid[668:668] } <= { N1051 };
    end 
    if(N1722) begin
      { valid[667:667] } <= { N1051 };
    end 
    if(N1721) begin
      { valid[666:666] } <= { N1051 };
    end 
    if(N1720) begin
      { valid[665:665] } <= { N1051 };
    end 
    if(N1719) begin
      { valid[664:664] } <= { N1051 };
    end 
    if(N1718) begin
      { valid[663:663] } <= { N1051 };
    end 
    if(N1717) begin
      { valid[662:662] } <= { N1051 };
    end 
    if(N1716) begin
      { valid[661:661] } <= { N1051 };
    end 
    if(N1715) begin
      { valid[660:660] } <= { N1051 };
    end 
    if(N1714) begin
      { valid[659:659] } <= { N1051 };
    end 
    if(N1713) begin
      { valid[658:658] } <= { N1051 };
    end 
    if(N1712) begin
      { valid[657:657] } <= { N1051 };
    end 
    if(N1711) begin
      { valid[656:656] } <= { N1051 };
    end 
    if(N1710) begin
      { valid[655:655] } <= { N1051 };
    end 
    if(N1709) begin
      { valid[654:654] } <= { N1051 };
    end 
    if(N1708) begin
      { valid[653:653] } <= { N1051 };
    end 
    if(N1707) begin
      { valid[652:652] } <= { N1051 };
    end 
    if(N1706) begin
      { valid[651:651] } <= { N1051 };
    end 
    if(N1705) begin
      { valid[650:650] } <= { N1051 };
    end 
    if(N1704) begin
      { valid[649:649] } <= { N1051 };
    end 
    if(N1703) begin
      { valid[648:648] } <= { N1051 };
    end 
    if(N1702) begin
      { valid[647:647] } <= { N1051 };
    end 
    if(N1701) begin
      { valid[646:646] } <= { N1051 };
    end 
    if(N1700) begin
      { valid[645:645] } <= { N1051 };
    end 
    if(N1699) begin
      { valid[644:644] } <= { N1051 };
    end 
    if(N1698) begin
      { valid[643:643] } <= { N1051 };
    end 
    if(N1697) begin
      { valid[642:642] } <= { N1051 };
    end 
    if(N1696) begin
      { valid[641:641] } <= { N1051 };
    end 
    if(N1695) begin
      { valid[640:640] } <= { N1051 };
    end 
    if(N1694) begin
      { valid[639:639] } <= { N1051 };
    end 
    if(N1693) begin
      { valid[638:638] } <= { N1051 };
    end 
    if(N1692) begin
      { valid[637:637] } <= { N1051 };
    end 
    if(N1691) begin
      { valid[636:636] } <= { N1051 };
    end 
    if(N1690) begin
      { valid[635:635] } <= { N1051 };
    end 
    if(N1689) begin
      { valid[634:634] } <= { N1051 };
    end 
    if(N1688) begin
      { valid[633:633] } <= { N1051 };
    end 
    if(N1687) begin
      { valid[632:632] } <= { N1051 };
    end 
    if(N1686) begin
      { valid[631:631] } <= { N1051 };
    end 
    if(N1685) begin
      { valid[630:630] } <= { N1051 };
    end 
    if(N1684) begin
      { valid[629:629] } <= { N1051 };
    end 
    if(N1683) begin
      { valid[628:628] } <= { N1051 };
    end 
    if(N1682) begin
      { valid[627:627] } <= { N1053 };
    end 
    if(N1681) begin
      { valid[626:626] } <= { N1053 };
    end 
    if(N1680) begin
      { valid[625:625] } <= { N1053 };
    end 
    if(N1679) begin
      { valid[624:624] } <= { N1053 };
    end 
    if(N1678) begin
      { valid[623:623] } <= { N1053 };
    end 
    if(N1677) begin
      { valid[622:622] } <= { N1053 };
    end 
    if(N1676) begin
      { valid[621:621] } <= { N1053 };
    end 
    if(N1675) begin
      { valid[620:620] } <= { N1053 };
    end 
    if(N1674) begin
      { valid[619:619] } <= { N1053 };
    end 
    if(N1673) begin
      { valid[618:618] } <= { N1053 };
    end 
    if(N1672) begin
      { valid[617:617] } <= { N1053 };
    end 
    if(N1671) begin
      { valid[616:616] } <= { N1053 };
    end 
    if(N1670) begin
      { valid[615:615] } <= { N1053 };
    end 
    if(N1669) begin
      { valid[614:614] } <= { N1053 };
    end 
    if(N1668) begin
      { valid[613:613] } <= { N1053 };
    end 
    if(N1667) begin
      { valid[612:612] } <= { N1053 };
    end 
    if(N1666) begin
      { valid[611:611] } <= { N1053 };
    end 
    if(N1665) begin
      { valid[610:610] } <= { N1053 };
    end 
    if(N1664) begin
      { valid[609:609] } <= { N1053 };
    end 
    if(N1663) begin
      { valid[608:608] } <= { N1053 };
    end 
    if(N1662) begin
      { valid[607:607] } <= { N1053 };
    end 
    if(N1661) begin
      { valid[606:606] } <= { N1053 };
    end 
    if(N1660) begin
      { valid[605:605] } <= { N1053 };
    end 
    if(N1659) begin
      { valid[604:604] } <= { N1053 };
    end 
    if(N1658) begin
      { valid[603:603] } <= { N1053 };
    end 
    if(N1657) begin
      { valid[602:602] } <= { N1053 };
    end 
    if(N1656) begin
      { valid[601:601] } <= { N1053 };
    end 
    if(N1655) begin
      { valid[600:600] } <= { N1053 };
    end 
    if(N1654) begin
      { valid[599:599] } <= { N1053 };
    end 
    if(N1653) begin
      { valid[598:598] } <= { N1053 };
    end 
    if(N1652) begin
      { valid[597:597] } <= { N1053 };
    end 
    if(N1651) begin
      { valid[596:596] } <= { N1053 };
    end 
    if(N1650) begin
      { valid[595:595] } <= { N1053 };
    end 
    if(N1649) begin
      { valid[594:594] } <= { N1053 };
    end 
    if(N1648) begin
      { valid[593:593] } <= { N1053 };
    end 
    if(N1647) begin
      { valid[592:592] } <= { N1053 };
    end 
    if(N1646) begin
      { valid[591:591] } <= { N1053 };
    end 
    if(N1645) begin
      { valid[590:590] } <= { N1053 };
    end 
    if(N1644) begin
      { valid[589:589] } <= { N1053 };
    end 
    if(N1643) begin
      { valid[588:588] } <= { N1053 };
    end 
    if(N1642) begin
      { valid[587:587] } <= { N1053 };
    end 
    if(N1641) begin
      { valid[586:586] } <= { N1053 };
    end 
    if(N1640) begin
      { valid[585:585] } <= { N1053 };
    end 
    if(N1639) begin
      { valid[584:584] } <= { N1053 };
    end 
    if(N1638) begin
      { valid[583:583] } <= { N1053 };
    end 
    if(N1637) begin
      { valid[582:582] } <= { N1053 };
    end 
    if(N1636) begin
      { valid[581:581] } <= { N1053 };
    end 
    if(N1635) begin
      { valid[580:580] } <= { N1053 };
    end 
    if(N1634) begin
      { valid[579:579] } <= { N1053 };
    end 
    if(N1633) begin
      { valid[578:578] } <= { N1053 };
    end 
    if(N1632) begin
      { valid[577:577] } <= { N1053 };
    end 
    if(N1631) begin
      { valid[576:576] } <= { N1053 };
    end 
    if(N1630) begin
      { valid[575:575] } <= { N1053 };
    end 
    if(N1629) begin
      { valid[574:574] } <= { N1053 };
    end 
    if(N1628) begin
      { valid[573:573] } <= { N1053 };
    end 
    if(N1627) begin
      { valid[572:572] } <= { N1053 };
    end 
    if(N1626) begin
      { valid[571:571] } <= { N1053 };
    end 
    if(N1625) begin
      { valid[570:570] } <= { N1053 };
    end 
    if(N1624) begin
      { valid[569:569] } <= { N1053 };
    end 
    if(N1623) begin
      { valid[568:568] } <= { N1053 };
    end 
    if(N1622) begin
      { valid[567:567] } <= { N1053 };
    end 
    if(N1621) begin
      { valid[566:566] } <= { N1053 };
    end 
    if(N1620) begin
      { valid[565:565] } <= { N1053 };
    end 
    if(N1619) begin
      { valid[564:564] } <= { N1053 };
    end 
    if(N1618) begin
      { valid[563:563] } <= { N1053 };
    end 
    if(N1617) begin
      { valid[562:562] } <= { N1053 };
    end 
    if(N1616) begin
      { valid[561:561] } <= { N1053 };
    end 
    if(N1615) begin
      { valid[560:560] } <= { N1053 };
    end 
    if(N1614) begin
      { valid[559:559] } <= { N1053 };
    end 
    if(N1613) begin
      { valid[558:558] } <= { N1053 };
    end 
    if(N1612) begin
      { valid[557:557] } <= { N1053 };
    end 
    if(N1611) begin
      { valid[556:556] } <= { N1053 };
    end 
    if(N1610) begin
      { valid[555:555] } <= { N1053 };
    end 
    if(N1609) begin
      { valid[554:554] } <= { N1053 };
    end 
    if(N1608) begin
      { valid[553:553] } <= { N1053 };
    end 
    if(N1607) begin
      { valid[552:552] } <= { N1053 };
    end 
    if(N1606) begin
      { valid[551:551] } <= { N1053 };
    end 
    if(N1605) begin
      { valid[550:550] } <= { N1053 };
    end 
    if(N1604) begin
      { valid[549:549] } <= { N1053 };
    end 
    if(N1603) begin
      { valid[548:548] } <= { N1053 };
    end 
    if(N1602) begin
      { valid[547:547] } <= { N1053 };
    end 
    if(N1601) begin
      { valid[546:546] } <= { N1053 };
    end 
    if(N1600) begin
      { valid[545:545] } <= { N1053 };
    end 
    if(N1599) begin
      { valid[544:544] } <= { N1053 };
    end 
    if(N1598) begin
      { valid[543:543] } <= { N1053 };
    end 
    if(N1597) begin
      { valid[542:542] } <= { N1053 };
    end 
    if(N1596) begin
      { valid[541:541] } <= { N1053 };
    end 
    if(N1595) begin
      { valid[540:540] } <= { N1053 };
    end 
    if(N1594) begin
      { valid[539:539] } <= { N1053 };
    end 
    if(N1593) begin
      { valid[538:538] } <= { N1053 };
    end 
    if(N1592) begin
      { valid[537:537] } <= { N1053 };
    end 
    if(N1591) begin
      { valid[536:536] } <= { N1053 };
    end 
    if(N1590) begin
      { valid[535:535] } <= { N1053 };
    end 
    if(N1589) begin
      { valid[534:534] } <= { N1053 };
    end 
    if(N1588) begin
      { valid[533:533] } <= { N1053 };
    end 
    if(N1587) begin
      { valid[532:532] } <= { N1053 };
    end 
    if(N1586) begin
      { valid[531:531] } <= { N1053 };
    end 
    if(N1585) begin
      { valid[530:530] } <= { N1053 };
    end 
    if(N1584) begin
      { valid[529:529] } <= { N1053 };
    end 
    if(N1583) begin
      { valid[528:528] } <= { N1055 };
    end 
    if(N1582) begin
      { valid[527:527] } <= { N1055 };
    end 
    if(N1581) begin
      { valid[526:526] } <= { N1055 };
    end 
    if(N1580) begin
      { valid[525:525] } <= { N1055 };
    end 
    if(N1579) begin
      { valid[524:524] } <= { N1055 };
    end 
    if(N1578) begin
      { valid[523:523] } <= { N1055 };
    end 
    if(N1577) begin
      { valid[522:522] } <= { N1055 };
    end 
    if(N1576) begin
      { valid[521:521] } <= { N1055 };
    end 
    if(N1575) begin
      { valid[520:520] } <= { N1055 };
    end 
    if(N1574) begin
      { valid[519:519] } <= { N1055 };
    end 
    if(N1573) begin
      { valid[518:518] } <= { N1055 };
    end 
    if(N1572) begin
      { valid[517:517] } <= { N1055 };
    end 
    if(N1571) begin
      { valid[516:516] } <= { N1055 };
    end 
    if(N1570) begin
      { valid[515:515] } <= { N1055 };
    end 
    if(N1569) begin
      { valid[514:514] } <= { N1055 };
    end 
    if(N1568) begin
      { valid[513:513] } <= { N1055 };
    end 
    if(N1567) begin
      { valid[512:512] } <= { N1055 };
    end 
    if(N1566) begin
      { valid[511:511] } <= { N1055 };
    end 
    if(N1565) begin
      { valid[510:510] } <= { N1055 };
    end 
    if(N1564) begin
      { valid[509:509] } <= { N1055 };
    end 
    if(N1563) begin
      { valid[508:508] } <= { N1055 };
    end 
    if(N1562) begin
      { valid[507:507] } <= { N1055 };
    end 
    if(N1561) begin
      { valid[506:506] } <= { N1055 };
    end 
    if(N1560) begin
      { valid[505:505] } <= { N1055 };
    end 
    if(N1559) begin
      { valid[504:504] } <= { N1055 };
    end 
    if(N1558) begin
      { valid[503:503] } <= { N1055 };
    end 
    if(N1557) begin
      { valid[502:502] } <= { N1055 };
    end 
    if(N1556) begin
      { valid[501:501] } <= { N1055 };
    end 
    if(N1555) begin
      { valid[500:500] } <= { N1055 };
    end 
    if(N1554) begin
      { valid[499:499] } <= { N1055 };
    end 
    if(N1553) begin
      { valid[498:498] } <= { N1055 };
    end 
    if(N1552) begin
      { valid[497:497] } <= { N1055 };
    end 
    if(N1551) begin
      { valid[496:496] } <= { N1055 };
    end 
    if(N1550) begin
      { valid[495:495] } <= { N1055 };
    end 
    if(N1549) begin
      { valid[494:494] } <= { N1055 };
    end 
    if(N1548) begin
      { valid[493:493] } <= { N1055 };
    end 
    if(N1547) begin
      { valid[492:492] } <= { N1055 };
    end 
    if(N1546) begin
      { valid[491:491] } <= { N1055 };
    end 
    if(N1545) begin
      { valid[490:490] } <= { N1055 };
    end 
    if(N1544) begin
      { valid[489:489] } <= { N1055 };
    end 
    if(N1543) begin
      { valid[488:488] } <= { N1055 };
    end 
    if(N1542) begin
      { valid[487:487] } <= { N1055 };
    end 
    if(N1541) begin
      { valid[486:486] } <= { N1055 };
    end 
    if(N1540) begin
      { valid[485:485] } <= { N1055 };
    end 
    if(N1539) begin
      { valid[484:484] } <= { N1055 };
    end 
    if(N1538) begin
      { valid[483:483] } <= { N1055 };
    end 
    if(N1537) begin
      { valid[482:482] } <= { N1055 };
    end 
    if(N1536) begin
      { valid[481:481] } <= { N1055 };
    end 
    if(N1535) begin
      { valid[480:480] } <= { N1055 };
    end 
    if(N1534) begin
      { valid[479:479] } <= { N1055 };
    end 
    if(N1533) begin
      { valid[478:478] } <= { N1055 };
    end 
    if(N1532) begin
      { valid[477:477] } <= { N1055 };
    end 
    if(N1531) begin
      { valid[476:476] } <= { N1055 };
    end 
    if(N1530) begin
      { valid[475:475] } <= { N1055 };
    end 
    if(N1529) begin
      { valid[474:474] } <= { N1055 };
    end 
    if(N1528) begin
      { valid[473:473] } <= { N1055 };
    end 
    if(N1527) begin
      { valid[472:472] } <= { N1055 };
    end 
    if(N1526) begin
      { valid[471:471] } <= { N1055 };
    end 
    if(N1525) begin
      { valid[470:470] } <= { N1055 };
    end 
    if(N1524) begin
      { valid[469:469] } <= { N1055 };
    end 
    if(N1523) begin
      { valid[468:468] } <= { N1055 };
    end 
    if(N1522) begin
      { valid[467:467] } <= { N1055 };
    end 
    if(N1521) begin
      { valid[466:466] } <= { N1055 };
    end 
    if(N1520) begin
      { valid[465:465] } <= { N1055 };
    end 
    if(N1519) begin
      { valid[464:464] } <= { N1055 };
    end 
    if(N1518) begin
      { valid[463:463] } <= { N1055 };
    end 
    if(N1517) begin
      { valid[462:462] } <= { N1055 };
    end 
    if(N1516) begin
      { valid[461:461] } <= { N1055 };
    end 
    if(N1515) begin
      { valid[460:460] } <= { N1055 };
    end 
    if(N1514) begin
      { valid[459:459] } <= { N1055 };
    end 
    if(N1513) begin
      { valid[458:458] } <= { N1055 };
    end 
    if(N1512) begin
      { valid[457:457] } <= { N1055 };
    end 
    if(N1511) begin
      { valid[456:456] } <= { N1055 };
    end 
    if(N1510) begin
      { valid[455:455] } <= { N1055 };
    end 
    if(N1509) begin
      { valid[454:454] } <= { N1055 };
    end 
    if(N1508) begin
      { valid[453:453] } <= { N1055 };
    end 
    if(N1507) begin
      { valid[452:452] } <= { N1055 };
    end 
    if(N1506) begin
      { valid[451:451] } <= { N1055 };
    end 
    if(N1505) begin
      { valid[450:450] } <= { N1055 };
    end 
    if(N1504) begin
      { valid[449:449] } <= { N1055 };
    end 
    if(N1503) begin
      { valid[448:448] } <= { N1055 };
    end 
    if(N1502) begin
      { valid[447:447] } <= { N1055 };
    end 
    if(N1501) begin
      { valid[446:446] } <= { N1055 };
    end 
    if(N1500) begin
      { valid[445:445] } <= { N1055 };
    end 
    if(N1499) begin
      { valid[444:444] } <= { N1055 };
    end 
    if(N1498) begin
      { valid[443:443] } <= { N1055 };
    end 
    if(N1497) begin
      { valid[442:442] } <= { N1055 };
    end 
    if(N1496) begin
      { valid[441:441] } <= { N1055 };
    end 
    if(N1495) begin
      { valid[440:440] } <= { N1055 };
    end 
    if(N1494) begin
      { valid[439:439] } <= { N1055 };
    end 
    if(N1493) begin
      { valid[438:438] } <= { N1055 };
    end 
    if(N1492) begin
      { valid[437:437] } <= { N1055 };
    end 
    if(N1491) begin
      { valid[436:436] } <= { N1055 };
    end 
    if(N1490) begin
      { valid[435:435] } <= { N1055 };
    end 
    if(N1489) begin
      { valid[434:434] } <= { N1055 };
    end 
    if(N1488) begin
      { valid[433:433] } <= { N1055 };
    end 
    if(N1487) begin
      { valid[432:432] } <= { N1055 };
    end 
    if(N1486) begin
      { valid[431:431] } <= { N1055 };
    end 
    if(N1485) begin
      { valid[430:430] } <= { N1055 };
    end 
    if(N1484) begin
      { valid[429:429] } <= { N1057 };
    end 
    if(N1483) begin
      { valid[428:428] } <= { N1057 };
    end 
    if(N1482) begin
      { valid[427:427] } <= { N1057 };
    end 
    if(N1481) begin
      { valid[426:426] } <= { N1057 };
    end 
    if(N1480) begin
      { valid[425:425] } <= { N1057 };
    end 
    if(N1479) begin
      { valid[424:424] } <= { N1057 };
    end 
    if(N1478) begin
      { valid[423:423] } <= { N1057 };
    end 
    if(N1477) begin
      { valid[422:422] } <= { N1057 };
    end 
    if(N1476) begin
      { valid[421:421] } <= { N1057 };
    end 
    if(N1475) begin
      { valid[420:420] } <= { N1057 };
    end 
    if(N1474) begin
      { valid[419:419] } <= { N1057 };
    end 
    if(N1473) begin
      { valid[418:418] } <= { N1057 };
    end 
    if(N1472) begin
      { valid[417:417] } <= { N1057 };
    end 
    if(N1471) begin
      { valid[416:416] } <= { N1057 };
    end 
    if(N1470) begin
      { valid[415:415] } <= { N1057 };
    end 
    if(N1469) begin
      { valid[414:414] } <= { N1057 };
    end 
    if(N1468) begin
      { valid[413:413] } <= { N1057 };
    end 
    if(N1467) begin
      { valid[412:412] } <= { N1057 };
    end 
    if(N1466) begin
      { valid[411:411] } <= { N1057 };
    end 
    if(N1465) begin
      { valid[410:410] } <= { N1057 };
    end 
    if(N1464) begin
      { valid[409:409] } <= { N1057 };
    end 
    if(N1463) begin
      { valid[408:408] } <= { N1057 };
    end 
    if(N1462) begin
      { valid[407:407] } <= { N1057 };
    end 
    if(N1461) begin
      { valid[406:406] } <= { N1057 };
    end 
    if(N1460) begin
      { valid[405:405] } <= { N1057 };
    end 
    if(N1459) begin
      { valid[404:404] } <= { N1057 };
    end 
    if(N1458) begin
      { valid[403:403] } <= { N1057 };
    end 
    if(N1457) begin
      { valid[402:402] } <= { N1057 };
    end 
    if(N1456) begin
      { valid[401:401] } <= { N1057 };
    end 
    if(N1455) begin
      { valid[400:400] } <= { N1057 };
    end 
    if(N1454) begin
      { valid[399:399] } <= { N1057 };
    end 
    if(N1453) begin
      { valid[398:398] } <= { N1057 };
    end 
    if(N1452) begin
      { valid[397:397] } <= { N1057 };
    end 
    if(N1451) begin
      { valid[396:396] } <= { N1057 };
    end 
    if(N1450) begin
      { valid[395:395] } <= { N1057 };
    end 
    if(N1449) begin
      { valid[394:394] } <= { N1057 };
    end 
    if(N1448) begin
      { valid[393:393] } <= { N1057 };
    end 
    if(N1447) begin
      { valid[392:392] } <= { N1057 };
    end 
    if(N1446) begin
      { valid[391:391] } <= { N1057 };
    end 
    if(N1445) begin
      { valid[390:390] } <= { N1057 };
    end 
    if(N1444) begin
      { valid[389:389] } <= { N1057 };
    end 
    if(N1443) begin
      { valid[388:388] } <= { N1057 };
    end 
    if(N1442) begin
      { valid[387:387] } <= { N1057 };
    end 
    if(N1441) begin
      { valid[386:386] } <= { N1057 };
    end 
    if(N1440) begin
      { valid[385:385] } <= { N1057 };
    end 
    if(N1439) begin
      { valid[384:384] } <= { N1057 };
    end 
    if(N1438) begin
      { valid[383:383] } <= { N1057 };
    end 
    if(N1437) begin
      { valid[382:382] } <= { N1057 };
    end 
    if(N1436) begin
      { valid[381:381] } <= { N1057 };
    end 
    if(N1435) begin
      { valid[380:380] } <= { N1057 };
    end 
    if(N1434) begin
      { valid[379:379] } <= { N1057 };
    end 
    if(N1433) begin
      { valid[378:378] } <= { N1057 };
    end 
    if(N1432) begin
      { valid[377:377] } <= { N1057 };
    end 
    if(N1431) begin
      { valid[376:376] } <= { N1057 };
    end 
    if(N1430) begin
      { valid[375:375] } <= { N1057 };
    end 
    if(N1429) begin
      { valid[374:374] } <= { N1057 };
    end 
    if(N1428) begin
      { valid[373:373] } <= { N1057 };
    end 
    if(N1427) begin
      { valid[372:372] } <= { N1057 };
    end 
    if(N1426) begin
      { valid[371:371] } <= { N1057 };
    end 
    if(N1425) begin
      { valid[370:370] } <= { N1057 };
    end 
    if(N1424) begin
      { valid[369:369] } <= { N1057 };
    end 
    if(N1423) begin
      { valid[368:368] } <= { N1057 };
    end 
    if(N1422) begin
      { valid[367:367] } <= { N1057 };
    end 
    if(N1421) begin
      { valid[366:366] } <= { N1057 };
    end 
    if(N1420) begin
      { valid[365:365] } <= { N1057 };
    end 
    if(N1419) begin
      { valid[364:364] } <= { N1057 };
    end 
    if(N1418) begin
      { valid[363:363] } <= { N1057 };
    end 
    if(N1417) begin
      { valid[362:362] } <= { N1057 };
    end 
    if(N1416) begin
      { valid[361:361] } <= { N1057 };
    end 
    if(N1415) begin
      { valid[360:360] } <= { N1057 };
    end 
    if(N1414) begin
      { valid[359:359] } <= { N1057 };
    end 
    if(N1413) begin
      { valid[358:358] } <= { N1057 };
    end 
    if(N1412) begin
      { valid[357:357] } <= { N1057 };
    end 
    if(N1411) begin
      { valid[356:356] } <= { N1057 };
    end 
    if(N1410) begin
      { valid[355:355] } <= { N1057 };
    end 
    if(N1409) begin
      { valid[354:354] } <= { N1057 };
    end 
    if(N1408) begin
      { valid[353:353] } <= { N1057 };
    end 
    if(N1407) begin
      { valid[352:352] } <= { N1057 };
    end 
    if(N1406) begin
      { valid[351:351] } <= { N1057 };
    end 
    if(N1405) begin
      { valid[350:350] } <= { N1057 };
    end 
    if(N1404) begin
      { valid[349:349] } <= { N1057 };
    end 
    if(N1403) begin
      { valid[348:348] } <= { N1057 };
    end 
    if(N1402) begin
      { valid[347:347] } <= { N1057 };
    end 
    if(N1401) begin
      { valid[346:346] } <= { N1057 };
    end 
    if(N1400) begin
      { valid[345:345] } <= { N1057 };
    end 
    if(N1399) begin
      { valid[344:344] } <= { N1057 };
    end 
    if(N1398) begin
      { valid[343:343] } <= { N1057 };
    end 
    if(N1397) begin
      { valid[342:342] } <= { N1057 };
    end 
    if(N1396) begin
      { valid[341:341] } <= { N1057 };
    end 
    if(N1395) begin
      { valid[340:340] } <= { N1057 };
    end 
    if(N1394) begin
      { valid[339:339] } <= { N1057 };
    end 
    if(N1393) begin
      { valid[338:338] } <= { N1057 };
    end 
    if(N1392) begin
      { valid[337:337] } <= { N1057 };
    end 
    if(N1391) begin
      { valid[336:336] } <= { N1057 };
    end 
    if(N1390) begin
      { valid[335:335] } <= { N1057 };
    end 
    if(N1389) begin
      { valid[334:334] } <= { N1057 };
    end 
    if(N1388) begin
      { valid[333:333] } <= { N1057 };
    end 
    if(N1387) begin
      { valid[332:332] } <= { N1057 };
    end 
    if(N1386) begin
      { valid[331:331] } <= { N1057 };
    end 
    if(N1385) begin
      { valid[330:330] } <= { N1059 };
    end 
    if(N1384) begin
      { valid[329:329] } <= { N1059 };
    end 
    if(N1383) begin
      { valid[328:328] } <= { N1059 };
    end 
    if(N1382) begin
      { valid[327:327] } <= { N1059 };
    end 
    if(N1381) begin
      { valid[326:326] } <= { N1059 };
    end 
    if(N1380) begin
      { valid[325:325] } <= { N1059 };
    end 
    if(N1379) begin
      { valid[324:324] } <= { N1059 };
    end 
    if(N1378) begin
      { valid[323:323] } <= { N1059 };
    end 
    if(N1377) begin
      { valid[322:322] } <= { N1059 };
    end 
    if(N1376) begin
      { valid[321:321] } <= { N1059 };
    end 
    if(N1375) begin
      { valid[320:320] } <= { N1059 };
    end 
    if(N1374) begin
      { valid[319:319] } <= { N1059 };
    end 
    if(N1373) begin
      { valid[318:318] } <= { N1059 };
    end 
    if(N1372) begin
      { valid[317:317] } <= { N1059 };
    end 
    if(N1371) begin
      { valid[316:316] } <= { N1059 };
    end 
    if(N1370) begin
      { valid[315:315] } <= { N1059 };
    end 
    if(N1369) begin
      { valid[314:314] } <= { N1059 };
    end 
    if(N1368) begin
      { valid[313:313] } <= { N1059 };
    end 
    if(N1367) begin
      { valid[312:312] } <= { N1059 };
    end 
    if(N1366) begin
      { valid[311:311] } <= { N1059 };
    end 
    if(N1365) begin
      { valid[310:310] } <= { N1059 };
    end 
    if(N1364) begin
      { valid[309:309] } <= { N1059 };
    end 
    if(N1363) begin
      { valid[308:308] } <= { N1059 };
    end 
    if(N1362) begin
      { valid[307:307] } <= { N1059 };
    end 
    if(N1361) begin
      { valid[306:306] } <= { N1059 };
    end 
    if(N1360) begin
      { valid[305:305] } <= { N1059 };
    end 
    if(N1359) begin
      { valid[304:304] } <= { N1059 };
    end 
    if(N1358) begin
      { valid[303:303] } <= { N1059 };
    end 
    if(N1357) begin
      { valid[302:302] } <= { N1059 };
    end 
    if(N1356) begin
      { valid[301:301] } <= { N1059 };
    end 
    if(N1355) begin
      { valid[300:300] } <= { N1059 };
    end 
    if(N1354) begin
      { valid[299:299] } <= { N1059 };
    end 
    if(N1353) begin
      { valid[298:298] } <= { N1059 };
    end 
    if(N1352) begin
      { valid[297:297] } <= { N1059 };
    end 
    if(N1351) begin
      { valid[296:296] } <= { N1059 };
    end 
    if(N1350) begin
      { valid[295:295] } <= { N1059 };
    end 
    if(N1349) begin
      { valid[294:294] } <= { N1059 };
    end 
    if(N1348) begin
      { valid[293:293] } <= { N1059 };
    end 
    if(N1347) begin
      { valid[292:292] } <= { N1059 };
    end 
    if(N1346) begin
      { valid[291:291] } <= { N1059 };
    end 
    if(N1345) begin
      { valid[290:290] } <= { N1059 };
    end 
    if(N1344) begin
      { valid[289:289] } <= { N1059 };
    end 
    if(N1343) begin
      { valid[288:288] } <= { N1059 };
    end 
    if(N1342) begin
      { valid[287:287] } <= { N1059 };
    end 
    if(N1341) begin
      { valid[286:286] } <= { N1059 };
    end 
    if(N1340) begin
      { valid[285:285] } <= { N1059 };
    end 
    if(N1339) begin
      { valid[284:284] } <= { N1059 };
    end 
    if(N1338) begin
      { valid[283:283] } <= { N1059 };
    end 
    if(N1337) begin
      { valid[282:282] } <= { N1059 };
    end 
    if(N1336) begin
      { valid[281:281] } <= { N1059 };
    end 
    if(N1335) begin
      { valid[280:280] } <= { N1059 };
    end 
    if(N1334) begin
      { valid[279:279] } <= { N1059 };
    end 
    if(N1333) begin
      { valid[278:278] } <= { N1059 };
    end 
    if(N1332) begin
      { valid[277:277] } <= { N1059 };
    end 
    if(N1331) begin
      { valid[276:276] } <= { N1059 };
    end 
    if(N1330) begin
      { valid[275:275] } <= { N1059 };
    end 
    if(N1329) begin
      { valid[274:274] } <= { N1059 };
    end 
    if(N1328) begin
      { valid[273:273] } <= { N1059 };
    end 
    if(N1327) begin
      { valid[272:272] } <= { N1059 };
    end 
    if(N1326) begin
      { valid[271:271] } <= { N1059 };
    end 
    if(N1325) begin
      { valid[270:270] } <= { N1059 };
    end 
    if(N1324) begin
      { valid[269:269] } <= { N1059 };
    end 
    if(N1323) begin
      { valid[268:268] } <= { N1059 };
    end 
    if(N1322) begin
      { valid[267:267] } <= { N1059 };
    end 
    if(N1321) begin
      { valid[266:266] } <= { N1059 };
    end 
    if(N1320) begin
      { valid[265:265] } <= { N1059 };
    end 
    if(N1319) begin
      { valid[264:264] } <= { N1059 };
    end 
    if(N1318) begin
      { valid[263:263] } <= { N1059 };
    end 
    if(N1317) begin
      { valid[262:262] } <= { N1059 };
    end 
    if(N1316) begin
      { valid[261:261] } <= { N1059 };
    end 
    if(N1315) begin
      { valid[260:260] } <= { N1059 };
    end 
    if(N1314) begin
      { valid[259:259] } <= { N1059 };
    end 
    if(N1313) begin
      { valid[258:258] } <= { N1059 };
    end 
    if(N1312) begin
      { valid[257:257] } <= { N1059 };
    end 
    if(N1311) begin
      { valid[256:256] } <= { N1059 };
    end 
    if(N1310) begin
      { valid[255:255] } <= { N1059 };
    end 
    if(N1309) begin
      { valid[254:254] } <= { N1059 };
    end 
    if(N1308) begin
      { valid[253:253] } <= { N1059 };
    end 
    if(N1307) begin
      { valid[252:252] } <= { N1059 };
    end 
    if(N1306) begin
      { valid[251:251] } <= { N1059 };
    end 
    if(N1305) begin
      { valid[250:250] } <= { N1059 };
    end 
    if(N1304) begin
      { valid[249:249] } <= { N1059 };
    end 
    if(N1303) begin
      { valid[248:248] } <= { N1059 };
    end 
    if(N1302) begin
      { valid[247:247] } <= { N1059 };
    end 
    if(N1301) begin
      { valid[246:246] } <= { N1059 };
    end 
    if(N1300) begin
      { valid[245:245] } <= { N1059 };
    end 
    if(N1299) begin
      { valid[244:244] } <= { N1059 };
    end 
    if(N1298) begin
      { valid[243:243] } <= { N1059 };
    end 
    if(N1297) begin
      { valid[242:242] } <= { N1059 };
    end 
    if(N1296) begin
      { valid[241:241] } <= { N1059 };
    end 
    if(N1295) begin
      { valid[240:240] } <= { N1059 };
    end 
    if(N1294) begin
      { valid[239:239] } <= { N1059 };
    end 
    if(N1293) begin
      { valid[238:238] } <= { N1059 };
    end 
    if(N1292) begin
      { valid[237:237] } <= { N1059 };
    end 
    if(N1291) begin
      { valid[236:236] } <= { N1059 };
    end 
    if(N1290) begin
      { valid[235:235] } <= { N1059 };
    end 
    if(N1289) begin
      { valid[234:234] } <= { N1059 };
    end 
    if(N1288) begin
      { valid[233:233] } <= { N1059 };
    end 
    if(N1287) begin
      { valid[232:232] } <= { N1059 };
    end 
    if(N1286) begin
      { valid[231:231] } <= { N1061 };
    end 
    if(N1285) begin
      { valid[230:230] } <= { N1061 };
    end 
    if(N1284) begin
      { valid[229:229] } <= { N1061 };
    end 
    if(N1283) begin
      { valid[228:228] } <= { N1061 };
    end 
    if(N1282) begin
      { valid[227:227] } <= { N1061 };
    end 
    if(N1281) begin
      { valid[226:226] } <= { N1061 };
    end 
    if(N1280) begin
      { valid[225:225] } <= { N1061 };
    end 
    if(N1279) begin
      { valid[224:224] } <= { N1061 };
    end 
    if(N1278) begin
      { valid[223:223] } <= { N1061 };
    end 
    if(N1277) begin
      { valid[222:222] } <= { N1061 };
    end 
    if(N1276) begin
      { valid[221:221] } <= { N1061 };
    end 
    if(N1275) begin
      { valid[220:220] } <= { N1061 };
    end 
    if(N1274) begin
      { valid[219:219] } <= { N1061 };
    end 
    if(N1273) begin
      { valid[218:218] } <= { N1061 };
    end 
    if(N1272) begin
      { valid[217:217] } <= { N1061 };
    end 
    if(N1271) begin
      { valid[216:216] } <= { N1061 };
    end 
    if(N1270) begin
      { valid[215:215] } <= { N1061 };
    end 
    if(N1269) begin
      { valid[214:214] } <= { N1061 };
    end 
    if(N1268) begin
      { valid[213:213] } <= { N1061 };
    end 
    if(N1267) begin
      { valid[212:212] } <= { N1061 };
    end 
    if(N1266) begin
      { valid[211:211] } <= { N1061 };
    end 
    if(N1265) begin
      { valid[210:210] } <= { N1061 };
    end 
    if(N1264) begin
      { valid[209:209] } <= { N1061 };
    end 
    if(N1263) begin
      { valid[208:208] } <= { N1061 };
    end 
    if(N1262) begin
      { valid[207:207] } <= { N1061 };
    end 
    if(N1261) begin
      { valid[206:206] } <= { N1061 };
    end 
    if(N1260) begin
      { valid[205:205] } <= { N1061 };
    end 
    if(N1259) begin
      { valid[204:204] } <= { N1061 };
    end 
    if(N1258) begin
      { valid[203:203] } <= { N1061 };
    end 
    if(N1257) begin
      { valid[202:202] } <= { N1061 };
    end 
    if(N1256) begin
      { valid[201:201] } <= { N1061 };
    end 
    if(N1255) begin
      { valid[200:200] } <= { N1061 };
    end 
    if(N1254) begin
      { valid[199:199] } <= { N1061 };
    end 
    if(N1253) begin
      { valid[198:198] } <= { N1061 };
    end 
    if(N1252) begin
      { valid[197:197] } <= { N1061 };
    end 
    if(N1251) begin
      { valid[196:196] } <= { N1061 };
    end 
    if(N1250) begin
      { valid[195:195] } <= { N1061 };
    end 
    if(N1249) begin
      { valid[194:194] } <= { N1061 };
    end 
    if(N1248) begin
      { valid[193:193] } <= { N1061 };
    end 
    if(N1247) begin
      { valid[192:192] } <= { N1061 };
    end 
    if(N1246) begin
      { valid[191:191] } <= { N1061 };
    end 
    if(N1245) begin
      { valid[190:190] } <= { N1061 };
    end 
    if(N1244) begin
      { valid[189:189] } <= { N1061 };
    end 
    if(N1243) begin
      { valid[188:188] } <= { N1061 };
    end 
    if(N1242) begin
      { valid[187:187] } <= { N1061 };
    end 
    if(N1241) begin
      { valid[186:186] } <= { N1061 };
    end 
    if(N1240) begin
      { valid[185:185] } <= { N1061 };
    end 
    if(N1239) begin
      { valid[184:184] } <= { N1061 };
    end 
    if(N1238) begin
      { valid[183:183] } <= { N1061 };
    end 
    if(N1237) begin
      { valid[182:182] } <= { N1061 };
    end 
    if(N1236) begin
      { valid[181:181] } <= { N1061 };
    end 
    if(N1235) begin
      { valid[180:180] } <= { N1061 };
    end 
    if(N1234) begin
      { valid[179:179] } <= { N1061 };
    end 
    if(N1233) begin
      { valid[178:178] } <= { N1061 };
    end 
    if(N1232) begin
      { valid[177:177] } <= { N1061 };
    end 
    if(N1231) begin
      { valid[176:176] } <= { N1061 };
    end 
    if(N1230) begin
      { valid[175:175] } <= { N1061 };
    end 
    if(N1229) begin
      { valid[174:174] } <= { N1061 };
    end 
    if(N1228) begin
      { valid[173:173] } <= { N1061 };
    end 
    if(N1227) begin
      { valid[172:172] } <= { N1061 };
    end 
    if(N1226) begin
      { valid[171:171] } <= { N1061 };
    end 
    if(N1225) begin
      { valid[170:170] } <= { N1061 };
    end 
    if(N1224) begin
      { valid[169:169] } <= { N1061 };
    end 
    if(N1223) begin
      { valid[168:168] } <= { N1061 };
    end 
    if(N1222) begin
      { valid[167:167] } <= { N1061 };
    end 
    if(N1221) begin
      { valid[166:166] } <= { N1061 };
    end 
    if(N1220) begin
      { valid[165:165] } <= { N1061 };
    end 
    if(N1219) begin
      { valid[164:164] } <= { N1061 };
    end 
    if(N1218) begin
      { valid[163:163] } <= { N1061 };
    end 
    if(N1217) begin
      { valid[162:162] } <= { N1061 };
    end 
    if(N1216) begin
      { valid[161:161] } <= { N1061 };
    end 
    if(N1215) begin
      { valid[160:160] } <= { N1061 };
    end 
    if(N1214) begin
      { valid[159:159] } <= { N1061 };
    end 
    if(N1213) begin
      { valid[158:158] } <= { N1061 };
    end 
    if(N1212) begin
      { valid[157:157] } <= { N1061 };
    end 
    if(N1211) begin
      { valid[156:156] } <= { N1061 };
    end 
    if(N1210) begin
      { valid[155:155] } <= { N1061 };
    end 
    if(N1209) begin
      { valid[154:154] } <= { N1061 };
    end 
    if(N1208) begin
      { valid[153:153] } <= { N1061 };
    end 
    if(N1207) begin
      { valid[152:152] } <= { N1061 };
    end 
    if(N1206) begin
      { valid[151:151] } <= { N1061 };
    end 
    if(N1205) begin
      { valid[150:150] } <= { N1061 };
    end 
    if(N1204) begin
      { valid[149:149] } <= { N1061 };
    end 
    if(N1203) begin
      { valid[148:148] } <= { N1061 };
    end 
    if(N1202) begin
      { valid[147:147] } <= { N1061 };
    end 
    if(N1201) begin
      { valid[146:146] } <= { N1061 };
    end 
    if(N1200) begin
      { valid[145:145] } <= { N1061 };
    end 
    if(N1199) begin
      { valid[144:144] } <= { N1061 };
    end 
    if(N1198) begin
      { valid[143:143] } <= { N1061 };
    end 
    if(N1197) begin
      { valid[142:142] } <= { N1061 };
    end 
    if(N1196) begin
      { valid[141:141] } <= { N1061 };
    end 
    if(N1195) begin
      { valid[140:140] } <= { N1061 };
    end 
    if(N1194) begin
      { valid[139:139] } <= { N1061 };
    end 
    if(N1193) begin
      { valid[138:138] } <= { N1061 };
    end 
    if(N1192) begin
      { valid[137:137] } <= { N1061 };
    end 
    if(N1191) begin
      { valid[136:136] } <= { N1061 };
    end 
    if(N1190) begin
      { valid[135:135] } <= { N1061 };
    end 
    if(N1189) begin
      { valid[134:134] } <= { N1061 };
    end 
    if(N1188) begin
      { valid[133:133] } <= { N1061 };
    end 
    if(N1187) begin
      { valid[132:132] } <= { N1063 };
    end 
    if(N1186) begin
      { valid[131:131] } <= { N1063 };
    end 
    if(N1185) begin
      { valid[130:130] } <= { N1063 };
    end 
    if(N1184) begin
      { valid[129:129] } <= { N1063 };
    end 
    if(N1183) begin
      { valid[128:128] } <= { N1063 };
    end 
    if(N1182) begin
      { valid[127:127] } <= { N1063 };
    end 
    if(N1181) begin
      { valid[126:126] } <= { N1063 };
    end 
    if(N1180) begin
      { valid[125:125] } <= { N1063 };
    end 
    if(N1179) begin
      { valid[124:124] } <= { N1063 };
    end 
    if(N1178) begin
      { valid[123:123] } <= { N1063 };
    end 
    if(N1177) begin
      { valid[122:122] } <= { N1063 };
    end 
    if(N1176) begin
      { valid[121:121] } <= { N1063 };
    end 
    if(N1175) begin
      { valid[120:120] } <= { N1063 };
    end 
    if(N1174) begin
      { valid[119:119] } <= { N1063 };
    end 
    if(N1173) begin
      { valid[118:118] } <= { N1063 };
    end 
    if(N1172) begin
      { valid[117:117] } <= { N1063 };
    end 
    if(N1171) begin
      { valid[116:116] } <= { N1063 };
    end 
    if(N1170) begin
      { valid[115:115] } <= { N1063 };
    end 
    if(N1169) begin
      { valid[114:114] } <= { N1063 };
    end 
    if(N1168) begin
      { valid[113:113] } <= { N1063 };
    end 
    if(N1167) begin
      { valid[112:112] } <= { N1063 };
    end 
    if(N1166) begin
      { valid[111:111] } <= { N1063 };
    end 
    if(N1165) begin
      { valid[110:110] } <= { N1063 };
    end 
    if(N1164) begin
      { valid[109:109] } <= { N1063 };
    end 
    if(N1163) begin
      { valid[108:108] } <= { N1063 };
    end 
    if(N1162) begin
      { valid[107:107] } <= { N1063 };
    end 
    if(N1161) begin
      { valid[106:106] } <= { N1063 };
    end 
    if(N1160) begin
      { valid[105:105] } <= { N1063 };
    end 
    if(N1159) begin
      { valid[104:104] } <= { N1063 };
    end 
    if(N1158) begin
      { valid[103:103] } <= { N1063 };
    end 
    if(N1157) begin
      { valid[102:102] } <= { N1063 };
    end 
    if(N1156) begin
      { valid[101:101] } <= { N1063 };
    end 
    if(N1155) begin
      { valid[100:100] } <= { N1063 };
    end 
    if(N1154) begin
      { valid[99:99] } <= { N1063 };
    end 
    if(N1153) begin
      { valid[98:98] } <= { N1063 };
    end 
    if(N1152) begin
      { valid[97:97] } <= { N1063 };
    end 
    if(N1151) begin
      { valid[96:96] } <= { N1063 };
    end 
    if(N1150) begin
      { valid[95:95] } <= { N1063 };
    end 
    if(N1149) begin
      { valid[94:94] } <= { N1063 };
    end 
    if(N1148) begin
      { valid[93:93] } <= { N1063 };
    end 
    if(N1147) begin
      { valid[92:92] } <= { N1063 };
    end 
    if(N1146) begin
      { valid[91:91] } <= { N1063 };
    end 
    if(N1145) begin
      { valid[90:90] } <= { N1063 };
    end 
    if(N1144) begin
      { valid[89:89] } <= { N1063 };
    end 
    if(N1143) begin
      { valid[88:88] } <= { N1063 };
    end 
    if(N1142) begin
      { valid[87:87] } <= { N1063 };
    end 
    if(N1141) begin
      { valid[86:86] } <= { N1063 };
    end 
    if(N1140) begin
      { valid[85:85] } <= { N1063 };
    end 
    if(N1139) begin
      { valid[84:84] } <= { N1063 };
    end 
    if(N1138) begin
      { valid[83:83] } <= { N1063 };
    end 
    if(N1137) begin
      { valid[82:82] } <= { N1063 };
    end 
    if(N1136) begin
      { valid[81:81] } <= { N1063 };
    end 
    if(N1135) begin
      { valid[80:80] } <= { N1063 };
    end 
    if(N1134) begin
      { valid[79:79] } <= { N1063 };
    end 
    if(N1133) begin
      { valid[78:78] } <= { N1063 };
    end 
    if(N1132) begin
      { valid[77:77] } <= { N1063 };
    end 
    if(N1131) begin
      { valid[76:76] } <= { N1063 };
    end 
    if(N1130) begin
      { valid[75:75] } <= { N1063 };
    end 
    if(N1129) begin
      { valid[74:74] } <= { N1063 };
    end 
    if(N1128) begin
      { valid[73:73] } <= { N1063 };
    end 
    if(N1127) begin
      { valid[72:72] } <= { N1063 };
    end 
    if(N1126) begin
      { valid[71:71] } <= { N1063 };
    end 
    if(N1125) begin
      { valid[70:70] } <= { N1063 };
    end 
    if(N1124) begin
      { valid[69:69] } <= { N1063 };
    end 
    if(N1123) begin
      { valid[68:68] } <= { N1063 };
    end 
    if(N1122) begin
      { valid[67:67] } <= { N1063 };
    end 
    if(N1121) begin
      { valid[66:66] } <= { N1063 };
    end 
    if(N1120) begin
      { valid[65:65] } <= { N1063 };
    end 
    if(N1119) begin
      { valid[64:64] } <= { N1063 };
    end 
    if(N1118) begin
      { valid[63:63] } <= { N1063 };
    end 
    if(N1117) begin
      { valid[62:62] } <= { N1063 };
    end 
    if(N1116) begin
      { valid[61:61] } <= { N1063 };
    end 
    if(N1115) begin
      { valid[60:60] } <= { N1063 };
    end 
    if(N1114) begin
      { valid[59:59] } <= { N1063 };
    end 
    if(N1113) begin
      { valid[58:58] } <= { N1063 };
    end 
    if(N1112) begin
      { valid[57:57] } <= { N1063 };
    end 
    if(N1111) begin
      { valid[56:56] } <= { N1063 };
    end 
    if(N1110) begin
      { valid[55:55] } <= { N1063 };
    end 
    if(N1109) begin
      { valid[54:54] } <= { N1063 };
    end 
    if(N1108) begin
      { valid[53:53] } <= { N1063 };
    end 
    if(N1107) begin
      { valid[52:52] } <= { N1063 };
    end 
    if(N1106) begin
      { valid[51:51] } <= { N1063 };
    end 
    if(N1105) begin
      { valid[50:50] } <= { N1063 };
    end 
    if(N1104) begin
      { valid[49:49] } <= { N1063 };
    end 
    if(N1103) begin
      { valid[48:48] } <= { N1063 };
    end 
    if(N1102) begin
      { valid[47:47] } <= { N1063 };
    end 
    if(N1101) begin
      { valid[46:46] } <= { N1063 };
    end 
    if(N1100) begin
      { valid[45:45] } <= { N1063 };
    end 
    if(N1099) begin
      { valid[44:44] } <= { N1063 };
    end 
    if(N1098) begin
      { valid[43:43] } <= { N1063 };
    end 
    if(N1097) begin
      { valid[42:42] } <= { N1063 };
    end 
    if(N1096) begin
      { valid[41:41] } <= { N1063 };
    end 
    if(N1095) begin
      { valid[40:40] } <= { N1063 };
    end 
    if(N1094) begin
      { valid[39:39] } <= { N1063 };
    end 
    if(N1093) begin
      { valid[38:38] } <= { N1063 };
    end 
    if(N1092) begin
      { valid[37:37] } <= { N1063 };
    end 
    if(N1091) begin
      { valid[36:36] } <= { N1063 };
    end 
    if(N1090) begin
      { valid[35:35] } <= { N1063 };
    end 
    if(N1089) begin
      { valid[34:34] } <= { N1063 };
    end 
    if(N1088) begin
      { valid[33:33] } <= { N1065 };
    end 
    if(N1087) begin
      { valid[32:32] } <= { N1065 };
    end 
    if(N1086) begin
      { valid[31:31] } <= { N1065 };
    end 
    if(N1085) begin
      { valid[30:30] } <= { N1065 };
    end 
    if(N1084) begin
      { valid[29:29] } <= { N1065 };
    end 
    if(N1083) begin
      { valid[28:28] } <= { N1065 };
    end 
    if(N1082) begin
      { valid[27:27] } <= { N1065 };
    end 
    if(N1081) begin
      { valid[26:26] } <= { N1065 };
    end 
    if(N1080) begin
      { valid[25:25] } <= { N1065 };
    end 
    if(N1079) begin
      { valid[24:24] } <= { N1065 };
    end 
    if(N1078) begin
      { valid[23:23] } <= { N1065 };
    end 
    if(N1077) begin
      { valid[22:22] } <= { N1065 };
    end 
    if(N1076) begin
      { valid[21:21] } <= { N1065 };
    end 
    if(N1075) begin
      { valid[20:20] } <= { N1065 };
    end 
    if(N1074) begin
      { valid[19:19] } <= { N1065 };
    end 
    if(N1073) begin
      { valid[18:18] } <= { N1065 };
    end 
    if(N1072) begin
      { valid[17:17] } <= { N1065 };
    end 
    if(N1071) begin
      { valid[16:16] } <= { N1065 };
    end 
    if(N1070) begin
      { valid[15:15] } <= { N1065 };
    end 
    if(N1069) begin
      { valid[14:14] } <= { N1065 };
    end 
    if(N1068) begin
      { valid[13:13] } <= { N1065 };
    end 
    if(N1067) begin
      { valid[12:12] } <= { N1065 };
    end 
    if(N1066) begin
      { valid[11:11] } <= { N1065 };
    end 
    if(N1064) begin
      { valid[10:10] } <= { N1065 };
    end 
    if(N1062) begin
      { valid[9:9] } <= { N1063 };
    end 
    if(N1060) begin
      { valid[8:8] } <= { N1061 };
    end 
    if(N1058) begin
      { valid[7:7] } <= { N1059 };
    end 
    if(N1056) begin
      { valid[6:6] } <= { N1057 };
    end 
    if(N1054) begin
      { valid[5:5] } <= { N1055 };
    end 
    if(N1052) begin
      { valid[4:4] } <= { N1053 };
    end 
    if(N1050) begin
      { valid[3:3] } <= { N1051 };
    end 
    if(N1048) begin
      { valid[2:2] } <= { N1049 };
    end 
    if(N1046) begin
      { valid[1:1] } <= { N1047 };
    end 
    if(N1044) begin
      { valid[0:0] } <= { N1045 };
    end 
  end


endmodule

