

module top
(
  data_i,
  sel_i,
  data_o
);

  input [1023:0] data_i;
  input [4:0] sel_i;
  output [1023:0] data_o;

  bsg_mux_butterfly
  wrapper
  (
    .data_i(data_i),
    .sel_i(sel_i),
    .data_o(data_o)
  );


endmodule



module bsg_swap_width_p32
(
  data_i,
  swap_i,
  data_o
);

  input [63:0] data_i;
  output [63:0] data_o;
  input swap_i;
  wire [63:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[31:0], data_i[63:32] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p64
(
  data_i,
  swap_i,
  data_o
);

  input [127:0] data_i;
  output [127:0] data_o;
  input swap_i;
  wire [127:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[63:0], data_i[127:64] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p128
(
  data_i,
  swap_i,
  data_o
);

  input [255:0] data_i;
  output [255:0] data_o;
  input swap_i;
  wire [255:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[127:0], data_i[255:128] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p256
(
  data_i,
  swap_i,
  data_o
);

  input [511:0] data_i;
  output [511:0] data_o;
  input swap_i;
  wire [511:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[255:0], data_i[511:256] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_swap_width_p512
(
  data_i,
  swap_i,
  data_o
);

  input [1023:0] data_i;
  output [1023:0] data_o;
  input swap_i;
  wire [1023:0] data_o;
  wire N0,N1,N2;
  assign data_o = (N0)? { data_i[511:0], data_i[1023:512] } : 
                  (N1)? data_i : 1'b0;
  assign N0 = swap_i;
  assign N1 = N2;
  assign N2 = ~swap_i;

endmodule



module bsg_mux_butterfly
(
  data_i,
  sel_i,
  data_o
);

  input [1023:0] data_i;
  input [4:0] sel_i;
  output [1023:0] data_o;
  wire [1023:0] data_o;
  wire data_stage_1__1023_,data_stage_1__1022_,data_stage_1__1021_,data_stage_1__1020_,
  data_stage_1__1019_,data_stage_1__1018_,data_stage_1__1017_,data_stage_1__1016_,
  data_stage_1__1015_,data_stage_1__1014_,data_stage_1__1013_,data_stage_1__1012_,
  data_stage_1__1011_,data_stage_1__1010_,data_stage_1__1009_,data_stage_1__1008_,
  data_stage_1__1007_,data_stage_1__1006_,data_stage_1__1005_,data_stage_1__1004_,
  data_stage_1__1003_,data_stage_1__1002_,data_stage_1__1001_,data_stage_1__1000_,
  data_stage_1__999_,data_stage_1__998_,data_stage_1__997_,data_stage_1__996_,
  data_stage_1__995_,data_stage_1__994_,data_stage_1__993_,data_stage_1__992_,
  data_stage_1__991_,data_stage_1__990_,data_stage_1__989_,data_stage_1__988_,
  data_stage_1__987_,data_stage_1__986_,data_stage_1__985_,data_stage_1__984_,
  data_stage_1__983_,data_stage_1__982_,data_stage_1__981_,data_stage_1__980_,data_stage_1__979_,
  data_stage_1__978_,data_stage_1__977_,data_stage_1__976_,data_stage_1__975_,
  data_stage_1__974_,data_stage_1__973_,data_stage_1__972_,data_stage_1__971_,
  data_stage_1__970_,data_stage_1__969_,data_stage_1__968_,data_stage_1__967_,
  data_stage_1__966_,data_stage_1__965_,data_stage_1__964_,data_stage_1__963_,
  data_stage_1__962_,data_stage_1__961_,data_stage_1__960_,data_stage_1__959_,data_stage_1__958_,
  data_stage_1__957_,data_stage_1__956_,data_stage_1__955_,data_stage_1__954_,
  data_stage_1__953_,data_stage_1__952_,data_stage_1__951_,data_stage_1__950_,
  data_stage_1__949_,data_stage_1__948_,data_stage_1__947_,data_stage_1__946_,
  data_stage_1__945_,data_stage_1__944_,data_stage_1__943_,data_stage_1__942_,
  data_stage_1__941_,data_stage_1__940_,data_stage_1__939_,data_stage_1__938_,data_stage_1__937_,
  data_stage_1__936_,data_stage_1__935_,data_stage_1__934_,data_stage_1__933_,
  data_stage_1__932_,data_stage_1__931_,data_stage_1__930_,data_stage_1__929_,
  data_stage_1__928_,data_stage_1__927_,data_stage_1__926_,data_stage_1__925_,
  data_stage_1__924_,data_stage_1__923_,data_stage_1__922_,data_stage_1__921_,data_stage_1__920_,
  data_stage_1__919_,data_stage_1__918_,data_stage_1__917_,data_stage_1__916_,
  data_stage_1__915_,data_stage_1__914_,data_stage_1__913_,data_stage_1__912_,
  data_stage_1__911_,data_stage_1__910_,data_stage_1__909_,data_stage_1__908_,
  data_stage_1__907_,data_stage_1__906_,data_stage_1__905_,data_stage_1__904_,
  data_stage_1__903_,data_stage_1__902_,data_stage_1__901_,data_stage_1__900_,data_stage_1__899_,
  data_stage_1__898_,data_stage_1__897_,data_stage_1__896_,data_stage_1__895_,
  data_stage_1__894_,data_stage_1__893_,data_stage_1__892_,data_stage_1__891_,
  data_stage_1__890_,data_stage_1__889_,data_stage_1__888_,data_stage_1__887_,
  data_stage_1__886_,data_stage_1__885_,data_stage_1__884_,data_stage_1__883_,
  data_stage_1__882_,data_stage_1__881_,data_stage_1__880_,data_stage_1__879_,data_stage_1__878_,
  data_stage_1__877_,data_stage_1__876_,data_stage_1__875_,data_stage_1__874_,
  data_stage_1__873_,data_stage_1__872_,data_stage_1__871_,data_stage_1__870_,
  data_stage_1__869_,data_stage_1__868_,data_stage_1__867_,data_stage_1__866_,
  data_stage_1__865_,data_stage_1__864_,data_stage_1__863_,data_stage_1__862_,
  data_stage_1__861_,data_stage_1__860_,data_stage_1__859_,data_stage_1__858_,data_stage_1__857_,
  data_stage_1__856_,data_stage_1__855_,data_stage_1__854_,data_stage_1__853_,
  data_stage_1__852_,data_stage_1__851_,data_stage_1__850_,data_stage_1__849_,
  data_stage_1__848_,data_stage_1__847_,data_stage_1__846_,data_stage_1__845_,
  data_stage_1__844_,data_stage_1__843_,data_stage_1__842_,data_stage_1__841_,data_stage_1__840_,
  data_stage_1__839_,data_stage_1__838_,data_stage_1__837_,data_stage_1__836_,
  data_stage_1__835_,data_stage_1__834_,data_stage_1__833_,data_stage_1__832_,
  data_stage_1__831_,data_stage_1__830_,data_stage_1__829_,data_stage_1__828_,
  data_stage_1__827_,data_stage_1__826_,data_stage_1__825_,data_stage_1__824_,
  data_stage_1__823_,data_stage_1__822_,data_stage_1__821_,data_stage_1__820_,data_stage_1__819_,
  data_stage_1__818_,data_stage_1__817_,data_stage_1__816_,data_stage_1__815_,
  data_stage_1__814_,data_stage_1__813_,data_stage_1__812_,data_stage_1__811_,
  data_stage_1__810_,data_stage_1__809_,data_stage_1__808_,data_stage_1__807_,
  data_stage_1__806_,data_stage_1__805_,data_stage_1__804_,data_stage_1__803_,
  data_stage_1__802_,data_stage_1__801_,data_stage_1__800_,data_stage_1__799_,data_stage_1__798_,
  data_stage_1__797_,data_stage_1__796_,data_stage_1__795_,data_stage_1__794_,
  data_stage_1__793_,data_stage_1__792_,data_stage_1__791_,data_stage_1__790_,
  data_stage_1__789_,data_stage_1__788_,data_stage_1__787_,data_stage_1__786_,
  data_stage_1__785_,data_stage_1__784_,data_stage_1__783_,data_stage_1__782_,
  data_stage_1__781_,data_stage_1__780_,data_stage_1__779_,data_stage_1__778_,data_stage_1__777_,
  data_stage_1__776_,data_stage_1__775_,data_stage_1__774_,data_stage_1__773_,
  data_stage_1__772_,data_stage_1__771_,data_stage_1__770_,data_stage_1__769_,
  data_stage_1__768_,data_stage_1__767_,data_stage_1__766_,data_stage_1__765_,
  data_stage_1__764_,data_stage_1__763_,data_stage_1__762_,data_stage_1__761_,data_stage_1__760_,
  data_stage_1__759_,data_stage_1__758_,data_stage_1__757_,data_stage_1__756_,
  data_stage_1__755_,data_stage_1__754_,data_stage_1__753_,data_stage_1__752_,
  data_stage_1__751_,data_stage_1__750_,data_stage_1__749_,data_stage_1__748_,
  data_stage_1__747_,data_stage_1__746_,data_stage_1__745_,data_stage_1__744_,
  data_stage_1__743_,data_stage_1__742_,data_stage_1__741_,data_stage_1__740_,data_stage_1__739_,
  data_stage_1__738_,data_stage_1__737_,data_stage_1__736_,data_stage_1__735_,
  data_stage_1__734_,data_stage_1__733_,data_stage_1__732_,data_stage_1__731_,
  data_stage_1__730_,data_stage_1__729_,data_stage_1__728_,data_stage_1__727_,
  data_stage_1__726_,data_stage_1__725_,data_stage_1__724_,data_stage_1__723_,
  data_stage_1__722_,data_stage_1__721_,data_stage_1__720_,data_stage_1__719_,data_stage_1__718_,
  data_stage_1__717_,data_stage_1__716_,data_stage_1__715_,data_stage_1__714_,
  data_stage_1__713_,data_stage_1__712_,data_stage_1__711_,data_stage_1__710_,
  data_stage_1__709_,data_stage_1__708_,data_stage_1__707_,data_stage_1__706_,
  data_stage_1__705_,data_stage_1__704_,data_stage_1__703_,data_stage_1__702_,
  data_stage_1__701_,data_stage_1__700_,data_stage_1__699_,data_stage_1__698_,data_stage_1__697_,
  data_stage_1__696_,data_stage_1__695_,data_stage_1__694_,data_stage_1__693_,
  data_stage_1__692_,data_stage_1__691_,data_stage_1__690_,data_stage_1__689_,
  data_stage_1__688_,data_stage_1__687_,data_stage_1__686_,data_stage_1__685_,
  data_stage_1__684_,data_stage_1__683_,data_stage_1__682_,data_stage_1__681_,data_stage_1__680_,
  data_stage_1__679_,data_stage_1__678_,data_stage_1__677_,data_stage_1__676_,
  data_stage_1__675_,data_stage_1__674_,data_stage_1__673_,data_stage_1__672_,
  data_stage_1__671_,data_stage_1__670_,data_stage_1__669_,data_stage_1__668_,
  data_stage_1__667_,data_stage_1__666_,data_stage_1__665_,data_stage_1__664_,
  data_stage_1__663_,data_stage_1__662_,data_stage_1__661_,data_stage_1__660_,data_stage_1__659_,
  data_stage_1__658_,data_stage_1__657_,data_stage_1__656_,data_stage_1__655_,
  data_stage_1__654_,data_stage_1__653_,data_stage_1__652_,data_stage_1__651_,
  data_stage_1__650_,data_stage_1__649_,data_stage_1__648_,data_stage_1__647_,
  data_stage_1__646_,data_stage_1__645_,data_stage_1__644_,data_stage_1__643_,
  data_stage_1__642_,data_stage_1__641_,data_stage_1__640_,data_stage_1__639_,data_stage_1__638_,
  data_stage_1__637_,data_stage_1__636_,data_stage_1__635_,data_stage_1__634_,
  data_stage_1__633_,data_stage_1__632_,data_stage_1__631_,data_stage_1__630_,
  data_stage_1__629_,data_stage_1__628_,data_stage_1__627_,data_stage_1__626_,
  data_stage_1__625_,data_stage_1__624_,data_stage_1__623_,data_stage_1__622_,
  data_stage_1__621_,data_stage_1__620_,data_stage_1__619_,data_stage_1__618_,data_stage_1__617_,
  data_stage_1__616_,data_stage_1__615_,data_stage_1__614_,data_stage_1__613_,
  data_stage_1__612_,data_stage_1__611_,data_stage_1__610_,data_stage_1__609_,
  data_stage_1__608_,data_stage_1__607_,data_stage_1__606_,data_stage_1__605_,
  data_stage_1__604_,data_stage_1__603_,data_stage_1__602_,data_stage_1__601_,data_stage_1__600_,
  data_stage_1__599_,data_stage_1__598_,data_stage_1__597_,data_stage_1__596_,
  data_stage_1__595_,data_stage_1__594_,data_stage_1__593_,data_stage_1__592_,
  data_stage_1__591_,data_stage_1__590_,data_stage_1__589_,data_stage_1__588_,
  data_stage_1__587_,data_stage_1__586_,data_stage_1__585_,data_stage_1__584_,
  data_stage_1__583_,data_stage_1__582_,data_stage_1__581_,data_stage_1__580_,data_stage_1__579_,
  data_stage_1__578_,data_stage_1__577_,data_stage_1__576_,data_stage_1__575_,
  data_stage_1__574_,data_stage_1__573_,data_stage_1__572_,data_stage_1__571_,
  data_stage_1__570_,data_stage_1__569_,data_stage_1__568_,data_stage_1__567_,
  data_stage_1__566_,data_stage_1__565_,data_stage_1__564_,data_stage_1__563_,
  data_stage_1__562_,data_stage_1__561_,data_stage_1__560_,data_stage_1__559_,data_stage_1__558_,
  data_stage_1__557_,data_stage_1__556_,data_stage_1__555_,data_stage_1__554_,
  data_stage_1__553_,data_stage_1__552_,data_stage_1__551_,data_stage_1__550_,
  data_stage_1__549_,data_stage_1__548_,data_stage_1__547_,data_stage_1__546_,
  data_stage_1__545_,data_stage_1__544_,data_stage_1__543_,data_stage_1__542_,
  data_stage_1__541_,data_stage_1__540_,data_stage_1__539_,data_stage_1__538_,data_stage_1__537_,
  data_stage_1__536_,data_stage_1__535_,data_stage_1__534_,data_stage_1__533_,
  data_stage_1__532_,data_stage_1__531_,data_stage_1__530_,data_stage_1__529_,
  data_stage_1__528_,data_stage_1__527_,data_stage_1__526_,data_stage_1__525_,
  data_stage_1__524_,data_stage_1__523_,data_stage_1__522_,data_stage_1__521_,data_stage_1__520_,
  data_stage_1__519_,data_stage_1__518_,data_stage_1__517_,data_stage_1__516_,
  data_stage_1__515_,data_stage_1__514_,data_stage_1__513_,data_stage_1__512_,
  data_stage_1__511_,data_stage_1__510_,data_stage_1__509_,data_stage_1__508_,
  data_stage_1__507_,data_stage_1__506_,data_stage_1__505_,data_stage_1__504_,
  data_stage_1__503_,data_stage_1__502_,data_stage_1__501_,data_stage_1__500_,data_stage_1__499_,
  data_stage_1__498_,data_stage_1__497_,data_stage_1__496_,data_stage_1__495_,
  data_stage_1__494_,data_stage_1__493_,data_stage_1__492_,data_stage_1__491_,
  data_stage_1__490_,data_stage_1__489_,data_stage_1__488_,data_stage_1__487_,
  data_stage_1__486_,data_stage_1__485_,data_stage_1__484_,data_stage_1__483_,
  data_stage_1__482_,data_stage_1__481_,data_stage_1__480_,data_stage_1__479_,data_stage_1__478_,
  data_stage_1__477_,data_stage_1__476_,data_stage_1__475_,data_stage_1__474_,
  data_stage_1__473_,data_stage_1__472_,data_stage_1__471_,data_stage_1__470_,
  data_stage_1__469_,data_stage_1__468_,data_stage_1__467_,data_stage_1__466_,
  data_stage_1__465_,data_stage_1__464_,data_stage_1__463_,data_stage_1__462_,
  data_stage_1__461_,data_stage_1__460_,data_stage_1__459_,data_stage_1__458_,data_stage_1__457_,
  data_stage_1__456_,data_stage_1__455_,data_stage_1__454_,data_stage_1__453_,
  data_stage_1__452_,data_stage_1__451_,data_stage_1__450_,data_stage_1__449_,
  data_stage_1__448_,data_stage_1__447_,data_stage_1__446_,data_stage_1__445_,
  data_stage_1__444_,data_stage_1__443_,data_stage_1__442_,data_stage_1__441_,data_stage_1__440_,
  data_stage_1__439_,data_stage_1__438_,data_stage_1__437_,data_stage_1__436_,
  data_stage_1__435_,data_stage_1__434_,data_stage_1__433_,data_stage_1__432_,
  data_stage_1__431_,data_stage_1__430_,data_stage_1__429_,data_stage_1__428_,
  data_stage_1__427_,data_stage_1__426_,data_stage_1__425_,data_stage_1__424_,
  data_stage_1__423_,data_stage_1__422_,data_stage_1__421_,data_stage_1__420_,data_stage_1__419_,
  data_stage_1__418_,data_stage_1__417_,data_stage_1__416_,data_stage_1__415_,
  data_stage_1__414_,data_stage_1__413_,data_stage_1__412_,data_stage_1__411_,
  data_stage_1__410_,data_stage_1__409_,data_stage_1__408_,data_stage_1__407_,
  data_stage_1__406_,data_stage_1__405_,data_stage_1__404_,data_stage_1__403_,
  data_stage_1__402_,data_stage_1__401_,data_stage_1__400_,data_stage_1__399_,data_stage_1__398_,
  data_stage_1__397_,data_stage_1__396_,data_stage_1__395_,data_stage_1__394_,
  data_stage_1__393_,data_stage_1__392_,data_stage_1__391_,data_stage_1__390_,
  data_stage_1__389_,data_stage_1__388_,data_stage_1__387_,data_stage_1__386_,
  data_stage_1__385_,data_stage_1__384_,data_stage_1__383_,data_stage_1__382_,
  data_stage_1__381_,data_stage_1__380_,data_stage_1__379_,data_stage_1__378_,data_stage_1__377_,
  data_stage_1__376_,data_stage_1__375_,data_stage_1__374_,data_stage_1__373_,
  data_stage_1__372_,data_stage_1__371_,data_stage_1__370_,data_stage_1__369_,
  data_stage_1__368_,data_stage_1__367_,data_stage_1__366_,data_stage_1__365_,
  data_stage_1__364_,data_stage_1__363_,data_stage_1__362_,data_stage_1__361_,data_stage_1__360_,
  data_stage_1__359_,data_stage_1__358_,data_stage_1__357_,data_stage_1__356_,
  data_stage_1__355_,data_stage_1__354_,data_stage_1__353_,data_stage_1__352_,
  data_stage_1__351_,data_stage_1__350_,data_stage_1__349_,data_stage_1__348_,
  data_stage_1__347_,data_stage_1__346_,data_stage_1__345_,data_stage_1__344_,
  data_stage_1__343_,data_stage_1__342_,data_stage_1__341_,data_stage_1__340_,data_stage_1__339_,
  data_stage_1__338_,data_stage_1__337_,data_stage_1__336_,data_stage_1__335_,
  data_stage_1__334_,data_stage_1__333_,data_stage_1__332_,data_stage_1__331_,
  data_stage_1__330_,data_stage_1__329_,data_stage_1__328_,data_stage_1__327_,
  data_stage_1__326_,data_stage_1__325_,data_stage_1__324_,data_stage_1__323_,
  data_stage_1__322_,data_stage_1__321_,data_stage_1__320_,data_stage_1__319_,data_stage_1__318_,
  data_stage_1__317_,data_stage_1__316_,data_stage_1__315_,data_stage_1__314_,
  data_stage_1__313_,data_stage_1__312_,data_stage_1__311_,data_stage_1__310_,
  data_stage_1__309_,data_stage_1__308_,data_stage_1__307_,data_stage_1__306_,
  data_stage_1__305_,data_stage_1__304_,data_stage_1__303_,data_stage_1__302_,
  data_stage_1__301_,data_stage_1__300_,data_stage_1__299_,data_stage_1__298_,data_stage_1__297_,
  data_stage_1__296_,data_stage_1__295_,data_stage_1__294_,data_stage_1__293_,
  data_stage_1__292_,data_stage_1__291_,data_stage_1__290_,data_stage_1__289_,
  data_stage_1__288_,data_stage_1__287_,data_stage_1__286_,data_stage_1__285_,
  data_stage_1__284_,data_stage_1__283_,data_stage_1__282_,data_stage_1__281_,data_stage_1__280_,
  data_stage_1__279_,data_stage_1__278_,data_stage_1__277_,data_stage_1__276_,
  data_stage_1__275_,data_stage_1__274_,data_stage_1__273_,data_stage_1__272_,
  data_stage_1__271_,data_stage_1__270_,data_stage_1__269_,data_stage_1__268_,
  data_stage_1__267_,data_stage_1__266_,data_stage_1__265_,data_stage_1__264_,
  data_stage_1__263_,data_stage_1__262_,data_stage_1__261_,data_stage_1__260_,data_stage_1__259_,
  data_stage_1__258_,data_stage_1__257_,data_stage_1__256_,data_stage_1__255_,
  data_stage_1__254_,data_stage_1__253_,data_stage_1__252_,data_stage_1__251_,
  data_stage_1__250_,data_stage_1__249_,data_stage_1__248_,data_stage_1__247_,
  data_stage_1__246_,data_stage_1__245_,data_stage_1__244_,data_stage_1__243_,
  data_stage_1__242_,data_stage_1__241_,data_stage_1__240_,data_stage_1__239_,data_stage_1__238_,
  data_stage_1__237_,data_stage_1__236_,data_stage_1__235_,data_stage_1__234_,
  data_stage_1__233_,data_stage_1__232_,data_stage_1__231_,data_stage_1__230_,
  data_stage_1__229_,data_stage_1__228_,data_stage_1__227_,data_stage_1__226_,
  data_stage_1__225_,data_stage_1__224_,data_stage_1__223_,data_stage_1__222_,
  data_stage_1__221_,data_stage_1__220_,data_stage_1__219_,data_stage_1__218_,data_stage_1__217_,
  data_stage_1__216_,data_stage_1__215_,data_stage_1__214_,data_stage_1__213_,
  data_stage_1__212_,data_stage_1__211_,data_stage_1__210_,data_stage_1__209_,
  data_stage_1__208_,data_stage_1__207_,data_stage_1__206_,data_stage_1__205_,
  data_stage_1__204_,data_stage_1__203_,data_stage_1__202_,data_stage_1__201_,data_stage_1__200_,
  data_stage_1__199_,data_stage_1__198_,data_stage_1__197_,data_stage_1__196_,
  data_stage_1__195_,data_stage_1__194_,data_stage_1__193_,data_stage_1__192_,
  data_stage_1__191_,data_stage_1__190_,data_stage_1__189_,data_stage_1__188_,
  data_stage_1__187_,data_stage_1__186_,data_stage_1__185_,data_stage_1__184_,
  data_stage_1__183_,data_stage_1__182_,data_stage_1__181_,data_stage_1__180_,data_stage_1__179_,
  data_stage_1__178_,data_stage_1__177_,data_stage_1__176_,data_stage_1__175_,
  data_stage_1__174_,data_stage_1__173_,data_stage_1__172_,data_stage_1__171_,
  data_stage_1__170_,data_stage_1__169_,data_stage_1__168_,data_stage_1__167_,
  data_stage_1__166_,data_stage_1__165_,data_stage_1__164_,data_stage_1__163_,
  data_stage_1__162_,data_stage_1__161_,data_stage_1__160_,data_stage_1__159_,data_stage_1__158_,
  data_stage_1__157_,data_stage_1__156_,data_stage_1__155_,data_stage_1__154_,
  data_stage_1__153_,data_stage_1__152_,data_stage_1__151_,data_stage_1__150_,
  data_stage_1__149_,data_stage_1__148_,data_stage_1__147_,data_stage_1__146_,
  data_stage_1__145_,data_stage_1__144_,data_stage_1__143_,data_stage_1__142_,
  data_stage_1__141_,data_stage_1__140_,data_stage_1__139_,data_stage_1__138_,data_stage_1__137_,
  data_stage_1__136_,data_stage_1__135_,data_stage_1__134_,data_stage_1__133_,
  data_stage_1__132_,data_stage_1__131_,data_stage_1__130_,data_stage_1__129_,
  data_stage_1__128_,data_stage_1__127_,data_stage_1__126_,data_stage_1__125_,
  data_stage_1__124_,data_stage_1__123_,data_stage_1__122_,data_stage_1__121_,data_stage_1__120_,
  data_stage_1__119_,data_stage_1__118_,data_stage_1__117_,data_stage_1__116_,
  data_stage_1__115_,data_stage_1__114_,data_stage_1__113_,data_stage_1__112_,
  data_stage_1__111_,data_stage_1__110_,data_stage_1__109_,data_stage_1__108_,
  data_stage_1__107_,data_stage_1__106_,data_stage_1__105_,data_stage_1__104_,
  data_stage_1__103_,data_stage_1__102_,data_stage_1__101_,data_stage_1__100_,data_stage_1__99_,
  data_stage_1__98_,data_stage_1__97_,data_stage_1__96_,data_stage_1__95_,
  data_stage_1__94_,data_stage_1__93_,data_stage_1__92_,data_stage_1__91_,data_stage_1__90_,
  data_stage_1__89_,data_stage_1__88_,data_stage_1__87_,data_stage_1__86_,
  data_stage_1__85_,data_stage_1__84_,data_stage_1__83_,data_stage_1__82_,
  data_stage_1__81_,data_stage_1__80_,data_stage_1__79_,data_stage_1__78_,data_stage_1__77_,
  data_stage_1__76_,data_stage_1__75_,data_stage_1__74_,data_stage_1__73_,
  data_stage_1__72_,data_stage_1__71_,data_stage_1__70_,data_stage_1__69_,data_stage_1__68_,
  data_stage_1__67_,data_stage_1__66_,data_stage_1__65_,data_stage_1__64_,
  data_stage_1__63_,data_stage_1__62_,data_stage_1__61_,data_stage_1__60_,data_stage_1__59_,
  data_stage_1__58_,data_stage_1__57_,data_stage_1__56_,data_stage_1__55_,
  data_stage_1__54_,data_stage_1__53_,data_stage_1__52_,data_stage_1__51_,data_stage_1__50_,
  data_stage_1__49_,data_stage_1__48_,data_stage_1__47_,data_stage_1__46_,
  data_stage_1__45_,data_stage_1__44_,data_stage_1__43_,data_stage_1__42_,
  data_stage_1__41_,data_stage_1__40_,data_stage_1__39_,data_stage_1__38_,data_stage_1__37_,
  data_stage_1__36_,data_stage_1__35_,data_stage_1__34_,data_stage_1__33_,
  data_stage_1__32_,data_stage_1__31_,data_stage_1__30_,data_stage_1__29_,data_stage_1__28_,
  data_stage_1__27_,data_stage_1__26_,data_stage_1__25_,data_stage_1__24_,
  data_stage_1__23_,data_stage_1__22_,data_stage_1__21_,data_stage_1__20_,data_stage_1__19_,
  data_stage_1__18_,data_stage_1__17_,data_stage_1__16_,data_stage_1__15_,
  data_stage_1__14_,data_stage_1__13_,data_stage_1__12_,data_stage_1__11_,data_stage_1__10_,
  data_stage_1__9_,data_stage_1__8_,data_stage_1__7_,data_stage_1__6_,
  data_stage_1__5_,data_stage_1__4_,data_stage_1__3_,data_stage_1__2_,data_stage_1__1_,
  data_stage_1__0_,data_stage_2__1023_,data_stage_2__1022_,data_stage_2__1021_,
  data_stage_2__1020_,data_stage_2__1019_,data_stage_2__1018_,data_stage_2__1017_,
  data_stage_2__1016_,data_stage_2__1015_,data_stage_2__1014_,data_stage_2__1013_,
  data_stage_2__1012_,data_stage_2__1011_,data_stage_2__1010_,data_stage_2__1009_,
  data_stage_2__1008_,data_stage_2__1007_,data_stage_2__1006_,data_stage_2__1005_,
  data_stage_2__1004_,data_stage_2__1003_,data_stage_2__1002_,data_stage_2__1001_,
  data_stage_2__1000_,data_stage_2__999_,data_stage_2__998_,data_stage_2__997_,
  data_stage_2__996_,data_stage_2__995_,data_stage_2__994_,data_stage_2__993_,
  data_stage_2__992_,data_stage_2__991_,data_stage_2__990_,data_stage_2__989_,data_stage_2__988_,
  data_stage_2__987_,data_stage_2__986_,data_stage_2__985_,data_stage_2__984_,
  data_stage_2__983_,data_stage_2__982_,data_stage_2__981_,data_stage_2__980_,
  data_stage_2__979_,data_stage_2__978_,data_stage_2__977_,data_stage_2__976_,
  data_stage_2__975_,data_stage_2__974_,data_stage_2__973_,data_stage_2__972_,
  data_stage_2__971_,data_stage_2__970_,data_stage_2__969_,data_stage_2__968_,data_stage_2__967_,
  data_stage_2__966_,data_stage_2__965_,data_stage_2__964_,data_stage_2__963_,
  data_stage_2__962_,data_stage_2__961_,data_stage_2__960_,data_stage_2__959_,
  data_stage_2__958_,data_stage_2__957_,data_stage_2__956_,data_stage_2__955_,
  data_stage_2__954_,data_stage_2__953_,data_stage_2__952_,data_stage_2__951_,data_stage_2__950_,
  data_stage_2__949_,data_stage_2__948_,data_stage_2__947_,data_stage_2__946_,
  data_stage_2__945_,data_stage_2__944_,data_stage_2__943_,data_stage_2__942_,
  data_stage_2__941_,data_stage_2__940_,data_stage_2__939_,data_stage_2__938_,
  data_stage_2__937_,data_stage_2__936_,data_stage_2__935_,data_stage_2__934_,
  data_stage_2__933_,data_stage_2__932_,data_stage_2__931_,data_stage_2__930_,data_stage_2__929_,
  data_stage_2__928_,data_stage_2__927_,data_stage_2__926_,data_stage_2__925_,
  data_stage_2__924_,data_stage_2__923_,data_stage_2__922_,data_stage_2__921_,
  data_stage_2__920_,data_stage_2__919_,data_stage_2__918_,data_stage_2__917_,
  data_stage_2__916_,data_stage_2__915_,data_stage_2__914_,data_stage_2__913_,
  data_stage_2__912_,data_stage_2__911_,data_stage_2__910_,data_stage_2__909_,data_stage_2__908_,
  data_stage_2__907_,data_stage_2__906_,data_stage_2__905_,data_stage_2__904_,
  data_stage_2__903_,data_stage_2__902_,data_stage_2__901_,data_stage_2__900_,
  data_stage_2__899_,data_stage_2__898_,data_stage_2__897_,data_stage_2__896_,
  data_stage_2__895_,data_stage_2__894_,data_stage_2__893_,data_stage_2__892_,
  data_stage_2__891_,data_stage_2__890_,data_stage_2__889_,data_stage_2__888_,data_stage_2__887_,
  data_stage_2__886_,data_stage_2__885_,data_stage_2__884_,data_stage_2__883_,
  data_stage_2__882_,data_stage_2__881_,data_stage_2__880_,data_stage_2__879_,
  data_stage_2__878_,data_stage_2__877_,data_stage_2__876_,data_stage_2__875_,
  data_stage_2__874_,data_stage_2__873_,data_stage_2__872_,data_stage_2__871_,data_stage_2__870_,
  data_stage_2__869_,data_stage_2__868_,data_stage_2__867_,data_stage_2__866_,
  data_stage_2__865_,data_stage_2__864_,data_stage_2__863_,data_stage_2__862_,
  data_stage_2__861_,data_stage_2__860_,data_stage_2__859_,data_stage_2__858_,
  data_stage_2__857_,data_stage_2__856_,data_stage_2__855_,data_stage_2__854_,
  data_stage_2__853_,data_stage_2__852_,data_stage_2__851_,data_stage_2__850_,data_stage_2__849_,
  data_stage_2__848_,data_stage_2__847_,data_stage_2__846_,data_stage_2__845_,
  data_stage_2__844_,data_stage_2__843_,data_stage_2__842_,data_stage_2__841_,
  data_stage_2__840_,data_stage_2__839_,data_stage_2__838_,data_stage_2__837_,
  data_stage_2__836_,data_stage_2__835_,data_stage_2__834_,data_stage_2__833_,
  data_stage_2__832_,data_stage_2__831_,data_stage_2__830_,data_stage_2__829_,data_stage_2__828_,
  data_stage_2__827_,data_stage_2__826_,data_stage_2__825_,data_stage_2__824_,
  data_stage_2__823_,data_stage_2__822_,data_stage_2__821_,data_stage_2__820_,
  data_stage_2__819_,data_stage_2__818_,data_stage_2__817_,data_stage_2__816_,
  data_stage_2__815_,data_stage_2__814_,data_stage_2__813_,data_stage_2__812_,
  data_stage_2__811_,data_stage_2__810_,data_stage_2__809_,data_stage_2__808_,data_stage_2__807_,
  data_stage_2__806_,data_stage_2__805_,data_stage_2__804_,data_stage_2__803_,
  data_stage_2__802_,data_stage_2__801_,data_stage_2__800_,data_stage_2__799_,
  data_stage_2__798_,data_stage_2__797_,data_stage_2__796_,data_stage_2__795_,
  data_stage_2__794_,data_stage_2__793_,data_stage_2__792_,data_stage_2__791_,data_stage_2__790_,
  data_stage_2__789_,data_stage_2__788_,data_stage_2__787_,data_stage_2__786_,
  data_stage_2__785_,data_stage_2__784_,data_stage_2__783_,data_stage_2__782_,
  data_stage_2__781_,data_stage_2__780_,data_stage_2__779_,data_stage_2__778_,
  data_stage_2__777_,data_stage_2__776_,data_stage_2__775_,data_stage_2__774_,
  data_stage_2__773_,data_stage_2__772_,data_stage_2__771_,data_stage_2__770_,data_stage_2__769_,
  data_stage_2__768_,data_stage_2__767_,data_stage_2__766_,data_stage_2__765_,
  data_stage_2__764_,data_stage_2__763_,data_stage_2__762_,data_stage_2__761_,
  data_stage_2__760_,data_stage_2__759_,data_stage_2__758_,data_stage_2__757_,
  data_stage_2__756_,data_stage_2__755_,data_stage_2__754_,data_stage_2__753_,
  data_stage_2__752_,data_stage_2__751_,data_stage_2__750_,data_stage_2__749_,data_stage_2__748_,
  data_stage_2__747_,data_stage_2__746_,data_stage_2__745_,data_stage_2__744_,
  data_stage_2__743_,data_stage_2__742_,data_stage_2__741_,data_stage_2__740_,
  data_stage_2__739_,data_stage_2__738_,data_stage_2__737_,data_stage_2__736_,
  data_stage_2__735_,data_stage_2__734_,data_stage_2__733_,data_stage_2__732_,
  data_stage_2__731_,data_stage_2__730_,data_stage_2__729_,data_stage_2__728_,data_stage_2__727_,
  data_stage_2__726_,data_stage_2__725_,data_stage_2__724_,data_stage_2__723_,
  data_stage_2__722_,data_stage_2__721_,data_stage_2__720_,data_stage_2__719_,
  data_stage_2__718_,data_stage_2__717_,data_stage_2__716_,data_stage_2__715_,
  data_stage_2__714_,data_stage_2__713_,data_stage_2__712_,data_stage_2__711_,data_stage_2__710_,
  data_stage_2__709_,data_stage_2__708_,data_stage_2__707_,data_stage_2__706_,
  data_stage_2__705_,data_stage_2__704_,data_stage_2__703_,data_stage_2__702_,
  data_stage_2__701_,data_stage_2__700_,data_stage_2__699_,data_stage_2__698_,
  data_stage_2__697_,data_stage_2__696_,data_stage_2__695_,data_stage_2__694_,
  data_stage_2__693_,data_stage_2__692_,data_stage_2__691_,data_stage_2__690_,data_stage_2__689_,
  data_stage_2__688_,data_stage_2__687_,data_stage_2__686_,data_stage_2__685_,
  data_stage_2__684_,data_stage_2__683_,data_stage_2__682_,data_stage_2__681_,
  data_stage_2__680_,data_stage_2__679_,data_stage_2__678_,data_stage_2__677_,
  data_stage_2__676_,data_stage_2__675_,data_stage_2__674_,data_stage_2__673_,
  data_stage_2__672_,data_stage_2__671_,data_stage_2__670_,data_stage_2__669_,data_stage_2__668_,
  data_stage_2__667_,data_stage_2__666_,data_stage_2__665_,data_stage_2__664_,
  data_stage_2__663_,data_stage_2__662_,data_stage_2__661_,data_stage_2__660_,
  data_stage_2__659_,data_stage_2__658_,data_stage_2__657_,data_stage_2__656_,
  data_stage_2__655_,data_stage_2__654_,data_stage_2__653_,data_stage_2__652_,
  data_stage_2__651_,data_stage_2__650_,data_stage_2__649_,data_stage_2__648_,data_stage_2__647_,
  data_stage_2__646_,data_stage_2__645_,data_stage_2__644_,data_stage_2__643_,
  data_stage_2__642_,data_stage_2__641_,data_stage_2__640_,data_stage_2__639_,
  data_stage_2__638_,data_stage_2__637_,data_stage_2__636_,data_stage_2__635_,
  data_stage_2__634_,data_stage_2__633_,data_stage_2__632_,data_stage_2__631_,data_stage_2__630_,
  data_stage_2__629_,data_stage_2__628_,data_stage_2__627_,data_stage_2__626_,
  data_stage_2__625_,data_stage_2__624_,data_stage_2__623_,data_stage_2__622_,
  data_stage_2__621_,data_stage_2__620_,data_stage_2__619_,data_stage_2__618_,
  data_stage_2__617_,data_stage_2__616_,data_stage_2__615_,data_stage_2__614_,
  data_stage_2__613_,data_stage_2__612_,data_stage_2__611_,data_stage_2__610_,data_stage_2__609_,
  data_stage_2__608_,data_stage_2__607_,data_stage_2__606_,data_stage_2__605_,
  data_stage_2__604_,data_stage_2__603_,data_stage_2__602_,data_stage_2__601_,
  data_stage_2__600_,data_stage_2__599_,data_stage_2__598_,data_stage_2__597_,
  data_stage_2__596_,data_stage_2__595_,data_stage_2__594_,data_stage_2__593_,
  data_stage_2__592_,data_stage_2__591_,data_stage_2__590_,data_stage_2__589_,data_stage_2__588_,
  data_stage_2__587_,data_stage_2__586_,data_stage_2__585_,data_stage_2__584_,
  data_stage_2__583_,data_stage_2__582_,data_stage_2__581_,data_stage_2__580_,
  data_stage_2__579_,data_stage_2__578_,data_stage_2__577_,data_stage_2__576_,
  data_stage_2__575_,data_stage_2__574_,data_stage_2__573_,data_stage_2__572_,
  data_stage_2__571_,data_stage_2__570_,data_stage_2__569_,data_stage_2__568_,data_stage_2__567_,
  data_stage_2__566_,data_stage_2__565_,data_stage_2__564_,data_stage_2__563_,
  data_stage_2__562_,data_stage_2__561_,data_stage_2__560_,data_stage_2__559_,
  data_stage_2__558_,data_stage_2__557_,data_stage_2__556_,data_stage_2__555_,
  data_stage_2__554_,data_stage_2__553_,data_stage_2__552_,data_stage_2__551_,data_stage_2__550_,
  data_stage_2__549_,data_stage_2__548_,data_stage_2__547_,data_stage_2__546_,
  data_stage_2__545_,data_stage_2__544_,data_stage_2__543_,data_stage_2__542_,
  data_stage_2__541_,data_stage_2__540_,data_stage_2__539_,data_stage_2__538_,
  data_stage_2__537_,data_stage_2__536_,data_stage_2__535_,data_stage_2__534_,
  data_stage_2__533_,data_stage_2__532_,data_stage_2__531_,data_stage_2__530_,data_stage_2__529_,
  data_stage_2__528_,data_stage_2__527_,data_stage_2__526_,data_stage_2__525_,
  data_stage_2__524_,data_stage_2__523_,data_stage_2__522_,data_stage_2__521_,
  data_stage_2__520_,data_stage_2__519_,data_stage_2__518_,data_stage_2__517_,
  data_stage_2__516_,data_stage_2__515_,data_stage_2__514_,data_stage_2__513_,
  data_stage_2__512_,data_stage_2__511_,data_stage_2__510_,data_stage_2__509_,data_stage_2__508_,
  data_stage_2__507_,data_stage_2__506_,data_stage_2__505_,data_stage_2__504_,
  data_stage_2__503_,data_stage_2__502_,data_stage_2__501_,data_stage_2__500_,
  data_stage_2__499_,data_stage_2__498_,data_stage_2__497_,data_stage_2__496_,
  data_stage_2__495_,data_stage_2__494_,data_stage_2__493_,data_stage_2__492_,
  data_stage_2__491_,data_stage_2__490_,data_stage_2__489_,data_stage_2__488_,data_stage_2__487_,
  data_stage_2__486_,data_stage_2__485_,data_stage_2__484_,data_stage_2__483_,
  data_stage_2__482_,data_stage_2__481_,data_stage_2__480_,data_stage_2__479_,
  data_stage_2__478_,data_stage_2__477_,data_stage_2__476_,data_stage_2__475_,
  data_stage_2__474_,data_stage_2__473_,data_stage_2__472_,data_stage_2__471_,data_stage_2__470_,
  data_stage_2__469_,data_stage_2__468_,data_stage_2__467_,data_stage_2__466_,
  data_stage_2__465_,data_stage_2__464_,data_stage_2__463_,data_stage_2__462_,
  data_stage_2__461_,data_stage_2__460_,data_stage_2__459_,data_stage_2__458_,
  data_stage_2__457_,data_stage_2__456_,data_stage_2__455_,data_stage_2__454_,
  data_stage_2__453_,data_stage_2__452_,data_stage_2__451_,data_stage_2__450_,data_stage_2__449_,
  data_stage_2__448_,data_stage_2__447_,data_stage_2__446_,data_stage_2__445_,
  data_stage_2__444_,data_stage_2__443_,data_stage_2__442_,data_stage_2__441_,
  data_stage_2__440_,data_stage_2__439_,data_stage_2__438_,data_stage_2__437_,
  data_stage_2__436_,data_stage_2__435_,data_stage_2__434_,data_stage_2__433_,
  data_stage_2__432_,data_stage_2__431_,data_stage_2__430_,data_stage_2__429_,data_stage_2__428_,
  data_stage_2__427_,data_stage_2__426_,data_stage_2__425_,data_stage_2__424_,
  data_stage_2__423_,data_stage_2__422_,data_stage_2__421_,data_stage_2__420_,
  data_stage_2__419_,data_stage_2__418_,data_stage_2__417_,data_stage_2__416_,
  data_stage_2__415_,data_stage_2__414_,data_stage_2__413_,data_stage_2__412_,
  data_stage_2__411_,data_stage_2__410_,data_stage_2__409_,data_stage_2__408_,data_stage_2__407_,
  data_stage_2__406_,data_stage_2__405_,data_stage_2__404_,data_stage_2__403_,
  data_stage_2__402_,data_stage_2__401_,data_stage_2__400_,data_stage_2__399_,
  data_stage_2__398_,data_stage_2__397_,data_stage_2__396_,data_stage_2__395_,
  data_stage_2__394_,data_stage_2__393_,data_stage_2__392_,data_stage_2__391_,data_stage_2__390_,
  data_stage_2__389_,data_stage_2__388_,data_stage_2__387_,data_stage_2__386_,
  data_stage_2__385_,data_stage_2__384_,data_stage_2__383_,data_stage_2__382_,
  data_stage_2__381_,data_stage_2__380_,data_stage_2__379_,data_stage_2__378_,
  data_stage_2__377_,data_stage_2__376_,data_stage_2__375_,data_stage_2__374_,
  data_stage_2__373_,data_stage_2__372_,data_stage_2__371_,data_stage_2__370_,data_stage_2__369_,
  data_stage_2__368_,data_stage_2__367_,data_stage_2__366_,data_stage_2__365_,
  data_stage_2__364_,data_stage_2__363_,data_stage_2__362_,data_stage_2__361_,
  data_stage_2__360_,data_stage_2__359_,data_stage_2__358_,data_stage_2__357_,
  data_stage_2__356_,data_stage_2__355_,data_stage_2__354_,data_stage_2__353_,
  data_stage_2__352_,data_stage_2__351_,data_stage_2__350_,data_stage_2__349_,data_stage_2__348_,
  data_stage_2__347_,data_stage_2__346_,data_stage_2__345_,data_stage_2__344_,
  data_stage_2__343_,data_stage_2__342_,data_stage_2__341_,data_stage_2__340_,
  data_stage_2__339_,data_stage_2__338_,data_stage_2__337_,data_stage_2__336_,
  data_stage_2__335_,data_stage_2__334_,data_stage_2__333_,data_stage_2__332_,
  data_stage_2__331_,data_stage_2__330_,data_stage_2__329_,data_stage_2__328_,data_stage_2__327_,
  data_stage_2__326_,data_stage_2__325_,data_stage_2__324_,data_stage_2__323_,
  data_stage_2__322_,data_stage_2__321_,data_stage_2__320_,data_stage_2__319_,
  data_stage_2__318_,data_stage_2__317_,data_stage_2__316_,data_stage_2__315_,
  data_stage_2__314_,data_stage_2__313_,data_stage_2__312_,data_stage_2__311_,data_stage_2__310_,
  data_stage_2__309_,data_stage_2__308_,data_stage_2__307_,data_stage_2__306_,
  data_stage_2__305_,data_stage_2__304_,data_stage_2__303_,data_stage_2__302_,
  data_stage_2__301_,data_stage_2__300_,data_stage_2__299_,data_stage_2__298_,
  data_stage_2__297_,data_stage_2__296_,data_stage_2__295_,data_stage_2__294_,
  data_stage_2__293_,data_stage_2__292_,data_stage_2__291_,data_stage_2__290_,data_stage_2__289_,
  data_stage_2__288_,data_stage_2__287_,data_stage_2__286_,data_stage_2__285_,
  data_stage_2__284_,data_stage_2__283_,data_stage_2__282_,data_stage_2__281_,
  data_stage_2__280_,data_stage_2__279_,data_stage_2__278_,data_stage_2__277_,
  data_stage_2__276_,data_stage_2__275_,data_stage_2__274_,data_stage_2__273_,
  data_stage_2__272_,data_stage_2__271_,data_stage_2__270_,data_stage_2__269_,data_stage_2__268_,
  data_stage_2__267_,data_stage_2__266_,data_stage_2__265_,data_stage_2__264_,
  data_stage_2__263_,data_stage_2__262_,data_stage_2__261_,data_stage_2__260_,
  data_stage_2__259_,data_stage_2__258_,data_stage_2__257_,data_stage_2__256_,
  data_stage_2__255_,data_stage_2__254_,data_stage_2__253_,data_stage_2__252_,
  data_stage_2__251_,data_stage_2__250_,data_stage_2__249_,data_stage_2__248_,data_stage_2__247_,
  data_stage_2__246_,data_stage_2__245_,data_stage_2__244_,data_stage_2__243_,
  data_stage_2__242_,data_stage_2__241_,data_stage_2__240_,data_stage_2__239_,
  data_stage_2__238_,data_stage_2__237_,data_stage_2__236_,data_stage_2__235_,
  data_stage_2__234_,data_stage_2__233_,data_stage_2__232_,data_stage_2__231_,data_stage_2__230_,
  data_stage_2__229_,data_stage_2__228_,data_stage_2__227_,data_stage_2__226_,
  data_stage_2__225_,data_stage_2__224_,data_stage_2__223_,data_stage_2__222_,
  data_stage_2__221_,data_stage_2__220_,data_stage_2__219_,data_stage_2__218_,
  data_stage_2__217_,data_stage_2__216_,data_stage_2__215_,data_stage_2__214_,
  data_stage_2__213_,data_stage_2__212_,data_stage_2__211_,data_stage_2__210_,data_stage_2__209_,
  data_stage_2__208_,data_stage_2__207_,data_stage_2__206_,data_stage_2__205_,
  data_stage_2__204_,data_stage_2__203_,data_stage_2__202_,data_stage_2__201_,
  data_stage_2__200_,data_stage_2__199_,data_stage_2__198_,data_stage_2__197_,
  data_stage_2__196_,data_stage_2__195_,data_stage_2__194_,data_stage_2__193_,
  data_stage_2__192_,data_stage_2__191_,data_stage_2__190_,data_stage_2__189_,data_stage_2__188_,
  data_stage_2__187_,data_stage_2__186_,data_stage_2__185_,data_stage_2__184_,
  data_stage_2__183_,data_stage_2__182_,data_stage_2__181_,data_stage_2__180_,
  data_stage_2__179_,data_stage_2__178_,data_stage_2__177_,data_stage_2__176_,
  data_stage_2__175_,data_stage_2__174_,data_stage_2__173_,data_stage_2__172_,
  data_stage_2__171_,data_stage_2__170_,data_stage_2__169_,data_stage_2__168_,data_stage_2__167_,
  data_stage_2__166_,data_stage_2__165_,data_stage_2__164_,data_stage_2__163_,
  data_stage_2__162_,data_stage_2__161_,data_stage_2__160_,data_stage_2__159_,
  data_stage_2__158_,data_stage_2__157_,data_stage_2__156_,data_stage_2__155_,
  data_stage_2__154_,data_stage_2__153_,data_stage_2__152_,data_stage_2__151_,data_stage_2__150_,
  data_stage_2__149_,data_stage_2__148_,data_stage_2__147_,data_stage_2__146_,
  data_stage_2__145_,data_stage_2__144_,data_stage_2__143_,data_stage_2__142_,
  data_stage_2__141_,data_stage_2__140_,data_stage_2__139_,data_stage_2__138_,
  data_stage_2__137_,data_stage_2__136_,data_stage_2__135_,data_stage_2__134_,
  data_stage_2__133_,data_stage_2__132_,data_stage_2__131_,data_stage_2__130_,data_stage_2__129_,
  data_stage_2__128_,data_stage_2__127_,data_stage_2__126_,data_stage_2__125_,
  data_stage_2__124_,data_stage_2__123_,data_stage_2__122_,data_stage_2__121_,
  data_stage_2__120_,data_stage_2__119_,data_stage_2__118_,data_stage_2__117_,
  data_stage_2__116_,data_stage_2__115_,data_stage_2__114_,data_stage_2__113_,
  data_stage_2__112_,data_stage_2__111_,data_stage_2__110_,data_stage_2__109_,data_stage_2__108_,
  data_stage_2__107_,data_stage_2__106_,data_stage_2__105_,data_stage_2__104_,
  data_stage_2__103_,data_stage_2__102_,data_stage_2__101_,data_stage_2__100_,
  data_stage_2__99_,data_stage_2__98_,data_stage_2__97_,data_stage_2__96_,data_stage_2__95_,
  data_stage_2__94_,data_stage_2__93_,data_stage_2__92_,data_stage_2__91_,
  data_stage_2__90_,data_stage_2__89_,data_stage_2__88_,data_stage_2__87_,
  data_stage_2__86_,data_stage_2__85_,data_stage_2__84_,data_stage_2__83_,data_stage_2__82_,
  data_stage_2__81_,data_stage_2__80_,data_stage_2__79_,data_stage_2__78_,
  data_stage_2__77_,data_stage_2__76_,data_stage_2__75_,data_stage_2__74_,data_stage_2__73_,
  data_stage_2__72_,data_stage_2__71_,data_stage_2__70_,data_stage_2__69_,
  data_stage_2__68_,data_stage_2__67_,data_stage_2__66_,data_stage_2__65_,data_stage_2__64_,
  data_stage_2__63_,data_stage_2__62_,data_stage_2__61_,data_stage_2__60_,
  data_stage_2__59_,data_stage_2__58_,data_stage_2__57_,data_stage_2__56_,data_stage_2__55_,
  data_stage_2__54_,data_stage_2__53_,data_stage_2__52_,data_stage_2__51_,
  data_stage_2__50_,data_stage_2__49_,data_stage_2__48_,data_stage_2__47_,
  data_stage_2__46_,data_stage_2__45_,data_stage_2__44_,data_stage_2__43_,data_stage_2__42_,
  data_stage_2__41_,data_stage_2__40_,data_stage_2__39_,data_stage_2__38_,
  data_stage_2__37_,data_stage_2__36_,data_stage_2__35_,data_stage_2__34_,data_stage_2__33_,
  data_stage_2__32_,data_stage_2__31_,data_stage_2__30_,data_stage_2__29_,
  data_stage_2__28_,data_stage_2__27_,data_stage_2__26_,data_stage_2__25_,data_stage_2__24_,
  data_stage_2__23_,data_stage_2__22_,data_stage_2__21_,data_stage_2__20_,
  data_stage_2__19_,data_stage_2__18_,data_stage_2__17_,data_stage_2__16_,data_stage_2__15_,
  data_stage_2__14_,data_stage_2__13_,data_stage_2__12_,data_stage_2__11_,
  data_stage_2__10_,data_stage_2__9_,data_stage_2__8_,data_stage_2__7_,data_stage_2__6_,
  data_stage_2__5_,data_stage_2__4_,data_stage_2__3_,data_stage_2__2_,
  data_stage_2__1_,data_stage_2__0_,data_stage_3__1023_,data_stage_3__1022_,data_stage_3__1021_,
  data_stage_3__1020_,data_stage_3__1019_,data_stage_3__1018_,data_stage_3__1017_,
  data_stage_3__1016_,data_stage_3__1015_,data_stage_3__1014_,data_stage_3__1013_,
  data_stage_3__1012_,data_stage_3__1011_,data_stage_3__1010_,data_stage_3__1009_,
  data_stage_3__1008_,data_stage_3__1007_,data_stage_3__1006_,data_stage_3__1005_,
  data_stage_3__1004_,data_stage_3__1003_,data_stage_3__1002_,data_stage_3__1001_,
  data_stage_3__1000_,data_stage_3__999_,data_stage_3__998_,data_stage_3__997_,
  data_stage_3__996_,data_stage_3__995_,data_stage_3__994_,data_stage_3__993_,
  data_stage_3__992_,data_stage_3__991_,data_stage_3__990_,data_stage_3__989_,
  data_stage_3__988_,data_stage_3__987_,data_stage_3__986_,data_stage_3__985_,
  data_stage_3__984_,data_stage_3__983_,data_stage_3__982_,data_stage_3__981_,data_stage_3__980_,
  data_stage_3__979_,data_stage_3__978_,data_stage_3__977_,data_stage_3__976_,
  data_stage_3__975_,data_stage_3__974_,data_stage_3__973_,data_stage_3__972_,
  data_stage_3__971_,data_stage_3__970_,data_stage_3__969_,data_stage_3__968_,
  data_stage_3__967_,data_stage_3__966_,data_stage_3__965_,data_stage_3__964_,
  data_stage_3__963_,data_stage_3__962_,data_stage_3__961_,data_stage_3__960_,data_stage_3__959_,
  data_stage_3__958_,data_stage_3__957_,data_stage_3__956_,data_stage_3__955_,
  data_stage_3__954_,data_stage_3__953_,data_stage_3__952_,data_stage_3__951_,
  data_stage_3__950_,data_stage_3__949_,data_stage_3__948_,data_stage_3__947_,
  data_stage_3__946_,data_stage_3__945_,data_stage_3__944_,data_stage_3__943_,
  data_stage_3__942_,data_stage_3__941_,data_stage_3__940_,data_stage_3__939_,data_stage_3__938_,
  data_stage_3__937_,data_stage_3__936_,data_stage_3__935_,data_stage_3__934_,
  data_stage_3__933_,data_stage_3__932_,data_stage_3__931_,data_stage_3__930_,
  data_stage_3__929_,data_stage_3__928_,data_stage_3__927_,data_stage_3__926_,
  data_stage_3__925_,data_stage_3__924_,data_stage_3__923_,data_stage_3__922_,
  data_stage_3__921_,data_stage_3__920_,data_stage_3__919_,data_stage_3__918_,data_stage_3__917_,
  data_stage_3__916_,data_stage_3__915_,data_stage_3__914_,data_stage_3__913_,
  data_stage_3__912_,data_stage_3__911_,data_stage_3__910_,data_stage_3__909_,
  data_stage_3__908_,data_stage_3__907_,data_stage_3__906_,data_stage_3__905_,
  data_stage_3__904_,data_stage_3__903_,data_stage_3__902_,data_stage_3__901_,data_stage_3__900_,
  data_stage_3__899_,data_stage_3__898_,data_stage_3__897_,data_stage_3__896_,
  data_stage_3__895_,data_stage_3__894_,data_stage_3__893_,data_stage_3__892_,
  data_stage_3__891_,data_stage_3__890_,data_stage_3__889_,data_stage_3__888_,
  data_stage_3__887_,data_stage_3__886_,data_stage_3__885_,data_stage_3__884_,
  data_stage_3__883_,data_stage_3__882_,data_stage_3__881_,data_stage_3__880_,data_stage_3__879_,
  data_stage_3__878_,data_stage_3__877_,data_stage_3__876_,data_stage_3__875_,
  data_stage_3__874_,data_stage_3__873_,data_stage_3__872_,data_stage_3__871_,
  data_stage_3__870_,data_stage_3__869_,data_stage_3__868_,data_stage_3__867_,
  data_stage_3__866_,data_stage_3__865_,data_stage_3__864_,data_stage_3__863_,
  data_stage_3__862_,data_stage_3__861_,data_stage_3__860_,data_stage_3__859_,data_stage_3__858_,
  data_stage_3__857_,data_stage_3__856_,data_stage_3__855_,data_stage_3__854_,
  data_stage_3__853_,data_stage_3__852_,data_stage_3__851_,data_stage_3__850_,
  data_stage_3__849_,data_stage_3__848_,data_stage_3__847_,data_stage_3__846_,
  data_stage_3__845_,data_stage_3__844_,data_stage_3__843_,data_stage_3__842_,
  data_stage_3__841_,data_stage_3__840_,data_stage_3__839_,data_stage_3__838_,data_stage_3__837_,
  data_stage_3__836_,data_stage_3__835_,data_stage_3__834_,data_stage_3__833_,
  data_stage_3__832_,data_stage_3__831_,data_stage_3__830_,data_stage_3__829_,
  data_stage_3__828_,data_stage_3__827_,data_stage_3__826_,data_stage_3__825_,
  data_stage_3__824_,data_stage_3__823_,data_stage_3__822_,data_stage_3__821_,data_stage_3__820_,
  data_stage_3__819_,data_stage_3__818_,data_stage_3__817_,data_stage_3__816_,
  data_stage_3__815_,data_stage_3__814_,data_stage_3__813_,data_stage_3__812_,
  data_stage_3__811_,data_stage_3__810_,data_stage_3__809_,data_stage_3__808_,
  data_stage_3__807_,data_stage_3__806_,data_stage_3__805_,data_stage_3__804_,
  data_stage_3__803_,data_stage_3__802_,data_stage_3__801_,data_stage_3__800_,data_stage_3__799_,
  data_stage_3__798_,data_stage_3__797_,data_stage_3__796_,data_stage_3__795_,
  data_stage_3__794_,data_stage_3__793_,data_stage_3__792_,data_stage_3__791_,
  data_stage_3__790_,data_stage_3__789_,data_stage_3__788_,data_stage_3__787_,
  data_stage_3__786_,data_stage_3__785_,data_stage_3__784_,data_stage_3__783_,
  data_stage_3__782_,data_stage_3__781_,data_stage_3__780_,data_stage_3__779_,data_stage_3__778_,
  data_stage_3__777_,data_stage_3__776_,data_stage_3__775_,data_stage_3__774_,
  data_stage_3__773_,data_stage_3__772_,data_stage_3__771_,data_stage_3__770_,
  data_stage_3__769_,data_stage_3__768_,data_stage_3__767_,data_stage_3__766_,
  data_stage_3__765_,data_stage_3__764_,data_stage_3__763_,data_stage_3__762_,
  data_stage_3__761_,data_stage_3__760_,data_stage_3__759_,data_stage_3__758_,data_stage_3__757_,
  data_stage_3__756_,data_stage_3__755_,data_stage_3__754_,data_stage_3__753_,
  data_stage_3__752_,data_stage_3__751_,data_stage_3__750_,data_stage_3__749_,
  data_stage_3__748_,data_stage_3__747_,data_stage_3__746_,data_stage_3__745_,
  data_stage_3__744_,data_stage_3__743_,data_stage_3__742_,data_stage_3__741_,data_stage_3__740_,
  data_stage_3__739_,data_stage_3__738_,data_stage_3__737_,data_stage_3__736_,
  data_stage_3__735_,data_stage_3__734_,data_stage_3__733_,data_stage_3__732_,
  data_stage_3__731_,data_stage_3__730_,data_stage_3__729_,data_stage_3__728_,
  data_stage_3__727_,data_stage_3__726_,data_stage_3__725_,data_stage_3__724_,
  data_stage_3__723_,data_stage_3__722_,data_stage_3__721_,data_stage_3__720_,data_stage_3__719_,
  data_stage_3__718_,data_stage_3__717_,data_stage_3__716_,data_stage_3__715_,
  data_stage_3__714_,data_stage_3__713_,data_stage_3__712_,data_stage_3__711_,
  data_stage_3__710_,data_stage_3__709_,data_stage_3__708_,data_stage_3__707_,
  data_stage_3__706_,data_stage_3__705_,data_stage_3__704_,data_stage_3__703_,
  data_stage_3__702_,data_stage_3__701_,data_stage_3__700_,data_stage_3__699_,data_stage_3__698_,
  data_stage_3__697_,data_stage_3__696_,data_stage_3__695_,data_stage_3__694_,
  data_stage_3__693_,data_stage_3__692_,data_stage_3__691_,data_stage_3__690_,
  data_stage_3__689_,data_stage_3__688_,data_stage_3__687_,data_stage_3__686_,
  data_stage_3__685_,data_stage_3__684_,data_stage_3__683_,data_stage_3__682_,
  data_stage_3__681_,data_stage_3__680_,data_stage_3__679_,data_stage_3__678_,data_stage_3__677_,
  data_stage_3__676_,data_stage_3__675_,data_stage_3__674_,data_stage_3__673_,
  data_stage_3__672_,data_stage_3__671_,data_stage_3__670_,data_stage_3__669_,
  data_stage_3__668_,data_stage_3__667_,data_stage_3__666_,data_stage_3__665_,
  data_stage_3__664_,data_stage_3__663_,data_stage_3__662_,data_stage_3__661_,data_stage_3__660_,
  data_stage_3__659_,data_stage_3__658_,data_stage_3__657_,data_stage_3__656_,
  data_stage_3__655_,data_stage_3__654_,data_stage_3__653_,data_stage_3__652_,
  data_stage_3__651_,data_stage_3__650_,data_stage_3__649_,data_stage_3__648_,
  data_stage_3__647_,data_stage_3__646_,data_stage_3__645_,data_stage_3__644_,
  data_stage_3__643_,data_stage_3__642_,data_stage_3__641_,data_stage_3__640_,data_stage_3__639_,
  data_stage_3__638_,data_stage_3__637_,data_stage_3__636_,data_stage_3__635_,
  data_stage_3__634_,data_stage_3__633_,data_stage_3__632_,data_stage_3__631_,
  data_stage_3__630_,data_stage_3__629_,data_stage_3__628_,data_stage_3__627_,
  data_stage_3__626_,data_stage_3__625_,data_stage_3__624_,data_stage_3__623_,
  data_stage_3__622_,data_stage_3__621_,data_stage_3__620_,data_stage_3__619_,data_stage_3__618_,
  data_stage_3__617_,data_stage_3__616_,data_stage_3__615_,data_stage_3__614_,
  data_stage_3__613_,data_stage_3__612_,data_stage_3__611_,data_stage_3__610_,
  data_stage_3__609_,data_stage_3__608_,data_stage_3__607_,data_stage_3__606_,
  data_stage_3__605_,data_stage_3__604_,data_stage_3__603_,data_stage_3__602_,
  data_stage_3__601_,data_stage_3__600_,data_stage_3__599_,data_stage_3__598_,data_stage_3__597_,
  data_stage_3__596_,data_stage_3__595_,data_stage_3__594_,data_stage_3__593_,
  data_stage_3__592_,data_stage_3__591_,data_stage_3__590_,data_stage_3__589_,
  data_stage_3__588_,data_stage_3__587_,data_stage_3__586_,data_stage_3__585_,
  data_stage_3__584_,data_stage_3__583_,data_stage_3__582_,data_stage_3__581_,data_stage_3__580_,
  data_stage_3__579_,data_stage_3__578_,data_stage_3__577_,data_stage_3__576_,
  data_stage_3__575_,data_stage_3__574_,data_stage_3__573_,data_stage_3__572_,
  data_stage_3__571_,data_stage_3__570_,data_stage_3__569_,data_stage_3__568_,
  data_stage_3__567_,data_stage_3__566_,data_stage_3__565_,data_stage_3__564_,
  data_stage_3__563_,data_stage_3__562_,data_stage_3__561_,data_stage_3__560_,data_stage_3__559_,
  data_stage_3__558_,data_stage_3__557_,data_stage_3__556_,data_stage_3__555_,
  data_stage_3__554_,data_stage_3__553_,data_stage_3__552_,data_stage_3__551_,
  data_stage_3__550_,data_stage_3__549_,data_stage_3__548_,data_stage_3__547_,
  data_stage_3__546_,data_stage_3__545_,data_stage_3__544_,data_stage_3__543_,
  data_stage_3__542_,data_stage_3__541_,data_stage_3__540_,data_stage_3__539_,data_stage_3__538_,
  data_stage_3__537_,data_stage_3__536_,data_stage_3__535_,data_stage_3__534_,
  data_stage_3__533_,data_stage_3__532_,data_stage_3__531_,data_stage_3__530_,
  data_stage_3__529_,data_stage_3__528_,data_stage_3__527_,data_stage_3__526_,
  data_stage_3__525_,data_stage_3__524_,data_stage_3__523_,data_stage_3__522_,
  data_stage_3__521_,data_stage_3__520_,data_stage_3__519_,data_stage_3__518_,data_stage_3__517_,
  data_stage_3__516_,data_stage_3__515_,data_stage_3__514_,data_stage_3__513_,
  data_stage_3__512_,data_stage_3__511_,data_stage_3__510_,data_stage_3__509_,
  data_stage_3__508_,data_stage_3__507_,data_stage_3__506_,data_stage_3__505_,
  data_stage_3__504_,data_stage_3__503_,data_stage_3__502_,data_stage_3__501_,data_stage_3__500_,
  data_stage_3__499_,data_stage_3__498_,data_stage_3__497_,data_stage_3__496_,
  data_stage_3__495_,data_stage_3__494_,data_stage_3__493_,data_stage_3__492_,
  data_stage_3__491_,data_stage_3__490_,data_stage_3__489_,data_stage_3__488_,
  data_stage_3__487_,data_stage_3__486_,data_stage_3__485_,data_stage_3__484_,
  data_stage_3__483_,data_stage_3__482_,data_stage_3__481_,data_stage_3__480_,data_stage_3__479_,
  data_stage_3__478_,data_stage_3__477_,data_stage_3__476_,data_stage_3__475_,
  data_stage_3__474_,data_stage_3__473_,data_stage_3__472_,data_stage_3__471_,
  data_stage_3__470_,data_stage_3__469_,data_stage_3__468_,data_stage_3__467_,
  data_stage_3__466_,data_stage_3__465_,data_stage_3__464_,data_stage_3__463_,
  data_stage_3__462_,data_stage_3__461_,data_stage_3__460_,data_stage_3__459_,data_stage_3__458_,
  data_stage_3__457_,data_stage_3__456_,data_stage_3__455_,data_stage_3__454_,
  data_stage_3__453_,data_stage_3__452_,data_stage_3__451_,data_stage_3__450_,
  data_stage_3__449_,data_stage_3__448_,data_stage_3__447_,data_stage_3__446_,
  data_stage_3__445_,data_stage_3__444_,data_stage_3__443_,data_stage_3__442_,
  data_stage_3__441_,data_stage_3__440_,data_stage_3__439_,data_stage_3__438_,data_stage_3__437_,
  data_stage_3__436_,data_stage_3__435_,data_stage_3__434_,data_stage_3__433_,
  data_stage_3__432_,data_stage_3__431_,data_stage_3__430_,data_stage_3__429_,
  data_stage_3__428_,data_stage_3__427_,data_stage_3__426_,data_stage_3__425_,
  data_stage_3__424_,data_stage_3__423_,data_stage_3__422_,data_stage_3__421_,data_stage_3__420_,
  data_stage_3__419_,data_stage_3__418_,data_stage_3__417_,data_stage_3__416_,
  data_stage_3__415_,data_stage_3__414_,data_stage_3__413_,data_stage_3__412_,
  data_stage_3__411_,data_stage_3__410_,data_stage_3__409_,data_stage_3__408_,
  data_stage_3__407_,data_stage_3__406_,data_stage_3__405_,data_stage_3__404_,
  data_stage_3__403_,data_stage_3__402_,data_stage_3__401_,data_stage_3__400_,data_stage_3__399_,
  data_stage_3__398_,data_stage_3__397_,data_stage_3__396_,data_stage_3__395_,
  data_stage_3__394_,data_stage_3__393_,data_stage_3__392_,data_stage_3__391_,
  data_stage_3__390_,data_stage_3__389_,data_stage_3__388_,data_stage_3__387_,
  data_stage_3__386_,data_stage_3__385_,data_stage_3__384_,data_stage_3__383_,
  data_stage_3__382_,data_stage_3__381_,data_stage_3__380_,data_stage_3__379_,data_stage_3__378_,
  data_stage_3__377_,data_stage_3__376_,data_stage_3__375_,data_stage_3__374_,
  data_stage_3__373_,data_stage_3__372_,data_stage_3__371_,data_stage_3__370_,
  data_stage_3__369_,data_stage_3__368_,data_stage_3__367_,data_stage_3__366_,
  data_stage_3__365_,data_stage_3__364_,data_stage_3__363_,data_stage_3__362_,
  data_stage_3__361_,data_stage_3__360_,data_stage_3__359_,data_stage_3__358_,data_stage_3__357_,
  data_stage_3__356_,data_stage_3__355_,data_stage_3__354_,data_stage_3__353_,
  data_stage_3__352_,data_stage_3__351_,data_stage_3__350_,data_stage_3__349_,
  data_stage_3__348_,data_stage_3__347_,data_stage_3__346_,data_stage_3__345_,
  data_stage_3__344_,data_stage_3__343_,data_stage_3__342_,data_stage_3__341_,data_stage_3__340_,
  data_stage_3__339_,data_stage_3__338_,data_stage_3__337_,data_stage_3__336_,
  data_stage_3__335_,data_stage_3__334_,data_stage_3__333_,data_stage_3__332_,
  data_stage_3__331_,data_stage_3__330_,data_stage_3__329_,data_stage_3__328_,
  data_stage_3__327_,data_stage_3__326_,data_stage_3__325_,data_stage_3__324_,
  data_stage_3__323_,data_stage_3__322_,data_stage_3__321_,data_stage_3__320_,data_stage_3__319_,
  data_stage_3__318_,data_stage_3__317_,data_stage_3__316_,data_stage_3__315_,
  data_stage_3__314_,data_stage_3__313_,data_stage_3__312_,data_stage_3__311_,
  data_stage_3__310_,data_stage_3__309_,data_stage_3__308_,data_stage_3__307_,
  data_stage_3__306_,data_stage_3__305_,data_stage_3__304_,data_stage_3__303_,
  data_stage_3__302_,data_stage_3__301_,data_stage_3__300_,data_stage_3__299_,data_stage_3__298_,
  data_stage_3__297_,data_stage_3__296_,data_stage_3__295_,data_stage_3__294_,
  data_stage_3__293_,data_stage_3__292_,data_stage_3__291_,data_stage_3__290_,
  data_stage_3__289_,data_stage_3__288_,data_stage_3__287_,data_stage_3__286_,
  data_stage_3__285_,data_stage_3__284_,data_stage_3__283_,data_stage_3__282_,
  data_stage_3__281_,data_stage_3__280_,data_stage_3__279_,data_stage_3__278_,data_stage_3__277_,
  data_stage_3__276_,data_stage_3__275_,data_stage_3__274_,data_stage_3__273_,
  data_stage_3__272_,data_stage_3__271_,data_stage_3__270_,data_stage_3__269_,
  data_stage_3__268_,data_stage_3__267_,data_stage_3__266_,data_stage_3__265_,
  data_stage_3__264_,data_stage_3__263_,data_stage_3__262_,data_stage_3__261_,data_stage_3__260_,
  data_stage_3__259_,data_stage_3__258_,data_stage_3__257_,data_stage_3__256_,
  data_stage_3__255_,data_stage_3__254_,data_stage_3__253_,data_stage_3__252_,
  data_stage_3__251_,data_stage_3__250_,data_stage_3__249_,data_stage_3__248_,
  data_stage_3__247_,data_stage_3__246_,data_stage_3__245_,data_stage_3__244_,
  data_stage_3__243_,data_stage_3__242_,data_stage_3__241_,data_stage_3__240_,data_stage_3__239_,
  data_stage_3__238_,data_stage_3__237_,data_stage_3__236_,data_stage_3__235_,
  data_stage_3__234_,data_stage_3__233_,data_stage_3__232_,data_stage_3__231_,
  data_stage_3__230_,data_stage_3__229_,data_stage_3__228_,data_stage_3__227_,
  data_stage_3__226_,data_stage_3__225_,data_stage_3__224_,data_stage_3__223_,
  data_stage_3__222_,data_stage_3__221_,data_stage_3__220_,data_stage_3__219_,data_stage_3__218_,
  data_stage_3__217_,data_stage_3__216_,data_stage_3__215_,data_stage_3__214_,
  data_stage_3__213_,data_stage_3__212_,data_stage_3__211_,data_stage_3__210_,
  data_stage_3__209_,data_stage_3__208_,data_stage_3__207_,data_stage_3__206_,
  data_stage_3__205_,data_stage_3__204_,data_stage_3__203_,data_stage_3__202_,
  data_stage_3__201_,data_stage_3__200_,data_stage_3__199_,data_stage_3__198_,data_stage_3__197_,
  data_stage_3__196_,data_stage_3__195_,data_stage_3__194_,data_stage_3__193_,
  data_stage_3__192_,data_stage_3__191_,data_stage_3__190_,data_stage_3__189_,
  data_stage_3__188_,data_stage_3__187_,data_stage_3__186_,data_stage_3__185_,
  data_stage_3__184_,data_stage_3__183_,data_stage_3__182_,data_stage_3__181_,data_stage_3__180_,
  data_stage_3__179_,data_stage_3__178_,data_stage_3__177_,data_stage_3__176_,
  data_stage_3__175_,data_stage_3__174_,data_stage_3__173_,data_stage_3__172_,
  data_stage_3__171_,data_stage_3__170_,data_stage_3__169_,data_stage_3__168_,
  data_stage_3__167_,data_stage_3__166_,data_stage_3__165_,data_stage_3__164_,
  data_stage_3__163_,data_stage_3__162_,data_stage_3__161_,data_stage_3__160_,data_stage_3__159_,
  data_stage_3__158_,data_stage_3__157_,data_stage_3__156_,data_stage_3__155_,
  data_stage_3__154_,data_stage_3__153_,data_stage_3__152_,data_stage_3__151_,
  data_stage_3__150_,data_stage_3__149_,data_stage_3__148_,data_stage_3__147_,
  data_stage_3__146_,data_stage_3__145_,data_stage_3__144_,data_stage_3__143_,
  data_stage_3__142_,data_stage_3__141_,data_stage_3__140_,data_stage_3__139_,data_stage_3__138_,
  data_stage_3__137_,data_stage_3__136_,data_stage_3__135_,data_stage_3__134_,
  data_stage_3__133_,data_stage_3__132_,data_stage_3__131_,data_stage_3__130_,
  data_stage_3__129_,data_stage_3__128_,data_stage_3__127_,data_stage_3__126_,
  data_stage_3__125_,data_stage_3__124_,data_stage_3__123_,data_stage_3__122_,
  data_stage_3__121_,data_stage_3__120_,data_stage_3__119_,data_stage_3__118_,data_stage_3__117_,
  data_stage_3__116_,data_stage_3__115_,data_stage_3__114_,data_stage_3__113_,
  data_stage_3__112_,data_stage_3__111_,data_stage_3__110_,data_stage_3__109_,
  data_stage_3__108_,data_stage_3__107_,data_stage_3__106_,data_stage_3__105_,
  data_stage_3__104_,data_stage_3__103_,data_stage_3__102_,data_stage_3__101_,data_stage_3__100_,
  data_stage_3__99_,data_stage_3__98_,data_stage_3__97_,data_stage_3__96_,
  data_stage_3__95_,data_stage_3__94_,data_stage_3__93_,data_stage_3__92_,
  data_stage_3__91_,data_stage_3__90_,data_stage_3__89_,data_stage_3__88_,data_stage_3__87_,
  data_stage_3__86_,data_stage_3__85_,data_stage_3__84_,data_stage_3__83_,
  data_stage_3__82_,data_stage_3__81_,data_stage_3__80_,data_stage_3__79_,data_stage_3__78_,
  data_stage_3__77_,data_stage_3__76_,data_stage_3__75_,data_stage_3__74_,
  data_stage_3__73_,data_stage_3__72_,data_stage_3__71_,data_stage_3__70_,data_stage_3__69_,
  data_stage_3__68_,data_stage_3__67_,data_stage_3__66_,data_stage_3__65_,
  data_stage_3__64_,data_stage_3__63_,data_stage_3__62_,data_stage_3__61_,data_stage_3__60_,
  data_stage_3__59_,data_stage_3__58_,data_stage_3__57_,data_stage_3__56_,
  data_stage_3__55_,data_stage_3__54_,data_stage_3__53_,data_stage_3__52_,
  data_stage_3__51_,data_stage_3__50_,data_stage_3__49_,data_stage_3__48_,data_stage_3__47_,
  data_stage_3__46_,data_stage_3__45_,data_stage_3__44_,data_stage_3__43_,
  data_stage_3__42_,data_stage_3__41_,data_stage_3__40_,data_stage_3__39_,data_stage_3__38_,
  data_stage_3__37_,data_stage_3__36_,data_stage_3__35_,data_stage_3__34_,
  data_stage_3__33_,data_stage_3__32_,data_stage_3__31_,data_stage_3__30_,data_stage_3__29_,
  data_stage_3__28_,data_stage_3__27_,data_stage_3__26_,data_stage_3__25_,
  data_stage_3__24_,data_stage_3__23_,data_stage_3__22_,data_stage_3__21_,data_stage_3__20_,
  data_stage_3__19_,data_stage_3__18_,data_stage_3__17_,data_stage_3__16_,
  data_stage_3__15_,data_stage_3__14_,data_stage_3__13_,data_stage_3__12_,
  data_stage_3__11_,data_stage_3__10_,data_stage_3__9_,data_stage_3__8_,data_stage_3__7_,
  data_stage_3__6_,data_stage_3__5_,data_stage_3__4_,data_stage_3__3_,data_stage_3__2_,
  data_stage_3__1_,data_stage_3__0_,data_stage_4__1023_,data_stage_4__1022_,
  data_stage_4__1021_,data_stage_4__1020_,data_stage_4__1019_,data_stage_4__1018_,
  data_stage_4__1017_,data_stage_4__1016_,data_stage_4__1015_,data_stage_4__1014_,
  data_stage_4__1013_,data_stage_4__1012_,data_stage_4__1011_,data_stage_4__1010_,
  data_stage_4__1009_,data_stage_4__1008_,data_stage_4__1007_,data_stage_4__1006_,
  data_stage_4__1005_,data_stage_4__1004_,data_stage_4__1003_,data_stage_4__1002_,
  data_stage_4__1001_,data_stage_4__1000_,data_stage_4__999_,data_stage_4__998_,
  data_stage_4__997_,data_stage_4__996_,data_stage_4__995_,data_stage_4__994_,
  data_stage_4__993_,data_stage_4__992_,data_stage_4__991_,data_stage_4__990_,data_stage_4__989_,
  data_stage_4__988_,data_stage_4__987_,data_stage_4__986_,data_stage_4__985_,
  data_stage_4__984_,data_stage_4__983_,data_stage_4__982_,data_stage_4__981_,
  data_stage_4__980_,data_stage_4__979_,data_stage_4__978_,data_stage_4__977_,
  data_stage_4__976_,data_stage_4__975_,data_stage_4__974_,data_stage_4__973_,
  data_stage_4__972_,data_stage_4__971_,data_stage_4__970_,data_stage_4__969_,data_stage_4__968_,
  data_stage_4__967_,data_stage_4__966_,data_stage_4__965_,data_stage_4__964_,
  data_stage_4__963_,data_stage_4__962_,data_stage_4__961_,data_stage_4__960_,
  data_stage_4__959_,data_stage_4__958_,data_stage_4__957_,data_stage_4__956_,
  data_stage_4__955_,data_stage_4__954_,data_stage_4__953_,data_stage_4__952_,
  data_stage_4__951_,data_stage_4__950_,data_stage_4__949_,data_stage_4__948_,data_stage_4__947_,
  data_stage_4__946_,data_stage_4__945_,data_stage_4__944_,data_stage_4__943_,
  data_stage_4__942_,data_stage_4__941_,data_stage_4__940_,data_stage_4__939_,
  data_stage_4__938_,data_stage_4__937_,data_stage_4__936_,data_stage_4__935_,
  data_stage_4__934_,data_stage_4__933_,data_stage_4__932_,data_stage_4__931_,data_stage_4__930_,
  data_stage_4__929_,data_stage_4__928_,data_stage_4__927_,data_stage_4__926_,
  data_stage_4__925_,data_stage_4__924_,data_stage_4__923_,data_stage_4__922_,
  data_stage_4__921_,data_stage_4__920_,data_stage_4__919_,data_stage_4__918_,
  data_stage_4__917_,data_stage_4__916_,data_stage_4__915_,data_stage_4__914_,
  data_stage_4__913_,data_stage_4__912_,data_stage_4__911_,data_stage_4__910_,data_stage_4__909_,
  data_stage_4__908_,data_stage_4__907_,data_stage_4__906_,data_stage_4__905_,
  data_stage_4__904_,data_stage_4__903_,data_stage_4__902_,data_stage_4__901_,
  data_stage_4__900_,data_stage_4__899_,data_stage_4__898_,data_stage_4__897_,
  data_stage_4__896_,data_stage_4__895_,data_stage_4__894_,data_stage_4__893_,
  data_stage_4__892_,data_stage_4__891_,data_stage_4__890_,data_stage_4__889_,data_stage_4__888_,
  data_stage_4__887_,data_stage_4__886_,data_stage_4__885_,data_stage_4__884_,
  data_stage_4__883_,data_stage_4__882_,data_stage_4__881_,data_stage_4__880_,
  data_stage_4__879_,data_stage_4__878_,data_stage_4__877_,data_stage_4__876_,
  data_stage_4__875_,data_stage_4__874_,data_stage_4__873_,data_stage_4__872_,
  data_stage_4__871_,data_stage_4__870_,data_stage_4__869_,data_stage_4__868_,data_stage_4__867_,
  data_stage_4__866_,data_stage_4__865_,data_stage_4__864_,data_stage_4__863_,
  data_stage_4__862_,data_stage_4__861_,data_stage_4__860_,data_stage_4__859_,
  data_stage_4__858_,data_stage_4__857_,data_stage_4__856_,data_stage_4__855_,
  data_stage_4__854_,data_stage_4__853_,data_stage_4__852_,data_stage_4__851_,data_stage_4__850_,
  data_stage_4__849_,data_stage_4__848_,data_stage_4__847_,data_stage_4__846_,
  data_stage_4__845_,data_stage_4__844_,data_stage_4__843_,data_stage_4__842_,
  data_stage_4__841_,data_stage_4__840_,data_stage_4__839_,data_stage_4__838_,
  data_stage_4__837_,data_stage_4__836_,data_stage_4__835_,data_stage_4__834_,
  data_stage_4__833_,data_stage_4__832_,data_stage_4__831_,data_stage_4__830_,data_stage_4__829_,
  data_stage_4__828_,data_stage_4__827_,data_stage_4__826_,data_stage_4__825_,
  data_stage_4__824_,data_stage_4__823_,data_stage_4__822_,data_stage_4__821_,
  data_stage_4__820_,data_stage_4__819_,data_stage_4__818_,data_stage_4__817_,
  data_stage_4__816_,data_stage_4__815_,data_stage_4__814_,data_stage_4__813_,
  data_stage_4__812_,data_stage_4__811_,data_stage_4__810_,data_stage_4__809_,data_stage_4__808_,
  data_stage_4__807_,data_stage_4__806_,data_stage_4__805_,data_stage_4__804_,
  data_stage_4__803_,data_stage_4__802_,data_stage_4__801_,data_stage_4__800_,
  data_stage_4__799_,data_stage_4__798_,data_stage_4__797_,data_stage_4__796_,
  data_stage_4__795_,data_stage_4__794_,data_stage_4__793_,data_stage_4__792_,
  data_stage_4__791_,data_stage_4__790_,data_stage_4__789_,data_stage_4__788_,data_stage_4__787_,
  data_stage_4__786_,data_stage_4__785_,data_stage_4__784_,data_stage_4__783_,
  data_stage_4__782_,data_stage_4__781_,data_stage_4__780_,data_stage_4__779_,
  data_stage_4__778_,data_stage_4__777_,data_stage_4__776_,data_stage_4__775_,
  data_stage_4__774_,data_stage_4__773_,data_stage_4__772_,data_stage_4__771_,data_stage_4__770_,
  data_stage_4__769_,data_stage_4__768_,data_stage_4__767_,data_stage_4__766_,
  data_stage_4__765_,data_stage_4__764_,data_stage_4__763_,data_stage_4__762_,
  data_stage_4__761_,data_stage_4__760_,data_stage_4__759_,data_stage_4__758_,
  data_stage_4__757_,data_stage_4__756_,data_stage_4__755_,data_stage_4__754_,
  data_stage_4__753_,data_stage_4__752_,data_stage_4__751_,data_stage_4__750_,data_stage_4__749_,
  data_stage_4__748_,data_stage_4__747_,data_stage_4__746_,data_stage_4__745_,
  data_stage_4__744_,data_stage_4__743_,data_stage_4__742_,data_stage_4__741_,
  data_stage_4__740_,data_stage_4__739_,data_stage_4__738_,data_stage_4__737_,
  data_stage_4__736_,data_stage_4__735_,data_stage_4__734_,data_stage_4__733_,
  data_stage_4__732_,data_stage_4__731_,data_stage_4__730_,data_stage_4__729_,data_stage_4__728_,
  data_stage_4__727_,data_stage_4__726_,data_stage_4__725_,data_stage_4__724_,
  data_stage_4__723_,data_stage_4__722_,data_stage_4__721_,data_stage_4__720_,
  data_stage_4__719_,data_stage_4__718_,data_stage_4__717_,data_stage_4__716_,
  data_stage_4__715_,data_stage_4__714_,data_stage_4__713_,data_stage_4__712_,
  data_stage_4__711_,data_stage_4__710_,data_stage_4__709_,data_stage_4__708_,data_stage_4__707_,
  data_stage_4__706_,data_stage_4__705_,data_stage_4__704_,data_stage_4__703_,
  data_stage_4__702_,data_stage_4__701_,data_stage_4__700_,data_stage_4__699_,
  data_stage_4__698_,data_stage_4__697_,data_stage_4__696_,data_stage_4__695_,
  data_stage_4__694_,data_stage_4__693_,data_stage_4__692_,data_stage_4__691_,data_stage_4__690_,
  data_stage_4__689_,data_stage_4__688_,data_stage_4__687_,data_stage_4__686_,
  data_stage_4__685_,data_stage_4__684_,data_stage_4__683_,data_stage_4__682_,
  data_stage_4__681_,data_stage_4__680_,data_stage_4__679_,data_stage_4__678_,
  data_stage_4__677_,data_stage_4__676_,data_stage_4__675_,data_stage_4__674_,
  data_stage_4__673_,data_stage_4__672_,data_stage_4__671_,data_stage_4__670_,data_stage_4__669_,
  data_stage_4__668_,data_stage_4__667_,data_stage_4__666_,data_stage_4__665_,
  data_stage_4__664_,data_stage_4__663_,data_stage_4__662_,data_stage_4__661_,
  data_stage_4__660_,data_stage_4__659_,data_stage_4__658_,data_stage_4__657_,
  data_stage_4__656_,data_stage_4__655_,data_stage_4__654_,data_stage_4__653_,
  data_stage_4__652_,data_stage_4__651_,data_stage_4__650_,data_stage_4__649_,data_stage_4__648_,
  data_stage_4__647_,data_stage_4__646_,data_stage_4__645_,data_stage_4__644_,
  data_stage_4__643_,data_stage_4__642_,data_stage_4__641_,data_stage_4__640_,
  data_stage_4__639_,data_stage_4__638_,data_stage_4__637_,data_stage_4__636_,
  data_stage_4__635_,data_stage_4__634_,data_stage_4__633_,data_stage_4__632_,
  data_stage_4__631_,data_stage_4__630_,data_stage_4__629_,data_stage_4__628_,data_stage_4__627_,
  data_stage_4__626_,data_stage_4__625_,data_stage_4__624_,data_stage_4__623_,
  data_stage_4__622_,data_stage_4__621_,data_stage_4__620_,data_stage_4__619_,
  data_stage_4__618_,data_stage_4__617_,data_stage_4__616_,data_stage_4__615_,
  data_stage_4__614_,data_stage_4__613_,data_stage_4__612_,data_stage_4__611_,data_stage_4__610_,
  data_stage_4__609_,data_stage_4__608_,data_stage_4__607_,data_stage_4__606_,
  data_stage_4__605_,data_stage_4__604_,data_stage_4__603_,data_stage_4__602_,
  data_stage_4__601_,data_stage_4__600_,data_stage_4__599_,data_stage_4__598_,
  data_stage_4__597_,data_stage_4__596_,data_stage_4__595_,data_stage_4__594_,
  data_stage_4__593_,data_stage_4__592_,data_stage_4__591_,data_stage_4__590_,data_stage_4__589_,
  data_stage_4__588_,data_stage_4__587_,data_stage_4__586_,data_stage_4__585_,
  data_stage_4__584_,data_stage_4__583_,data_stage_4__582_,data_stage_4__581_,
  data_stage_4__580_,data_stage_4__579_,data_stage_4__578_,data_stage_4__577_,
  data_stage_4__576_,data_stage_4__575_,data_stage_4__574_,data_stage_4__573_,
  data_stage_4__572_,data_stage_4__571_,data_stage_4__570_,data_stage_4__569_,data_stage_4__568_,
  data_stage_4__567_,data_stage_4__566_,data_stage_4__565_,data_stage_4__564_,
  data_stage_4__563_,data_stage_4__562_,data_stage_4__561_,data_stage_4__560_,
  data_stage_4__559_,data_stage_4__558_,data_stage_4__557_,data_stage_4__556_,
  data_stage_4__555_,data_stage_4__554_,data_stage_4__553_,data_stage_4__552_,
  data_stage_4__551_,data_stage_4__550_,data_stage_4__549_,data_stage_4__548_,data_stage_4__547_,
  data_stage_4__546_,data_stage_4__545_,data_stage_4__544_,data_stage_4__543_,
  data_stage_4__542_,data_stage_4__541_,data_stage_4__540_,data_stage_4__539_,
  data_stage_4__538_,data_stage_4__537_,data_stage_4__536_,data_stage_4__535_,
  data_stage_4__534_,data_stage_4__533_,data_stage_4__532_,data_stage_4__531_,data_stage_4__530_,
  data_stage_4__529_,data_stage_4__528_,data_stage_4__527_,data_stage_4__526_,
  data_stage_4__525_,data_stage_4__524_,data_stage_4__523_,data_stage_4__522_,
  data_stage_4__521_,data_stage_4__520_,data_stage_4__519_,data_stage_4__518_,
  data_stage_4__517_,data_stage_4__516_,data_stage_4__515_,data_stage_4__514_,
  data_stage_4__513_,data_stage_4__512_,data_stage_4__511_,data_stage_4__510_,data_stage_4__509_,
  data_stage_4__508_,data_stage_4__507_,data_stage_4__506_,data_stage_4__505_,
  data_stage_4__504_,data_stage_4__503_,data_stage_4__502_,data_stage_4__501_,
  data_stage_4__500_,data_stage_4__499_,data_stage_4__498_,data_stage_4__497_,
  data_stage_4__496_,data_stage_4__495_,data_stage_4__494_,data_stage_4__493_,
  data_stage_4__492_,data_stage_4__491_,data_stage_4__490_,data_stage_4__489_,data_stage_4__488_,
  data_stage_4__487_,data_stage_4__486_,data_stage_4__485_,data_stage_4__484_,
  data_stage_4__483_,data_stage_4__482_,data_stage_4__481_,data_stage_4__480_,
  data_stage_4__479_,data_stage_4__478_,data_stage_4__477_,data_stage_4__476_,
  data_stage_4__475_,data_stage_4__474_,data_stage_4__473_,data_stage_4__472_,
  data_stage_4__471_,data_stage_4__470_,data_stage_4__469_,data_stage_4__468_,data_stage_4__467_,
  data_stage_4__466_,data_stage_4__465_,data_stage_4__464_,data_stage_4__463_,
  data_stage_4__462_,data_stage_4__461_,data_stage_4__460_,data_stage_4__459_,
  data_stage_4__458_,data_stage_4__457_,data_stage_4__456_,data_stage_4__455_,
  data_stage_4__454_,data_stage_4__453_,data_stage_4__452_,data_stage_4__451_,data_stage_4__450_,
  data_stage_4__449_,data_stage_4__448_,data_stage_4__447_,data_stage_4__446_,
  data_stage_4__445_,data_stage_4__444_,data_stage_4__443_,data_stage_4__442_,
  data_stage_4__441_,data_stage_4__440_,data_stage_4__439_,data_stage_4__438_,
  data_stage_4__437_,data_stage_4__436_,data_stage_4__435_,data_stage_4__434_,
  data_stage_4__433_,data_stage_4__432_,data_stage_4__431_,data_stage_4__430_,data_stage_4__429_,
  data_stage_4__428_,data_stage_4__427_,data_stage_4__426_,data_stage_4__425_,
  data_stage_4__424_,data_stage_4__423_,data_stage_4__422_,data_stage_4__421_,
  data_stage_4__420_,data_stage_4__419_,data_stage_4__418_,data_stage_4__417_,
  data_stage_4__416_,data_stage_4__415_,data_stage_4__414_,data_stage_4__413_,
  data_stage_4__412_,data_stage_4__411_,data_stage_4__410_,data_stage_4__409_,data_stage_4__408_,
  data_stage_4__407_,data_stage_4__406_,data_stage_4__405_,data_stage_4__404_,
  data_stage_4__403_,data_stage_4__402_,data_stage_4__401_,data_stage_4__400_,
  data_stage_4__399_,data_stage_4__398_,data_stage_4__397_,data_stage_4__396_,
  data_stage_4__395_,data_stage_4__394_,data_stage_4__393_,data_stage_4__392_,
  data_stage_4__391_,data_stage_4__390_,data_stage_4__389_,data_stage_4__388_,data_stage_4__387_,
  data_stage_4__386_,data_stage_4__385_,data_stage_4__384_,data_stage_4__383_,
  data_stage_4__382_,data_stage_4__381_,data_stage_4__380_,data_stage_4__379_,
  data_stage_4__378_,data_stage_4__377_,data_stage_4__376_,data_stage_4__375_,
  data_stage_4__374_,data_stage_4__373_,data_stage_4__372_,data_stage_4__371_,data_stage_4__370_,
  data_stage_4__369_,data_stage_4__368_,data_stage_4__367_,data_stage_4__366_,
  data_stage_4__365_,data_stage_4__364_,data_stage_4__363_,data_stage_4__362_,
  data_stage_4__361_,data_stage_4__360_,data_stage_4__359_,data_stage_4__358_,
  data_stage_4__357_,data_stage_4__356_,data_stage_4__355_,data_stage_4__354_,
  data_stage_4__353_,data_stage_4__352_,data_stage_4__351_,data_stage_4__350_,data_stage_4__349_,
  data_stage_4__348_,data_stage_4__347_,data_stage_4__346_,data_stage_4__345_,
  data_stage_4__344_,data_stage_4__343_,data_stage_4__342_,data_stage_4__341_,
  data_stage_4__340_,data_stage_4__339_,data_stage_4__338_,data_stage_4__337_,
  data_stage_4__336_,data_stage_4__335_,data_stage_4__334_,data_stage_4__333_,
  data_stage_4__332_,data_stage_4__331_,data_stage_4__330_,data_stage_4__329_,data_stage_4__328_,
  data_stage_4__327_,data_stage_4__326_,data_stage_4__325_,data_stage_4__324_,
  data_stage_4__323_,data_stage_4__322_,data_stage_4__321_,data_stage_4__320_,
  data_stage_4__319_,data_stage_4__318_,data_stage_4__317_,data_stage_4__316_,
  data_stage_4__315_,data_stage_4__314_,data_stage_4__313_,data_stage_4__312_,
  data_stage_4__311_,data_stage_4__310_,data_stage_4__309_,data_stage_4__308_,data_stage_4__307_,
  data_stage_4__306_,data_stage_4__305_,data_stage_4__304_,data_stage_4__303_,
  data_stage_4__302_,data_stage_4__301_,data_stage_4__300_,data_stage_4__299_,
  data_stage_4__298_,data_stage_4__297_,data_stage_4__296_,data_stage_4__295_,
  data_stage_4__294_,data_stage_4__293_,data_stage_4__292_,data_stage_4__291_,data_stage_4__290_,
  data_stage_4__289_,data_stage_4__288_,data_stage_4__287_,data_stage_4__286_,
  data_stage_4__285_,data_stage_4__284_,data_stage_4__283_,data_stage_4__282_,
  data_stage_4__281_,data_stage_4__280_,data_stage_4__279_,data_stage_4__278_,
  data_stage_4__277_,data_stage_4__276_,data_stage_4__275_,data_stage_4__274_,
  data_stage_4__273_,data_stage_4__272_,data_stage_4__271_,data_stage_4__270_,data_stage_4__269_,
  data_stage_4__268_,data_stage_4__267_,data_stage_4__266_,data_stage_4__265_,
  data_stage_4__264_,data_stage_4__263_,data_stage_4__262_,data_stage_4__261_,
  data_stage_4__260_,data_stage_4__259_,data_stage_4__258_,data_stage_4__257_,
  data_stage_4__256_,data_stage_4__255_,data_stage_4__254_,data_stage_4__253_,
  data_stage_4__252_,data_stage_4__251_,data_stage_4__250_,data_stage_4__249_,data_stage_4__248_,
  data_stage_4__247_,data_stage_4__246_,data_stage_4__245_,data_stage_4__244_,
  data_stage_4__243_,data_stage_4__242_,data_stage_4__241_,data_stage_4__240_,
  data_stage_4__239_,data_stage_4__238_,data_stage_4__237_,data_stage_4__236_,
  data_stage_4__235_,data_stage_4__234_,data_stage_4__233_,data_stage_4__232_,
  data_stage_4__231_,data_stage_4__230_,data_stage_4__229_,data_stage_4__228_,data_stage_4__227_,
  data_stage_4__226_,data_stage_4__225_,data_stage_4__224_,data_stage_4__223_,
  data_stage_4__222_,data_stage_4__221_,data_stage_4__220_,data_stage_4__219_,
  data_stage_4__218_,data_stage_4__217_,data_stage_4__216_,data_stage_4__215_,
  data_stage_4__214_,data_stage_4__213_,data_stage_4__212_,data_stage_4__211_,data_stage_4__210_,
  data_stage_4__209_,data_stage_4__208_,data_stage_4__207_,data_stage_4__206_,
  data_stage_4__205_,data_stage_4__204_,data_stage_4__203_,data_stage_4__202_,
  data_stage_4__201_,data_stage_4__200_,data_stage_4__199_,data_stage_4__198_,
  data_stage_4__197_,data_stage_4__196_,data_stage_4__195_,data_stage_4__194_,
  data_stage_4__193_,data_stage_4__192_,data_stage_4__191_,data_stage_4__190_,data_stage_4__189_,
  data_stage_4__188_,data_stage_4__187_,data_stage_4__186_,data_stage_4__185_,
  data_stage_4__184_,data_stage_4__183_,data_stage_4__182_,data_stage_4__181_,
  data_stage_4__180_,data_stage_4__179_,data_stage_4__178_,data_stage_4__177_,
  data_stage_4__176_,data_stage_4__175_,data_stage_4__174_,data_stage_4__173_,
  data_stage_4__172_,data_stage_4__171_,data_stage_4__170_,data_stage_4__169_,data_stage_4__168_,
  data_stage_4__167_,data_stage_4__166_,data_stage_4__165_,data_stage_4__164_,
  data_stage_4__163_,data_stage_4__162_,data_stage_4__161_,data_stage_4__160_,
  data_stage_4__159_,data_stage_4__158_,data_stage_4__157_,data_stage_4__156_,
  data_stage_4__155_,data_stage_4__154_,data_stage_4__153_,data_stage_4__152_,
  data_stage_4__151_,data_stage_4__150_,data_stage_4__149_,data_stage_4__148_,data_stage_4__147_,
  data_stage_4__146_,data_stage_4__145_,data_stage_4__144_,data_stage_4__143_,
  data_stage_4__142_,data_stage_4__141_,data_stage_4__140_,data_stage_4__139_,
  data_stage_4__138_,data_stage_4__137_,data_stage_4__136_,data_stage_4__135_,
  data_stage_4__134_,data_stage_4__133_,data_stage_4__132_,data_stage_4__131_,data_stage_4__130_,
  data_stage_4__129_,data_stage_4__128_,data_stage_4__127_,data_stage_4__126_,
  data_stage_4__125_,data_stage_4__124_,data_stage_4__123_,data_stage_4__122_,
  data_stage_4__121_,data_stage_4__120_,data_stage_4__119_,data_stage_4__118_,
  data_stage_4__117_,data_stage_4__116_,data_stage_4__115_,data_stage_4__114_,
  data_stage_4__113_,data_stage_4__112_,data_stage_4__111_,data_stage_4__110_,data_stage_4__109_,
  data_stage_4__108_,data_stage_4__107_,data_stage_4__106_,data_stage_4__105_,
  data_stage_4__104_,data_stage_4__103_,data_stage_4__102_,data_stage_4__101_,
  data_stage_4__100_,data_stage_4__99_,data_stage_4__98_,data_stage_4__97_,
  data_stage_4__96_,data_stage_4__95_,data_stage_4__94_,data_stage_4__93_,data_stage_4__92_,
  data_stage_4__91_,data_stage_4__90_,data_stage_4__89_,data_stage_4__88_,
  data_stage_4__87_,data_stage_4__86_,data_stage_4__85_,data_stage_4__84_,data_stage_4__83_,
  data_stage_4__82_,data_stage_4__81_,data_stage_4__80_,data_stage_4__79_,
  data_stage_4__78_,data_stage_4__77_,data_stage_4__76_,data_stage_4__75_,data_stage_4__74_,
  data_stage_4__73_,data_stage_4__72_,data_stage_4__71_,data_stage_4__70_,
  data_stage_4__69_,data_stage_4__68_,data_stage_4__67_,data_stage_4__66_,data_stage_4__65_,
  data_stage_4__64_,data_stage_4__63_,data_stage_4__62_,data_stage_4__61_,
  data_stage_4__60_,data_stage_4__59_,data_stage_4__58_,data_stage_4__57_,
  data_stage_4__56_,data_stage_4__55_,data_stage_4__54_,data_stage_4__53_,data_stage_4__52_,
  data_stage_4__51_,data_stage_4__50_,data_stage_4__49_,data_stage_4__48_,
  data_stage_4__47_,data_stage_4__46_,data_stage_4__45_,data_stage_4__44_,data_stage_4__43_,
  data_stage_4__42_,data_stage_4__41_,data_stage_4__40_,data_stage_4__39_,
  data_stage_4__38_,data_stage_4__37_,data_stage_4__36_,data_stage_4__35_,data_stage_4__34_,
  data_stage_4__33_,data_stage_4__32_,data_stage_4__31_,data_stage_4__30_,
  data_stage_4__29_,data_stage_4__28_,data_stage_4__27_,data_stage_4__26_,data_stage_4__25_,
  data_stage_4__24_,data_stage_4__23_,data_stage_4__22_,data_stage_4__21_,
  data_stage_4__20_,data_stage_4__19_,data_stage_4__18_,data_stage_4__17_,
  data_stage_4__16_,data_stage_4__15_,data_stage_4__14_,data_stage_4__13_,data_stage_4__12_,
  data_stage_4__11_,data_stage_4__10_,data_stage_4__9_,data_stage_4__8_,
  data_stage_4__7_,data_stage_4__6_,data_stage_4__5_,data_stage_4__4_,data_stage_4__3_,
  data_stage_4__2_,data_stage_4__1_,data_stage_4__0_;

  bsg_swap_width_p32
  mux_stage_0__mux_swap_0__swap_inst
  (
    .data_i(data_i[63:0]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_1__swap_inst
  (
    .data_i(data_i[127:64]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_2__swap_inst
  (
    .data_i(data_i[191:128]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_3__swap_inst
  (
    .data_i(data_i[255:192]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_4__swap_inst
  (
    .data_i(data_i[319:256]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_5__swap_inst
  (
    .data_i(data_i[383:320]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_6__swap_inst
  (
    .data_i(data_i[447:384]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_7__swap_inst
  (
    .data_i(data_i[511:448]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_8__swap_inst
  (
    .data_i(data_i[575:512]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__575_, data_stage_1__574_, data_stage_1__573_, data_stage_1__572_, data_stage_1__571_, data_stage_1__570_, data_stage_1__569_, data_stage_1__568_, data_stage_1__567_, data_stage_1__566_, data_stage_1__565_, data_stage_1__564_, data_stage_1__563_, data_stage_1__562_, data_stage_1__561_, data_stage_1__560_, data_stage_1__559_, data_stage_1__558_, data_stage_1__557_, data_stage_1__556_, data_stage_1__555_, data_stage_1__554_, data_stage_1__553_, data_stage_1__552_, data_stage_1__551_, data_stage_1__550_, data_stage_1__549_, data_stage_1__548_, data_stage_1__547_, data_stage_1__546_, data_stage_1__545_, data_stage_1__544_, data_stage_1__543_, data_stage_1__542_, data_stage_1__541_, data_stage_1__540_, data_stage_1__539_, data_stage_1__538_, data_stage_1__537_, data_stage_1__536_, data_stage_1__535_, data_stage_1__534_, data_stage_1__533_, data_stage_1__532_, data_stage_1__531_, data_stage_1__530_, data_stage_1__529_, data_stage_1__528_, data_stage_1__527_, data_stage_1__526_, data_stage_1__525_, data_stage_1__524_, data_stage_1__523_, data_stage_1__522_, data_stage_1__521_, data_stage_1__520_, data_stage_1__519_, data_stage_1__518_, data_stage_1__517_, data_stage_1__516_, data_stage_1__515_, data_stage_1__514_, data_stage_1__513_, data_stage_1__512_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_9__swap_inst
  (
    .data_i(data_i[639:576]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__639_, data_stage_1__638_, data_stage_1__637_, data_stage_1__636_, data_stage_1__635_, data_stage_1__634_, data_stage_1__633_, data_stage_1__632_, data_stage_1__631_, data_stage_1__630_, data_stage_1__629_, data_stage_1__628_, data_stage_1__627_, data_stage_1__626_, data_stage_1__625_, data_stage_1__624_, data_stage_1__623_, data_stage_1__622_, data_stage_1__621_, data_stage_1__620_, data_stage_1__619_, data_stage_1__618_, data_stage_1__617_, data_stage_1__616_, data_stage_1__615_, data_stage_1__614_, data_stage_1__613_, data_stage_1__612_, data_stage_1__611_, data_stage_1__610_, data_stage_1__609_, data_stage_1__608_, data_stage_1__607_, data_stage_1__606_, data_stage_1__605_, data_stage_1__604_, data_stage_1__603_, data_stage_1__602_, data_stage_1__601_, data_stage_1__600_, data_stage_1__599_, data_stage_1__598_, data_stage_1__597_, data_stage_1__596_, data_stage_1__595_, data_stage_1__594_, data_stage_1__593_, data_stage_1__592_, data_stage_1__591_, data_stage_1__590_, data_stage_1__589_, data_stage_1__588_, data_stage_1__587_, data_stage_1__586_, data_stage_1__585_, data_stage_1__584_, data_stage_1__583_, data_stage_1__582_, data_stage_1__581_, data_stage_1__580_, data_stage_1__579_, data_stage_1__578_, data_stage_1__577_, data_stage_1__576_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_10__swap_inst
  (
    .data_i(data_i[703:640]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__703_, data_stage_1__702_, data_stage_1__701_, data_stage_1__700_, data_stage_1__699_, data_stage_1__698_, data_stage_1__697_, data_stage_1__696_, data_stage_1__695_, data_stage_1__694_, data_stage_1__693_, data_stage_1__692_, data_stage_1__691_, data_stage_1__690_, data_stage_1__689_, data_stage_1__688_, data_stage_1__687_, data_stage_1__686_, data_stage_1__685_, data_stage_1__684_, data_stage_1__683_, data_stage_1__682_, data_stage_1__681_, data_stage_1__680_, data_stage_1__679_, data_stage_1__678_, data_stage_1__677_, data_stage_1__676_, data_stage_1__675_, data_stage_1__674_, data_stage_1__673_, data_stage_1__672_, data_stage_1__671_, data_stage_1__670_, data_stage_1__669_, data_stage_1__668_, data_stage_1__667_, data_stage_1__666_, data_stage_1__665_, data_stage_1__664_, data_stage_1__663_, data_stage_1__662_, data_stage_1__661_, data_stage_1__660_, data_stage_1__659_, data_stage_1__658_, data_stage_1__657_, data_stage_1__656_, data_stage_1__655_, data_stage_1__654_, data_stage_1__653_, data_stage_1__652_, data_stage_1__651_, data_stage_1__650_, data_stage_1__649_, data_stage_1__648_, data_stage_1__647_, data_stage_1__646_, data_stage_1__645_, data_stage_1__644_, data_stage_1__643_, data_stage_1__642_, data_stage_1__641_, data_stage_1__640_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_11__swap_inst
  (
    .data_i(data_i[767:704]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__767_, data_stage_1__766_, data_stage_1__765_, data_stage_1__764_, data_stage_1__763_, data_stage_1__762_, data_stage_1__761_, data_stage_1__760_, data_stage_1__759_, data_stage_1__758_, data_stage_1__757_, data_stage_1__756_, data_stage_1__755_, data_stage_1__754_, data_stage_1__753_, data_stage_1__752_, data_stage_1__751_, data_stage_1__750_, data_stage_1__749_, data_stage_1__748_, data_stage_1__747_, data_stage_1__746_, data_stage_1__745_, data_stage_1__744_, data_stage_1__743_, data_stage_1__742_, data_stage_1__741_, data_stage_1__740_, data_stage_1__739_, data_stage_1__738_, data_stage_1__737_, data_stage_1__736_, data_stage_1__735_, data_stage_1__734_, data_stage_1__733_, data_stage_1__732_, data_stage_1__731_, data_stage_1__730_, data_stage_1__729_, data_stage_1__728_, data_stage_1__727_, data_stage_1__726_, data_stage_1__725_, data_stage_1__724_, data_stage_1__723_, data_stage_1__722_, data_stage_1__721_, data_stage_1__720_, data_stage_1__719_, data_stage_1__718_, data_stage_1__717_, data_stage_1__716_, data_stage_1__715_, data_stage_1__714_, data_stage_1__713_, data_stage_1__712_, data_stage_1__711_, data_stage_1__710_, data_stage_1__709_, data_stage_1__708_, data_stage_1__707_, data_stage_1__706_, data_stage_1__705_, data_stage_1__704_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_12__swap_inst
  (
    .data_i(data_i[831:768]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__831_, data_stage_1__830_, data_stage_1__829_, data_stage_1__828_, data_stage_1__827_, data_stage_1__826_, data_stage_1__825_, data_stage_1__824_, data_stage_1__823_, data_stage_1__822_, data_stage_1__821_, data_stage_1__820_, data_stage_1__819_, data_stage_1__818_, data_stage_1__817_, data_stage_1__816_, data_stage_1__815_, data_stage_1__814_, data_stage_1__813_, data_stage_1__812_, data_stage_1__811_, data_stage_1__810_, data_stage_1__809_, data_stage_1__808_, data_stage_1__807_, data_stage_1__806_, data_stage_1__805_, data_stage_1__804_, data_stage_1__803_, data_stage_1__802_, data_stage_1__801_, data_stage_1__800_, data_stage_1__799_, data_stage_1__798_, data_stage_1__797_, data_stage_1__796_, data_stage_1__795_, data_stage_1__794_, data_stage_1__793_, data_stage_1__792_, data_stage_1__791_, data_stage_1__790_, data_stage_1__789_, data_stage_1__788_, data_stage_1__787_, data_stage_1__786_, data_stage_1__785_, data_stage_1__784_, data_stage_1__783_, data_stage_1__782_, data_stage_1__781_, data_stage_1__780_, data_stage_1__779_, data_stage_1__778_, data_stage_1__777_, data_stage_1__776_, data_stage_1__775_, data_stage_1__774_, data_stage_1__773_, data_stage_1__772_, data_stage_1__771_, data_stage_1__770_, data_stage_1__769_, data_stage_1__768_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_13__swap_inst
  (
    .data_i(data_i[895:832]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__895_, data_stage_1__894_, data_stage_1__893_, data_stage_1__892_, data_stage_1__891_, data_stage_1__890_, data_stage_1__889_, data_stage_1__888_, data_stage_1__887_, data_stage_1__886_, data_stage_1__885_, data_stage_1__884_, data_stage_1__883_, data_stage_1__882_, data_stage_1__881_, data_stage_1__880_, data_stage_1__879_, data_stage_1__878_, data_stage_1__877_, data_stage_1__876_, data_stage_1__875_, data_stage_1__874_, data_stage_1__873_, data_stage_1__872_, data_stage_1__871_, data_stage_1__870_, data_stage_1__869_, data_stage_1__868_, data_stage_1__867_, data_stage_1__866_, data_stage_1__865_, data_stage_1__864_, data_stage_1__863_, data_stage_1__862_, data_stage_1__861_, data_stage_1__860_, data_stage_1__859_, data_stage_1__858_, data_stage_1__857_, data_stage_1__856_, data_stage_1__855_, data_stage_1__854_, data_stage_1__853_, data_stage_1__852_, data_stage_1__851_, data_stage_1__850_, data_stage_1__849_, data_stage_1__848_, data_stage_1__847_, data_stage_1__846_, data_stage_1__845_, data_stage_1__844_, data_stage_1__843_, data_stage_1__842_, data_stage_1__841_, data_stage_1__840_, data_stage_1__839_, data_stage_1__838_, data_stage_1__837_, data_stage_1__836_, data_stage_1__835_, data_stage_1__834_, data_stage_1__833_, data_stage_1__832_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_14__swap_inst
  (
    .data_i(data_i[959:896]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__959_, data_stage_1__958_, data_stage_1__957_, data_stage_1__956_, data_stage_1__955_, data_stage_1__954_, data_stage_1__953_, data_stage_1__952_, data_stage_1__951_, data_stage_1__950_, data_stage_1__949_, data_stage_1__948_, data_stage_1__947_, data_stage_1__946_, data_stage_1__945_, data_stage_1__944_, data_stage_1__943_, data_stage_1__942_, data_stage_1__941_, data_stage_1__940_, data_stage_1__939_, data_stage_1__938_, data_stage_1__937_, data_stage_1__936_, data_stage_1__935_, data_stage_1__934_, data_stage_1__933_, data_stage_1__932_, data_stage_1__931_, data_stage_1__930_, data_stage_1__929_, data_stage_1__928_, data_stage_1__927_, data_stage_1__926_, data_stage_1__925_, data_stage_1__924_, data_stage_1__923_, data_stage_1__922_, data_stage_1__921_, data_stage_1__920_, data_stage_1__919_, data_stage_1__918_, data_stage_1__917_, data_stage_1__916_, data_stage_1__915_, data_stage_1__914_, data_stage_1__913_, data_stage_1__912_, data_stage_1__911_, data_stage_1__910_, data_stage_1__909_, data_stage_1__908_, data_stage_1__907_, data_stage_1__906_, data_stage_1__905_, data_stage_1__904_, data_stage_1__903_, data_stage_1__902_, data_stage_1__901_, data_stage_1__900_, data_stage_1__899_, data_stage_1__898_, data_stage_1__897_, data_stage_1__896_ })
  );


  bsg_swap_width_p32
  mux_stage_0__mux_swap_15__swap_inst
  (
    .data_i(data_i[1023:960]),
    .swap_i(sel_i[0]),
    .data_o({ data_stage_1__1023_, data_stage_1__1022_, data_stage_1__1021_, data_stage_1__1020_, data_stage_1__1019_, data_stage_1__1018_, data_stage_1__1017_, data_stage_1__1016_, data_stage_1__1015_, data_stage_1__1014_, data_stage_1__1013_, data_stage_1__1012_, data_stage_1__1011_, data_stage_1__1010_, data_stage_1__1009_, data_stage_1__1008_, data_stage_1__1007_, data_stage_1__1006_, data_stage_1__1005_, data_stage_1__1004_, data_stage_1__1003_, data_stage_1__1002_, data_stage_1__1001_, data_stage_1__1000_, data_stage_1__999_, data_stage_1__998_, data_stage_1__997_, data_stage_1__996_, data_stage_1__995_, data_stage_1__994_, data_stage_1__993_, data_stage_1__992_, data_stage_1__991_, data_stage_1__990_, data_stage_1__989_, data_stage_1__988_, data_stage_1__987_, data_stage_1__986_, data_stage_1__985_, data_stage_1__984_, data_stage_1__983_, data_stage_1__982_, data_stage_1__981_, data_stage_1__980_, data_stage_1__979_, data_stage_1__978_, data_stage_1__977_, data_stage_1__976_, data_stage_1__975_, data_stage_1__974_, data_stage_1__973_, data_stage_1__972_, data_stage_1__971_, data_stage_1__970_, data_stage_1__969_, data_stage_1__968_, data_stage_1__967_, data_stage_1__966_, data_stage_1__965_, data_stage_1__964_, data_stage_1__963_, data_stage_1__962_, data_stage_1__961_, data_stage_1__960_ })
  );


  bsg_swap_width_p64
  mux_stage_1__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_1__127_, data_stage_1__126_, data_stage_1__125_, data_stage_1__124_, data_stage_1__123_, data_stage_1__122_, data_stage_1__121_, data_stage_1__120_, data_stage_1__119_, data_stage_1__118_, data_stage_1__117_, data_stage_1__116_, data_stage_1__115_, data_stage_1__114_, data_stage_1__113_, data_stage_1__112_, data_stage_1__111_, data_stage_1__110_, data_stage_1__109_, data_stage_1__108_, data_stage_1__107_, data_stage_1__106_, data_stage_1__105_, data_stage_1__104_, data_stage_1__103_, data_stage_1__102_, data_stage_1__101_, data_stage_1__100_, data_stage_1__99_, data_stage_1__98_, data_stage_1__97_, data_stage_1__96_, data_stage_1__95_, data_stage_1__94_, data_stage_1__93_, data_stage_1__92_, data_stage_1__91_, data_stage_1__90_, data_stage_1__89_, data_stage_1__88_, data_stage_1__87_, data_stage_1__86_, data_stage_1__85_, data_stage_1__84_, data_stage_1__83_, data_stage_1__82_, data_stage_1__81_, data_stage_1__80_, data_stage_1__79_, data_stage_1__78_, data_stage_1__77_, data_stage_1__76_, data_stage_1__75_, data_stage_1__74_, data_stage_1__73_, data_stage_1__72_, data_stage_1__71_, data_stage_1__70_, data_stage_1__69_, data_stage_1__68_, data_stage_1__67_, data_stage_1__66_, data_stage_1__65_, data_stage_1__64_, data_stage_1__63_, data_stage_1__62_, data_stage_1__61_, data_stage_1__60_, data_stage_1__59_, data_stage_1__58_, data_stage_1__57_, data_stage_1__56_, data_stage_1__55_, data_stage_1__54_, data_stage_1__53_, data_stage_1__52_, data_stage_1__51_, data_stage_1__50_, data_stage_1__49_, data_stage_1__48_, data_stage_1__47_, data_stage_1__46_, data_stage_1__45_, data_stage_1__44_, data_stage_1__43_, data_stage_1__42_, data_stage_1__41_, data_stage_1__40_, data_stage_1__39_, data_stage_1__38_, data_stage_1__37_, data_stage_1__36_, data_stage_1__35_, data_stage_1__34_, data_stage_1__33_, data_stage_1__32_, data_stage_1__31_, data_stage_1__30_, data_stage_1__29_, data_stage_1__28_, data_stage_1__27_, data_stage_1__26_, data_stage_1__25_, data_stage_1__24_, data_stage_1__23_, data_stage_1__22_, data_stage_1__21_, data_stage_1__20_, data_stage_1__19_, data_stage_1__18_, data_stage_1__17_, data_stage_1__16_, data_stage_1__15_, data_stage_1__14_, data_stage_1__13_, data_stage_1__12_, data_stage_1__11_, data_stage_1__10_, data_stage_1__9_, data_stage_1__8_, data_stage_1__7_, data_stage_1__6_, data_stage_1__5_, data_stage_1__4_, data_stage_1__3_, data_stage_1__2_, data_stage_1__1_, data_stage_1__0_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ })
  );


  bsg_swap_width_p64
  mux_stage_1__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_1__255_, data_stage_1__254_, data_stage_1__253_, data_stage_1__252_, data_stage_1__251_, data_stage_1__250_, data_stage_1__249_, data_stage_1__248_, data_stage_1__247_, data_stage_1__246_, data_stage_1__245_, data_stage_1__244_, data_stage_1__243_, data_stage_1__242_, data_stage_1__241_, data_stage_1__240_, data_stage_1__239_, data_stage_1__238_, data_stage_1__237_, data_stage_1__236_, data_stage_1__235_, data_stage_1__234_, data_stage_1__233_, data_stage_1__232_, data_stage_1__231_, data_stage_1__230_, data_stage_1__229_, data_stage_1__228_, data_stage_1__227_, data_stage_1__226_, data_stage_1__225_, data_stage_1__224_, data_stage_1__223_, data_stage_1__222_, data_stage_1__221_, data_stage_1__220_, data_stage_1__219_, data_stage_1__218_, data_stage_1__217_, data_stage_1__216_, data_stage_1__215_, data_stage_1__214_, data_stage_1__213_, data_stage_1__212_, data_stage_1__211_, data_stage_1__210_, data_stage_1__209_, data_stage_1__208_, data_stage_1__207_, data_stage_1__206_, data_stage_1__205_, data_stage_1__204_, data_stage_1__203_, data_stage_1__202_, data_stage_1__201_, data_stage_1__200_, data_stage_1__199_, data_stage_1__198_, data_stage_1__197_, data_stage_1__196_, data_stage_1__195_, data_stage_1__194_, data_stage_1__193_, data_stage_1__192_, data_stage_1__191_, data_stage_1__190_, data_stage_1__189_, data_stage_1__188_, data_stage_1__187_, data_stage_1__186_, data_stage_1__185_, data_stage_1__184_, data_stage_1__183_, data_stage_1__182_, data_stage_1__181_, data_stage_1__180_, data_stage_1__179_, data_stage_1__178_, data_stage_1__177_, data_stage_1__176_, data_stage_1__175_, data_stage_1__174_, data_stage_1__173_, data_stage_1__172_, data_stage_1__171_, data_stage_1__170_, data_stage_1__169_, data_stage_1__168_, data_stage_1__167_, data_stage_1__166_, data_stage_1__165_, data_stage_1__164_, data_stage_1__163_, data_stage_1__162_, data_stage_1__161_, data_stage_1__160_, data_stage_1__159_, data_stage_1__158_, data_stage_1__157_, data_stage_1__156_, data_stage_1__155_, data_stage_1__154_, data_stage_1__153_, data_stage_1__152_, data_stage_1__151_, data_stage_1__150_, data_stage_1__149_, data_stage_1__148_, data_stage_1__147_, data_stage_1__146_, data_stage_1__145_, data_stage_1__144_, data_stage_1__143_, data_stage_1__142_, data_stage_1__141_, data_stage_1__140_, data_stage_1__139_, data_stage_1__138_, data_stage_1__137_, data_stage_1__136_, data_stage_1__135_, data_stage_1__134_, data_stage_1__133_, data_stage_1__132_, data_stage_1__131_, data_stage_1__130_, data_stage_1__129_, data_stage_1__128_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_ })
  );


  bsg_swap_width_p64
  mux_stage_1__mux_swap_2__swap_inst
  (
    .data_i({ data_stage_1__383_, data_stage_1__382_, data_stage_1__381_, data_stage_1__380_, data_stage_1__379_, data_stage_1__378_, data_stage_1__377_, data_stage_1__376_, data_stage_1__375_, data_stage_1__374_, data_stage_1__373_, data_stage_1__372_, data_stage_1__371_, data_stage_1__370_, data_stage_1__369_, data_stage_1__368_, data_stage_1__367_, data_stage_1__366_, data_stage_1__365_, data_stage_1__364_, data_stage_1__363_, data_stage_1__362_, data_stage_1__361_, data_stage_1__360_, data_stage_1__359_, data_stage_1__358_, data_stage_1__357_, data_stage_1__356_, data_stage_1__355_, data_stage_1__354_, data_stage_1__353_, data_stage_1__352_, data_stage_1__351_, data_stage_1__350_, data_stage_1__349_, data_stage_1__348_, data_stage_1__347_, data_stage_1__346_, data_stage_1__345_, data_stage_1__344_, data_stage_1__343_, data_stage_1__342_, data_stage_1__341_, data_stage_1__340_, data_stage_1__339_, data_stage_1__338_, data_stage_1__337_, data_stage_1__336_, data_stage_1__335_, data_stage_1__334_, data_stage_1__333_, data_stage_1__332_, data_stage_1__331_, data_stage_1__330_, data_stage_1__329_, data_stage_1__328_, data_stage_1__327_, data_stage_1__326_, data_stage_1__325_, data_stage_1__324_, data_stage_1__323_, data_stage_1__322_, data_stage_1__321_, data_stage_1__320_, data_stage_1__319_, data_stage_1__318_, data_stage_1__317_, data_stage_1__316_, data_stage_1__315_, data_stage_1__314_, data_stage_1__313_, data_stage_1__312_, data_stage_1__311_, data_stage_1__310_, data_stage_1__309_, data_stage_1__308_, data_stage_1__307_, data_stage_1__306_, data_stage_1__305_, data_stage_1__304_, data_stage_1__303_, data_stage_1__302_, data_stage_1__301_, data_stage_1__300_, data_stage_1__299_, data_stage_1__298_, data_stage_1__297_, data_stage_1__296_, data_stage_1__295_, data_stage_1__294_, data_stage_1__293_, data_stage_1__292_, data_stage_1__291_, data_stage_1__290_, data_stage_1__289_, data_stage_1__288_, data_stage_1__287_, data_stage_1__286_, data_stage_1__285_, data_stage_1__284_, data_stage_1__283_, data_stage_1__282_, data_stage_1__281_, data_stage_1__280_, data_stage_1__279_, data_stage_1__278_, data_stage_1__277_, data_stage_1__276_, data_stage_1__275_, data_stage_1__274_, data_stage_1__273_, data_stage_1__272_, data_stage_1__271_, data_stage_1__270_, data_stage_1__269_, data_stage_1__268_, data_stage_1__267_, data_stage_1__266_, data_stage_1__265_, data_stage_1__264_, data_stage_1__263_, data_stage_1__262_, data_stage_1__261_, data_stage_1__260_, data_stage_1__259_, data_stage_1__258_, data_stage_1__257_, data_stage_1__256_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_ })
  );


  bsg_swap_width_p64
  mux_stage_1__mux_swap_3__swap_inst
  (
    .data_i({ data_stage_1__511_, data_stage_1__510_, data_stage_1__509_, data_stage_1__508_, data_stage_1__507_, data_stage_1__506_, data_stage_1__505_, data_stage_1__504_, data_stage_1__503_, data_stage_1__502_, data_stage_1__501_, data_stage_1__500_, data_stage_1__499_, data_stage_1__498_, data_stage_1__497_, data_stage_1__496_, data_stage_1__495_, data_stage_1__494_, data_stage_1__493_, data_stage_1__492_, data_stage_1__491_, data_stage_1__490_, data_stage_1__489_, data_stage_1__488_, data_stage_1__487_, data_stage_1__486_, data_stage_1__485_, data_stage_1__484_, data_stage_1__483_, data_stage_1__482_, data_stage_1__481_, data_stage_1__480_, data_stage_1__479_, data_stage_1__478_, data_stage_1__477_, data_stage_1__476_, data_stage_1__475_, data_stage_1__474_, data_stage_1__473_, data_stage_1__472_, data_stage_1__471_, data_stage_1__470_, data_stage_1__469_, data_stage_1__468_, data_stage_1__467_, data_stage_1__466_, data_stage_1__465_, data_stage_1__464_, data_stage_1__463_, data_stage_1__462_, data_stage_1__461_, data_stage_1__460_, data_stage_1__459_, data_stage_1__458_, data_stage_1__457_, data_stage_1__456_, data_stage_1__455_, data_stage_1__454_, data_stage_1__453_, data_stage_1__452_, data_stage_1__451_, data_stage_1__450_, data_stage_1__449_, data_stage_1__448_, data_stage_1__447_, data_stage_1__446_, data_stage_1__445_, data_stage_1__444_, data_stage_1__443_, data_stage_1__442_, data_stage_1__441_, data_stage_1__440_, data_stage_1__439_, data_stage_1__438_, data_stage_1__437_, data_stage_1__436_, data_stage_1__435_, data_stage_1__434_, data_stage_1__433_, data_stage_1__432_, data_stage_1__431_, data_stage_1__430_, data_stage_1__429_, data_stage_1__428_, data_stage_1__427_, data_stage_1__426_, data_stage_1__425_, data_stage_1__424_, data_stage_1__423_, data_stage_1__422_, data_stage_1__421_, data_stage_1__420_, data_stage_1__419_, data_stage_1__418_, data_stage_1__417_, data_stage_1__416_, data_stage_1__415_, data_stage_1__414_, data_stage_1__413_, data_stage_1__412_, data_stage_1__411_, data_stage_1__410_, data_stage_1__409_, data_stage_1__408_, data_stage_1__407_, data_stage_1__406_, data_stage_1__405_, data_stage_1__404_, data_stage_1__403_, data_stage_1__402_, data_stage_1__401_, data_stage_1__400_, data_stage_1__399_, data_stage_1__398_, data_stage_1__397_, data_stage_1__396_, data_stage_1__395_, data_stage_1__394_, data_stage_1__393_, data_stage_1__392_, data_stage_1__391_, data_stage_1__390_, data_stage_1__389_, data_stage_1__388_, data_stage_1__387_, data_stage_1__386_, data_stage_1__385_, data_stage_1__384_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_ })
  );


  bsg_swap_width_p64
  mux_stage_1__mux_swap_4__swap_inst
  (
    .data_i({ data_stage_1__639_, data_stage_1__638_, data_stage_1__637_, data_stage_1__636_, data_stage_1__635_, data_stage_1__634_, data_stage_1__633_, data_stage_1__632_, data_stage_1__631_, data_stage_1__630_, data_stage_1__629_, data_stage_1__628_, data_stage_1__627_, data_stage_1__626_, data_stage_1__625_, data_stage_1__624_, data_stage_1__623_, data_stage_1__622_, data_stage_1__621_, data_stage_1__620_, data_stage_1__619_, data_stage_1__618_, data_stage_1__617_, data_stage_1__616_, data_stage_1__615_, data_stage_1__614_, data_stage_1__613_, data_stage_1__612_, data_stage_1__611_, data_stage_1__610_, data_stage_1__609_, data_stage_1__608_, data_stage_1__607_, data_stage_1__606_, data_stage_1__605_, data_stage_1__604_, data_stage_1__603_, data_stage_1__602_, data_stage_1__601_, data_stage_1__600_, data_stage_1__599_, data_stage_1__598_, data_stage_1__597_, data_stage_1__596_, data_stage_1__595_, data_stage_1__594_, data_stage_1__593_, data_stage_1__592_, data_stage_1__591_, data_stage_1__590_, data_stage_1__589_, data_stage_1__588_, data_stage_1__587_, data_stage_1__586_, data_stage_1__585_, data_stage_1__584_, data_stage_1__583_, data_stage_1__582_, data_stage_1__581_, data_stage_1__580_, data_stage_1__579_, data_stage_1__578_, data_stage_1__577_, data_stage_1__576_, data_stage_1__575_, data_stage_1__574_, data_stage_1__573_, data_stage_1__572_, data_stage_1__571_, data_stage_1__570_, data_stage_1__569_, data_stage_1__568_, data_stage_1__567_, data_stage_1__566_, data_stage_1__565_, data_stage_1__564_, data_stage_1__563_, data_stage_1__562_, data_stage_1__561_, data_stage_1__560_, data_stage_1__559_, data_stage_1__558_, data_stage_1__557_, data_stage_1__556_, data_stage_1__555_, data_stage_1__554_, data_stage_1__553_, data_stage_1__552_, data_stage_1__551_, data_stage_1__550_, data_stage_1__549_, data_stage_1__548_, data_stage_1__547_, data_stage_1__546_, data_stage_1__545_, data_stage_1__544_, data_stage_1__543_, data_stage_1__542_, data_stage_1__541_, data_stage_1__540_, data_stage_1__539_, data_stage_1__538_, data_stage_1__537_, data_stage_1__536_, data_stage_1__535_, data_stage_1__534_, data_stage_1__533_, data_stage_1__532_, data_stage_1__531_, data_stage_1__530_, data_stage_1__529_, data_stage_1__528_, data_stage_1__527_, data_stage_1__526_, data_stage_1__525_, data_stage_1__524_, data_stage_1__523_, data_stage_1__522_, data_stage_1__521_, data_stage_1__520_, data_stage_1__519_, data_stage_1__518_, data_stage_1__517_, data_stage_1__516_, data_stage_1__515_, data_stage_1__514_, data_stage_1__513_, data_stage_1__512_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__639_, data_stage_2__638_, data_stage_2__637_, data_stage_2__636_, data_stage_2__635_, data_stage_2__634_, data_stage_2__633_, data_stage_2__632_, data_stage_2__631_, data_stage_2__630_, data_stage_2__629_, data_stage_2__628_, data_stage_2__627_, data_stage_2__626_, data_stage_2__625_, data_stage_2__624_, data_stage_2__623_, data_stage_2__622_, data_stage_2__621_, data_stage_2__620_, data_stage_2__619_, data_stage_2__618_, data_stage_2__617_, data_stage_2__616_, data_stage_2__615_, data_stage_2__614_, data_stage_2__613_, data_stage_2__612_, data_stage_2__611_, data_stage_2__610_, data_stage_2__609_, data_stage_2__608_, data_stage_2__607_, data_stage_2__606_, data_stage_2__605_, data_stage_2__604_, data_stage_2__603_, data_stage_2__602_, data_stage_2__601_, data_stage_2__600_, data_stage_2__599_, data_stage_2__598_, data_stage_2__597_, data_stage_2__596_, data_stage_2__595_, data_stage_2__594_, data_stage_2__593_, data_stage_2__592_, data_stage_2__591_, data_stage_2__590_, data_stage_2__589_, data_stage_2__588_, data_stage_2__587_, data_stage_2__586_, data_stage_2__585_, data_stage_2__584_, data_stage_2__583_, data_stage_2__582_, data_stage_2__581_, data_stage_2__580_, data_stage_2__579_, data_stage_2__578_, data_stage_2__577_, data_stage_2__576_, data_stage_2__575_, data_stage_2__574_, data_stage_2__573_, data_stage_2__572_, data_stage_2__571_, data_stage_2__570_, data_stage_2__569_, data_stage_2__568_, data_stage_2__567_, data_stage_2__566_, data_stage_2__565_, data_stage_2__564_, data_stage_2__563_, data_stage_2__562_, data_stage_2__561_, data_stage_2__560_, data_stage_2__559_, data_stage_2__558_, data_stage_2__557_, data_stage_2__556_, data_stage_2__555_, data_stage_2__554_, data_stage_2__553_, data_stage_2__552_, data_stage_2__551_, data_stage_2__550_, data_stage_2__549_, data_stage_2__548_, data_stage_2__547_, data_stage_2__546_, data_stage_2__545_, data_stage_2__544_, data_stage_2__543_, data_stage_2__542_, data_stage_2__541_, data_stage_2__540_, data_stage_2__539_, data_stage_2__538_, data_stage_2__537_, data_stage_2__536_, data_stage_2__535_, data_stage_2__534_, data_stage_2__533_, data_stage_2__532_, data_stage_2__531_, data_stage_2__530_, data_stage_2__529_, data_stage_2__528_, data_stage_2__527_, data_stage_2__526_, data_stage_2__525_, data_stage_2__524_, data_stage_2__523_, data_stage_2__522_, data_stage_2__521_, data_stage_2__520_, data_stage_2__519_, data_stage_2__518_, data_stage_2__517_, data_stage_2__516_, data_stage_2__515_, data_stage_2__514_, data_stage_2__513_, data_stage_2__512_ })
  );


  bsg_swap_width_p64
  mux_stage_1__mux_swap_5__swap_inst
  (
    .data_i({ data_stage_1__767_, data_stage_1__766_, data_stage_1__765_, data_stage_1__764_, data_stage_1__763_, data_stage_1__762_, data_stage_1__761_, data_stage_1__760_, data_stage_1__759_, data_stage_1__758_, data_stage_1__757_, data_stage_1__756_, data_stage_1__755_, data_stage_1__754_, data_stage_1__753_, data_stage_1__752_, data_stage_1__751_, data_stage_1__750_, data_stage_1__749_, data_stage_1__748_, data_stage_1__747_, data_stage_1__746_, data_stage_1__745_, data_stage_1__744_, data_stage_1__743_, data_stage_1__742_, data_stage_1__741_, data_stage_1__740_, data_stage_1__739_, data_stage_1__738_, data_stage_1__737_, data_stage_1__736_, data_stage_1__735_, data_stage_1__734_, data_stage_1__733_, data_stage_1__732_, data_stage_1__731_, data_stage_1__730_, data_stage_1__729_, data_stage_1__728_, data_stage_1__727_, data_stage_1__726_, data_stage_1__725_, data_stage_1__724_, data_stage_1__723_, data_stage_1__722_, data_stage_1__721_, data_stage_1__720_, data_stage_1__719_, data_stage_1__718_, data_stage_1__717_, data_stage_1__716_, data_stage_1__715_, data_stage_1__714_, data_stage_1__713_, data_stage_1__712_, data_stage_1__711_, data_stage_1__710_, data_stage_1__709_, data_stage_1__708_, data_stage_1__707_, data_stage_1__706_, data_stage_1__705_, data_stage_1__704_, data_stage_1__703_, data_stage_1__702_, data_stage_1__701_, data_stage_1__700_, data_stage_1__699_, data_stage_1__698_, data_stage_1__697_, data_stage_1__696_, data_stage_1__695_, data_stage_1__694_, data_stage_1__693_, data_stage_1__692_, data_stage_1__691_, data_stage_1__690_, data_stage_1__689_, data_stage_1__688_, data_stage_1__687_, data_stage_1__686_, data_stage_1__685_, data_stage_1__684_, data_stage_1__683_, data_stage_1__682_, data_stage_1__681_, data_stage_1__680_, data_stage_1__679_, data_stage_1__678_, data_stage_1__677_, data_stage_1__676_, data_stage_1__675_, data_stage_1__674_, data_stage_1__673_, data_stage_1__672_, data_stage_1__671_, data_stage_1__670_, data_stage_1__669_, data_stage_1__668_, data_stage_1__667_, data_stage_1__666_, data_stage_1__665_, data_stage_1__664_, data_stage_1__663_, data_stage_1__662_, data_stage_1__661_, data_stage_1__660_, data_stage_1__659_, data_stage_1__658_, data_stage_1__657_, data_stage_1__656_, data_stage_1__655_, data_stage_1__654_, data_stage_1__653_, data_stage_1__652_, data_stage_1__651_, data_stage_1__650_, data_stage_1__649_, data_stage_1__648_, data_stage_1__647_, data_stage_1__646_, data_stage_1__645_, data_stage_1__644_, data_stage_1__643_, data_stage_1__642_, data_stage_1__641_, data_stage_1__640_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__767_, data_stage_2__766_, data_stage_2__765_, data_stage_2__764_, data_stage_2__763_, data_stage_2__762_, data_stage_2__761_, data_stage_2__760_, data_stage_2__759_, data_stage_2__758_, data_stage_2__757_, data_stage_2__756_, data_stage_2__755_, data_stage_2__754_, data_stage_2__753_, data_stage_2__752_, data_stage_2__751_, data_stage_2__750_, data_stage_2__749_, data_stage_2__748_, data_stage_2__747_, data_stage_2__746_, data_stage_2__745_, data_stage_2__744_, data_stage_2__743_, data_stage_2__742_, data_stage_2__741_, data_stage_2__740_, data_stage_2__739_, data_stage_2__738_, data_stage_2__737_, data_stage_2__736_, data_stage_2__735_, data_stage_2__734_, data_stage_2__733_, data_stage_2__732_, data_stage_2__731_, data_stage_2__730_, data_stage_2__729_, data_stage_2__728_, data_stage_2__727_, data_stage_2__726_, data_stage_2__725_, data_stage_2__724_, data_stage_2__723_, data_stage_2__722_, data_stage_2__721_, data_stage_2__720_, data_stage_2__719_, data_stage_2__718_, data_stage_2__717_, data_stage_2__716_, data_stage_2__715_, data_stage_2__714_, data_stage_2__713_, data_stage_2__712_, data_stage_2__711_, data_stage_2__710_, data_stage_2__709_, data_stage_2__708_, data_stage_2__707_, data_stage_2__706_, data_stage_2__705_, data_stage_2__704_, data_stage_2__703_, data_stage_2__702_, data_stage_2__701_, data_stage_2__700_, data_stage_2__699_, data_stage_2__698_, data_stage_2__697_, data_stage_2__696_, data_stage_2__695_, data_stage_2__694_, data_stage_2__693_, data_stage_2__692_, data_stage_2__691_, data_stage_2__690_, data_stage_2__689_, data_stage_2__688_, data_stage_2__687_, data_stage_2__686_, data_stage_2__685_, data_stage_2__684_, data_stage_2__683_, data_stage_2__682_, data_stage_2__681_, data_stage_2__680_, data_stage_2__679_, data_stage_2__678_, data_stage_2__677_, data_stage_2__676_, data_stage_2__675_, data_stage_2__674_, data_stage_2__673_, data_stage_2__672_, data_stage_2__671_, data_stage_2__670_, data_stage_2__669_, data_stage_2__668_, data_stage_2__667_, data_stage_2__666_, data_stage_2__665_, data_stage_2__664_, data_stage_2__663_, data_stage_2__662_, data_stage_2__661_, data_stage_2__660_, data_stage_2__659_, data_stage_2__658_, data_stage_2__657_, data_stage_2__656_, data_stage_2__655_, data_stage_2__654_, data_stage_2__653_, data_stage_2__652_, data_stage_2__651_, data_stage_2__650_, data_stage_2__649_, data_stage_2__648_, data_stage_2__647_, data_stage_2__646_, data_stage_2__645_, data_stage_2__644_, data_stage_2__643_, data_stage_2__642_, data_stage_2__641_, data_stage_2__640_ })
  );


  bsg_swap_width_p64
  mux_stage_1__mux_swap_6__swap_inst
  (
    .data_i({ data_stage_1__895_, data_stage_1__894_, data_stage_1__893_, data_stage_1__892_, data_stage_1__891_, data_stage_1__890_, data_stage_1__889_, data_stage_1__888_, data_stage_1__887_, data_stage_1__886_, data_stage_1__885_, data_stage_1__884_, data_stage_1__883_, data_stage_1__882_, data_stage_1__881_, data_stage_1__880_, data_stage_1__879_, data_stage_1__878_, data_stage_1__877_, data_stage_1__876_, data_stage_1__875_, data_stage_1__874_, data_stage_1__873_, data_stage_1__872_, data_stage_1__871_, data_stage_1__870_, data_stage_1__869_, data_stage_1__868_, data_stage_1__867_, data_stage_1__866_, data_stage_1__865_, data_stage_1__864_, data_stage_1__863_, data_stage_1__862_, data_stage_1__861_, data_stage_1__860_, data_stage_1__859_, data_stage_1__858_, data_stage_1__857_, data_stage_1__856_, data_stage_1__855_, data_stage_1__854_, data_stage_1__853_, data_stage_1__852_, data_stage_1__851_, data_stage_1__850_, data_stage_1__849_, data_stage_1__848_, data_stage_1__847_, data_stage_1__846_, data_stage_1__845_, data_stage_1__844_, data_stage_1__843_, data_stage_1__842_, data_stage_1__841_, data_stage_1__840_, data_stage_1__839_, data_stage_1__838_, data_stage_1__837_, data_stage_1__836_, data_stage_1__835_, data_stage_1__834_, data_stage_1__833_, data_stage_1__832_, data_stage_1__831_, data_stage_1__830_, data_stage_1__829_, data_stage_1__828_, data_stage_1__827_, data_stage_1__826_, data_stage_1__825_, data_stage_1__824_, data_stage_1__823_, data_stage_1__822_, data_stage_1__821_, data_stage_1__820_, data_stage_1__819_, data_stage_1__818_, data_stage_1__817_, data_stage_1__816_, data_stage_1__815_, data_stage_1__814_, data_stage_1__813_, data_stage_1__812_, data_stage_1__811_, data_stage_1__810_, data_stage_1__809_, data_stage_1__808_, data_stage_1__807_, data_stage_1__806_, data_stage_1__805_, data_stage_1__804_, data_stage_1__803_, data_stage_1__802_, data_stage_1__801_, data_stage_1__800_, data_stage_1__799_, data_stage_1__798_, data_stage_1__797_, data_stage_1__796_, data_stage_1__795_, data_stage_1__794_, data_stage_1__793_, data_stage_1__792_, data_stage_1__791_, data_stage_1__790_, data_stage_1__789_, data_stage_1__788_, data_stage_1__787_, data_stage_1__786_, data_stage_1__785_, data_stage_1__784_, data_stage_1__783_, data_stage_1__782_, data_stage_1__781_, data_stage_1__780_, data_stage_1__779_, data_stage_1__778_, data_stage_1__777_, data_stage_1__776_, data_stage_1__775_, data_stage_1__774_, data_stage_1__773_, data_stage_1__772_, data_stage_1__771_, data_stage_1__770_, data_stage_1__769_, data_stage_1__768_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__895_, data_stage_2__894_, data_stage_2__893_, data_stage_2__892_, data_stage_2__891_, data_stage_2__890_, data_stage_2__889_, data_stage_2__888_, data_stage_2__887_, data_stage_2__886_, data_stage_2__885_, data_stage_2__884_, data_stage_2__883_, data_stage_2__882_, data_stage_2__881_, data_stage_2__880_, data_stage_2__879_, data_stage_2__878_, data_stage_2__877_, data_stage_2__876_, data_stage_2__875_, data_stage_2__874_, data_stage_2__873_, data_stage_2__872_, data_stage_2__871_, data_stage_2__870_, data_stage_2__869_, data_stage_2__868_, data_stage_2__867_, data_stage_2__866_, data_stage_2__865_, data_stage_2__864_, data_stage_2__863_, data_stage_2__862_, data_stage_2__861_, data_stage_2__860_, data_stage_2__859_, data_stage_2__858_, data_stage_2__857_, data_stage_2__856_, data_stage_2__855_, data_stage_2__854_, data_stage_2__853_, data_stage_2__852_, data_stage_2__851_, data_stage_2__850_, data_stage_2__849_, data_stage_2__848_, data_stage_2__847_, data_stage_2__846_, data_stage_2__845_, data_stage_2__844_, data_stage_2__843_, data_stage_2__842_, data_stage_2__841_, data_stage_2__840_, data_stage_2__839_, data_stage_2__838_, data_stage_2__837_, data_stage_2__836_, data_stage_2__835_, data_stage_2__834_, data_stage_2__833_, data_stage_2__832_, data_stage_2__831_, data_stage_2__830_, data_stage_2__829_, data_stage_2__828_, data_stage_2__827_, data_stage_2__826_, data_stage_2__825_, data_stage_2__824_, data_stage_2__823_, data_stage_2__822_, data_stage_2__821_, data_stage_2__820_, data_stage_2__819_, data_stage_2__818_, data_stage_2__817_, data_stage_2__816_, data_stage_2__815_, data_stage_2__814_, data_stage_2__813_, data_stage_2__812_, data_stage_2__811_, data_stage_2__810_, data_stage_2__809_, data_stage_2__808_, data_stage_2__807_, data_stage_2__806_, data_stage_2__805_, data_stage_2__804_, data_stage_2__803_, data_stage_2__802_, data_stage_2__801_, data_stage_2__800_, data_stage_2__799_, data_stage_2__798_, data_stage_2__797_, data_stage_2__796_, data_stage_2__795_, data_stage_2__794_, data_stage_2__793_, data_stage_2__792_, data_stage_2__791_, data_stage_2__790_, data_stage_2__789_, data_stage_2__788_, data_stage_2__787_, data_stage_2__786_, data_stage_2__785_, data_stage_2__784_, data_stage_2__783_, data_stage_2__782_, data_stage_2__781_, data_stage_2__780_, data_stage_2__779_, data_stage_2__778_, data_stage_2__777_, data_stage_2__776_, data_stage_2__775_, data_stage_2__774_, data_stage_2__773_, data_stage_2__772_, data_stage_2__771_, data_stage_2__770_, data_stage_2__769_, data_stage_2__768_ })
  );


  bsg_swap_width_p64
  mux_stage_1__mux_swap_7__swap_inst
  (
    .data_i({ data_stage_1__1023_, data_stage_1__1022_, data_stage_1__1021_, data_stage_1__1020_, data_stage_1__1019_, data_stage_1__1018_, data_stage_1__1017_, data_stage_1__1016_, data_stage_1__1015_, data_stage_1__1014_, data_stage_1__1013_, data_stage_1__1012_, data_stage_1__1011_, data_stage_1__1010_, data_stage_1__1009_, data_stage_1__1008_, data_stage_1__1007_, data_stage_1__1006_, data_stage_1__1005_, data_stage_1__1004_, data_stage_1__1003_, data_stage_1__1002_, data_stage_1__1001_, data_stage_1__1000_, data_stage_1__999_, data_stage_1__998_, data_stage_1__997_, data_stage_1__996_, data_stage_1__995_, data_stage_1__994_, data_stage_1__993_, data_stage_1__992_, data_stage_1__991_, data_stage_1__990_, data_stage_1__989_, data_stage_1__988_, data_stage_1__987_, data_stage_1__986_, data_stage_1__985_, data_stage_1__984_, data_stage_1__983_, data_stage_1__982_, data_stage_1__981_, data_stage_1__980_, data_stage_1__979_, data_stage_1__978_, data_stage_1__977_, data_stage_1__976_, data_stage_1__975_, data_stage_1__974_, data_stage_1__973_, data_stage_1__972_, data_stage_1__971_, data_stage_1__970_, data_stage_1__969_, data_stage_1__968_, data_stage_1__967_, data_stage_1__966_, data_stage_1__965_, data_stage_1__964_, data_stage_1__963_, data_stage_1__962_, data_stage_1__961_, data_stage_1__960_, data_stage_1__959_, data_stage_1__958_, data_stage_1__957_, data_stage_1__956_, data_stage_1__955_, data_stage_1__954_, data_stage_1__953_, data_stage_1__952_, data_stage_1__951_, data_stage_1__950_, data_stage_1__949_, data_stage_1__948_, data_stage_1__947_, data_stage_1__946_, data_stage_1__945_, data_stage_1__944_, data_stage_1__943_, data_stage_1__942_, data_stage_1__941_, data_stage_1__940_, data_stage_1__939_, data_stage_1__938_, data_stage_1__937_, data_stage_1__936_, data_stage_1__935_, data_stage_1__934_, data_stage_1__933_, data_stage_1__932_, data_stage_1__931_, data_stage_1__930_, data_stage_1__929_, data_stage_1__928_, data_stage_1__927_, data_stage_1__926_, data_stage_1__925_, data_stage_1__924_, data_stage_1__923_, data_stage_1__922_, data_stage_1__921_, data_stage_1__920_, data_stage_1__919_, data_stage_1__918_, data_stage_1__917_, data_stage_1__916_, data_stage_1__915_, data_stage_1__914_, data_stage_1__913_, data_stage_1__912_, data_stage_1__911_, data_stage_1__910_, data_stage_1__909_, data_stage_1__908_, data_stage_1__907_, data_stage_1__906_, data_stage_1__905_, data_stage_1__904_, data_stage_1__903_, data_stage_1__902_, data_stage_1__901_, data_stage_1__900_, data_stage_1__899_, data_stage_1__898_, data_stage_1__897_, data_stage_1__896_ }),
    .swap_i(sel_i[1]),
    .data_o({ data_stage_2__1023_, data_stage_2__1022_, data_stage_2__1021_, data_stage_2__1020_, data_stage_2__1019_, data_stage_2__1018_, data_stage_2__1017_, data_stage_2__1016_, data_stage_2__1015_, data_stage_2__1014_, data_stage_2__1013_, data_stage_2__1012_, data_stage_2__1011_, data_stage_2__1010_, data_stage_2__1009_, data_stage_2__1008_, data_stage_2__1007_, data_stage_2__1006_, data_stage_2__1005_, data_stage_2__1004_, data_stage_2__1003_, data_stage_2__1002_, data_stage_2__1001_, data_stage_2__1000_, data_stage_2__999_, data_stage_2__998_, data_stage_2__997_, data_stage_2__996_, data_stage_2__995_, data_stage_2__994_, data_stage_2__993_, data_stage_2__992_, data_stage_2__991_, data_stage_2__990_, data_stage_2__989_, data_stage_2__988_, data_stage_2__987_, data_stage_2__986_, data_stage_2__985_, data_stage_2__984_, data_stage_2__983_, data_stage_2__982_, data_stage_2__981_, data_stage_2__980_, data_stage_2__979_, data_stage_2__978_, data_stage_2__977_, data_stage_2__976_, data_stage_2__975_, data_stage_2__974_, data_stage_2__973_, data_stage_2__972_, data_stage_2__971_, data_stage_2__970_, data_stage_2__969_, data_stage_2__968_, data_stage_2__967_, data_stage_2__966_, data_stage_2__965_, data_stage_2__964_, data_stage_2__963_, data_stage_2__962_, data_stage_2__961_, data_stage_2__960_, data_stage_2__959_, data_stage_2__958_, data_stage_2__957_, data_stage_2__956_, data_stage_2__955_, data_stage_2__954_, data_stage_2__953_, data_stage_2__952_, data_stage_2__951_, data_stage_2__950_, data_stage_2__949_, data_stage_2__948_, data_stage_2__947_, data_stage_2__946_, data_stage_2__945_, data_stage_2__944_, data_stage_2__943_, data_stage_2__942_, data_stage_2__941_, data_stage_2__940_, data_stage_2__939_, data_stage_2__938_, data_stage_2__937_, data_stage_2__936_, data_stage_2__935_, data_stage_2__934_, data_stage_2__933_, data_stage_2__932_, data_stage_2__931_, data_stage_2__930_, data_stage_2__929_, data_stage_2__928_, data_stage_2__927_, data_stage_2__926_, data_stage_2__925_, data_stage_2__924_, data_stage_2__923_, data_stage_2__922_, data_stage_2__921_, data_stage_2__920_, data_stage_2__919_, data_stage_2__918_, data_stage_2__917_, data_stage_2__916_, data_stage_2__915_, data_stage_2__914_, data_stage_2__913_, data_stage_2__912_, data_stage_2__911_, data_stage_2__910_, data_stage_2__909_, data_stage_2__908_, data_stage_2__907_, data_stage_2__906_, data_stage_2__905_, data_stage_2__904_, data_stage_2__903_, data_stage_2__902_, data_stage_2__901_, data_stage_2__900_, data_stage_2__899_, data_stage_2__898_, data_stage_2__897_, data_stage_2__896_ })
  );


  bsg_swap_width_p128
  mux_stage_2__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_2__255_, data_stage_2__254_, data_stage_2__253_, data_stage_2__252_, data_stage_2__251_, data_stage_2__250_, data_stage_2__249_, data_stage_2__248_, data_stage_2__247_, data_stage_2__246_, data_stage_2__245_, data_stage_2__244_, data_stage_2__243_, data_stage_2__242_, data_stage_2__241_, data_stage_2__240_, data_stage_2__239_, data_stage_2__238_, data_stage_2__237_, data_stage_2__236_, data_stage_2__235_, data_stage_2__234_, data_stage_2__233_, data_stage_2__232_, data_stage_2__231_, data_stage_2__230_, data_stage_2__229_, data_stage_2__228_, data_stage_2__227_, data_stage_2__226_, data_stage_2__225_, data_stage_2__224_, data_stage_2__223_, data_stage_2__222_, data_stage_2__221_, data_stage_2__220_, data_stage_2__219_, data_stage_2__218_, data_stage_2__217_, data_stage_2__216_, data_stage_2__215_, data_stage_2__214_, data_stage_2__213_, data_stage_2__212_, data_stage_2__211_, data_stage_2__210_, data_stage_2__209_, data_stage_2__208_, data_stage_2__207_, data_stage_2__206_, data_stage_2__205_, data_stage_2__204_, data_stage_2__203_, data_stage_2__202_, data_stage_2__201_, data_stage_2__200_, data_stage_2__199_, data_stage_2__198_, data_stage_2__197_, data_stage_2__196_, data_stage_2__195_, data_stage_2__194_, data_stage_2__193_, data_stage_2__192_, data_stage_2__191_, data_stage_2__190_, data_stage_2__189_, data_stage_2__188_, data_stage_2__187_, data_stage_2__186_, data_stage_2__185_, data_stage_2__184_, data_stage_2__183_, data_stage_2__182_, data_stage_2__181_, data_stage_2__180_, data_stage_2__179_, data_stage_2__178_, data_stage_2__177_, data_stage_2__176_, data_stage_2__175_, data_stage_2__174_, data_stage_2__173_, data_stage_2__172_, data_stage_2__171_, data_stage_2__170_, data_stage_2__169_, data_stage_2__168_, data_stage_2__167_, data_stage_2__166_, data_stage_2__165_, data_stage_2__164_, data_stage_2__163_, data_stage_2__162_, data_stage_2__161_, data_stage_2__160_, data_stage_2__159_, data_stage_2__158_, data_stage_2__157_, data_stage_2__156_, data_stage_2__155_, data_stage_2__154_, data_stage_2__153_, data_stage_2__152_, data_stage_2__151_, data_stage_2__150_, data_stage_2__149_, data_stage_2__148_, data_stage_2__147_, data_stage_2__146_, data_stage_2__145_, data_stage_2__144_, data_stage_2__143_, data_stage_2__142_, data_stage_2__141_, data_stage_2__140_, data_stage_2__139_, data_stage_2__138_, data_stage_2__137_, data_stage_2__136_, data_stage_2__135_, data_stage_2__134_, data_stage_2__133_, data_stage_2__132_, data_stage_2__131_, data_stage_2__130_, data_stage_2__129_, data_stage_2__128_, data_stage_2__127_, data_stage_2__126_, data_stage_2__125_, data_stage_2__124_, data_stage_2__123_, data_stage_2__122_, data_stage_2__121_, data_stage_2__120_, data_stage_2__119_, data_stage_2__118_, data_stage_2__117_, data_stage_2__116_, data_stage_2__115_, data_stage_2__114_, data_stage_2__113_, data_stage_2__112_, data_stage_2__111_, data_stage_2__110_, data_stage_2__109_, data_stage_2__108_, data_stage_2__107_, data_stage_2__106_, data_stage_2__105_, data_stage_2__104_, data_stage_2__103_, data_stage_2__102_, data_stage_2__101_, data_stage_2__100_, data_stage_2__99_, data_stage_2__98_, data_stage_2__97_, data_stage_2__96_, data_stage_2__95_, data_stage_2__94_, data_stage_2__93_, data_stage_2__92_, data_stage_2__91_, data_stage_2__90_, data_stage_2__89_, data_stage_2__88_, data_stage_2__87_, data_stage_2__86_, data_stage_2__85_, data_stage_2__84_, data_stage_2__83_, data_stage_2__82_, data_stage_2__81_, data_stage_2__80_, data_stage_2__79_, data_stage_2__78_, data_stage_2__77_, data_stage_2__76_, data_stage_2__75_, data_stage_2__74_, data_stage_2__73_, data_stage_2__72_, data_stage_2__71_, data_stage_2__70_, data_stage_2__69_, data_stage_2__68_, data_stage_2__67_, data_stage_2__66_, data_stage_2__65_, data_stage_2__64_, data_stage_2__63_, data_stage_2__62_, data_stage_2__61_, data_stage_2__60_, data_stage_2__59_, data_stage_2__58_, data_stage_2__57_, data_stage_2__56_, data_stage_2__55_, data_stage_2__54_, data_stage_2__53_, data_stage_2__52_, data_stage_2__51_, data_stage_2__50_, data_stage_2__49_, data_stage_2__48_, data_stage_2__47_, data_stage_2__46_, data_stage_2__45_, data_stage_2__44_, data_stage_2__43_, data_stage_2__42_, data_stage_2__41_, data_stage_2__40_, data_stage_2__39_, data_stage_2__38_, data_stage_2__37_, data_stage_2__36_, data_stage_2__35_, data_stage_2__34_, data_stage_2__33_, data_stage_2__32_, data_stage_2__31_, data_stage_2__30_, data_stage_2__29_, data_stage_2__28_, data_stage_2__27_, data_stage_2__26_, data_stage_2__25_, data_stage_2__24_, data_stage_2__23_, data_stage_2__22_, data_stage_2__21_, data_stage_2__20_, data_stage_2__19_, data_stage_2__18_, data_stage_2__17_, data_stage_2__16_, data_stage_2__15_, data_stage_2__14_, data_stage_2__13_, data_stage_2__12_, data_stage_2__11_, data_stage_2__10_, data_stage_2__9_, data_stage_2__8_, data_stage_2__7_, data_stage_2__6_, data_stage_2__5_, data_stage_2__4_, data_stage_2__3_, data_stage_2__2_, data_stage_2__1_, data_stage_2__0_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__255_, data_stage_3__254_, data_stage_3__253_, data_stage_3__252_, data_stage_3__251_, data_stage_3__250_, data_stage_3__249_, data_stage_3__248_, data_stage_3__247_, data_stage_3__246_, data_stage_3__245_, data_stage_3__244_, data_stage_3__243_, data_stage_3__242_, data_stage_3__241_, data_stage_3__240_, data_stage_3__239_, data_stage_3__238_, data_stage_3__237_, data_stage_3__236_, data_stage_3__235_, data_stage_3__234_, data_stage_3__233_, data_stage_3__232_, data_stage_3__231_, data_stage_3__230_, data_stage_3__229_, data_stage_3__228_, data_stage_3__227_, data_stage_3__226_, data_stage_3__225_, data_stage_3__224_, data_stage_3__223_, data_stage_3__222_, data_stage_3__221_, data_stage_3__220_, data_stage_3__219_, data_stage_3__218_, data_stage_3__217_, data_stage_3__216_, data_stage_3__215_, data_stage_3__214_, data_stage_3__213_, data_stage_3__212_, data_stage_3__211_, data_stage_3__210_, data_stage_3__209_, data_stage_3__208_, data_stage_3__207_, data_stage_3__206_, data_stage_3__205_, data_stage_3__204_, data_stage_3__203_, data_stage_3__202_, data_stage_3__201_, data_stage_3__200_, data_stage_3__199_, data_stage_3__198_, data_stage_3__197_, data_stage_3__196_, data_stage_3__195_, data_stage_3__194_, data_stage_3__193_, data_stage_3__192_, data_stage_3__191_, data_stage_3__190_, data_stage_3__189_, data_stage_3__188_, data_stage_3__187_, data_stage_3__186_, data_stage_3__185_, data_stage_3__184_, data_stage_3__183_, data_stage_3__182_, data_stage_3__181_, data_stage_3__180_, data_stage_3__179_, data_stage_3__178_, data_stage_3__177_, data_stage_3__176_, data_stage_3__175_, data_stage_3__174_, data_stage_3__173_, data_stage_3__172_, data_stage_3__171_, data_stage_3__170_, data_stage_3__169_, data_stage_3__168_, data_stage_3__167_, data_stage_3__166_, data_stage_3__165_, data_stage_3__164_, data_stage_3__163_, data_stage_3__162_, data_stage_3__161_, data_stage_3__160_, data_stage_3__159_, data_stage_3__158_, data_stage_3__157_, data_stage_3__156_, data_stage_3__155_, data_stage_3__154_, data_stage_3__153_, data_stage_3__152_, data_stage_3__151_, data_stage_3__150_, data_stage_3__149_, data_stage_3__148_, data_stage_3__147_, data_stage_3__146_, data_stage_3__145_, data_stage_3__144_, data_stage_3__143_, data_stage_3__142_, data_stage_3__141_, data_stage_3__140_, data_stage_3__139_, data_stage_3__138_, data_stage_3__137_, data_stage_3__136_, data_stage_3__135_, data_stage_3__134_, data_stage_3__133_, data_stage_3__132_, data_stage_3__131_, data_stage_3__130_, data_stage_3__129_, data_stage_3__128_, data_stage_3__127_, data_stage_3__126_, data_stage_3__125_, data_stage_3__124_, data_stage_3__123_, data_stage_3__122_, data_stage_3__121_, data_stage_3__120_, data_stage_3__119_, data_stage_3__118_, data_stage_3__117_, data_stage_3__116_, data_stage_3__115_, data_stage_3__114_, data_stage_3__113_, data_stage_3__112_, data_stage_3__111_, data_stage_3__110_, data_stage_3__109_, data_stage_3__108_, data_stage_3__107_, data_stage_3__106_, data_stage_3__105_, data_stage_3__104_, data_stage_3__103_, data_stage_3__102_, data_stage_3__101_, data_stage_3__100_, data_stage_3__99_, data_stage_3__98_, data_stage_3__97_, data_stage_3__96_, data_stage_3__95_, data_stage_3__94_, data_stage_3__93_, data_stage_3__92_, data_stage_3__91_, data_stage_3__90_, data_stage_3__89_, data_stage_3__88_, data_stage_3__87_, data_stage_3__86_, data_stage_3__85_, data_stage_3__84_, data_stage_3__83_, data_stage_3__82_, data_stage_3__81_, data_stage_3__80_, data_stage_3__79_, data_stage_3__78_, data_stage_3__77_, data_stage_3__76_, data_stage_3__75_, data_stage_3__74_, data_stage_3__73_, data_stage_3__72_, data_stage_3__71_, data_stage_3__70_, data_stage_3__69_, data_stage_3__68_, data_stage_3__67_, data_stage_3__66_, data_stage_3__65_, data_stage_3__64_, data_stage_3__63_, data_stage_3__62_, data_stage_3__61_, data_stage_3__60_, data_stage_3__59_, data_stage_3__58_, data_stage_3__57_, data_stage_3__56_, data_stage_3__55_, data_stage_3__54_, data_stage_3__53_, data_stage_3__52_, data_stage_3__51_, data_stage_3__50_, data_stage_3__49_, data_stage_3__48_, data_stage_3__47_, data_stage_3__46_, data_stage_3__45_, data_stage_3__44_, data_stage_3__43_, data_stage_3__42_, data_stage_3__41_, data_stage_3__40_, data_stage_3__39_, data_stage_3__38_, data_stage_3__37_, data_stage_3__36_, data_stage_3__35_, data_stage_3__34_, data_stage_3__33_, data_stage_3__32_, data_stage_3__31_, data_stage_3__30_, data_stage_3__29_, data_stage_3__28_, data_stage_3__27_, data_stage_3__26_, data_stage_3__25_, data_stage_3__24_, data_stage_3__23_, data_stage_3__22_, data_stage_3__21_, data_stage_3__20_, data_stage_3__19_, data_stage_3__18_, data_stage_3__17_, data_stage_3__16_, data_stage_3__15_, data_stage_3__14_, data_stage_3__13_, data_stage_3__12_, data_stage_3__11_, data_stage_3__10_, data_stage_3__9_, data_stage_3__8_, data_stage_3__7_, data_stage_3__6_, data_stage_3__5_, data_stage_3__4_, data_stage_3__3_, data_stage_3__2_, data_stage_3__1_, data_stage_3__0_ })
  );


  bsg_swap_width_p128
  mux_stage_2__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_2__511_, data_stage_2__510_, data_stage_2__509_, data_stage_2__508_, data_stage_2__507_, data_stage_2__506_, data_stage_2__505_, data_stage_2__504_, data_stage_2__503_, data_stage_2__502_, data_stage_2__501_, data_stage_2__500_, data_stage_2__499_, data_stage_2__498_, data_stage_2__497_, data_stage_2__496_, data_stage_2__495_, data_stage_2__494_, data_stage_2__493_, data_stage_2__492_, data_stage_2__491_, data_stage_2__490_, data_stage_2__489_, data_stage_2__488_, data_stage_2__487_, data_stage_2__486_, data_stage_2__485_, data_stage_2__484_, data_stage_2__483_, data_stage_2__482_, data_stage_2__481_, data_stage_2__480_, data_stage_2__479_, data_stage_2__478_, data_stage_2__477_, data_stage_2__476_, data_stage_2__475_, data_stage_2__474_, data_stage_2__473_, data_stage_2__472_, data_stage_2__471_, data_stage_2__470_, data_stage_2__469_, data_stage_2__468_, data_stage_2__467_, data_stage_2__466_, data_stage_2__465_, data_stage_2__464_, data_stage_2__463_, data_stage_2__462_, data_stage_2__461_, data_stage_2__460_, data_stage_2__459_, data_stage_2__458_, data_stage_2__457_, data_stage_2__456_, data_stage_2__455_, data_stage_2__454_, data_stage_2__453_, data_stage_2__452_, data_stage_2__451_, data_stage_2__450_, data_stage_2__449_, data_stage_2__448_, data_stage_2__447_, data_stage_2__446_, data_stage_2__445_, data_stage_2__444_, data_stage_2__443_, data_stage_2__442_, data_stage_2__441_, data_stage_2__440_, data_stage_2__439_, data_stage_2__438_, data_stage_2__437_, data_stage_2__436_, data_stage_2__435_, data_stage_2__434_, data_stage_2__433_, data_stage_2__432_, data_stage_2__431_, data_stage_2__430_, data_stage_2__429_, data_stage_2__428_, data_stage_2__427_, data_stage_2__426_, data_stage_2__425_, data_stage_2__424_, data_stage_2__423_, data_stage_2__422_, data_stage_2__421_, data_stage_2__420_, data_stage_2__419_, data_stage_2__418_, data_stage_2__417_, data_stage_2__416_, data_stage_2__415_, data_stage_2__414_, data_stage_2__413_, data_stage_2__412_, data_stage_2__411_, data_stage_2__410_, data_stage_2__409_, data_stage_2__408_, data_stage_2__407_, data_stage_2__406_, data_stage_2__405_, data_stage_2__404_, data_stage_2__403_, data_stage_2__402_, data_stage_2__401_, data_stage_2__400_, data_stage_2__399_, data_stage_2__398_, data_stage_2__397_, data_stage_2__396_, data_stage_2__395_, data_stage_2__394_, data_stage_2__393_, data_stage_2__392_, data_stage_2__391_, data_stage_2__390_, data_stage_2__389_, data_stage_2__388_, data_stage_2__387_, data_stage_2__386_, data_stage_2__385_, data_stage_2__384_, data_stage_2__383_, data_stage_2__382_, data_stage_2__381_, data_stage_2__380_, data_stage_2__379_, data_stage_2__378_, data_stage_2__377_, data_stage_2__376_, data_stage_2__375_, data_stage_2__374_, data_stage_2__373_, data_stage_2__372_, data_stage_2__371_, data_stage_2__370_, data_stage_2__369_, data_stage_2__368_, data_stage_2__367_, data_stage_2__366_, data_stage_2__365_, data_stage_2__364_, data_stage_2__363_, data_stage_2__362_, data_stage_2__361_, data_stage_2__360_, data_stage_2__359_, data_stage_2__358_, data_stage_2__357_, data_stage_2__356_, data_stage_2__355_, data_stage_2__354_, data_stage_2__353_, data_stage_2__352_, data_stage_2__351_, data_stage_2__350_, data_stage_2__349_, data_stage_2__348_, data_stage_2__347_, data_stage_2__346_, data_stage_2__345_, data_stage_2__344_, data_stage_2__343_, data_stage_2__342_, data_stage_2__341_, data_stage_2__340_, data_stage_2__339_, data_stage_2__338_, data_stage_2__337_, data_stage_2__336_, data_stage_2__335_, data_stage_2__334_, data_stage_2__333_, data_stage_2__332_, data_stage_2__331_, data_stage_2__330_, data_stage_2__329_, data_stage_2__328_, data_stage_2__327_, data_stage_2__326_, data_stage_2__325_, data_stage_2__324_, data_stage_2__323_, data_stage_2__322_, data_stage_2__321_, data_stage_2__320_, data_stage_2__319_, data_stage_2__318_, data_stage_2__317_, data_stage_2__316_, data_stage_2__315_, data_stage_2__314_, data_stage_2__313_, data_stage_2__312_, data_stage_2__311_, data_stage_2__310_, data_stage_2__309_, data_stage_2__308_, data_stage_2__307_, data_stage_2__306_, data_stage_2__305_, data_stage_2__304_, data_stage_2__303_, data_stage_2__302_, data_stage_2__301_, data_stage_2__300_, data_stage_2__299_, data_stage_2__298_, data_stage_2__297_, data_stage_2__296_, data_stage_2__295_, data_stage_2__294_, data_stage_2__293_, data_stage_2__292_, data_stage_2__291_, data_stage_2__290_, data_stage_2__289_, data_stage_2__288_, data_stage_2__287_, data_stage_2__286_, data_stage_2__285_, data_stage_2__284_, data_stage_2__283_, data_stage_2__282_, data_stage_2__281_, data_stage_2__280_, data_stage_2__279_, data_stage_2__278_, data_stage_2__277_, data_stage_2__276_, data_stage_2__275_, data_stage_2__274_, data_stage_2__273_, data_stage_2__272_, data_stage_2__271_, data_stage_2__270_, data_stage_2__269_, data_stage_2__268_, data_stage_2__267_, data_stage_2__266_, data_stage_2__265_, data_stage_2__264_, data_stage_2__263_, data_stage_2__262_, data_stage_2__261_, data_stage_2__260_, data_stage_2__259_, data_stage_2__258_, data_stage_2__257_, data_stage_2__256_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__511_, data_stage_3__510_, data_stage_3__509_, data_stage_3__508_, data_stage_3__507_, data_stage_3__506_, data_stage_3__505_, data_stage_3__504_, data_stage_3__503_, data_stage_3__502_, data_stage_3__501_, data_stage_3__500_, data_stage_3__499_, data_stage_3__498_, data_stage_3__497_, data_stage_3__496_, data_stage_3__495_, data_stage_3__494_, data_stage_3__493_, data_stage_3__492_, data_stage_3__491_, data_stage_3__490_, data_stage_3__489_, data_stage_3__488_, data_stage_3__487_, data_stage_3__486_, data_stage_3__485_, data_stage_3__484_, data_stage_3__483_, data_stage_3__482_, data_stage_3__481_, data_stage_3__480_, data_stage_3__479_, data_stage_3__478_, data_stage_3__477_, data_stage_3__476_, data_stage_3__475_, data_stage_3__474_, data_stage_3__473_, data_stage_3__472_, data_stage_3__471_, data_stage_3__470_, data_stage_3__469_, data_stage_3__468_, data_stage_3__467_, data_stage_3__466_, data_stage_3__465_, data_stage_3__464_, data_stage_3__463_, data_stage_3__462_, data_stage_3__461_, data_stage_3__460_, data_stage_3__459_, data_stage_3__458_, data_stage_3__457_, data_stage_3__456_, data_stage_3__455_, data_stage_3__454_, data_stage_3__453_, data_stage_3__452_, data_stage_3__451_, data_stage_3__450_, data_stage_3__449_, data_stage_3__448_, data_stage_3__447_, data_stage_3__446_, data_stage_3__445_, data_stage_3__444_, data_stage_3__443_, data_stage_3__442_, data_stage_3__441_, data_stage_3__440_, data_stage_3__439_, data_stage_3__438_, data_stage_3__437_, data_stage_3__436_, data_stage_3__435_, data_stage_3__434_, data_stage_3__433_, data_stage_3__432_, data_stage_3__431_, data_stage_3__430_, data_stage_3__429_, data_stage_3__428_, data_stage_3__427_, data_stage_3__426_, data_stage_3__425_, data_stage_3__424_, data_stage_3__423_, data_stage_3__422_, data_stage_3__421_, data_stage_3__420_, data_stage_3__419_, data_stage_3__418_, data_stage_3__417_, data_stage_3__416_, data_stage_3__415_, data_stage_3__414_, data_stage_3__413_, data_stage_3__412_, data_stage_3__411_, data_stage_3__410_, data_stage_3__409_, data_stage_3__408_, data_stage_3__407_, data_stage_3__406_, data_stage_3__405_, data_stage_3__404_, data_stage_3__403_, data_stage_3__402_, data_stage_3__401_, data_stage_3__400_, data_stage_3__399_, data_stage_3__398_, data_stage_3__397_, data_stage_3__396_, data_stage_3__395_, data_stage_3__394_, data_stage_3__393_, data_stage_3__392_, data_stage_3__391_, data_stage_3__390_, data_stage_3__389_, data_stage_3__388_, data_stage_3__387_, data_stage_3__386_, data_stage_3__385_, data_stage_3__384_, data_stage_3__383_, data_stage_3__382_, data_stage_3__381_, data_stage_3__380_, data_stage_3__379_, data_stage_3__378_, data_stage_3__377_, data_stage_3__376_, data_stage_3__375_, data_stage_3__374_, data_stage_3__373_, data_stage_3__372_, data_stage_3__371_, data_stage_3__370_, data_stage_3__369_, data_stage_3__368_, data_stage_3__367_, data_stage_3__366_, data_stage_3__365_, data_stage_3__364_, data_stage_3__363_, data_stage_3__362_, data_stage_3__361_, data_stage_3__360_, data_stage_3__359_, data_stage_3__358_, data_stage_3__357_, data_stage_3__356_, data_stage_3__355_, data_stage_3__354_, data_stage_3__353_, data_stage_3__352_, data_stage_3__351_, data_stage_3__350_, data_stage_3__349_, data_stage_3__348_, data_stage_3__347_, data_stage_3__346_, data_stage_3__345_, data_stage_3__344_, data_stage_3__343_, data_stage_3__342_, data_stage_3__341_, data_stage_3__340_, data_stage_3__339_, data_stage_3__338_, data_stage_3__337_, data_stage_3__336_, data_stage_3__335_, data_stage_3__334_, data_stage_3__333_, data_stage_3__332_, data_stage_3__331_, data_stage_3__330_, data_stage_3__329_, data_stage_3__328_, data_stage_3__327_, data_stage_3__326_, data_stage_3__325_, data_stage_3__324_, data_stage_3__323_, data_stage_3__322_, data_stage_3__321_, data_stage_3__320_, data_stage_3__319_, data_stage_3__318_, data_stage_3__317_, data_stage_3__316_, data_stage_3__315_, data_stage_3__314_, data_stage_3__313_, data_stage_3__312_, data_stage_3__311_, data_stage_3__310_, data_stage_3__309_, data_stage_3__308_, data_stage_3__307_, data_stage_3__306_, data_stage_3__305_, data_stage_3__304_, data_stage_3__303_, data_stage_3__302_, data_stage_3__301_, data_stage_3__300_, data_stage_3__299_, data_stage_3__298_, data_stage_3__297_, data_stage_3__296_, data_stage_3__295_, data_stage_3__294_, data_stage_3__293_, data_stage_3__292_, data_stage_3__291_, data_stage_3__290_, data_stage_3__289_, data_stage_3__288_, data_stage_3__287_, data_stage_3__286_, data_stage_3__285_, data_stage_3__284_, data_stage_3__283_, data_stage_3__282_, data_stage_3__281_, data_stage_3__280_, data_stage_3__279_, data_stage_3__278_, data_stage_3__277_, data_stage_3__276_, data_stage_3__275_, data_stage_3__274_, data_stage_3__273_, data_stage_3__272_, data_stage_3__271_, data_stage_3__270_, data_stage_3__269_, data_stage_3__268_, data_stage_3__267_, data_stage_3__266_, data_stage_3__265_, data_stage_3__264_, data_stage_3__263_, data_stage_3__262_, data_stage_3__261_, data_stage_3__260_, data_stage_3__259_, data_stage_3__258_, data_stage_3__257_, data_stage_3__256_ })
  );


  bsg_swap_width_p128
  mux_stage_2__mux_swap_2__swap_inst
  (
    .data_i({ data_stage_2__767_, data_stage_2__766_, data_stage_2__765_, data_stage_2__764_, data_stage_2__763_, data_stage_2__762_, data_stage_2__761_, data_stage_2__760_, data_stage_2__759_, data_stage_2__758_, data_stage_2__757_, data_stage_2__756_, data_stage_2__755_, data_stage_2__754_, data_stage_2__753_, data_stage_2__752_, data_stage_2__751_, data_stage_2__750_, data_stage_2__749_, data_stage_2__748_, data_stage_2__747_, data_stage_2__746_, data_stage_2__745_, data_stage_2__744_, data_stage_2__743_, data_stage_2__742_, data_stage_2__741_, data_stage_2__740_, data_stage_2__739_, data_stage_2__738_, data_stage_2__737_, data_stage_2__736_, data_stage_2__735_, data_stage_2__734_, data_stage_2__733_, data_stage_2__732_, data_stage_2__731_, data_stage_2__730_, data_stage_2__729_, data_stage_2__728_, data_stage_2__727_, data_stage_2__726_, data_stage_2__725_, data_stage_2__724_, data_stage_2__723_, data_stage_2__722_, data_stage_2__721_, data_stage_2__720_, data_stage_2__719_, data_stage_2__718_, data_stage_2__717_, data_stage_2__716_, data_stage_2__715_, data_stage_2__714_, data_stage_2__713_, data_stage_2__712_, data_stage_2__711_, data_stage_2__710_, data_stage_2__709_, data_stage_2__708_, data_stage_2__707_, data_stage_2__706_, data_stage_2__705_, data_stage_2__704_, data_stage_2__703_, data_stage_2__702_, data_stage_2__701_, data_stage_2__700_, data_stage_2__699_, data_stage_2__698_, data_stage_2__697_, data_stage_2__696_, data_stage_2__695_, data_stage_2__694_, data_stage_2__693_, data_stage_2__692_, data_stage_2__691_, data_stage_2__690_, data_stage_2__689_, data_stage_2__688_, data_stage_2__687_, data_stage_2__686_, data_stage_2__685_, data_stage_2__684_, data_stage_2__683_, data_stage_2__682_, data_stage_2__681_, data_stage_2__680_, data_stage_2__679_, data_stage_2__678_, data_stage_2__677_, data_stage_2__676_, data_stage_2__675_, data_stage_2__674_, data_stage_2__673_, data_stage_2__672_, data_stage_2__671_, data_stage_2__670_, data_stage_2__669_, data_stage_2__668_, data_stage_2__667_, data_stage_2__666_, data_stage_2__665_, data_stage_2__664_, data_stage_2__663_, data_stage_2__662_, data_stage_2__661_, data_stage_2__660_, data_stage_2__659_, data_stage_2__658_, data_stage_2__657_, data_stage_2__656_, data_stage_2__655_, data_stage_2__654_, data_stage_2__653_, data_stage_2__652_, data_stage_2__651_, data_stage_2__650_, data_stage_2__649_, data_stage_2__648_, data_stage_2__647_, data_stage_2__646_, data_stage_2__645_, data_stage_2__644_, data_stage_2__643_, data_stage_2__642_, data_stage_2__641_, data_stage_2__640_, data_stage_2__639_, data_stage_2__638_, data_stage_2__637_, data_stage_2__636_, data_stage_2__635_, data_stage_2__634_, data_stage_2__633_, data_stage_2__632_, data_stage_2__631_, data_stage_2__630_, data_stage_2__629_, data_stage_2__628_, data_stage_2__627_, data_stage_2__626_, data_stage_2__625_, data_stage_2__624_, data_stage_2__623_, data_stage_2__622_, data_stage_2__621_, data_stage_2__620_, data_stage_2__619_, data_stage_2__618_, data_stage_2__617_, data_stage_2__616_, data_stage_2__615_, data_stage_2__614_, data_stage_2__613_, data_stage_2__612_, data_stage_2__611_, data_stage_2__610_, data_stage_2__609_, data_stage_2__608_, data_stage_2__607_, data_stage_2__606_, data_stage_2__605_, data_stage_2__604_, data_stage_2__603_, data_stage_2__602_, data_stage_2__601_, data_stage_2__600_, data_stage_2__599_, data_stage_2__598_, data_stage_2__597_, data_stage_2__596_, data_stage_2__595_, data_stage_2__594_, data_stage_2__593_, data_stage_2__592_, data_stage_2__591_, data_stage_2__590_, data_stage_2__589_, data_stage_2__588_, data_stage_2__587_, data_stage_2__586_, data_stage_2__585_, data_stage_2__584_, data_stage_2__583_, data_stage_2__582_, data_stage_2__581_, data_stage_2__580_, data_stage_2__579_, data_stage_2__578_, data_stage_2__577_, data_stage_2__576_, data_stage_2__575_, data_stage_2__574_, data_stage_2__573_, data_stage_2__572_, data_stage_2__571_, data_stage_2__570_, data_stage_2__569_, data_stage_2__568_, data_stage_2__567_, data_stage_2__566_, data_stage_2__565_, data_stage_2__564_, data_stage_2__563_, data_stage_2__562_, data_stage_2__561_, data_stage_2__560_, data_stage_2__559_, data_stage_2__558_, data_stage_2__557_, data_stage_2__556_, data_stage_2__555_, data_stage_2__554_, data_stage_2__553_, data_stage_2__552_, data_stage_2__551_, data_stage_2__550_, data_stage_2__549_, data_stage_2__548_, data_stage_2__547_, data_stage_2__546_, data_stage_2__545_, data_stage_2__544_, data_stage_2__543_, data_stage_2__542_, data_stage_2__541_, data_stage_2__540_, data_stage_2__539_, data_stage_2__538_, data_stage_2__537_, data_stage_2__536_, data_stage_2__535_, data_stage_2__534_, data_stage_2__533_, data_stage_2__532_, data_stage_2__531_, data_stage_2__530_, data_stage_2__529_, data_stage_2__528_, data_stage_2__527_, data_stage_2__526_, data_stage_2__525_, data_stage_2__524_, data_stage_2__523_, data_stage_2__522_, data_stage_2__521_, data_stage_2__520_, data_stage_2__519_, data_stage_2__518_, data_stage_2__517_, data_stage_2__516_, data_stage_2__515_, data_stage_2__514_, data_stage_2__513_, data_stage_2__512_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__767_, data_stage_3__766_, data_stage_3__765_, data_stage_3__764_, data_stage_3__763_, data_stage_3__762_, data_stage_3__761_, data_stage_3__760_, data_stage_3__759_, data_stage_3__758_, data_stage_3__757_, data_stage_3__756_, data_stage_3__755_, data_stage_3__754_, data_stage_3__753_, data_stage_3__752_, data_stage_3__751_, data_stage_3__750_, data_stage_3__749_, data_stage_3__748_, data_stage_3__747_, data_stage_3__746_, data_stage_3__745_, data_stage_3__744_, data_stage_3__743_, data_stage_3__742_, data_stage_3__741_, data_stage_3__740_, data_stage_3__739_, data_stage_3__738_, data_stage_3__737_, data_stage_3__736_, data_stage_3__735_, data_stage_3__734_, data_stage_3__733_, data_stage_3__732_, data_stage_3__731_, data_stage_3__730_, data_stage_3__729_, data_stage_3__728_, data_stage_3__727_, data_stage_3__726_, data_stage_3__725_, data_stage_3__724_, data_stage_3__723_, data_stage_3__722_, data_stage_3__721_, data_stage_3__720_, data_stage_3__719_, data_stage_3__718_, data_stage_3__717_, data_stage_3__716_, data_stage_3__715_, data_stage_3__714_, data_stage_3__713_, data_stage_3__712_, data_stage_3__711_, data_stage_3__710_, data_stage_3__709_, data_stage_3__708_, data_stage_3__707_, data_stage_3__706_, data_stage_3__705_, data_stage_3__704_, data_stage_3__703_, data_stage_3__702_, data_stage_3__701_, data_stage_3__700_, data_stage_3__699_, data_stage_3__698_, data_stage_3__697_, data_stage_3__696_, data_stage_3__695_, data_stage_3__694_, data_stage_3__693_, data_stage_3__692_, data_stage_3__691_, data_stage_3__690_, data_stage_3__689_, data_stage_3__688_, data_stage_3__687_, data_stage_3__686_, data_stage_3__685_, data_stage_3__684_, data_stage_3__683_, data_stage_3__682_, data_stage_3__681_, data_stage_3__680_, data_stage_3__679_, data_stage_3__678_, data_stage_3__677_, data_stage_3__676_, data_stage_3__675_, data_stage_3__674_, data_stage_3__673_, data_stage_3__672_, data_stage_3__671_, data_stage_3__670_, data_stage_3__669_, data_stage_3__668_, data_stage_3__667_, data_stage_3__666_, data_stage_3__665_, data_stage_3__664_, data_stage_3__663_, data_stage_3__662_, data_stage_3__661_, data_stage_3__660_, data_stage_3__659_, data_stage_3__658_, data_stage_3__657_, data_stage_3__656_, data_stage_3__655_, data_stage_3__654_, data_stage_3__653_, data_stage_3__652_, data_stage_3__651_, data_stage_3__650_, data_stage_3__649_, data_stage_3__648_, data_stage_3__647_, data_stage_3__646_, data_stage_3__645_, data_stage_3__644_, data_stage_3__643_, data_stage_3__642_, data_stage_3__641_, data_stage_3__640_, data_stage_3__639_, data_stage_3__638_, data_stage_3__637_, data_stage_3__636_, data_stage_3__635_, data_stage_3__634_, data_stage_3__633_, data_stage_3__632_, data_stage_3__631_, data_stage_3__630_, data_stage_3__629_, data_stage_3__628_, data_stage_3__627_, data_stage_3__626_, data_stage_3__625_, data_stage_3__624_, data_stage_3__623_, data_stage_3__622_, data_stage_3__621_, data_stage_3__620_, data_stage_3__619_, data_stage_3__618_, data_stage_3__617_, data_stage_3__616_, data_stage_3__615_, data_stage_3__614_, data_stage_3__613_, data_stage_3__612_, data_stage_3__611_, data_stage_3__610_, data_stage_3__609_, data_stage_3__608_, data_stage_3__607_, data_stage_3__606_, data_stage_3__605_, data_stage_3__604_, data_stage_3__603_, data_stage_3__602_, data_stage_3__601_, data_stage_3__600_, data_stage_3__599_, data_stage_3__598_, data_stage_3__597_, data_stage_3__596_, data_stage_3__595_, data_stage_3__594_, data_stage_3__593_, data_stage_3__592_, data_stage_3__591_, data_stage_3__590_, data_stage_3__589_, data_stage_3__588_, data_stage_3__587_, data_stage_3__586_, data_stage_3__585_, data_stage_3__584_, data_stage_3__583_, data_stage_3__582_, data_stage_3__581_, data_stage_3__580_, data_stage_3__579_, data_stage_3__578_, data_stage_3__577_, data_stage_3__576_, data_stage_3__575_, data_stage_3__574_, data_stage_3__573_, data_stage_3__572_, data_stage_3__571_, data_stage_3__570_, data_stage_3__569_, data_stage_3__568_, data_stage_3__567_, data_stage_3__566_, data_stage_3__565_, data_stage_3__564_, data_stage_3__563_, data_stage_3__562_, data_stage_3__561_, data_stage_3__560_, data_stage_3__559_, data_stage_3__558_, data_stage_3__557_, data_stage_3__556_, data_stage_3__555_, data_stage_3__554_, data_stage_3__553_, data_stage_3__552_, data_stage_3__551_, data_stage_3__550_, data_stage_3__549_, data_stage_3__548_, data_stage_3__547_, data_stage_3__546_, data_stage_3__545_, data_stage_3__544_, data_stage_3__543_, data_stage_3__542_, data_stage_3__541_, data_stage_3__540_, data_stage_3__539_, data_stage_3__538_, data_stage_3__537_, data_stage_3__536_, data_stage_3__535_, data_stage_3__534_, data_stage_3__533_, data_stage_3__532_, data_stage_3__531_, data_stage_3__530_, data_stage_3__529_, data_stage_3__528_, data_stage_3__527_, data_stage_3__526_, data_stage_3__525_, data_stage_3__524_, data_stage_3__523_, data_stage_3__522_, data_stage_3__521_, data_stage_3__520_, data_stage_3__519_, data_stage_3__518_, data_stage_3__517_, data_stage_3__516_, data_stage_3__515_, data_stage_3__514_, data_stage_3__513_, data_stage_3__512_ })
  );


  bsg_swap_width_p128
  mux_stage_2__mux_swap_3__swap_inst
  (
    .data_i({ data_stage_2__1023_, data_stage_2__1022_, data_stage_2__1021_, data_stage_2__1020_, data_stage_2__1019_, data_stage_2__1018_, data_stage_2__1017_, data_stage_2__1016_, data_stage_2__1015_, data_stage_2__1014_, data_stage_2__1013_, data_stage_2__1012_, data_stage_2__1011_, data_stage_2__1010_, data_stage_2__1009_, data_stage_2__1008_, data_stage_2__1007_, data_stage_2__1006_, data_stage_2__1005_, data_stage_2__1004_, data_stage_2__1003_, data_stage_2__1002_, data_stage_2__1001_, data_stage_2__1000_, data_stage_2__999_, data_stage_2__998_, data_stage_2__997_, data_stage_2__996_, data_stage_2__995_, data_stage_2__994_, data_stage_2__993_, data_stage_2__992_, data_stage_2__991_, data_stage_2__990_, data_stage_2__989_, data_stage_2__988_, data_stage_2__987_, data_stage_2__986_, data_stage_2__985_, data_stage_2__984_, data_stage_2__983_, data_stage_2__982_, data_stage_2__981_, data_stage_2__980_, data_stage_2__979_, data_stage_2__978_, data_stage_2__977_, data_stage_2__976_, data_stage_2__975_, data_stage_2__974_, data_stage_2__973_, data_stage_2__972_, data_stage_2__971_, data_stage_2__970_, data_stage_2__969_, data_stage_2__968_, data_stage_2__967_, data_stage_2__966_, data_stage_2__965_, data_stage_2__964_, data_stage_2__963_, data_stage_2__962_, data_stage_2__961_, data_stage_2__960_, data_stage_2__959_, data_stage_2__958_, data_stage_2__957_, data_stage_2__956_, data_stage_2__955_, data_stage_2__954_, data_stage_2__953_, data_stage_2__952_, data_stage_2__951_, data_stage_2__950_, data_stage_2__949_, data_stage_2__948_, data_stage_2__947_, data_stage_2__946_, data_stage_2__945_, data_stage_2__944_, data_stage_2__943_, data_stage_2__942_, data_stage_2__941_, data_stage_2__940_, data_stage_2__939_, data_stage_2__938_, data_stage_2__937_, data_stage_2__936_, data_stage_2__935_, data_stage_2__934_, data_stage_2__933_, data_stage_2__932_, data_stage_2__931_, data_stage_2__930_, data_stage_2__929_, data_stage_2__928_, data_stage_2__927_, data_stage_2__926_, data_stage_2__925_, data_stage_2__924_, data_stage_2__923_, data_stage_2__922_, data_stage_2__921_, data_stage_2__920_, data_stage_2__919_, data_stage_2__918_, data_stage_2__917_, data_stage_2__916_, data_stage_2__915_, data_stage_2__914_, data_stage_2__913_, data_stage_2__912_, data_stage_2__911_, data_stage_2__910_, data_stage_2__909_, data_stage_2__908_, data_stage_2__907_, data_stage_2__906_, data_stage_2__905_, data_stage_2__904_, data_stage_2__903_, data_stage_2__902_, data_stage_2__901_, data_stage_2__900_, data_stage_2__899_, data_stage_2__898_, data_stage_2__897_, data_stage_2__896_, data_stage_2__895_, data_stage_2__894_, data_stage_2__893_, data_stage_2__892_, data_stage_2__891_, data_stage_2__890_, data_stage_2__889_, data_stage_2__888_, data_stage_2__887_, data_stage_2__886_, data_stage_2__885_, data_stage_2__884_, data_stage_2__883_, data_stage_2__882_, data_stage_2__881_, data_stage_2__880_, data_stage_2__879_, data_stage_2__878_, data_stage_2__877_, data_stage_2__876_, data_stage_2__875_, data_stage_2__874_, data_stage_2__873_, data_stage_2__872_, data_stage_2__871_, data_stage_2__870_, data_stage_2__869_, data_stage_2__868_, data_stage_2__867_, data_stage_2__866_, data_stage_2__865_, data_stage_2__864_, data_stage_2__863_, data_stage_2__862_, data_stage_2__861_, data_stage_2__860_, data_stage_2__859_, data_stage_2__858_, data_stage_2__857_, data_stage_2__856_, data_stage_2__855_, data_stage_2__854_, data_stage_2__853_, data_stage_2__852_, data_stage_2__851_, data_stage_2__850_, data_stage_2__849_, data_stage_2__848_, data_stage_2__847_, data_stage_2__846_, data_stage_2__845_, data_stage_2__844_, data_stage_2__843_, data_stage_2__842_, data_stage_2__841_, data_stage_2__840_, data_stage_2__839_, data_stage_2__838_, data_stage_2__837_, data_stage_2__836_, data_stage_2__835_, data_stage_2__834_, data_stage_2__833_, data_stage_2__832_, data_stage_2__831_, data_stage_2__830_, data_stage_2__829_, data_stage_2__828_, data_stage_2__827_, data_stage_2__826_, data_stage_2__825_, data_stage_2__824_, data_stage_2__823_, data_stage_2__822_, data_stage_2__821_, data_stage_2__820_, data_stage_2__819_, data_stage_2__818_, data_stage_2__817_, data_stage_2__816_, data_stage_2__815_, data_stage_2__814_, data_stage_2__813_, data_stage_2__812_, data_stage_2__811_, data_stage_2__810_, data_stage_2__809_, data_stage_2__808_, data_stage_2__807_, data_stage_2__806_, data_stage_2__805_, data_stage_2__804_, data_stage_2__803_, data_stage_2__802_, data_stage_2__801_, data_stage_2__800_, data_stage_2__799_, data_stage_2__798_, data_stage_2__797_, data_stage_2__796_, data_stage_2__795_, data_stage_2__794_, data_stage_2__793_, data_stage_2__792_, data_stage_2__791_, data_stage_2__790_, data_stage_2__789_, data_stage_2__788_, data_stage_2__787_, data_stage_2__786_, data_stage_2__785_, data_stage_2__784_, data_stage_2__783_, data_stage_2__782_, data_stage_2__781_, data_stage_2__780_, data_stage_2__779_, data_stage_2__778_, data_stage_2__777_, data_stage_2__776_, data_stage_2__775_, data_stage_2__774_, data_stage_2__773_, data_stage_2__772_, data_stage_2__771_, data_stage_2__770_, data_stage_2__769_, data_stage_2__768_ }),
    .swap_i(sel_i[2]),
    .data_o({ data_stage_3__1023_, data_stage_3__1022_, data_stage_3__1021_, data_stage_3__1020_, data_stage_3__1019_, data_stage_3__1018_, data_stage_3__1017_, data_stage_3__1016_, data_stage_3__1015_, data_stage_3__1014_, data_stage_3__1013_, data_stage_3__1012_, data_stage_3__1011_, data_stage_3__1010_, data_stage_3__1009_, data_stage_3__1008_, data_stage_3__1007_, data_stage_3__1006_, data_stage_3__1005_, data_stage_3__1004_, data_stage_3__1003_, data_stage_3__1002_, data_stage_3__1001_, data_stage_3__1000_, data_stage_3__999_, data_stage_3__998_, data_stage_3__997_, data_stage_3__996_, data_stage_3__995_, data_stage_3__994_, data_stage_3__993_, data_stage_3__992_, data_stage_3__991_, data_stage_3__990_, data_stage_3__989_, data_stage_3__988_, data_stage_3__987_, data_stage_3__986_, data_stage_3__985_, data_stage_3__984_, data_stage_3__983_, data_stage_3__982_, data_stage_3__981_, data_stage_3__980_, data_stage_3__979_, data_stage_3__978_, data_stage_3__977_, data_stage_3__976_, data_stage_3__975_, data_stage_3__974_, data_stage_3__973_, data_stage_3__972_, data_stage_3__971_, data_stage_3__970_, data_stage_3__969_, data_stage_3__968_, data_stage_3__967_, data_stage_3__966_, data_stage_3__965_, data_stage_3__964_, data_stage_3__963_, data_stage_3__962_, data_stage_3__961_, data_stage_3__960_, data_stage_3__959_, data_stage_3__958_, data_stage_3__957_, data_stage_3__956_, data_stage_3__955_, data_stage_3__954_, data_stage_3__953_, data_stage_3__952_, data_stage_3__951_, data_stage_3__950_, data_stage_3__949_, data_stage_3__948_, data_stage_3__947_, data_stage_3__946_, data_stage_3__945_, data_stage_3__944_, data_stage_3__943_, data_stage_3__942_, data_stage_3__941_, data_stage_3__940_, data_stage_3__939_, data_stage_3__938_, data_stage_3__937_, data_stage_3__936_, data_stage_3__935_, data_stage_3__934_, data_stage_3__933_, data_stage_3__932_, data_stage_3__931_, data_stage_3__930_, data_stage_3__929_, data_stage_3__928_, data_stage_3__927_, data_stage_3__926_, data_stage_3__925_, data_stage_3__924_, data_stage_3__923_, data_stage_3__922_, data_stage_3__921_, data_stage_3__920_, data_stage_3__919_, data_stage_3__918_, data_stage_3__917_, data_stage_3__916_, data_stage_3__915_, data_stage_3__914_, data_stage_3__913_, data_stage_3__912_, data_stage_3__911_, data_stage_3__910_, data_stage_3__909_, data_stage_3__908_, data_stage_3__907_, data_stage_3__906_, data_stage_3__905_, data_stage_3__904_, data_stage_3__903_, data_stage_3__902_, data_stage_3__901_, data_stage_3__900_, data_stage_3__899_, data_stage_3__898_, data_stage_3__897_, data_stage_3__896_, data_stage_3__895_, data_stage_3__894_, data_stage_3__893_, data_stage_3__892_, data_stage_3__891_, data_stage_3__890_, data_stage_3__889_, data_stage_3__888_, data_stage_3__887_, data_stage_3__886_, data_stage_3__885_, data_stage_3__884_, data_stage_3__883_, data_stage_3__882_, data_stage_3__881_, data_stage_3__880_, data_stage_3__879_, data_stage_3__878_, data_stage_3__877_, data_stage_3__876_, data_stage_3__875_, data_stage_3__874_, data_stage_3__873_, data_stage_3__872_, data_stage_3__871_, data_stage_3__870_, data_stage_3__869_, data_stage_3__868_, data_stage_3__867_, data_stage_3__866_, data_stage_3__865_, data_stage_3__864_, data_stage_3__863_, data_stage_3__862_, data_stage_3__861_, data_stage_3__860_, data_stage_3__859_, data_stage_3__858_, data_stage_3__857_, data_stage_3__856_, data_stage_3__855_, data_stage_3__854_, data_stage_3__853_, data_stage_3__852_, data_stage_3__851_, data_stage_3__850_, data_stage_3__849_, data_stage_3__848_, data_stage_3__847_, data_stage_3__846_, data_stage_3__845_, data_stage_3__844_, data_stage_3__843_, data_stage_3__842_, data_stage_3__841_, data_stage_3__840_, data_stage_3__839_, data_stage_3__838_, data_stage_3__837_, data_stage_3__836_, data_stage_3__835_, data_stage_3__834_, data_stage_3__833_, data_stage_3__832_, data_stage_3__831_, data_stage_3__830_, data_stage_3__829_, data_stage_3__828_, data_stage_3__827_, data_stage_3__826_, data_stage_3__825_, data_stage_3__824_, data_stage_3__823_, data_stage_3__822_, data_stage_3__821_, data_stage_3__820_, data_stage_3__819_, data_stage_3__818_, data_stage_3__817_, data_stage_3__816_, data_stage_3__815_, data_stage_3__814_, data_stage_3__813_, data_stage_3__812_, data_stage_3__811_, data_stage_3__810_, data_stage_3__809_, data_stage_3__808_, data_stage_3__807_, data_stage_3__806_, data_stage_3__805_, data_stage_3__804_, data_stage_3__803_, data_stage_3__802_, data_stage_3__801_, data_stage_3__800_, data_stage_3__799_, data_stage_3__798_, data_stage_3__797_, data_stage_3__796_, data_stage_3__795_, data_stage_3__794_, data_stage_3__793_, data_stage_3__792_, data_stage_3__791_, data_stage_3__790_, data_stage_3__789_, data_stage_3__788_, data_stage_3__787_, data_stage_3__786_, data_stage_3__785_, data_stage_3__784_, data_stage_3__783_, data_stage_3__782_, data_stage_3__781_, data_stage_3__780_, data_stage_3__779_, data_stage_3__778_, data_stage_3__777_, data_stage_3__776_, data_stage_3__775_, data_stage_3__774_, data_stage_3__773_, data_stage_3__772_, data_stage_3__771_, data_stage_3__770_, data_stage_3__769_, data_stage_3__768_ })
  );


  bsg_swap_width_p256
  mux_stage_3__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_3__511_, data_stage_3__510_, data_stage_3__509_, data_stage_3__508_, data_stage_3__507_, data_stage_3__506_, data_stage_3__505_, data_stage_3__504_, data_stage_3__503_, data_stage_3__502_, data_stage_3__501_, data_stage_3__500_, data_stage_3__499_, data_stage_3__498_, data_stage_3__497_, data_stage_3__496_, data_stage_3__495_, data_stage_3__494_, data_stage_3__493_, data_stage_3__492_, data_stage_3__491_, data_stage_3__490_, data_stage_3__489_, data_stage_3__488_, data_stage_3__487_, data_stage_3__486_, data_stage_3__485_, data_stage_3__484_, data_stage_3__483_, data_stage_3__482_, data_stage_3__481_, data_stage_3__480_, data_stage_3__479_, data_stage_3__478_, data_stage_3__477_, data_stage_3__476_, data_stage_3__475_, data_stage_3__474_, data_stage_3__473_, data_stage_3__472_, data_stage_3__471_, data_stage_3__470_, data_stage_3__469_, data_stage_3__468_, data_stage_3__467_, data_stage_3__466_, data_stage_3__465_, data_stage_3__464_, data_stage_3__463_, data_stage_3__462_, data_stage_3__461_, data_stage_3__460_, data_stage_3__459_, data_stage_3__458_, data_stage_3__457_, data_stage_3__456_, data_stage_3__455_, data_stage_3__454_, data_stage_3__453_, data_stage_3__452_, data_stage_3__451_, data_stage_3__450_, data_stage_3__449_, data_stage_3__448_, data_stage_3__447_, data_stage_3__446_, data_stage_3__445_, data_stage_3__444_, data_stage_3__443_, data_stage_3__442_, data_stage_3__441_, data_stage_3__440_, data_stage_3__439_, data_stage_3__438_, data_stage_3__437_, data_stage_3__436_, data_stage_3__435_, data_stage_3__434_, data_stage_3__433_, data_stage_3__432_, data_stage_3__431_, data_stage_3__430_, data_stage_3__429_, data_stage_3__428_, data_stage_3__427_, data_stage_3__426_, data_stage_3__425_, data_stage_3__424_, data_stage_3__423_, data_stage_3__422_, data_stage_3__421_, data_stage_3__420_, data_stage_3__419_, data_stage_3__418_, data_stage_3__417_, data_stage_3__416_, data_stage_3__415_, data_stage_3__414_, data_stage_3__413_, data_stage_3__412_, data_stage_3__411_, data_stage_3__410_, data_stage_3__409_, data_stage_3__408_, data_stage_3__407_, data_stage_3__406_, data_stage_3__405_, data_stage_3__404_, data_stage_3__403_, data_stage_3__402_, data_stage_3__401_, data_stage_3__400_, data_stage_3__399_, data_stage_3__398_, data_stage_3__397_, data_stage_3__396_, data_stage_3__395_, data_stage_3__394_, data_stage_3__393_, data_stage_3__392_, data_stage_3__391_, data_stage_3__390_, data_stage_3__389_, data_stage_3__388_, data_stage_3__387_, data_stage_3__386_, data_stage_3__385_, data_stage_3__384_, data_stage_3__383_, data_stage_3__382_, data_stage_3__381_, data_stage_3__380_, data_stage_3__379_, data_stage_3__378_, data_stage_3__377_, data_stage_3__376_, data_stage_3__375_, data_stage_3__374_, data_stage_3__373_, data_stage_3__372_, data_stage_3__371_, data_stage_3__370_, data_stage_3__369_, data_stage_3__368_, data_stage_3__367_, data_stage_3__366_, data_stage_3__365_, data_stage_3__364_, data_stage_3__363_, data_stage_3__362_, data_stage_3__361_, data_stage_3__360_, data_stage_3__359_, data_stage_3__358_, data_stage_3__357_, data_stage_3__356_, data_stage_3__355_, data_stage_3__354_, data_stage_3__353_, data_stage_3__352_, data_stage_3__351_, data_stage_3__350_, data_stage_3__349_, data_stage_3__348_, data_stage_3__347_, data_stage_3__346_, data_stage_3__345_, data_stage_3__344_, data_stage_3__343_, data_stage_3__342_, data_stage_3__341_, data_stage_3__340_, data_stage_3__339_, data_stage_3__338_, data_stage_3__337_, data_stage_3__336_, data_stage_3__335_, data_stage_3__334_, data_stage_3__333_, data_stage_3__332_, data_stage_3__331_, data_stage_3__330_, data_stage_3__329_, data_stage_3__328_, data_stage_3__327_, data_stage_3__326_, data_stage_3__325_, data_stage_3__324_, data_stage_3__323_, data_stage_3__322_, data_stage_3__321_, data_stage_3__320_, data_stage_3__319_, data_stage_3__318_, data_stage_3__317_, data_stage_3__316_, data_stage_3__315_, data_stage_3__314_, data_stage_3__313_, data_stage_3__312_, data_stage_3__311_, data_stage_3__310_, data_stage_3__309_, data_stage_3__308_, data_stage_3__307_, data_stage_3__306_, data_stage_3__305_, data_stage_3__304_, data_stage_3__303_, data_stage_3__302_, data_stage_3__301_, data_stage_3__300_, data_stage_3__299_, data_stage_3__298_, data_stage_3__297_, data_stage_3__296_, data_stage_3__295_, data_stage_3__294_, data_stage_3__293_, data_stage_3__292_, data_stage_3__291_, data_stage_3__290_, data_stage_3__289_, data_stage_3__288_, data_stage_3__287_, data_stage_3__286_, data_stage_3__285_, data_stage_3__284_, data_stage_3__283_, data_stage_3__282_, data_stage_3__281_, data_stage_3__280_, data_stage_3__279_, data_stage_3__278_, data_stage_3__277_, data_stage_3__276_, data_stage_3__275_, data_stage_3__274_, data_stage_3__273_, data_stage_3__272_, data_stage_3__271_, data_stage_3__270_, data_stage_3__269_, data_stage_3__268_, data_stage_3__267_, data_stage_3__266_, data_stage_3__265_, data_stage_3__264_, data_stage_3__263_, data_stage_3__262_, data_stage_3__261_, data_stage_3__260_, data_stage_3__259_, data_stage_3__258_, data_stage_3__257_, data_stage_3__256_, data_stage_3__255_, data_stage_3__254_, data_stage_3__253_, data_stage_3__252_, data_stage_3__251_, data_stage_3__250_, data_stage_3__249_, data_stage_3__248_, data_stage_3__247_, data_stage_3__246_, data_stage_3__245_, data_stage_3__244_, data_stage_3__243_, data_stage_3__242_, data_stage_3__241_, data_stage_3__240_, data_stage_3__239_, data_stage_3__238_, data_stage_3__237_, data_stage_3__236_, data_stage_3__235_, data_stage_3__234_, data_stage_3__233_, data_stage_3__232_, data_stage_3__231_, data_stage_3__230_, data_stage_3__229_, data_stage_3__228_, data_stage_3__227_, data_stage_3__226_, data_stage_3__225_, data_stage_3__224_, data_stage_3__223_, data_stage_3__222_, data_stage_3__221_, data_stage_3__220_, data_stage_3__219_, data_stage_3__218_, data_stage_3__217_, data_stage_3__216_, data_stage_3__215_, data_stage_3__214_, data_stage_3__213_, data_stage_3__212_, data_stage_3__211_, data_stage_3__210_, data_stage_3__209_, data_stage_3__208_, data_stage_3__207_, data_stage_3__206_, data_stage_3__205_, data_stage_3__204_, data_stage_3__203_, data_stage_3__202_, data_stage_3__201_, data_stage_3__200_, data_stage_3__199_, data_stage_3__198_, data_stage_3__197_, data_stage_3__196_, data_stage_3__195_, data_stage_3__194_, data_stage_3__193_, data_stage_3__192_, data_stage_3__191_, data_stage_3__190_, data_stage_3__189_, data_stage_3__188_, data_stage_3__187_, data_stage_3__186_, data_stage_3__185_, data_stage_3__184_, data_stage_3__183_, data_stage_3__182_, data_stage_3__181_, data_stage_3__180_, data_stage_3__179_, data_stage_3__178_, data_stage_3__177_, data_stage_3__176_, data_stage_3__175_, data_stage_3__174_, data_stage_3__173_, data_stage_3__172_, data_stage_3__171_, data_stage_3__170_, data_stage_3__169_, data_stage_3__168_, data_stage_3__167_, data_stage_3__166_, data_stage_3__165_, data_stage_3__164_, data_stage_3__163_, data_stage_3__162_, data_stage_3__161_, data_stage_3__160_, data_stage_3__159_, data_stage_3__158_, data_stage_3__157_, data_stage_3__156_, data_stage_3__155_, data_stage_3__154_, data_stage_3__153_, data_stage_3__152_, data_stage_3__151_, data_stage_3__150_, data_stage_3__149_, data_stage_3__148_, data_stage_3__147_, data_stage_3__146_, data_stage_3__145_, data_stage_3__144_, data_stage_3__143_, data_stage_3__142_, data_stage_3__141_, data_stage_3__140_, data_stage_3__139_, data_stage_3__138_, data_stage_3__137_, data_stage_3__136_, data_stage_3__135_, data_stage_3__134_, data_stage_3__133_, data_stage_3__132_, data_stage_3__131_, data_stage_3__130_, data_stage_3__129_, data_stage_3__128_, data_stage_3__127_, data_stage_3__126_, data_stage_3__125_, data_stage_3__124_, data_stage_3__123_, data_stage_3__122_, data_stage_3__121_, data_stage_3__120_, data_stage_3__119_, data_stage_3__118_, data_stage_3__117_, data_stage_3__116_, data_stage_3__115_, data_stage_3__114_, data_stage_3__113_, data_stage_3__112_, data_stage_3__111_, data_stage_3__110_, data_stage_3__109_, data_stage_3__108_, data_stage_3__107_, data_stage_3__106_, data_stage_3__105_, data_stage_3__104_, data_stage_3__103_, data_stage_3__102_, data_stage_3__101_, data_stage_3__100_, data_stage_3__99_, data_stage_3__98_, data_stage_3__97_, data_stage_3__96_, data_stage_3__95_, data_stage_3__94_, data_stage_3__93_, data_stage_3__92_, data_stage_3__91_, data_stage_3__90_, data_stage_3__89_, data_stage_3__88_, data_stage_3__87_, data_stage_3__86_, data_stage_3__85_, data_stage_3__84_, data_stage_3__83_, data_stage_3__82_, data_stage_3__81_, data_stage_3__80_, data_stage_3__79_, data_stage_3__78_, data_stage_3__77_, data_stage_3__76_, data_stage_3__75_, data_stage_3__74_, data_stage_3__73_, data_stage_3__72_, data_stage_3__71_, data_stage_3__70_, data_stage_3__69_, data_stage_3__68_, data_stage_3__67_, data_stage_3__66_, data_stage_3__65_, data_stage_3__64_, data_stage_3__63_, data_stage_3__62_, data_stage_3__61_, data_stage_3__60_, data_stage_3__59_, data_stage_3__58_, data_stage_3__57_, data_stage_3__56_, data_stage_3__55_, data_stage_3__54_, data_stage_3__53_, data_stage_3__52_, data_stage_3__51_, data_stage_3__50_, data_stage_3__49_, data_stage_3__48_, data_stage_3__47_, data_stage_3__46_, data_stage_3__45_, data_stage_3__44_, data_stage_3__43_, data_stage_3__42_, data_stage_3__41_, data_stage_3__40_, data_stage_3__39_, data_stage_3__38_, data_stage_3__37_, data_stage_3__36_, data_stage_3__35_, data_stage_3__34_, data_stage_3__33_, data_stage_3__32_, data_stage_3__31_, data_stage_3__30_, data_stage_3__29_, data_stage_3__28_, data_stage_3__27_, data_stage_3__26_, data_stage_3__25_, data_stage_3__24_, data_stage_3__23_, data_stage_3__22_, data_stage_3__21_, data_stage_3__20_, data_stage_3__19_, data_stage_3__18_, data_stage_3__17_, data_stage_3__16_, data_stage_3__15_, data_stage_3__14_, data_stage_3__13_, data_stage_3__12_, data_stage_3__11_, data_stage_3__10_, data_stage_3__9_, data_stage_3__8_, data_stage_3__7_, data_stage_3__6_, data_stage_3__5_, data_stage_3__4_, data_stage_3__3_, data_stage_3__2_, data_stage_3__1_, data_stage_3__0_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__511_, data_stage_4__510_, data_stage_4__509_, data_stage_4__508_, data_stage_4__507_, data_stage_4__506_, data_stage_4__505_, data_stage_4__504_, data_stage_4__503_, data_stage_4__502_, data_stage_4__501_, data_stage_4__500_, data_stage_4__499_, data_stage_4__498_, data_stage_4__497_, data_stage_4__496_, data_stage_4__495_, data_stage_4__494_, data_stage_4__493_, data_stage_4__492_, data_stage_4__491_, data_stage_4__490_, data_stage_4__489_, data_stage_4__488_, data_stage_4__487_, data_stage_4__486_, data_stage_4__485_, data_stage_4__484_, data_stage_4__483_, data_stage_4__482_, data_stage_4__481_, data_stage_4__480_, data_stage_4__479_, data_stage_4__478_, data_stage_4__477_, data_stage_4__476_, data_stage_4__475_, data_stage_4__474_, data_stage_4__473_, data_stage_4__472_, data_stage_4__471_, data_stage_4__470_, data_stage_4__469_, data_stage_4__468_, data_stage_4__467_, data_stage_4__466_, data_stage_4__465_, data_stage_4__464_, data_stage_4__463_, data_stage_4__462_, data_stage_4__461_, data_stage_4__460_, data_stage_4__459_, data_stage_4__458_, data_stage_4__457_, data_stage_4__456_, data_stage_4__455_, data_stage_4__454_, data_stage_4__453_, data_stage_4__452_, data_stage_4__451_, data_stage_4__450_, data_stage_4__449_, data_stage_4__448_, data_stage_4__447_, data_stage_4__446_, data_stage_4__445_, data_stage_4__444_, data_stage_4__443_, data_stage_4__442_, data_stage_4__441_, data_stage_4__440_, data_stage_4__439_, data_stage_4__438_, data_stage_4__437_, data_stage_4__436_, data_stage_4__435_, data_stage_4__434_, data_stage_4__433_, data_stage_4__432_, data_stage_4__431_, data_stage_4__430_, data_stage_4__429_, data_stage_4__428_, data_stage_4__427_, data_stage_4__426_, data_stage_4__425_, data_stage_4__424_, data_stage_4__423_, data_stage_4__422_, data_stage_4__421_, data_stage_4__420_, data_stage_4__419_, data_stage_4__418_, data_stage_4__417_, data_stage_4__416_, data_stage_4__415_, data_stage_4__414_, data_stage_4__413_, data_stage_4__412_, data_stage_4__411_, data_stage_4__410_, data_stage_4__409_, data_stage_4__408_, data_stage_4__407_, data_stage_4__406_, data_stage_4__405_, data_stage_4__404_, data_stage_4__403_, data_stage_4__402_, data_stage_4__401_, data_stage_4__400_, data_stage_4__399_, data_stage_4__398_, data_stage_4__397_, data_stage_4__396_, data_stage_4__395_, data_stage_4__394_, data_stage_4__393_, data_stage_4__392_, data_stage_4__391_, data_stage_4__390_, data_stage_4__389_, data_stage_4__388_, data_stage_4__387_, data_stage_4__386_, data_stage_4__385_, data_stage_4__384_, data_stage_4__383_, data_stage_4__382_, data_stage_4__381_, data_stage_4__380_, data_stage_4__379_, data_stage_4__378_, data_stage_4__377_, data_stage_4__376_, data_stage_4__375_, data_stage_4__374_, data_stage_4__373_, data_stage_4__372_, data_stage_4__371_, data_stage_4__370_, data_stage_4__369_, data_stage_4__368_, data_stage_4__367_, data_stage_4__366_, data_stage_4__365_, data_stage_4__364_, data_stage_4__363_, data_stage_4__362_, data_stage_4__361_, data_stage_4__360_, data_stage_4__359_, data_stage_4__358_, data_stage_4__357_, data_stage_4__356_, data_stage_4__355_, data_stage_4__354_, data_stage_4__353_, data_stage_4__352_, data_stage_4__351_, data_stage_4__350_, data_stage_4__349_, data_stage_4__348_, data_stage_4__347_, data_stage_4__346_, data_stage_4__345_, data_stage_4__344_, data_stage_4__343_, data_stage_4__342_, data_stage_4__341_, data_stage_4__340_, data_stage_4__339_, data_stage_4__338_, data_stage_4__337_, data_stage_4__336_, data_stage_4__335_, data_stage_4__334_, data_stage_4__333_, data_stage_4__332_, data_stage_4__331_, data_stage_4__330_, data_stage_4__329_, data_stage_4__328_, data_stage_4__327_, data_stage_4__326_, data_stage_4__325_, data_stage_4__324_, data_stage_4__323_, data_stage_4__322_, data_stage_4__321_, data_stage_4__320_, data_stage_4__319_, data_stage_4__318_, data_stage_4__317_, data_stage_4__316_, data_stage_4__315_, data_stage_4__314_, data_stage_4__313_, data_stage_4__312_, data_stage_4__311_, data_stage_4__310_, data_stage_4__309_, data_stage_4__308_, data_stage_4__307_, data_stage_4__306_, data_stage_4__305_, data_stage_4__304_, data_stage_4__303_, data_stage_4__302_, data_stage_4__301_, data_stage_4__300_, data_stage_4__299_, data_stage_4__298_, data_stage_4__297_, data_stage_4__296_, data_stage_4__295_, data_stage_4__294_, data_stage_4__293_, data_stage_4__292_, data_stage_4__291_, data_stage_4__290_, data_stage_4__289_, data_stage_4__288_, data_stage_4__287_, data_stage_4__286_, data_stage_4__285_, data_stage_4__284_, data_stage_4__283_, data_stage_4__282_, data_stage_4__281_, data_stage_4__280_, data_stage_4__279_, data_stage_4__278_, data_stage_4__277_, data_stage_4__276_, data_stage_4__275_, data_stage_4__274_, data_stage_4__273_, data_stage_4__272_, data_stage_4__271_, data_stage_4__270_, data_stage_4__269_, data_stage_4__268_, data_stage_4__267_, data_stage_4__266_, data_stage_4__265_, data_stage_4__264_, data_stage_4__263_, data_stage_4__262_, data_stage_4__261_, data_stage_4__260_, data_stage_4__259_, data_stage_4__258_, data_stage_4__257_, data_stage_4__256_, data_stage_4__255_, data_stage_4__254_, data_stage_4__253_, data_stage_4__252_, data_stage_4__251_, data_stage_4__250_, data_stage_4__249_, data_stage_4__248_, data_stage_4__247_, data_stage_4__246_, data_stage_4__245_, data_stage_4__244_, data_stage_4__243_, data_stage_4__242_, data_stage_4__241_, data_stage_4__240_, data_stage_4__239_, data_stage_4__238_, data_stage_4__237_, data_stage_4__236_, data_stage_4__235_, data_stage_4__234_, data_stage_4__233_, data_stage_4__232_, data_stage_4__231_, data_stage_4__230_, data_stage_4__229_, data_stage_4__228_, data_stage_4__227_, data_stage_4__226_, data_stage_4__225_, data_stage_4__224_, data_stage_4__223_, data_stage_4__222_, data_stage_4__221_, data_stage_4__220_, data_stage_4__219_, data_stage_4__218_, data_stage_4__217_, data_stage_4__216_, data_stage_4__215_, data_stage_4__214_, data_stage_4__213_, data_stage_4__212_, data_stage_4__211_, data_stage_4__210_, data_stage_4__209_, data_stage_4__208_, data_stage_4__207_, data_stage_4__206_, data_stage_4__205_, data_stage_4__204_, data_stage_4__203_, data_stage_4__202_, data_stage_4__201_, data_stage_4__200_, data_stage_4__199_, data_stage_4__198_, data_stage_4__197_, data_stage_4__196_, data_stage_4__195_, data_stage_4__194_, data_stage_4__193_, data_stage_4__192_, data_stage_4__191_, data_stage_4__190_, data_stage_4__189_, data_stage_4__188_, data_stage_4__187_, data_stage_4__186_, data_stage_4__185_, data_stage_4__184_, data_stage_4__183_, data_stage_4__182_, data_stage_4__181_, data_stage_4__180_, data_stage_4__179_, data_stage_4__178_, data_stage_4__177_, data_stage_4__176_, data_stage_4__175_, data_stage_4__174_, data_stage_4__173_, data_stage_4__172_, data_stage_4__171_, data_stage_4__170_, data_stage_4__169_, data_stage_4__168_, data_stage_4__167_, data_stage_4__166_, data_stage_4__165_, data_stage_4__164_, data_stage_4__163_, data_stage_4__162_, data_stage_4__161_, data_stage_4__160_, data_stage_4__159_, data_stage_4__158_, data_stage_4__157_, data_stage_4__156_, data_stage_4__155_, data_stage_4__154_, data_stage_4__153_, data_stage_4__152_, data_stage_4__151_, data_stage_4__150_, data_stage_4__149_, data_stage_4__148_, data_stage_4__147_, data_stage_4__146_, data_stage_4__145_, data_stage_4__144_, data_stage_4__143_, data_stage_4__142_, data_stage_4__141_, data_stage_4__140_, data_stage_4__139_, data_stage_4__138_, data_stage_4__137_, data_stage_4__136_, data_stage_4__135_, data_stage_4__134_, data_stage_4__133_, data_stage_4__132_, data_stage_4__131_, data_stage_4__130_, data_stage_4__129_, data_stage_4__128_, data_stage_4__127_, data_stage_4__126_, data_stage_4__125_, data_stage_4__124_, data_stage_4__123_, data_stage_4__122_, data_stage_4__121_, data_stage_4__120_, data_stage_4__119_, data_stage_4__118_, data_stage_4__117_, data_stage_4__116_, data_stage_4__115_, data_stage_4__114_, data_stage_4__113_, data_stage_4__112_, data_stage_4__111_, data_stage_4__110_, data_stage_4__109_, data_stage_4__108_, data_stage_4__107_, data_stage_4__106_, data_stage_4__105_, data_stage_4__104_, data_stage_4__103_, data_stage_4__102_, data_stage_4__101_, data_stage_4__100_, data_stage_4__99_, data_stage_4__98_, data_stage_4__97_, data_stage_4__96_, data_stage_4__95_, data_stage_4__94_, data_stage_4__93_, data_stage_4__92_, data_stage_4__91_, data_stage_4__90_, data_stage_4__89_, data_stage_4__88_, data_stage_4__87_, data_stage_4__86_, data_stage_4__85_, data_stage_4__84_, data_stage_4__83_, data_stage_4__82_, data_stage_4__81_, data_stage_4__80_, data_stage_4__79_, data_stage_4__78_, data_stage_4__77_, data_stage_4__76_, data_stage_4__75_, data_stage_4__74_, data_stage_4__73_, data_stage_4__72_, data_stage_4__71_, data_stage_4__70_, data_stage_4__69_, data_stage_4__68_, data_stage_4__67_, data_stage_4__66_, data_stage_4__65_, data_stage_4__64_, data_stage_4__63_, data_stage_4__62_, data_stage_4__61_, data_stage_4__60_, data_stage_4__59_, data_stage_4__58_, data_stage_4__57_, data_stage_4__56_, data_stage_4__55_, data_stage_4__54_, data_stage_4__53_, data_stage_4__52_, data_stage_4__51_, data_stage_4__50_, data_stage_4__49_, data_stage_4__48_, data_stage_4__47_, data_stage_4__46_, data_stage_4__45_, data_stage_4__44_, data_stage_4__43_, data_stage_4__42_, data_stage_4__41_, data_stage_4__40_, data_stage_4__39_, data_stage_4__38_, data_stage_4__37_, data_stage_4__36_, data_stage_4__35_, data_stage_4__34_, data_stage_4__33_, data_stage_4__32_, data_stage_4__31_, data_stage_4__30_, data_stage_4__29_, data_stage_4__28_, data_stage_4__27_, data_stage_4__26_, data_stage_4__25_, data_stage_4__24_, data_stage_4__23_, data_stage_4__22_, data_stage_4__21_, data_stage_4__20_, data_stage_4__19_, data_stage_4__18_, data_stage_4__17_, data_stage_4__16_, data_stage_4__15_, data_stage_4__14_, data_stage_4__13_, data_stage_4__12_, data_stage_4__11_, data_stage_4__10_, data_stage_4__9_, data_stage_4__8_, data_stage_4__7_, data_stage_4__6_, data_stage_4__5_, data_stage_4__4_, data_stage_4__3_, data_stage_4__2_, data_stage_4__1_, data_stage_4__0_ })
  );


  bsg_swap_width_p256
  mux_stage_3__mux_swap_1__swap_inst
  (
    .data_i({ data_stage_3__1023_, data_stage_3__1022_, data_stage_3__1021_, data_stage_3__1020_, data_stage_3__1019_, data_stage_3__1018_, data_stage_3__1017_, data_stage_3__1016_, data_stage_3__1015_, data_stage_3__1014_, data_stage_3__1013_, data_stage_3__1012_, data_stage_3__1011_, data_stage_3__1010_, data_stage_3__1009_, data_stage_3__1008_, data_stage_3__1007_, data_stage_3__1006_, data_stage_3__1005_, data_stage_3__1004_, data_stage_3__1003_, data_stage_3__1002_, data_stage_3__1001_, data_stage_3__1000_, data_stage_3__999_, data_stage_3__998_, data_stage_3__997_, data_stage_3__996_, data_stage_3__995_, data_stage_3__994_, data_stage_3__993_, data_stage_3__992_, data_stage_3__991_, data_stage_3__990_, data_stage_3__989_, data_stage_3__988_, data_stage_3__987_, data_stage_3__986_, data_stage_3__985_, data_stage_3__984_, data_stage_3__983_, data_stage_3__982_, data_stage_3__981_, data_stage_3__980_, data_stage_3__979_, data_stage_3__978_, data_stage_3__977_, data_stage_3__976_, data_stage_3__975_, data_stage_3__974_, data_stage_3__973_, data_stage_3__972_, data_stage_3__971_, data_stage_3__970_, data_stage_3__969_, data_stage_3__968_, data_stage_3__967_, data_stage_3__966_, data_stage_3__965_, data_stage_3__964_, data_stage_3__963_, data_stage_3__962_, data_stage_3__961_, data_stage_3__960_, data_stage_3__959_, data_stage_3__958_, data_stage_3__957_, data_stage_3__956_, data_stage_3__955_, data_stage_3__954_, data_stage_3__953_, data_stage_3__952_, data_stage_3__951_, data_stage_3__950_, data_stage_3__949_, data_stage_3__948_, data_stage_3__947_, data_stage_3__946_, data_stage_3__945_, data_stage_3__944_, data_stage_3__943_, data_stage_3__942_, data_stage_3__941_, data_stage_3__940_, data_stage_3__939_, data_stage_3__938_, data_stage_3__937_, data_stage_3__936_, data_stage_3__935_, data_stage_3__934_, data_stage_3__933_, data_stage_3__932_, data_stage_3__931_, data_stage_3__930_, data_stage_3__929_, data_stage_3__928_, data_stage_3__927_, data_stage_3__926_, data_stage_3__925_, data_stage_3__924_, data_stage_3__923_, data_stage_3__922_, data_stage_3__921_, data_stage_3__920_, data_stage_3__919_, data_stage_3__918_, data_stage_3__917_, data_stage_3__916_, data_stage_3__915_, data_stage_3__914_, data_stage_3__913_, data_stage_3__912_, data_stage_3__911_, data_stage_3__910_, data_stage_3__909_, data_stage_3__908_, data_stage_3__907_, data_stage_3__906_, data_stage_3__905_, data_stage_3__904_, data_stage_3__903_, data_stage_3__902_, data_stage_3__901_, data_stage_3__900_, data_stage_3__899_, data_stage_3__898_, data_stage_3__897_, data_stage_3__896_, data_stage_3__895_, data_stage_3__894_, data_stage_3__893_, data_stage_3__892_, data_stage_3__891_, data_stage_3__890_, data_stage_3__889_, data_stage_3__888_, data_stage_3__887_, data_stage_3__886_, data_stage_3__885_, data_stage_3__884_, data_stage_3__883_, data_stage_3__882_, data_stage_3__881_, data_stage_3__880_, data_stage_3__879_, data_stage_3__878_, data_stage_3__877_, data_stage_3__876_, data_stage_3__875_, data_stage_3__874_, data_stage_3__873_, data_stage_3__872_, data_stage_3__871_, data_stage_3__870_, data_stage_3__869_, data_stage_3__868_, data_stage_3__867_, data_stage_3__866_, data_stage_3__865_, data_stage_3__864_, data_stage_3__863_, data_stage_3__862_, data_stage_3__861_, data_stage_3__860_, data_stage_3__859_, data_stage_3__858_, data_stage_3__857_, data_stage_3__856_, data_stage_3__855_, data_stage_3__854_, data_stage_3__853_, data_stage_3__852_, data_stage_3__851_, data_stage_3__850_, data_stage_3__849_, data_stage_3__848_, data_stage_3__847_, data_stage_3__846_, data_stage_3__845_, data_stage_3__844_, data_stage_3__843_, data_stage_3__842_, data_stage_3__841_, data_stage_3__840_, data_stage_3__839_, data_stage_3__838_, data_stage_3__837_, data_stage_3__836_, data_stage_3__835_, data_stage_3__834_, data_stage_3__833_, data_stage_3__832_, data_stage_3__831_, data_stage_3__830_, data_stage_3__829_, data_stage_3__828_, data_stage_3__827_, data_stage_3__826_, data_stage_3__825_, data_stage_3__824_, data_stage_3__823_, data_stage_3__822_, data_stage_3__821_, data_stage_3__820_, data_stage_3__819_, data_stage_3__818_, data_stage_3__817_, data_stage_3__816_, data_stage_3__815_, data_stage_3__814_, data_stage_3__813_, data_stage_3__812_, data_stage_3__811_, data_stage_3__810_, data_stage_3__809_, data_stage_3__808_, data_stage_3__807_, data_stage_3__806_, data_stage_3__805_, data_stage_3__804_, data_stage_3__803_, data_stage_3__802_, data_stage_3__801_, data_stage_3__800_, data_stage_3__799_, data_stage_3__798_, data_stage_3__797_, data_stage_3__796_, data_stage_3__795_, data_stage_3__794_, data_stage_3__793_, data_stage_3__792_, data_stage_3__791_, data_stage_3__790_, data_stage_3__789_, data_stage_3__788_, data_stage_3__787_, data_stage_3__786_, data_stage_3__785_, data_stage_3__784_, data_stage_3__783_, data_stage_3__782_, data_stage_3__781_, data_stage_3__780_, data_stage_3__779_, data_stage_3__778_, data_stage_3__777_, data_stage_3__776_, data_stage_3__775_, data_stage_3__774_, data_stage_3__773_, data_stage_3__772_, data_stage_3__771_, data_stage_3__770_, data_stage_3__769_, data_stage_3__768_, data_stage_3__767_, data_stage_3__766_, data_stage_3__765_, data_stage_3__764_, data_stage_3__763_, data_stage_3__762_, data_stage_3__761_, data_stage_3__760_, data_stage_3__759_, data_stage_3__758_, data_stage_3__757_, data_stage_3__756_, data_stage_3__755_, data_stage_3__754_, data_stage_3__753_, data_stage_3__752_, data_stage_3__751_, data_stage_3__750_, data_stage_3__749_, data_stage_3__748_, data_stage_3__747_, data_stage_3__746_, data_stage_3__745_, data_stage_3__744_, data_stage_3__743_, data_stage_3__742_, data_stage_3__741_, data_stage_3__740_, data_stage_3__739_, data_stage_3__738_, data_stage_3__737_, data_stage_3__736_, data_stage_3__735_, data_stage_3__734_, data_stage_3__733_, data_stage_3__732_, data_stage_3__731_, data_stage_3__730_, data_stage_3__729_, data_stage_3__728_, data_stage_3__727_, data_stage_3__726_, data_stage_3__725_, data_stage_3__724_, data_stage_3__723_, data_stage_3__722_, data_stage_3__721_, data_stage_3__720_, data_stage_3__719_, data_stage_3__718_, data_stage_3__717_, data_stage_3__716_, data_stage_3__715_, data_stage_3__714_, data_stage_3__713_, data_stage_3__712_, data_stage_3__711_, data_stage_3__710_, data_stage_3__709_, data_stage_3__708_, data_stage_3__707_, data_stage_3__706_, data_stage_3__705_, data_stage_3__704_, data_stage_3__703_, data_stage_3__702_, data_stage_3__701_, data_stage_3__700_, data_stage_3__699_, data_stage_3__698_, data_stage_3__697_, data_stage_3__696_, data_stage_3__695_, data_stage_3__694_, data_stage_3__693_, data_stage_3__692_, data_stage_3__691_, data_stage_3__690_, data_stage_3__689_, data_stage_3__688_, data_stage_3__687_, data_stage_3__686_, data_stage_3__685_, data_stage_3__684_, data_stage_3__683_, data_stage_3__682_, data_stage_3__681_, data_stage_3__680_, data_stage_3__679_, data_stage_3__678_, data_stage_3__677_, data_stage_3__676_, data_stage_3__675_, data_stage_3__674_, data_stage_3__673_, data_stage_3__672_, data_stage_3__671_, data_stage_3__670_, data_stage_3__669_, data_stage_3__668_, data_stage_3__667_, data_stage_3__666_, data_stage_3__665_, data_stage_3__664_, data_stage_3__663_, data_stage_3__662_, data_stage_3__661_, data_stage_3__660_, data_stage_3__659_, data_stage_3__658_, data_stage_3__657_, data_stage_3__656_, data_stage_3__655_, data_stage_3__654_, data_stage_3__653_, data_stage_3__652_, data_stage_3__651_, data_stage_3__650_, data_stage_3__649_, data_stage_3__648_, data_stage_3__647_, data_stage_3__646_, data_stage_3__645_, data_stage_3__644_, data_stage_3__643_, data_stage_3__642_, data_stage_3__641_, data_stage_3__640_, data_stage_3__639_, data_stage_3__638_, data_stage_3__637_, data_stage_3__636_, data_stage_3__635_, data_stage_3__634_, data_stage_3__633_, data_stage_3__632_, data_stage_3__631_, data_stage_3__630_, data_stage_3__629_, data_stage_3__628_, data_stage_3__627_, data_stage_3__626_, data_stage_3__625_, data_stage_3__624_, data_stage_3__623_, data_stage_3__622_, data_stage_3__621_, data_stage_3__620_, data_stage_3__619_, data_stage_3__618_, data_stage_3__617_, data_stage_3__616_, data_stage_3__615_, data_stage_3__614_, data_stage_3__613_, data_stage_3__612_, data_stage_3__611_, data_stage_3__610_, data_stage_3__609_, data_stage_3__608_, data_stage_3__607_, data_stage_3__606_, data_stage_3__605_, data_stage_3__604_, data_stage_3__603_, data_stage_3__602_, data_stage_3__601_, data_stage_3__600_, data_stage_3__599_, data_stage_3__598_, data_stage_3__597_, data_stage_3__596_, data_stage_3__595_, data_stage_3__594_, data_stage_3__593_, data_stage_3__592_, data_stage_3__591_, data_stage_3__590_, data_stage_3__589_, data_stage_3__588_, data_stage_3__587_, data_stage_3__586_, data_stage_3__585_, data_stage_3__584_, data_stage_3__583_, data_stage_3__582_, data_stage_3__581_, data_stage_3__580_, data_stage_3__579_, data_stage_3__578_, data_stage_3__577_, data_stage_3__576_, data_stage_3__575_, data_stage_3__574_, data_stage_3__573_, data_stage_3__572_, data_stage_3__571_, data_stage_3__570_, data_stage_3__569_, data_stage_3__568_, data_stage_3__567_, data_stage_3__566_, data_stage_3__565_, data_stage_3__564_, data_stage_3__563_, data_stage_3__562_, data_stage_3__561_, data_stage_3__560_, data_stage_3__559_, data_stage_3__558_, data_stage_3__557_, data_stage_3__556_, data_stage_3__555_, data_stage_3__554_, data_stage_3__553_, data_stage_3__552_, data_stage_3__551_, data_stage_3__550_, data_stage_3__549_, data_stage_3__548_, data_stage_3__547_, data_stage_3__546_, data_stage_3__545_, data_stage_3__544_, data_stage_3__543_, data_stage_3__542_, data_stage_3__541_, data_stage_3__540_, data_stage_3__539_, data_stage_3__538_, data_stage_3__537_, data_stage_3__536_, data_stage_3__535_, data_stage_3__534_, data_stage_3__533_, data_stage_3__532_, data_stage_3__531_, data_stage_3__530_, data_stage_3__529_, data_stage_3__528_, data_stage_3__527_, data_stage_3__526_, data_stage_3__525_, data_stage_3__524_, data_stage_3__523_, data_stage_3__522_, data_stage_3__521_, data_stage_3__520_, data_stage_3__519_, data_stage_3__518_, data_stage_3__517_, data_stage_3__516_, data_stage_3__515_, data_stage_3__514_, data_stage_3__513_, data_stage_3__512_ }),
    .swap_i(sel_i[3]),
    .data_o({ data_stage_4__1023_, data_stage_4__1022_, data_stage_4__1021_, data_stage_4__1020_, data_stage_4__1019_, data_stage_4__1018_, data_stage_4__1017_, data_stage_4__1016_, data_stage_4__1015_, data_stage_4__1014_, data_stage_4__1013_, data_stage_4__1012_, data_stage_4__1011_, data_stage_4__1010_, data_stage_4__1009_, data_stage_4__1008_, data_stage_4__1007_, data_stage_4__1006_, data_stage_4__1005_, data_stage_4__1004_, data_stage_4__1003_, data_stage_4__1002_, data_stage_4__1001_, data_stage_4__1000_, data_stage_4__999_, data_stage_4__998_, data_stage_4__997_, data_stage_4__996_, data_stage_4__995_, data_stage_4__994_, data_stage_4__993_, data_stage_4__992_, data_stage_4__991_, data_stage_4__990_, data_stage_4__989_, data_stage_4__988_, data_stage_4__987_, data_stage_4__986_, data_stage_4__985_, data_stage_4__984_, data_stage_4__983_, data_stage_4__982_, data_stage_4__981_, data_stage_4__980_, data_stage_4__979_, data_stage_4__978_, data_stage_4__977_, data_stage_4__976_, data_stage_4__975_, data_stage_4__974_, data_stage_4__973_, data_stage_4__972_, data_stage_4__971_, data_stage_4__970_, data_stage_4__969_, data_stage_4__968_, data_stage_4__967_, data_stage_4__966_, data_stage_4__965_, data_stage_4__964_, data_stage_4__963_, data_stage_4__962_, data_stage_4__961_, data_stage_4__960_, data_stage_4__959_, data_stage_4__958_, data_stage_4__957_, data_stage_4__956_, data_stage_4__955_, data_stage_4__954_, data_stage_4__953_, data_stage_4__952_, data_stage_4__951_, data_stage_4__950_, data_stage_4__949_, data_stage_4__948_, data_stage_4__947_, data_stage_4__946_, data_stage_4__945_, data_stage_4__944_, data_stage_4__943_, data_stage_4__942_, data_stage_4__941_, data_stage_4__940_, data_stage_4__939_, data_stage_4__938_, data_stage_4__937_, data_stage_4__936_, data_stage_4__935_, data_stage_4__934_, data_stage_4__933_, data_stage_4__932_, data_stage_4__931_, data_stage_4__930_, data_stage_4__929_, data_stage_4__928_, data_stage_4__927_, data_stage_4__926_, data_stage_4__925_, data_stage_4__924_, data_stage_4__923_, data_stage_4__922_, data_stage_4__921_, data_stage_4__920_, data_stage_4__919_, data_stage_4__918_, data_stage_4__917_, data_stage_4__916_, data_stage_4__915_, data_stage_4__914_, data_stage_4__913_, data_stage_4__912_, data_stage_4__911_, data_stage_4__910_, data_stage_4__909_, data_stage_4__908_, data_stage_4__907_, data_stage_4__906_, data_stage_4__905_, data_stage_4__904_, data_stage_4__903_, data_stage_4__902_, data_stage_4__901_, data_stage_4__900_, data_stage_4__899_, data_stage_4__898_, data_stage_4__897_, data_stage_4__896_, data_stage_4__895_, data_stage_4__894_, data_stage_4__893_, data_stage_4__892_, data_stage_4__891_, data_stage_4__890_, data_stage_4__889_, data_stage_4__888_, data_stage_4__887_, data_stage_4__886_, data_stage_4__885_, data_stage_4__884_, data_stage_4__883_, data_stage_4__882_, data_stage_4__881_, data_stage_4__880_, data_stage_4__879_, data_stage_4__878_, data_stage_4__877_, data_stage_4__876_, data_stage_4__875_, data_stage_4__874_, data_stage_4__873_, data_stage_4__872_, data_stage_4__871_, data_stage_4__870_, data_stage_4__869_, data_stage_4__868_, data_stage_4__867_, data_stage_4__866_, data_stage_4__865_, data_stage_4__864_, data_stage_4__863_, data_stage_4__862_, data_stage_4__861_, data_stage_4__860_, data_stage_4__859_, data_stage_4__858_, data_stage_4__857_, data_stage_4__856_, data_stage_4__855_, data_stage_4__854_, data_stage_4__853_, data_stage_4__852_, data_stage_4__851_, data_stage_4__850_, data_stage_4__849_, data_stage_4__848_, data_stage_4__847_, data_stage_4__846_, data_stage_4__845_, data_stage_4__844_, data_stage_4__843_, data_stage_4__842_, data_stage_4__841_, data_stage_4__840_, data_stage_4__839_, data_stage_4__838_, data_stage_4__837_, data_stage_4__836_, data_stage_4__835_, data_stage_4__834_, data_stage_4__833_, data_stage_4__832_, data_stage_4__831_, data_stage_4__830_, data_stage_4__829_, data_stage_4__828_, data_stage_4__827_, data_stage_4__826_, data_stage_4__825_, data_stage_4__824_, data_stage_4__823_, data_stage_4__822_, data_stage_4__821_, data_stage_4__820_, data_stage_4__819_, data_stage_4__818_, data_stage_4__817_, data_stage_4__816_, data_stage_4__815_, data_stage_4__814_, data_stage_4__813_, data_stage_4__812_, data_stage_4__811_, data_stage_4__810_, data_stage_4__809_, data_stage_4__808_, data_stage_4__807_, data_stage_4__806_, data_stage_4__805_, data_stage_4__804_, data_stage_4__803_, data_stage_4__802_, data_stage_4__801_, data_stage_4__800_, data_stage_4__799_, data_stage_4__798_, data_stage_4__797_, data_stage_4__796_, data_stage_4__795_, data_stage_4__794_, data_stage_4__793_, data_stage_4__792_, data_stage_4__791_, data_stage_4__790_, data_stage_4__789_, data_stage_4__788_, data_stage_4__787_, data_stage_4__786_, data_stage_4__785_, data_stage_4__784_, data_stage_4__783_, data_stage_4__782_, data_stage_4__781_, data_stage_4__780_, data_stage_4__779_, data_stage_4__778_, data_stage_4__777_, data_stage_4__776_, data_stage_4__775_, data_stage_4__774_, data_stage_4__773_, data_stage_4__772_, data_stage_4__771_, data_stage_4__770_, data_stage_4__769_, data_stage_4__768_, data_stage_4__767_, data_stage_4__766_, data_stage_4__765_, data_stage_4__764_, data_stage_4__763_, data_stage_4__762_, data_stage_4__761_, data_stage_4__760_, data_stage_4__759_, data_stage_4__758_, data_stage_4__757_, data_stage_4__756_, data_stage_4__755_, data_stage_4__754_, data_stage_4__753_, data_stage_4__752_, data_stage_4__751_, data_stage_4__750_, data_stage_4__749_, data_stage_4__748_, data_stage_4__747_, data_stage_4__746_, data_stage_4__745_, data_stage_4__744_, data_stage_4__743_, data_stage_4__742_, data_stage_4__741_, data_stage_4__740_, data_stage_4__739_, data_stage_4__738_, data_stage_4__737_, data_stage_4__736_, data_stage_4__735_, data_stage_4__734_, data_stage_4__733_, data_stage_4__732_, data_stage_4__731_, data_stage_4__730_, data_stage_4__729_, data_stage_4__728_, data_stage_4__727_, data_stage_4__726_, data_stage_4__725_, data_stage_4__724_, data_stage_4__723_, data_stage_4__722_, data_stage_4__721_, data_stage_4__720_, data_stage_4__719_, data_stage_4__718_, data_stage_4__717_, data_stage_4__716_, data_stage_4__715_, data_stage_4__714_, data_stage_4__713_, data_stage_4__712_, data_stage_4__711_, data_stage_4__710_, data_stage_4__709_, data_stage_4__708_, data_stage_4__707_, data_stage_4__706_, data_stage_4__705_, data_stage_4__704_, data_stage_4__703_, data_stage_4__702_, data_stage_4__701_, data_stage_4__700_, data_stage_4__699_, data_stage_4__698_, data_stage_4__697_, data_stage_4__696_, data_stage_4__695_, data_stage_4__694_, data_stage_4__693_, data_stage_4__692_, data_stage_4__691_, data_stage_4__690_, data_stage_4__689_, data_stage_4__688_, data_stage_4__687_, data_stage_4__686_, data_stage_4__685_, data_stage_4__684_, data_stage_4__683_, data_stage_4__682_, data_stage_4__681_, data_stage_4__680_, data_stage_4__679_, data_stage_4__678_, data_stage_4__677_, data_stage_4__676_, data_stage_4__675_, data_stage_4__674_, data_stage_4__673_, data_stage_4__672_, data_stage_4__671_, data_stage_4__670_, data_stage_4__669_, data_stage_4__668_, data_stage_4__667_, data_stage_4__666_, data_stage_4__665_, data_stage_4__664_, data_stage_4__663_, data_stage_4__662_, data_stage_4__661_, data_stage_4__660_, data_stage_4__659_, data_stage_4__658_, data_stage_4__657_, data_stage_4__656_, data_stage_4__655_, data_stage_4__654_, data_stage_4__653_, data_stage_4__652_, data_stage_4__651_, data_stage_4__650_, data_stage_4__649_, data_stage_4__648_, data_stage_4__647_, data_stage_4__646_, data_stage_4__645_, data_stage_4__644_, data_stage_4__643_, data_stage_4__642_, data_stage_4__641_, data_stage_4__640_, data_stage_4__639_, data_stage_4__638_, data_stage_4__637_, data_stage_4__636_, data_stage_4__635_, data_stage_4__634_, data_stage_4__633_, data_stage_4__632_, data_stage_4__631_, data_stage_4__630_, data_stage_4__629_, data_stage_4__628_, data_stage_4__627_, data_stage_4__626_, data_stage_4__625_, data_stage_4__624_, data_stage_4__623_, data_stage_4__622_, data_stage_4__621_, data_stage_4__620_, data_stage_4__619_, data_stage_4__618_, data_stage_4__617_, data_stage_4__616_, data_stage_4__615_, data_stage_4__614_, data_stage_4__613_, data_stage_4__612_, data_stage_4__611_, data_stage_4__610_, data_stage_4__609_, data_stage_4__608_, data_stage_4__607_, data_stage_4__606_, data_stage_4__605_, data_stage_4__604_, data_stage_4__603_, data_stage_4__602_, data_stage_4__601_, data_stage_4__600_, data_stage_4__599_, data_stage_4__598_, data_stage_4__597_, data_stage_4__596_, data_stage_4__595_, data_stage_4__594_, data_stage_4__593_, data_stage_4__592_, data_stage_4__591_, data_stage_4__590_, data_stage_4__589_, data_stage_4__588_, data_stage_4__587_, data_stage_4__586_, data_stage_4__585_, data_stage_4__584_, data_stage_4__583_, data_stage_4__582_, data_stage_4__581_, data_stage_4__580_, data_stage_4__579_, data_stage_4__578_, data_stage_4__577_, data_stage_4__576_, data_stage_4__575_, data_stage_4__574_, data_stage_4__573_, data_stage_4__572_, data_stage_4__571_, data_stage_4__570_, data_stage_4__569_, data_stage_4__568_, data_stage_4__567_, data_stage_4__566_, data_stage_4__565_, data_stage_4__564_, data_stage_4__563_, data_stage_4__562_, data_stage_4__561_, data_stage_4__560_, data_stage_4__559_, data_stage_4__558_, data_stage_4__557_, data_stage_4__556_, data_stage_4__555_, data_stage_4__554_, data_stage_4__553_, data_stage_4__552_, data_stage_4__551_, data_stage_4__550_, data_stage_4__549_, data_stage_4__548_, data_stage_4__547_, data_stage_4__546_, data_stage_4__545_, data_stage_4__544_, data_stage_4__543_, data_stage_4__542_, data_stage_4__541_, data_stage_4__540_, data_stage_4__539_, data_stage_4__538_, data_stage_4__537_, data_stage_4__536_, data_stage_4__535_, data_stage_4__534_, data_stage_4__533_, data_stage_4__532_, data_stage_4__531_, data_stage_4__530_, data_stage_4__529_, data_stage_4__528_, data_stage_4__527_, data_stage_4__526_, data_stage_4__525_, data_stage_4__524_, data_stage_4__523_, data_stage_4__522_, data_stage_4__521_, data_stage_4__520_, data_stage_4__519_, data_stage_4__518_, data_stage_4__517_, data_stage_4__516_, data_stage_4__515_, data_stage_4__514_, data_stage_4__513_, data_stage_4__512_ })
  );


  bsg_swap_width_p512
  mux_stage_4__mux_swap_0__swap_inst
  (
    .data_i({ data_stage_4__1023_, data_stage_4__1022_, data_stage_4__1021_, data_stage_4__1020_, data_stage_4__1019_, data_stage_4__1018_, data_stage_4__1017_, data_stage_4__1016_, data_stage_4__1015_, data_stage_4__1014_, data_stage_4__1013_, data_stage_4__1012_, data_stage_4__1011_, data_stage_4__1010_, data_stage_4__1009_, data_stage_4__1008_, data_stage_4__1007_, data_stage_4__1006_, data_stage_4__1005_, data_stage_4__1004_, data_stage_4__1003_, data_stage_4__1002_, data_stage_4__1001_, data_stage_4__1000_, data_stage_4__999_, data_stage_4__998_, data_stage_4__997_, data_stage_4__996_, data_stage_4__995_, data_stage_4__994_, data_stage_4__993_, data_stage_4__992_, data_stage_4__991_, data_stage_4__990_, data_stage_4__989_, data_stage_4__988_, data_stage_4__987_, data_stage_4__986_, data_stage_4__985_, data_stage_4__984_, data_stage_4__983_, data_stage_4__982_, data_stage_4__981_, data_stage_4__980_, data_stage_4__979_, data_stage_4__978_, data_stage_4__977_, data_stage_4__976_, data_stage_4__975_, data_stage_4__974_, data_stage_4__973_, data_stage_4__972_, data_stage_4__971_, data_stage_4__970_, data_stage_4__969_, data_stage_4__968_, data_stage_4__967_, data_stage_4__966_, data_stage_4__965_, data_stage_4__964_, data_stage_4__963_, data_stage_4__962_, data_stage_4__961_, data_stage_4__960_, data_stage_4__959_, data_stage_4__958_, data_stage_4__957_, data_stage_4__956_, data_stage_4__955_, data_stage_4__954_, data_stage_4__953_, data_stage_4__952_, data_stage_4__951_, data_stage_4__950_, data_stage_4__949_, data_stage_4__948_, data_stage_4__947_, data_stage_4__946_, data_stage_4__945_, data_stage_4__944_, data_stage_4__943_, data_stage_4__942_, data_stage_4__941_, data_stage_4__940_, data_stage_4__939_, data_stage_4__938_, data_stage_4__937_, data_stage_4__936_, data_stage_4__935_, data_stage_4__934_, data_stage_4__933_, data_stage_4__932_, data_stage_4__931_, data_stage_4__930_, data_stage_4__929_, data_stage_4__928_, data_stage_4__927_, data_stage_4__926_, data_stage_4__925_, data_stage_4__924_, data_stage_4__923_, data_stage_4__922_, data_stage_4__921_, data_stage_4__920_, data_stage_4__919_, data_stage_4__918_, data_stage_4__917_, data_stage_4__916_, data_stage_4__915_, data_stage_4__914_, data_stage_4__913_, data_stage_4__912_, data_stage_4__911_, data_stage_4__910_, data_stage_4__909_, data_stage_4__908_, data_stage_4__907_, data_stage_4__906_, data_stage_4__905_, data_stage_4__904_, data_stage_4__903_, data_stage_4__902_, data_stage_4__901_, data_stage_4__900_, data_stage_4__899_, data_stage_4__898_, data_stage_4__897_, data_stage_4__896_, data_stage_4__895_, data_stage_4__894_, data_stage_4__893_, data_stage_4__892_, data_stage_4__891_, data_stage_4__890_, data_stage_4__889_, data_stage_4__888_, data_stage_4__887_, data_stage_4__886_, data_stage_4__885_, data_stage_4__884_, data_stage_4__883_, data_stage_4__882_, data_stage_4__881_, data_stage_4__880_, data_stage_4__879_, data_stage_4__878_, data_stage_4__877_, data_stage_4__876_, data_stage_4__875_, data_stage_4__874_, data_stage_4__873_, data_stage_4__872_, data_stage_4__871_, data_stage_4__870_, data_stage_4__869_, data_stage_4__868_, data_stage_4__867_, data_stage_4__866_, data_stage_4__865_, data_stage_4__864_, data_stage_4__863_, data_stage_4__862_, data_stage_4__861_, data_stage_4__860_, data_stage_4__859_, data_stage_4__858_, data_stage_4__857_, data_stage_4__856_, data_stage_4__855_, data_stage_4__854_, data_stage_4__853_, data_stage_4__852_, data_stage_4__851_, data_stage_4__850_, data_stage_4__849_, data_stage_4__848_, data_stage_4__847_, data_stage_4__846_, data_stage_4__845_, data_stage_4__844_, data_stage_4__843_, data_stage_4__842_, data_stage_4__841_, data_stage_4__840_, data_stage_4__839_, data_stage_4__838_, data_stage_4__837_, data_stage_4__836_, data_stage_4__835_, data_stage_4__834_, data_stage_4__833_, data_stage_4__832_, data_stage_4__831_, data_stage_4__830_, data_stage_4__829_, data_stage_4__828_, data_stage_4__827_, data_stage_4__826_, data_stage_4__825_, data_stage_4__824_, data_stage_4__823_, data_stage_4__822_, data_stage_4__821_, data_stage_4__820_, data_stage_4__819_, data_stage_4__818_, data_stage_4__817_, data_stage_4__816_, data_stage_4__815_, data_stage_4__814_, data_stage_4__813_, data_stage_4__812_, data_stage_4__811_, data_stage_4__810_, data_stage_4__809_, data_stage_4__808_, data_stage_4__807_, data_stage_4__806_, data_stage_4__805_, data_stage_4__804_, data_stage_4__803_, data_stage_4__802_, data_stage_4__801_, data_stage_4__800_, data_stage_4__799_, data_stage_4__798_, data_stage_4__797_, data_stage_4__796_, data_stage_4__795_, data_stage_4__794_, data_stage_4__793_, data_stage_4__792_, data_stage_4__791_, data_stage_4__790_, data_stage_4__789_, data_stage_4__788_, data_stage_4__787_, data_stage_4__786_, data_stage_4__785_, data_stage_4__784_, data_stage_4__783_, data_stage_4__782_, data_stage_4__781_, data_stage_4__780_, data_stage_4__779_, data_stage_4__778_, data_stage_4__777_, data_stage_4__776_, data_stage_4__775_, data_stage_4__774_, data_stage_4__773_, data_stage_4__772_, data_stage_4__771_, data_stage_4__770_, data_stage_4__769_, data_stage_4__768_, data_stage_4__767_, data_stage_4__766_, data_stage_4__765_, data_stage_4__764_, data_stage_4__763_, data_stage_4__762_, data_stage_4__761_, data_stage_4__760_, data_stage_4__759_, data_stage_4__758_, data_stage_4__757_, data_stage_4__756_, data_stage_4__755_, data_stage_4__754_, data_stage_4__753_, data_stage_4__752_, data_stage_4__751_, data_stage_4__750_, data_stage_4__749_, data_stage_4__748_, data_stage_4__747_, data_stage_4__746_, data_stage_4__745_, data_stage_4__744_, data_stage_4__743_, data_stage_4__742_, data_stage_4__741_, data_stage_4__740_, data_stage_4__739_, data_stage_4__738_, data_stage_4__737_, data_stage_4__736_, data_stage_4__735_, data_stage_4__734_, data_stage_4__733_, data_stage_4__732_, data_stage_4__731_, data_stage_4__730_, data_stage_4__729_, data_stage_4__728_, data_stage_4__727_, data_stage_4__726_, data_stage_4__725_, data_stage_4__724_, data_stage_4__723_, data_stage_4__722_, data_stage_4__721_, data_stage_4__720_, data_stage_4__719_, data_stage_4__718_, data_stage_4__717_, data_stage_4__716_, data_stage_4__715_, data_stage_4__714_, data_stage_4__713_, data_stage_4__712_, data_stage_4__711_, data_stage_4__710_, data_stage_4__709_, data_stage_4__708_, data_stage_4__707_, data_stage_4__706_, data_stage_4__705_, data_stage_4__704_, data_stage_4__703_, data_stage_4__702_, data_stage_4__701_, data_stage_4__700_, data_stage_4__699_, data_stage_4__698_, data_stage_4__697_, data_stage_4__696_, data_stage_4__695_, data_stage_4__694_, data_stage_4__693_, data_stage_4__692_, data_stage_4__691_, data_stage_4__690_, data_stage_4__689_, data_stage_4__688_, data_stage_4__687_, data_stage_4__686_, data_stage_4__685_, data_stage_4__684_, data_stage_4__683_, data_stage_4__682_, data_stage_4__681_, data_stage_4__680_, data_stage_4__679_, data_stage_4__678_, data_stage_4__677_, data_stage_4__676_, data_stage_4__675_, data_stage_4__674_, data_stage_4__673_, data_stage_4__672_, data_stage_4__671_, data_stage_4__670_, data_stage_4__669_, data_stage_4__668_, data_stage_4__667_, data_stage_4__666_, data_stage_4__665_, data_stage_4__664_, data_stage_4__663_, data_stage_4__662_, data_stage_4__661_, data_stage_4__660_, data_stage_4__659_, data_stage_4__658_, data_stage_4__657_, data_stage_4__656_, data_stage_4__655_, data_stage_4__654_, data_stage_4__653_, data_stage_4__652_, data_stage_4__651_, data_stage_4__650_, data_stage_4__649_, data_stage_4__648_, data_stage_4__647_, data_stage_4__646_, data_stage_4__645_, data_stage_4__644_, data_stage_4__643_, data_stage_4__642_, data_stage_4__641_, data_stage_4__640_, data_stage_4__639_, data_stage_4__638_, data_stage_4__637_, data_stage_4__636_, data_stage_4__635_, data_stage_4__634_, data_stage_4__633_, data_stage_4__632_, data_stage_4__631_, data_stage_4__630_, data_stage_4__629_, data_stage_4__628_, data_stage_4__627_, data_stage_4__626_, data_stage_4__625_, data_stage_4__624_, data_stage_4__623_, data_stage_4__622_, data_stage_4__621_, data_stage_4__620_, data_stage_4__619_, data_stage_4__618_, data_stage_4__617_, data_stage_4__616_, data_stage_4__615_, data_stage_4__614_, data_stage_4__613_, data_stage_4__612_, data_stage_4__611_, data_stage_4__610_, data_stage_4__609_, data_stage_4__608_, data_stage_4__607_, data_stage_4__606_, data_stage_4__605_, data_stage_4__604_, data_stage_4__603_, data_stage_4__602_, data_stage_4__601_, data_stage_4__600_, data_stage_4__599_, data_stage_4__598_, data_stage_4__597_, data_stage_4__596_, data_stage_4__595_, data_stage_4__594_, data_stage_4__593_, data_stage_4__592_, data_stage_4__591_, data_stage_4__590_, data_stage_4__589_, data_stage_4__588_, data_stage_4__587_, data_stage_4__586_, data_stage_4__585_, data_stage_4__584_, data_stage_4__583_, data_stage_4__582_, data_stage_4__581_, data_stage_4__580_, data_stage_4__579_, data_stage_4__578_, data_stage_4__577_, data_stage_4__576_, data_stage_4__575_, data_stage_4__574_, data_stage_4__573_, data_stage_4__572_, data_stage_4__571_, data_stage_4__570_, data_stage_4__569_, data_stage_4__568_, data_stage_4__567_, data_stage_4__566_, data_stage_4__565_, data_stage_4__564_, data_stage_4__563_, data_stage_4__562_, data_stage_4__561_, data_stage_4__560_, data_stage_4__559_, data_stage_4__558_, data_stage_4__557_, data_stage_4__556_, data_stage_4__555_, data_stage_4__554_, data_stage_4__553_, data_stage_4__552_, data_stage_4__551_, data_stage_4__550_, data_stage_4__549_, data_stage_4__548_, data_stage_4__547_, data_stage_4__546_, data_stage_4__545_, data_stage_4__544_, data_stage_4__543_, data_stage_4__542_, data_stage_4__541_, data_stage_4__540_, data_stage_4__539_, data_stage_4__538_, data_stage_4__537_, data_stage_4__536_, data_stage_4__535_, data_stage_4__534_, data_stage_4__533_, data_stage_4__532_, data_stage_4__531_, data_stage_4__530_, data_stage_4__529_, data_stage_4__528_, data_stage_4__527_, data_stage_4__526_, data_stage_4__525_, data_stage_4__524_, data_stage_4__523_, data_stage_4__522_, data_stage_4__521_, data_stage_4__520_, data_stage_4__519_, data_stage_4__518_, data_stage_4__517_, data_stage_4__516_, data_stage_4__515_, data_stage_4__514_, data_stage_4__513_, data_stage_4__512_, data_stage_4__511_, data_stage_4__510_, data_stage_4__509_, data_stage_4__508_, data_stage_4__507_, data_stage_4__506_, data_stage_4__505_, data_stage_4__504_, data_stage_4__503_, data_stage_4__502_, data_stage_4__501_, data_stage_4__500_, data_stage_4__499_, data_stage_4__498_, data_stage_4__497_, data_stage_4__496_, data_stage_4__495_, data_stage_4__494_, data_stage_4__493_, data_stage_4__492_, data_stage_4__491_, data_stage_4__490_, data_stage_4__489_, data_stage_4__488_, data_stage_4__487_, data_stage_4__486_, data_stage_4__485_, data_stage_4__484_, data_stage_4__483_, data_stage_4__482_, data_stage_4__481_, data_stage_4__480_, data_stage_4__479_, data_stage_4__478_, data_stage_4__477_, data_stage_4__476_, data_stage_4__475_, data_stage_4__474_, data_stage_4__473_, data_stage_4__472_, data_stage_4__471_, data_stage_4__470_, data_stage_4__469_, data_stage_4__468_, data_stage_4__467_, data_stage_4__466_, data_stage_4__465_, data_stage_4__464_, data_stage_4__463_, data_stage_4__462_, data_stage_4__461_, data_stage_4__460_, data_stage_4__459_, data_stage_4__458_, data_stage_4__457_, data_stage_4__456_, data_stage_4__455_, data_stage_4__454_, data_stage_4__453_, data_stage_4__452_, data_stage_4__451_, data_stage_4__450_, data_stage_4__449_, data_stage_4__448_, data_stage_4__447_, data_stage_4__446_, data_stage_4__445_, data_stage_4__444_, data_stage_4__443_, data_stage_4__442_, data_stage_4__441_, data_stage_4__440_, data_stage_4__439_, data_stage_4__438_, data_stage_4__437_, data_stage_4__436_, data_stage_4__435_, data_stage_4__434_, data_stage_4__433_, data_stage_4__432_, data_stage_4__431_, data_stage_4__430_, data_stage_4__429_, data_stage_4__428_, data_stage_4__427_, data_stage_4__426_, data_stage_4__425_, data_stage_4__424_, data_stage_4__423_, data_stage_4__422_, data_stage_4__421_, data_stage_4__420_, data_stage_4__419_, data_stage_4__418_, data_stage_4__417_, data_stage_4__416_, data_stage_4__415_, data_stage_4__414_, data_stage_4__413_, data_stage_4__412_, data_stage_4__411_, data_stage_4__410_, data_stage_4__409_, data_stage_4__408_, data_stage_4__407_, data_stage_4__406_, data_stage_4__405_, data_stage_4__404_, data_stage_4__403_, data_stage_4__402_, data_stage_4__401_, data_stage_4__400_, data_stage_4__399_, data_stage_4__398_, data_stage_4__397_, data_stage_4__396_, data_stage_4__395_, data_stage_4__394_, data_stage_4__393_, data_stage_4__392_, data_stage_4__391_, data_stage_4__390_, data_stage_4__389_, data_stage_4__388_, data_stage_4__387_, data_stage_4__386_, data_stage_4__385_, data_stage_4__384_, data_stage_4__383_, data_stage_4__382_, data_stage_4__381_, data_stage_4__380_, data_stage_4__379_, data_stage_4__378_, data_stage_4__377_, data_stage_4__376_, data_stage_4__375_, data_stage_4__374_, data_stage_4__373_, data_stage_4__372_, data_stage_4__371_, data_stage_4__370_, data_stage_4__369_, data_stage_4__368_, data_stage_4__367_, data_stage_4__366_, data_stage_4__365_, data_stage_4__364_, data_stage_4__363_, data_stage_4__362_, data_stage_4__361_, data_stage_4__360_, data_stage_4__359_, data_stage_4__358_, data_stage_4__357_, data_stage_4__356_, data_stage_4__355_, data_stage_4__354_, data_stage_4__353_, data_stage_4__352_, data_stage_4__351_, data_stage_4__350_, data_stage_4__349_, data_stage_4__348_, data_stage_4__347_, data_stage_4__346_, data_stage_4__345_, data_stage_4__344_, data_stage_4__343_, data_stage_4__342_, data_stage_4__341_, data_stage_4__340_, data_stage_4__339_, data_stage_4__338_, data_stage_4__337_, data_stage_4__336_, data_stage_4__335_, data_stage_4__334_, data_stage_4__333_, data_stage_4__332_, data_stage_4__331_, data_stage_4__330_, data_stage_4__329_, data_stage_4__328_, data_stage_4__327_, data_stage_4__326_, data_stage_4__325_, data_stage_4__324_, data_stage_4__323_, data_stage_4__322_, data_stage_4__321_, data_stage_4__320_, data_stage_4__319_, data_stage_4__318_, data_stage_4__317_, data_stage_4__316_, data_stage_4__315_, data_stage_4__314_, data_stage_4__313_, data_stage_4__312_, data_stage_4__311_, data_stage_4__310_, data_stage_4__309_, data_stage_4__308_, data_stage_4__307_, data_stage_4__306_, data_stage_4__305_, data_stage_4__304_, data_stage_4__303_, data_stage_4__302_, data_stage_4__301_, data_stage_4__300_, data_stage_4__299_, data_stage_4__298_, data_stage_4__297_, data_stage_4__296_, data_stage_4__295_, data_stage_4__294_, data_stage_4__293_, data_stage_4__292_, data_stage_4__291_, data_stage_4__290_, data_stage_4__289_, data_stage_4__288_, data_stage_4__287_, data_stage_4__286_, data_stage_4__285_, data_stage_4__284_, data_stage_4__283_, data_stage_4__282_, data_stage_4__281_, data_stage_4__280_, data_stage_4__279_, data_stage_4__278_, data_stage_4__277_, data_stage_4__276_, data_stage_4__275_, data_stage_4__274_, data_stage_4__273_, data_stage_4__272_, data_stage_4__271_, data_stage_4__270_, data_stage_4__269_, data_stage_4__268_, data_stage_4__267_, data_stage_4__266_, data_stage_4__265_, data_stage_4__264_, data_stage_4__263_, data_stage_4__262_, data_stage_4__261_, data_stage_4__260_, data_stage_4__259_, data_stage_4__258_, data_stage_4__257_, data_stage_4__256_, data_stage_4__255_, data_stage_4__254_, data_stage_4__253_, data_stage_4__252_, data_stage_4__251_, data_stage_4__250_, data_stage_4__249_, data_stage_4__248_, data_stage_4__247_, data_stage_4__246_, data_stage_4__245_, data_stage_4__244_, data_stage_4__243_, data_stage_4__242_, data_stage_4__241_, data_stage_4__240_, data_stage_4__239_, data_stage_4__238_, data_stage_4__237_, data_stage_4__236_, data_stage_4__235_, data_stage_4__234_, data_stage_4__233_, data_stage_4__232_, data_stage_4__231_, data_stage_4__230_, data_stage_4__229_, data_stage_4__228_, data_stage_4__227_, data_stage_4__226_, data_stage_4__225_, data_stage_4__224_, data_stage_4__223_, data_stage_4__222_, data_stage_4__221_, data_stage_4__220_, data_stage_4__219_, data_stage_4__218_, data_stage_4__217_, data_stage_4__216_, data_stage_4__215_, data_stage_4__214_, data_stage_4__213_, data_stage_4__212_, data_stage_4__211_, data_stage_4__210_, data_stage_4__209_, data_stage_4__208_, data_stage_4__207_, data_stage_4__206_, data_stage_4__205_, data_stage_4__204_, data_stage_4__203_, data_stage_4__202_, data_stage_4__201_, data_stage_4__200_, data_stage_4__199_, data_stage_4__198_, data_stage_4__197_, data_stage_4__196_, data_stage_4__195_, data_stage_4__194_, data_stage_4__193_, data_stage_4__192_, data_stage_4__191_, data_stage_4__190_, data_stage_4__189_, data_stage_4__188_, data_stage_4__187_, data_stage_4__186_, data_stage_4__185_, data_stage_4__184_, data_stage_4__183_, data_stage_4__182_, data_stage_4__181_, data_stage_4__180_, data_stage_4__179_, data_stage_4__178_, data_stage_4__177_, data_stage_4__176_, data_stage_4__175_, data_stage_4__174_, data_stage_4__173_, data_stage_4__172_, data_stage_4__171_, data_stage_4__170_, data_stage_4__169_, data_stage_4__168_, data_stage_4__167_, data_stage_4__166_, data_stage_4__165_, data_stage_4__164_, data_stage_4__163_, data_stage_4__162_, data_stage_4__161_, data_stage_4__160_, data_stage_4__159_, data_stage_4__158_, data_stage_4__157_, data_stage_4__156_, data_stage_4__155_, data_stage_4__154_, data_stage_4__153_, data_stage_4__152_, data_stage_4__151_, data_stage_4__150_, data_stage_4__149_, data_stage_4__148_, data_stage_4__147_, data_stage_4__146_, data_stage_4__145_, data_stage_4__144_, data_stage_4__143_, data_stage_4__142_, data_stage_4__141_, data_stage_4__140_, data_stage_4__139_, data_stage_4__138_, data_stage_4__137_, data_stage_4__136_, data_stage_4__135_, data_stage_4__134_, data_stage_4__133_, data_stage_4__132_, data_stage_4__131_, data_stage_4__130_, data_stage_4__129_, data_stage_4__128_, data_stage_4__127_, data_stage_4__126_, data_stage_4__125_, data_stage_4__124_, data_stage_4__123_, data_stage_4__122_, data_stage_4__121_, data_stage_4__120_, data_stage_4__119_, data_stage_4__118_, data_stage_4__117_, data_stage_4__116_, data_stage_4__115_, data_stage_4__114_, data_stage_4__113_, data_stage_4__112_, data_stage_4__111_, data_stage_4__110_, data_stage_4__109_, data_stage_4__108_, data_stage_4__107_, data_stage_4__106_, data_stage_4__105_, data_stage_4__104_, data_stage_4__103_, data_stage_4__102_, data_stage_4__101_, data_stage_4__100_, data_stage_4__99_, data_stage_4__98_, data_stage_4__97_, data_stage_4__96_, data_stage_4__95_, data_stage_4__94_, data_stage_4__93_, data_stage_4__92_, data_stage_4__91_, data_stage_4__90_, data_stage_4__89_, data_stage_4__88_, data_stage_4__87_, data_stage_4__86_, data_stage_4__85_, data_stage_4__84_, data_stage_4__83_, data_stage_4__82_, data_stage_4__81_, data_stage_4__80_, data_stage_4__79_, data_stage_4__78_, data_stage_4__77_, data_stage_4__76_, data_stage_4__75_, data_stage_4__74_, data_stage_4__73_, data_stage_4__72_, data_stage_4__71_, data_stage_4__70_, data_stage_4__69_, data_stage_4__68_, data_stage_4__67_, data_stage_4__66_, data_stage_4__65_, data_stage_4__64_, data_stage_4__63_, data_stage_4__62_, data_stage_4__61_, data_stage_4__60_, data_stage_4__59_, data_stage_4__58_, data_stage_4__57_, data_stage_4__56_, data_stage_4__55_, data_stage_4__54_, data_stage_4__53_, data_stage_4__52_, data_stage_4__51_, data_stage_4__50_, data_stage_4__49_, data_stage_4__48_, data_stage_4__47_, data_stage_4__46_, data_stage_4__45_, data_stage_4__44_, data_stage_4__43_, data_stage_4__42_, data_stage_4__41_, data_stage_4__40_, data_stage_4__39_, data_stage_4__38_, data_stage_4__37_, data_stage_4__36_, data_stage_4__35_, data_stage_4__34_, data_stage_4__33_, data_stage_4__32_, data_stage_4__31_, data_stage_4__30_, data_stage_4__29_, data_stage_4__28_, data_stage_4__27_, data_stage_4__26_, data_stage_4__25_, data_stage_4__24_, data_stage_4__23_, data_stage_4__22_, data_stage_4__21_, data_stage_4__20_, data_stage_4__19_, data_stage_4__18_, data_stage_4__17_, data_stage_4__16_, data_stage_4__15_, data_stage_4__14_, data_stage_4__13_, data_stage_4__12_, data_stage_4__11_, data_stage_4__10_, data_stage_4__9_, data_stage_4__8_, data_stage_4__7_, data_stage_4__6_, data_stage_4__5_, data_stage_4__4_, data_stage_4__3_, data_stage_4__2_, data_stage_4__1_, data_stage_4__0_ }),
    .swap_i(sel_i[4]),
    .data_o(data_o)
  );


endmodule

